
module psi_BMR_b10000_n2 ( p_input, o );
  input [19999:0] p_input;
  output [9999:0] o;


  AND U1 ( .A(p_input[9]), .B(p_input[10009]), .Z(o[9]) );
  AND U2 ( .A(p_input[99]), .B(p_input[10099]), .Z(o[99]) );
  AND U3 ( .A(p_input[999]), .B(p_input[10999]), .Z(o[999]) );
  AND U4 ( .A(p_input[9999]), .B(p_input[19999]), .Z(o[9999]) );
  AND U5 ( .A(p_input[9998]), .B(p_input[19998]), .Z(o[9998]) );
  AND U6 ( .A(p_input[9997]), .B(p_input[19997]), .Z(o[9997]) );
  AND U7 ( .A(p_input[9996]), .B(p_input[19996]), .Z(o[9996]) );
  AND U8 ( .A(p_input[9995]), .B(p_input[19995]), .Z(o[9995]) );
  AND U9 ( .A(p_input[9994]), .B(p_input[19994]), .Z(o[9994]) );
  AND U10 ( .A(p_input[9993]), .B(p_input[19993]), .Z(o[9993]) );
  AND U11 ( .A(p_input[9992]), .B(p_input[19992]), .Z(o[9992]) );
  AND U12 ( .A(p_input[9991]), .B(p_input[19991]), .Z(o[9991]) );
  AND U13 ( .A(p_input[9990]), .B(p_input[19990]), .Z(o[9990]) );
  AND U14 ( .A(p_input[998]), .B(p_input[10998]), .Z(o[998]) );
  AND U15 ( .A(p_input[9989]), .B(p_input[19989]), .Z(o[9989]) );
  AND U16 ( .A(p_input[9988]), .B(p_input[19988]), .Z(o[9988]) );
  AND U17 ( .A(p_input[9987]), .B(p_input[19987]), .Z(o[9987]) );
  AND U18 ( .A(p_input[9986]), .B(p_input[19986]), .Z(o[9986]) );
  AND U19 ( .A(p_input[9985]), .B(p_input[19985]), .Z(o[9985]) );
  AND U20 ( .A(p_input[9984]), .B(p_input[19984]), .Z(o[9984]) );
  AND U21 ( .A(p_input[9983]), .B(p_input[19983]), .Z(o[9983]) );
  AND U22 ( .A(p_input[9982]), .B(p_input[19982]), .Z(o[9982]) );
  AND U23 ( .A(p_input[9981]), .B(p_input[19981]), .Z(o[9981]) );
  AND U24 ( .A(p_input[9980]), .B(p_input[19980]), .Z(o[9980]) );
  AND U25 ( .A(p_input[997]), .B(p_input[10997]), .Z(o[997]) );
  AND U26 ( .A(p_input[9979]), .B(p_input[19979]), .Z(o[9979]) );
  AND U27 ( .A(p_input[9978]), .B(p_input[19978]), .Z(o[9978]) );
  AND U28 ( .A(p_input[9977]), .B(p_input[19977]), .Z(o[9977]) );
  AND U29 ( .A(p_input[9976]), .B(p_input[19976]), .Z(o[9976]) );
  AND U30 ( .A(p_input[9975]), .B(p_input[19975]), .Z(o[9975]) );
  AND U31 ( .A(p_input[9974]), .B(p_input[19974]), .Z(o[9974]) );
  AND U32 ( .A(p_input[9973]), .B(p_input[19973]), .Z(o[9973]) );
  AND U33 ( .A(p_input[9972]), .B(p_input[19972]), .Z(o[9972]) );
  AND U34 ( .A(p_input[9971]), .B(p_input[19971]), .Z(o[9971]) );
  AND U35 ( .A(p_input[9970]), .B(p_input[19970]), .Z(o[9970]) );
  AND U36 ( .A(p_input[996]), .B(p_input[10996]), .Z(o[996]) );
  AND U37 ( .A(p_input[9969]), .B(p_input[19969]), .Z(o[9969]) );
  AND U38 ( .A(p_input[9968]), .B(p_input[19968]), .Z(o[9968]) );
  AND U39 ( .A(p_input[9967]), .B(p_input[19967]), .Z(o[9967]) );
  AND U40 ( .A(p_input[9966]), .B(p_input[19966]), .Z(o[9966]) );
  AND U41 ( .A(p_input[9965]), .B(p_input[19965]), .Z(o[9965]) );
  AND U42 ( .A(p_input[9964]), .B(p_input[19964]), .Z(o[9964]) );
  AND U43 ( .A(p_input[9963]), .B(p_input[19963]), .Z(o[9963]) );
  AND U44 ( .A(p_input[9962]), .B(p_input[19962]), .Z(o[9962]) );
  AND U45 ( .A(p_input[9961]), .B(p_input[19961]), .Z(o[9961]) );
  AND U46 ( .A(p_input[9960]), .B(p_input[19960]), .Z(o[9960]) );
  AND U47 ( .A(p_input[995]), .B(p_input[10995]), .Z(o[995]) );
  AND U48 ( .A(p_input[9959]), .B(p_input[19959]), .Z(o[9959]) );
  AND U49 ( .A(p_input[9958]), .B(p_input[19958]), .Z(o[9958]) );
  AND U50 ( .A(p_input[9957]), .B(p_input[19957]), .Z(o[9957]) );
  AND U51 ( .A(p_input[9956]), .B(p_input[19956]), .Z(o[9956]) );
  AND U52 ( .A(p_input[9955]), .B(p_input[19955]), .Z(o[9955]) );
  AND U53 ( .A(p_input[9954]), .B(p_input[19954]), .Z(o[9954]) );
  AND U54 ( .A(p_input[9953]), .B(p_input[19953]), .Z(o[9953]) );
  AND U55 ( .A(p_input[9952]), .B(p_input[19952]), .Z(o[9952]) );
  AND U56 ( .A(p_input[9951]), .B(p_input[19951]), .Z(o[9951]) );
  AND U57 ( .A(p_input[9950]), .B(p_input[19950]), .Z(o[9950]) );
  AND U58 ( .A(p_input[994]), .B(p_input[10994]), .Z(o[994]) );
  AND U59 ( .A(p_input[9949]), .B(p_input[19949]), .Z(o[9949]) );
  AND U60 ( .A(p_input[9948]), .B(p_input[19948]), .Z(o[9948]) );
  AND U61 ( .A(p_input[9947]), .B(p_input[19947]), .Z(o[9947]) );
  AND U62 ( .A(p_input[9946]), .B(p_input[19946]), .Z(o[9946]) );
  AND U63 ( .A(p_input[9945]), .B(p_input[19945]), .Z(o[9945]) );
  AND U64 ( .A(p_input[9944]), .B(p_input[19944]), .Z(o[9944]) );
  AND U65 ( .A(p_input[9943]), .B(p_input[19943]), .Z(o[9943]) );
  AND U66 ( .A(p_input[9942]), .B(p_input[19942]), .Z(o[9942]) );
  AND U67 ( .A(p_input[9941]), .B(p_input[19941]), .Z(o[9941]) );
  AND U68 ( .A(p_input[9940]), .B(p_input[19940]), .Z(o[9940]) );
  AND U69 ( .A(p_input[993]), .B(p_input[10993]), .Z(o[993]) );
  AND U70 ( .A(p_input[9939]), .B(p_input[19939]), .Z(o[9939]) );
  AND U71 ( .A(p_input[9938]), .B(p_input[19938]), .Z(o[9938]) );
  AND U72 ( .A(p_input[9937]), .B(p_input[19937]), .Z(o[9937]) );
  AND U73 ( .A(p_input[9936]), .B(p_input[19936]), .Z(o[9936]) );
  AND U74 ( .A(p_input[9935]), .B(p_input[19935]), .Z(o[9935]) );
  AND U75 ( .A(p_input[9934]), .B(p_input[19934]), .Z(o[9934]) );
  AND U76 ( .A(p_input[9933]), .B(p_input[19933]), .Z(o[9933]) );
  AND U77 ( .A(p_input[9932]), .B(p_input[19932]), .Z(o[9932]) );
  AND U78 ( .A(p_input[9931]), .B(p_input[19931]), .Z(o[9931]) );
  AND U79 ( .A(p_input[9930]), .B(p_input[19930]), .Z(o[9930]) );
  AND U80 ( .A(p_input[992]), .B(p_input[10992]), .Z(o[992]) );
  AND U81 ( .A(p_input[9929]), .B(p_input[19929]), .Z(o[9929]) );
  AND U82 ( .A(p_input[9928]), .B(p_input[19928]), .Z(o[9928]) );
  AND U83 ( .A(p_input[9927]), .B(p_input[19927]), .Z(o[9927]) );
  AND U84 ( .A(p_input[9926]), .B(p_input[19926]), .Z(o[9926]) );
  AND U85 ( .A(p_input[9925]), .B(p_input[19925]), .Z(o[9925]) );
  AND U86 ( .A(p_input[9924]), .B(p_input[19924]), .Z(o[9924]) );
  AND U87 ( .A(p_input[9923]), .B(p_input[19923]), .Z(o[9923]) );
  AND U88 ( .A(p_input[9922]), .B(p_input[19922]), .Z(o[9922]) );
  AND U89 ( .A(p_input[9921]), .B(p_input[19921]), .Z(o[9921]) );
  AND U90 ( .A(p_input[9920]), .B(p_input[19920]), .Z(o[9920]) );
  AND U91 ( .A(p_input[991]), .B(p_input[10991]), .Z(o[991]) );
  AND U92 ( .A(p_input[9919]), .B(p_input[19919]), .Z(o[9919]) );
  AND U93 ( .A(p_input[9918]), .B(p_input[19918]), .Z(o[9918]) );
  AND U94 ( .A(p_input[9917]), .B(p_input[19917]), .Z(o[9917]) );
  AND U95 ( .A(p_input[9916]), .B(p_input[19916]), .Z(o[9916]) );
  AND U96 ( .A(p_input[9915]), .B(p_input[19915]), .Z(o[9915]) );
  AND U97 ( .A(p_input[9914]), .B(p_input[19914]), .Z(o[9914]) );
  AND U98 ( .A(p_input[9913]), .B(p_input[19913]), .Z(o[9913]) );
  AND U99 ( .A(p_input[9912]), .B(p_input[19912]), .Z(o[9912]) );
  AND U100 ( .A(p_input[9911]), .B(p_input[19911]), .Z(o[9911]) );
  AND U101 ( .A(p_input[9910]), .B(p_input[19910]), .Z(o[9910]) );
  AND U102 ( .A(p_input[990]), .B(p_input[10990]), .Z(o[990]) );
  AND U103 ( .A(p_input[9909]), .B(p_input[19909]), .Z(o[9909]) );
  AND U104 ( .A(p_input[9908]), .B(p_input[19908]), .Z(o[9908]) );
  AND U105 ( .A(p_input[9907]), .B(p_input[19907]), .Z(o[9907]) );
  AND U106 ( .A(p_input[9906]), .B(p_input[19906]), .Z(o[9906]) );
  AND U107 ( .A(p_input[9905]), .B(p_input[19905]), .Z(o[9905]) );
  AND U108 ( .A(p_input[9904]), .B(p_input[19904]), .Z(o[9904]) );
  AND U109 ( .A(p_input[9903]), .B(p_input[19903]), .Z(o[9903]) );
  AND U110 ( .A(p_input[9902]), .B(p_input[19902]), .Z(o[9902]) );
  AND U111 ( .A(p_input[9901]), .B(p_input[19901]), .Z(o[9901]) );
  AND U112 ( .A(p_input[9900]), .B(p_input[19900]), .Z(o[9900]) );
  AND U113 ( .A(p_input[98]), .B(p_input[10098]), .Z(o[98]) );
  AND U114 ( .A(p_input[989]), .B(p_input[10989]), .Z(o[989]) );
  AND U115 ( .A(p_input[9899]), .B(p_input[19899]), .Z(o[9899]) );
  AND U116 ( .A(p_input[9898]), .B(p_input[19898]), .Z(o[9898]) );
  AND U117 ( .A(p_input[9897]), .B(p_input[19897]), .Z(o[9897]) );
  AND U118 ( .A(p_input[9896]), .B(p_input[19896]), .Z(o[9896]) );
  AND U119 ( .A(p_input[9895]), .B(p_input[19895]), .Z(o[9895]) );
  AND U120 ( .A(p_input[9894]), .B(p_input[19894]), .Z(o[9894]) );
  AND U121 ( .A(p_input[9893]), .B(p_input[19893]), .Z(o[9893]) );
  AND U122 ( .A(p_input[9892]), .B(p_input[19892]), .Z(o[9892]) );
  AND U123 ( .A(p_input[9891]), .B(p_input[19891]), .Z(o[9891]) );
  AND U124 ( .A(p_input[9890]), .B(p_input[19890]), .Z(o[9890]) );
  AND U125 ( .A(p_input[988]), .B(p_input[10988]), .Z(o[988]) );
  AND U126 ( .A(p_input[9889]), .B(p_input[19889]), .Z(o[9889]) );
  AND U127 ( .A(p_input[9888]), .B(p_input[19888]), .Z(o[9888]) );
  AND U128 ( .A(p_input[9887]), .B(p_input[19887]), .Z(o[9887]) );
  AND U129 ( .A(p_input[9886]), .B(p_input[19886]), .Z(o[9886]) );
  AND U130 ( .A(p_input[9885]), .B(p_input[19885]), .Z(o[9885]) );
  AND U131 ( .A(p_input[9884]), .B(p_input[19884]), .Z(o[9884]) );
  AND U132 ( .A(p_input[9883]), .B(p_input[19883]), .Z(o[9883]) );
  AND U133 ( .A(p_input[9882]), .B(p_input[19882]), .Z(o[9882]) );
  AND U134 ( .A(p_input[9881]), .B(p_input[19881]), .Z(o[9881]) );
  AND U135 ( .A(p_input[9880]), .B(p_input[19880]), .Z(o[9880]) );
  AND U136 ( .A(p_input[987]), .B(p_input[10987]), .Z(o[987]) );
  AND U137 ( .A(p_input[9879]), .B(p_input[19879]), .Z(o[9879]) );
  AND U138 ( .A(p_input[9878]), .B(p_input[19878]), .Z(o[9878]) );
  AND U139 ( .A(p_input[9877]), .B(p_input[19877]), .Z(o[9877]) );
  AND U140 ( .A(p_input[9876]), .B(p_input[19876]), .Z(o[9876]) );
  AND U141 ( .A(p_input[9875]), .B(p_input[19875]), .Z(o[9875]) );
  AND U142 ( .A(p_input[9874]), .B(p_input[19874]), .Z(o[9874]) );
  AND U143 ( .A(p_input[9873]), .B(p_input[19873]), .Z(o[9873]) );
  AND U144 ( .A(p_input[9872]), .B(p_input[19872]), .Z(o[9872]) );
  AND U145 ( .A(p_input[9871]), .B(p_input[19871]), .Z(o[9871]) );
  AND U146 ( .A(p_input[9870]), .B(p_input[19870]), .Z(o[9870]) );
  AND U147 ( .A(p_input[986]), .B(p_input[10986]), .Z(o[986]) );
  AND U148 ( .A(p_input[9869]), .B(p_input[19869]), .Z(o[9869]) );
  AND U149 ( .A(p_input[9868]), .B(p_input[19868]), .Z(o[9868]) );
  AND U150 ( .A(p_input[9867]), .B(p_input[19867]), .Z(o[9867]) );
  AND U151 ( .A(p_input[9866]), .B(p_input[19866]), .Z(o[9866]) );
  AND U152 ( .A(p_input[9865]), .B(p_input[19865]), .Z(o[9865]) );
  AND U153 ( .A(p_input[9864]), .B(p_input[19864]), .Z(o[9864]) );
  AND U154 ( .A(p_input[9863]), .B(p_input[19863]), .Z(o[9863]) );
  AND U155 ( .A(p_input[9862]), .B(p_input[19862]), .Z(o[9862]) );
  AND U156 ( .A(p_input[9861]), .B(p_input[19861]), .Z(o[9861]) );
  AND U157 ( .A(p_input[9860]), .B(p_input[19860]), .Z(o[9860]) );
  AND U158 ( .A(p_input[985]), .B(p_input[10985]), .Z(o[985]) );
  AND U159 ( .A(p_input[9859]), .B(p_input[19859]), .Z(o[9859]) );
  AND U160 ( .A(p_input[9858]), .B(p_input[19858]), .Z(o[9858]) );
  AND U161 ( .A(p_input[9857]), .B(p_input[19857]), .Z(o[9857]) );
  AND U162 ( .A(p_input[9856]), .B(p_input[19856]), .Z(o[9856]) );
  AND U163 ( .A(p_input[9855]), .B(p_input[19855]), .Z(o[9855]) );
  AND U164 ( .A(p_input[9854]), .B(p_input[19854]), .Z(o[9854]) );
  AND U165 ( .A(p_input[9853]), .B(p_input[19853]), .Z(o[9853]) );
  AND U166 ( .A(p_input[9852]), .B(p_input[19852]), .Z(o[9852]) );
  AND U167 ( .A(p_input[9851]), .B(p_input[19851]), .Z(o[9851]) );
  AND U168 ( .A(p_input[9850]), .B(p_input[19850]), .Z(o[9850]) );
  AND U169 ( .A(p_input[984]), .B(p_input[10984]), .Z(o[984]) );
  AND U170 ( .A(p_input[9849]), .B(p_input[19849]), .Z(o[9849]) );
  AND U171 ( .A(p_input[9848]), .B(p_input[19848]), .Z(o[9848]) );
  AND U172 ( .A(p_input[9847]), .B(p_input[19847]), .Z(o[9847]) );
  AND U173 ( .A(p_input[9846]), .B(p_input[19846]), .Z(o[9846]) );
  AND U174 ( .A(p_input[9845]), .B(p_input[19845]), .Z(o[9845]) );
  AND U175 ( .A(p_input[9844]), .B(p_input[19844]), .Z(o[9844]) );
  AND U176 ( .A(p_input[9843]), .B(p_input[19843]), .Z(o[9843]) );
  AND U177 ( .A(p_input[9842]), .B(p_input[19842]), .Z(o[9842]) );
  AND U178 ( .A(p_input[9841]), .B(p_input[19841]), .Z(o[9841]) );
  AND U179 ( .A(p_input[9840]), .B(p_input[19840]), .Z(o[9840]) );
  AND U180 ( .A(p_input[983]), .B(p_input[10983]), .Z(o[983]) );
  AND U181 ( .A(p_input[9839]), .B(p_input[19839]), .Z(o[9839]) );
  AND U182 ( .A(p_input[9838]), .B(p_input[19838]), .Z(o[9838]) );
  AND U183 ( .A(p_input[9837]), .B(p_input[19837]), .Z(o[9837]) );
  AND U184 ( .A(p_input[9836]), .B(p_input[19836]), .Z(o[9836]) );
  AND U185 ( .A(p_input[9835]), .B(p_input[19835]), .Z(o[9835]) );
  AND U186 ( .A(p_input[9834]), .B(p_input[19834]), .Z(o[9834]) );
  AND U187 ( .A(p_input[9833]), .B(p_input[19833]), .Z(o[9833]) );
  AND U188 ( .A(p_input[9832]), .B(p_input[19832]), .Z(o[9832]) );
  AND U189 ( .A(p_input[9831]), .B(p_input[19831]), .Z(o[9831]) );
  AND U190 ( .A(p_input[9830]), .B(p_input[19830]), .Z(o[9830]) );
  AND U191 ( .A(p_input[982]), .B(p_input[10982]), .Z(o[982]) );
  AND U192 ( .A(p_input[9829]), .B(p_input[19829]), .Z(o[9829]) );
  AND U193 ( .A(p_input[9828]), .B(p_input[19828]), .Z(o[9828]) );
  AND U194 ( .A(p_input[9827]), .B(p_input[19827]), .Z(o[9827]) );
  AND U195 ( .A(p_input[9826]), .B(p_input[19826]), .Z(o[9826]) );
  AND U196 ( .A(p_input[9825]), .B(p_input[19825]), .Z(o[9825]) );
  AND U197 ( .A(p_input[9824]), .B(p_input[19824]), .Z(o[9824]) );
  AND U198 ( .A(p_input[9823]), .B(p_input[19823]), .Z(o[9823]) );
  AND U199 ( .A(p_input[9822]), .B(p_input[19822]), .Z(o[9822]) );
  AND U200 ( .A(p_input[9821]), .B(p_input[19821]), .Z(o[9821]) );
  AND U201 ( .A(p_input[9820]), .B(p_input[19820]), .Z(o[9820]) );
  AND U202 ( .A(p_input[981]), .B(p_input[10981]), .Z(o[981]) );
  AND U203 ( .A(p_input[9819]), .B(p_input[19819]), .Z(o[9819]) );
  AND U204 ( .A(p_input[9818]), .B(p_input[19818]), .Z(o[9818]) );
  AND U205 ( .A(p_input[9817]), .B(p_input[19817]), .Z(o[9817]) );
  AND U206 ( .A(p_input[9816]), .B(p_input[19816]), .Z(o[9816]) );
  AND U207 ( .A(p_input[9815]), .B(p_input[19815]), .Z(o[9815]) );
  AND U208 ( .A(p_input[9814]), .B(p_input[19814]), .Z(o[9814]) );
  AND U209 ( .A(p_input[9813]), .B(p_input[19813]), .Z(o[9813]) );
  AND U210 ( .A(p_input[9812]), .B(p_input[19812]), .Z(o[9812]) );
  AND U211 ( .A(p_input[9811]), .B(p_input[19811]), .Z(o[9811]) );
  AND U212 ( .A(p_input[9810]), .B(p_input[19810]), .Z(o[9810]) );
  AND U213 ( .A(p_input[980]), .B(p_input[10980]), .Z(o[980]) );
  AND U214 ( .A(p_input[9809]), .B(p_input[19809]), .Z(o[9809]) );
  AND U215 ( .A(p_input[9808]), .B(p_input[19808]), .Z(o[9808]) );
  AND U216 ( .A(p_input[9807]), .B(p_input[19807]), .Z(o[9807]) );
  AND U217 ( .A(p_input[9806]), .B(p_input[19806]), .Z(o[9806]) );
  AND U218 ( .A(p_input[9805]), .B(p_input[19805]), .Z(o[9805]) );
  AND U219 ( .A(p_input[9804]), .B(p_input[19804]), .Z(o[9804]) );
  AND U220 ( .A(p_input[9803]), .B(p_input[19803]), .Z(o[9803]) );
  AND U221 ( .A(p_input[9802]), .B(p_input[19802]), .Z(o[9802]) );
  AND U222 ( .A(p_input[9801]), .B(p_input[19801]), .Z(o[9801]) );
  AND U223 ( .A(p_input[9800]), .B(p_input[19800]), .Z(o[9800]) );
  AND U224 ( .A(p_input[97]), .B(p_input[10097]), .Z(o[97]) );
  AND U225 ( .A(p_input[979]), .B(p_input[10979]), .Z(o[979]) );
  AND U226 ( .A(p_input[9799]), .B(p_input[19799]), .Z(o[9799]) );
  AND U227 ( .A(p_input[9798]), .B(p_input[19798]), .Z(o[9798]) );
  AND U228 ( .A(p_input[9797]), .B(p_input[19797]), .Z(o[9797]) );
  AND U229 ( .A(p_input[9796]), .B(p_input[19796]), .Z(o[9796]) );
  AND U230 ( .A(p_input[9795]), .B(p_input[19795]), .Z(o[9795]) );
  AND U231 ( .A(p_input[9794]), .B(p_input[19794]), .Z(o[9794]) );
  AND U232 ( .A(p_input[9793]), .B(p_input[19793]), .Z(o[9793]) );
  AND U233 ( .A(p_input[9792]), .B(p_input[19792]), .Z(o[9792]) );
  AND U234 ( .A(p_input[9791]), .B(p_input[19791]), .Z(o[9791]) );
  AND U235 ( .A(p_input[9790]), .B(p_input[19790]), .Z(o[9790]) );
  AND U236 ( .A(p_input[978]), .B(p_input[10978]), .Z(o[978]) );
  AND U237 ( .A(p_input[9789]), .B(p_input[19789]), .Z(o[9789]) );
  AND U238 ( .A(p_input[9788]), .B(p_input[19788]), .Z(o[9788]) );
  AND U239 ( .A(p_input[9787]), .B(p_input[19787]), .Z(o[9787]) );
  AND U240 ( .A(p_input[9786]), .B(p_input[19786]), .Z(o[9786]) );
  AND U241 ( .A(p_input[9785]), .B(p_input[19785]), .Z(o[9785]) );
  AND U242 ( .A(p_input[9784]), .B(p_input[19784]), .Z(o[9784]) );
  AND U243 ( .A(p_input[9783]), .B(p_input[19783]), .Z(o[9783]) );
  AND U244 ( .A(p_input[9782]), .B(p_input[19782]), .Z(o[9782]) );
  AND U245 ( .A(p_input[9781]), .B(p_input[19781]), .Z(o[9781]) );
  AND U246 ( .A(p_input[9780]), .B(p_input[19780]), .Z(o[9780]) );
  AND U247 ( .A(p_input[977]), .B(p_input[10977]), .Z(o[977]) );
  AND U248 ( .A(p_input[9779]), .B(p_input[19779]), .Z(o[9779]) );
  AND U249 ( .A(p_input[9778]), .B(p_input[19778]), .Z(o[9778]) );
  AND U250 ( .A(p_input[9777]), .B(p_input[19777]), .Z(o[9777]) );
  AND U251 ( .A(p_input[9776]), .B(p_input[19776]), .Z(o[9776]) );
  AND U252 ( .A(p_input[9775]), .B(p_input[19775]), .Z(o[9775]) );
  AND U253 ( .A(p_input[9774]), .B(p_input[19774]), .Z(o[9774]) );
  AND U254 ( .A(p_input[9773]), .B(p_input[19773]), .Z(o[9773]) );
  AND U255 ( .A(p_input[9772]), .B(p_input[19772]), .Z(o[9772]) );
  AND U256 ( .A(p_input[9771]), .B(p_input[19771]), .Z(o[9771]) );
  AND U257 ( .A(p_input[9770]), .B(p_input[19770]), .Z(o[9770]) );
  AND U258 ( .A(p_input[976]), .B(p_input[10976]), .Z(o[976]) );
  AND U259 ( .A(p_input[9769]), .B(p_input[19769]), .Z(o[9769]) );
  AND U260 ( .A(p_input[9768]), .B(p_input[19768]), .Z(o[9768]) );
  AND U261 ( .A(p_input[9767]), .B(p_input[19767]), .Z(o[9767]) );
  AND U262 ( .A(p_input[9766]), .B(p_input[19766]), .Z(o[9766]) );
  AND U263 ( .A(p_input[9765]), .B(p_input[19765]), .Z(o[9765]) );
  AND U264 ( .A(p_input[9764]), .B(p_input[19764]), .Z(o[9764]) );
  AND U265 ( .A(p_input[9763]), .B(p_input[19763]), .Z(o[9763]) );
  AND U266 ( .A(p_input[9762]), .B(p_input[19762]), .Z(o[9762]) );
  AND U267 ( .A(p_input[9761]), .B(p_input[19761]), .Z(o[9761]) );
  AND U268 ( .A(p_input[9760]), .B(p_input[19760]), .Z(o[9760]) );
  AND U269 ( .A(p_input[975]), .B(p_input[10975]), .Z(o[975]) );
  AND U270 ( .A(p_input[9759]), .B(p_input[19759]), .Z(o[9759]) );
  AND U271 ( .A(p_input[9758]), .B(p_input[19758]), .Z(o[9758]) );
  AND U272 ( .A(p_input[9757]), .B(p_input[19757]), .Z(o[9757]) );
  AND U273 ( .A(p_input[9756]), .B(p_input[19756]), .Z(o[9756]) );
  AND U274 ( .A(p_input[9755]), .B(p_input[19755]), .Z(o[9755]) );
  AND U275 ( .A(p_input[9754]), .B(p_input[19754]), .Z(o[9754]) );
  AND U276 ( .A(p_input[9753]), .B(p_input[19753]), .Z(o[9753]) );
  AND U277 ( .A(p_input[9752]), .B(p_input[19752]), .Z(o[9752]) );
  AND U278 ( .A(p_input[9751]), .B(p_input[19751]), .Z(o[9751]) );
  AND U279 ( .A(p_input[9750]), .B(p_input[19750]), .Z(o[9750]) );
  AND U280 ( .A(p_input[974]), .B(p_input[10974]), .Z(o[974]) );
  AND U281 ( .A(p_input[9749]), .B(p_input[19749]), .Z(o[9749]) );
  AND U282 ( .A(p_input[9748]), .B(p_input[19748]), .Z(o[9748]) );
  AND U283 ( .A(p_input[9747]), .B(p_input[19747]), .Z(o[9747]) );
  AND U284 ( .A(p_input[9746]), .B(p_input[19746]), .Z(o[9746]) );
  AND U285 ( .A(p_input[9745]), .B(p_input[19745]), .Z(o[9745]) );
  AND U286 ( .A(p_input[9744]), .B(p_input[19744]), .Z(o[9744]) );
  AND U287 ( .A(p_input[9743]), .B(p_input[19743]), .Z(o[9743]) );
  AND U288 ( .A(p_input[9742]), .B(p_input[19742]), .Z(o[9742]) );
  AND U289 ( .A(p_input[9741]), .B(p_input[19741]), .Z(o[9741]) );
  AND U290 ( .A(p_input[9740]), .B(p_input[19740]), .Z(o[9740]) );
  AND U291 ( .A(p_input[973]), .B(p_input[10973]), .Z(o[973]) );
  AND U292 ( .A(p_input[9739]), .B(p_input[19739]), .Z(o[9739]) );
  AND U293 ( .A(p_input[9738]), .B(p_input[19738]), .Z(o[9738]) );
  AND U294 ( .A(p_input[9737]), .B(p_input[19737]), .Z(o[9737]) );
  AND U295 ( .A(p_input[9736]), .B(p_input[19736]), .Z(o[9736]) );
  AND U296 ( .A(p_input[9735]), .B(p_input[19735]), .Z(o[9735]) );
  AND U297 ( .A(p_input[9734]), .B(p_input[19734]), .Z(o[9734]) );
  AND U298 ( .A(p_input[9733]), .B(p_input[19733]), .Z(o[9733]) );
  AND U299 ( .A(p_input[9732]), .B(p_input[19732]), .Z(o[9732]) );
  AND U300 ( .A(p_input[9731]), .B(p_input[19731]), .Z(o[9731]) );
  AND U301 ( .A(p_input[9730]), .B(p_input[19730]), .Z(o[9730]) );
  AND U302 ( .A(p_input[972]), .B(p_input[10972]), .Z(o[972]) );
  AND U303 ( .A(p_input[9729]), .B(p_input[19729]), .Z(o[9729]) );
  AND U304 ( .A(p_input[9728]), .B(p_input[19728]), .Z(o[9728]) );
  AND U305 ( .A(p_input[9727]), .B(p_input[19727]), .Z(o[9727]) );
  AND U306 ( .A(p_input[9726]), .B(p_input[19726]), .Z(o[9726]) );
  AND U307 ( .A(p_input[9725]), .B(p_input[19725]), .Z(o[9725]) );
  AND U308 ( .A(p_input[9724]), .B(p_input[19724]), .Z(o[9724]) );
  AND U309 ( .A(p_input[9723]), .B(p_input[19723]), .Z(o[9723]) );
  AND U310 ( .A(p_input[9722]), .B(p_input[19722]), .Z(o[9722]) );
  AND U311 ( .A(p_input[9721]), .B(p_input[19721]), .Z(o[9721]) );
  AND U312 ( .A(p_input[9720]), .B(p_input[19720]), .Z(o[9720]) );
  AND U313 ( .A(p_input[971]), .B(p_input[10971]), .Z(o[971]) );
  AND U314 ( .A(p_input[9719]), .B(p_input[19719]), .Z(o[9719]) );
  AND U315 ( .A(p_input[9718]), .B(p_input[19718]), .Z(o[9718]) );
  AND U316 ( .A(p_input[9717]), .B(p_input[19717]), .Z(o[9717]) );
  AND U317 ( .A(p_input[9716]), .B(p_input[19716]), .Z(o[9716]) );
  AND U318 ( .A(p_input[9715]), .B(p_input[19715]), .Z(o[9715]) );
  AND U319 ( .A(p_input[9714]), .B(p_input[19714]), .Z(o[9714]) );
  AND U320 ( .A(p_input[9713]), .B(p_input[19713]), .Z(o[9713]) );
  AND U321 ( .A(p_input[9712]), .B(p_input[19712]), .Z(o[9712]) );
  AND U322 ( .A(p_input[9711]), .B(p_input[19711]), .Z(o[9711]) );
  AND U323 ( .A(p_input[9710]), .B(p_input[19710]), .Z(o[9710]) );
  AND U324 ( .A(p_input[970]), .B(p_input[10970]), .Z(o[970]) );
  AND U325 ( .A(p_input[9709]), .B(p_input[19709]), .Z(o[9709]) );
  AND U326 ( .A(p_input[9708]), .B(p_input[19708]), .Z(o[9708]) );
  AND U327 ( .A(p_input[9707]), .B(p_input[19707]), .Z(o[9707]) );
  AND U328 ( .A(p_input[9706]), .B(p_input[19706]), .Z(o[9706]) );
  AND U329 ( .A(p_input[9705]), .B(p_input[19705]), .Z(o[9705]) );
  AND U330 ( .A(p_input[9704]), .B(p_input[19704]), .Z(o[9704]) );
  AND U331 ( .A(p_input[9703]), .B(p_input[19703]), .Z(o[9703]) );
  AND U332 ( .A(p_input[9702]), .B(p_input[19702]), .Z(o[9702]) );
  AND U333 ( .A(p_input[9701]), .B(p_input[19701]), .Z(o[9701]) );
  AND U334 ( .A(p_input[9700]), .B(p_input[19700]), .Z(o[9700]) );
  AND U335 ( .A(p_input[96]), .B(p_input[10096]), .Z(o[96]) );
  AND U336 ( .A(p_input[969]), .B(p_input[10969]), .Z(o[969]) );
  AND U337 ( .A(p_input[9699]), .B(p_input[19699]), .Z(o[9699]) );
  AND U338 ( .A(p_input[9698]), .B(p_input[19698]), .Z(o[9698]) );
  AND U339 ( .A(p_input[9697]), .B(p_input[19697]), .Z(o[9697]) );
  AND U340 ( .A(p_input[9696]), .B(p_input[19696]), .Z(o[9696]) );
  AND U341 ( .A(p_input[9695]), .B(p_input[19695]), .Z(o[9695]) );
  AND U342 ( .A(p_input[9694]), .B(p_input[19694]), .Z(o[9694]) );
  AND U343 ( .A(p_input[9693]), .B(p_input[19693]), .Z(o[9693]) );
  AND U344 ( .A(p_input[9692]), .B(p_input[19692]), .Z(o[9692]) );
  AND U345 ( .A(p_input[9691]), .B(p_input[19691]), .Z(o[9691]) );
  AND U346 ( .A(p_input[9690]), .B(p_input[19690]), .Z(o[9690]) );
  AND U347 ( .A(p_input[968]), .B(p_input[10968]), .Z(o[968]) );
  AND U348 ( .A(p_input[9689]), .B(p_input[19689]), .Z(o[9689]) );
  AND U349 ( .A(p_input[9688]), .B(p_input[19688]), .Z(o[9688]) );
  AND U350 ( .A(p_input[9687]), .B(p_input[19687]), .Z(o[9687]) );
  AND U351 ( .A(p_input[9686]), .B(p_input[19686]), .Z(o[9686]) );
  AND U352 ( .A(p_input[9685]), .B(p_input[19685]), .Z(o[9685]) );
  AND U353 ( .A(p_input[9684]), .B(p_input[19684]), .Z(o[9684]) );
  AND U354 ( .A(p_input[9683]), .B(p_input[19683]), .Z(o[9683]) );
  AND U355 ( .A(p_input[9682]), .B(p_input[19682]), .Z(o[9682]) );
  AND U356 ( .A(p_input[9681]), .B(p_input[19681]), .Z(o[9681]) );
  AND U357 ( .A(p_input[9680]), .B(p_input[19680]), .Z(o[9680]) );
  AND U358 ( .A(p_input[967]), .B(p_input[10967]), .Z(o[967]) );
  AND U359 ( .A(p_input[9679]), .B(p_input[19679]), .Z(o[9679]) );
  AND U360 ( .A(p_input[9678]), .B(p_input[19678]), .Z(o[9678]) );
  AND U361 ( .A(p_input[9677]), .B(p_input[19677]), .Z(o[9677]) );
  AND U362 ( .A(p_input[9676]), .B(p_input[19676]), .Z(o[9676]) );
  AND U363 ( .A(p_input[9675]), .B(p_input[19675]), .Z(o[9675]) );
  AND U364 ( .A(p_input[9674]), .B(p_input[19674]), .Z(o[9674]) );
  AND U365 ( .A(p_input[9673]), .B(p_input[19673]), .Z(o[9673]) );
  AND U366 ( .A(p_input[9672]), .B(p_input[19672]), .Z(o[9672]) );
  AND U367 ( .A(p_input[9671]), .B(p_input[19671]), .Z(o[9671]) );
  AND U368 ( .A(p_input[9670]), .B(p_input[19670]), .Z(o[9670]) );
  AND U369 ( .A(p_input[966]), .B(p_input[10966]), .Z(o[966]) );
  AND U370 ( .A(p_input[9669]), .B(p_input[19669]), .Z(o[9669]) );
  AND U371 ( .A(p_input[9668]), .B(p_input[19668]), .Z(o[9668]) );
  AND U372 ( .A(p_input[9667]), .B(p_input[19667]), .Z(o[9667]) );
  AND U373 ( .A(p_input[9666]), .B(p_input[19666]), .Z(o[9666]) );
  AND U374 ( .A(p_input[9665]), .B(p_input[19665]), .Z(o[9665]) );
  AND U375 ( .A(p_input[9664]), .B(p_input[19664]), .Z(o[9664]) );
  AND U376 ( .A(p_input[9663]), .B(p_input[19663]), .Z(o[9663]) );
  AND U377 ( .A(p_input[9662]), .B(p_input[19662]), .Z(o[9662]) );
  AND U378 ( .A(p_input[9661]), .B(p_input[19661]), .Z(o[9661]) );
  AND U379 ( .A(p_input[9660]), .B(p_input[19660]), .Z(o[9660]) );
  AND U380 ( .A(p_input[965]), .B(p_input[10965]), .Z(o[965]) );
  AND U381 ( .A(p_input[9659]), .B(p_input[19659]), .Z(o[9659]) );
  AND U382 ( .A(p_input[9658]), .B(p_input[19658]), .Z(o[9658]) );
  AND U383 ( .A(p_input[9657]), .B(p_input[19657]), .Z(o[9657]) );
  AND U384 ( .A(p_input[9656]), .B(p_input[19656]), .Z(o[9656]) );
  AND U385 ( .A(p_input[9655]), .B(p_input[19655]), .Z(o[9655]) );
  AND U386 ( .A(p_input[9654]), .B(p_input[19654]), .Z(o[9654]) );
  AND U387 ( .A(p_input[9653]), .B(p_input[19653]), .Z(o[9653]) );
  AND U388 ( .A(p_input[9652]), .B(p_input[19652]), .Z(o[9652]) );
  AND U389 ( .A(p_input[9651]), .B(p_input[19651]), .Z(o[9651]) );
  AND U390 ( .A(p_input[9650]), .B(p_input[19650]), .Z(o[9650]) );
  AND U391 ( .A(p_input[964]), .B(p_input[10964]), .Z(o[964]) );
  AND U392 ( .A(p_input[9649]), .B(p_input[19649]), .Z(o[9649]) );
  AND U393 ( .A(p_input[9648]), .B(p_input[19648]), .Z(o[9648]) );
  AND U394 ( .A(p_input[9647]), .B(p_input[19647]), .Z(o[9647]) );
  AND U395 ( .A(p_input[9646]), .B(p_input[19646]), .Z(o[9646]) );
  AND U396 ( .A(p_input[9645]), .B(p_input[19645]), .Z(o[9645]) );
  AND U397 ( .A(p_input[9644]), .B(p_input[19644]), .Z(o[9644]) );
  AND U398 ( .A(p_input[9643]), .B(p_input[19643]), .Z(o[9643]) );
  AND U399 ( .A(p_input[9642]), .B(p_input[19642]), .Z(o[9642]) );
  AND U400 ( .A(p_input[9641]), .B(p_input[19641]), .Z(o[9641]) );
  AND U401 ( .A(p_input[9640]), .B(p_input[19640]), .Z(o[9640]) );
  AND U402 ( .A(p_input[963]), .B(p_input[10963]), .Z(o[963]) );
  AND U403 ( .A(p_input[9639]), .B(p_input[19639]), .Z(o[9639]) );
  AND U404 ( .A(p_input[9638]), .B(p_input[19638]), .Z(o[9638]) );
  AND U405 ( .A(p_input[9637]), .B(p_input[19637]), .Z(o[9637]) );
  AND U406 ( .A(p_input[9636]), .B(p_input[19636]), .Z(o[9636]) );
  AND U407 ( .A(p_input[9635]), .B(p_input[19635]), .Z(o[9635]) );
  AND U408 ( .A(p_input[9634]), .B(p_input[19634]), .Z(o[9634]) );
  AND U409 ( .A(p_input[9633]), .B(p_input[19633]), .Z(o[9633]) );
  AND U410 ( .A(p_input[9632]), .B(p_input[19632]), .Z(o[9632]) );
  AND U411 ( .A(p_input[9631]), .B(p_input[19631]), .Z(o[9631]) );
  AND U412 ( .A(p_input[9630]), .B(p_input[19630]), .Z(o[9630]) );
  AND U413 ( .A(p_input[962]), .B(p_input[10962]), .Z(o[962]) );
  AND U414 ( .A(p_input[9629]), .B(p_input[19629]), .Z(o[9629]) );
  AND U415 ( .A(p_input[9628]), .B(p_input[19628]), .Z(o[9628]) );
  AND U416 ( .A(p_input[9627]), .B(p_input[19627]), .Z(o[9627]) );
  AND U417 ( .A(p_input[9626]), .B(p_input[19626]), .Z(o[9626]) );
  AND U418 ( .A(p_input[9625]), .B(p_input[19625]), .Z(o[9625]) );
  AND U419 ( .A(p_input[9624]), .B(p_input[19624]), .Z(o[9624]) );
  AND U420 ( .A(p_input[9623]), .B(p_input[19623]), .Z(o[9623]) );
  AND U421 ( .A(p_input[9622]), .B(p_input[19622]), .Z(o[9622]) );
  AND U422 ( .A(p_input[9621]), .B(p_input[19621]), .Z(o[9621]) );
  AND U423 ( .A(p_input[9620]), .B(p_input[19620]), .Z(o[9620]) );
  AND U424 ( .A(p_input[961]), .B(p_input[10961]), .Z(o[961]) );
  AND U425 ( .A(p_input[9619]), .B(p_input[19619]), .Z(o[9619]) );
  AND U426 ( .A(p_input[9618]), .B(p_input[19618]), .Z(o[9618]) );
  AND U427 ( .A(p_input[9617]), .B(p_input[19617]), .Z(o[9617]) );
  AND U428 ( .A(p_input[9616]), .B(p_input[19616]), .Z(o[9616]) );
  AND U429 ( .A(p_input[9615]), .B(p_input[19615]), .Z(o[9615]) );
  AND U430 ( .A(p_input[9614]), .B(p_input[19614]), .Z(o[9614]) );
  AND U431 ( .A(p_input[9613]), .B(p_input[19613]), .Z(o[9613]) );
  AND U432 ( .A(p_input[9612]), .B(p_input[19612]), .Z(o[9612]) );
  AND U433 ( .A(p_input[9611]), .B(p_input[19611]), .Z(o[9611]) );
  AND U434 ( .A(p_input[9610]), .B(p_input[19610]), .Z(o[9610]) );
  AND U435 ( .A(p_input[960]), .B(p_input[10960]), .Z(o[960]) );
  AND U436 ( .A(p_input[9609]), .B(p_input[19609]), .Z(o[9609]) );
  AND U437 ( .A(p_input[9608]), .B(p_input[19608]), .Z(o[9608]) );
  AND U438 ( .A(p_input[9607]), .B(p_input[19607]), .Z(o[9607]) );
  AND U439 ( .A(p_input[9606]), .B(p_input[19606]), .Z(o[9606]) );
  AND U440 ( .A(p_input[9605]), .B(p_input[19605]), .Z(o[9605]) );
  AND U441 ( .A(p_input[9604]), .B(p_input[19604]), .Z(o[9604]) );
  AND U442 ( .A(p_input[9603]), .B(p_input[19603]), .Z(o[9603]) );
  AND U443 ( .A(p_input[9602]), .B(p_input[19602]), .Z(o[9602]) );
  AND U444 ( .A(p_input[9601]), .B(p_input[19601]), .Z(o[9601]) );
  AND U445 ( .A(p_input[9600]), .B(p_input[19600]), .Z(o[9600]) );
  AND U446 ( .A(p_input[95]), .B(p_input[10095]), .Z(o[95]) );
  AND U447 ( .A(p_input[959]), .B(p_input[10959]), .Z(o[959]) );
  AND U448 ( .A(p_input[9599]), .B(p_input[19599]), .Z(o[9599]) );
  AND U449 ( .A(p_input[9598]), .B(p_input[19598]), .Z(o[9598]) );
  AND U450 ( .A(p_input[9597]), .B(p_input[19597]), .Z(o[9597]) );
  AND U451 ( .A(p_input[9596]), .B(p_input[19596]), .Z(o[9596]) );
  AND U452 ( .A(p_input[9595]), .B(p_input[19595]), .Z(o[9595]) );
  AND U453 ( .A(p_input[9594]), .B(p_input[19594]), .Z(o[9594]) );
  AND U454 ( .A(p_input[9593]), .B(p_input[19593]), .Z(o[9593]) );
  AND U455 ( .A(p_input[9592]), .B(p_input[19592]), .Z(o[9592]) );
  AND U456 ( .A(p_input[9591]), .B(p_input[19591]), .Z(o[9591]) );
  AND U457 ( .A(p_input[9590]), .B(p_input[19590]), .Z(o[9590]) );
  AND U458 ( .A(p_input[958]), .B(p_input[10958]), .Z(o[958]) );
  AND U459 ( .A(p_input[9589]), .B(p_input[19589]), .Z(o[9589]) );
  AND U460 ( .A(p_input[9588]), .B(p_input[19588]), .Z(o[9588]) );
  AND U461 ( .A(p_input[9587]), .B(p_input[19587]), .Z(o[9587]) );
  AND U462 ( .A(p_input[9586]), .B(p_input[19586]), .Z(o[9586]) );
  AND U463 ( .A(p_input[9585]), .B(p_input[19585]), .Z(o[9585]) );
  AND U464 ( .A(p_input[9584]), .B(p_input[19584]), .Z(o[9584]) );
  AND U465 ( .A(p_input[9583]), .B(p_input[19583]), .Z(o[9583]) );
  AND U466 ( .A(p_input[9582]), .B(p_input[19582]), .Z(o[9582]) );
  AND U467 ( .A(p_input[9581]), .B(p_input[19581]), .Z(o[9581]) );
  AND U468 ( .A(p_input[9580]), .B(p_input[19580]), .Z(o[9580]) );
  AND U469 ( .A(p_input[957]), .B(p_input[10957]), .Z(o[957]) );
  AND U470 ( .A(p_input[9579]), .B(p_input[19579]), .Z(o[9579]) );
  AND U471 ( .A(p_input[9578]), .B(p_input[19578]), .Z(o[9578]) );
  AND U472 ( .A(p_input[9577]), .B(p_input[19577]), .Z(o[9577]) );
  AND U473 ( .A(p_input[9576]), .B(p_input[19576]), .Z(o[9576]) );
  AND U474 ( .A(p_input[9575]), .B(p_input[19575]), .Z(o[9575]) );
  AND U475 ( .A(p_input[9574]), .B(p_input[19574]), .Z(o[9574]) );
  AND U476 ( .A(p_input[9573]), .B(p_input[19573]), .Z(o[9573]) );
  AND U477 ( .A(p_input[9572]), .B(p_input[19572]), .Z(o[9572]) );
  AND U478 ( .A(p_input[9571]), .B(p_input[19571]), .Z(o[9571]) );
  AND U479 ( .A(p_input[9570]), .B(p_input[19570]), .Z(o[9570]) );
  AND U480 ( .A(p_input[956]), .B(p_input[10956]), .Z(o[956]) );
  AND U481 ( .A(p_input[9569]), .B(p_input[19569]), .Z(o[9569]) );
  AND U482 ( .A(p_input[9568]), .B(p_input[19568]), .Z(o[9568]) );
  AND U483 ( .A(p_input[9567]), .B(p_input[19567]), .Z(o[9567]) );
  AND U484 ( .A(p_input[9566]), .B(p_input[19566]), .Z(o[9566]) );
  AND U485 ( .A(p_input[9565]), .B(p_input[19565]), .Z(o[9565]) );
  AND U486 ( .A(p_input[9564]), .B(p_input[19564]), .Z(o[9564]) );
  AND U487 ( .A(p_input[9563]), .B(p_input[19563]), .Z(o[9563]) );
  AND U488 ( .A(p_input[9562]), .B(p_input[19562]), .Z(o[9562]) );
  AND U489 ( .A(p_input[9561]), .B(p_input[19561]), .Z(o[9561]) );
  AND U490 ( .A(p_input[9560]), .B(p_input[19560]), .Z(o[9560]) );
  AND U491 ( .A(p_input[955]), .B(p_input[10955]), .Z(o[955]) );
  AND U492 ( .A(p_input[9559]), .B(p_input[19559]), .Z(o[9559]) );
  AND U493 ( .A(p_input[9558]), .B(p_input[19558]), .Z(o[9558]) );
  AND U494 ( .A(p_input[9557]), .B(p_input[19557]), .Z(o[9557]) );
  AND U495 ( .A(p_input[9556]), .B(p_input[19556]), .Z(o[9556]) );
  AND U496 ( .A(p_input[9555]), .B(p_input[19555]), .Z(o[9555]) );
  AND U497 ( .A(p_input[9554]), .B(p_input[19554]), .Z(o[9554]) );
  AND U498 ( .A(p_input[9553]), .B(p_input[19553]), .Z(o[9553]) );
  AND U499 ( .A(p_input[9552]), .B(p_input[19552]), .Z(o[9552]) );
  AND U500 ( .A(p_input[9551]), .B(p_input[19551]), .Z(o[9551]) );
  AND U501 ( .A(p_input[9550]), .B(p_input[19550]), .Z(o[9550]) );
  AND U502 ( .A(p_input[954]), .B(p_input[10954]), .Z(o[954]) );
  AND U503 ( .A(p_input[9549]), .B(p_input[19549]), .Z(o[9549]) );
  AND U504 ( .A(p_input[9548]), .B(p_input[19548]), .Z(o[9548]) );
  AND U505 ( .A(p_input[9547]), .B(p_input[19547]), .Z(o[9547]) );
  AND U506 ( .A(p_input[9546]), .B(p_input[19546]), .Z(o[9546]) );
  AND U507 ( .A(p_input[9545]), .B(p_input[19545]), .Z(o[9545]) );
  AND U508 ( .A(p_input[9544]), .B(p_input[19544]), .Z(o[9544]) );
  AND U509 ( .A(p_input[9543]), .B(p_input[19543]), .Z(o[9543]) );
  AND U510 ( .A(p_input[9542]), .B(p_input[19542]), .Z(o[9542]) );
  AND U511 ( .A(p_input[9541]), .B(p_input[19541]), .Z(o[9541]) );
  AND U512 ( .A(p_input[9540]), .B(p_input[19540]), .Z(o[9540]) );
  AND U513 ( .A(p_input[953]), .B(p_input[10953]), .Z(o[953]) );
  AND U514 ( .A(p_input[9539]), .B(p_input[19539]), .Z(o[9539]) );
  AND U515 ( .A(p_input[9538]), .B(p_input[19538]), .Z(o[9538]) );
  AND U516 ( .A(p_input[9537]), .B(p_input[19537]), .Z(o[9537]) );
  AND U517 ( .A(p_input[9536]), .B(p_input[19536]), .Z(o[9536]) );
  AND U518 ( .A(p_input[9535]), .B(p_input[19535]), .Z(o[9535]) );
  AND U519 ( .A(p_input[9534]), .B(p_input[19534]), .Z(o[9534]) );
  AND U520 ( .A(p_input[9533]), .B(p_input[19533]), .Z(o[9533]) );
  AND U521 ( .A(p_input[9532]), .B(p_input[19532]), .Z(o[9532]) );
  AND U522 ( .A(p_input[9531]), .B(p_input[19531]), .Z(o[9531]) );
  AND U523 ( .A(p_input[9530]), .B(p_input[19530]), .Z(o[9530]) );
  AND U524 ( .A(p_input[952]), .B(p_input[10952]), .Z(o[952]) );
  AND U525 ( .A(p_input[9529]), .B(p_input[19529]), .Z(o[9529]) );
  AND U526 ( .A(p_input[9528]), .B(p_input[19528]), .Z(o[9528]) );
  AND U527 ( .A(p_input[9527]), .B(p_input[19527]), .Z(o[9527]) );
  AND U528 ( .A(p_input[9526]), .B(p_input[19526]), .Z(o[9526]) );
  AND U529 ( .A(p_input[9525]), .B(p_input[19525]), .Z(o[9525]) );
  AND U530 ( .A(p_input[9524]), .B(p_input[19524]), .Z(o[9524]) );
  AND U531 ( .A(p_input[9523]), .B(p_input[19523]), .Z(o[9523]) );
  AND U532 ( .A(p_input[9522]), .B(p_input[19522]), .Z(o[9522]) );
  AND U533 ( .A(p_input[9521]), .B(p_input[19521]), .Z(o[9521]) );
  AND U534 ( .A(p_input[9520]), .B(p_input[19520]), .Z(o[9520]) );
  AND U535 ( .A(p_input[951]), .B(p_input[10951]), .Z(o[951]) );
  AND U536 ( .A(p_input[9519]), .B(p_input[19519]), .Z(o[9519]) );
  AND U537 ( .A(p_input[9518]), .B(p_input[19518]), .Z(o[9518]) );
  AND U538 ( .A(p_input[9517]), .B(p_input[19517]), .Z(o[9517]) );
  AND U539 ( .A(p_input[9516]), .B(p_input[19516]), .Z(o[9516]) );
  AND U540 ( .A(p_input[9515]), .B(p_input[19515]), .Z(o[9515]) );
  AND U541 ( .A(p_input[9514]), .B(p_input[19514]), .Z(o[9514]) );
  AND U542 ( .A(p_input[9513]), .B(p_input[19513]), .Z(o[9513]) );
  AND U543 ( .A(p_input[9512]), .B(p_input[19512]), .Z(o[9512]) );
  AND U544 ( .A(p_input[9511]), .B(p_input[19511]), .Z(o[9511]) );
  AND U545 ( .A(p_input[9510]), .B(p_input[19510]), .Z(o[9510]) );
  AND U546 ( .A(p_input[950]), .B(p_input[10950]), .Z(o[950]) );
  AND U547 ( .A(p_input[9509]), .B(p_input[19509]), .Z(o[9509]) );
  AND U548 ( .A(p_input[9508]), .B(p_input[19508]), .Z(o[9508]) );
  AND U549 ( .A(p_input[9507]), .B(p_input[19507]), .Z(o[9507]) );
  AND U550 ( .A(p_input[9506]), .B(p_input[19506]), .Z(o[9506]) );
  AND U551 ( .A(p_input[9505]), .B(p_input[19505]), .Z(o[9505]) );
  AND U552 ( .A(p_input[9504]), .B(p_input[19504]), .Z(o[9504]) );
  AND U553 ( .A(p_input[9503]), .B(p_input[19503]), .Z(o[9503]) );
  AND U554 ( .A(p_input[9502]), .B(p_input[19502]), .Z(o[9502]) );
  AND U555 ( .A(p_input[9501]), .B(p_input[19501]), .Z(o[9501]) );
  AND U556 ( .A(p_input[9500]), .B(p_input[19500]), .Z(o[9500]) );
  AND U557 ( .A(p_input[94]), .B(p_input[10094]), .Z(o[94]) );
  AND U558 ( .A(p_input[949]), .B(p_input[10949]), .Z(o[949]) );
  AND U559 ( .A(p_input[9499]), .B(p_input[19499]), .Z(o[9499]) );
  AND U560 ( .A(p_input[9498]), .B(p_input[19498]), .Z(o[9498]) );
  AND U561 ( .A(p_input[9497]), .B(p_input[19497]), .Z(o[9497]) );
  AND U562 ( .A(p_input[9496]), .B(p_input[19496]), .Z(o[9496]) );
  AND U563 ( .A(p_input[9495]), .B(p_input[19495]), .Z(o[9495]) );
  AND U564 ( .A(p_input[9494]), .B(p_input[19494]), .Z(o[9494]) );
  AND U565 ( .A(p_input[9493]), .B(p_input[19493]), .Z(o[9493]) );
  AND U566 ( .A(p_input[9492]), .B(p_input[19492]), .Z(o[9492]) );
  AND U567 ( .A(p_input[9491]), .B(p_input[19491]), .Z(o[9491]) );
  AND U568 ( .A(p_input[9490]), .B(p_input[19490]), .Z(o[9490]) );
  AND U569 ( .A(p_input[948]), .B(p_input[10948]), .Z(o[948]) );
  AND U570 ( .A(p_input[9489]), .B(p_input[19489]), .Z(o[9489]) );
  AND U571 ( .A(p_input[9488]), .B(p_input[19488]), .Z(o[9488]) );
  AND U572 ( .A(p_input[9487]), .B(p_input[19487]), .Z(o[9487]) );
  AND U573 ( .A(p_input[9486]), .B(p_input[19486]), .Z(o[9486]) );
  AND U574 ( .A(p_input[9485]), .B(p_input[19485]), .Z(o[9485]) );
  AND U575 ( .A(p_input[9484]), .B(p_input[19484]), .Z(o[9484]) );
  AND U576 ( .A(p_input[9483]), .B(p_input[19483]), .Z(o[9483]) );
  AND U577 ( .A(p_input[9482]), .B(p_input[19482]), .Z(o[9482]) );
  AND U578 ( .A(p_input[9481]), .B(p_input[19481]), .Z(o[9481]) );
  AND U579 ( .A(p_input[9480]), .B(p_input[19480]), .Z(o[9480]) );
  AND U580 ( .A(p_input[947]), .B(p_input[10947]), .Z(o[947]) );
  AND U581 ( .A(p_input[9479]), .B(p_input[19479]), .Z(o[9479]) );
  AND U582 ( .A(p_input[9478]), .B(p_input[19478]), .Z(o[9478]) );
  AND U583 ( .A(p_input[9477]), .B(p_input[19477]), .Z(o[9477]) );
  AND U584 ( .A(p_input[9476]), .B(p_input[19476]), .Z(o[9476]) );
  AND U585 ( .A(p_input[9475]), .B(p_input[19475]), .Z(o[9475]) );
  AND U586 ( .A(p_input[9474]), .B(p_input[19474]), .Z(o[9474]) );
  AND U587 ( .A(p_input[9473]), .B(p_input[19473]), .Z(o[9473]) );
  AND U588 ( .A(p_input[9472]), .B(p_input[19472]), .Z(o[9472]) );
  AND U589 ( .A(p_input[9471]), .B(p_input[19471]), .Z(o[9471]) );
  AND U590 ( .A(p_input[9470]), .B(p_input[19470]), .Z(o[9470]) );
  AND U591 ( .A(p_input[946]), .B(p_input[10946]), .Z(o[946]) );
  AND U592 ( .A(p_input[9469]), .B(p_input[19469]), .Z(o[9469]) );
  AND U593 ( .A(p_input[9468]), .B(p_input[19468]), .Z(o[9468]) );
  AND U594 ( .A(p_input[9467]), .B(p_input[19467]), .Z(o[9467]) );
  AND U595 ( .A(p_input[9466]), .B(p_input[19466]), .Z(o[9466]) );
  AND U596 ( .A(p_input[9465]), .B(p_input[19465]), .Z(o[9465]) );
  AND U597 ( .A(p_input[9464]), .B(p_input[19464]), .Z(o[9464]) );
  AND U598 ( .A(p_input[9463]), .B(p_input[19463]), .Z(o[9463]) );
  AND U599 ( .A(p_input[9462]), .B(p_input[19462]), .Z(o[9462]) );
  AND U600 ( .A(p_input[9461]), .B(p_input[19461]), .Z(o[9461]) );
  AND U601 ( .A(p_input[9460]), .B(p_input[19460]), .Z(o[9460]) );
  AND U602 ( .A(p_input[945]), .B(p_input[10945]), .Z(o[945]) );
  AND U603 ( .A(p_input[9459]), .B(p_input[19459]), .Z(o[9459]) );
  AND U604 ( .A(p_input[9458]), .B(p_input[19458]), .Z(o[9458]) );
  AND U605 ( .A(p_input[9457]), .B(p_input[19457]), .Z(o[9457]) );
  AND U606 ( .A(p_input[9456]), .B(p_input[19456]), .Z(o[9456]) );
  AND U607 ( .A(p_input[9455]), .B(p_input[19455]), .Z(o[9455]) );
  AND U608 ( .A(p_input[9454]), .B(p_input[19454]), .Z(o[9454]) );
  AND U609 ( .A(p_input[9453]), .B(p_input[19453]), .Z(o[9453]) );
  AND U610 ( .A(p_input[9452]), .B(p_input[19452]), .Z(o[9452]) );
  AND U611 ( .A(p_input[9451]), .B(p_input[19451]), .Z(o[9451]) );
  AND U612 ( .A(p_input[9450]), .B(p_input[19450]), .Z(o[9450]) );
  AND U613 ( .A(p_input[944]), .B(p_input[10944]), .Z(o[944]) );
  AND U614 ( .A(p_input[9449]), .B(p_input[19449]), .Z(o[9449]) );
  AND U615 ( .A(p_input[9448]), .B(p_input[19448]), .Z(o[9448]) );
  AND U616 ( .A(p_input[9447]), .B(p_input[19447]), .Z(o[9447]) );
  AND U617 ( .A(p_input[9446]), .B(p_input[19446]), .Z(o[9446]) );
  AND U618 ( .A(p_input[9445]), .B(p_input[19445]), .Z(o[9445]) );
  AND U619 ( .A(p_input[9444]), .B(p_input[19444]), .Z(o[9444]) );
  AND U620 ( .A(p_input[9443]), .B(p_input[19443]), .Z(o[9443]) );
  AND U621 ( .A(p_input[9442]), .B(p_input[19442]), .Z(o[9442]) );
  AND U622 ( .A(p_input[9441]), .B(p_input[19441]), .Z(o[9441]) );
  AND U623 ( .A(p_input[9440]), .B(p_input[19440]), .Z(o[9440]) );
  AND U624 ( .A(p_input[943]), .B(p_input[10943]), .Z(o[943]) );
  AND U625 ( .A(p_input[9439]), .B(p_input[19439]), .Z(o[9439]) );
  AND U626 ( .A(p_input[9438]), .B(p_input[19438]), .Z(o[9438]) );
  AND U627 ( .A(p_input[9437]), .B(p_input[19437]), .Z(o[9437]) );
  AND U628 ( .A(p_input[9436]), .B(p_input[19436]), .Z(o[9436]) );
  AND U629 ( .A(p_input[9435]), .B(p_input[19435]), .Z(o[9435]) );
  AND U630 ( .A(p_input[9434]), .B(p_input[19434]), .Z(o[9434]) );
  AND U631 ( .A(p_input[9433]), .B(p_input[19433]), .Z(o[9433]) );
  AND U632 ( .A(p_input[9432]), .B(p_input[19432]), .Z(o[9432]) );
  AND U633 ( .A(p_input[9431]), .B(p_input[19431]), .Z(o[9431]) );
  AND U634 ( .A(p_input[9430]), .B(p_input[19430]), .Z(o[9430]) );
  AND U635 ( .A(p_input[942]), .B(p_input[10942]), .Z(o[942]) );
  AND U636 ( .A(p_input[9429]), .B(p_input[19429]), .Z(o[9429]) );
  AND U637 ( .A(p_input[9428]), .B(p_input[19428]), .Z(o[9428]) );
  AND U638 ( .A(p_input[9427]), .B(p_input[19427]), .Z(o[9427]) );
  AND U639 ( .A(p_input[9426]), .B(p_input[19426]), .Z(o[9426]) );
  AND U640 ( .A(p_input[9425]), .B(p_input[19425]), .Z(o[9425]) );
  AND U641 ( .A(p_input[9424]), .B(p_input[19424]), .Z(o[9424]) );
  AND U642 ( .A(p_input[9423]), .B(p_input[19423]), .Z(o[9423]) );
  AND U643 ( .A(p_input[9422]), .B(p_input[19422]), .Z(o[9422]) );
  AND U644 ( .A(p_input[9421]), .B(p_input[19421]), .Z(o[9421]) );
  AND U645 ( .A(p_input[9420]), .B(p_input[19420]), .Z(o[9420]) );
  AND U646 ( .A(p_input[941]), .B(p_input[10941]), .Z(o[941]) );
  AND U647 ( .A(p_input[9419]), .B(p_input[19419]), .Z(o[9419]) );
  AND U648 ( .A(p_input[9418]), .B(p_input[19418]), .Z(o[9418]) );
  AND U649 ( .A(p_input[9417]), .B(p_input[19417]), .Z(o[9417]) );
  AND U650 ( .A(p_input[9416]), .B(p_input[19416]), .Z(o[9416]) );
  AND U651 ( .A(p_input[9415]), .B(p_input[19415]), .Z(o[9415]) );
  AND U652 ( .A(p_input[9414]), .B(p_input[19414]), .Z(o[9414]) );
  AND U653 ( .A(p_input[9413]), .B(p_input[19413]), .Z(o[9413]) );
  AND U654 ( .A(p_input[9412]), .B(p_input[19412]), .Z(o[9412]) );
  AND U655 ( .A(p_input[9411]), .B(p_input[19411]), .Z(o[9411]) );
  AND U656 ( .A(p_input[9410]), .B(p_input[19410]), .Z(o[9410]) );
  AND U657 ( .A(p_input[940]), .B(p_input[10940]), .Z(o[940]) );
  AND U658 ( .A(p_input[9409]), .B(p_input[19409]), .Z(o[9409]) );
  AND U659 ( .A(p_input[9408]), .B(p_input[19408]), .Z(o[9408]) );
  AND U660 ( .A(p_input[9407]), .B(p_input[19407]), .Z(o[9407]) );
  AND U661 ( .A(p_input[9406]), .B(p_input[19406]), .Z(o[9406]) );
  AND U662 ( .A(p_input[9405]), .B(p_input[19405]), .Z(o[9405]) );
  AND U663 ( .A(p_input[9404]), .B(p_input[19404]), .Z(o[9404]) );
  AND U664 ( .A(p_input[9403]), .B(p_input[19403]), .Z(o[9403]) );
  AND U665 ( .A(p_input[9402]), .B(p_input[19402]), .Z(o[9402]) );
  AND U666 ( .A(p_input[9401]), .B(p_input[19401]), .Z(o[9401]) );
  AND U667 ( .A(p_input[9400]), .B(p_input[19400]), .Z(o[9400]) );
  AND U668 ( .A(p_input[93]), .B(p_input[10093]), .Z(o[93]) );
  AND U669 ( .A(p_input[939]), .B(p_input[10939]), .Z(o[939]) );
  AND U670 ( .A(p_input[9399]), .B(p_input[19399]), .Z(o[9399]) );
  AND U671 ( .A(p_input[9398]), .B(p_input[19398]), .Z(o[9398]) );
  AND U672 ( .A(p_input[9397]), .B(p_input[19397]), .Z(o[9397]) );
  AND U673 ( .A(p_input[9396]), .B(p_input[19396]), .Z(o[9396]) );
  AND U674 ( .A(p_input[9395]), .B(p_input[19395]), .Z(o[9395]) );
  AND U675 ( .A(p_input[9394]), .B(p_input[19394]), .Z(o[9394]) );
  AND U676 ( .A(p_input[9393]), .B(p_input[19393]), .Z(o[9393]) );
  AND U677 ( .A(p_input[9392]), .B(p_input[19392]), .Z(o[9392]) );
  AND U678 ( .A(p_input[9391]), .B(p_input[19391]), .Z(o[9391]) );
  AND U679 ( .A(p_input[9390]), .B(p_input[19390]), .Z(o[9390]) );
  AND U680 ( .A(p_input[938]), .B(p_input[10938]), .Z(o[938]) );
  AND U681 ( .A(p_input[9389]), .B(p_input[19389]), .Z(o[9389]) );
  AND U682 ( .A(p_input[9388]), .B(p_input[19388]), .Z(o[9388]) );
  AND U683 ( .A(p_input[9387]), .B(p_input[19387]), .Z(o[9387]) );
  AND U684 ( .A(p_input[9386]), .B(p_input[19386]), .Z(o[9386]) );
  AND U685 ( .A(p_input[9385]), .B(p_input[19385]), .Z(o[9385]) );
  AND U686 ( .A(p_input[9384]), .B(p_input[19384]), .Z(o[9384]) );
  AND U687 ( .A(p_input[9383]), .B(p_input[19383]), .Z(o[9383]) );
  AND U688 ( .A(p_input[9382]), .B(p_input[19382]), .Z(o[9382]) );
  AND U689 ( .A(p_input[9381]), .B(p_input[19381]), .Z(o[9381]) );
  AND U690 ( .A(p_input[9380]), .B(p_input[19380]), .Z(o[9380]) );
  AND U691 ( .A(p_input[937]), .B(p_input[10937]), .Z(o[937]) );
  AND U692 ( .A(p_input[9379]), .B(p_input[19379]), .Z(o[9379]) );
  AND U693 ( .A(p_input[9378]), .B(p_input[19378]), .Z(o[9378]) );
  AND U694 ( .A(p_input[9377]), .B(p_input[19377]), .Z(o[9377]) );
  AND U695 ( .A(p_input[9376]), .B(p_input[19376]), .Z(o[9376]) );
  AND U696 ( .A(p_input[9375]), .B(p_input[19375]), .Z(o[9375]) );
  AND U697 ( .A(p_input[9374]), .B(p_input[19374]), .Z(o[9374]) );
  AND U698 ( .A(p_input[9373]), .B(p_input[19373]), .Z(o[9373]) );
  AND U699 ( .A(p_input[9372]), .B(p_input[19372]), .Z(o[9372]) );
  AND U700 ( .A(p_input[9371]), .B(p_input[19371]), .Z(o[9371]) );
  AND U701 ( .A(p_input[9370]), .B(p_input[19370]), .Z(o[9370]) );
  AND U702 ( .A(p_input[936]), .B(p_input[10936]), .Z(o[936]) );
  AND U703 ( .A(p_input[9369]), .B(p_input[19369]), .Z(o[9369]) );
  AND U704 ( .A(p_input[9368]), .B(p_input[19368]), .Z(o[9368]) );
  AND U705 ( .A(p_input[9367]), .B(p_input[19367]), .Z(o[9367]) );
  AND U706 ( .A(p_input[9366]), .B(p_input[19366]), .Z(o[9366]) );
  AND U707 ( .A(p_input[9365]), .B(p_input[19365]), .Z(o[9365]) );
  AND U708 ( .A(p_input[9364]), .B(p_input[19364]), .Z(o[9364]) );
  AND U709 ( .A(p_input[9363]), .B(p_input[19363]), .Z(o[9363]) );
  AND U710 ( .A(p_input[9362]), .B(p_input[19362]), .Z(o[9362]) );
  AND U711 ( .A(p_input[9361]), .B(p_input[19361]), .Z(o[9361]) );
  AND U712 ( .A(p_input[9360]), .B(p_input[19360]), .Z(o[9360]) );
  AND U713 ( .A(p_input[935]), .B(p_input[10935]), .Z(o[935]) );
  AND U714 ( .A(p_input[9359]), .B(p_input[19359]), .Z(o[9359]) );
  AND U715 ( .A(p_input[9358]), .B(p_input[19358]), .Z(o[9358]) );
  AND U716 ( .A(p_input[9357]), .B(p_input[19357]), .Z(o[9357]) );
  AND U717 ( .A(p_input[9356]), .B(p_input[19356]), .Z(o[9356]) );
  AND U718 ( .A(p_input[9355]), .B(p_input[19355]), .Z(o[9355]) );
  AND U719 ( .A(p_input[9354]), .B(p_input[19354]), .Z(o[9354]) );
  AND U720 ( .A(p_input[9353]), .B(p_input[19353]), .Z(o[9353]) );
  AND U721 ( .A(p_input[9352]), .B(p_input[19352]), .Z(o[9352]) );
  AND U722 ( .A(p_input[9351]), .B(p_input[19351]), .Z(o[9351]) );
  AND U723 ( .A(p_input[9350]), .B(p_input[19350]), .Z(o[9350]) );
  AND U724 ( .A(p_input[934]), .B(p_input[10934]), .Z(o[934]) );
  AND U725 ( .A(p_input[9349]), .B(p_input[19349]), .Z(o[9349]) );
  AND U726 ( .A(p_input[9348]), .B(p_input[19348]), .Z(o[9348]) );
  AND U727 ( .A(p_input[9347]), .B(p_input[19347]), .Z(o[9347]) );
  AND U728 ( .A(p_input[9346]), .B(p_input[19346]), .Z(o[9346]) );
  AND U729 ( .A(p_input[9345]), .B(p_input[19345]), .Z(o[9345]) );
  AND U730 ( .A(p_input[9344]), .B(p_input[19344]), .Z(o[9344]) );
  AND U731 ( .A(p_input[9343]), .B(p_input[19343]), .Z(o[9343]) );
  AND U732 ( .A(p_input[9342]), .B(p_input[19342]), .Z(o[9342]) );
  AND U733 ( .A(p_input[9341]), .B(p_input[19341]), .Z(o[9341]) );
  AND U734 ( .A(p_input[9340]), .B(p_input[19340]), .Z(o[9340]) );
  AND U735 ( .A(p_input[933]), .B(p_input[10933]), .Z(o[933]) );
  AND U736 ( .A(p_input[9339]), .B(p_input[19339]), .Z(o[9339]) );
  AND U737 ( .A(p_input[9338]), .B(p_input[19338]), .Z(o[9338]) );
  AND U738 ( .A(p_input[9337]), .B(p_input[19337]), .Z(o[9337]) );
  AND U739 ( .A(p_input[9336]), .B(p_input[19336]), .Z(o[9336]) );
  AND U740 ( .A(p_input[9335]), .B(p_input[19335]), .Z(o[9335]) );
  AND U741 ( .A(p_input[9334]), .B(p_input[19334]), .Z(o[9334]) );
  AND U742 ( .A(p_input[9333]), .B(p_input[19333]), .Z(o[9333]) );
  AND U743 ( .A(p_input[9332]), .B(p_input[19332]), .Z(o[9332]) );
  AND U744 ( .A(p_input[9331]), .B(p_input[19331]), .Z(o[9331]) );
  AND U745 ( .A(p_input[9330]), .B(p_input[19330]), .Z(o[9330]) );
  AND U746 ( .A(p_input[932]), .B(p_input[10932]), .Z(o[932]) );
  AND U747 ( .A(p_input[9329]), .B(p_input[19329]), .Z(o[9329]) );
  AND U748 ( .A(p_input[9328]), .B(p_input[19328]), .Z(o[9328]) );
  AND U749 ( .A(p_input[9327]), .B(p_input[19327]), .Z(o[9327]) );
  AND U750 ( .A(p_input[9326]), .B(p_input[19326]), .Z(o[9326]) );
  AND U751 ( .A(p_input[9325]), .B(p_input[19325]), .Z(o[9325]) );
  AND U752 ( .A(p_input[9324]), .B(p_input[19324]), .Z(o[9324]) );
  AND U753 ( .A(p_input[9323]), .B(p_input[19323]), .Z(o[9323]) );
  AND U754 ( .A(p_input[9322]), .B(p_input[19322]), .Z(o[9322]) );
  AND U755 ( .A(p_input[9321]), .B(p_input[19321]), .Z(o[9321]) );
  AND U756 ( .A(p_input[9320]), .B(p_input[19320]), .Z(o[9320]) );
  AND U757 ( .A(p_input[931]), .B(p_input[10931]), .Z(o[931]) );
  AND U758 ( .A(p_input[9319]), .B(p_input[19319]), .Z(o[9319]) );
  AND U759 ( .A(p_input[9318]), .B(p_input[19318]), .Z(o[9318]) );
  AND U760 ( .A(p_input[9317]), .B(p_input[19317]), .Z(o[9317]) );
  AND U761 ( .A(p_input[9316]), .B(p_input[19316]), .Z(o[9316]) );
  AND U762 ( .A(p_input[9315]), .B(p_input[19315]), .Z(o[9315]) );
  AND U763 ( .A(p_input[9314]), .B(p_input[19314]), .Z(o[9314]) );
  AND U764 ( .A(p_input[9313]), .B(p_input[19313]), .Z(o[9313]) );
  AND U765 ( .A(p_input[9312]), .B(p_input[19312]), .Z(o[9312]) );
  AND U766 ( .A(p_input[9311]), .B(p_input[19311]), .Z(o[9311]) );
  AND U767 ( .A(p_input[9310]), .B(p_input[19310]), .Z(o[9310]) );
  AND U768 ( .A(p_input[930]), .B(p_input[10930]), .Z(o[930]) );
  AND U769 ( .A(p_input[9309]), .B(p_input[19309]), .Z(o[9309]) );
  AND U770 ( .A(p_input[9308]), .B(p_input[19308]), .Z(o[9308]) );
  AND U771 ( .A(p_input[9307]), .B(p_input[19307]), .Z(o[9307]) );
  AND U772 ( .A(p_input[9306]), .B(p_input[19306]), .Z(o[9306]) );
  AND U773 ( .A(p_input[9305]), .B(p_input[19305]), .Z(o[9305]) );
  AND U774 ( .A(p_input[9304]), .B(p_input[19304]), .Z(o[9304]) );
  AND U775 ( .A(p_input[9303]), .B(p_input[19303]), .Z(o[9303]) );
  AND U776 ( .A(p_input[9302]), .B(p_input[19302]), .Z(o[9302]) );
  AND U777 ( .A(p_input[9301]), .B(p_input[19301]), .Z(o[9301]) );
  AND U778 ( .A(p_input[9300]), .B(p_input[19300]), .Z(o[9300]) );
  AND U779 ( .A(p_input[92]), .B(p_input[10092]), .Z(o[92]) );
  AND U780 ( .A(p_input[929]), .B(p_input[10929]), .Z(o[929]) );
  AND U781 ( .A(p_input[9299]), .B(p_input[19299]), .Z(o[9299]) );
  AND U782 ( .A(p_input[9298]), .B(p_input[19298]), .Z(o[9298]) );
  AND U783 ( .A(p_input[9297]), .B(p_input[19297]), .Z(o[9297]) );
  AND U784 ( .A(p_input[9296]), .B(p_input[19296]), .Z(o[9296]) );
  AND U785 ( .A(p_input[9295]), .B(p_input[19295]), .Z(o[9295]) );
  AND U786 ( .A(p_input[9294]), .B(p_input[19294]), .Z(o[9294]) );
  AND U787 ( .A(p_input[9293]), .B(p_input[19293]), .Z(o[9293]) );
  AND U788 ( .A(p_input[9292]), .B(p_input[19292]), .Z(o[9292]) );
  AND U789 ( .A(p_input[9291]), .B(p_input[19291]), .Z(o[9291]) );
  AND U790 ( .A(p_input[9290]), .B(p_input[19290]), .Z(o[9290]) );
  AND U791 ( .A(p_input[928]), .B(p_input[10928]), .Z(o[928]) );
  AND U792 ( .A(p_input[9289]), .B(p_input[19289]), .Z(o[9289]) );
  AND U793 ( .A(p_input[9288]), .B(p_input[19288]), .Z(o[9288]) );
  AND U794 ( .A(p_input[9287]), .B(p_input[19287]), .Z(o[9287]) );
  AND U795 ( .A(p_input[9286]), .B(p_input[19286]), .Z(o[9286]) );
  AND U796 ( .A(p_input[9285]), .B(p_input[19285]), .Z(o[9285]) );
  AND U797 ( .A(p_input[9284]), .B(p_input[19284]), .Z(o[9284]) );
  AND U798 ( .A(p_input[9283]), .B(p_input[19283]), .Z(o[9283]) );
  AND U799 ( .A(p_input[9282]), .B(p_input[19282]), .Z(o[9282]) );
  AND U800 ( .A(p_input[9281]), .B(p_input[19281]), .Z(o[9281]) );
  AND U801 ( .A(p_input[9280]), .B(p_input[19280]), .Z(o[9280]) );
  AND U802 ( .A(p_input[927]), .B(p_input[10927]), .Z(o[927]) );
  AND U803 ( .A(p_input[9279]), .B(p_input[19279]), .Z(o[9279]) );
  AND U804 ( .A(p_input[9278]), .B(p_input[19278]), .Z(o[9278]) );
  AND U805 ( .A(p_input[9277]), .B(p_input[19277]), .Z(o[9277]) );
  AND U806 ( .A(p_input[9276]), .B(p_input[19276]), .Z(o[9276]) );
  AND U807 ( .A(p_input[9275]), .B(p_input[19275]), .Z(o[9275]) );
  AND U808 ( .A(p_input[9274]), .B(p_input[19274]), .Z(o[9274]) );
  AND U809 ( .A(p_input[9273]), .B(p_input[19273]), .Z(o[9273]) );
  AND U810 ( .A(p_input[9272]), .B(p_input[19272]), .Z(o[9272]) );
  AND U811 ( .A(p_input[9271]), .B(p_input[19271]), .Z(o[9271]) );
  AND U812 ( .A(p_input[9270]), .B(p_input[19270]), .Z(o[9270]) );
  AND U813 ( .A(p_input[926]), .B(p_input[10926]), .Z(o[926]) );
  AND U814 ( .A(p_input[9269]), .B(p_input[19269]), .Z(o[9269]) );
  AND U815 ( .A(p_input[9268]), .B(p_input[19268]), .Z(o[9268]) );
  AND U816 ( .A(p_input[9267]), .B(p_input[19267]), .Z(o[9267]) );
  AND U817 ( .A(p_input[9266]), .B(p_input[19266]), .Z(o[9266]) );
  AND U818 ( .A(p_input[9265]), .B(p_input[19265]), .Z(o[9265]) );
  AND U819 ( .A(p_input[9264]), .B(p_input[19264]), .Z(o[9264]) );
  AND U820 ( .A(p_input[9263]), .B(p_input[19263]), .Z(o[9263]) );
  AND U821 ( .A(p_input[9262]), .B(p_input[19262]), .Z(o[9262]) );
  AND U822 ( .A(p_input[9261]), .B(p_input[19261]), .Z(o[9261]) );
  AND U823 ( .A(p_input[9260]), .B(p_input[19260]), .Z(o[9260]) );
  AND U824 ( .A(p_input[925]), .B(p_input[10925]), .Z(o[925]) );
  AND U825 ( .A(p_input[9259]), .B(p_input[19259]), .Z(o[9259]) );
  AND U826 ( .A(p_input[9258]), .B(p_input[19258]), .Z(o[9258]) );
  AND U827 ( .A(p_input[9257]), .B(p_input[19257]), .Z(o[9257]) );
  AND U828 ( .A(p_input[9256]), .B(p_input[19256]), .Z(o[9256]) );
  AND U829 ( .A(p_input[9255]), .B(p_input[19255]), .Z(o[9255]) );
  AND U830 ( .A(p_input[9254]), .B(p_input[19254]), .Z(o[9254]) );
  AND U831 ( .A(p_input[9253]), .B(p_input[19253]), .Z(o[9253]) );
  AND U832 ( .A(p_input[9252]), .B(p_input[19252]), .Z(o[9252]) );
  AND U833 ( .A(p_input[9251]), .B(p_input[19251]), .Z(o[9251]) );
  AND U834 ( .A(p_input[9250]), .B(p_input[19250]), .Z(o[9250]) );
  AND U835 ( .A(p_input[924]), .B(p_input[10924]), .Z(o[924]) );
  AND U836 ( .A(p_input[9249]), .B(p_input[19249]), .Z(o[9249]) );
  AND U837 ( .A(p_input[9248]), .B(p_input[19248]), .Z(o[9248]) );
  AND U838 ( .A(p_input[9247]), .B(p_input[19247]), .Z(o[9247]) );
  AND U839 ( .A(p_input[9246]), .B(p_input[19246]), .Z(o[9246]) );
  AND U840 ( .A(p_input[9245]), .B(p_input[19245]), .Z(o[9245]) );
  AND U841 ( .A(p_input[9244]), .B(p_input[19244]), .Z(o[9244]) );
  AND U842 ( .A(p_input[9243]), .B(p_input[19243]), .Z(o[9243]) );
  AND U843 ( .A(p_input[9242]), .B(p_input[19242]), .Z(o[9242]) );
  AND U844 ( .A(p_input[9241]), .B(p_input[19241]), .Z(o[9241]) );
  AND U845 ( .A(p_input[9240]), .B(p_input[19240]), .Z(o[9240]) );
  AND U846 ( .A(p_input[923]), .B(p_input[10923]), .Z(o[923]) );
  AND U847 ( .A(p_input[9239]), .B(p_input[19239]), .Z(o[9239]) );
  AND U848 ( .A(p_input[9238]), .B(p_input[19238]), .Z(o[9238]) );
  AND U849 ( .A(p_input[9237]), .B(p_input[19237]), .Z(o[9237]) );
  AND U850 ( .A(p_input[9236]), .B(p_input[19236]), .Z(o[9236]) );
  AND U851 ( .A(p_input[9235]), .B(p_input[19235]), .Z(o[9235]) );
  AND U852 ( .A(p_input[9234]), .B(p_input[19234]), .Z(o[9234]) );
  AND U853 ( .A(p_input[9233]), .B(p_input[19233]), .Z(o[9233]) );
  AND U854 ( .A(p_input[9232]), .B(p_input[19232]), .Z(o[9232]) );
  AND U855 ( .A(p_input[9231]), .B(p_input[19231]), .Z(o[9231]) );
  AND U856 ( .A(p_input[9230]), .B(p_input[19230]), .Z(o[9230]) );
  AND U857 ( .A(p_input[922]), .B(p_input[10922]), .Z(o[922]) );
  AND U858 ( .A(p_input[9229]), .B(p_input[19229]), .Z(o[9229]) );
  AND U859 ( .A(p_input[9228]), .B(p_input[19228]), .Z(o[9228]) );
  AND U860 ( .A(p_input[9227]), .B(p_input[19227]), .Z(o[9227]) );
  AND U861 ( .A(p_input[9226]), .B(p_input[19226]), .Z(o[9226]) );
  AND U862 ( .A(p_input[9225]), .B(p_input[19225]), .Z(o[9225]) );
  AND U863 ( .A(p_input[9224]), .B(p_input[19224]), .Z(o[9224]) );
  AND U864 ( .A(p_input[9223]), .B(p_input[19223]), .Z(o[9223]) );
  AND U865 ( .A(p_input[9222]), .B(p_input[19222]), .Z(o[9222]) );
  AND U866 ( .A(p_input[9221]), .B(p_input[19221]), .Z(o[9221]) );
  AND U867 ( .A(p_input[9220]), .B(p_input[19220]), .Z(o[9220]) );
  AND U868 ( .A(p_input[921]), .B(p_input[10921]), .Z(o[921]) );
  AND U869 ( .A(p_input[9219]), .B(p_input[19219]), .Z(o[9219]) );
  AND U870 ( .A(p_input[9218]), .B(p_input[19218]), .Z(o[9218]) );
  AND U871 ( .A(p_input[9217]), .B(p_input[19217]), .Z(o[9217]) );
  AND U872 ( .A(p_input[9216]), .B(p_input[19216]), .Z(o[9216]) );
  AND U873 ( .A(p_input[9215]), .B(p_input[19215]), .Z(o[9215]) );
  AND U874 ( .A(p_input[9214]), .B(p_input[19214]), .Z(o[9214]) );
  AND U875 ( .A(p_input[9213]), .B(p_input[19213]), .Z(o[9213]) );
  AND U876 ( .A(p_input[9212]), .B(p_input[19212]), .Z(o[9212]) );
  AND U877 ( .A(p_input[9211]), .B(p_input[19211]), .Z(o[9211]) );
  AND U878 ( .A(p_input[9210]), .B(p_input[19210]), .Z(o[9210]) );
  AND U879 ( .A(p_input[920]), .B(p_input[10920]), .Z(o[920]) );
  AND U880 ( .A(p_input[9209]), .B(p_input[19209]), .Z(o[9209]) );
  AND U881 ( .A(p_input[9208]), .B(p_input[19208]), .Z(o[9208]) );
  AND U882 ( .A(p_input[9207]), .B(p_input[19207]), .Z(o[9207]) );
  AND U883 ( .A(p_input[9206]), .B(p_input[19206]), .Z(o[9206]) );
  AND U884 ( .A(p_input[9205]), .B(p_input[19205]), .Z(o[9205]) );
  AND U885 ( .A(p_input[9204]), .B(p_input[19204]), .Z(o[9204]) );
  AND U886 ( .A(p_input[9203]), .B(p_input[19203]), .Z(o[9203]) );
  AND U887 ( .A(p_input[9202]), .B(p_input[19202]), .Z(o[9202]) );
  AND U888 ( .A(p_input[9201]), .B(p_input[19201]), .Z(o[9201]) );
  AND U889 ( .A(p_input[9200]), .B(p_input[19200]), .Z(o[9200]) );
  AND U890 ( .A(p_input[91]), .B(p_input[10091]), .Z(o[91]) );
  AND U891 ( .A(p_input[919]), .B(p_input[10919]), .Z(o[919]) );
  AND U892 ( .A(p_input[9199]), .B(p_input[19199]), .Z(o[9199]) );
  AND U893 ( .A(p_input[9198]), .B(p_input[19198]), .Z(o[9198]) );
  AND U894 ( .A(p_input[9197]), .B(p_input[19197]), .Z(o[9197]) );
  AND U895 ( .A(p_input[9196]), .B(p_input[19196]), .Z(o[9196]) );
  AND U896 ( .A(p_input[9195]), .B(p_input[19195]), .Z(o[9195]) );
  AND U897 ( .A(p_input[9194]), .B(p_input[19194]), .Z(o[9194]) );
  AND U898 ( .A(p_input[9193]), .B(p_input[19193]), .Z(o[9193]) );
  AND U899 ( .A(p_input[9192]), .B(p_input[19192]), .Z(o[9192]) );
  AND U900 ( .A(p_input[9191]), .B(p_input[19191]), .Z(o[9191]) );
  AND U901 ( .A(p_input[9190]), .B(p_input[19190]), .Z(o[9190]) );
  AND U902 ( .A(p_input[918]), .B(p_input[10918]), .Z(o[918]) );
  AND U903 ( .A(p_input[9189]), .B(p_input[19189]), .Z(o[9189]) );
  AND U904 ( .A(p_input[9188]), .B(p_input[19188]), .Z(o[9188]) );
  AND U905 ( .A(p_input[9187]), .B(p_input[19187]), .Z(o[9187]) );
  AND U906 ( .A(p_input[9186]), .B(p_input[19186]), .Z(o[9186]) );
  AND U907 ( .A(p_input[9185]), .B(p_input[19185]), .Z(o[9185]) );
  AND U908 ( .A(p_input[9184]), .B(p_input[19184]), .Z(o[9184]) );
  AND U909 ( .A(p_input[9183]), .B(p_input[19183]), .Z(o[9183]) );
  AND U910 ( .A(p_input[9182]), .B(p_input[19182]), .Z(o[9182]) );
  AND U911 ( .A(p_input[9181]), .B(p_input[19181]), .Z(o[9181]) );
  AND U912 ( .A(p_input[9180]), .B(p_input[19180]), .Z(o[9180]) );
  AND U913 ( .A(p_input[917]), .B(p_input[10917]), .Z(o[917]) );
  AND U914 ( .A(p_input[9179]), .B(p_input[19179]), .Z(o[9179]) );
  AND U915 ( .A(p_input[9178]), .B(p_input[19178]), .Z(o[9178]) );
  AND U916 ( .A(p_input[9177]), .B(p_input[19177]), .Z(o[9177]) );
  AND U917 ( .A(p_input[9176]), .B(p_input[19176]), .Z(o[9176]) );
  AND U918 ( .A(p_input[9175]), .B(p_input[19175]), .Z(o[9175]) );
  AND U919 ( .A(p_input[9174]), .B(p_input[19174]), .Z(o[9174]) );
  AND U920 ( .A(p_input[9173]), .B(p_input[19173]), .Z(o[9173]) );
  AND U921 ( .A(p_input[9172]), .B(p_input[19172]), .Z(o[9172]) );
  AND U922 ( .A(p_input[9171]), .B(p_input[19171]), .Z(o[9171]) );
  AND U923 ( .A(p_input[9170]), .B(p_input[19170]), .Z(o[9170]) );
  AND U924 ( .A(p_input[916]), .B(p_input[10916]), .Z(o[916]) );
  AND U925 ( .A(p_input[9169]), .B(p_input[19169]), .Z(o[9169]) );
  AND U926 ( .A(p_input[9168]), .B(p_input[19168]), .Z(o[9168]) );
  AND U927 ( .A(p_input[9167]), .B(p_input[19167]), .Z(o[9167]) );
  AND U928 ( .A(p_input[9166]), .B(p_input[19166]), .Z(o[9166]) );
  AND U929 ( .A(p_input[9165]), .B(p_input[19165]), .Z(o[9165]) );
  AND U930 ( .A(p_input[9164]), .B(p_input[19164]), .Z(o[9164]) );
  AND U931 ( .A(p_input[9163]), .B(p_input[19163]), .Z(o[9163]) );
  AND U932 ( .A(p_input[9162]), .B(p_input[19162]), .Z(o[9162]) );
  AND U933 ( .A(p_input[9161]), .B(p_input[19161]), .Z(o[9161]) );
  AND U934 ( .A(p_input[9160]), .B(p_input[19160]), .Z(o[9160]) );
  AND U935 ( .A(p_input[915]), .B(p_input[10915]), .Z(o[915]) );
  AND U936 ( .A(p_input[9159]), .B(p_input[19159]), .Z(o[9159]) );
  AND U937 ( .A(p_input[9158]), .B(p_input[19158]), .Z(o[9158]) );
  AND U938 ( .A(p_input[9157]), .B(p_input[19157]), .Z(o[9157]) );
  AND U939 ( .A(p_input[9156]), .B(p_input[19156]), .Z(o[9156]) );
  AND U940 ( .A(p_input[9155]), .B(p_input[19155]), .Z(o[9155]) );
  AND U941 ( .A(p_input[9154]), .B(p_input[19154]), .Z(o[9154]) );
  AND U942 ( .A(p_input[9153]), .B(p_input[19153]), .Z(o[9153]) );
  AND U943 ( .A(p_input[9152]), .B(p_input[19152]), .Z(o[9152]) );
  AND U944 ( .A(p_input[9151]), .B(p_input[19151]), .Z(o[9151]) );
  AND U945 ( .A(p_input[9150]), .B(p_input[19150]), .Z(o[9150]) );
  AND U946 ( .A(p_input[914]), .B(p_input[10914]), .Z(o[914]) );
  AND U947 ( .A(p_input[9149]), .B(p_input[19149]), .Z(o[9149]) );
  AND U948 ( .A(p_input[9148]), .B(p_input[19148]), .Z(o[9148]) );
  AND U949 ( .A(p_input[9147]), .B(p_input[19147]), .Z(o[9147]) );
  AND U950 ( .A(p_input[9146]), .B(p_input[19146]), .Z(o[9146]) );
  AND U951 ( .A(p_input[9145]), .B(p_input[19145]), .Z(o[9145]) );
  AND U952 ( .A(p_input[9144]), .B(p_input[19144]), .Z(o[9144]) );
  AND U953 ( .A(p_input[9143]), .B(p_input[19143]), .Z(o[9143]) );
  AND U954 ( .A(p_input[9142]), .B(p_input[19142]), .Z(o[9142]) );
  AND U955 ( .A(p_input[9141]), .B(p_input[19141]), .Z(o[9141]) );
  AND U956 ( .A(p_input[9140]), .B(p_input[19140]), .Z(o[9140]) );
  AND U957 ( .A(p_input[913]), .B(p_input[10913]), .Z(o[913]) );
  AND U958 ( .A(p_input[9139]), .B(p_input[19139]), .Z(o[9139]) );
  AND U959 ( .A(p_input[9138]), .B(p_input[19138]), .Z(o[9138]) );
  AND U960 ( .A(p_input[9137]), .B(p_input[19137]), .Z(o[9137]) );
  AND U961 ( .A(p_input[9136]), .B(p_input[19136]), .Z(o[9136]) );
  AND U962 ( .A(p_input[9135]), .B(p_input[19135]), .Z(o[9135]) );
  AND U963 ( .A(p_input[9134]), .B(p_input[19134]), .Z(o[9134]) );
  AND U964 ( .A(p_input[9133]), .B(p_input[19133]), .Z(o[9133]) );
  AND U965 ( .A(p_input[9132]), .B(p_input[19132]), .Z(o[9132]) );
  AND U966 ( .A(p_input[9131]), .B(p_input[19131]), .Z(o[9131]) );
  AND U967 ( .A(p_input[9130]), .B(p_input[19130]), .Z(o[9130]) );
  AND U968 ( .A(p_input[912]), .B(p_input[10912]), .Z(o[912]) );
  AND U969 ( .A(p_input[9129]), .B(p_input[19129]), .Z(o[9129]) );
  AND U970 ( .A(p_input[9128]), .B(p_input[19128]), .Z(o[9128]) );
  AND U971 ( .A(p_input[9127]), .B(p_input[19127]), .Z(o[9127]) );
  AND U972 ( .A(p_input[9126]), .B(p_input[19126]), .Z(o[9126]) );
  AND U973 ( .A(p_input[9125]), .B(p_input[19125]), .Z(o[9125]) );
  AND U974 ( .A(p_input[9124]), .B(p_input[19124]), .Z(o[9124]) );
  AND U975 ( .A(p_input[9123]), .B(p_input[19123]), .Z(o[9123]) );
  AND U976 ( .A(p_input[9122]), .B(p_input[19122]), .Z(o[9122]) );
  AND U977 ( .A(p_input[9121]), .B(p_input[19121]), .Z(o[9121]) );
  AND U978 ( .A(p_input[9120]), .B(p_input[19120]), .Z(o[9120]) );
  AND U979 ( .A(p_input[911]), .B(p_input[10911]), .Z(o[911]) );
  AND U980 ( .A(p_input[9119]), .B(p_input[19119]), .Z(o[9119]) );
  AND U981 ( .A(p_input[9118]), .B(p_input[19118]), .Z(o[9118]) );
  AND U982 ( .A(p_input[9117]), .B(p_input[19117]), .Z(o[9117]) );
  AND U983 ( .A(p_input[9116]), .B(p_input[19116]), .Z(o[9116]) );
  AND U984 ( .A(p_input[9115]), .B(p_input[19115]), .Z(o[9115]) );
  AND U985 ( .A(p_input[9114]), .B(p_input[19114]), .Z(o[9114]) );
  AND U986 ( .A(p_input[9113]), .B(p_input[19113]), .Z(o[9113]) );
  AND U987 ( .A(p_input[9112]), .B(p_input[19112]), .Z(o[9112]) );
  AND U988 ( .A(p_input[9111]), .B(p_input[19111]), .Z(o[9111]) );
  AND U989 ( .A(p_input[9110]), .B(p_input[19110]), .Z(o[9110]) );
  AND U990 ( .A(p_input[910]), .B(p_input[10910]), .Z(o[910]) );
  AND U991 ( .A(p_input[9109]), .B(p_input[19109]), .Z(o[9109]) );
  AND U992 ( .A(p_input[9108]), .B(p_input[19108]), .Z(o[9108]) );
  AND U993 ( .A(p_input[9107]), .B(p_input[19107]), .Z(o[9107]) );
  AND U994 ( .A(p_input[9106]), .B(p_input[19106]), .Z(o[9106]) );
  AND U995 ( .A(p_input[9105]), .B(p_input[19105]), .Z(o[9105]) );
  AND U996 ( .A(p_input[9104]), .B(p_input[19104]), .Z(o[9104]) );
  AND U997 ( .A(p_input[9103]), .B(p_input[19103]), .Z(o[9103]) );
  AND U998 ( .A(p_input[9102]), .B(p_input[19102]), .Z(o[9102]) );
  AND U999 ( .A(p_input[9101]), .B(p_input[19101]), .Z(o[9101]) );
  AND U1000 ( .A(p_input[9100]), .B(p_input[19100]), .Z(o[9100]) );
  AND U1001 ( .A(p_input[90]), .B(p_input[10090]), .Z(o[90]) );
  AND U1002 ( .A(p_input[909]), .B(p_input[10909]), .Z(o[909]) );
  AND U1003 ( .A(p_input[9099]), .B(p_input[19099]), .Z(o[9099]) );
  AND U1004 ( .A(p_input[9098]), .B(p_input[19098]), .Z(o[9098]) );
  AND U1005 ( .A(p_input[9097]), .B(p_input[19097]), .Z(o[9097]) );
  AND U1006 ( .A(p_input[9096]), .B(p_input[19096]), .Z(o[9096]) );
  AND U1007 ( .A(p_input[9095]), .B(p_input[19095]), .Z(o[9095]) );
  AND U1008 ( .A(p_input[9094]), .B(p_input[19094]), .Z(o[9094]) );
  AND U1009 ( .A(p_input[9093]), .B(p_input[19093]), .Z(o[9093]) );
  AND U1010 ( .A(p_input[9092]), .B(p_input[19092]), .Z(o[9092]) );
  AND U1011 ( .A(p_input[9091]), .B(p_input[19091]), .Z(o[9091]) );
  AND U1012 ( .A(p_input[9090]), .B(p_input[19090]), .Z(o[9090]) );
  AND U1013 ( .A(p_input[908]), .B(p_input[10908]), .Z(o[908]) );
  AND U1014 ( .A(p_input[9089]), .B(p_input[19089]), .Z(o[9089]) );
  AND U1015 ( .A(p_input[9088]), .B(p_input[19088]), .Z(o[9088]) );
  AND U1016 ( .A(p_input[9087]), .B(p_input[19087]), .Z(o[9087]) );
  AND U1017 ( .A(p_input[9086]), .B(p_input[19086]), .Z(o[9086]) );
  AND U1018 ( .A(p_input[9085]), .B(p_input[19085]), .Z(o[9085]) );
  AND U1019 ( .A(p_input[9084]), .B(p_input[19084]), .Z(o[9084]) );
  AND U1020 ( .A(p_input[9083]), .B(p_input[19083]), .Z(o[9083]) );
  AND U1021 ( .A(p_input[9082]), .B(p_input[19082]), .Z(o[9082]) );
  AND U1022 ( .A(p_input[9081]), .B(p_input[19081]), .Z(o[9081]) );
  AND U1023 ( .A(p_input[9080]), .B(p_input[19080]), .Z(o[9080]) );
  AND U1024 ( .A(p_input[907]), .B(p_input[10907]), .Z(o[907]) );
  AND U1025 ( .A(p_input[9079]), .B(p_input[19079]), .Z(o[9079]) );
  AND U1026 ( .A(p_input[9078]), .B(p_input[19078]), .Z(o[9078]) );
  AND U1027 ( .A(p_input[9077]), .B(p_input[19077]), .Z(o[9077]) );
  AND U1028 ( .A(p_input[9076]), .B(p_input[19076]), .Z(o[9076]) );
  AND U1029 ( .A(p_input[9075]), .B(p_input[19075]), .Z(o[9075]) );
  AND U1030 ( .A(p_input[9074]), .B(p_input[19074]), .Z(o[9074]) );
  AND U1031 ( .A(p_input[9073]), .B(p_input[19073]), .Z(o[9073]) );
  AND U1032 ( .A(p_input[9072]), .B(p_input[19072]), .Z(o[9072]) );
  AND U1033 ( .A(p_input[9071]), .B(p_input[19071]), .Z(o[9071]) );
  AND U1034 ( .A(p_input[9070]), .B(p_input[19070]), .Z(o[9070]) );
  AND U1035 ( .A(p_input[906]), .B(p_input[10906]), .Z(o[906]) );
  AND U1036 ( .A(p_input[9069]), .B(p_input[19069]), .Z(o[9069]) );
  AND U1037 ( .A(p_input[9068]), .B(p_input[19068]), .Z(o[9068]) );
  AND U1038 ( .A(p_input[9067]), .B(p_input[19067]), .Z(o[9067]) );
  AND U1039 ( .A(p_input[9066]), .B(p_input[19066]), .Z(o[9066]) );
  AND U1040 ( .A(p_input[9065]), .B(p_input[19065]), .Z(o[9065]) );
  AND U1041 ( .A(p_input[9064]), .B(p_input[19064]), .Z(o[9064]) );
  AND U1042 ( .A(p_input[9063]), .B(p_input[19063]), .Z(o[9063]) );
  AND U1043 ( .A(p_input[9062]), .B(p_input[19062]), .Z(o[9062]) );
  AND U1044 ( .A(p_input[9061]), .B(p_input[19061]), .Z(o[9061]) );
  AND U1045 ( .A(p_input[9060]), .B(p_input[19060]), .Z(o[9060]) );
  AND U1046 ( .A(p_input[905]), .B(p_input[10905]), .Z(o[905]) );
  AND U1047 ( .A(p_input[9059]), .B(p_input[19059]), .Z(o[9059]) );
  AND U1048 ( .A(p_input[9058]), .B(p_input[19058]), .Z(o[9058]) );
  AND U1049 ( .A(p_input[9057]), .B(p_input[19057]), .Z(o[9057]) );
  AND U1050 ( .A(p_input[9056]), .B(p_input[19056]), .Z(o[9056]) );
  AND U1051 ( .A(p_input[9055]), .B(p_input[19055]), .Z(o[9055]) );
  AND U1052 ( .A(p_input[9054]), .B(p_input[19054]), .Z(o[9054]) );
  AND U1053 ( .A(p_input[9053]), .B(p_input[19053]), .Z(o[9053]) );
  AND U1054 ( .A(p_input[9052]), .B(p_input[19052]), .Z(o[9052]) );
  AND U1055 ( .A(p_input[9051]), .B(p_input[19051]), .Z(o[9051]) );
  AND U1056 ( .A(p_input[9050]), .B(p_input[19050]), .Z(o[9050]) );
  AND U1057 ( .A(p_input[904]), .B(p_input[10904]), .Z(o[904]) );
  AND U1058 ( .A(p_input[9049]), .B(p_input[19049]), .Z(o[9049]) );
  AND U1059 ( .A(p_input[9048]), .B(p_input[19048]), .Z(o[9048]) );
  AND U1060 ( .A(p_input[9047]), .B(p_input[19047]), .Z(o[9047]) );
  AND U1061 ( .A(p_input[9046]), .B(p_input[19046]), .Z(o[9046]) );
  AND U1062 ( .A(p_input[9045]), .B(p_input[19045]), .Z(o[9045]) );
  AND U1063 ( .A(p_input[9044]), .B(p_input[19044]), .Z(o[9044]) );
  AND U1064 ( .A(p_input[9043]), .B(p_input[19043]), .Z(o[9043]) );
  AND U1065 ( .A(p_input[9042]), .B(p_input[19042]), .Z(o[9042]) );
  AND U1066 ( .A(p_input[9041]), .B(p_input[19041]), .Z(o[9041]) );
  AND U1067 ( .A(p_input[9040]), .B(p_input[19040]), .Z(o[9040]) );
  AND U1068 ( .A(p_input[903]), .B(p_input[10903]), .Z(o[903]) );
  AND U1069 ( .A(p_input[9039]), .B(p_input[19039]), .Z(o[9039]) );
  AND U1070 ( .A(p_input[9038]), .B(p_input[19038]), .Z(o[9038]) );
  AND U1071 ( .A(p_input[9037]), .B(p_input[19037]), .Z(o[9037]) );
  AND U1072 ( .A(p_input[9036]), .B(p_input[19036]), .Z(o[9036]) );
  AND U1073 ( .A(p_input[9035]), .B(p_input[19035]), .Z(o[9035]) );
  AND U1074 ( .A(p_input[9034]), .B(p_input[19034]), .Z(o[9034]) );
  AND U1075 ( .A(p_input[9033]), .B(p_input[19033]), .Z(o[9033]) );
  AND U1076 ( .A(p_input[9032]), .B(p_input[19032]), .Z(o[9032]) );
  AND U1077 ( .A(p_input[9031]), .B(p_input[19031]), .Z(o[9031]) );
  AND U1078 ( .A(p_input[9030]), .B(p_input[19030]), .Z(o[9030]) );
  AND U1079 ( .A(p_input[902]), .B(p_input[10902]), .Z(o[902]) );
  AND U1080 ( .A(p_input[9029]), .B(p_input[19029]), .Z(o[9029]) );
  AND U1081 ( .A(p_input[9028]), .B(p_input[19028]), .Z(o[9028]) );
  AND U1082 ( .A(p_input[9027]), .B(p_input[19027]), .Z(o[9027]) );
  AND U1083 ( .A(p_input[9026]), .B(p_input[19026]), .Z(o[9026]) );
  AND U1084 ( .A(p_input[9025]), .B(p_input[19025]), .Z(o[9025]) );
  AND U1085 ( .A(p_input[9024]), .B(p_input[19024]), .Z(o[9024]) );
  AND U1086 ( .A(p_input[9023]), .B(p_input[19023]), .Z(o[9023]) );
  AND U1087 ( .A(p_input[9022]), .B(p_input[19022]), .Z(o[9022]) );
  AND U1088 ( .A(p_input[9021]), .B(p_input[19021]), .Z(o[9021]) );
  AND U1089 ( .A(p_input[9020]), .B(p_input[19020]), .Z(o[9020]) );
  AND U1090 ( .A(p_input[901]), .B(p_input[10901]), .Z(o[901]) );
  AND U1091 ( .A(p_input[9019]), .B(p_input[19019]), .Z(o[9019]) );
  AND U1092 ( .A(p_input[9018]), .B(p_input[19018]), .Z(o[9018]) );
  AND U1093 ( .A(p_input[9017]), .B(p_input[19017]), .Z(o[9017]) );
  AND U1094 ( .A(p_input[9016]), .B(p_input[19016]), .Z(o[9016]) );
  AND U1095 ( .A(p_input[9015]), .B(p_input[19015]), .Z(o[9015]) );
  AND U1096 ( .A(p_input[9014]), .B(p_input[19014]), .Z(o[9014]) );
  AND U1097 ( .A(p_input[9013]), .B(p_input[19013]), .Z(o[9013]) );
  AND U1098 ( .A(p_input[9012]), .B(p_input[19012]), .Z(o[9012]) );
  AND U1099 ( .A(p_input[9011]), .B(p_input[19011]), .Z(o[9011]) );
  AND U1100 ( .A(p_input[9010]), .B(p_input[19010]), .Z(o[9010]) );
  AND U1101 ( .A(p_input[900]), .B(p_input[10900]), .Z(o[900]) );
  AND U1102 ( .A(p_input[9009]), .B(p_input[19009]), .Z(o[9009]) );
  AND U1103 ( .A(p_input[9008]), .B(p_input[19008]), .Z(o[9008]) );
  AND U1104 ( .A(p_input[9007]), .B(p_input[19007]), .Z(o[9007]) );
  AND U1105 ( .A(p_input[9006]), .B(p_input[19006]), .Z(o[9006]) );
  AND U1106 ( .A(p_input[9005]), .B(p_input[19005]), .Z(o[9005]) );
  AND U1107 ( .A(p_input[9004]), .B(p_input[19004]), .Z(o[9004]) );
  AND U1108 ( .A(p_input[9003]), .B(p_input[19003]), .Z(o[9003]) );
  AND U1109 ( .A(p_input[9002]), .B(p_input[19002]), .Z(o[9002]) );
  AND U1110 ( .A(p_input[9001]), .B(p_input[19001]), .Z(o[9001]) );
  AND U1111 ( .A(p_input[9000]), .B(p_input[19000]), .Z(o[9000]) );
  AND U1112 ( .A(p_input[8]), .B(p_input[10008]), .Z(o[8]) );
  AND U1113 ( .A(p_input[89]), .B(p_input[10089]), .Z(o[89]) );
  AND U1114 ( .A(p_input[899]), .B(p_input[10899]), .Z(o[899]) );
  AND U1115 ( .A(p_input[8999]), .B(p_input[18999]), .Z(o[8999]) );
  AND U1116 ( .A(p_input[8998]), .B(p_input[18998]), .Z(o[8998]) );
  AND U1117 ( .A(p_input[8997]), .B(p_input[18997]), .Z(o[8997]) );
  AND U1118 ( .A(p_input[8996]), .B(p_input[18996]), .Z(o[8996]) );
  AND U1119 ( .A(p_input[8995]), .B(p_input[18995]), .Z(o[8995]) );
  AND U1120 ( .A(p_input[8994]), .B(p_input[18994]), .Z(o[8994]) );
  AND U1121 ( .A(p_input[8993]), .B(p_input[18993]), .Z(o[8993]) );
  AND U1122 ( .A(p_input[8992]), .B(p_input[18992]), .Z(o[8992]) );
  AND U1123 ( .A(p_input[8991]), .B(p_input[18991]), .Z(o[8991]) );
  AND U1124 ( .A(p_input[8990]), .B(p_input[18990]), .Z(o[8990]) );
  AND U1125 ( .A(p_input[898]), .B(p_input[10898]), .Z(o[898]) );
  AND U1126 ( .A(p_input[8989]), .B(p_input[18989]), .Z(o[8989]) );
  AND U1127 ( .A(p_input[8988]), .B(p_input[18988]), .Z(o[8988]) );
  AND U1128 ( .A(p_input[8987]), .B(p_input[18987]), .Z(o[8987]) );
  AND U1129 ( .A(p_input[8986]), .B(p_input[18986]), .Z(o[8986]) );
  AND U1130 ( .A(p_input[8985]), .B(p_input[18985]), .Z(o[8985]) );
  AND U1131 ( .A(p_input[8984]), .B(p_input[18984]), .Z(o[8984]) );
  AND U1132 ( .A(p_input[8983]), .B(p_input[18983]), .Z(o[8983]) );
  AND U1133 ( .A(p_input[8982]), .B(p_input[18982]), .Z(o[8982]) );
  AND U1134 ( .A(p_input[8981]), .B(p_input[18981]), .Z(o[8981]) );
  AND U1135 ( .A(p_input[8980]), .B(p_input[18980]), .Z(o[8980]) );
  AND U1136 ( .A(p_input[897]), .B(p_input[10897]), .Z(o[897]) );
  AND U1137 ( .A(p_input[8979]), .B(p_input[18979]), .Z(o[8979]) );
  AND U1138 ( .A(p_input[8978]), .B(p_input[18978]), .Z(o[8978]) );
  AND U1139 ( .A(p_input[8977]), .B(p_input[18977]), .Z(o[8977]) );
  AND U1140 ( .A(p_input[8976]), .B(p_input[18976]), .Z(o[8976]) );
  AND U1141 ( .A(p_input[8975]), .B(p_input[18975]), .Z(o[8975]) );
  AND U1142 ( .A(p_input[8974]), .B(p_input[18974]), .Z(o[8974]) );
  AND U1143 ( .A(p_input[8973]), .B(p_input[18973]), .Z(o[8973]) );
  AND U1144 ( .A(p_input[8972]), .B(p_input[18972]), .Z(o[8972]) );
  AND U1145 ( .A(p_input[8971]), .B(p_input[18971]), .Z(o[8971]) );
  AND U1146 ( .A(p_input[8970]), .B(p_input[18970]), .Z(o[8970]) );
  AND U1147 ( .A(p_input[896]), .B(p_input[10896]), .Z(o[896]) );
  AND U1148 ( .A(p_input[8969]), .B(p_input[18969]), .Z(o[8969]) );
  AND U1149 ( .A(p_input[8968]), .B(p_input[18968]), .Z(o[8968]) );
  AND U1150 ( .A(p_input[8967]), .B(p_input[18967]), .Z(o[8967]) );
  AND U1151 ( .A(p_input[8966]), .B(p_input[18966]), .Z(o[8966]) );
  AND U1152 ( .A(p_input[8965]), .B(p_input[18965]), .Z(o[8965]) );
  AND U1153 ( .A(p_input[8964]), .B(p_input[18964]), .Z(o[8964]) );
  AND U1154 ( .A(p_input[8963]), .B(p_input[18963]), .Z(o[8963]) );
  AND U1155 ( .A(p_input[8962]), .B(p_input[18962]), .Z(o[8962]) );
  AND U1156 ( .A(p_input[8961]), .B(p_input[18961]), .Z(o[8961]) );
  AND U1157 ( .A(p_input[8960]), .B(p_input[18960]), .Z(o[8960]) );
  AND U1158 ( .A(p_input[895]), .B(p_input[10895]), .Z(o[895]) );
  AND U1159 ( .A(p_input[8959]), .B(p_input[18959]), .Z(o[8959]) );
  AND U1160 ( .A(p_input[8958]), .B(p_input[18958]), .Z(o[8958]) );
  AND U1161 ( .A(p_input[8957]), .B(p_input[18957]), .Z(o[8957]) );
  AND U1162 ( .A(p_input[8956]), .B(p_input[18956]), .Z(o[8956]) );
  AND U1163 ( .A(p_input[8955]), .B(p_input[18955]), .Z(o[8955]) );
  AND U1164 ( .A(p_input[8954]), .B(p_input[18954]), .Z(o[8954]) );
  AND U1165 ( .A(p_input[8953]), .B(p_input[18953]), .Z(o[8953]) );
  AND U1166 ( .A(p_input[8952]), .B(p_input[18952]), .Z(o[8952]) );
  AND U1167 ( .A(p_input[8951]), .B(p_input[18951]), .Z(o[8951]) );
  AND U1168 ( .A(p_input[8950]), .B(p_input[18950]), .Z(o[8950]) );
  AND U1169 ( .A(p_input[894]), .B(p_input[10894]), .Z(o[894]) );
  AND U1170 ( .A(p_input[8949]), .B(p_input[18949]), .Z(o[8949]) );
  AND U1171 ( .A(p_input[8948]), .B(p_input[18948]), .Z(o[8948]) );
  AND U1172 ( .A(p_input[8947]), .B(p_input[18947]), .Z(o[8947]) );
  AND U1173 ( .A(p_input[8946]), .B(p_input[18946]), .Z(o[8946]) );
  AND U1174 ( .A(p_input[8945]), .B(p_input[18945]), .Z(o[8945]) );
  AND U1175 ( .A(p_input[8944]), .B(p_input[18944]), .Z(o[8944]) );
  AND U1176 ( .A(p_input[8943]), .B(p_input[18943]), .Z(o[8943]) );
  AND U1177 ( .A(p_input[8942]), .B(p_input[18942]), .Z(o[8942]) );
  AND U1178 ( .A(p_input[8941]), .B(p_input[18941]), .Z(o[8941]) );
  AND U1179 ( .A(p_input[8940]), .B(p_input[18940]), .Z(o[8940]) );
  AND U1180 ( .A(p_input[893]), .B(p_input[10893]), .Z(o[893]) );
  AND U1181 ( .A(p_input[8939]), .B(p_input[18939]), .Z(o[8939]) );
  AND U1182 ( .A(p_input[8938]), .B(p_input[18938]), .Z(o[8938]) );
  AND U1183 ( .A(p_input[8937]), .B(p_input[18937]), .Z(o[8937]) );
  AND U1184 ( .A(p_input[8936]), .B(p_input[18936]), .Z(o[8936]) );
  AND U1185 ( .A(p_input[8935]), .B(p_input[18935]), .Z(o[8935]) );
  AND U1186 ( .A(p_input[8934]), .B(p_input[18934]), .Z(o[8934]) );
  AND U1187 ( .A(p_input[8933]), .B(p_input[18933]), .Z(o[8933]) );
  AND U1188 ( .A(p_input[8932]), .B(p_input[18932]), .Z(o[8932]) );
  AND U1189 ( .A(p_input[8931]), .B(p_input[18931]), .Z(o[8931]) );
  AND U1190 ( .A(p_input[8930]), .B(p_input[18930]), .Z(o[8930]) );
  AND U1191 ( .A(p_input[892]), .B(p_input[10892]), .Z(o[892]) );
  AND U1192 ( .A(p_input[8929]), .B(p_input[18929]), .Z(o[8929]) );
  AND U1193 ( .A(p_input[8928]), .B(p_input[18928]), .Z(o[8928]) );
  AND U1194 ( .A(p_input[8927]), .B(p_input[18927]), .Z(o[8927]) );
  AND U1195 ( .A(p_input[8926]), .B(p_input[18926]), .Z(o[8926]) );
  AND U1196 ( .A(p_input[8925]), .B(p_input[18925]), .Z(o[8925]) );
  AND U1197 ( .A(p_input[8924]), .B(p_input[18924]), .Z(o[8924]) );
  AND U1198 ( .A(p_input[8923]), .B(p_input[18923]), .Z(o[8923]) );
  AND U1199 ( .A(p_input[8922]), .B(p_input[18922]), .Z(o[8922]) );
  AND U1200 ( .A(p_input[8921]), .B(p_input[18921]), .Z(o[8921]) );
  AND U1201 ( .A(p_input[8920]), .B(p_input[18920]), .Z(o[8920]) );
  AND U1202 ( .A(p_input[891]), .B(p_input[10891]), .Z(o[891]) );
  AND U1203 ( .A(p_input[8919]), .B(p_input[18919]), .Z(o[8919]) );
  AND U1204 ( .A(p_input[8918]), .B(p_input[18918]), .Z(o[8918]) );
  AND U1205 ( .A(p_input[8917]), .B(p_input[18917]), .Z(o[8917]) );
  AND U1206 ( .A(p_input[8916]), .B(p_input[18916]), .Z(o[8916]) );
  AND U1207 ( .A(p_input[8915]), .B(p_input[18915]), .Z(o[8915]) );
  AND U1208 ( .A(p_input[8914]), .B(p_input[18914]), .Z(o[8914]) );
  AND U1209 ( .A(p_input[8913]), .B(p_input[18913]), .Z(o[8913]) );
  AND U1210 ( .A(p_input[8912]), .B(p_input[18912]), .Z(o[8912]) );
  AND U1211 ( .A(p_input[8911]), .B(p_input[18911]), .Z(o[8911]) );
  AND U1212 ( .A(p_input[8910]), .B(p_input[18910]), .Z(o[8910]) );
  AND U1213 ( .A(p_input[890]), .B(p_input[10890]), .Z(o[890]) );
  AND U1214 ( .A(p_input[8909]), .B(p_input[18909]), .Z(o[8909]) );
  AND U1215 ( .A(p_input[8908]), .B(p_input[18908]), .Z(o[8908]) );
  AND U1216 ( .A(p_input[8907]), .B(p_input[18907]), .Z(o[8907]) );
  AND U1217 ( .A(p_input[8906]), .B(p_input[18906]), .Z(o[8906]) );
  AND U1218 ( .A(p_input[8905]), .B(p_input[18905]), .Z(o[8905]) );
  AND U1219 ( .A(p_input[8904]), .B(p_input[18904]), .Z(o[8904]) );
  AND U1220 ( .A(p_input[8903]), .B(p_input[18903]), .Z(o[8903]) );
  AND U1221 ( .A(p_input[8902]), .B(p_input[18902]), .Z(o[8902]) );
  AND U1222 ( .A(p_input[8901]), .B(p_input[18901]), .Z(o[8901]) );
  AND U1223 ( .A(p_input[8900]), .B(p_input[18900]), .Z(o[8900]) );
  AND U1224 ( .A(p_input[88]), .B(p_input[10088]), .Z(o[88]) );
  AND U1225 ( .A(p_input[889]), .B(p_input[10889]), .Z(o[889]) );
  AND U1226 ( .A(p_input[8899]), .B(p_input[18899]), .Z(o[8899]) );
  AND U1227 ( .A(p_input[8898]), .B(p_input[18898]), .Z(o[8898]) );
  AND U1228 ( .A(p_input[8897]), .B(p_input[18897]), .Z(o[8897]) );
  AND U1229 ( .A(p_input[8896]), .B(p_input[18896]), .Z(o[8896]) );
  AND U1230 ( .A(p_input[8895]), .B(p_input[18895]), .Z(o[8895]) );
  AND U1231 ( .A(p_input[8894]), .B(p_input[18894]), .Z(o[8894]) );
  AND U1232 ( .A(p_input[8893]), .B(p_input[18893]), .Z(o[8893]) );
  AND U1233 ( .A(p_input[8892]), .B(p_input[18892]), .Z(o[8892]) );
  AND U1234 ( .A(p_input[8891]), .B(p_input[18891]), .Z(o[8891]) );
  AND U1235 ( .A(p_input[8890]), .B(p_input[18890]), .Z(o[8890]) );
  AND U1236 ( .A(p_input[888]), .B(p_input[10888]), .Z(o[888]) );
  AND U1237 ( .A(p_input[8889]), .B(p_input[18889]), .Z(o[8889]) );
  AND U1238 ( .A(p_input[8888]), .B(p_input[18888]), .Z(o[8888]) );
  AND U1239 ( .A(p_input[8887]), .B(p_input[18887]), .Z(o[8887]) );
  AND U1240 ( .A(p_input[8886]), .B(p_input[18886]), .Z(o[8886]) );
  AND U1241 ( .A(p_input[8885]), .B(p_input[18885]), .Z(o[8885]) );
  AND U1242 ( .A(p_input[8884]), .B(p_input[18884]), .Z(o[8884]) );
  AND U1243 ( .A(p_input[8883]), .B(p_input[18883]), .Z(o[8883]) );
  AND U1244 ( .A(p_input[8882]), .B(p_input[18882]), .Z(o[8882]) );
  AND U1245 ( .A(p_input[8881]), .B(p_input[18881]), .Z(o[8881]) );
  AND U1246 ( .A(p_input[8880]), .B(p_input[18880]), .Z(o[8880]) );
  AND U1247 ( .A(p_input[887]), .B(p_input[10887]), .Z(o[887]) );
  AND U1248 ( .A(p_input[8879]), .B(p_input[18879]), .Z(o[8879]) );
  AND U1249 ( .A(p_input[8878]), .B(p_input[18878]), .Z(o[8878]) );
  AND U1250 ( .A(p_input[8877]), .B(p_input[18877]), .Z(o[8877]) );
  AND U1251 ( .A(p_input[8876]), .B(p_input[18876]), .Z(o[8876]) );
  AND U1252 ( .A(p_input[8875]), .B(p_input[18875]), .Z(o[8875]) );
  AND U1253 ( .A(p_input[8874]), .B(p_input[18874]), .Z(o[8874]) );
  AND U1254 ( .A(p_input[8873]), .B(p_input[18873]), .Z(o[8873]) );
  AND U1255 ( .A(p_input[8872]), .B(p_input[18872]), .Z(o[8872]) );
  AND U1256 ( .A(p_input[8871]), .B(p_input[18871]), .Z(o[8871]) );
  AND U1257 ( .A(p_input[8870]), .B(p_input[18870]), .Z(o[8870]) );
  AND U1258 ( .A(p_input[886]), .B(p_input[10886]), .Z(o[886]) );
  AND U1259 ( .A(p_input[8869]), .B(p_input[18869]), .Z(o[8869]) );
  AND U1260 ( .A(p_input[8868]), .B(p_input[18868]), .Z(o[8868]) );
  AND U1261 ( .A(p_input[8867]), .B(p_input[18867]), .Z(o[8867]) );
  AND U1262 ( .A(p_input[8866]), .B(p_input[18866]), .Z(o[8866]) );
  AND U1263 ( .A(p_input[8865]), .B(p_input[18865]), .Z(o[8865]) );
  AND U1264 ( .A(p_input[8864]), .B(p_input[18864]), .Z(o[8864]) );
  AND U1265 ( .A(p_input[8863]), .B(p_input[18863]), .Z(o[8863]) );
  AND U1266 ( .A(p_input[8862]), .B(p_input[18862]), .Z(o[8862]) );
  AND U1267 ( .A(p_input[8861]), .B(p_input[18861]), .Z(o[8861]) );
  AND U1268 ( .A(p_input[8860]), .B(p_input[18860]), .Z(o[8860]) );
  AND U1269 ( .A(p_input[885]), .B(p_input[10885]), .Z(o[885]) );
  AND U1270 ( .A(p_input[8859]), .B(p_input[18859]), .Z(o[8859]) );
  AND U1271 ( .A(p_input[8858]), .B(p_input[18858]), .Z(o[8858]) );
  AND U1272 ( .A(p_input[8857]), .B(p_input[18857]), .Z(o[8857]) );
  AND U1273 ( .A(p_input[8856]), .B(p_input[18856]), .Z(o[8856]) );
  AND U1274 ( .A(p_input[8855]), .B(p_input[18855]), .Z(o[8855]) );
  AND U1275 ( .A(p_input[8854]), .B(p_input[18854]), .Z(o[8854]) );
  AND U1276 ( .A(p_input[8853]), .B(p_input[18853]), .Z(o[8853]) );
  AND U1277 ( .A(p_input[8852]), .B(p_input[18852]), .Z(o[8852]) );
  AND U1278 ( .A(p_input[8851]), .B(p_input[18851]), .Z(o[8851]) );
  AND U1279 ( .A(p_input[8850]), .B(p_input[18850]), .Z(o[8850]) );
  AND U1280 ( .A(p_input[884]), .B(p_input[10884]), .Z(o[884]) );
  AND U1281 ( .A(p_input[8849]), .B(p_input[18849]), .Z(o[8849]) );
  AND U1282 ( .A(p_input[8848]), .B(p_input[18848]), .Z(o[8848]) );
  AND U1283 ( .A(p_input[8847]), .B(p_input[18847]), .Z(o[8847]) );
  AND U1284 ( .A(p_input[8846]), .B(p_input[18846]), .Z(o[8846]) );
  AND U1285 ( .A(p_input[8845]), .B(p_input[18845]), .Z(o[8845]) );
  AND U1286 ( .A(p_input[8844]), .B(p_input[18844]), .Z(o[8844]) );
  AND U1287 ( .A(p_input[8843]), .B(p_input[18843]), .Z(o[8843]) );
  AND U1288 ( .A(p_input[8842]), .B(p_input[18842]), .Z(o[8842]) );
  AND U1289 ( .A(p_input[8841]), .B(p_input[18841]), .Z(o[8841]) );
  AND U1290 ( .A(p_input[8840]), .B(p_input[18840]), .Z(o[8840]) );
  AND U1291 ( .A(p_input[883]), .B(p_input[10883]), .Z(o[883]) );
  AND U1292 ( .A(p_input[8839]), .B(p_input[18839]), .Z(o[8839]) );
  AND U1293 ( .A(p_input[8838]), .B(p_input[18838]), .Z(o[8838]) );
  AND U1294 ( .A(p_input[8837]), .B(p_input[18837]), .Z(o[8837]) );
  AND U1295 ( .A(p_input[8836]), .B(p_input[18836]), .Z(o[8836]) );
  AND U1296 ( .A(p_input[8835]), .B(p_input[18835]), .Z(o[8835]) );
  AND U1297 ( .A(p_input[8834]), .B(p_input[18834]), .Z(o[8834]) );
  AND U1298 ( .A(p_input[8833]), .B(p_input[18833]), .Z(o[8833]) );
  AND U1299 ( .A(p_input[8832]), .B(p_input[18832]), .Z(o[8832]) );
  AND U1300 ( .A(p_input[8831]), .B(p_input[18831]), .Z(o[8831]) );
  AND U1301 ( .A(p_input[8830]), .B(p_input[18830]), .Z(o[8830]) );
  AND U1302 ( .A(p_input[882]), .B(p_input[10882]), .Z(o[882]) );
  AND U1303 ( .A(p_input[8829]), .B(p_input[18829]), .Z(o[8829]) );
  AND U1304 ( .A(p_input[8828]), .B(p_input[18828]), .Z(o[8828]) );
  AND U1305 ( .A(p_input[8827]), .B(p_input[18827]), .Z(o[8827]) );
  AND U1306 ( .A(p_input[8826]), .B(p_input[18826]), .Z(o[8826]) );
  AND U1307 ( .A(p_input[8825]), .B(p_input[18825]), .Z(o[8825]) );
  AND U1308 ( .A(p_input[8824]), .B(p_input[18824]), .Z(o[8824]) );
  AND U1309 ( .A(p_input[8823]), .B(p_input[18823]), .Z(o[8823]) );
  AND U1310 ( .A(p_input[8822]), .B(p_input[18822]), .Z(o[8822]) );
  AND U1311 ( .A(p_input[8821]), .B(p_input[18821]), .Z(o[8821]) );
  AND U1312 ( .A(p_input[8820]), .B(p_input[18820]), .Z(o[8820]) );
  AND U1313 ( .A(p_input[881]), .B(p_input[10881]), .Z(o[881]) );
  AND U1314 ( .A(p_input[8819]), .B(p_input[18819]), .Z(o[8819]) );
  AND U1315 ( .A(p_input[8818]), .B(p_input[18818]), .Z(o[8818]) );
  AND U1316 ( .A(p_input[8817]), .B(p_input[18817]), .Z(o[8817]) );
  AND U1317 ( .A(p_input[8816]), .B(p_input[18816]), .Z(o[8816]) );
  AND U1318 ( .A(p_input[8815]), .B(p_input[18815]), .Z(o[8815]) );
  AND U1319 ( .A(p_input[8814]), .B(p_input[18814]), .Z(o[8814]) );
  AND U1320 ( .A(p_input[8813]), .B(p_input[18813]), .Z(o[8813]) );
  AND U1321 ( .A(p_input[8812]), .B(p_input[18812]), .Z(o[8812]) );
  AND U1322 ( .A(p_input[8811]), .B(p_input[18811]), .Z(o[8811]) );
  AND U1323 ( .A(p_input[8810]), .B(p_input[18810]), .Z(o[8810]) );
  AND U1324 ( .A(p_input[880]), .B(p_input[10880]), .Z(o[880]) );
  AND U1325 ( .A(p_input[8809]), .B(p_input[18809]), .Z(o[8809]) );
  AND U1326 ( .A(p_input[8808]), .B(p_input[18808]), .Z(o[8808]) );
  AND U1327 ( .A(p_input[8807]), .B(p_input[18807]), .Z(o[8807]) );
  AND U1328 ( .A(p_input[8806]), .B(p_input[18806]), .Z(o[8806]) );
  AND U1329 ( .A(p_input[8805]), .B(p_input[18805]), .Z(o[8805]) );
  AND U1330 ( .A(p_input[8804]), .B(p_input[18804]), .Z(o[8804]) );
  AND U1331 ( .A(p_input[8803]), .B(p_input[18803]), .Z(o[8803]) );
  AND U1332 ( .A(p_input[8802]), .B(p_input[18802]), .Z(o[8802]) );
  AND U1333 ( .A(p_input[8801]), .B(p_input[18801]), .Z(o[8801]) );
  AND U1334 ( .A(p_input[8800]), .B(p_input[18800]), .Z(o[8800]) );
  AND U1335 ( .A(p_input[87]), .B(p_input[10087]), .Z(o[87]) );
  AND U1336 ( .A(p_input[879]), .B(p_input[10879]), .Z(o[879]) );
  AND U1337 ( .A(p_input[8799]), .B(p_input[18799]), .Z(o[8799]) );
  AND U1338 ( .A(p_input[8798]), .B(p_input[18798]), .Z(o[8798]) );
  AND U1339 ( .A(p_input[8797]), .B(p_input[18797]), .Z(o[8797]) );
  AND U1340 ( .A(p_input[8796]), .B(p_input[18796]), .Z(o[8796]) );
  AND U1341 ( .A(p_input[8795]), .B(p_input[18795]), .Z(o[8795]) );
  AND U1342 ( .A(p_input[8794]), .B(p_input[18794]), .Z(o[8794]) );
  AND U1343 ( .A(p_input[8793]), .B(p_input[18793]), .Z(o[8793]) );
  AND U1344 ( .A(p_input[8792]), .B(p_input[18792]), .Z(o[8792]) );
  AND U1345 ( .A(p_input[8791]), .B(p_input[18791]), .Z(o[8791]) );
  AND U1346 ( .A(p_input[8790]), .B(p_input[18790]), .Z(o[8790]) );
  AND U1347 ( .A(p_input[878]), .B(p_input[10878]), .Z(o[878]) );
  AND U1348 ( .A(p_input[8789]), .B(p_input[18789]), .Z(o[8789]) );
  AND U1349 ( .A(p_input[8788]), .B(p_input[18788]), .Z(o[8788]) );
  AND U1350 ( .A(p_input[8787]), .B(p_input[18787]), .Z(o[8787]) );
  AND U1351 ( .A(p_input[8786]), .B(p_input[18786]), .Z(o[8786]) );
  AND U1352 ( .A(p_input[8785]), .B(p_input[18785]), .Z(o[8785]) );
  AND U1353 ( .A(p_input[8784]), .B(p_input[18784]), .Z(o[8784]) );
  AND U1354 ( .A(p_input[8783]), .B(p_input[18783]), .Z(o[8783]) );
  AND U1355 ( .A(p_input[8782]), .B(p_input[18782]), .Z(o[8782]) );
  AND U1356 ( .A(p_input[8781]), .B(p_input[18781]), .Z(o[8781]) );
  AND U1357 ( .A(p_input[8780]), .B(p_input[18780]), .Z(o[8780]) );
  AND U1358 ( .A(p_input[877]), .B(p_input[10877]), .Z(o[877]) );
  AND U1359 ( .A(p_input[8779]), .B(p_input[18779]), .Z(o[8779]) );
  AND U1360 ( .A(p_input[8778]), .B(p_input[18778]), .Z(o[8778]) );
  AND U1361 ( .A(p_input[8777]), .B(p_input[18777]), .Z(o[8777]) );
  AND U1362 ( .A(p_input[8776]), .B(p_input[18776]), .Z(o[8776]) );
  AND U1363 ( .A(p_input[8775]), .B(p_input[18775]), .Z(o[8775]) );
  AND U1364 ( .A(p_input[8774]), .B(p_input[18774]), .Z(o[8774]) );
  AND U1365 ( .A(p_input[8773]), .B(p_input[18773]), .Z(o[8773]) );
  AND U1366 ( .A(p_input[8772]), .B(p_input[18772]), .Z(o[8772]) );
  AND U1367 ( .A(p_input[8771]), .B(p_input[18771]), .Z(o[8771]) );
  AND U1368 ( .A(p_input[8770]), .B(p_input[18770]), .Z(o[8770]) );
  AND U1369 ( .A(p_input[876]), .B(p_input[10876]), .Z(o[876]) );
  AND U1370 ( .A(p_input[8769]), .B(p_input[18769]), .Z(o[8769]) );
  AND U1371 ( .A(p_input[8768]), .B(p_input[18768]), .Z(o[8768]) );
  AND U1372 ( .A(p_input[8767]), .B(p_input[18767]), .Z(o[8767]) );
  AND U1373 ( .A(p_input[8766]), .B(p_input[18766]), .Z(o[8766]) );
  AND U1374 ( .A(p_input[8765]), .B(p_input[18765]), .Z(o[8765]) );
  AND U1375 ( .A(p_input[8764]), .B(p_input[18764]), .Z(o[8764]) );
  AND U1376 ( .A(p_input[8763]), .B(p_input[18763]), .Z(o[8763]) );
  AND U1377 ( .A(p_input[8762]), .B(p_input[18762]), .Z(o[8762]) );
  AND U1378 ( .A(p_input[8761]), .B(p_input[18761]), .Z(o[8761]) );
  AND U1379 ( .A(p_input[8760]), .B(p_input[18760]), .Z(o[8760]) );
  AND U1380 ( .A(p_input[875]), .B(p_input[10875]), .Z(o[875]) );
  AND U1381 ( .A(p_input[8759]), .B(p_input[18759]), .Z(o[8759]) );
  AND U1382 ( .A(p_input[8758]), .B(p_input[18758]), .Z(o[8758]) );
  AND U1383 ( .A(p_input[8757]), .B(p_input[18757]), .Z(o[8757]) );
  AND U1384 ( .A(p_input[8756]), .B(p_input[18756]), .Z(o[8756]) );
  AND U1385 ( .A(p_input[8755]), .B(p_input[18755]), .Z(o[8755]) );
  AND U1386 ( .A(p_input[8754]), .B(p_input[18754]), .Z(o[8754]) );
  AND U1387 ( .A(p_input[8753]), .B(p_input[18753]), .Z(o[8753]) );
  AND U1388 ( .A(p_input[8752]), .B(p_input[18752]), .Z(o[8752]) );
  AND U1389 ( .A(p_input[8751]), .B(p_input[18751]), .Z(o[8751]) );
  AND U1390 ( .A(p_input[8750]), .B(p_input[18750]), .Z(o[8750]) );
  AND U1391 ( .A(p_input[874]), .B(p_input[10874]), .Z(o[874]) );
  AND U1392 ( .A(p_input[8749]), .B(p_input[18749]), .Z(o[8749]) );
  AND U1393 ( .A(p_input[8748]), .B(p_input[18748]), .Z(o[8748]) );
  AND U1394 ( .A(p_input[8747]), .B(p_input[18747]), .Z(o[8747]) );
  AND U1395 ( .A(p_input[8746]), .B(p_input[18746]), .Z(o[8746]) );
  AND U1396 ( .A(p_input[8745]), .B(p_input[18745]), .Z(o[8745]) );
  AND U1397 ( .A(p_input[8744]), .B(p_input[18744]), .Z(o[8744]) );
  AND U1398 ( .A(p_input[8743]), .B(p_input[18743]), .Z(o[8743]) );
  AND U1399 ( .A(p_input[8742]), .B(p_input[18742]), .Z(o[8742]) );
  AND U1400 ( .A(p_input[8741]), .B(p_input[18741]), .Z(o[8741]) );
  AND U1401 ( .A(p_input[8740]), .B(p_input[18740]), .Z(o[8740]) );
  AND U1402 ( .A(p_input[873]), .B(p_input[10873]), .Z(o[873]) );
  AND U1403 ( .A(p_input[8739]), .B(p_input[18739]), .Z(o[8739]) );
  AND U1404 ( .A(p_input[8738]), .B(p_input[18738]), .Z(o[8738]) );
  AND U1405 ( .A(p_input[8737]), .B(p_input[18737]), .Z(o[8737]) );
  AND U1406 ( .A(p_input[8736]), .B(p_input[18736]), .Z(o[8736]) );
  AND U1407 ( .A(p_input[8735]), .B(p_input[18735]), .Z(o[8735]) );
  AND U1408 ( .A(p_input[8734]), .B(p_input[18734]), .Z(o[8734]) );
  AND U1409 ( .A(p_input[8733]), .B(p_input[18733]), .Z(o[8733]) );
  AND U1410 ( .A(p_input[8732]), .B(p_input[18732]), .Z(o[8732]) );
  AND U1411 ( .A(p_input[8731]), .B(p_input[18731]), .Z(o[8731]) );
  AND U1412 ( .A(p_input[8730]), .B(p_input[18730]), .Z(o[8730]) );
  AND U1413 ( .A(p_input[872]), .B(p_input[10872]), .Z(o[872]) );
  AND U1414 ( .A(p_input[8729]), .B(p_input[18729]), .Z(o[8729]) );
  AND U1415 ( .A(p_input[8728]), .B(p_input[18728]), .Z(o[8728]) );
  AND U1416 ( .A(p_input[8727]), .B(p_input[18727]), .Z(o[8727]) );
  AND U1417 ( .A(p_input[8726]), .B(p_input[18726]), .Z(o[8726]) );
  AND U1418 ( .A(p_input[8725]), .B(p_input[18725]), .Z(o[8725]) );
  AND U1419 ( .A(p_input[8724]), .B(p_input[18724]), .Z(o[8724]) );
  AND U1420 ( .A(p_input[8723]), .B(p_input[18723]), .Z(o[8723]) );
  AND U1421 ( .A(p_input[8722]), .B(p_input[18722]), .Z(o[8722]) );
  AND U1422 ( .A(p_input[8721]), .B(p_input[18721]), .Z(o[8721]) );
  AND U1423 ( .A(p_input[8720]), .B(p_input[18720]), .Z(o[8720]) );
  AND U1424 ( .A(p_input[871]), .B(p_input[10871]), .Z(o[871]) );
  AND U1425 ( .A(p_input[8719]), .B(p_input[18719]), .Z(o[8719]) );
  AND U1426 ( .A(p_input[8718]), .B(p_input[18718]), .Z(o[8718]) );
  AND U1427 ( .A(p_input[8717]), .B(p_input[18717]), .Z(o[8717]) );
  AND U1428 ( .A(p_input[8716]), .B(p_input[18716]), .Z(o[8716]) );
  AND U1429 ( .A(p_input[8715]), .B(p_input[18715]), .Z(o[8715]) );
  AND U1430 ( .A(p_input[8714]), .B(p_input[18714]), .Z(o[8714]) );
  AND U1431 ( .A(p_input[8713]), .B(p_input[18713]), .Z(o[8713]) );
  AND U1432 ( .A(p_input[8712]), .B(p_input[18712]), .Z(o[8712]) );
  AND U1433 ( .A(p_input[8711]), .B(p_input[18711]), .Z(o[8711]) );
  AND U1434 ( .A(p_input[8710]), .B(p_input[18710]), .Z(o[8710]) );
  AND U1435 ( .A(p_input[870]), .B(p_input[10870]), .Z(o[870]) );
  AND U1436 ( .A(p_input[8709]), .B(p_input[18709]), .Z(o[8709]) );
  AND U1437 ( .A(p_input[8708]), .B(p_input[18708]), .Z(o[8708]) );
  AND U1438 ( .A(p_input[8707]), .B(p_input[18707]), .Z(o[8707]) );
  AND U1439 ( .A(p_input[8706]), .B(p_input[18706]), .Z(o[8706]) );
  AND U1440 ( .A(p_input[8705]), .B(p_input[18705]), .Z(o[8705]) );
  AND U1441 ( .A(p_input[8704]), .B(p_input[18704]), .Z(o[8704]) );
  AND U1442 ( .A(p_input[8703]), .B(p_input[18703]), .Z(o[8703]) );
  AND U1443 ( .A(p_input[8702]), .B(p_input[18702]), .Z(o[8702]) );
  AND U1444 ( .A(p_input[8701]), .B(p_input[18701]), .Z(o[8701]) );
  AND U1445 ( .A(p_input[8700]), .B(p_input[18700]), .Z(o[8700]) );
  AND U1446 ( .A(p_input[86]), .B(p_input[10086]), .Z(o[86]) );
  AND U1447 ( .A(p_input[869]), .B(p_input[10869]), .Z(o[869]) );
  AND U1448 ( .A(p_input[8699]), .B(p_input[18699]), .Z(o[8699]) );
  AND U1449 ( .A(p_input[8698]), .B(p_input[18698]), .Z(o[8698]) );
  AND U1450 ( .A(p_input[8697]), .B(p_input[18697]), .Z(o[8697]) );
  AND U1451 ( .A(p_input[8696]), .B(p_input[18696]), .Z(o[8696]) );
  AND U1452 ( .A(p_input[8695]), .B(p_input[18695]), .Z(o[8695]) );
  AND U1453 ( .A(p_input[8694]), .B(p_input[18694]), .Z(o[8694]) );
  AND U1454 ( .A(p_input[8693]), .B(p_input[18693]), .Z(o[8693]) );
  AND U1455 ( .A(p_input[8692]), .B(p_input[18692]), .Z(o[8692]) );
  AND U1456 ( .A(p_input[8691]), .B(p_input[18691]), .Z(o[8691]) );
  AND U1457 ( .A(p_input[8690]), .B(p_input[18690]), .Z(o[8690]) );
  AND U1458 ( .A(p_input[868]), .B(p_input[10868]), .Z(o[868]) );
  AND U1459 ( .A(p_input[8689]), .B(p_input[18689]), .Z(o[8689]) );
  AND U1460 ( .A(p_input[8688]), .B(p_input[18688]), .Z(o[8688]) );
  AND U1461 ( .A(p_input[8687]), .B(p_input[18687]), .Z(o[8687]) );
  AND U1462 ( .A(p_input[8686]), .B(p_input[18686]), .Z(o[8686]) );
  AND U1463 ( .A(p_input[8685]), .B(p_input[18685]), .Z(o[8685]) );
  AND U1464 ( .A(p_input[8684]), .B(p_input[18684]), .Z(o[8684]) );
  AND U1465 ( .A(p_input[8683]), .B(p_input[18683]), .Z(o[8683]) );
  AND U1466 ( .A(p_input[8682]), .B(p_input[18682]), .Z(o[8682]) );
  AND U1467 ( .A(p_input[8681]), .B(p_input[18681]), .Z(o[8681]) );
  AND U1468 ( .A(p_input[8680]), .B(p_input[18680]), .Z(o[8680]) );
  AND U1469 ( .A(p_input[867]), .B(p_input[10867]), .Z(o[867]) );
  AND U1470 ( .A(p_input[8679]), .B(p_input[18679]), .Z(o[8679]) );
  AND U1471 ( .A(p_input[8678]), .B(p_input[18678]), .Z(o[8678]) );
  AND U1472 ( .A(p_input[8677]), .B(p_input[18677]), .Z(o[8677]) );
  AND U1473 ( .A(p_input[8676]), .B(p_input[18676]), .Z(o[8676]) );
  AND U1474 ( .A(p_input[8675]), .B(p_input[18675]), .Z(o[8675]) );
  AND U1475 ( .A(p_input[8674]), .B(p_input[18674]), .Z(o[8674]) );
  AND U1476 ( .A(p_input[8673]), .B(p_input[18673]), .Z(o[8673]) );
  AND U1477 ( .A(p_input[8672]), .B(p_input[18672]), .Z(o[8672]) );
  AND U1478 ( .A(p_input[8671]), .B(p_input[18671]), .Z(o[8671]) );
  AND U1479 ( .A(p_input[8670]), .B(p_input[18670]), .Z(o[8670]) );
  AND U1480 ( .A(p_input[866]), .B(p_input[10866]), .Z(o[866]) );
  AND U1481 ( .A(p_input[8669]), .B(p_input[18669]), .Z(o[8669]) );
  AND U1482 ( .A(p_input[8668]), .B(p_input[18668]), .Z(o[8668]) );
  AND U1483 ( .A(p_input[8667]), .B(p_input[18667]), .Z(o[8667]) );
  AND U1484 ( .A(p_input[8666]), .B(p_input[18666]), .Z(o[8666]) );
  AND U1485 ( .A(p_input[8665]), .B(p_input[18665]), .Z(o[8665]) );
  AND U1486 ( .A(p_input[8664]), .B(p_input[18664]), .Z(o[8664]) );
  AND U1487 ( .A(p_input[8663]), .B(p_input[18663]), .Z(o[8663]) );
  AND U1488 ( .A(p_input[8662]), .B(p_input[18662]), .Z(o[8662]) );
  AND U1489 ( .A(p_input[8661]), .B(p_input[18661]), .Z(o[8661]) );
  AND U1490 ( .A(p_input[8660]), .B(p_input[18660]), .Z(o[8660]) );
  AND U1491 ( .A(p_input[865]), .B(p_input[10865]), .Z(o[865]) );
  AND U1492 ( .A(p_input[8659]), .B(p_input[18659]), .Z(o[8659]) );
  AND U1493 ( .A(p_input[8658]), .B(p_input[18658]), .Z(o[8658]) );
  AND U1494 ( .A(p_input[8657]), .B(p_input[18657]), .Z(o[8657]) );
  AND U1495 ( .A(p_input[8656]), .B(p_input[18656]), .Z(o[8656]) );
  AND U1496 ( .A(p_input[8655]), .B(p_input[18655]), .Z(o[8655]) );
  AND U1497 ( .A(p_input[8654]), .B(p_input[18654]), .Z(o[8654]) );
  AND U1498 ( .A(p_input[8653]), .B(p_input[18653]), .Z(o[8653]) );
  AND U1499 ( .A(p_input[8652]), .B(p_input[18652]), .Z(o[8652]) );
  AND U1500 ( .A(p_input[8651]), .B(p_input[18651]), .Z(o[8651]) );
  AND U1501 ( .A(p_input[8650]), .B(p_input[18650]), .Z(o[8650]) );
  AND U1502 ( .A(p_input[864]), .B(p_input[10864]), .Z(o[864]) );
  AND U1503 ( .A(p_input[8649]), .B(p_input[18649]), .Z(o[8649]) );
  AND U1504 ( .A(p_input[8648]), .B(p_input[18648]), .Z(o[8648]) );
  AND U1505 ( .A(p_input[8647]), .B(p_input[18647]), .Z(o[8647]) );
  AND U1506 ( .A(p_input[8646]), .B(p_input[18646]), .Z(o[8646]) );
  AND U1507 ( .A(p_input[8645]), .B(p_input[18645]), .Z(o[8645]) );
  AND U1508 ( .A(p_input[8644]), .B(p_input[18644]), .Z(o[8644]) );
  AND U1509 ( .A(p_input[8643]), .B(p_input[18643]), .Z(o[8643]) );
  AND U1510 ( .A(p_input[8642]), .B(p_input[18642]), .Z(o[8642]) );
  AND U1511 ( .A(p_input[8641]), .B(p_input[18641]), .Z(o[8641]) );
  AND U1512 ( .A(p_input[8640]), .B(p_input[18640]), .Z(o[8640]) );
  AND U1513 ( .A(p_input[863]), .B(p_input[10863]), .Z(o[863]) );
  AND U1514 ( .A(p_input[8639]), .B(p_input[18639]), .Z(o[8639]) );
  AND U1515 ( .A(p_input[8638]), .B(p_input[18638]), .Z(o[8638]) );
  AND U1516 ( .A(p_input[8637]), .B(p_input[18637]), .Z(o[8637]) );
  AND U1517 ( .A(p_input[8636]), .B(p_input[18636]), .Z(o[8636]) );
  AND U1518 ( .A(p_input[8635]), .B(p_input[18635]), .Z(o[8635]) );
  AND U1519 ( .A(p_input[8634]), .B(p_input[18634]), .Z(o[8634]) );
  AND U1520 ( .A(p_input[8633]), .B(p_input[18633]), .Z(o[8633]) );
  AND U1521 ( .A(p_input[8632]), .B(p_input[18632]), .Z(o[8632]) );
  AND U1522 ( .A(p_input[8631]), .B(p_input[18631]), .Z(o[8631]) );
  AND U1523 ( .A(p_input[8630]), .B(p_input[18630]), .Z(o[8630]) );
  AND U1524 ( .A(p_input[862]), .B(p_input[10862]), .Z(o[862]) );
  AND U1525 ( .A(p_input[8629]), .B(p_input[18629]), .Z(o[8629]) );
  AND U1526 ( .A(p_input[8628]), .B(p_input[18628]), .Z(o[8628]) );
  AND U1527 ( .A(p_input[8627]), .B(p_input[18627]), .Z(o[8627]) );
  AND U1528 ( .A(p_input[8626]), .B(p_input[18626]), .Z(o[8626]) );
  AND U1529 ( .A(p_input[8625]), .B(p_input[18625]), .Z(o[8625]) );
  AND U1530 ( .A(p_input[8624]), .B(p_input[18624]), .Z(o[8624]) );
  AND U1531 ( .A(p_input[8623]), .B(p_input[18623]), .Z(o[8623]) );
  AND U1532 ( .A(p_input[8622]), .B(p_input[18622]), .Z(o[8622]) );
  AND U1533 ( .A(p_input[8621]), .B(p_input[18621]), .Z(o[8621]) );
  AND U1534 ( .A(p_input[8620]), .B(p_input[18620]), .Z(o[8620]) );
  AND U1535 ( .A(p_input[861]), .B(p_input[10861]), .Z(o[861]) );
  AND U1536 ( .A(p_input[8619]), .B(p_input[18619]), .Z(o[8619]) );
  AND U1537 ( .A(p_input[8618]), .B(p_input[18618]), .Z(o[8618]) );
  AND U1538 ( .A(p_input[8617]), .B(p_input[18617]), .Z(o[8617]) );
  AND U1539 ( .A(p_input[8616]), .B(p_input[18616]), .Z(o[8616]) );
  AND U1540 ( .A(p_input[8615]), .B(p_input[18615]), .Z(o[8615]) );
  AND U1541 ( .A(p_input[8614]), .B(p_input[18614]), .Z(o[8614]) );
  AND U1542 ( .A(p_input[8613]), .B(p_input[18613]), .Z(o[8613]) );
  AND U1543 ( .A(p_input[8612]), .B(p_input[18612]), .Z(o[8612]) );
  AND U1544 ( .A(p_input[8611]), .B(p_input[18611]), .Z(o[8611]) );
  AND U1545 ( .A(p_input[8610]), .B(p_input[18610]), .Z(o[8610]) );
  AND U1546 ( .A(p_input[860]), .B(p_input[10860]), .Z(o[860]) );
  AND U1547 ( .A(p_input[8609]), .B(p_input[18609]), .Z(o[8609]) );
  AND U1548 ( .A(p_input[8608]), .B(p_input[18608]), .Z(o[8608]) );
  AND U1549 ( .A(p_input[8607]), .B(p_input[18607]), .Z(o[8607]) );
  AND U1550 ( .A(p_input[8606]), .B(p_input[18606]), .Z(o[8606]) );
  AND U1551 ( .A(p_input[8605]), .B(p_input[18605]), .Z(o[8605]) );
  AND U1552 ( .A(p_input[8604]), .B(p_input[18604]), .Z(o[8604]) );
  AND U1553 ( .A(p_input[8603]), .B(p_input[18603]), .Z(o[8603]) );
  AND U1554 ( .A(p_input[8602]), .B(p_input[18602]), .Z(o[8602]) );
  AND U1555 ( .A(p_input[8601]), .B(p_input[18601]), .Z(o[8601]) );
  AND U1556 ( .A(p_input[8600]), .B(p_input[18600]), .Z(o[8600]) );
  AND U1557 ( .A(p_input[85]), .B(p_input[10085]), .Z(o[85]) );
  AND U1558 ( .A(p_input[859]), .B(p_input[10859]), .Z(o[859]) );
  AND U1559 ( .A(p_input[8599]), .B(p_input[18599]), .Z(o[8599]) );
  AND U1560 ( .A(p_input[8598]), .B(p_input[18598]), .Z(o[8598]) );
  AND U1561 ( .A(p_input[8597]), .B(p_input[18597]), .Z(o[8597]) );
  AND U1562 ( .A(p_input[8596]), .B(p_input[18596]), .Z(o[8596]) );
  AND U1563 ( .A(p_input[8595]), .B(p_input[18595]), .Z(o[8595]) );
  AND U1564 ( .A(p_input[8594]), .B(p_input[18594]), .Z(o[8594]) );
  AND U1565 ( .A(p_input[8593]), .B(p_input[18593]), .Z(o[8593]) );
  AND U1566 ( .A(p_input[8592]), .B(p_input[18592]), .Z(o[8592]) );
  AND U1567 ( .A(p_input[8591]), .B(p_input[18591]), .Z(o[8591]) );
  AND U1568 ( .A(p_input[8590]), .B(p_input[18590]), .Z(o[8590]) );
  AND U1569 ( .A(p_input[858]), .B(p_input[10858]), .Z(o[858]) );
  AND U1570 ( .A(p_input[8589]), .B(p_input[18589]), .Z(o[8589]) );
  AND U1571 ( .A(p_input[8588]), .B(p_input[18588]), .Z(o[8588]) );
  AND U1572 ( .A(p_input[8587]), .B(p_input[18587]), .Z(o[8587]) );
  AND U1573 ( .A(p_input[8586]), .B(p_input[18586]), .Z(o[8586]) );
  AND U1574 ( .A(p_input[8585]), .B(p_input[18585]), .Z(o[8585]) );
  AND U1575 ( .A(p_input[8584]), .B(p_input[18584]), .Z(o[8584]) );
  AND U1576 ( .A(p_input[8583]), .B(p_input[18583]), .Z(o[8583]) );
  AND U1577 ( .A(p_input[8582]), .B(p_input[18582]), .Z(o[8582]) );
  AND U1578 ( .A(p_input[8581]), .B(p_input[18581]), .Z(o[8581]) );
  AND U1579 ( .A(p_input[8580]), .B(p_input[18580]), .Z(o[8580]) );
  AND U1580 ( .A(p_input[857]), .B(p_input[10857]), .Z(o[857]) );
  AND U1581 ( .A(p_input[8579]), .B(p_input[18579]), .Z(o[8579]) );
  AND U1582 ( .A(p_input[8578]), .B(p_input[18578]), .Z(o[8578]) );
  AND U1583 ( .A(p_input[8577]), .B(p_input[18577]), .Z(o[8577]) );
  AND U1584 ( .A(p_input[8576]), .B(p_input[18576]), .Z(o[8576]) );
  AND U1585 ( .A(p_input[8575]), .B(p_input[18575]), .Z(o[8575]) );
  AND U1586 ( .A(p_input[8574]), .B(p_input[18574]), .Z(o[8574]) );
  AND U1587 ( .A(p_input[8573]), .B(p_input[18573]), .Z(o[8573]) );
  AND U1588 ( .A(p_input[8572]), .B(p_input[18572]), .Z(o[8572]) );
  AND U1589 ( .A(p_input[8571]), .B(p_input[18571]), .Z(o[8571]) );
  AND U1590 ( .A(p_input[8570]), .B(p_input[18570]), .Z(o[8570]) );
  AND U1591 ( .A(p_input[856]), .B(p_input[10856]), .Z(o[856]) );
  AND U1592 ( .A(p_input[8569]), .B(p_input[18569]), .Z(o[8569]) );
  AND U1593 ( .A(p_input[8568]), .B(p_input[18568]), .Z(o[8568]) );
  AND U1594 ( .A(p_input[8567]), .B(p_input[18567]), .Z(o[8567]) );
  AND U1595 ( .A(p_input[8566]), .B(p_input[18566]), .Z(o[8566]) );
  AND U1596 ( .A(p_input[8565]), .B(p_input[18565]), .Z(o[8565]) );
  AND U1597 ( .A(p_input[8564]), .B(p_input[18564]), .Z(o[8564]) );
  AND U1598 ( .A(p_input[8563]), .B(p_input[18563]), .Z(o[8563]) );
  AND U1599 ( .A(p_input[8562]), .B(p_input[18562]), .Z(o[8562]) );
  AND U1600 ( .A(p_input[8561]), .B(p_input[18561]), .Z(o[8561]) );
  AND U1601 ( .A(p_input[8560]), .B(p_input[18560]), .Z(o[8560]) );
  AND U1602 ( .A(p_input[855]), .B(p_input[10855]), .Z(o[855]) );
  AND U1603 ( .A(p_input[8559]), .B(p_input[18559]), .Z(o[8559]) );
  AND U1604 ( .A(p_input[8558]), .B(p_input[18558]), .Z(o[8558]) );
  AND U1605 ( .A(p_input[8557]), .B(p_input[18557]), .Z(o[8557]) );
  AND U1606 ( .A(p_input[8556]), .B(p_input[18556]), .Z(o[8556]) );
  AND U1607 ( .A(p_input[8555]), .B(p_input[18555]), .Z(o[8555]) );
  AND U1608 ( .A(p_input[8554]), .B(p_input[18554]), .Z(o[8554]) );
  AND U1609 ( .A(p_input[8553]), .B(p_input[18553]), .Z(o[8553]) );
  AND U1610 ( .A(p_input[8552]), .B(p_input[18552]), .Z(o[8552]) );
  AND U1611 ( .A(p_input[8551]), .B(p_input[18551]), .Z(o[8551]) );
  AND U1612 ( .A(p_input[8550]), .B(p_input[18550]), .Z(o[8550]) );
  AND U1613 ( .A(p_input[854]), .B(p_input[10854]), .Z(o[854]) );
  AND U1614 ( .A(p_input[8549]), .B(p_input[18549]), .Z(o[8549]) );
  AND U1615 ( .A(p_input[8548]), .B(p_input[18548]), .Z(o[8548]) );
  AND U1616 ( .A(p_input[8547]), .B(p_input[18547]), .Z(o[8547]) );
  AND U1617 ( .A(p_input[8546]), .B(p_input[18546]), .Z(o[8546]) );
  AND U1618 ( .A(p_input[8545]), .B(p_input[18545]), .Z(o[8545]) );
  AND U1619 ( .A(p_input[8544]), .B(p_input[18544]), .Z(o[8544]) );
  AND U1620 ( .A(p_input[8543]), .B(p_input[18543]), .Z(o[8543]) );
  AND U1621 ( .A(p_input[8542]), .B(p_input[18542]), .Z(o[8542]) );
  AND U1622 ( .A(p_input[8541]), .B(p_input[18541]), .Z(o[8541]) );
  AND U1623 ( .A(p_input[8540]), .B(p_input[18540]), .Z(o[8540]) );
  AND U1624 ( .A(p_input[853]), .B(p_input[10853]), .Z(o[853]) );
  AND U1625 ( .A(p_input[8539]), .B(p_input[18539]), .Z(o[8539]) );
  AND U1626 ( .A(p_input[8538]), .B(p_input[18538]), .Z(o[8538]) );
  AND U1627 ( .A(p_input[8537]), .B(p_input[18537]), .Z(o[8537]) );
  AND U1628 ( .A(p_input[8536]), .B(p_input[18536]), .Z(o[8536]) );
  AND U1629 ( .A(p_input[8535]), .B(p_input[18535]), .Z(o[8535]) );
  AND U1630 ( .A(p_input[8534]), .B(p_input[18534]), .Z(o[8534]) );
  AND U1631 ( .A(p_input[8533]), .B(p_input[18533]), .Z(o[8533]) );
  AND U1632 ( .A(p_input[8532]), .B(p_input[18532]), .Z(o[8532]) );
  AND U1633 ( .A(p_input[8531]), .B(p_input[18531]), .Z(o[8531]) );
  AND U1634 ( .A(p_input[8530]), .B(p_input[18530]), .Z(o[8530]) );
  AND U1635 ( .A(p_input[852]), .B(p_input[10852]), .Z(o[852]) );
  AND U1636 ( .A(p_input[8529]), .B(p_input[18529]), .Z(o[8529]) );
  AND U1637 ( .A(p_input[8528]), .B(p_input[18528]), .Z(o[8528]) );
  AND U1638 ( .A(p_input[8527]), .B(p_input[18527]), .Z(o[8527]) );
  AND U1639 ( .A(p_input[8526]), .B(p_input[18526]), .Z(o[8526]) );
  AND U1640 ( .A(p_input[8525]), .B(p_input[18525]), .Z(o[8525]) );
  AND U1641 ( .A(p_input[8524]), .B(p_input[18524]), .Z(o[8524]) );
  AND U1642 ( .A(p_input[8523]), .B(p_input[18523]), .Z(o[8523]) );
  AND U1643 ( .A(p_input[8522]), .B(p_input[18522]), .Z(o[8522]) );
  AND U1644 ( .A(p_input[8521]), .B(p_input[18521]), .Z(o[8521]) );
  AND U1645 ( .A(p_input[8520]), .B(p_input[18520]), .Z(o[8520]) );
  AND U1646 ( .A(p_input[851]), .B(p_input[10851]), .Z(o[851]) );
  AND U1647 ( .A(p_input[8519]), .B(p_input[18519]), .Z(o[8519]) );
  AND U1648 ( .A(p_input[8518]), .B(p_input[18518]), .Z(o[8518]) );
  AND U1649 ( .A(p_input[8517]), .B(p_input[18517]), .Z(o[8517]) );
  AND U1650 ( .A(p_input[8516]), .B(p_input[18516]), .Z(o[8516]) );
  AND U1651 ( .A(p_input[8515]), .B(p_input[18515]), .Z(o[8515]) );
  AND U1652 ( .A(p_input[8514]), .B(p_input[18514]), .Z(o[8514]) );
  AND U1653 ( .A(p_input[8513]), .B(p_input[18513]), .Z(o[8513]) );
  AND U1654 ( .A(p_input[8512]), .B(p_input[18512]), .Z(o[8512]) );
  AND U1655 ( .A(p_input[8511]), .B(p_input[18511]), .Z(o[8511]) );
  AND U1656 ( .A(p_input[8510]), .B(p_input[18510]), .Z(o[8510]) );
  AND U1657 ( .A(p_input[850]), .B(p_input[10850]), .Z(o[850]) );
  AND U1658 ( .A(p_input[8509]), .B(p_input[18509]), .Z(o[8509]) );
  AND U1659 ( .A(p_input[8508]), .B(p_input[18508]), .Z(o[8508]) );
  AND U1660 ( .A(p_input[8507]), .B(p_input[18507]), .Z(o[8507]) );
  AND U1661 ( .A(p_input[8506]), .B(p_input[18506]), .Z(o[8506]) );
  AND U1662 ( .A(p_input[8505]), .B(p_input[18505]), .Z(o[8505]) );
  AND U1663 ( .A(p_input[8504]), .B(p_input[18504]), .Z(o[8504]) );
  AND U1664 ( .A(p_input[8503]), .B(p_input[18503]), .Z(o[8503]) );
  AND U1665 ( .A(p_input[8502]), .B(p_input[18502]), .Z(o[8502]) );
  AND U1666 ( .A(p_input[8501]), .B(p_input[18501]), .Z(o[8501]) );
  AND U1667 ( .A(p_input[8500]), .B(p_input[18500]), .Z(o[8500]) );
  AND U1668 ( .A(p_input[84]), .B(p_input[10084]), .Z(o[84]) );
  AND U1669 ( .A(p_input[849]), .B(p_input[10849]), .Z(o[849]) );
  AND U1670 ( .A(p_input[8499]), .B(p_input[18499]), .Z(o[8499]) );
  AND U1671 ( .A(p_input[8498]), .B(p_input[18498]), .Z(o[8498]) );
  AND U1672 ( .A(p_input[8497]), .B(p_input[18497]), .Z(o[8497]) );
  AND U1673 ( .A(p_input[8496]), .B(p_input[18496]), .Z(o[8496]) );
  AND U1674 ( .A(p_input[8495]), .B(p_input[18495]), .Z(o[8495]) );
  AND U1675 ( .A(p_input[8494]), .B(p_input[18494]), .Z(o[8494]) );
  AND U1676 ( .A(p_input[8493]), .B(p_input[18493]), .Z(o[8493]) );
  AND U1677 ( .A(p_input[8492]), .B(p_input[18492]), .Z(o[8492]) );
  AND U1678 ( .A(p_input[8491]), .B(p_input[18491]), .Z(o[8491]) );
  AND U1679 ( .A(p_input[8490]), .B(p_input[18490]), .Z(o[8490]) );
  AND U1680 ( .A(p_input[848]), .B(p_input[10848]), .Z(o[848]) );
  AND U1681 ( .A(p_input[8489]), .B(p_input[18489]), .Z(o[8489]) );
  AND U1682 ( .A(p_input[8488]), .B(p_input[18488]), .Z(o[8488]) );
  AND U1683 ( .A(p_input[8487]), .B(p_input[18487]), .Z(o[8487]) );
  AND U1684 ( .A(p_input[8486]), .B(p_input[18486]), .Z(o[8486]) );
  AND U1685 ( .A(p_input[8485]), .B(p_input[18485]), .Z(o[8485]) );
  AND U1686 ( .A(p_input[8484]), .B(p_input[18484]), .Z(o[8484]) );
  AND U1687 ( .A(p_input[8483]), .B(p_input[18483]), .Z(o[8483]) );
  AND U1688 ( .A(p_input[8482]), .B(p_input[18482]), .Z(o[8482]) );
  AND U1689 ( .A(p_input[8481]), .B(p_input[18481]), .Z(o[8481]) );
  AND U1690 ( .A(p_input[8480]), .B(p_input[18480]), .Z(o[8480]) );
  AND U1691 ( .A(p_input[847]), .B(p_input[10847]), .Z(o[847]) );
  AND U1692 ( .A(p_input[8479]), .B(p_input[18479]), .Z(o[8479]) );
  AND U1693 ( .A(p_input[8478]), .B(p_input[18478]), .Z(o[8478]) );
  AND U1694 ( .A(p_input[8477]), .B(p_input[18477]), .Z(o[8477]) );
  AND U1695 ( .A(p_input[8476]), .B(p_input[18476]), .Z(o[8476]) );
  AND U1696 ( .A(p_input[8475]), .B(p_input[18475]), .Z(o[8475]) );
  AND U1697 ( .A(p_input[8474]), .B(p_input[18474]), .Z(o[8474]) );
  AND U1698 ( .A(p_input[8473]), .B(p_input[18473]), .Z(o[8473]) );
  AND U1699 ( .A(p_input[8472]), .B(p_input[18472]), .Z(o[8472]) );
  AND U1700 ( .A(p_input[8471]), .B(p_input[18471]), .Z(o[8471]) );
  AND U1701 ( .A(p_input[8470]), .B(p_input[18470]), .Z(o[8470]) );
  AND U1702 ( .A(p_input[846]), .B(p_input[10846]), .Z(o[846]) );
  AND U1703 ( .A(p_input[8469]), .B(p_input[18469]), .Z(o[8469]) );
  AND U1704 ( .A(p_input[8468]), .B(p_input[18468]), .Z(o[8468]) );
  AND U1705 ( .A(p_input[8467]), .B(p_input[18467]), .Z(o[8467]) );
  AND U1706 ( .A(p_input[8466]), .B(p_input[18466]), .Z(o[8466]) );
  AND U1707 ( .A(p_input[8465]), .B(p_input[18465]), .Z(o[8465]) );
  AND U1708 ( .A(p_input[8464]), .B(p_input[18464]), .Z(o[8464]) );
  AND U1709 ( .A(p_input[8463]), .B(p_input[18463]), .Z(o[8463]) );
  AND U1710 ( .A(p_input[8462]), .B(p_input[18462]), .Z(o[8462]) );
  AND U1711 ( .A(p_input[8461]), .B(p_input[18461]), .Z(o[8461]) );
  AND U1712 ( .A(p_input[8460]), .B(p_input[18460]), .Z(o[8460]) );
  AND U1713 ( .A(p_input[845]), .B(p_input[10845]), .Z(o[845]) );
  AND U1714 ( .A(p_input[8459]), .B(p_input[18459]), .Z(o[8459]) );
  AND U1715 ( .A(p_input[8458]), .B(p_input[18458]), .Z(o[8458]) );
  AND U1716 ( .A(p_input[8457]), .B(p_input[18457]), .Z(o[8457]) );
  AND U1717 ( .A(p_input[8456]), .B(p_input[18456]), .Z(o[8456]) );
  AND U1718 ( .A(p_input[8455]), .B(p_input[18455]), .Z(o[8455]) );
  AND U1719 ( .A(p_input[8454]), .B(p_input[18454]), .Z(o[8454]) );
  AND U1720 ( .A(p_input[8453]), .B(p_input[18453]), .Z(o[8453]) );
  AND U1721 ( .A(p_input[8452]), .B(p_input[18452]), .Z(o[8452]) );
  AND U1722 ( .A(p_input[8451]), .B(p_input[18451]), .Z(o[8451]) );
  AND U1723 ( .A(p_input[8450]), .B(p_input[18450]), .Z(o[8450]) );
  AND U1724 ( .A(p_input[844]), .B(p_input[10844]), .Z(o[844]) );
  AND U1725 ( .A(p_input[8449]), .B(p_input[18449]), .Z(o[8449]) );
  AND U1726 ( .A(p_input[8448]), .B(p_input[18448]), .Z(o[8448]) );
  AND U1727 ( .A(p_input[8447]), .B(p_input[18447]), .Z(o[8447]) );
  AND U1728 ( .A(p_input[8446]), .B(p_input[18446]), .Z(o[8446]) );
  AND U1729 ( .A(p_input[8445]), .B(p_input[18445]), .Z(o[8445]) );
  AND U1730 ( .A(p_input[8444]), .B(p_input[18444]), .Z(o[8444]) );
  AND U1731 ( .A(p_input[8443]), .B(p_input[18443]), .Z(o[8443]) );
  AND U1732 ( .A(p_input[8442]), .B(p_input[18442]), .Z(o[8442]) );
  AND U1733 ( .A(p_input[8441]), .B(p_input[18441]), .Z(o[8441]) );
  AND U1734 ( .A(p_input[8440]), .B(p_input[18440]), .Z(o[8440]) );
  AND U1735 ( .A(p_input[843]), .B(p_input[10843]), .Z(o[843]) );
  AND U1736 ( .A(p_input[8439]), .B(p_input[18439]), .Z(o[8439]) );
  AND U1737 ( .A(p_input[8438]), .B(p_input[18438]), .Z(o[8438]) );
  AND U1738 ( .A(p_input[8437]), .B(p_input[18437]), .Z(o[8437]) );
  AND U1739 ( .A(p_input[8436]), .B(p_input[18436]), .Z(o[8436]) );
  AND U1740 ( .A(p_input[8435]), .B(p_input[18435]), .Z(o[8435]) );
  AND U1741 ( .A(p_input[8434]), .B(p_input[18434]), .Z(o[8434]) );
  AND U1742 ( .A(p_input[8433]), .B(p_input[18433]), .Z(o[8433]) );
  AND U1743 ( .A(p_input[8432]), .B(p_input[18432]), .Z(o[8432]) );
  AND U1744 ( .A(p_input[8431]), .B(p_input[18431]), .Z(o[8431]) );
  AND U1745 ( .A(p_input[8430]), .B(p_input[18430]), .Z(o[8430]) );
  AND U1746 ( .A(p_input[842]), .B(p_input[10842]), .Z(o[842]) );
  AND U1747 ( .A(p_input[8429]), .B(p_input[18429]), .Z(o[8429]) );
  AND U1748 ( .A(p_input[8428]), .B(p_input[18428]), .Z(o[8428]) );
  AND U1749 ( .A(p_input[8427]), .B(p_input[18427]), .Z(o[8427]) );
  AND U1750 ( .A(p_input[8426]), .B(p_input[18426]), .Z(o[8426]) );
  AND U1751 ( .A(p_input[8425]), .B(p_input[18425]), .Z(o[8425]) );
  AND U1752 ( .A(p_input[8424]), .B(p_input[18424]), .Z(o[8424]) );
  AND U1753 ( .A(p_input[8423]), .B(p_input[18423]), .Z(o[8423]) );
  AND U1754 ( .A(p_input[8422]), .B(p_input[18422]), .Z(o[8422]) );
  AND U1755 ( .A(p_input[8421]), .B(p_input[18421]), .Z(o[8421]) );
  AND U1756 ( .A(p_input[8420]), .B(p_input[18420]), .Z(o[8420]) );
  AND U1757 ( .A(p_input[841]), .B(p_input[10841]), .Z(o[841]) );
  AND U1758 ( .A(p_input[8419]), .B(p_input[18419]), .Z(o[8419]) );
  AND U1759 ( .A(p_input[8418]), .B(p_input[18418]), .Z(o[8418]) );
  AND U1760 ( .A(p_input[8417]), .B(p_input[18417]), .Z(o[8417]) );
  AND U1761 ( .A(p_input[8416]), .B(p_input[18416]), .Z(o[8416]) );
  AND U1762 ( .A(p_input[8415]), .B(p_input[18415]), .Z(o[8415]) );
  AND U1763 ( .A(p_input[8414]), .B(p_input[18414]), .Z(o[8414]) );
  AND U1764 ( .A(p_input[8413]), .B(p_input[18413]), .Z(o[8413]) );
  AND U1765 ( .A(p_input[8412]), .B(p_input[18412]), .Z(o[8412]) );
  AND U1766 ( .A(p_input[8411]), .B(p_input[18411]), .Z(o[8411]) );
  AND U1767 ( .A(p_input[8410]), .B(p_input[18410]), .Z(o[8410]) );
  AND U1768 ( .A(p_input[840]), .B(p_input[10840]), .Z(o[840]) );
  AND U1769 ( .A(p_input[8409]), .B(p_input[18409]), .Z(o[8409]) );
  AND U1770 ( .A(p_input[8408]), .B(p_input[18408]), .Z(o[8408]) );
  AND U1771 ( .A(p_input[8407]), .B(p_input[18407]), .Z(o[8407]) );
  AND U1772 ( .A(p_input[8406]), .B(p_input[18406]), .Z(o[8406]) );
  AND U1773 ( .A(p_input[8405]), .B(p_input[18405]), .Z(o[8405]) );
  AND U1774 ( .A(p_input[8404]), .B(p_input[18404]), .Z(o[8404]) );
  AND U1775 ( .A(p_input[8403]), .B(p_input[18403]), .Z(o[8403]) );
  AND U1776 ( .A(p_input[8402]), .B(p_input[18402]), .Z(o[8402]) );
  AND U1777 ( .A(p_input[8401]), .B(p_input[18401]), .Z(o[8401]) );
  AND U1778 ( .A(p_input[8400]), .B(p_input[18400]), .Z(o[8400]) );
  AND U1779 ( .A(p_input[83]), .B(p_input[10083]), .Z(o[83]) );
  AND U1780 ( .A(p_input[839]), .B(p_input[10839]), .Z(o[839]) );
  AND U1781 ( .A(p_input[8399]), .B(p_input[18399]), .Z(o[8399]) );
  AND U1782 ( .A(p_input[8398]), .B(p_input[18398]), .Z(o[8398]) );
  AND U1783 ( .A(p_input[8397]), .B(p_input[18397]), .Z(o[8397]) );
  AND U1784 ( .A(p_input[8396]), .B(p_input[18396]), .Z(o[8396]) );
  AND U1785 ( .A(p_input[8395]), .B(p_input[18395]), .Z(o[8395]) );
  AND U1786 ( .A(p_input[8394]), .B(p_input[18394]), .Z(o[8394]) );
  AND U1787 ( .A(p_input[8393]), .B(p_input[18393]), .Z(o[8393]) );
  AND U1788 ( .A(p_input[8392]), .B(p_input[18392]), .Z(o[8392]) );
  AND U1789 ( .A(p_input[8391]), .B(p_input[18391]), .Z(o[8391]) );
  AND U1790 ( .A(p_input[8390]), .B(p_input[18390]), .Z(o[8390]) );
  AND U1791 ( .A(p_input[838]), .B(p_input[10838]), .Z(o[838]) );
  AND U1792 ( .A(p_input[8389]), .B(p_input[18389]), .Z(o[8389]) );
  AND U1793 ( .A(p_input[8388]), .B(p_input[18388]), .Z(o[8388]) );
  AND U1794 ( .A(p_input[8387]), .B(p_input[18387]), .Z(o[8387]) );
  AND U1795 ( .A(p_input[8386]), .B(p_input[18386]), .Z(o[8386]) );
  AND U1796 ( .A(p_input[8385]), .B(p_input[18385]), .Z(o[8385]) );
  AND U1797 ( .A(p_input[8384]), .B(p_input[18384]), .Z(o[8384]) );
  AND U1798 ( .A(p_input[8383]), .B(p_input[18383]), .Z(o[8383]) );
  AND U1799 ( .A(p_input[8382]), .B(p_input[18382]), .Z(o[8382]) );
  AND U1800 ( .A(p_input[8381]), .B(p_input[18381]), .Z(o[8381]) );
  AND U1801 ( .A(p_input[8380]), .B(p_input[18380]), .Z(o[8380]) );
  AND U1802 ( .A(p_input[837]), .B(p_input[10837]), .Z(o[837]) );
  AND U1803 ( .A(p_input[8379]), .B(p_input[18379]), .Z(o[8379]) );
  AND U1804 ( .A(p_input[8378]), .B(p_input[18378]), .Z(o[8378]) );
  AND U1805 ( .A(p_input[8377]), .B(p_input[18377]), .Z(o[8377]) );
  AND U1806 ( .A(p_input[8376]), .B(p_input[18376]), .Z(o[8376]) );
  AND U1807 ( .A(p_input[8375]), .B(p_input[18375]), .Z(o[8375]) );
  AND U1808 ( .A(p_input[8374]), .B(p_input[18374]), .Z(o[8374]) );
  AND U1809 ( .A(p_input[8373]), .B(p_input[18373]), .Z(o[8373]) );
  AND U1810 ( .A(p_input[8372]), .B(p_input[18372]), .Z(o[8372]) );
  AND U1811 ( .A(p_input[8371]), .B(p_input[18371]), .Z(o[8371]) );
  AND U1812 ( .A(p_input[8370]), .B(p_input[18370]), .Z(o[8370]) );
  AND U1813 ( .A(p_input[836]), .B(p_input[10836]), .Z(o[836]) );
  AND U1814 ( .A(p_input[8369]), .B(p_input[18369]), .Z(o[8369]) );
  AND U1815 ( .A(p_input[8368]), .B(p_input[18368]), .Z(o[8368]) );
  AND U1816 ( .A(p_input[8367]), .B(p_input[18367]), .Z(o[8367]) );
  AND U1817 ( .A(p_input[8366]), .B(p_input[18366]), .Z(o[8366]) );
  AND U1818 ( .A(p_input[8365]), .B(p_input[18365]), .Z(o[8365]) );
  AND U1819 ( .A(p_input[8364]), .B(p_input[18364]), .Z(o[8364]) );
  AND U1820 ( .A(p_input[8363]), .B(p_input[18363]), .Z(o[8363]) );
  AND U1821 ( .A(p_input[8362]), .B(p_input[18362]), .Z(o[8362]) );
  AND U1822 ( .A(p_input[8361]), .B(p_input[18361]), .Z(o[8361]) );
  AND U1823 ( .A(p_input[8360]), .B(p_input[18360]), .Z(o[8360]) );
  AND U1824 ( .A(p_input[835]), .B(p_input[10835]), .Z(o[835]) );
  AND U1825 ( .A(p_input[8359]), .B(p_input[18359]), .Z(o[8359]) );
  AND U1826 ( .A(p_input[8358]), .B(p_input[18358]), .Z(o[8358]) );
  AND U1827 ( .A(p_input[8357]), .B(p_input[18357]), .Z(o[8357]) );
  AND U1828 ( .A(p_input[8356]), .B(p_input[18356]), .Z(o[8356]) );
  AND U1829 ( .A(p_input[8355]), .B(p_input[18355]), .Z(o[8355]) );
  AND U1830 ( .A(p_input[8354]), .B(p_input[18354]), .Z(o[8354]) );
  AND U1831 ( .A(p_input[8353]), .B(p_input[18353]), .Z(o[8353]) );
  AND U1832 ( .A(p_input[8352]), .B(p_input[18352]), .Z(o[8352]) );
  AND U1833 ( .A(p_input[8351]), .B(p_input[18351]), .Z(o[8351]) );
  AND U1834 ( .A(p_input[8350]), .B(p_input[18350]), .Z(o[8350]) );
  AND U1835 ( .A(p_input[834]), .B(p_input[10834]), .Z(o[834]) );
  AND U1836 ( .A(p_input[8349]), .B(p_input[18349]), .Z(o[8349]) );
  AND U1837 ( .A(p_input[8348]), .B(p_input[18348]), .Z(o[8348]) );
  AND U1838 ( .A(p_input[8347]), .B(p_input[18347]), .Z(o[8347]) );
  AND U1839 ( .A(p_input[8346]), .B(p_input[18346]), .Z(o[8346]) );
  AND U1840 ( .A(p_input[8345]), .B(p_input[18345]), .Z(o[8345]) );
  AND U1841 ( .A(p_input[8344]), .B(p_input[18344]), .Z(o[8344]) );
  AND U1842 ( .A(p_input[8343]), .B(p_input[18343]), .Z(o[8343]) );
  AND U1843 ( .A(p_input[8342]), .B(p_input[18342]), .Z(o[8342]) );
  AND U1844 ( .A(p_input[8341]), .B(p_input[18341]), .Z(o[8341]) );
  AND U1845 ( .A(p_input[8340]), .B(p_input[18340]), .Z(o[8340]) );
  AND U1846 ( .A(p_input[833]), .B(p_input[10833]), .Z(o[833]) );
  AND U1847 ( .A(p_input[8339]), .B(p_input[18339]), .Z(o[8339]) );
  AND U1848 ( .A(p_input[8338]), .B(p_input[18338]), .Z(o[8338]) );
  AND U1849 ( .A(p_input[8337]), .B(p_input[18337]), .Z(o[8337]) );
  AND U1850 ( .A(p_input[8336]), .B(p_input[18336]), .Z(o[8336]) );
  AND U1851 ( .A(p_input[8335]), .B(p_input[18335]), .Z(o[8335]) );
  AND U1852 ( .A(p_input[8334]), .B(p_input[18334]), .Z(o[8334]) );
  AND U1853 ( .A(p_input[8333]), .B(p_input[18333]), .Z(o[8333]) );
  AND U1854 ( .A(p_input[8332]), .B(p_input[18332]), .Z(o[8332]) );
  AND U1855 ( .A(p_input[8331]), .B(p_input[18331]), .Z(o[8331]) );
  AND U1856 ( .A(p_input[8330]), .B(p_input[18330]), .Z(o[8330]) );
  AND U1857 ( .A(p_input[832]), .B(p_input[10832]), .Z(o[832]) );
  AND U1858 ( .A(p_input[8329]), .B(p_input[18329]), .Z(o[8329]) );
  AND U1859 ( .A(p_input[8328]), .B(p_input[18328]), .Z(o[8328]) );
  AND U1860 ( .A(p_input[8327]), .B(p_input[18327]), .Z(o[8327]) );
  AND U1861 ( .A(p_input[8326]), .B(p_input[18326]), .Z(o[8326]) );
  AND U1862 ( .A(p_input[8325]), .B(p_input[18325]), .Z(o[8325]) );
  AND U1863 ( .A(p_input[8324]), .B(p_input[18324]), .Z(o[8324]) );
  AND U1864 ( .A(p_input[8323]), .B(p_input[18323]), .Z(o[8323]) );
  AND U1865 ( .A(p_input[8322]), .B(p_input[18322]), .Z(o[8322]) );
  AND U1866 ( .A(p_input[8321]), .B(p_input[18321]), .Z(o[8321]) );
  AND U1867 ( .A(p_input[8320]), .B(p_input[18320]), .Z(o[8320]) );
  AND U1868 ( .A(p_input[831]), .B(p_input[10831]), .Z(o[831]) );
  AND U1869 ( .A(p_input[8319]), .B(p_input[18319]), .Z(o[8319]) );
  AND U1870 ( .A(p_input[8318]), .B(p_input[18318]), .Z(o[8318]) );
  AND U1871 ( .A(p_input[8317]), .B(p_input[18317]), .Z(o[8317]) );
  AND U1872 ( .A(p_input[8316]), .B(p_input[18316]), .Z(o[8316]) );
  AND U1873 ( .A(p_input[8315]), .B(p_input[18315]), .Z(o[8315]) );
  AND U1874 ( .A(p_input[8314]), .B(p_input[18314]), .Z(o[8314]) );
  AND U1875 ( .A(p_input[8313]), .B(p_input[18313]), .Z(o[8313]) );
  AND U1876 ( .A(p_input[8312]), .B(p_input[18312]), .Z(o[8312]) );
  AND U1877 ( .A(p_input[8311]), .B(p_input[18311]), .Z(o[8311]) );
  AND U1878 ( .A(p_input[8310]), .B(p_input[18310]), .Z(o[8310]) );
  AND U1879 ( .A(p_input[830]), .B(p_input[10830]), .Z(o[830]) );
  AND U1880 ( .A(p_input[8309]), .B(p_input[18309]), .Z(o[8309]) );
  AND U1881 ( .A(p_input[8308]), .B(p_input[18308]), .Z(o[8308]) );
  AND U1882 ( .A(p_input[8307]), .B(p_input[18307]), .Z(o[8307]) );
  AND U1883 ( .A(p_input[8306]), .B(p_input[18306]), .Z(o[8306]) );
  AND U1884 ( .A(p_input[8305]), .B(p_input[18305]), .Z(o[8305]) );
  AND U1885 ( .A(p_input[8304]), .B(p_input[18304]), .Z(o[8304]) );
  AND U1886 ( .A(p_input[8303]), .B(p_input[18303]), .Z(o[8303]) );
  AND U1887 ( .A(p_input[8302]), .B(p_input[18302]), .Z(o[8302]) );
  AND U1888 ( .A(p_input[8301]), .B(p_input[18301]), .Z(o[8301]) );
  AND U1889 ( .A(p_input[8300]), .B(p_input[18300]), .Z(o[8300]) );
  AND U1890 ( .A(p_input[82]), .B(p_input[10082]), .Z(o[82]) );
  AND U1891 ( .A(p_input[829]), .B(p_input[10829]), .Z(o[829]) );
  AND U1892 ( .A(p_input[8299]), .B(p_input[18299]), .Z(o[8299]) );
  AND U1893 ( .A(p_input[8298]), .B(p_input[18298]), .Z(o[8298]) );
  AND U1894 ( .A(p_input[8297]), .B(p_input[18297]), .Z(o[8297]) );
  AND U1895 ( .A(p_input[8296]), .B(p_input[18296]), .Z(o[8296]) );
  AND U1896 ( .A(p_input[8295]), .B(p_input[18295]), .Z(o[8295]) );
  AND U1897 ( .A(p_input[8294]), .B(p_input[18294]), .Z(o[8294]) );
  AND U1898 ( .A(p_input[8293]), .B(p_input[18293]), .Z(o[8293]) );
  AND U1899 ( .A(p_input[8292]), .B(p_input[18292]), .Z(o[8292]) );
  AND U1900 ( .A(p_input[8291]), .B(p_input[18291]), .Z(o[8291]) );
  AND U1901 ( .A(p_input[8290]), .B(p_input[18290]), .Z(o[8290]) );
  AND U1902 ( .A(p_input[828]), .B(p_input[10828]), .Z(o[828]) );
  AND U1903 ( .A(p_input[8289]), .B(p_input[18289]), .Z(o[8289]) );
  AND U1904 ( .A(p_input[8288]), .B(p_input[18288]), .Z(o[8288]) );
  AND U1905 ( .A(p_input[8287]), .B(p_input[18287]), .Z(o[8287]) );
  AND U1906 ( .A(p_input[8286]), .B(p_input[18286]), .Z(o[8286]) );
  AND U1907 ( .A(p_input[8285]), .B(p_input[18285]), .Z(o[8285]) );
  AND U1908 ( .A(p_input[8284]), .B(p_input[18284]), .Z(o[8284]) );
  AND U1909 ( .A(p_input[8283]), .B(p_input[18283]), .Z(o[8283]) );
  AND U1910 ( .A(p_input[8282]), .B(p_input[18282]), .Z(o[8282]) );
  AND U1911 ( .A(p_input[8281]), .B(p_input[18281]), .Z(o[8281]) );
  AND U1912 ( .A(p_input[8280]), .B(p_input[18280]), .Z(o[8280]) );
  AND U1913 ( .A(p_input[827]), .B(p_input[10827]), .Z(o[827]) );
  AND U1914 ( .A(p_input[8279]), .B(p_input[18279]), .Z(o[8279]) );
  AND U1915 ( .A(p_input[8278]), .B(p_input[18278]), .Z(o[8278]) );
  AND U1916 ( .A(p_input[8277]), .B(p_input[18277]), .Z(o[8277]) );
  AND U1917 ( .A(p_input[8276]), .B(p_input[18276]), .Z(o[8276]) );
  AND U1918 ( .A(p_input[8275]), .B(p_input[18275]), .Z(o[8275]) );
  AND U1919 ( .A(p_input[8274]), .B(p_input[18274]), .Z(o[8274]) );
  AND U1920 ( .A(p_input[8273]), .B(p_input[18273]), .Z(o[8273]) );
  AND U1921 ( .A(p_input[8272]), .B(p_input[18272]), .Z(o[8272]) );
  AND U1922 ( .A(p_input[8271]), .B(p_input[18271]), .Z(o[8271]) );
  AND U1923 ( .A(p_input[8270]), .B(p_input[18270]), .Z(o[8270]) );
  AND U1924 ( .A(p_input[826]), .B(p_input[10826]), .Z(o[826]) );
  AND U1925 ( .A(p_input[8269]), .B(p_input[18269]), .Z(o[8269]) );
  AND U1926 ( .A(p_input[8268]), .B(p_input[18268]), .Z(o[8268]) );
  AND U1927 ( .A(p_input[8267]), .B(p_input[18267]), .Z(o[8267]) );
  AND U1928 ( .A(p_input[8266]), .B(p_input[18266]), .Z(o[8266]) );
  AND U1929 ( .A(p_input[8265]), .B(p_input[18265]), .Z(o[8265]) );
  AND U1930 ( .A(p_input[8264]), .B(p_input[18264]), .Z(o[8264]) );
  AND U1931 ( .A(p_input[8263]), .B(p_input[18263]), .Z(o[8263]) );
  AND U1932 ( .A(p_input[8262]), .B(p_input[18262]), .Z(o[8262]) );
  AND U1933 ( .A(p_input[8261]), .B(p_input[18261]), .Z(o[8261]) );
  AND U1934 ( .A(p_input[8260]), .B(p_input[18260]), .Z(o[8260]) );
  AND U1935 ( .A(p_input[825]), .B(p_input[10825]), .Z(o[825]) );
  AND U1936 ( .A(p_input[8259]), .B(p_input[18259]), .Z(o[8259]) );
  AND U1937 ( .A(p_input[8258]), .B(p_input[18258]), .Z(o[8258]) );
  AND U1938 ( .A(p_input[8257]), .B(p_input[18257]), .Z(o[8257]) );
  AND U1939 ( .A(p_input[8256]), .B(p_input[18256]), .Z(o[8256]) );
  AND U1940 ( .A(p_input[8255]), .B(p_input[18255]), .Z(o[8255]) );
  AND U1941 ( .A(p_input[8254]), .B(p_input[18254]), .Z(o[8254]) );
  AND U1942 ( .A(p_input[8253]), .B(p_input[18253]), .Z(o[8253]) );
  AND U1943 ( .A(p_input[8252]), .B(p_input[18252]), .Z(o[8252]) );
  AND U1944 ( .A(p_input[8251]), .B(p_input[18251]), .Z(o[8251]) );
  AND U1945 ( .A(p_input[8250]), .B(p_input[18250]), .Z(o[8250]) );
  AND U1946 ( .A(p_input[824]), .B(p_input[10824]), .Z(o[824]) );
  AND U1947 ( .A(p_input[8249]), .B(p_input[18249]), .Z(o[8249]) );
  AND U1948 ( .A(p_input[8248]), .B(p_input[18248]), .Z(o[8248]) );
  AND U1949 ( .A(p_input[8247]), .B(p_input[18247]), .Z(o[8247]) );
  AND U1950 ( .A(p_input[8246]), .B(p_input[18246]), .Z(o[8246]) );
  AND U1951 ( .A(p_input[8245]), .B(p_input[18245]), .Z(o[8245]) );
  AND U1952 ( .A(p_input[8244]), .B(p_input[18244]), .Z(o[8244]) );
  AND U1953 ( .A(p_input[8243]), .B(p_input[18243]), .Z(o[8243]) );
  AND U1954 ( .A(p_input[8242]), .B(p_input[18242]), .Z(o[8242]) );
  AND U1955 ( .A(p_input[8241]), .B(p_input[18241]), .Z(o[8241]) );
  AND U1956 ( .A(p_input[8240]), .B(p_input[18240]), .Z(o[8240]) );
  AND U1957 ( .A(p_input[823]), .B(p_input[10823]), .Z(o[823]) );
  AND U1958 ( .A(p_input[8239]), .B(p_input[18239]), .Z(o[8239]) );
  AND U1959 ( .A(p_input[8238]), .B(p_input[18238]), .Z(o[8238]) );
  AND U1960 ( .A(p_input[8237]), .B(p_input[18237]), .Z(o[8237]) );
  AND U1961 ( .A(p_input[8236]), .B(p_input[18236]), .Z(o[8236]) );
  AND U1962 ( .A(p_input[8235]), .B(p_input[18235]), .Z(o[8235]) );
  AND U1963 ( .A(p_input[8234]), .B(p_input[18234]), .Z(o[8234]) );
  AND U1964 ( .A(p_input[8233]), .B(p_input[18233]), .Z(o[8233]) );
  AND U1965 ( .A(p_input[8232]), .B(p_input[18232]), .Z(o[8232]) );
  AND U1966 ( .A(p_input[8231]), .B(p_input[18231]), .Z(o[8231]) );
  AND U1967 ( .A(p_input[8230]), .B(p_input[18230]), .Z(o[8230]) );
  AND U1968 ( .A(p_input[822]), .B(p_input[10822]), .Z(o[822]) );
  AND U1969 ( .A(p_input[8229]), .B(p_input[18229]), .Z(o[8229]) );
  AND U1970 ( .A(p_input[8228]), .B(p_input[18228]), .Z(o[8228]) );
  AND U1971 ( .A(p_input[8227]), .B(p_input[18227]), .Z(o[8227]) );
  AND U1972 ( .A(p_input[8226]), .B(p_input[18226]), .Z(o[8226]) );
  AND U1973 ( .A(p_input[8225]), .B(p_input[18225]), .Z(o[8225]) );
  AND U1974 ( .A(p_input[8224]), .B(p_input[18224]), .Z(o[8224]) );
  AND U1975 ( .A(p_input[8223]), .B(p_input[18223]), .Z(o[8223]) );
  AND U1976 ( .A(p_input[8222]), .B(p_input[18222]), .Z(o[8222]) );
  AND U1977 ( .A(p_input[8221]), .B(p_input[18221]), .Z(o[8221]) );
  AND U1978 ( .A(p_input[8220]), .B(p_input[18220]), .Z(o[8220]) );
  AND U1979 ( .A(p_input[821]), .B(p_input[10821]), .Z(o[821]) );
  AND U1980 ( .A(p_input[8219]), .B(p_input[18219]), .Z(o[8219]) );
  AND U1981 ( .A(p_input[8218]), .B(p_input[18218]), .Z(o[8218]) );
  AND U1982 ( .A(p_input[8217]), .B(p_input[18217]), .Z(o[8217]) );
  AND U1983 ( .A(p_input[8216]), .B(p_input[18216]), .Z(o[8216]) );
  AND U1984 ( .A(p_input[8215]), .B(p_input[18215]), .Z(o[8215]) );
  AND U1985 ( .A(p_input[8214]), .B(p_input[18214]), .Z(o[8214]) );
  AND U1986 ( .A(p_input[8213]), .B(p_input[18213]), .Z(o[8213]) );
  AND U1987 ( .A(p_input[8212]), .B(p_input[18212]), .Z(o[8212]) );
  AND U1988 ( .A(p_input[8211]), .B(p_input[18211]), .Z(o[8211]) );
  AND U1989 ( .A(p_input[8210]), .B(p_input[18210]), .Z(o[8210]) );
  AND U1990 ( .A(p_input[820]), .B(p_input[10820]), .Z(o[820]) );
  AND U1991 ( .A(p_input[8209]), .B(p_input[18209]), .Z(o[8209]) );
  AND U1992 ( .A(p_input[8208]), .B(p_input[18208]), .Z(o[8208]) );
  AND U1993 ( .A(p_input[8207]), .B(p_input[18207]), .Z(o[8207]) );
  AND U1994 ( .A(p_input[8206]), .B(p_input[18206]), .Z(o[8206]) );
  AND U1995 ( .A(p_input[8205]), .B(p_input[18205]), .Z(o[8205]) );
  AND U1996 ( .A(p_input[8204]), .B(p_input[18204]), .Z(o[8204]) );
  AND U1997 ( .A(p_input[8203]), .B(p_input[18203]), .Z(o[8203]) );
  AND U1998 ( .A(p_input[8202]), .B(p_input[18202]), .Z(o[8202]) );
  AND U1999 ( .A(p_input[8201]), .B(p_input[18201]), .Z(o[8201]) );
  AND U2000 ( .A(p_input[8200]), .B(p_input[18200]), .Z(o[8200]) );
  AND U2001 ( .A(p_input[81]), .B(p_input[10081]), .Z(o[81]) );
  AND U2002 ( .A(p_input[819]), .B(p_input[10819]), .Z(o[819]) );
  AND U2003 ( .A(p_input[8199]), .B(p_input[18199]), .Z(o[8199]) );
  AND U2004 ( .A(p_input[8198]), .B(p_input[18198]), .Z(o[8198]) );
  AND U2005 ( .A(p_input[8197]), .B(p_input[18197]), .Z(o[8197]) );
  AND U2006 ( .A(p_input[8196]), .B(p_input[18196]), .Z(o[8196]) );
  AND U2007 ( .A(p_input[8195]), .B(p_input[18195]), .Z(o[8195]) );
  AND U2008 ( .A(p_input[8194]), .B(p_input[18194]), .Z(o[8194]) );
  AND U2009 ( .A(p_input[8193]), .B(p_input[18193]), .Z(o[8193]) );
  AND U2010 ( .A(p_input[8192]), .B(p_input[18192]), .Z(o[8192]) );
  AND U2011 ( .A(p_input[8191]), .B(p_input[18191]), .Z(o[8191]) );
  AND U2012 ( .A(p_input[8190]), .B(p_input[18190]), .Z(o[8190]) );
  AND U2013 ( .A(p_input[818]), .B(p_input[10818]), .Z(o[818]) );
  AND U2014 ( .A(p_input[8189]), .B(p_input[18189]), .Z(o[8189]) );
  AND U2015 ( .A(p_input[8188]), .B(p_input[18188]), .Z(o[8188]) );
  AND U2016 ( .A(p_input[8187]), .B(p_input[18187]), .Z(o[8187]) );
  AND U2017 ( .A(p_input[8186]), .B(p_input[18186]), .Z(o[8186]) );
  AND U2018 ( .A(p_input[8185]), .B(p_input[18185]), .Z(o[8185]) );
  AND U2019 ( .A(p_input[8184]), .B(p_input[18184]), .Z(o[8184]) );
  AND U2020 ( .A(p_input[8183]), .B(p_input[18183]), .Z(o[8183]) );
  AND U2021 ( .A(p_input[8182]), .B(p_input[18182]), .Z(o[8182]) );
  AND U2022 ( .A(p_input[8181]), .B(p_input[18181]), .Z(o[8181]) );
  AND U2023 ( .A(p_input[8180]), .B(p_input[18180]), .Z(o[8180]) );
  AND U2024 ( .A(p_input[817]), .B(p_input[10817]), .Z(o[817]) );
  AND U2025 ( .A(p_input[8179]), .B(p_input[18179]), .Z(o[8179]) );
  AND U2026 ( .A(p_input[8178]), .B(p_input[18178]), .Z(o[8178]) );
  AND U2027 ( .A(p_input[8177]), .B(p_input[18177]), .Z(o[8177]) );
  AND U2028 ( .A(p_input[8176]), .B(p_input[18176]), .Z(o[8176]) );
  AND U2029 ( .A(p_input[8175]), .B(p_input[18175]), .Z(o[8175]) );
  AND U2030 ( .A(p_input[8174]), .B(p_input[18174]), .Z(o[8174]) );
  AND U2031 ( .A(p_input[8173]), .B(p_input[18173]), .Z(o[8173]) );
  AND U2032 ( .A(p_input[8172]), .B(p_input[18172]), .Z(o[8172]) );
  AND U2033 ( .A(p_input[8171]), .B(p_input[18171]), .Z(o[8171]) );
  AND U2034 ( .A(p_input[8170]), .B(p_input[18170]), .Z(o[8170]) );
  AND U2035 ( .A(p_input[816]), .B(p_input[10816]), .Z(o[816]) );
  AND U2036 ( .A(p_input[8169]), .B(p_input[18169]), .Z(o[8169]) );
  AND U2037 ( .A(p_input[8168]), .B(p_input[18168]), .Z(o[8168]) );
  AND U2038 ( .A(p_input[8167]), .B(p_input[18167]), .Z(o[8167]) );
  AND U2039 ( .A(p_input[8166]), .B(p_input[18166]), .Z(o[8166]) );
  AND U2040 ( .A(p_input[8165]), .B(p_input[18165]), .Z(o[8165]) );
  AND U2041 ( .A(p_input[8164]), .B(p_input[18164]), .Z(o[8164]) );
  AND U2042 ( .A(p_input[8163]), .B(p_input[18163]), .Z(o[8163]) );
  AND U2043 ( .A(p_input[8162]), .B(p_input[18162]), .Z(o[8162]) );
  AND U2044 ( .A(p_input[8161]), .B(p_input[18161]), .Z(o[8161]) );
  AND U2045 ( .A(p_input[8160]), .B(p_input[18160]), .Z(o[8160]) );
  AND U2046 ( .A(p_input[815]), .B(p_input[10815]), .Z(o[815]) );
  AND U2047 ( .A(p_input[8159]), .B(p_input[18159]), .Z(o[8159]) );
  AND U2048 ( .A(p_input[8158]), .B(p_input[18158]), .Z(o[8158]) );
  AND U2049 ( .A(p_input[8157]), .B(p_input[18157]), .Z(o[8157]) );
  AND U2050 ( .A(p_input[8156]), .B(p_input[18156]), .Z(o[8156]) );
  AND U2051 ( .A(p_input[8155]), .B(p_input[18155]), .Z(o[8155]) );
  AND U2052 ( .A(p_input[8154]), .B(p_input[18154]), .Z(o[8154]) );
  AND U2053 ( .A(p_input[8153]), .B(p_input[18153]), .Z(o[8153]) );
  AND U2054 ( .A(p_input[8152]), .B(p_input[18152]), .Z(o[8152]) );
  AND U2055 ( .A(p_input[8151]), .B(p_input[18151]), .Z(o[8151]) );
  AND U2056 ( .A(p_input[8150]), .B(p_input[18150]), .Z(o[8150]) );
  AND U2057 ( .A(p_input[814]), .B(p_input[10814]), .Z(o[814]) );
  AND U2058 ( .A(p_input[8149]), .B(p_input[18149]), .Z(o[8149]) );
  AND U2059 ( .A(p_input[8148]), .B(p_input[18148]), .Z(o[8148]) );
  AND U2060 ( .A(p_input[8147]), .B(p_input[18147]), .Z(o[8147]) );
  AND U2061 ( .A(p_input[8146]), .B(p_input[18146]), .Z(o[8146]) );
  AND U2062 ( .A(p_input[8145]), .B(p_input[18145]), .Z(o[8145]) );
  AND U2063 ( .A(p_input[8144]), .B(p_input[18144]), .Z(o[8144]) );
  AND U2064 ( .A(p_input[8143]), .B(p_input[18143]), .Z(o[8143]) );
  AND U2065 ( .A(p_input[8142]), .B(p_input[18142]), .Z(o[8142]) );
  AND U2066 ( .A(p_input[8141]), .B(p_input[18141]), .Z(o[8141]) );
  AND U2067 ( .A(p_input[8140]), .B(p_input[18140]), .Z(o[8140]) );
  AND U2068 ( .A(p_input[813]), .B(p_input[10813]), .Z(o[813]) );
  AND U2069 ( .A(p_input[8139]), .B(p_input[18139]), .Z(o[8139]) );
  AND U2070 ( .A(p_input[8138]), .B(p_input[18138]), .Z(o[8138]) );
  AND U2071 ( .A(p_input[8137]), .B(p_input[18137]), .Z(o[8137]) );
  AND U2072 ( .A(p_input[8136]), .B(p_input[18136]), .Z(o[8136]) );
  AND U2073 ( .A(p_input[8135]), .B(p_input[18135]), .Z(o[8135]) );
  AND U2074 ( .A(p_input[8134]), .B(p_input[18134]), .Z(o[8134]) );
  AND U2075 ( .A(p_input[8133]), .B(p_input[18133]), .Z(o[8133]) );
  AND U2076 ( .A(p_input[8132]), .B(p_input[18132]), .Z(o[8132]) );
  AND U2077 ( .A(p_input[8131]), .B(p_input[18131]), .Z(o[8131]) );
  AND U2078 ( .A(p_input[8130]), .B(p_input[18130]), .Z(o[8130]) );
  AND U2079 ( .A(p_input[812]), .B(p_input[10812]), .Z(o[812]) );
  AND U2080 ( .A(p_input[8129]), .B(p_input[18129]), .Z(o[8129]) );
  AND U2081 ( .A(p_input[8128]), .B(p_input[18128]), .Z(o[8128]) );
  AND U2082 ( .A(p_input[8127]), .B(p_input[18127]), .Z(o[8127]) );
  AND U2083 ( .A(p_input[8126]), .B(p_input[18126]), .Z(o[8126]) );
  AND U2084 ( .A(p_input[8125]), .B(p_input[18125]), .Z(o[8125]) );
  AND U2085 ( .A(p_input[8124]), .B(p_input[18124]), .Z(o[8124]) );
  AND U2086 ( .A(p_input[8123]), .B(p_input[18123]), .Z(o[8123]) );
  AND U2087 ( .A(p_input[8122]), .B(p_input[18122]), .Z(o[8122]) );
  AND U2088 ( .A(p_input[8121]), .B(p_input[18121]), .Z(o[8121]) );
  AND U2089 ( .A(p_input[8120]), .B(p_input[18120]), .Z(o[8120]) );
  AND U2090 ( .A(p_input[811]), .B(p_input[10811]), .Z(o[811]) );
  AND U2091 ( .A(p_input[8119]), .B(p_input[18119]), .Z(o[8119]) );
  AND U2092 ( .A(p_input[8118]), .B(p_input[18118]), .Z(o[8118]) );
  AND U2093 ( .A(p_input[8117]), .B(p_input[18117]), .Z(o[8117]) );
  AND U2094 ( .A(p_input[8116]), .B(p_input[18116]), .Z(o[8116]) );
  AND U2095 ( .A(p_input[8115]), .B(p_input[18115]), .Z(o[8115]) );
  AND U2096 ( .A(p_input[8114]), .B(p_input[18114]), .Z(o[8114]) );
  AND U2097 ( .A(p_input[8113]), .B(p_input[18113]), .Z(o[8113]) );
  AND U2098 ( .A(p_input[8112]), .B(p_input[18112]), .Z(o[8112]) );
  AND U2099 ( .A(p_input[8111]), .B(p_input[18111]), .Z(o[8111]) );
  AND U2100 ( .A(p_input[8110]), .B(p_input[18110]), .Z(o[8110]) );
  AND U2101 ( .A(p_input[810]), .B(p_input[10810]), .Z(o[810]) );
  AND U2102 ( .A(p_input[8109]), .B(p_input[18109]), .Z(o[8109]) );
  AND U2103 ( .A(p_input[8108]), .B(p_input[18108]), .Z(o[8108]) );
  AND U2104 ( .A(p_input[8107]), .B(p_input[18107]), .Z(o[8107]) );
  AND U2105 ( .A(p_input[8106]), .B(p_input[18106]), .Z(o[8106]) );
  AND U2106 ( .A(p_input[8105]), .B(p_input[18105]), .Z(o[8105]) );
  AND U2107 ( .A(p_input[8104]), .B(p_input[18104]), .Z(o[8104]) );
  AND U2108 ( .A(p_input[8103]), .B(p_input[18103]), .Z(o[8103]) );
  AND U2109 ( .A(p_input[8102]), .B(p_input[18102]), .Z(o[8102]) );
  AND U2110 ( .A(p_input[8101]), .B(p_input[18101]), .Z(o[8101]) );
  AND U2111 ( .A(p_input[8100]), .B(p_input[18100]), .Z(o[8100]) );
  AND U2112 ( .A(p_input[80]), .B(p_input[10080]), .Z(o[80]) );
  AND U2113 ( .A(p_input[809]), .B(p_input[10809]), .Z(o[809]) );
  AND U2114 ( .A(p_input[8099]), .B(p_input[18099]), .Z(o[8099]) );
  AND U2115 ( .A(p_input[8098]), .B(p_input[18098]), .Z(o[8098]) );
  AND U2116 ( .A(p_input[8097]), .B(p_input[18097]), .Z(o[8097]) );
  AND U2117 ( .A(p_input[8096]), .B(p_input[18096]), .Z(o[8096]) );
  AND U2118 ( .A(p_input[8095]), .B(p_input[18095]), .Z(o[8095]) );
  AND U2119 ( .A(p_input[8094]), .B(p_input[18094]), .Z(o[8094]) );
  AND U2120 ( .A(p_input[8093]), .B(p_input[18093]), .Z(o[8093]) );
  AND U2121 ( .A(p_input[8092]), .B(p_input[18092]), .Z(o[8092]) );
  AND U2122 ( .A(p_input[8091]), .B(p_input[18091]), .Z(o[8091]) );
  AND U2123 ( .A(p_input[8090]), .B(p_input[18090]), .Z(o[8090]) );
  AND U2124 ( .A(p_input[808]), .B(p_input[10808]), .Z(o[808]) );
  AND U2125 ( .A(p_input[8089]), .B(p_input[18089]), .Z(o[8089]) );
  AND U2126 ( .A(p_input[8088]), .B(p_input[18088]), .Z(o[8088]) );
  AND U2127 ( .A(p_input[8087]), .B(p_input[18087]), .Z(o[8087]) );
  AND U2128 ( .A(p_input[8086]), .B(p_input[18086]), .Z(o[8086]) );
  AND U2129 ( .A(p_input[8085]), .B(p_input[18085]), .Z(o[8085]) );
  AND U2130 ( .A(p_input[8084]), .B(p_input[18084]), .Z(o[8084]) );
  AND U2131 ( .A(p_input[8083]), .B(p_input[18083]), .Z(o[8083]) );
  AND U2132 ( .A(p_input[8082]), .B(p_input[18082]), .Z(o[8082]) );
  AND U2133 ( .A(p_input[8081]), .B(p_input[18081]), .Z(o[8081]) );
  AND U2134 ( .A(p_input[8080]), .B(p_input[18080]), .Z(o[8080]) );
  AND U2135 ( .A(p_input[807]), .B(p_input[10807]), .Z(o[807]) );
  AND U2136 ( .A(p_input[8079]), .B(p_input[18079]), .Z(o[8079]) );
  AND U2137 ( .A(p_input[8078]), .B(p_input[18078]), .Z(o[8078]) );
  AND U2138 ( .A(p_input[8077]), .B(p_input[18077]), .Z(o[8077]) );
  AND U2139 ( .A(p_input[8076]), .B(p_input[18076]), .Z(o[8076]) );
  AND U2140 ( .A(p_input[8075]), .B(p_input[18075]), .Z(o[8075]) );
  AND U2141 ( .A(p_input[8074]), .B(p_input[18074]), .Z(o[8074]) );
  AND U2142 ( .A(p_input[8073]), .B(p_input[18073]), .Z(o[8073]) );
  AND U2143 ( .A(p_input[8072]), .B(p_input[18072]), .Z(o[8072]) );
  AND U2144 ( .A(p_input[8071]), .B(p_input[18071]), .Z(o[8071]) );
  AND U2145 ( .A(p_input[8070]), .B(p_input[18070]), .Z(o[8070]) );
  AND U2146 ( .A(p_input[806]), .B(p_input[10806]), .Z(o[806]) );
  AND U2147 ( .A(p_input[8069]), .B(p_input[18069]), .Z(o[8069]) );
  AND U2148 ( .A(p_input[8068]), .B(p_input[18068]), .Z(o[8068]) );
  AND U2149 ( .A(p_input[8067]), .B(p_input[18067]), .Z(o[8067]) );
  AND U2150 ( .A(p_input[8066]), .B(p_input[18066]), .Z(o[8066]) );
  AND U2151 ( .A(p_input[8065]), .B(p_input[18065]), .Z(o[8065]) );
  AND U2152 ( .A(p_input[8064]), .B(p_input[18064]), .Z(o[8064]) );
  AND U2153 ( .A(p_input[8063]), .B(p_input[18063]), .Z(o[8063]) );
  AND U2154 ( .A(p_input[8062]), .B(p_input[18062]), .Z(o[8062]) );
  AND U2155 ( .A(p_input[8061]), .B(p_input[18061]), .Z(o[8061]) );
  AND U2156 ( .A(p_input[8060]), .B(p_input[18060]), .Z(o[8060]) );
  AND U2157 ( .A(p_input[805]), .B(p_input[10805]), .Z(o[805]) );
  AND U2158 ( .A(p_input[8059]), .B(p_input[18059]), .Z(o[8059]) );
  AND U2159 ( .A(p_input[8058]), .B(p_input[18058]), .Z(o[8058]) );
  AND U2160 ( .A(p_input[8057]), .B(p_input[18057]), .Z(o[8057]) );
  AND U2161 ( .A(p_input[8056]), .B(p_input[18056]), .Z(o[8056]) );
  AND U2162 ( .A(p_input[8055]), .B(p_input[18055]), .Z(o[8055]) );
  AND U2163 ( .A(p_input[8054]), .B(p_input[18054]), .Z(o[8054]) );
  AND U2164 ( .A(p_input[8053]), .B(p_input[18053]), .Z(o[8053]) );
  AND U2165 ( .A(p_input[8052]), .B(p_input[18052]), .Z(o[8052]) );
  AND U2166 ( .A(p_input[8051]), .B(p_input[18051]), .Z(o[8051]) );
  AND U2167 ( .A(p_input[8050]), .B(p_input[18050]), .Z(o[8050]) );
  AND U2168 ( .A(p_input[804]), .B(p_input[10804]), .Z(o[804]) );
  AND U2169 ( .A(p_input[8049]), .B(p_input[18049]), .Z(o[8049]) );
  AND U2170 ( .A(p_input[8048]), .B(p_input[18048]), .Z(o[8048]) );
  AND U2171 ( .A(p_input[8047]), .B(p_input[18047]), .Z(o[8047]) );
  AND U2172 ( .A(p_input[8046]), .B(p_input[18046]), .Z(o[8046]) );
  AND U2173 ( .A(p_input[8045]), .B(p_input[18045]), .Z(o[8045]) );
  AND U2174 ( .A(p_input[8044]), .B(p_input[18044]), .Z(o[8044]) );
  AND U2175 ( .A(p_input[8043]), .B(p_input[18043]), .Z(o[8043]) );
  AND U2176 ( .A(p_input[8042]), .B(p_input[18042]), .Z(o[8042]) );
  AND U2177 ( .A(p_input[8041]), .B(p_input[18041]), .Z(o[8041]) );
  AND U2178 ( .A(p_input[8040]), .B(p_input[18040]), .Z(o[8040]) );
  AND U2179 ( .A(p_input[803]), .B(p_input[10803]), .Z(o[803]) );
  AND U2180 ( .A(p_input[8039]), .B(p_input[18039]), .Z(o[8039]) );
  AND U2181 ( .A(p_input[8038]), .B(p_input[18038]), .Z(o[8038]) );
  AND U2182 ( .A(p_input[8037]), .B(p_input[18037]), .Z(o[8037]) );
  AND U2183 ( .A(p_input[8036]), .B(p_input[18036]), .Z(o[8036]) );
  AND U2184 ( .A(p_input[8035]), .B(p_input[18035]), .Z(o[8035]) );
  AND U2185 ( .A(p_input[8034]), .B(p_input[18034]), .Z(o[8034]) );
  AND U2186 ( .A(p_input[8033]), .B(p_input[18033]), .Z(o[8033]) );
  AND U2187 ( .A(p_input[8032]), .B(p_input[18032]), .Z(o[8032]) );
  AND U2188 ( .A(p_input[8031]), .B(p_input[18031]), .Z(o[8031]) );
  AND U2189 ( .A(p_input[8030]), .B(p_input[18030]), .Z(o[8030]) );
  AND U2190 ( .A(p_input[802]), .B(p_input[10802]), .Z(o[802]) );
  AND U2191 ( .A(p_input[8029]), .B(p_input[18029]), .Z(o[8029]) );
  AND U2192 ( .A(p_input[8028]), .B(p_input[18028]), .Z(o[8028]) );
  AND U2193 ( .A(p_input[8027]), .B(p_input[18027]), .Z(o[8027]) );
  AND U2194 ( .A(p_input[8026]), .B(p_input[18026]), .Z(o[8026]) );
  AND U2195 ( .A(p_input[8025]), .B(p_input[18025]), .Z(o[8025]) );
  AND U2196 ( .A(p_input[8024]), .B(p_input[18024]), .Z(o[8024]) );
  AND U2197 ( .A(p_input[8023]), .B(p_input[18023]), .Z(o[8023]) );
  AND U2198 ( .A(p_input[8022]), .B(p_input[18022]), .Z(o[8022]) );
  AND U2199 ( .A(p_input[8021]), .B(p_input[18021]), .Z(o[8021]) );
  AND U2200 ( .A(p_input[8020]), .B(p_input[18020]), .Z(o[8020]) );
  AND U2201 ( .A(p_input[801]), .B(p_input[10801]), .Z(o[801]) );
  AND U2202 ( .A(p_input[8019]), .B(p_input[18019]), .Z(o[8019]) );
  AND U2203 ( .A(p_input[8018]), .B(p_input[18018]), .Z(o[8018]) );
  AND U2204 ( .A(p_input[8017]), .B(p_input[18017]), .Z(o[8017]) );
  AND U2205 ( .A(p_input[8016]), .B(p_input[18016]), .Z(o[8016]) );
  AND U2206 ( .A(p_input[8015]), .B(p_input[18015]), .Z(o[8015]) );
  AND U2207 ( .A(p_input[8014]), .B(p_input[18014]), .Z(o[8014]) );
  AND U2208 ( .A(p_input[8013]), .B(p_input[18013]), .Z(o[8013]) );
  AND U2209 ( .A(p_input[8012]), .B(p_input[18012]), .Z(o[8012]) );
  AND U2210 ( .A(p_input[8011]), .B(p_input[18011]), .Z(o[8011]) );
  AND U2211 ( .A(p_input[8010]), .B(p_input[18010]), .Z(o[8010]) );
  AND U2212 ( .A(p_input[800]), .B(p_input[10800]), .Z(o[800]) );
  AND U2213 ( .A(p_input[8009]), .B(p_input[18009]), .Z(o[8009]) );
  AND U2214 ( .A(p_input[8008]), .B(p_input[18008]), .Z(o[8008]) );
  AND U2215 ( .A(p_input[8007]), .B(p_input[18007]), .Z(o[8007]) );
  AND U2216 ( .A(p_input[8006]), .B(p_input[18006]), .Z(o[8006]) );
  AND U2217 ( .A(p_input[8005]), .B(p_input[18005]), .Z(o[8005]) );
  AND U2218 ( .A(p_input[8004]), .B(p_input[18004]), .Z(o[8004]) );
  AND U2219 ( .A(p_input[8003]), .B(p_input[18003]), .Z(o[8003]) );
  AND U2220 ( .A(p_input[8002]), .B(p_input[18002]), .Z(o[8002]) );
  AND U2221 ( .A(p_input[8001]), .B(p_input[18001]), .Z(o[8001]) );
  AND U2222 ( .A(p_input[8000]), .B(p_input[18000]), .Z(o[8000]) );
  AND U2223 ( .A(p_input[7]), .B(p_input[10007]), .Z(o[7]) );
  AND U2224 ( .A(p_input[79]), .B(p_input[10079]), .Z(o[79]) );
  AND U2225 ( .A(p_input[799]), .B(p_input[10799]), .Z(o[799]) );
  AND U2226 ( .A(p_input[7999]), .B(p_input[17999]), .Z(o[7999]) );
  AND U2227 ( .A(p_input[7998]), .B(p_input[17998]), .Z(o[7998]) );
  AND U2228 ( .A(p_input[7997]), .B(p_input[17997]), .Z(o[7997]) );
  AND U2229 ( .A(p_input[7996]), .B(p_input[17996]), .Z(o[7996]) );
  AND U2230 ( .A(p_input[7995]), .B(p_input[17995]), .Z(o[7995]) );
  AND U2231 ( .A(p_input[7994]), .B(p_input[17994]), .Z(o[7994]) );
  AND U2232 ( .A(p_input[7993]), .B(p_input[17993]), .Z(o[7993]) );
  AND U2233 ( .A(p_input[7992]), .B(p_input[17992]), .Z(o[7992]) );
  AND U2234 ( .A(p_input[7991]), .B(p_input[17991]), .Z(o[7991]) );
  AND U2235 ( .A(p_input[7990]), .B(p_input[17990]), .Z(o[7990]) );
  AND U2236 ( .A(p_input[798]), .B(p_input[10798]), .Z(o[798]) );
  AND U2237 ( .A(p_input[7989]), .B(p_input[17989]), .Z(o[7989]) );
  AND U2238 ( .A(p_input[7988]), .B(p_input[17988]), .Z(o[7988]) );
  AND U2239 ( .A(p_input[7987]), .B(p_input[17987]), .Z(o[7987]) );
  AND U2240 ( .A(p_input[7986]), .B(p_input[17986]), .Z(o[7986]) );
  AND U2241 ( .A(p_input[7985]), .B(p_input[17985]), .Z(o[7985]) );
  AND U2242 ( .A(p_input[7984]), .B(p_input[17984]), .Z(o[7984]) );
  AND U2243 ( .A(p_input[7983]), .B(p_input[17983]), .Z(o[7983]) );
  AND U2244 ( .A(p_input[7982]), .B(p_input[17982]), .Z(o[7982]) );
  AND U2245 ( .A(p_input[7981]), .B(p_input[17981]), .Z(o[7981]) );
  AND U2246 ( .A(p_input[7980]), .B(p_input[17980]), .Z(o[7980]) );
  AND U2247 ( .A(p_input[797]), .B(p_input[10797]), .Z(o[797]) );
  AND U2248 ( .A(p_input[7979]), .B(p_input[17979]), .Z(o[7979]) );
  AND U2249 ( .A(p_input[7978]), .B(p_input[17978]), .Z(o[7978]) );
  AND U2250 ( .A(p_input[7977]), .B(p_input[17977]), .Z(o[7977]) );
  AND U2251 ( .A(p_input[7976]), .B(p_input[17976]), .Z(o[7976]) );
  AND U2252 ( .A(p_input[7975]), .B(p_input[17975]), .Z(o[7975]) );
  AND U2253 ( .A(p_input[7974]), .B(p_input[17974]), .Z(o[7974]) );
  AND U2254 ( .A(p_input[7973]), .B(p_input[17973]), .Z(o[7973]) );
  AND U2255 ( .A(p_input[7972]), .B(p_input[17972]), .Z(o[7972]) );
  AND U2256 ( .A(p_input[7971]), .B(p_input[17971]), .Z(o[7971]) );
  AND U2257 ( .A(p_input[7970]), .B(p_input[17970]), .Z(o[7970]) );
  AND U2258 ( .A(p_input[796]), .B(p_input[10796]), .Z(o[796]) );
  AND U2259 ( .A(p_input[7969]), .B(p_input[17969]), .Z(o[7969]) );
  AND U2260 ( .A(p_input[7968]), .B(p_input[17968]), .Z(o[7968]) );
  AND U2261 ( .A(p_input[7967]), .B(p_input[17967]), .Z(o[7967]) );
  AND U2262 ( .A(p_input[7966]), .B(p_input[17966]), .Z(o[7966]) );
  AND U2263 ( .A(p_input[7965]), .B(p_input[17965]), .Z(o[7965]) );
  AND U2264 ( .A(p_input[7964]), .B(p_input[17964]), .Z(o[7964]) );
  AND U2265 ( .A(p_input[7963]), .B(p_input[17963]), .Z(o[7963]) );
  AND U2266 ( .A(p_input[7962]), .B(p_input[17962]), .Z(o[7962]) );
  AND U2267 ( .A(p_input[7961]), .B(p_input[17961]), .Z(o[7961]) );
  AND U2268 ( .A(p_input[7960]), .B(p_input[17960]), .Z(o[7960]) );
  AND U2269 ( .A(p_input[795]), .B(p_input[10795]), .Z(o[795]) );
  AND U2270 ( .A(p_input[7959]), .B(p_input[17959]), .Z(o[7959]) );
  AND U2271 ( .A(p_input[7958]), .B(p_input[17958]), .Z(o[7958]) );
  AND U2272 ( .A(p_input[7957]), .B(p_input[17957]), .Z(o[7957]) );
  AND U2273 ( .A(p_input[7956]), .B(p_input[17956]), .Z(o[7956]) );
  AND U2274 ( .A(p_input[7955]), .B(p_input[17955]), .Z(o[7955]) );
  AND U2275 ( .A(p_input[7954]), .B(p_input[17954]), .Z(o[7954]) );
  AND U2276 ( .A(p_input[7953]), .B(p_input[17953]), .Z(o[7953]) );
  AND U2277 ( .A(p_input[7952]), .B(p_input[17952]), .Z(o[7952]) );
  AND U2278 ( .A(p_input[7951]), .B(p_input[17951]), .Z(o[7951]) );
  AND U2279 ( .A(p_input[7950]), .B(p_input[17950]), .Z(o[7950]) );
  AND U2280 ( .A(p_input[794]), .B(p_input[10794]), .Z(o[794]) );
  AND U2281 ( .A(p_input[7949]), .B(p_input[17949]), .Z(o[7949]) );
  AND U2282 ( .A(p_input[7948]), .B(p_input[17948]), .Z(o[7948]) );
  AND U2283 ( .A(p_input[7947]), .B(p_input[17947]), .Z(o[7947]) );
  AND U2284 ( .A(p_input[7946]), .B(p_input[17946]), .Z(o[7946]) );
  AND U2285 ( .A(p_input[7945]), .B(p_input[17945]), .Z(o[7945]) );
  AND U2286 ( .A(p_input[7944]), .B(p_input[17944]), .Z(o[7944]) );
  AND U2287 ( .A(p_input[7943]), .B(p_input[17943]), .Z(o[7943]) );
  AND U2288 ( .A(p_input[7942]), .B(p_input[17942]), .Z(o[7942]) );
  AND U2289 ( .A(p_input[7941]), .B(p_input[17941]), .Z(o[7941]) );
  AND U2290 ( .A(p_input[7940]), .B(p_input[17940]), .Z(o[7940]) );
  AND U2291 ( .A(p_input[793]), .B(p_input[10793]), .Z(o[793]) );
  AND U2292 ( .A(p_input[7939]), .B(p_input[17939]), .Z(o[7939]) );
  AND U2293 ( .A(p_input[7938]), .B(p_input[17938]), .Z(o[7938]) );
  AND U2294 ( .A(p_input[7937]), .B(p_input[17937]), .Z(o[7937]) );
  AND U2295 ( .A(p_input[7936]), .B(p_input[17936]), .Z(o[7936]) );
  AND U2296 ( .A(p_input[7935]), .B(p_input[17935]), .Z(o[7935]) );
  AND U2297 ( .A(p_input[7934]), .B(p_input[17934]), .Z(o[7934]) );
  AND U2298 ( .A(p_input[7933]), .B(p_input[17933]), .Z(o[7933]) );
  AND U2299 ( .A(p_input[7932]), .B(p_input[17932]), .Z(o[7932]) );
  AND U2300 ( .A(p_input[7931]), .B(p_input[17931]), .Z(o[7931]) );
  AND U2301 ( .A(p_input[7930]), .B(p_input[17930]), .Z(o[7930]) );
  AND U2302 ( .A(p_input[792]), .B(p_input[10792]), .Z(o[792]) );
  AND U2303 ( .A(p_input[7929]), .B(p_input[17929]), .Z(o[7929]) );
  AND U2304 ( .A(p_input[7928]), .B(p_input[17928]), .Z(o[7928]) );
  AND U2305 ( .A(p_input[7927]), .B(p_input[17927]), .Z(o[7927]) );
  AND U2306 ( .A(p_input[7926]), .B(p_input[17926]), .Z(o[7926]) );
  AND U2307 ( .A(p_input[7925]), .B(p_input[17925]), .Z(o[7925]) );
  AND U2308 ( .A(p_input[7924]), .B(p_input[17924]), .Z(o[7924]) );
  AND U2309 ( .A(p_input[7923]), .B(p_input[17923]), .Z(o[7923]) );
  AND U2310 ( .A(p_input[7922]), .B(p_input[17922]), .Z(o[7922]) );
  AND U2311 ( .A(p_input[7921]), .B(p_input[17921]), .Z(o[7921]) );
  AND U2312 ( .A(p_input[7920]), .B(p_input[17920]), .Z(o[7920]) );
  AND U2313 ( .A(p_input[791]), .B(p_input[10791]), .Z(o[791]) );
  AND U2314 ( .A(p_input[7919]), .B(p_input[17919]), .Z(o[7919]) );
  AND U2315 ( .A(p_input[7918]), .B(p_input[17918]), .Z(o[7918]) );
  AND U2316 ( .A(p_input[7917]), .B(p_input[17917]), .Z(o[7917]) );
  AND U2317 ( .A(p_input[7916]), .B(p_input[17916]), .Z(o[7916]) );
  AND U2318 ( .A(p_input[7915]), .B(p_input[17915]), .Z(o[7915]) );
  AND U2319 ( .A(p_input[7914]), .B(p_input[17914]), .Z(o[7914]) );
  AND U2320 ( .A(p_input[7913]), .B(p_input[17913]), .Z(o[7913]) );
  AND U2321 ( .A(p_input[7912]), .B(p_input[17912]), .Z(o[7912]) );
  AND U2322 ( .A(p_input[7911]), .B(p_input[17911]), .Z(o[7911]) );
  AND U2323 ( .A(p_input[7910]), .B(p_input[17910]), .Z(o[7910]) );
  AND U2324 ( .A(p_input[790]), .B(p_input[10790]), .Z(o[790]) );
  AND U2325 ( .A(p_input[7909]), .B(p_input[17909]), .Z(o[7909]) );
  AND U2326 ( .A(p_input[7908]), .B(p_input[17908]), .Z(o[7908]) );
  AND U2327 ( .A(p_input[7907]), .B(p_input[17907]), .Z(o[7907]) );
  AND U2328 ( .A(p_input[7906]), .B(p_input[17906]), .Z(o[7906]) );
  AND U2329 ( .A(p_input[7905]), .B(p_input[17905]), .Z(o[7905]) );
  AND U2330 ( .A(p_input[7904]), .B(p_input[17904]), .Z(o[7904]) );
  AND U2331 ( .A(p_input[7903]), .B(p_input[17903]), .Z(o[7903]) );
  AND U2332 ( .A(p_input[7902]), .B(p_input[17902]), .Z(o[7902]) );
  AND U2333 ( .A(p_input[7901]), .B(p_input[17901]), .Z(o[7901]) );
  AND U2334 ( .A(p_input[7900]), .B(p_input[17900]), .Z(o[7900]) );
  AND U2335 ( .A(p_input[78]), .B(p_input[10078]), .Z(o[78]) );
  AND U2336 ( .A(p_input[789]), .B(p_input[10789]), .Z(o[789]) );
  AND U2337 ( .A(p_input[7899]), .B(p_input[17899]), .Z(o[7899]) );
  AND U2338 ( .A(p_input[7898]), .B(p_input[17898]), .Z(o[7898]) );
  AND U2339 ( .A(p_input[7897]), .B(p_input[17897]), .Z(o[7897]) );
  AND U2340 ( .A(p_input[7896]), .B(p_input[17896]), .Z(o[7896]) );
  AND U2341 ( .A(p_input[7895]), .B(p_input[17895]), .Z(o[7895]) );
  AND U2342 ( .A(p_input[7894]), .B(p_input[17894]), .Z(o[7894]) );
  AND U2343 ( .A(p_input[7893]), .B(p_input[17893]), .Z(o[7893]) );
  AND U2344 ( .A(p_input[7892]), .B(p_input[17892]), .Z(o[7892]) );
  AND U2345 ( .A(p_input[7891]), .B(p_input[17891]), .Z(o[7891]) );
  AND U2346 ( .A(p_input[7890]), .B(p_input[17890]), .Z(o[7890]) );
  AND U2347 ( .A(p_input[788]), .B(p_input[10788]), .Z(o[788]) );
  AND U2348 ( .A(p_input[7889]), .B(p_input[17889]), .Z(o[7889]) );
  AND U2349 ( .A(p_input[7888]), .B(p_input[17888]), .Z(o[7888]) );
  AND U2350 ( .A(p_input[7887]), .B(p_input[17887]), .Z(o[7887]) );
  AND U2351 ( .A(p_input[7886]), .B(p_input[17886]), .Z(o[7886]) );
  AND U2352 ( .A(p_input[7885]), .B(p_input[17885]), .Z(o[7885]) );
  AND U2353 ( .A(p_input[7884]), .B(p_input[17884]), .Z(o[7884]) );
  AND U2354 ( .A(p_input[7883]), .B(p_input[17883]), .Z(o[7883]) );
  AND U2355 ( .A(p_input[7882]), .B(p_input[17882]), .Z(o[7882]) );
  AND U2356 ( .A(p_input[7881]), .B(p_input[17881]), .Z(o[7881]) );
  AND U2357 ( .A(p_input[7880]), .B(p_input[17880]), .Z(o[7880]) );
  AND U2358 ( .A(p_input[787]), .B(p_input[10787]), .Z(o[787]) );
  AND U2359 ( .A(p_input[7879]), .B(p_input[17879]), .Z(o[7879]) );
  AND U2360 ( .A(p_input[7878]), .B(p_input[17878]), .Z(o[7878]) );
  AND U2361 ( .A(p_input[7877]), .B(p_input[17877]), .Z(o[7877]) );
  AND U2362 ( .A(p_input[7876]), .B(p_input[17876]), .Z(o[7876]) );
  AND U2363 ( .A(p_input[7875]), .B(p_input[17875]), .Z(o[7875]) );
  AND U2364 ( .A(p_input[7874]), .B(p_input[17874]), .Z(o[7874]) );
  AND U2365 ( .A(p_input[7873]), .B(p_input[17873]), .Z(o[7873]) );
  AND U2366 ( .A(p_input[7872]), .B(p_input[17872]), .Z(o[7872]) );
  AND U2367 ( .A(p_input[7871]), .B(p_input[17871]), .Z(o[7871]) );
  AND U2368 ( .A(p_input[7870]), .B(p_input[17870]), .Z(o[7870]) );
  AND U2369 ( .A(p_input[786]), .B(p_input[10786]), .Z(o[786]) );
  AND U2370 ( .A(p_input[7869]), .B(p_input[17869]), .Z(o[7869]) );
  AND U2371 ( .A(p_input[7868]), .B(p_input[17868]), .Z(o[7868]) );
  AND U2372 ( .A(p_input[7867]), .B(p_input[17867]), .Z(o[7867]) );
  AND U2373 ( .A(p_input[7866]), .B(p_input[17866]), .Z(o[7866]) );
  AND U2374 ( .A(p_input[7865]), .B(p_input[17865]), .Z(o[7865]) );
  AND U2375 ( .A(p_input[7864]), .B(p_input[17864]), .Z(o[7864]) );
  AND U2376 ( .A(p_input[7863]), .B(p_input[17863]), .Z(o[7863]) );
  AND U2377 ( .A(p_input[7862]), .B(p_input[17862]), .Z(o[7862]) );
  AND U2378 ( .A(p_input[7861]), .B(p_input[17861]), .Z(o[7861]) );
  AND U2379 ( .A(p_input[7860]), .B(p_input[17860]), .Z(o[7860]) );
  AND U2380 ( .A(p_input[785]), .B(p_input[10785]), .Z(o[785]) );
  AND U2381 ( .A(p_input[7859]), .B(p_input[17859]), .Z(o[7859]) );
  AND U2382 ( .A(p_input[7858]), .B(p_input[17858]), .Z(o[7858]) );
  AND U2383 ( .A(p_input[7857]), .B(p_input[17857]), .Z(o[7857]) );
  AND U2384 ( .A(p_input[7856]), .B(p_input[17856]), .Z(o[7856]) );
  AND U2385 ( .A(p_input[7855]), .B(p_input[17855]), .Z(o[7855]) );
  AND U2386 ( .A(p_input[7854]), .B(p_input[17854]), .Z(o[7854]) );
  AND U2387 ( .A(p_input[7853]), .B(p_input[17853]), .Z(o[7853]) );
  AND U2388 ( .A(p_input[7852]), .B(p_input[17852]), .Z(o[7852]) );
  AND U2389 ( .A(p_input[7851]), .B(p_input[17851]), .Z(o[7851]) );
  AND U2390 ( .A(p_input[7850]), .B(p_input[17850]), .Z(o[7850]) );
  AND U2391 ( .A(p_input[784]), .B(p_input[10784]), .Z(o[784]) );
  AND U2392 ( .A(p_input[7849]), .B(p_input[17849]), .Z(o[7849]) );
  AND U2393 ( .A(p_input[7848]), .B(p_input[17848]), .Z(o[7848]) );
  AND U2394 ( .A(p_input[7847]), .B(p_input[17847]), .Z(o[7847]) );
  AND U2395 ( .A(p_input[7846]), .B(p_input[17846]), .Z(o[7846]) );
  AND U2396 ( .A(p_input[7845]), .B(p_input[17845]), .Z(o[7845]) );
  AND U2397 ( .A(p_input[7844]), .B(p_input[17844]), .Z(o[7844]) );
  AND U2398 ( .A(p_input[7843]), .B(p_input[17843]), .Z(o[7843]) );
  AND U2399 ( .A(p_input[7842]), .B(p_input[17842]), .Z(o[7842]) );
  AND U2400 ( .A(p_input[7841]), .B(p_input[17841]), .Z(o[7841]) );
  AND U2401 ( .A(p_input[7840]), .B(p_input[17840]), .Z(o[7840]) );
  AND U2402 ( .A(p_input[783]), .B(p_input[10783]), .Z(o[783]) );
  AND U2403 ( .A(p_input[7839]), .B(p_input[17839]), .Z(o[7839]) );
  AND U2404 ( .A(p_input[7838]), .B(p_input[17838]), .Z(o[7838]) );
  AND U2405 ( .A(p_input[7837]), .B(p_input[17837]), .Z(o[7837]) );
  AND U2406 ( .A(p_input[7836]), .B(p_input[17836]), .Z(o[7836]) );
  AND U2407 ( .A(p_input[7835]), .B(p_input[17835]), .Z(o[7835]) );
  AND U2408 ( .A(p_input[7834]), .B(p_input[17834]), .Z(o[7834]) );
  AND U2409 ( .A(p_input[7833]), .B(p_input[17833]), .Z(o[7833]) );
  AND U2410 ( .A(p_input[7832]), .B(p_input[17832]), .Z(o[7832]) );
  AND U2411 ( .A(p_input[7831]), .B(p_input[17831]), .Z(o[7831]) );
  AND U2412 ( .A(p_input[7830]), .B(p_input[17830]), .Z(o[7830]) );
  AND U2413 ( .A(p_input[782]), .B(p_input[10782]), .Z(o[782]) );
  AND U2414 ( .A(p_input[7829]), .B(p_input[17829]), .Z(o[7829]) );
  AND U2415 ( .A(p_input[7828]), .B(p_input[17828]), .Z(o[7828]) );
  AND U2416 ( .A(p_input[7827]), .B(p_input[17827]), .Z(o[7827]) );
  AND U2417 ( .A(p_input[7826]), .B(p_input[17826]), .Z(o[7826]) );
  AND U2418 ( .A(p_input[7825]), .B(p_input[17825]), .Z(o[7825]) );
  AND U2419 ( .A(p_input[7824]), .B(p_input[17824]), .Z(o[7824]) );
  AND U2420 ( .A(p_input[7823]), .B(p_input[17823]), .Z(o[7823]) );
  AND U2421 ( .A(p_input[7822]), .B(p_input[17822]), .Z(o[7822]) );
  AND U2422 ( .A(p_input[7821]), .B(p_input[17821]), .Z(o[7821]) );
  AND U2423 ( .A(p_input[7820]), .B(p_input[17820]), .Z(o[7820]) );
  AND U2424 ( .A(p_input[781]), .B(p_input[10781]), .Z(o[781]) );
  AND U2425 ( .A(p_input[7819]), .B(p_input[17819]), .Z(o[7819]) );
  AND U2426 ( .A(p_input[7818]), .B(p_input[17818]), .Z(o[7818]) );
  AND U2427 ( .A(p_input[7817]), .B(p_input[17817]), .Z(o[7817]) );
  AND U2428 ( .A(p_input[7816]), .B(p_input[17816]), .Z(o[7816]) );
  AND U2429 ( .A(p_input[7815]), .B(p_input[17815]), .Z(o[7815]) );
  AND U2430 ( .A(p_input[7814]), .B(p_input[17814]), .Z(o[7814]) );
  AND U2431 ( .A(p_input[7813]), .B(p_input[17813]), .Z(o[7813]) );
  AND U2432 ( .A(p_input[7812]), .B(p_input[17812]), .Z(o[7812]) );
  AND U2433 ( .A(p_input[7811]), .B(p_input[17811]), .Z(o[7811]) );
  AND U2434 ( .A(p_input[7810]), .B(p_input[17810]), .Z(o[7810]) );
  AND U2435 ( .A(p_input[780]), .B(p_input[10780]), .Z(o[780]) );
  AND U2436 ( .A(p_input[7809]), .B(p_input[17809]), .Z(o[7809]) );
  AND U2437 ( .A(p_input[7808]), .B(p_input[17808]), .Z(o[7808]) );
  AND U2438 ( .A(p_input[7807]), .B(p_input[17807]), .Z(o[7807]) );
  AND U2439 ( .A(p_input[7806]), .B(p_input[17806]), .Z(o[7806]) );
  AND U2440 ( .A(p_input[7805]), .B(p_input[17805]), .Z(o[7805]) );
  AND U2441 ( .A(p_input[7804]), .B(p_input[17804]), .Z(o[7804]) );
  AND U2442 ( .A(p_input[7803]), .B(p_input[17803]), .Z(o[7803]) );
  AND U2443 ( .A(p_input[7802]), .B(p_input[17802]), .Z(o[7802]) );
  AND U2444 ( .A(p_input[7801]), .B(p_input[17801]), .Z(o[7801]) );
  AND U2445 ( .A(p_input[7800]), .B(p_input[17800]), .Z(o[7800]) );
  AND U2446 ( .A(p_input[77]), .B(p_input[10077]), .Z(o[77]) );
  AND U2447 ( .A(p_input[779]), .B(p_input[10779]), .Z(o[779]) );
  AND U2448 ( .A(p_input[7799]), .B(p_input[17799]), .Z(o[7799]) );
  AND U2449 ( .A(p_input[7798]), .B(p_input[17798]), .Z(o[7798]) );
  AND U2450 ( .A(p_input[7797]), .B(p_input[17797]), .Z(o[7797]) );
  AND U2451 ( .A(p_input[7796]), .B(p_input[17796]), .Z(o[7796]) );
  AND U2452 ( .A(p_input[7795]), .B(p_input[17795]), .Z(o[7795]) );
  AND U2453 ( .A(p_input[7794]), .B(p_input[17794]), .Z(o[7794]) );
  AND U2454 ( .A(p_input[7793]), .B(p_input[17793]), .Z(o[7793]) );
  AND U2455 ( .A(p_input[7792]), .B(p_input[17792]), .Z(o[7792]) );
  AND U2456 ( .A(p_input[7791]), .B(p_input[17791]), .Z(o[7791]) );
  AND U2457 ( .A(p_input[7790]), .B(p_input[17790]), .Z(o[7790]) );
  AND U2458 ( .A(p_input[778]), .B(p_input[10778]), .Z(o[778]) );
  AND U2459 ( .A(p_input[7789]), .B(p_input[17789]), .Z(o[7789]) );
  AND U2460 ( .A(p_input[7788]), .B(p_input[17788]), .Z(o[7788]) );
  AND U2461 ( .A(p_input[7787]), .B(p_input[17787]), .Z(o[7787]) );
  AND U2462 ( .A(p_input[7786]), .B(p_input[17786]), .Z(o[7786]) );
  AND U2463 ( .A(p_input[7785]), .B(p_input[17785]), .Z(o[7785]) );
  AND U2464 ( .A(p_input[7784]), .B(p_input[17784]), .Z(o[7784]) );
  AND U2465 ( .A(p_input[7783]), .B(p_input[17783]), .Z(o[7783]) );
  AND U2466 ( .A(p_input[7782]), .B(p_input[17782]), .Z(o[7782]) );
  AND U2467 ( .A(p_input[7781]), .B(p_input[17781]), .Z(o[7781]) );
  AND U2468 ( .A(p_input[7780]), .B(p_input[17780]), .Z(o[7780]) );
  AND U2469 ( .A(p_input[777]), .B(p_input[10777]), .Z(o[777]) );
  AND U2470 ( .A(p_input[7779]), .B(p_input[17779]), .Z(o[7779]) );
  AND U2471 ( .A(p_input[7778]), .B(p_input[17778]), .Z(o[7778]) );
  AND U2472 ( .A(p_input[7777]), .B(p_input[17777]), .Z(o[7777]) );
  AND U2473 ( .A(p_input[7776]), .B(p_input[17776]), .Z(o[7776]) );
  AND U2474 ( .A(p_input[7775]), .B(p_input[17775]), .Z(o[7775]) );
  AND U2475 ( .A(p_input[7774]), .B(p_input[17774]), .Z(o[7774]) );
  AND U2476 ( .A(p_input[7773]), .B(p_input[17773]), .Z(o[7773]) );
  AND U2477 ( .A(p_input[7772]), .B(p_input[17772]), .Z(o[7772]) );
  AND U2478 ( .A(p_input[7771]), .B(p_input[17771]), .Z(o[7771]) );
  AND U2479 ( .A(p_input[7770]), .B(p_input[17770]), .Z(o[7770]) );
  AND U2480 ( .A(p_input[776]), .B(p_input[10776]), .Z(o[776]) );
  AND U2481 ( .A(p_input[7769]), .B(p_input[17769]), .Z(o[7769]) );
  AND U2482 ( .A(p_input[7768]), .B(p_input[17768]), .Z(o[7768]) );
  AND U2483 ( .A(p_input[7767]), .B(p_input[17767]), .Z(o[7767]) );
  AND U2484 ( .A(p_input[7766]), .B(p_input[17766]), .Z(o[7766]) );
  AND U2485 ( .A(p_input[7765]), .B(p_input[17765]), .Z(o[7765]) );
  AND U2486 ( .A(p_input[7764]), .B(p_input[17764]), .Z(o[7764]) );
  AND U2487 ( .A(p_input[7763]), .B(p_input[17763]), .Z(o[7763]) );
  AND U2488 ( .A(p_input[7762]), .B(p_input[17762]), .Z(o[7762]) );
  AND U2489 ( .A(p_input[7761]), .B(p_input[17761]), .Z(o[7761]) );
  AND U2490 ( .A(p_input[7760]), .B(p_input[17760]), .Z(o[7760]) );
  AND U2491 ( .A(p_input[775]), .B(p_input[10775]), .Z(o[775]) );
  AND U2492 ( .A(p_input[7759]), .B(p_input[17759]), .Z(o[7759]) );
  AND U2493 ( .A(p_input[7758]), .B(p_input[17758]), .Z(o[7758]) );
  AND U2494 ( .A(p_input[7757]), .B(p_input[17757]), .Z(o[7757]) );
  AND U2495 ( .A(p_input[7756]), .B(p_input[17756]), .Z(o[7756]) );
  AND U2496 ( .A(p_input[7755]), .B(p_input[17755]), .Z(o[7755]) );
  AND U2497 ( .A(p_input[7754]), .B(p_input[17754]), .Z(o[7754]) );
  AND U2498 ( .A(p_input[7753]), .B(p_input[17753]), .Z(o[7753]) );
  AND U2499 ( .A(p_input[7752]), .B(p_input[17752]), .Z(o[7752]) );
  AND U2500 ( .A(p_input[7751]), .B(p_input[17751]), .Z(o[7751]) );
  AND U2501 ( .A(p_input[7750]), .B(p_input[17750]), .Z(o[7750]) );
  AND U2502 ( .A(p_input[774]), .B(p_input[10774]), .Z(o[774]) );
  AND U2503 ( .A(p_input[7749]), .B(p_input[17749]), .Z(o[7749]) );
  AND U2504 ( .A(p_input[7748]), .B(p_input[17748]), .Z(o[7748]) );
  AND U2505 ( .A(p_input[7747]), .B(p_input[17747]), .Z(o[7747]) );
  AND U2506 ( .A(p_input[7746]), .B(p_input[17746]), .Z(o[7746]) );
  AND U2507 ( .A(p_input[7745]), .B(p_input[17745]), .Z(o[7745]) );
  AND U2508 ( .A(p_input[7744]), .B(p_input[17744]), .Z(o[7744]) );
  AND U2509 ( .A(p_input[7743]), .B(p_input[17743]), .Z(o[7743]) );
  AND U2510 ( .A(p_input[7742]), .B(p_input[17742]), .Z(o[7742]) );
  AND U2511 ( .A(p_input[7741]), .B(p_input[17741]), .Z(o[7741]) );
  AND U2512 ( .A(p_input[7740]), .B(p_input[17740]), .Z(o[7740]) );
  AND U2513 ( .A(p_input[773]), .B(p_input[10773]), .Z(o[773]) );
  AND U2514 ( .A(p_input[7739]), .B(p_input[17739]), .Z(o[7739]) );
  AND U2515 ( .A(p_input[7738]), .B(p_input[17738]), .Z(o[7738]) );
  AND U2516 ( .A(p_input[7737]), .B(p_input[17737]), .Z(o[7737]) );
  AND U2517 ( .A(p_input[7736]), .B(p_input[17736]), .Z(o[7736]) );
  AND U2518 ( .A(p_input[7735]), .B(p_input[17735]), .Z(o[7735]) );
  AND U2519 ( .A(p_input[7734]), .B(p_input[17734]), .Z(o[7734]) );
  AND U2520 ( .A(p_input[7733]), .B(p_input[17733]), .Z(o[7733]) );
  AND U2521 ( .A(p_input[7732]), .B(p_input[17732]), .Z(o[7732]) );
  AND U2522 ( .A(p_input[7731]), .B(p_input[17731]), .Z(o[7731]) );
  AND U2523 ( .A(p_input[7730]), .B(p_input[17730]), .Z(o[7730]) );
  AND U2524 ( .A(p_input[772]), .B(p_input[10772]), .Z(o[772]) );
  AND U2525 ( .A(p_input[7729]), .B(p_input[17729]), .Z(o[7729]) );
  AND U2526 ( .A(p_input[7728]), .B(p_input[17728]), .Z(o[7728]) );
  AND U2527 ( .A(p_input[7727]), .B(p_input[17727]), .Z(o[7727]) );
  AND U2528 ( .A(p_input[7726]), .B(p_input[17726]), .Z(o[7726]) );
  AND U2529 ( .A(p_input[7725]), .B(p_input[17725]), .Z(o[7725]) );
  AND U2530 ( .A(p_input[7724]), .B(p_input[17724]), .Z(o[7724]) );
  AND U2531 ( .A(p_input[7723]), .B(p_input[17723]), .Z(o[7723]) );
  AND U2532 ( .A(p_input[7722]), .B(p_input[17722]), .Z(o[7722]) );
  AND U2533 ( .A(p_input[7721]), .B(p_input[17721]), .Z(o[7721]) );
  AND U2534 ( .A(p_input[7720]), .B(p_input[17720]), .Z(o[7720]) );
  AND U2535 ( .A(p_input[771]), .B(p_input[10771]), .Z(o[771]) );
  AND U2536 ( .A(p_input[7719]), .B(p_input[17719]), .Z(o[7719]) );
  AND U2537 ( .A(p_input[7718]), .B(p_input[17718]), .Z(o[7718]) );
  AND U2538 ( .A(p_input[7717]), .B(p_input[17717]), .Z(o[7717]) );
  AND U2539 ( .A(p_input[7716]), .B(p_input[17716]), .Z(o[7716]) );
  AND U2540 ( .A(p_input[7715]), .B(p_input[17715]), .Z(o[7715]) );
  AND U2541 ( .A(p_input[7714]), .B(p_input[17714]), .Z(o[7714]) );
  AND U2542 ( .A(p_input[7713]), .B(p_input[17713]), .Z(o[7713]) );
  AND U2543 ( .A(p_input[7712]), .B(p_input[17712]), .Z(o[7712]) );
  AND U2544 ( .A(p_input[7711]), .B(p_input[17711]), .Z(o[7711]) );
  AND U2545 ( .A(p_input[7710]), .B(p_input[17710]), .Z(o[7710]) );
  AND U2546 ( .A(p_input[770]), .B(p_input[10770]), .Z(o[770]) );
  AND U2547 ( .A(p_input[7709]), .B(p_input[17709]), .Z(o[7709]) );
  AND U2548 ( .A(p_input[7708]), .B(p_input[17708]), .Z(o[7708]) );
  AND U2549 ( .A(p_input[7707]), .B(p_input[17707]), .Z(o[7707]) );
  AND U2550 ( .A(p_input[7706]), .B(p_input[17706]), .Z(o[7706]) );
  AND U2551 ( .A(p_input[7705]), .B(p_input[17705]), .Z(o[7705]) );
  AND U2552 ( .A(p_input[7704]), .B(p_input[17704]), .Z(o[7704]) );
  AND U2553 ( .A(p_input[7703]), .B(p_input[17703]), .Z(o[7703]) );
  AND U2554 ( .A(p_input[7702]), .B(p_input[17702]), .Z(o[7702]) );
  AND U2555 ( .A(p_input[7701]), .B(p_input[17701]), .Z(o[7701]) );
  AND U2556 ( .A(p_input[7700]), .B(p_input[17700]), .Z(o[7700]) );
  AND U2557 ( .A(p_input[76]), .B(p_input[10076]), .Z(o[76]) );
  AND U2558 ( .A(p_input[769]), .B(p_input[10769]), .Z(o[769]) );
  AND U2559 ( .A(p_input[7699]), .B(p_input[17699]), .Z(o[7699]) );
  AND U2560 ( .A(p_input[7698]), .B(p_input[17698]), .Z(o[7698]) );
  AND U2561 ( .A(p_input[7697]), .B(p_input[17697]), .Z(o[7697]) );
  AND U2562 ( .A(p_input[7696]), .B(p_input[17696]), .Z(o[7696]) );
  AND U2563 ( .A(p_input[7695]), .B(p_input[17695]), .Z(o[7695]) );
  AND U2564 ( .A(p_input[7694]), .B(p_input[17694]), .Z(o[7694]) );
  AND U2565 ( .A(p_input[7693]), .B(p_input[17693]), .Z(o[7693]) );
  AND U2566 ( .A(p_input[7692]), .B(p_input[17692]), .Z(o[7692]) );
  AND U2567 ( .A(p_input[7691]), .B(p_input[17691]), .Z(o[7691]) );
  AND U2568 ( .A(p_input[7690]), .B(p_input[17690]), .Z(o[7690]) );
  AND U2569 ( .A(p_input[768]), .B(p_input[10768]), .Z(o[768]) );
  AND U2570 ( .A(p_input[7689]), .B(p_input[17689]), .Z(o[7689]) );
  AND U2571 ( .A(p_input[7688]), .B(p_input[17688]), .Z(o[7688]) );
  AND U2572 ( .A(p_input[7687]), .B(p_input[17687]), .Z(o[7687]) );
  AND U2573 ( .A(p_input[7686]), .B(p_input[17686]), .Z(o[7686]) );
  AND U2574 ( .A(p_input[7685]), .B(p_input[17685]), .Z(o[7685]) );
  AND U2575 ( .A(p_input[7684]), .B(p_input[17684]), .Z(o[7684]) );
  AND U2576 ( .A(p_input[7683]), .B(p_input[17683]), .Z(o[7683]) );
  AND U2577 ( .A(p_input[7682]), .B(p_input[17682]), .Z(o[7682]) );
  AND U2578 ( .A(p_input[7681]), .B(p_input[17681]), .Z(o[7681]) );
  AND U2579 ( .A(p_input[7680]), .B(p_input[17680]), .Z(o[7680]) );
  AND U2580 ( .A(p_input[767]), .B(p_input[10767]), .Z(o[767]) );
  AND U2581 ( .A(p_input[7679]), .B(p_input[17679]), .Z(o[7679]) );
  AND U2582 ( .A(p_input[7678]), .B(p_input[17678]), .Z(o[7678]) );
  AND U2583 ( .A(p_input[7677]), .B(p_input[17677]), .Z(o[7677]) );
  AND U2584 ( .A(p_input[7676]), .B(p_input[17676]), .Z(o[7676]) );
  AND U2585 ( .A(p_input[7675]), .B(p_input[17675]), .Z(o[7675]) );
  AND U2586 ( .A(p_input[7674]), .B(p_input[17674]), .Z(o[7674]) );
  AND U2587 ( .A(p_input[7673]), .B(p_input[17673]), .Z(o[7673]) );
  AND U2588 ( .A(p_input[7672]), .B(p_input[17672]), .Z(o[7672]) );
  AND U2589 ( .A(p_input[7671]), .B(p_input[17671]), .Z(o[7671]) );
  AND U2590 ( .A(p_input[7670]), .B(p_input[17670]), .Z(o[7670]) );
  AND U2591 ( .A(p_input[766]), .B(p_input[10766]), .Z(o[766]) );
  AND U2592 ( .A(p_input[7669]), .B(p_input[17669]), .Z(o[7669]) );
  AND U2593 ( .A(p_input[7668]), .B(p_input[17668]), .Z(o[7668]) );
  AND U2594 ( .A(p_input[7667]), .B(p_input[17667]), .Z(o[7667]) );
  AND U2595 ( .A(p_input[7666]), .B(p_input[17666]), .Z(o[7666]) );
  AND U2596 ( .A(p_input[7665]), .B(p_input[17665]), .Z(o[7665]) );
  AND U2597 ( .A(p_input[7664]), .B(p_input[17664]), .Z(o[7664]) );
  AND U2598 ( .A(p_input[7663]), .B(p_input[17663]), .Z(o[7663]) );
  AND U2599 ( .A(p_input[7662]), .B(p_input[17662]), .Z(o[7662]) );
  AND U2600 ( .A(p_input[7661]), .B(p_input[17661]), .Z(o[7661]) );
  AND U2601 ( .A(p_input[7660]), .B(p_input[17660]), .Z(o[7660]) );
  AND U2602 ( .A(p_input[765]), .B(p_input[10765]), .Z(o[765]) );
  AND U2603 ( .A(p_input[7659]), .B(p_input[17659]), .Z(o[7659]) );
  AND U2604 ( .A(p_input[7658]), .B(p_input[17658]), .Z(o[7658]) );
  AND U2605 ( .A(p_input[7657]), .B(p_input[17657]), .Z(o[7657]) );
  AND U2606 ( .A(p_input[7656]), .B(p_input[17656]), .Z(o[7656]) );
  AND U2607 ( .A(p_input[7655]), .B(p_input[17655]), .Z(o[7655]) );
  AND U2608 ( .A(p_input[7654]), .B(p_input[17654]), .Z(o[7654]) );
  AND U2609 ( .A(p_input[7653]), .B(p_input[17653]), .Z(o[7653]) );
  AND U2610 ( .A(p_input[7652]), .B(p_input[17652]), .Z(o[7652]) );
  AND U2611 ( .A(p_input[7651]), .B(p_input[17651]), .Z(o[7651]) );
  AND U2612 ( .A(p_input[7650]), .B(p_input[17650]), .Z(o[7650]) );
  AND U2613 ( .A(p_input[764]), .B(p_input[10764]), .Z(o[764]) );
  AND U2614 ( .A(p_input[7649]), .B(p_input[17649]), .Z(o[7649]) );
  AND U2615 ( .A(p_input[7648]), .B(p_input[17648]), .Z(o[7648]) );
  AND U2616 ( .A(p_input[7647]), .B(p_input[17647]), .Z(o[7647]) );
  AND U2617 ( .A(p_input[7646]), .B(p_input[17646]), .Z(o[7646]) );
  AND U2618 ( .A(p_input[7645]), .B(p_input[17645]), .Z(o[7645]) );
  AND U2619 ( .A(p_input[7644]), .B(p_input[17644]), .Z(o[7644]) );
  AND U2620 ( .A(p_input[7643]), .B(p_input[17643]), .Z(o[7643]) );
  AND U2621 ( .A(p_input[7642]), .B(p_input[17642]), .Z(o[7642]) );
  AND U2622 ( .A(p_input[7641]), .B(p_input[17641]), .Z(o[7641]) );
  AND U2623 ( .A(p_input[7640]), .B(p_input[17640]), .Z(o[7640]) );
  AND U2624 ( .A(p_input[763]), .B(p_input[10763]), .Z(o[763]) );
  AND U2625 ( .A(p_input[7639]), .B(p_input[17639]), .Z(o[7639]) );
  AND U2626 ( .A(p_input[7638]), .B(p_input[17638]), .Z(o[7638]) );
  AND U2627 ( .A(p_input[7637]), .B(p_input[17637]), .Z(o[7637]) );
  AND U2628 ( .A(p_input[7636]), .B(p_input[17636]), .Z(o[7636]) );
  AND U2629 ( .A(p_input[7635]), .B(p_input[17635]), .Z(o[7635]) );
  AND U2630 ( .A(p_input[7634]), .B(p_input[17634]), .Z(o[7634]) );
  AND U2631 ( .A(p_input[7633]), .B(p_input[17633]), .Z(o[7633]) );
  AND U2632 ( .A(p_input[7632]), .B(p_input[17632]), .Z(o[7632]) );
  AND U2633 ( .A(p_input[7631]), .B(p_input[17631]), .Z(o[7631]) );
  AND U2634 ( .A(p_input[7630]), .B(p_input[17630]), .Z(o[7630]) );
  AND U2635 ( .A(p_input[762]), .B(p_input[10762]), .Z(o[762]) );
  AND U2636 ( .A(p_input[7629]), .B(p_input[17629]), .Z(o[7629]) );
  AND U2637 ( .A(p_input[7628]), .B(p_input[17628]), .Z(o[7628]) );
  AND U2638 ( .A(p_input[7627]), .B(p_input[17627]), .Z(o[7627]) );
  AND U2639 ( .A(p_input[7626]), .B(p_input[17626]), .Z(o[7626]) );
  AND U2640 ( .A(p_input[7625]), .B(p_input[17625]), .Z(o[7625]) );
  AND U2641 ( .A(p_input[7624]), .B(p_input[17624]), .Z(o[7624]) );
  AND U2642 ( .A(p_input[7623]), .B(p_input[17623]), .Z(o[7623]) );
  AND U2643 ( .A(p_input[7622]), .B(p_input[17622]), .Z(o[7622]) );
  AND U2644 ( .A(p_input[7621]), .B(p_input[17621]), .Z(o[7621]) );
  AND U2645 ( .A(p_input[7620]), .B(p_input[17620]), .Z(o[7620]) );
  AND U2646 ( .A(p_input[761]), .B(p_input[10761]), .Z(o[761]) );
  AND U2647 ( .A(p_input[7619]), .B(p_input[17619]), .Z(o[7619]) );
  AND U2648 ( .A(p_input[7618]), .B(p_input[17618]), .Z(o[7618]) );
  AND U2649 ( .A(p_input[7617]), .B(p_input[17617]), .Z(o[7617]) );
  AND U2650 ( .A(p_input[7616]), .B(p_input[17616]), .Z(o[7616]) );
  AND U2651 ( .A(p_input[7615]), .B(p_input[17615]), .Z(o[7615]) );
  AND U2652 ( .A(p_input[7614]), .B(p_input[17614]), .Z(o[7614]) );
  AND U2653 ( .A(p_input[7613]), .B(p_input[17613]), .Z(o[7613]) );
  AND U2654 ( .A(p_input[7612]), .B(p_input[17612]), .Z(o[7612]) );
  AND U2655 ( .A(p_input[7611]), .B(p_input[17611]), .Z(o[7611]) );
  AND U2656 ( .A(p_input[7610]), .B(p_input[17610]), .Z(o[7610]) );
  AND U2657 ( .A(p_input[760]), .B(p_input[10760]), .Z(o[760]) );
  AND U2658 ( .A(p_input[7609]), .B(p_input[17609]), .Z(o[7609]) );
  AND U2659 ( .A(p_input[7608]), .B(p_input[17608]), .Z(o[7608]) );
  AND U2660 ( .A(p_input[7607]), .B(p_input[17607]), .Z(o[7607]) );
  AND U2661 ( .A(p_input[7606]), .B(p_input[17606]), .Z(o[7606]) );
  AND U2662 ( .A(p_input[7605]), .B(p_input[17605]), .Z(o[7605]) );
  AND U2663 ( .A(p_input[7604]), .B(p_input[17604]), .Z(o[7604]) );
  AND U2664 ( .A(p_input[7603]), .B(p_input[17603]), .Z(o[7603]) );
  AND U2665 ( .A(p_input[7602]), .B(p_input[17602]), .Z(o[7602]) );
  AND U2666 ( .A(p_input[7601]), .B(p_input[17601]), .Z(o[7601]) );
  AND U2667 ( .A(p_input[7600]), .B(p_input[17600]), .Z(o[7600]) );
  AND U2668 ( .A(p_input[75]), .B(p_input[10075]), .Z(o[75]) );
  AND U2669 ( .A(p_input[759]), .B(p_input[10759]), .Z(o[759]) );
  AND U2670 ( .A(p_input[7599]), .B(p_input[17599]), .Z(o[7599]) );
  AND U2671 ( .A(p_input[7598]), .B(p_input[17598]), .Z(o[7598]) );
  AND U2672 ( .A(p_input[7597]), .B(p_input[17597]), .Z(o[7597]) );
  AND U2673 ( .A(p_input[7596]), .B(p_input[17596]), .Z(o[7596]) );
  AND U2674 ( .A(p_input[7595]), .B(p_input[17595]), .Z(o[7595]) );
  AND U2675 ( .A(p_input[7594]), .B(p_input[17594]), .Z(o[7594]) );
  AND U2676 ( .A(p_input[7593]), .B(p_input[17593]), .Z(o[7593]) );
  AND U2677 ( .A(p_input[7592]), .B(p_input[17592]), .Z(o[7592]) );
  AND U2678 ( .A(p_input[7591]), .B(p_input[17591]), .Z(o[7591]) );
  AND U2679 ( .A(p_input[7590]), .B(p_input[17590]), .Z(o[7590]) );
  AND U2680 ( .A(p_input[758]), .B(p_input[10758]), .Z(o[758]) );
  AND U2681 ( .A(p_input[7589]), .B(p_input[17589]), .Z(o[7589]) );
  AND U2682 ( .A(p_input[7588]), .B(p_input[17588]), .Z(o[7588]) );
  AND U2683 ( .A(p_input[7587]), .B(p_input[17587]), .Z(o[7587]) );
  AND U2684 ( .A(p_input[7586]), .B(p_input[17586]), .Z(o[7586]) );
  AND U2685 ( .A(p_input[7585]), .B(p_input[17585]), .Z(o[7585]) );
  AND U2686 ( .A(p_input[7584]), .B(p_input[17584]), .Z(o[7584]) );
  AND U2687 ( .A(p_input[7583]), .B(p_input[17583]), .Z(o[7583]) );
  AND U2688 ( .A(p_input[7582]), .B(p_input[17582]), .Z(o[7582]) );
  AND U2689 ( .A(p_input[7581]), .B(p_input[17581]), .Z(o[7581]) );
  AND U2690 ( .A(p_input[7580]), .B(p_input[17580]), .Z(o[7580]) );
  AND U2691 ( .A(p_input[757]), .B(p_input[10757]), .Z(o[757]) );
  AND U2692 ( .A(p_input[7579]), .B(p_input[17579]), .Z(o[7579]) );
  AND U2693 ( .A(p_input[7578]), .B(p_input[17578]), .Z(o[7578]) );
  AND U2694 ( .A(p_input[7577]), .B(p_input[17577]), .Z(o[7577]) );
  AND U2695 ( .A(p_input[7576]), .B(p_input[17576]), .Z(o[7576]) );
  AND U2696 ( .A(p_input[7575]), .B(p_input[17575]), .Z(o[7575]) );
  AND U2697 ( .A(p_input[7574]), .B(p_input[17574]), .Z(o[7574]) );
  AND U2698 ( .A(p_input[7573]), .B(p_input[17573]), .Z(o[7573]) );
  AND U2699 ( .A(p_input[7572]), .B(p_input[17572]), .Z(o[7572]) );
  AND U2700 ( .A(p_input[7571]), .B(p_input[17571]), .Z(o[7571]) );
  AND U2701 ( .A(p_input[7570]), .B(p_input[17570]), .Z(o[7570]) );
  AND U2702 ( .A(p_input[756]), .B(p_input[10756]), .Z(o[756]) );
  AND U2703 ( .A(p_input[7569]), .B(p_input[17569]), .Z(o[7569]) );
  AND U2704 ( .A(p_input[7568]), .B(p_input[17568]), .Z(o[7568]) );
  AND U2705 ( .A(p_input[7567]), .B(p_input[17567]), .Z(o[7567]) );
  AND U2706 ( .A(p_input[7566]), .B(p_input[17566]), .Z(o[7566]) );
  AND U2707 ( .A(p_input[7565]), .B(p_input[17565]), .Z(o[7565]) );
  AND U2708 ( .A(p_input[7564]), .B(p_input[17564]), .Z(o[7564]) );
  AND U2709 ( .A(p_input[7563]), .B(p_input[17563]), .Z(o[7563]) );
  AND U2710 ( .A(p_input[7562]), .B(p_input[17562]), .Z(o[7562]) );
  AND U2711 ( .A(p_input[7561]), .B(p_input[17561]), .Z(o[7561]) );
  AND U2712 ( .A(p_input[7560]), .B(p_input[17560]), .Z(o[7560]) );
  AND U2713 ( .A(p_input[755]), .B(p_input[10755]), .Z(o[755]) );
  AND U2714 ( .A(p_input[7559]), .B(p_input[17559]), .Z(o[7559]) );
  AND U2715 ( .A(p_input[7558]), .B(p_input[17558]), .Z(o[7558]) );
  AND U2716 ( .A(p_input[7557]), .B(p_input[17557]), .Z(o[7557]) );
  AND U2717 ( .A(p_input[7556]), .B(p_input[17556]), .Z(o[7556]) );
  AND U2718 ( .A(p_input[7555]), .B(p_input[17555]), .Z(o[7555]) );
  AND U2719 ( .A(p_input[7554]), .B(p_input[17554]), .Z(o[7554]) );
  AND U2720 ( .A(p_input[7553]), .B(p_input[17553]), .Z(o[7553]) );
  AND U2721 ( .A(p_input[7552]), .B(p_input[17552]), .Z(o[7552]) );
  AND U2722 ( .A(p_input[7551]), .B(p_input[17551]), .Z(o[7551]) );
  AND U2723 ( .A(p_input[7550]), .B(p_input[17550]), .Z(o[7550]) );
  AND U2724 ( .A(p_input[754]), .B(p_input[10754]), .Z(o[754]) );
  AND U2725 ( .A(p_input[7549]), .B(p_input[17549]), .Z(o[7549]) );
  AND U2726 ( .A(p_input[7548]), .B(p_input[17548]), .Z(o[7548]) );
  AND U2727 ( .A(p_input[7547]), .B(p_input[17547]), .Z(o[7547]) );
  AND U2728 ( .A(p_input[7546]), .B(p_input[17546]), .Z(o[7546]) );
  AND U2729 ( .A(p_input[7545]), .B(p_input[17545]), .Z(o[7545]) );
  AND U2730 ( .A(p_input[7544]), .B(p_input[17544]), .Z(o[7544]) );
  AND U2731 ( .A(p_input[7543]), .B(p_input[17543]), .Z(o[7543]) );
  AND U2732 ( .A(p_input[7542]), .B(p_input[17542]), .Z(o[7542]) );
  AND U2733 ( .A(p_input[7541]), .B(p_input[17541]), .Z(o[7541]) );
  AND U2734 ( .A(p_input[7540]), .B(p_input[17540]), .Z(o[7540]) );
  AND U2735 ( .A(p_input[753]), .B(p_input[10753]), .Z(o[753]) );
  AND U2736 ( .A(p_input[7539]), .B(p_input[17539]), .Z(o[7539]) );
  AND U2737 ( .A(p_input[7538]), .B(p_input[17538]), .Z(o[7538]) );
  AND U2738 ( .A(p_input[7537]), .B(p_input[17537]), .Z(o[7537]) );
  AND U2739 ( .A(p_input[7536]), .B(p_input[17536]), .Z(o[7536]) );
  AND U2740 ( .A(p_input[7535]), .B(p_input[17535]), .Z(o[7535]) );
  AND U2741 ( .A(p_input[7534]), .B(p_input[17534]), .Z(o[7534]) );
  AND U2742 ( .A(p_input[7533]), .B(p_input[17533]), .Z(o[7533]) );
  AND U2743 ( .A(p_input[7532]), .B(p_input[17532]), .Z(o[7532]) );
  AND U2744 ( .A(p_input[7531]), .B(p_input[17531]), .Z(o[7531]) );
  AND U2745 ( .A(p_input[7530]), .B(p_input[17530]), .Z(o[7530]) );
  AND U2746 ( .A(p_input[752]), .B(p_input[10752]), .Z(o[752]) );
  AND U2747 ( .A(p_input[7529]), .B(p_input[17529]), .Z(o[7529]) );
  AND U2748 ( .A(p_input[7528]), .B(p_input[17528]), .Z(o[7528]) );
  AND U2749 ( .A(p_input[7527]), .B(p_input[17527]), .Z(o[7527]) );
  AND U2750 ( .A(p_input[7526]), .B(p_input[17526]), .Z(o[7526]) );
  AND U2751 ( .A(p_input[7525]), .B(p_input[17525]), .Z(o[7525]) );
  AND U2752 ( .A(p_input[7524]), .B(p_input[17524]), .Z(o[7524]) );
  AND U2753 ( .A(p_input[7523]), .B(p_input[17523]), .Z(o[7523]) );
  AND U2754 ( .A(p_input[7522]), .B(p_input[17522]), .Z(o[7522]) );
  AND U2755 ( .A(p_input[7521]), .B(p_input[17521]), .Z(o[7521]) );
  AND U2756 ( .A(p_input[7520]), .B(p_input[17520]), .Z(o[7520]) );
  AND U2757 ( .A(p_input[751]), .B(p_input[10751]), .Z(o[751]) );
  AND U2758 ( .A(p_input[7519]), .B(p_input[17519]), .Z(o[7519]) );
  AND U2759 ( .A(p_input[7518]), .B(p_input[17518]), .Z(o[7518]) );
  AND U2760 ( .A(p_input[7517]), .B(p_input[17517]), .Z(o[7517]) );
  AND U2761 ( .A(p_input[7516]), .B(p_input[17516]), .Z(o[7516]) );
  AND U2762 ( .A(p_input[7515]), .B(p_input[17515]), .Z(o[7515]) );
  AND U2763 ( .A(p_input[7514]), .B(p_input[17514]), .Z(o[7514]) );
  AND U2764 ( .A(p_input[7513]), .B(p_input[17513]), .Z(o[7513]) );
  AND U2765 ( .A(p_input[7512]), .B(p_input[17512]), .Z(o[7512]) );
  AND U2766 ( .A(p_input[7511]), .B(p_input[17511]), .Z(o[7511]) );
  AND U2767 ( .A(p_input[7510]), .B(p_input[17510]), .Z(o[7510]) );
  AND U2768 ( .A(p_input[750]), .B(p_input[10750]), .Z(o[750]) );
  AND U2769 ( .A(p_input[7509]), .B(p_input[17509]), .Z(o[7509]) );
  AND U2770 ( .A(p_input[7508]), .B(p_input[17508]), .Z(o[7508]) );
  AND U2771 ( .A(p_input[7507]), .B(p_input[17507]), .Z(o[7507]) );
  AND U2772 ( .A(p_input[7506]), .B(p_input[17506]), .Z(o[7506]) );
  AND U2773 ( .A(p_input[7505]), .B(p_input[17505]), .Z(o[7505]) );
  AND U2774 ( .A(p_input[7504]), .B(p_input[17504]), .Z(o[7504]) );
  AND U2775 ( .A(p_input[7503]), .B(p_input[17503]), .Z(o[7503]) );
  AND U2776 ( .A(p_input[7502]), .B(p_input[17502]), .Z(o[7502]) );
  AND U2777 ( .A(p_input[7501]), .B(p_input[17501]), .Z(o[7501]) );
  AND U2778 ( .A(p_input[7500]), .B(p_input[17500]), .Z(o[7500]) );
  AND U2779 ( .A(p_input[74]), .B(p_input[10074]), .Z(o[74]) );
  AND U2780 ( .A(p_input[749]), .B(p_input[10749]), .Z(o[749]) );
  AND U2781 ( .A(p_input[7499]), .B(p_input[17499]), .Z(o[7499]) );
  AND U2782 ( .A(p_input[7498]), .B(p_input[17498]), .Z(o[7498]) );
  AND U2783 ( .A(p_input[7497]), .B(p_input[17497]), .Z(o[7497]) );
  AND U2784 ( .A(p_input[7496]), .B(p_input[17496]), .Z(o[7496]) );
  AND U2785 ( .A(p_input[7495]), .B(p_input[17495]), .Z(o[7495]) );
  AND U2786 ( .A(p_input[7494]), .B(p_input[17494]), .Z(o[7494]) );
  AND U2787 ( .A(p_input[7493]), .B(p_input[17493]), .Z(o[7493]) );
  AND U2788 ( .A(p_input[7492]), .B(p_input[17492]), .Z(o[7492]) );
  AND U2789 ( .A(p_input[7491]), .B(p_input[17491]), .Z(o[7491]) );
  AND U2790 ( .A(p_input[7490]), .B(p_input[17490]), .Z(o[7490]) );
  AND U2791 ( .A(p_input[748]), .B(p_input[10748]), .Z(o[748]) );
  AND U2792 ( .A(p_input[7489]), .B(p_input[17489]), .Z(o[7489]) );
  AND U2793 ( .A(p_input[7488]), .B(p_input[17488]), .Z(o[7488]) );
  AND U2794 ( .A(p_input[7487]), .B(p_input[17487]), .Z(o[7487]) );
  AND U2795 ( .A(p_input[7486]), .B(p_input[17486]), .Z(o[7486]) );
  AND U2796 ( .A(p_input[7485]), .B(p_input[17485]), .Z(o[7485]) );
  AND U2797 ( .A(p_input[7484]), .B(p_input[17484]), .Z(o[7484]) );
  AND U2798 ( .A(p_input[7483]), .B(p_input[17483]), .Z(o[7483]) );
  AND U2799 ( .A(p_input[7482]), .B(p_input[17482]), .Z(o[7482]) );
  AND U2800 ( .A(p_input[7481]), .B(p_input[17481]), .Z(o[7481]) );
  AND U2801 ( .A(p_input[7480]), .B(p_input[17480]), .Z(o[7480]) );
  AND U2802 ( .A(p_input[747]), .B(p_input[10747]), .Z(o[747]) );
  AND U2803 ( .A(p_input[7479]), .B(p_input[17479]), .Z(o[7479]) );
  AND U2804 ( .A(p_input[7478]), .B(p_input[17478]), .Z(o[7478]) );
  AND U2805 ( .A(p_input[7477]), .B(p_input[17477]), .Z(o[7477]) );
  AND U2806 ( .A(p_input[7476]), .B(p_input[17476]), .Z(o[7476]) );
  AND U2807 ( .A(p_input[7475]), .B(p_input[17475]), .Z(o[7475]) );
  AND U2808 ( .A(p_input[7474]), .B(p_input[17474]), .Z(o[7474]) );
  AND U2809 ( .A(p_input[7473]), .B(p_input[17473]), .Z(o[7473]) );
  AND U2810 ( .A(p_input[7472]), .B(p_input[17472]), .Z(o[7472]) );
  AND U2811 ( .A(p_input[7471]), .B(p_input[17471]), .Z(o[7471]) );
  AND U2812 ( .A(p_input[7470]), .B(p_input[17470]), .Z(o[7470]) );
  AND U2813 ( .A(p_input[746]), .B(p_input[10746]), .Z(o[746]) );
  AND U2814 ( .A(p_input[7469]), .B(p_input[17469]), .Z(o[7469]) );
  AND U2815 ( .A(p_input[7468]), .B(p_input[17468]), .Z(o[7468]) );
  AND U2816 ( .A(p_input[7467]), .B(p_input[17467]), .Z(o[7467]) );
  AND U2817 ( .A(p_input[7466]), .B(p_input[17466]), .Z(o[7466]) );
  AND U2818 ( .A(p_input[7465]), .B(p_input[17465]), .Z(o[7465]) );
  AND U2819 ( .A(p_input[7464]), .B(p_input[17464]), .Z(o[7464]) );
  AND U2820 ( .A(p_input[7463]), .B(p_input[17463]), .Z(o[7463]) );
  AND U2821 ( .A(p_input[7462]), .B(p_input[17462]), .Z(o[7462]) );
  AND U2822 ( .A(p_input[7461]), .B(p_input[17461]), .Z(o[7461]) );
  AND U2823 ( .A(p_input[7460]), .B(p_input[17460]), .Z(o[7460]) );
  AND U2824 ( .A(p_input[745]), .B(p_input[10745]), .Z(o[745]) );
  AND U2825 ( .A(p_input[7459]), .B(p_input[17459]), .Z(o[7459]) );
  AND U2826 ( .A(p_input[7458]), .B(p_input[17458]), .Z(o[7458]) );
  AND U2827 ( .A(p_input[7457]), .B(p_input[17457]), .Z(o[7457]) );
  AND U2828 ( .A(p_input[7456]), .B(p_input[17456]), .Z(o[7456]) );
  AND U2829 ( .A(p_input[7455]), .B(p_input[17455]), .Z(o[7455]) );
  AND U2830 ( .A(p_input[7454]), .B(p_input[17454]), .Z(o[7454]) );
  AND U2831 ( .A(p_input[7453]), .B(p_input[17453]), .Z(o[7453]) );
  AND U2832 ( .A(p_input[7452]), .B(p_input[17452]), .Z(o[7452]) );
  AND U2833 ( .A(p_input[7451]), .B(p_input[17451]), .Z(o[7451]) );
  AND U2834 ( .A(p_input[7450]), .B(p_input[17450]), .Z(o[7450]) );
  AND U2835 ( .A(p_input[744]), .B(p_input[10744]), .Z(o[744]) );
  AND U2836 ( .A(p_input[7449]), .B(p_input[17449]), .Z(o[7449]) );
  AND U2837 ( .A(p_input[7448]), .B(p_input[17448]), .Z(o[7448]) );
  AND U2838 ( .A(p_input[7447]), .B(p_input[17447]), .Z(o[7447]) );
  AND U2839 ( .A(p_input[7446]), .B(p_input[17446]), .Z(o[7446]) );
  AND U2840 ( .A(p_input[7445]), .B(p_input[17445]), .Z(o[7445]) );
  AND U2841 ( .A(p_input[7444]), .B(p_input[17444]), .Z(o[7444]) );
  AND U2842 ( .A(p_input[7443]), .B(p_input[17443]), .Z(o[7443]) );
  AND U2843 ( .A(p_input[7442]), .B(p_input[17442]), .Z(o[7442]) );
  AND U2844 ( .A(p_input[7441]), .B(p_input[17441]), .Z(o[7441]) );
  AND U2845 ( .A(p_input[7440]), .B(p_input[17440]), .Z(o[7440]) );
  AND U2846 ( .A(p_input[743]), .B(p_input[10743]), .Z(o[743]) );
  AND U2847 ( .A(p_input[7439]), .B(p_input[17439]), .Z(o[7439]) );
  AND U2848 ( .A(p_input[7438]), .B(p_input[17438]), .Z(o[7438]) );
  AND U2849 ( .A(p_input[7437]), .B(p_input[17437]), .Z(o[7437]) );
  AND U2850 ( .A(p_input[7436]), .B(p_input[17436]), .Z(o[7436]) );
  AND U2851 ( .A(p_input[7435]), .B(p_input[17435]), .Z(o[7435]) );
  AND U2852 ( .A(p_input[7434]), .B(p_input[17434]), .Z(o[7434]) );
  AND U2853 ( .A(p_input[7433]), .B(p_input[17433]), .Z(o[7433]) );
  AND U2854 ( .A(p_input[7432]), .B(p_input[17432]), .Z(o[7432]) );
  AND U2855 ( .A(p_input[7431]), .B(p_input[17431]), .Z(o[7431]) );
  AND U2856 ( .A(p_input[7430]), .B(p_input[17430]), .Z(o[7430]) );
  AND U2857 ( .A(p_input[742]), .B(p_input[10742]), .Z(o[742]) );
  AND U2858 ( .A(p_input[7429]), .B(p_input[17429]), .Z(o[7429]) );
  AND U2859 ( .A(p_input[7428]), .B(p_input[17428]), .Z(o[7428]) );
  AND U2860 ( .A(p_input[7427]), .B(p_input[17427]), .Z(o[7427]) );
  AND U2861 ( .A(p_input[7426]), .B(p_input[17426]), .Z(o[7426]) );
  AND U2862 ( .A(p_input[7425]), .B(p_input[17425]), .Z(o[7425]) );
  AND U2863 ( .A(p_input[7424]), .B(p_input[17424]), .Z(o[7424]) );
  AND U2864 ( .A(p_input[7423]), .B(p_input[17423]), .Z(o[7423]) );
  AND U2865 ( .A(p_input[7422]), .B(p_input[17422]), .Z(o[7422]) );
  AND U2866 ( .A(p_input[7421]), .B(p_input[17421]), .Z(o[7421]) );
  AND U2867 ( .A(p_input[7420]), .B(p_input[17420]), .Z(o[7420]) );
  AND U2868 ( .A(p_input[741]), .B(p_input[10741]), .Z(o[741]) );
  AND U2869 ( .A(p_input[7419]), .B(p_input[17419]), .Z(o[7419]) );
  AND U2870 ( .A(p_input[7418]), .B(p_input[17418]), .Z(o[7418]) );
  AND U2871 ( .A(p_input[7417]), .B(p_input[17417]), .Z(o[7417]) );
  AND U2872 ( .A(p_input[7416]), .B(p_input[17416]), .Z(o[7416]) );
  AND U2873 ( .A(p_input[7415]), .B(p_input[17415]), .Z(o[7415]) );
  AND U2874 ( .A(p_input[7414]), .B(p_input[17414]), .Z(o[7414]) );
  AND U2875 ( .A(p_input[7413]), .B(p_input[17413]), .Z(o[7413]) );
  AND U2876 ( .A(p_input[7412]), .B(p_input[17412]), .Z(o[7412]) );
  AND U2877 ( .A(p_input[7411]), .B(p_input[17411]), .Z(o[7411]) );
  AND U2878 ( .A(p_input[7410]), .B(p_input[17410]), .Z(o[7410]) );
  AND U2879 ( .A(p_input[740]), .B(p_input[10740]), .Z(o[740]) );
  AND U2880 ( .A(p_input[7409]), .B(p_input[17409]), .Z(o[7409]) );
  AND U2881 ( .A(p_input[7408]), .B(p_input[17408]), .Z(o[7408]) );
  AND U2882 ( .A(p_input[7407]), .B(p_input[17407]), .Z(o[7407]) );
  AND U2883 ( .A(p_input[7406]), .B(p_input[17406]), .Z(o[7406]) );
  AND U2884 ( .A(p_input[7405]), .B(p_input[17405]), .Z(o[7405]) );
  AND U2885 ( .A(p_input[7404]), .B(p_input[17404]), .Z(o[7404]) );
  AND U2886 ( .A(p_input[7403]), .B(p_input[17403]), .Z(o[7403]) );
  AND U2887 ( .A(p_input[7402]), .B(p_input[17402]), .Z(o[7402]) );
  AND U2888 ( .A(p_input[7401]), .B(p_input[17401]), .Z(o[7401]) );
  AND U2889 ( .A(p_input[7400]), .B(p_input[17400]), .Z(o[7400]) );
  AND U2890 ( .A(p_input[73]), .B(p_input[10073]), .Z(o[73]) );
  AND U2891 ( .A(p_input[739]), .B(p_input[10739]), .Z(o[739]) );
  AND U2892 ( .A(p_input[7399]), .B(p_input[17399]), .Z(o[7399]) );
  AND U2893 ( .A(p_input[7398]), .B(p_input[17398]), .Z(o[7398]) );
  AND U2894 ( .A(p_input[7397]), .B(p_input[17397]), .Z(o[7397]) );
  AND U2895 ( .A(p_input[7396]), .B(p_input[17396]), .Z(o[7396]) );
  AND U2896 ( .A(p_input[7395]), .B(p_input[17395]), .Z(o[7395]) );
  AND U2897 ( .A(p_input[7394]), .B(p_input[17394]), .Z(o[7394]) );
  AND U2898 ( .A(p_input[7393]), .B(p_input[17393]), .Z(o[7393]) );
  AND U2899 ( .A(p_input[7392]), .B(p_input[17392]), .Z(o[7392]) );
  AND U2900 ( .A(p_input[7391]), .B(p_input[17391]), .Z(o[7391]) );
  AND U2901 ( .A(p_input[7390]), .B(p_input[17390]), .Z(o[7390]) );
  AND U2902 ( .A(p_input[738]), .B(p_input[10738]), .Z(o[738]) );
  AND U2903 ( .A(p_input[7389]), .B(p_input[17389]), .Z(o[7389]) );
  AND U2904 ( .A(p_input[7388]), .B(p_input[17388]), .Z(o[7388]) );
  AND U2905 ( .A(p_input[7387]), .B(p_input[17387]), .Z(o[7387]) );
  AND U2906 ( .A(p_input[7386]), .B(p_input[17386]), .Z(o[7386]) );
  AND U2907 ( .A(p_input[7385]), .B(p_input[17385]), .Z(o[7385]) );
  AND U2908 ( .A(p_input[7384]), .B(p_input[17384]), .Z(o[7384]) );
  AND U2909 ( .A(p_input[7383]), .B(p_input[17383]), .Z(o[7383]) );
  AND U2910 ( .A(p_input[7382]), .B(p_input[17382]), .Z(o[7382]) );
  AND U2911 ( .A(p_input[7381]), .B(p_input[17381]), .Z(o[7381]) );
  AND U2912 ( .A(p_input[7380]), .B(p_input[17380]), .Z(o[7380]) );
  AND U2913 ( .A(p_input[737]), .B(p_input[10737]), .Z(o[737]) );
  AND U2914 ( .A(p_input[7379]), .B(p_input[17379]), .Z(o[7379]) );
  AND U2915 ( .A(p_input[7378]), .B(p_input[17378]), .Z(o[7378]) );
  AND U2916 ( .A(p_input[7377]), .B(p_input[17377]), .Z(o[7377]) );
  AND U2917 ( .A(p_input[7376]), .B(p_input[17376]), .Z(o[7376]) );
  AND U2918 ( .A(p_input[7375]), .B(p_input[17375]), .Z(o[7375]) );
  AND U2919 ( .A(p_input[7374]), .B(p_input[17374]), .Z(o[7374]) );
  AND U2920 ( .A(p_input[7373]), .B(p_input[17373]), .Z(o[7373]) );
  AND U2921 ( .A(p_input[7372]), .B(p_input[17372]), .Z(o[7372]) );
  AND U2922 ( .A(p_input[7371]), .B(p_input[17371]), .Z(o[7371]) );
  AND U2923 ( .A(p_input[7370]), .B(p_input[17370]), .Z(o[7370]) );
  AND U2924 ( .A(p_input[736]), .B(p_input[10736]), .Z(o[736]) );
  AND U2925 ( .A(p_input[7369]), .B(p_input[17369]), .Z(o[7369]) );
  AND U2926 ( .A(p_input[7368]), .B(p_input[17368]), .Z(o[7368]) );
  AND U2927 ( .A(p_input[7367]), .B(p_input[17367]), .Z(o[7367]) );
  AND U2928 ( .A(p_input[7366]), .B(p_input[17366]), .Z(o[7366]) );
  AND U2929 ( .A(p_input[7365]), .B(p_input[17365]), .Z(o[7365]) );
  AND U2930 ( .A(p_input[7364]), .B(p_input[17364]), .Z(o[7364]) );
  AND U2931 ( .A(p_input[7363]), .B(p_input[17363]), .Z(o[7363]) );
  AND U2932 ( .A(p_input[7362]), .B(p_input[17362]), .Z(o[7362]) );
  AND U2933 ( .A(p_input[7361]), .B(p_input[17361]), .Z(o[7361]) );
  AND U2934 ( .A(p_input[7360]), .B(p_input[17360]), .Z(o[7360]) );
  AND U2935 ( .A(p_input[735]), .B(p_input[10735]), .Z(o[735]) );
  AND U2936 ( .A(p_input[7359]), .B(p_input[17359]), .Z(o[7359]) );
  AND U2937 ( .A(p_input[7358]), .B(p_input[17358]), .Z(o[7358]) );
  AND U2938 ( .A(p_input[7357]), .B(p_input[17357]), .Z(o[7357]) );
  AND U2939 ( .A(p_input[7356]), .B(p_input[17356]), .Z(o[7356]) );
  AND U2940 ( .A(p_input[7355]), .B(p_input[17355]), .Z(o[7355]) );
  AND U2941 ( .A(p_input[7354]), .B(p_input[17354]), .Z(o[7354]) );
  AND U2942 ( .A(p_input[7353]), .B(p_input[17353]), .Z(o[7353]) );
  AND U2943 ( .A(p_input[7352]), .B(p_input[17352]), .Z(o[7352]) );
  AND U2944 ( .A(p_input[7351]), .B(p_input[17351]), .Z(o[7351]) );
  AND U2945 ( .A(p_input[7350]), .B(p_input[17350]), .Z(o[7350]) );
  AND U2946 ( .A(p_input[734]), .B(p_input[10734]), .Z(o[734]) );
  AND U2947 ( .A(p_input[7349]), .B(p_input[17349]), .Z(o[7349]) );
  AND U2948 ( .A(p_input[7348]), .B(p_input[17348]), .Z(o[7348]) );
  AND U2949 ( .A(p_input[7347]), .B(p_input[17347]), .Z(o[7347]) );
  AND U2950 ( .A(p_input[7346]), .B(p_input[17346]), .Z(o[7346]) );
  AND U2951 ( .A(p_input[7345]), .B(p_input[17345]), .Z(o[7345]) );
  AND U2952 ( .A(p_input[7344]), .B(p_input[17344]), .Z(o[7344]) );
  AND U2953 ( .A(p_input[7343]), .B(p_input[17343]), .Z(o[7343]) );
  AND U2954 ( .A(p_input[7342]), .B(p_input[17342]), .Z(o[7342]) );
  AND U2955 ( .A(p_input[7341]), .B(p_input[17341]), .Z(o[7341]) );
  AND U2956 ( .A(p_input[7340]), .B(p_input[17340]), .Z(o[7340]) );
  AND U2957 ( .A(p_input[733]), .B(p_input[10733]), .Z(o[733]) );
  AND U2958 ( .A(p_input[7339]), .B(p_input[17339]), .Z(o[7339]) );
  AND U2959 ( .A(p_input[7338]), .B(p_input[17338]), .Z(o[7338]) );
  AND U2960 ( .A(p_input[7337]), .B(p_input[17337]), .Z(o[7337]) );
  AND U2961 ( .A(p_input[7336]), .B(p_input[17336]), .Z(o[7336]) );
  AND U2962 ( .A(p_input[7335]), .B(p_input[17335]), .Z(o[7335]) );
  AND U2963 ( .A(p_input[7334]), .B(p_input[17334]), .Z(o[7334]) );
  AND U2964 ( .A(p_input[7333]), .B(p_input[17333]), .Z(o[7333]) );
  AND U2965 ( .A(p_input[7332]), .B(p_input[17332]), .Z(o[7332]) );
  AND U2966 ( .A(p_input[7331]), .B(p_input[17331]), .Z(o[7331]) );
  AND U2967 ( .A(p_input[7330]), .B(p_input[17330]), .Z(o[7330]) );
  AND U2968 ( .A(p_input[732]), .B(p_input[10732]), .Z(o[732]) );
  AND U2969 ( .A(p_input[7329]), .B(p_input[17329]), .Z(o[7329]) );
  AND U2970 ( .A(p_input[7328]), .B(p_input[17328]), .Z(o[7328]) );
  AND U2971 ( .A(p_input[7327]), .B(p_input[17327]), .Z(o[7327]) );
  AND U2972 ( .A(p_input[7326]), .B(p_input[17326]), .Z(o[7326]) );
  AND U2973 ( .A(p_input[7325]), .B(p_input[17325]), .Z(o[7325]) );
  AND U2974 ( .A(p_input[7324]), .B(p_input[17324]), .Z(o[7324]) );
  AND U2975 ( .A(p_input[7323]), .B(p_input[17323]), .Z(o[7323]) );
  AND U2976 ( .A(p_input[7322]), .B(p_input[17322]), .Z(o[7322]) );
  AND U2977 ( .A(p_input[7321]), .B(p_input[17321]), .Z(o[7321]) );
  AND U2978 ( .A(p_input[7320]), .B(p_input[17320]), .Z(o[7320]) );
  AND U2979 ( .A(p_input[731]), .B(p_input[10731]), .Z(o[731]) );
  AND U2980 ( .A(p_input[7319]), .B(p_input[17319]), .Z(o[7319]) );
  AND U2981 ( .A(p_input[7318]), .B(p_input[17318]), .Z(o[7318]) );
  AND U2982 ( .A(p_input[7317]), .B(p_input[17317]), .Z(o[7317]) );
  AND U2983 ( .A(p_input[7316]), .B(p_input[17316]), .Z(o[7316]) );
  AND U2984 ( .A(p_input[7315]), .B(p_input[17315]), .Z(o[7315]) );
  AND U2985 ( .A(p_input[7314]), .B(p_input[17314]), .Z(o[7314]) );
  AND U2986 ( .A(p_input[7313]), .B(p_input[17313]), .Z(o[7313]) );
  AND U2987 ( .A(p_input[7312]), .B(p_input[17312]), .Z(o[7312]) );
  AND U2988 ( .A(p_input[7311]), .B(p_input[17311]), .Z(o[7311]) );
  AND U2989 ( .A(p_input[7310]), .B(p_input[17310]), .Z(o[7310]) );
  AND U2990 ( .A(p_input[730]), .B(p_input[10730]), .Z(o[730]) );
  AND U2991 ( .A(p_input[7309]), .B(p_input[17309]), .Z(o[7309]) );
  AND U2992 ( .A(p_input[7308]), .B(p_input[17308]), .Z(o[7308]) );
  AND U2993 ( .A(p_input[7307]), .B(p_input[17307]), .Z(o[7307]) );
  AND U2994 ( .A(p_input[7306]), .B(p_input[17306]), .Z(o[7306]) );
  AND U2995 ( .A(p_input[7305]), .B(p_input[17305]), .Z(o[7305]) );
  AND U2996 ( .A(p_input[7304]), .B(p_input[17304]), .Z(o[7304]) );
  AND U2997 ( .A(p_input[7303]), .B(p_input[17303]), .Z(o[7303]) );
  AND U2998 ( .A(p_input[7302]), .B(p_input[17302]), .Z(o[7302]) );
  AND U2999 ( .A(p_input[7301]), .B(p_input[17301]), .Z(o[7301]) );
  AND U3000 ( .A(p_input[7300]), .B(p_input[17300]), .Z(o[7300]) );
  AND U3001 ( .A(p_input[72]), .B(p_input[10072]), .Z(o[72]) );
  AND U3002 ( .A(p_input[729]), .B(p_input[10729]), .Z(o[729]) );
  AND U3003 ( .A(p_input[7299]), .B(p_input[17299]), .Z(o[7299]) );
  AND U3004 ( .A(p_input[7298]), .B(p_input[17298]), .Z(o[7298]) );
  AND U3005 ( .A(p_input[7297]), .B(p_input[17297]), .Z(o[7297]) );
  AND U3006 ( .A(p_input[7296]), .B(p_input[17296]), .Z(o[7296]) );
  AND U3007 ( .A(p_input[7295]), .B(p_input[17295]), .Z(o[7295]) );
  AND U3008 ( .A(p_input[7294]), .B(p_input[17294]), .Z(o[7294]) );
  AND U3009 ( .A(p_input[7293]), .B(p_input[17293]), .Z(o[7293]) );
  AND U3010 ( .A(p_input[7292]), .B(p_input[17292]), .Z(o[7292]) );
  AND U3011 ( .A(p_input[7291]), .B(p_input[17291]), .Z(o[7291]) );
  AND U3012 ( .A(p_input[7290]), .B(p_input[17290]), .Z(o[7290]) );
  AND U3013 ( .A(p_input[728]), .B(p_input[10728]), .Z(o[728]) );
  AND U3014 ( .A(p_input[7289]), .B(p_input[17289]), .Z(o[7289]) );
  AND U3015 ( .A(p_input[7288]), .B(p_input[17288]), .Z(o[7288]) );
  AND U3016 ( .A(p_input[7287]), .B(p_input[17287]), .Z(o[7287]) );
  AND U3017 ( .A(p_input[7286]), .B(p_input[17286]), .Z(o[7286]) );
  AND U3018 ( .A(p_input[7285]), .B(p_input[17285]), .Z(o[7285]) );
  AND U3019 ( .A(p_input[7284]), .B(p_input[17284]), .Z(o[7284]) );
  AND U3020 ( .A(p_input[7283]), .B(p_input[17283]), .Z(o[7283]) );
  AND U3021 ( .A(p_input[7282]), .B(p_input[17282]), .Z(o[7282]) );
  AND U3022 ( .A(p_input[7281]), .B(p_input[17281]), .Z(o[7281]) );
  AND U3023 ( .A(p_input[7280]), .B(p_input[17280]), .Z(o[7280]) );
  AND U3024 ( .A(p_input[727]), .B(p_input[10727]), .Z(o[727]) );
  AND U3025 ( .A(p_input[7279]), .B(p_input[17279]), .Z(o[7279]) );
  AND U3026 ( .A(p_input[7278]), .B(p_input[17278]), .Z(o[7278]) );
  AND U3027 ( .A(p_input[7277]), .B(p_input[17277]), .Z(o[7277]) );
  AND U3028 ( .A(p_input[7276]), .B(p_input[17276]), .Z(o[7276]) );
  AND U3029 ( .A(p_input[7275]), .B(p_input[17275]), .Z(o[7275]) );
  AND U3030 ( .A(p_input[7274]), .B(p_input[17274]), .Z(o[7274]) );
  AND U3031 ( .A(p_input[7273]), .B(p_input[17273]), .Z(o[7273]) );
  AND U3032 ( .A(p_input[7272]), .B(p_input[17272]), .Z(o[7272]) );
  AND U3033 ( .A(p_input[7271]), .B(p_input[17271]), .Z(o[7271]) );
  AND U3034 ( .A(p_input[7270]), .B(p_input[17270]), .Z(o[7270]) );
  AND U3035 ( .A(p_input[726]), .B(p_input[10726]), .Z(o[726]) );
  AND U3036 ( .A(p_input[7269]), .B(p_input[17269]), .Z(o[7269]) );
  AND U3037 ( .A(p_input[7268]), .B(p_input[17268]), .Z(o[7268]) );
  AND U3038 ( .A(p_input[7267]), .B(p_input[17267]), .Z(o[7267]) );
  AND U3039 ( .A(p_input[7266]), .B(p_input[17266]), .Z(o[7266]) );
  AND U3040 ( .A(p_input[7265]), .B(p_input[17265]), .Z(o[7265]) );
  AND U3041 ( .A(p_input[7264]), .B(p_input[17264]), .Z(o[7264]) );
  AND U3042 ( .A(p_input[7263]), .B(p_input[17263]), .Z(o[7263]) );
  AND U3043 ( .A(p_input[7262]), .B(p_input[17262]), .Z(o[7262]) );
  AND U3044 ( .A(p_input[7261]), .B(p_input[17261]), .Z(o[7261]) );
  AND U3045 ( .A(p_input[7260]), .B(p_input[17260]), .Z(o[7260]) );
  AND U3046 ( .A(p_input[725]), .B(p_input[10725]), .Z(o[725]) );
  AND U3047 ( .A(p_input[7259]), .B(p_input[17259]), .Z(o[7259]) );
  AND U3048 ( .A(p_input[7258]), .B(p_input[17258]), .Z(o[7258]) );
  AND U3049 ( .A(p_input[7257]), .B(p_input[17257]), .Z(o[7257]) );
  AND U3050 ( .A(p_input[7256]), .B(p_input[17256]), .Z(o[7256]) );
  AND U3051 ( .A(p_input[7255]), .B(p_input[17255]), .Z(o[7255]) );
  AND U3052 ( .A(p_input[7254]), .B(p_input[17254]), .Z(o[7254]) );
  AND U3053 ( .A(p_input[7253]), .B(p_input[17253]), .Z(o[7253]) );
  AND U3054 ( .A(p_input[7252]), .B(p_input[17252]), .Z(o[7252]) );
  AND U3055 ( .A(p_input[7251]), .B(p_input[17251]), .Z(o[7251]) );
  AND U3056 ( .A(p_input[7250]), .B(p_input[17250]), .Z(o[7250]) );
  AND U3057 ( .A(p_input[724]), .B(p_input[10724]), .Z(o[724]) );
  AND U3058 ( .A(p_input[7249]), .B(p_input[17249]), .Z(o[7249]) );
  AND U3059 ( .A(p_input[7248]), .B(p_input[17248]), .Z(o[7248]) );
  AND U3060 ( .A(p_input[7247]), .B(p_input[17247]), .Z(o[7247]) );
  AND U3061 ( .A(p_input[7246]), .B(p_input[17246]), .Z(o[7246]) );
  AND U3062 ( .A(p_input[7245]), .B(p_input[17245]), .Z(o[7245]) );
  AND U3063 ( .A(p_input[7244]), .B(p_input[17244]), .Z(o[7244]) );
  AND U3064 ( .A(p_input[7243]), .B(p_input[17243]), .Z(o[7243]) );
  AND U3065 ( .A(p_input[7242]), .B(p_input[17242]), .Z(o[7242]) );
  AND U3066 ( .A(p_input[7241]), .B(p_input[17241]), .Z(o[7241]) );
  AND U3067 ( .A(p_input[7240]), .B(p_input[17240]), .Z(o[7240]) );
  AND U3068 ( .A(p_input[723]), .B(p_input[10723]), .Z(o[723]) );
  AND U3069 ( .A(p_input[7239]), .B(p_input[17239]), .Z(o[7239]) );
  AND U3070 ( .A(p_input[7238]), .B(p_input[17238]), .Z(o[7238]) );
  AND U3071 ( .A(p_input[7237]), .B(p_input[17237]), .Z(o[7237]) );
  AND U3072 ( .A(p_input[7236]), .B(p_input[17236]), .Z(o[7236]) );
  AND U3073 ( .A(p_input[7235]), .B(p_input[17235]), .Z(o[7235]) );
  AND U3074 ( .A(p_input[7234]), .B(p_input[17234]), .Z(o[7234]) );
  AND U3075 ( .A(p_input[7233]), .B(p_input[17233]), .Z(o[7233]) );
  AND U3076 ( .A(p_input[7232]), .B(p_input[17232]), .Z(o[7232]) );
  AND U3077 ( .A(p_input[7231]), .B(p_input[17231]), .Z(o[7231]) );
  AND U3078 ( .A(p_input[7230]), .B(p_input[17230]), .Z(o[7230]) );
  AND U3079 ( .A(p_input[722]), .B(p_input[10722]), .Z(o[722]) );
  AND U3080 ( .A(p_input[7229]), .B(p_input[17229]), .Z(o[7229]) );
  AND U3081 ( .A(p_input[7228]), .B(p_input[17228]), .Z(o[7228]) );
  AND U3082 ( .A(p_input[7227]), .B(p_input[17227]), .Z(o[7227]) );
  AND U3083 ( .A(p_input[7226]), .B(p_input[17226]), .Z(o[7226]) );
  AND U3084 ( .A(p_input[7225]), .B(p_input[17225]), .Z(o[7225]) );
  AND U3085 ( .A(p_input[7224]), .B(p_input[17224]), .Z(o[7224]) );
  AND U3086 ( .A(p_input[7223]), .B(p_input[17223]), .Z(o[7223]) );
  AND U3087 ( .A(p_input[7222]), .B(p_input[17222]), .Z(o[7222]) );
  AND U3088 ( .A(p_input[7221]), .B(p_input[17221]), .Z(o[7221]) );
  AND U3089 ( .A(p_input[7220]), .B(p_input[17220]), .Z(o[7220]) );
  AND U3090 ( .A(p_input[721]), .B(p_input[10721]), .Z(o[721]) );
  AND U3091 ( .A(p_input[7219]), .B(p_input[17219]), .Z(o[7219]) );
  AND U3092 ( .A(p_input[7218]), .B(p_input[17218]), .Z(o[7218]) );
  AND U3093 ( .A(p_input[7217]), .B(p_input[17217]), .Z(o[7217]) );
  AND U3094 ( .A(p_input[7216]), .B(p_input[17216]), .Z(o[7216]) );
  AND U3095 ( .A(p_input[7215]), .B(p_input[17215]), .Z(o[7215]) );
  AND U3096 ( .A(p_input[7214]), .B(p_input[17214]), .Z(o[7214]) );
  AND U3097 ( .A(p_input[7213]), .B(p_input[17213]), .Z(o[7213]) );
  AND U3098 ( .A(p_input[7212]), .B(p_input[17212]), .Z(o[7212]) );
  AND U3099 ( .A(p_input[7211]), .B(p_input[17211]), .Z(o[7211]) );
  AND U3100 ( .A(p_input[7210]), .B(p_input[17210]), .Z(o[7210]) );
  AND U3101 ( .A(p_input[720]), .B(p_input[10720]), .Z(o[720]) );
  AND U3102 ( .A(p_input[7209]), .B(p_input[17209]), .Z(o[7209]) );
  AND U3103 ( .A(p_input[7208]), .B(p_input[17208]), .Z(o[7208]) );
  AND U3104 ( .A(p_input[7207]), .B(p_input[17207]), .Z(o[7207]) );
  AND U3105 ( .A(p_input[7206]), .B(p_input[17206]), .Z(o[7206]) );
  AND U3106 ( .A(p_input[7205]), .B(p_input[17205]), .Z(o[7205]) );
  AND U3107 ( .A(p_input[7204]), .B(p_input[17204]), .Z(o[7204]) );
  AND U3108 ( .A(p_input[7203]), .B(p_input[17203]), .Z(o[7203]) );
  AND U3109 ( .A(p_input[7202]), .B(p_input[17202]), .Z(o[7202]) );
  AND U3110 ( .A(p_input[7201]), .B(p_input[17201]), .Z(o[7201]) );
  AND U3111 ( .A(p_input[7200]), .B(p_input[17200]), .Z(o[7200]) );
  AND U3112 ( .A(p_input[71]), .B(p_input[10071]), .Z(o[71]) );
  AND U3113 ( .A(p_input[719]), .B(p_input[10719]), .Z(o[719]) );
  AND U3114 ( .A(p_input[7199]), .B(p_input[17199]), .Z(o[7199]) );
  AND U3115 ( .A(p_input[7198]), .B(p_input[17198]), .Z(o[7198]) );
  AND U3116 ( .A(p_input[7197]), .B(p_input[17197]), .Z(o[7197]) );
  AND U3117 ( .A(p_input[7196]), .B(p_input[17196]), .Z(o[7196]) );
  AND U3118 ( .A(p_input[7195]), .B(p_input[17195]), .Z(o[7195]) );
  AND U3119 ( .A(p_input[7194]), .B(p_input[17194]), .Z(o[7194]) );
  AND U3120 ( .A(p_input[7193]), .B(p_input[17193]), .Z(o[7193]) );
  AND U3121 ( .A(p_input[7192]), .B(p_input[17192]), .Z(o[7192]) );
  AND U3122 ( .A(p_input[7191]), .B(p_input[17191]), .Z(o[7191]) );
  AND U3123 ( .A(p_input[7190]), .B(p_input[17190]), .Z(o[7190]) );
  AND U3124 ( .A(p_input[718]), .B(p_input[10718]), .Z(o[718]) );
  AND U3125 ( .A(p_input[7189]), .B(p_input[17189]), .Z(o[7189]) );
  AND U3126 ( .A(p_input[7188]), .B(p_input[17188]), .Z(o[7188]) );
  AND U3127 ( .A(p_input[7187]), .B(p_input[17187]), .Z(o[7187]) );
  AND U3128 ( .A(p_input[7186]), .B(p_input[17186]), .Z(o[7186]) );
  AND U3129 ( .A(p_input[7185]), .B(p_input[17185]), .Z(o[7185]) );
  AND U3130 ( .A(p_input[7184]), .B(p_input[17184]), .Z(o[7184]) );
  AND U3131 ( .A(p_input[7183]), .B(p_input[17183]), .Z(o[7183]) );
  AND U3132 ( .A(p_input[7182]), .B(p_input[17182]), .Z(o[7182]) );
  AND U3133 ( .A(p_input[7181]), .B(p_input[17181]), .Z(o[7181]) );
  AND U3134 ( .A(p_input[7180]), .B(p_input[17180]), .Z(o[7180]) );
  AND U3135 ( .A(p_input[717]), .B(p_input[10717]), .Z(o[717]) );
  AND U3136 ( .A(p_input[7179]), .B(p_input[17179]), .Z(o[7179]) );
  AND U3137 ( .A(p_input[7178]), .B(p_input[17178]), .Z(o[7178]) );
  AND U3138 ( .A(p_input[7177]), .B(p_input[17177]), .Z(o[7177]) );
  AND U3139 ( .A(p_input[7176]), .B(p_input[17176]), .Z(o[7176]) );
  AND U3140 ( .A(p_input[7175]), .B(p_input[17175]), .Z(o[7175]) );
  AND U3141 ( .A(p_input[7174]), .B(p_input[17174]), .Z(o[7174]) );
  AND U3142 ( .A(p_input[7173]), .B(p_input[17173]), .Z(o[7173]) );
  AND U3143 ( .A(p_input[7172]), .B(p_input[17172]), .Z(o[7172]) );
  AND U3144 ( .A(p_input[7171]), .B(p_input[17171]), .Z(o[7171]) );
  AND U3145 ( .A(p_input[7170]), .B(p_input[17170]), .Z(o[7170]) );
  AND U3146 ( .A(p_input[716]), .B(p_input[10716]), .Z(o[716]) );
  AND U3147 ( .A(p_input[7169]), .B(p_input[17169]), .Z(o[7169]) );
  AND U3148 ( .A(p_input[7168]), .B(p_input[17168]), .Z(o[7168]) );
  AND U3149 ( .A(p_input[7167]), .B(p_input[17167]), .Z(o[7167]) );
  AND U3150 ( .A(p_input[7166]), .B(p_input[17166]), .Z(o[7166]) );
  AND U3151 ( .A(p_input[7165]), .B(p_input[17165]), .Z(o[7165]) );
  AND U3152 ( .A(p_input[7164]), .B(p_input[17164]), .Z(o[7164]) );
  AND U3153 ( .A(p_input[7163]), .B(p_input[17163]), .Z(o[7163]) );
  AND U3154 ( .A(p_input[7162]), .B(p_input[17162]), .Z(o[7162]) );
  AND U3155 ( .A(p_input[7161]), .B(p_input[17161]), .Z(o[7161]) );
  AND U3156 ( .A(p_input[7160]), .B(p_input[17160]), .Z(o[7160]) );
  AND U3157 ( .A(p_input[715]), .B(p_input[10715]), .Z(o[715]) );
  AND U3158 ( .A(p_input[7159]), .B(p_input[17159]), .Z(o[7159]) );
  AND U3159 ( .A(p_input[7158]), .B(p_input[17158]), .Z(o[7158]) );
  AND U3160 ( .A(p_input[7157]), .B(p_input[17157]), .Z(o[7157]) );
  AND U3161 ( .A(p_input[7156]), .B(p_input[17156]), .Z(o[7156]) );
  AND U3162 ( .A(p_input[7155]), .B(p_input[17155]), .Z(o[7155]) );
  AND U3163 ( .A(p_input[7154]), .B(p_input[17154]), .Z(o[7154]) );
  AND U3164 ( .A(p_input[7153]), .B(p_input[17153]), .Z(o[7153]) );
  AND U3165 ( .A(p_input[7152]), .B(p_input[17152]), .Z(o[7152]) );
  AND U3166 ( .A(p_input[7151]), .B(p_input[17151]), .Z(o[7151]) );
  AND U3167 ( .A(p_input[7150]), .B(p_input[17150]), .Z(o[7150]) );
  AND U3168 ( .A(p_input[714]), .B(p_input[10714]), .Z(o[714]) );
  AND U3169 ( .A(p_input[7149]), .B(p_input[17149]), .Z(o[7149]) );
  AND U3170 ( .A(p_input[7148]), .B(p_input[17148]), .Z(o[7148]) );
  AND U3171 ( .A(p_input[7147]), .B(p_input[17147]), .Z(o[7147]) );
  AND U3172 ( .A(p_input[7146]), .B(p_input[17146]), .Z(o[7146]) );
  AND U3173 ( .A(p_input[7145]), .B(p_input[17145]), .Z(o[7145]) );
  AND U3174 ( .A(p_input[7144]), .B(p_input[17144]), .Z(o[7144]) );
  AND U3175 ( .A(p_input[7143]), .B(p_input[17143]), .Z(o[7143]) );
  AND U3176 ( .A(p_input[7142]), .B(p_input[17142]), .Z(o[7142]) );
  AND U3177 ( .A(p_input[7141]), .B(p_input[17141]), .Z(o[7141]) );
  AND U3178 ( .A(p_input[7140]), .B(p_input[17140]), .Z(o[7140]) );
  AND U3179 ( .A(p_input[713]), .B(p_input[10713]), .Z(o[713]) );
  AND U3180 ( .A(p_input[7139]), .B(p_input[17139]), .Z(o[7139]) );
  AND U3181 ( .A(p_input[7138]), .B(p_input[17138]), .Z(o[7138]) );
  AND U3182 ( .A(p_input[7137]), .B(p_input[17137]), .Z(o[7137]) );
  AND U3183 ( .A(p_input[7136]), .B(p_input[17136]), .Z(o[7136]) );
  AND U3184 ( .A(p_input[7135]), .B(p_input[17135]), .Z(o[7135]) );
  AND U3185 ( .A(p_input[7134]), .B(p_input[17134]), .Z(o[7134]) );
  AND U3186 ( .A(p_input[7133]), .B(p_input[17133]), .Z(o[7133]) );
  AND U3187 ( .A(p_input[7132]), .B(p_input[17132]), .Z(o[7132]) );
  AND U3188 ( .A(p_input[7131]), .B(p_input[17131]), .Z(o[7131]) );
  AND U3189 ( .A(p_input[7130]), .B(p_input[17130]), .Z(o[7130]) );
  AND U3190 ( .A(p_input[712]), .B(p_input[10712]), .Z(o[712]) );
  AND U3191 ( .A(p_input[7129]), .B(p_input[17129]), .Z(o[7129]) );
  AND U3192 ( .A(p_input[7128]), .B(p_input[17128]), .Z(o[7128]) );
  AND U3193 ( .A(p_input[7127]), .B(p_input[17127]), .Z(o[7127]) );
  AND U3194 ( .A(p_input[7126]), .B(p_input[17126]), .Z(o[7126]) );
  AND U3195 ( .A(p_input[7125]), .B(p_input[17125]), .Z(o[7125]) );
  AND U3196 ( .A(p_input[7124]), .B(p_input[17124]), .Z(o[7124]) );
  AND U3197 ( .A(p_input[7123]), .B(p_input[17123]), .Z(o[7123]) );
  AND U3198 ( .A(p_input[7122]), .B(p_input[17122]), .Z(o[7122]) );
  AND U3199 ( .A(p_input[7121]), .B(p_input[17121]), .Z(o[7121]) );
  AND U3200 ( .A(p_input[7120]), .B(p_input[17120]), .Z(o[7120]) );
  AND U3201 ( .A(p_input[711]), .B(p_input[10711]), .Z(o[711]) );
  AND U3202 ( .A(p_input[7119]), .B(p_input[17119]), .Z(o[7119]) );
  AND U3203 ( .A(p_input[7118]), .B(p_input[17118]), .Z(o[7118]) );
  AND U3204 ( .A(p_input[7117]), .B(p_input[17117]), .Z(o[7117]) );
  AND U3205 ( .A(p_input[7116]), .B(p_input[17116]), .Z(o[7116]) );
  AND U3206 ( .A(p_input[7115]), .B(p_input[17115]), .Z(o[7115]) );
  AND U3207 ( .A(p_input[7114]), .B(p_input[17114]), .Z(o[7114]) );
  AND U3208 ( .A(p_input[7113]), .B(p_input[17113]), .Z(o[7113]) );
  AND U3209 ( .A(p_input[7112]), .B(p_input[17112]), .Z(o[7112]) );
  AND U3210 ( .A(p_input[7111]), .B(p_input[17111]), .Z(o[7111]) );
  AND U3211 ( .A(p_input[7110]), .B(p_input[17110]), .Z(o[7110]) );
  AND U3212 ( .A(p_input[710]), .B(p_input[10710]), .Z(o[710]) );
  AND U3213 ( .A(p_input[7109]), .B(p_input[17109]), .Z(o[7109]) );
  AND U3214 ( .A(p_input[7108]), .B(p_input[17108]), .Z(o[7108]) );
  AND U3215 ( .A(p_input[7107]), .B(p_input[17107]), .Z(o[7107]) );
  AND U3216 ( .A(p_input[7106]), .B(p_input[17106]), .Z(o[7106]) );
  AND U3217 ( .A(p_input[7105]), .B(p_input[17105]), .Z(o[7105]) );
  AND U3218 ( .A(p_input[7104]), .B(p_input[17104]), .Z(o[7104]) );
  AND U3219 ( .A(p_input[7103]), .B(p_input[17103]), .Z(o[7103]) );
  AND U3220 ( .A(p_input[7102]), .B(p_input[17102]), .Z(o[7102]) );
  AND U3221 ( .A(p_input[7101]), .B(p_input[17101]), .Z(o[7101]) );
  AND U3222 ( .A(p_input[7100]), .B(p_input[17100]), .Z(o[7100]) );
  AND U3223 ( .A(p_input[70]), .B(p_input[10070]), .Z(o[70]) );
  AND U3224 ( .A(p_input[709]), .B(p_input[10709]), .Z(o[709]) );
  AND U3225 ( .A(p_input[7099]), .B(p_input[17099]), .Z(o[7099]) );
  AND U3226 ( .A(p_input[7098]), .B(p_input[17098]), .Z(o[7098]) );
  AND U3227 ( .A(p_input[7097]), .B(p_input[17097]), .Z(o[7097]) );
  AND U3228 ( .A(p_input[7096]), .B(p_input[17096]), .Z(o[7096]) );
  AND U3229 ( .A(p_input[7095]), .B(p_input[17095]), .Z(o[7095]) );
  AND U3230 ( .A(p_input[7094]), .B(p_input[17094]), .Z(o[7094]) );
  AND U3231 ( .A(p_input[7093]), .B(p_input[17093]), .Z(o[7093]) );
  AND U3232 ( .A(p_input[7092]), .B(p_input[17092]), .Z(o[7092]) );
  AND U3233 ( .A(p_input[7091]), .B(p_input[17091]), .Z(o[7091]) );
  AND U3234 ( .A(p_input[7090]), .B(p_input[17090]), .Z(o[7090]) );
  AND U3235 ( .A(p_input[708]), .B(p_input[10708]), .Z(o[708]) );
  AND U3236 ( .A(p_input[7089]), .B(p_input[17089]), .Z(o[7089]) );
  AND U3237 ( .A(p_input[7088]), .B(p_input[17088]), .Z(o[7088]) );
  AND U3238 ( .A(p_input[7087]), .B(p_input[17087]), .Z(o[7087]) );
  AND U3239 ( .A(p_input[7086]), .B(p_input[17086]), .Z(o[7086]) );
  AND U3240 ( .A(p_input[7085]), .B(p_input[17085]), .Z(o[7085]) );
  AND U3241 ( .A(p_input[7084]), .B(p_input[17084]), .Z(o[7084]) );
  AND U3242 ( .A(p_input[7083]), .B(p_input[17083]), .Z(o[7083]) );
  AND U3243 ( .A(p_input[7082]), .B(p_input[17082]), .Z(o[7082]) );
  AND U3244 ( .A(p_input[7081]), .B(p_input[17081]), .Z(o[7081]) );
  AND U3245 ( .A(p_input[7080]), .B(p_input[17080]), .Z(o[7080]) );
  AND U3246 ( .A(p_input[707]), .B(p_input[10707]), .Z(o[707]) );
  AND U3247 ( .A(p_input[7079]), .B(p_input[17079]), .Z(o[7079]) );
  AND U3248 ( .A(p_input[7078]), .B(p_input[17078]), .Z(o[7078]) );
  AND U3249 ( .A(p_input[7077]), .B(p_input[17077]), .Z(o[7077]) );
  AND U3250 ( .A(p_input[7076]), .B(p_input[17076]), .Z(o[7076]) );
  AND U3251 ( .A(p_input[7075]), .B(p_input[17075]), .Z(o[7075]) );
  AND U3252 ( .A(p_input[7074]), .B(p_input[17074]), .Z(o[7074]) );
  AND U3253 ( .A(p_input[7073]), .B(p_input[17073]), .Z(o[7073]) );
  AND U3254 ( .A(p_input[7072]), .B(p_input[17072]), .Z(o[7072]) );
  AND U3255 ( .A(p_input[7071]), .B(p_input[17071]), .Z(o[7071]) );
  AND U3256 ( .A(p_input[7070]), .B(p_input[17070]), .Z(o[7070]) );
  AND U3257 ( .A(p_input[706]), .B(p_input[10706]), .Z(o[706]) );
  AND U3258 ( .A(p_input[7069]), .B(p_input[17069]), .Z(o[7069]) );
  AND U3259 ( .A(p_input[7068]), .B(p_input[17068]), .Z(o[7068]) );
  AND U3260 ( .A(p_input[7067]), .B(p_input[17067]), .Z(o[7067]) );
  AND U3261 ( .A(p_input[7066]), .B(p_input[17066]), .Z(o[7066]) );
  AND U3262 ( .A(p_input[7065]), .B(p_input[17065]), .Z(o[7065]) );
  AND U3263 ( .A(p_input[7064]), .B(p_input[17064]), .Z(o[7064]) );
  AND U3264 ( .A(p_input[7063]), .B(p_input[17063]), .Z(o[7063]) );
  AND U3265 ( .A(p_input[7062]), .B(p_input[17062]), .Z(o[7062]) );
  AND U3266 ( .A(p_input[7061]), .B(p_input[17061]), .Z(o[7061]) );
  AND U3267 ( .A(p_input[7060]), .B(p_input[17060]), .Z(o[7060]) );
  AND U3268 ( .A(p_input[705]), .B(p_input[10705]), .Z(o[705]) );
  AND U3269 ( .A(p_input[7059]), .B(p_input[17059]), .Z(o[7059]) );
  AND U3270 ( .A(p_input[7058]), .B(p_input[17058]), .Z(o[7058]) );
  AND U3271 ( .A(p_input[7057]), .B(p_input[17057]), .Z(o[7057]) );
  AND U3272 ( .A(p_input[7056]), .B(p_input[17056]), .Z(o[7056]) );
  AND U3273 ( .A(p_input[7055]), .B(p_input[17055]), .Z(o[7055]) );
  AND U3274 ( .A(p_input[7054]), .B(p_input[17054]), .Z(o[7054]) );
  AND U3275 ( .A(p_input[7053]), .B(p_input[17053]), .Z(o[7053]) );
  AND U3276 ( .A(p_input[7052]), .B(p_input[17052]), .Z(o[7052]) );
  AND U3277 ( .A(p_input[7051]), .B(p_input[17051]), .Z(o[7051]) );
  AND U3278 ( .A(p_input[7050]), .B(p_input[17050]), .Z(o[7050]) );
  AND U3279 ( .A(p_input[704]), .B(p_input[10704]), .Z(o[704]) );
  AND U3280 ( .A(p_input[7049]), .B(p_input[17049]), .Z(o[7049]) );
  AND U3281 ( .A(p_input[7048]), .B(p_input[17048]), .Z(o[7048]) );
  AND U3282 ( .A(p_input[7047]), .B(p_input[17047]), .Z(o[7047]) );
  AND U3283 ( .A(p_input[7046]), .B(p_input[17046]), .Z(o[7046]) );
  AND U3284 ( .A(p_input[7045]), .B(p_input[17045]), .Z(o[7045]) );
  AND U3285 ( .A(p_input[7044]), .B(p_input[17044]), .Z(o[7044]) );
  AND U3286 ( .A(p_input[7043]), .B(p_input[17043]), .Z(o[7043]) );
  AND U3287 ( .A(p_input[7042]), .B(p_input[17042]), .Z(o[7042]) );
  AND U3288 ( .A(p_input[7041]), .B(p_input[17041]), .Z(o[7041]) );
  AND U3289 ( .A(p_input[7040]), .B(p_input[17040]), .Z(o[7040]) );
  AND U3290 ( .A(p_input[703]), .B(p_input[10703]), .Z(o[703]) );
  AND U3291 ( .A(p_input[7039]), .B(p_input[17039]), .Z(o[7039]) );
  AND U3292 ( .A(p_input[7038]), .B(p_input[17038]), .Z(o[7038]) );
  AND U3293 ( .A(p_input[7037]), .B(p_input[17037]), .Z(o[7037]) );
  AND U3294 ( .A(p_input[7036]), .B(p_input[17036]), .Z(o[7036]) );
  AND U3295 ( .A(p_input[7035]), .B(p_input[17035]), .Z(o[7035]) );
  AND U3296 ( .A(p_input[7034]), .B(p_input[17034]), .Z(o[7034]) );
  AND U3297 ( .A(p_input[7033]), .B(p_input[17033]), .Z(o[7033]) );
  AND U3298 ( .A(p_input[7032]), .B(p_input[17032]), .Z(o[7032]) );
  AND U3299 ( .A(p_input[7031]), .B(p_input[17031]), .Z(o[7031]) );
  AND U3300 ( .A(p_input[7030]), .B(p_input[17030]), .Z(o[7030]) );
  AND U3301 ( .A(p_input[702]), .B(p_input[10702]), .Z(o[702]) );
  AND U3302 ( .A(p_input[7029]), .B(p_input[17029]), .Z(o[7029]) );
  AND U3303 ( .A(p_input[7028]), .B(p_input[17028]), .Z(o[7028]) );
  AND U3304 ( .A(p_input[7027]), .B(p_input[17027]), .Z(o[7027]) );
  AND U3305 ( .A(p_input[7026]), .B(p_input[17026]), .Z(o[7026]) );
  AND U3306 ( .A(p_input[7025]), .B(p_input[17025]), .Z(o[7025]) );
  AND U3307 ( .A(p_input[7024]), .B(p_input[17024]), .Z(o[7024]) );
  AND U3308 ( .A(p_input[7023]), .B(p_input[17023]), .Z(o[7023]) );
  AND U3309 ( .A(p_input[7022]), .B(p_input[17022]), .Z(o[7022]) );
  AND U3310 ( .A(p_input[7021]), .B(p_input[17021]), .Z(o[7021]) );
  AND U3311 ( .A(p_input[7020]), .B(p_input[17020]), .Z(o[7020]) );
  AND U3312 ( .A(p_input[701]), .B(p_input[10701]), .Z(o[701]) );
  AND U3313 ( .A(p_input[7019]), .B(p_input[17019]), .Z(o[7019]) );
  AND U3314 ( .A(p_input[7018]), .B(p_input[17018]), .Z(o[7018]) );
  AND U3315 ( .A(p_input[7017]), .B(p_input[17017]), .Z(o[7017]) );
  AND U3316 ( .A(p_input[7016]), .B(p_input[17016]), .Z(o[7016]) );
  AND U3317 ( .A(p_input[7015]), .B(p_input[17015]), .Z(o[7015]) );
  AND U3318 ( .A(p_input[7014]), .B(p_input[17014]), .Z(o[7014]) );
  AND U3319 ( .A(p_input[7013]), .B(p_input[17013]), .Z(o[7013]) );
  AND U3320 ( .A(p_input[7012]), .B(p_input[17012]), .Z(o[7012]) );
  AND U3321 ( .A(p_input[7011]), .B(p_input[17011]), .Z(o[7011]) );
  AND U3322 ( .A(p_input[7010]), .B(p_input[17010]), .Z(o[7010]) );
  AND U3323 ( .A(p_input[700]), .B(p_input[10700]), .Z(o[700]) );
  AND U3324 ( .A(p_input[7009]), .B(p_input[17009]), .Z(o[7009]) );
  AND U3325 ( .A(p_input[7008]), .B(p_input[17008]), .Z(o[7008]) );
  AND U3326 ( .A(p_input[7007]), .B(p_input[17007]), .Z(o[7007]) );
  AND U3327 ( .A(p_input[7006]), .B(p_input[17006]), .Z(o[7006]) );
  AND U3328 ( .A(p_input[7005]), .B(p_input[17005]), .Z(o[7005]) );
  AND U3329 ( .A(p_input[7004]), .B(p_input[17004]), .Z(o[7004]) );
  AND U3330 ( .A(p_input[7003]), .B(p_input[17003]), .Z(o[7003]) );
  AND U3331 ( .A(p_input[7002]), .B(p_input[17002]), .Z(o[7002]) );
  AND U3332 ( .A(p_input[7001]), .B(p_input[17001]), .Z(o[7001]) );
  AND U3333 ( .A(p_input[7000]), .B(p_input[17000]), .Z(o[7000]) );
  AND U3334 ( .A(p_input[6]), .B(p_input[10006]), .Z(o[6]) );
  AND U3335 ( .A(p_input[69]), .B(p_input[10069]), .Z(o[69]) );
  AND U3336 ( .A(p_input[699]), .B(p_input[10699]), .Z(o[699]) );
  AND U3337 ( .A(p_input[6999]), .B(p_input[16999]), .Z(o[6999]) );
  AND U3338 ( .A(p_input[6998]), .B(p_input[16998]), .Z(o[6998]) );
  AND U3339 ( .A(p_input[6997]), .B(p_input[16997]), .Z(o[6997]) );
  AND U3340 ( .A(p_input[6996]), .B(p_input[16996]), .Z(o[6996]) );
  AND U3341 ( .A(p_input[6995]), .B(p_input[16995]), .Z(o[6995]) );
  AND U3342 ( .A(p_input[6994]), .B(p_input[16994]), .Z(o[6994]) );
  AND U3343 ( .A(p_input[6993]), .B(p_input[16993]), .Z(o[6993]) );
  AND U3344 ( .A(p_input[6992]), .B(p_input[16992]), .Z(o[6992]) );
  AND U3345 ( .A(p_input[6991]), .B(p_input[16991]), .Z(o[6991]) );
  AND U3346 ( .A(p_input[6990]), .B(p_input[16990]), .Z(o[6990]) );
  AND U3347 ( .A(p_input[698]), .B(p_input[10698]), .Z(o[698]) );
  AND U3348 ( .A(p_input[6989]), .B(p_input[16989]), .Z(o[6989]) );
  AND U3349 ( .A(p_input[6988]), .B(p_input[16988]), .Z(o[6988]) );
  AND U3350 ( .A(p_input[6987]), .B(p_input[16987]), .Z(o[6987]) );
  AND U3351 ( .A(p_input[6986]), .B(p_input[16986]), .Z(o[6986]) );
  AND U3352 ( .A(p_input[6985]), .B(p_input[16985]), .Z(o[6985]) );
  AND U3353 ( .A(p_input[6984]), .B(p_input[16984]), .Z(o[6984]) );
  AND U3354 ( .A(p_input[6983]), .B(p_input[16983]), .Z(o[6983]) );
  AND U3355 ( .A(p_input[6982]), .B(p_input[16982]), .Z(o[6982]) );
  AND U3356 ( .A(p_input[6981]), .B(p_input[16981]), .Z(o[6981]) );
  AND U3357 ( .A(p_input[6980]), .B(p_input[16980]), .Z(o[6980]) );
  AND U3358 ( .A(p_input[697]), .B(p_input[10697]), .Z(o[697]) );
  AND U3359 ( .A(p_input[6979]), .B(p_input[16979]), .Z(o[6979]) );
  AND U3360 ( .A(p_input[6978]), .B(p_input[16978]), .Z(o[6978]) );
  AND U3361 ( .A(p_input[6977]), .B(p_input[16977]), .Z(o[6977]) );
  AND U3362 ( .A(p_input[6976]), .B(p_input[16976]), .Z(o[6976]) );
  AND U3363 ( .A(p_input[6975]), .B(p_input[16975]), .Z(o[6975]) );
  AND U3364 ( .A(p_input[6974]), .B(p_input[16974]), .Z(o[6974]) );
  AND U3365 ( .A(p_input[6973]), .B(p_input[16973]), .Z(o[6973]) );
  AND U3366 ( .A(p_input[6972]), .B(p_input[16972]), .Z(o[6972]) );
  AND U3367 ( .A(p_input[6971]), .B(p_input[16971]), .Z(o[6971]) );
  AND U3368 ( .A(p_input[6970]), .B(p_input[16970]), .Z(o[6970]) );
  AND U3369 ( .A(p_input[696]), .B(p_input[10696]), .Z(o[696]) );
  AND U3370 ( .A(p_input[6969]), .B(p_input[16969]), .Z(o[6969]) );
  AND U3371 ( .A(p_input[6968]), .B(p_input[16968]), .Z(o[6968]) );
  AND U3372 ( .A(p_input[6967]), .B(p_input[16967]), .Z(o[6967]) );
  AND U3373 ( .A(p_input[6966]), .B(p_input[16966]), .Z(o[6966]) );
  AND U3374 ( .A(p_input[6965]), .B(p_input[16965]), .Z(o[6965]) );
  AND U3375 ( .A(p_input[6964]), .B(p_input[16964]), .Z(o[6964]) );
  AND U3376 ( .A(p_input[6963]), .B(p_input[16963]), .Z(o[6963]) );
  AND U3377 ( .A(p_input[6962]), .B(p_input[16962]), .Z(o[6962]) );
  AND U3378 ( .A(p_input[6961]), .B(p_input[16961]), .Z(o[6961]) );
  AND U3379 ( .A(p_input[6960]), .B(p_input[16960]), .Z(o[6960]) );
  AND U3380 ( .A(p_input[695]), .B(p_input[10695]), .Z(o[695]) );
  AND U3381 ( .A(p_input[6959]), .B(p_input[16959]), .Z(o[6959]) );
  AND U3382 ( .A(p_input[6958]), .B(p_input[16958]), .Z(o[6958]) );
  AND U3383 ( .A(p_input[6957]), .B(p_input[16957]), .Z(o[6957]) );
  AND U3384 ( .A(p_input[6956]), .B(p_input[16956]), .Z(o[6956]) );
  AND U3385 ( .A(p_input[6955]), .B(p_input[16955]), .Z(o[6955]) );
  AND U3386 ( .A(p_input[6954]), .B(p_input[16954]), .Z(o[6954]) );
  AND U3387 ( .A(p_input[6953]), .B(p_input[16953]), .Z(o[6953]) );
  AND U3388 ( .A(p_input[6952]), .B(p_input[16952]), .Z(o[6952]) );
  AND U3389 ( .A(p_input[6951]), .B(p_input[16951]), .Z(o[6951]) );
  AND U3390 ( .A(p_input[6950]), .B(p_input[16950]), .Z(o[6950]) );
  AND U3391 ( .A(p_input[694]), .B(p_input[10694]), .Z(o[694]) );
  AND U3392 ( .A(p_input[6949]), .B(p_input[16949]), .Z(o[6949]) );
  AND U3393 ( .A(p_input[6948]), .B(p_input[16948]), .Z(o[6948]) );
  AND U3394 ( .A(p_input[6947]), .B(p_input[16947]), .Z(o[6947]) );
  AND U3395 ( .A(p_input[6946]), .B(p_input[16946]), .Z(o[6946]) );
  AND U3396 ( .A(p_input[6945]), .B(p_input[16945]), .Z(o[6945]) );
  AND U3397 ( .A(p_input[6944]), .B(p_input[16944]), .Z(o[6944]) );
  AND U3398 ( .A(p_input[6943]), .B(p_input[16943]), .Z(o[6943]) );
  AND U3399 ( .A(p_input[6942]), .B(p_input[16942]), .Z(o[6942]) );
  AND U3400 ( .A(p_input[6941]), .B(p_input[16941]), .Z(o[6941]) );
  AND U3401 ( .A(p_input[6940]), .B(p_input[16940]), .Z(o[6940]) );
  AND U3402 ( .A(p_input[693]), .B(p_input[10693]), .Z(o[693]) );
  AND U3403 ( .A(p_input[6939]), .B(p_input[16939]), .Z(o[6939]) );
  AND U3404 ( .A(p_input[6938]), .B(p_input[16938]), .Z(o[6938]) );
  AND U3405 ( .A(p_input[6937]), .B(p_input[16937]), .Z(o[6937]) );
  AND U3406 ( .A(p_input[6936]), .B(p_input[16936]), .Z(o[6936]) );
  AND U3407 ( .A(p_input[6935]), .B(p_input[16935]), .Z(o[6935]) );
  AND U3408 ( .A(p_input[6934]), .B(p_input[16934]), .Z(o[6934]) );
  AND U3409 ( .A(p_input[6933]), .B(p_input[16933]), .Z(o[6933]) );
  AND U3410 ( .A(p_input[6932]), .B(p_input[16932]), .Z(o[6932]) );
  AND U3411 ( .A(p_input[6931]), .B(p_input[16931]), .Z(o[6931]) );
  AND U3412 ( .A(p_input[6930]), .B(p_input[16930]), .Z(o[6930]) );
  AND U3413 ( .A(p_input[692]), .B(p_input[10692]), .Z(o[692]) );
  AND U3414 ( .A(p_input[6929]), .B(p_input[16929]), .Z(o[6929]) );
  AND U3415 ( .A(p_input[6928]), .B(p_input[16928]), .Z(o[6928]) );
  AND U3416 ( .A(p_input[6927]), .B(p_input[16927]), .Z(o[6927]) );
  AND U3417 ( .A(p_input[6926]), .B(p_input[16926]), .Z(o[6926]) );
  AND U3418 ( .A(p_input[6925]), .B(p_input[16925]), .Z(o[6925]) );
  AND U3419 ( .A(p_input[6924]), .B(p_input[16924]), .Z(o[6924]) );
  AND U3420 ( .A(p_input[6923]), .B(p_input[16923]), .Z(o[6923]) );
  AND U3421 ( .A(p_input[6922]), .B(p_input[16922]), .Z(o[6922]) );
  AND U3422 ( .A(p_input[6921]), .B(p_input[16921]), .Z(o[6921]) );
  AND U3423 ( .A(p_input[6920]), .B(p_input[16920]), .Z(o[6920]) );
  AND U3424 ( .A(p_input[691]), .B(p_input[10691]), .Z(o[691]) );
  AND U3425 ( .A(p_input[6919]), .B(p_input[16919]), .Z(o[6919]) );
  AND U3426 ( .A(p_input[6918]), .B(p_input[16918]), .Z(o[6918]) );
  AND U3427 ( .A(p_input[6917]), .B(p_input[16917]), .Z(o[6917]) );
  AND U3428 ( .A(p_input[6916]), .B(p_input[16916]), .Z(o[6916]) );
  AND U3429 ( .A(p_input[6915]), .B(p_input[16915]), .Z(o[6915]) );
  AND U3430 ( .A(p_input[6914]), .B(p_input[16914]), .Z(o[6914]) );
  AND U3431 ( .A(p_input[6913]), .B(p_input[16913]), .Z(o[6913]) );
  AND U3432 ( .A(p_input[6912]), .B(p_input[16912]), .Z(o[6912]) );
  AND U3433 ( .A(p_input[6911]), .B(p_input[16911]), .Z(o[6911]) );
  AND U3434 ( .A(p_input[6910]), .B(p_input[16910]), .Z(o[6910]) );
  AND U3435 ( .A(p_input[690]), .B(p_input[10690]), .Z(o[690]) );
  AND U3436 ( .A(p_input[6909]), .B(p_input[16909]), .Z(o[6909]) );
  AND U3437 ( .A(p_input[6908]), .B(p_input[16908]), .Z(o[6908]) );
  AND U3438 ( .A(p_input[6907]), .B(p_input[16907]), .Z(o[6907]) );
  AND U3439 ( .A(p_input[6906]), .B(p_input[16906]), .Z(o[6906]) );
  AND U3440 ( .A(p_input[6905]), .B(p_input[16905]), .Z(o[6905]) );
  AND U3441 ( .A(p_input[6904]), .B(p_input[16904]), .Z(o[6904]) );
  AND U3442 ( .A(p_input[6903]), .B(p_input[16903]), .Z(o[6903]) );
  AND U3443 ( .A(p_input[6902]), .B(p_input[16902]), .Z(o[6902]) );
  AND U3444 ( .A(p_input[6901]), .B(p_input[16901]), .Z(o[6901]) );
  AND U3445 ( .A(p_input[6900]), .B(p_input[16900]), .Z(o[6900]) );
  AND U3446 ( .A(p_input[68]), .B(p_input[10068]), .Z(o[68]) );
  AND U3447 ( .A(p_input[689]), .B(p_input[10689]), .Z(o[689]) );
  AND U3448 ( .A(p_input[6899]), .B(p_input[16899]), .Z(o[6899]) );
  AND U3449 ( .A(p_input[6898]), .B(p_input[16898]), .Z(o[6898]) );
  AND U3450 ( .A(p_input[6897]), .B(p_input[16897]), .Z(o[6897]) );
  AND U3451 ( .A(p_input[6896]), .B(p_input[16896]), .Z(o[6896]) );
  AND U3452 ( .A(p_input[6895]), .B(p_input[16895]), .Z(o[6895]) );
  AND U3453 ( .A(p_input[6894]), .B(p_input[16894]), .Z(o[6894]) );
  AND U3454 ( .A(p_input[6893]), .B(p_input[16893]), .Z(o[6893]) );
  AND U3455 ( .A(p_input[6892]), .B(p_input[16892]), .Z(o[6892]) );
  AND U3456 ( .A(p_input[6891]), .B(p_input[16891]), .Z(o[6891]) );
  AND U3457 ( .A(p_input[6890]), .B(p_input[16890]), .Z(o[6890]) );
  AND U3458 ( .A(p_input[688]), .B(p_input[10688]), .Z(o[688]) );
  AND U3459 ( .A(p_input[6889]), .B(p_input[16889]), .Z(o[6889]) );
  AND U3460 ( .A(p_input[6888]), .B(p_input[16888]), .Z(o[6888]) );
  AND U3461 ( .A(p_input[6887]), .B(p_input[16887]), .Z(o[6887]) );
  AND U3462 ( .A(p_input[6886]), .B(p_input[16886]), .Z(o[6886]) );
  AND U3463 ( .A(p_input[6885]), .B(p_input[16885]), .Z(o[6885]) );
  AND U3464 ( .A(p_input[6884]), .B(p_input[16884]), .Z(o[6884]) );
  AND U3465 ( .A(p_input[6883]), .B(p_input[16883]), .Z(o[6883]) );
  AND U3466 ( .A(p_input[6882]), .B(p_input[16882]), .Z(o[6882]) );
  AND U3467 ( .A(p_input[6881]), .B(p_input[16881]), .Z(o[6881]) );
  AND U3468 ( .A(p_input[6880]), .B(p_input[16880]), .Z(o[6880]) );
  AND U3469 ( .A(p_input[687]), .B(p_input[10687]), .Z(o[687]) );
  AND U3470 ( .A(p_input[6879]), .B(p_input[16879]), .Z(o[6879]) );
  AND U3471 ( .A(p_input[6878]), .B(p_input[16878]), .Z(o[6878]) );
  AND U3472 ( .A(p_input[6877]), .B(p_input[16877]), .Z(o[6877]) );
  AND U3473 ( .A(p_input[6876]), .B(p_input[16876]), .Z(o[6876]) );
  AND U3474 ( .A(p_input[6875]), .B(p_input[16875]), .Z(o[6875]) );
  AND U3475 ( .A(p_input[6874]), .B(p_input[16874]), .Z(o[6874]) );
  AND U3476 ( .A(p_input[6873]), .B(p_input[16873]), .Z(o[6873]) );
  AND U3477 ( .A(p_input[6872]), .B(p_input[16872]), .Z(o[6872]) );
  AND U3478 ( .A(p_input[6871]), .B(p_input[16871]), .Z(o[6871]) );
  AND U3479 ( .A(p_input[6870]), .B(p_input[16870]), .Z(o[6870]) );
  AND U3480 ( .A(p_input[686]), .B(p_input[10686]), .Z(o[686]) );
  AND U3481 ( .A(p_input[6869]), .B(p_input[16869]), .Z(o[6869]) );
  AND U3482 ( .A(p_input[6868]), .B(p_input[16868]), .Z(o[6868]) );
  AND U3483 ( .A(p_input[6867]), .B(p_input[16867]), .Z(o[6867]) );
  AND U3484 ( .A(p_input[6866]), .B(p_input[16866]), .Z(o[6866]) );
  AND U3485 ( .A(p_input[6865]), .B(p_input[16865]), .Z(o[6865]) );
  AND U3486 ( .A(p_input[6864]), .B(p_input[16864]), .Z(o[6864]) );
  AND U3487 ( .A(p_input[6863]), .B(p_input[16863]), .Z(o[6863]) );
  AND U3488 ( .A(p_input[6862]), .B(p_input[16862]), .Z(o[6862]) );
  AND U3489 ( .A(p_input[6861]), .B(p_input[16861]), .Z(o[6861]) );
  AND U3490 ( .A(p_input[6860]), .B(p_input[16860]), .Z(o[6860]) );
  AND U3491 ( .A(p_input[685]), .B(p_input[10685]), .Z(o[685]) );
  AND U3492 ( .A(p_input[6859]), .B(p_input[16859]), .Z(o[6859]) );
  AND U3493 ( .A(p_input[6858]), .B(p_input[16858]), .Z(o[6858]) );
  AND U3494 ( .A(p_input[6857]), .B(p_input[16857]), .Z(o[6857]) );
  AND U3495 ( .A(p_input[6856]), .B(p_input[16856]), .Z(o[6856]) );
  AND U3496 ( .A(p_input[6855]), .B(p_input[16855]), .Z(o[6855]) );
  AND U3497 ( .A(p_input[6854]), .B(p_input[16854]), .Z(o[6854]) );
  AND U3498 ( .A(p_input[6853]), .B(p_input[16853]), .Z(o[6853]) );
  AND U3499 ( .A(p_input[6852]), .B(p_input[16852]), .Z(o[6852]) );
  AND U3500 ( .A(p_input[6851]), .B(p_input[16851]), .Z(o[6851]) );
  AND U3501 ( .A(p_input[6850]), .B(p_input[16850]), .Z(o[6850]) );
  AND U3502 ( .A(p_input[684]), .B(p_input[10684]), .Z(o[684]) );
  AND U3503 ( .A(p_input[6849]), .B(p_input[16849]), .Z(o[6849]) );
  AND U3504 ( .A(p_input[6848]), .B(p_input[16848]), .Z(o[6848]) );
  AND U3505 ( .A(p_input[6847]), .B(p_input[16847]), .Z(o[6847]) );
  AND U3506 ( .A(p_input[6846]), .B(p_input[16846]), .Z(o[6846]) );
  AND U3507 ( .A(p_input[6845]), .B(p_input[16845]), .Z(o[6845]) );
  AND U3508 ( .A(p_input[6844]), .B(p_input[16844]), .Z(o[6844]) );
  AND U3509 ( .A(p_input[6843]), .B(p_input[16843]), .Z(o[6843]) );
  AND U3510 ( .A(p_input[6842]), .B(p_input[16842]), .Z(o[6842]) );
  AND U3511 ( .A(p_input[6841]), .B(p_input[16841]), .Z(o[6841]) );
  AND U3512 ( .A(p_input[6840]), .B(p_input[16840]), .Z(o[6840]) );
  AND U3513 ( .A(p_input[683]), .B(p_input[10683]), .Z(o[683]) );
  AND U3514 ( .A(p_input[6839]), .B(p_input[16839]), .Z(o[6839]) );
  AND U3515 ( .A(p_input[6838]), .B(p_input[16838]), .Z(o[6838]) );
  AND U3516 ( .A(p_input[6837]), .B(p_input[16837]), .Z(o[6837]) );
  AND U3517 ( .A(p_input[6836]), .B(p_input[16836]), .Z(o[6836]) );
  AND U3518 ( .A(p_input[6835]), .B(p_input[16835]), .Z(o[6835]) );
  AND U3519 ( .A(p_input[6834]), .B(p_input[16834]), .Z(o[6834]) );
  AND U3520 ( .A(p_input[6833]), .B(p_input[16833]), .Z(o[6833]) );
  AND U3521 ( .A(p_input[6832]), .B(p_input[16832]), .Z(o[6832]) );
  AND U3522 ( .A(p_input[6831]), .B(p_input[16831]), .Z(o[6831]) );
  AND U3523 ( .A(p_input[6830]), .B(p_input[16830]), .Z(o[6830]) );
  AND U3524 ( .A(p_input[682]), .B(p_input[10682]), .Z(o[682]) );
  AND U3525 ( .A(p_input[6829]), .B(p_input[16829]), .Z(o[6829]) );
  AND U3526 ( .A(p_input[6828]), .B(p_input[16828]), .Z(o[6828]) );
  AND U3527 ( .A(p_input[6827]), .B(p_input[16827]), .Z(o[6827]) );
  AND U3528 ( .A(p_input[6826]), .B(p_input[16826]), .Z(o[6826]) );
  AND U3529 ( .A(p_input[6825]), .B(p_input[16825]), .Z(o[6825]) );
  AND U3530 ( .A(p_input[6824]), .B(p_input[16824]), .Z(o[6824]) );
  AND U3531 ( .A(p_input[6823]), .B(p_input[16823]), .Z(o[6823]) );
  AND U3532 ( .A(p_input[6822]), .B(p_input[16822]), .Z(o[6822]) );
  AND U3533 ( .A(p_input[6821]), .B(p_input[16821]), .Z(o[6821]) );
  AND U3534 ( .A(p_input[6820]), .B(p_input[16820]), .Z(o[6820]) );
  AND U3535 ( .A(p_input[681]), .B(p_input[10681]), .Z(o[681]) );
  AND U3536 ( .A(p_input[6819]), .B(p_input[16819]), .Z(o[6819]) );
  AND U3537 ( .A(p_input[6818]), .B(p_input[16818]), .Z(o[6818]) );
  AND U3538 ( .A(p_input[6817]), .B(p_input[16817]), .Z(o[6817]) );
  AND U3539 ( .A(p_input[6816]), .B(p_input[16816]), .Z(o[6816]) );
  AND U3540 ( .A(p_input[6815]), .B(p_input[16815]), .Z(o[6815]) );
  AND U3541 ( .A(p_input[6814]), .B(p_input[16814]), .Z(o[6814]) );
  AND U3542 ( .A(p_input[6813]), .B(p_input[16813]), .Z(o[6813]) );
  AND U3543 ( .A(p_input[6812]), .B(p_input[16812]), .Z(o[6812]) );
  AND U3544 ( .A(p_input[6811]), .B(p_input[16811]), .Z(o[6811]) );
  AND U3545 ( .A(p_input[6810]), .B(p_input[16810]), .Z(o[6810]) );
  AND U3546 ( .A(p_input[680]), .B(p_input[10680]), .Z(o[680]) );
  AND U3547 ( .A(p_input[6809]), .B(p_input[16809]), .Z(o[6809]) );
  AND U3548 ( .A(p_input[6808]), .B(p_input[16808]), .Z(o[6808]) );
  AND U3549 ( .A(p_input[6807]), .B(p_input[16807]), .Z(o[6807]) );
  AND U3550 ( .A(p_input[6806]), .B(p_input[16806]), .Z(o[6806]) );
  AND U3551 ( .A(p_input[6805]), .B(p_input[16805]), .Z(o[6805]) );
  AND U3552 ( .A(p_input[6804]), .B(p_input[16804]), .Z(o[6804]) );
  AND U3553 ( .A(p_input[6803]), .B(p_input[16803]), .Z(o[6803]) );
  AND U3554 ( .A(p_input[6802]), .B(p_input[16802]), .Z(o[6802]) );
  AND U3555 ( .A(p_input[6801]), .B(p_input[16801]), .Z(o[6801]) );
  AND U3556 ( .A(p_input[6800]), .B(p_input[16800]), .Z(o[6800]) );
  AND U3557 ( .A(p_input[67]), .B(p_input[10067]), .Z(o[67]) );
  AND U3558 ( .A(p_input[679]), .B(p_input[10679]), .Z(o[679]) );
  AND U3559 ( .A(p_input[6799]), .B(p_input[16799]), .Z(o[6799]) );
  AND U3560 ( .A(p_input[6798]), .B(p_input[16798]), .Z(o[6798]) );
  AND U3561 ( .A(p_input[6797]), .B(p_input[16797]), .Z(o[6797]) );
  AND U3562 ( .A(p_input[6796]), .B(p_input[16796]), .Z(o[6796]) );
  AND U3563 ( .A(p_input[6795]), .B(p_input[16795]), .Z(o[6795]) );
  AND U3564 ( .A(p_input[6794]), .B(p_input[16794]), .Z(o[6794]) );
  AND U3565 ( .A(p_input[6793]), .B(p_input[16793]), .Z(o[6793]) );
  AND U3566 ( .A(p_input[6792]), .B(p_input[16792]), .Z(o[6792]) );
  AND U3567 ( .A(p_input[6791]), .B(p_input[16791]), .Z(o[6791]) );
  AND U3568 ( .A(p_input[6790]), .B(p_input[16790]), .Z(o[6790]) );
  AND U3569 ( .A(p_input[678]), .B(p_input[10678]), .Z(o[678]) );
  AND U3570 ( .A(p_input[6789]), .B(p_input[16789]), .Z(o[6789]) );
  AND U3571 ( .A(p_input[6788]), .B(p_input[16788]), .Z(o[6788]) );
  AND U3572 ( .A(p_input[6787]), .B(p_input[16787]), .Z(o[6787]) );
  AND U3573 ( .A(p_input[6786]), .B(p_input[16786]), .Z(o[6786]) );
  AND U3574 ( .A(p_input[6785]), .B(p_input[16785]), .Z(o[6785]) );
  AND U3575 ( .A(p_input[6784]), .B(p_input[16784]), .Z(o[6784]) );
  AND U3576 ( .A(p_input[6783]), .B(p_input[16783]), .Z(o[6783]) );
  AND U3577 ( .A(p_input[6782]), .B(p_input[16782]), .Z(o[6782]) );
  AND U3578 ( .A(p_input[6781]), .B(p_input[16781]), .Z(o[6781]) );
  AND U3579 ( .A(p_input[6780]), .B(p_input[16780]), .Z(o[6780]) );
  AND U3580 ( .A(p_input[677]), .B(p_input[10677]), .Z(o[677]) );
  AND U3581 ( .A(p_input[6779]), .B(p_input[16779]), .Z(o[6779]) );
  AND U3582 ( .A(p_input[6778]), .B(p_input[16778]), .Z(o[6778]) );
  AND U3583 ( .A(p_input[6777]), .B(p_input[16777]), .Z(o[6777]) );
  AND U3584 ( .A(p_input[6776]), .B(p_input[16776]), .Z(o[6776]) );
  AND U3585 ( .A(p_input[6775]), .B(p_input[16775]), .Z(o[6775]) );
  AND U3586 ( .A(p_input[6774]), .B(p_input[16774]), .Z(o[6774]) );
  AND U3587 ( .A(p_input[6773]), .B(p_input[16773]), .Z(o[6773]) );
  AND U3588 ( .A(p_input[6772]), .B(p_input[16772]), .Z(o[6772]) );
  AND U3589 ( .A(p_input[6771]), .B(p_input[16771]), .Z(o[6771]) );
  AND U3590 ( .A(p_input[6770]), .B(p_input[16770]), .Z(o[6770]) );
  AND U3591 ( .A(p_input[676]), .B(p_input[10676]), .Z(o[676]) );
  AND U3592 ( .A(p_input[6769]), .B(p_input[16769]), .Z(o[6769]) );
  AND U3593 ( .A(p_input[6768]), .B(p_input[16768]), .Z(o[6768]) );
  AND U3594 ( .A(p_input[6767]), .B(p_input[16767]), .Z(o[6767]) );
  AND U3595 ( .A(p_input[6766]), .B(p_input[16766]), .Z(o[6766]) );
  AND U3596 ( .A(p_input[6765]), .B(p_input[16765]), .Z(o[6765]) );
  AND U3597 ( .A(p_input[6764]), .B(p_input[16764]), .Z(o[6764]) );
  AND U3598 ( .A(p_input[6763]), .B(p_input[16763]), .Z(o[6763]) );
  AND U3599 ( .A(p_input[6762]), .B(p_input[16762]), .Z(o[6762]) );
  AND U3600 ( .A(p_input[6761]), .B(p_input[16761]), .Z(o[6761]) );
  AND U3601 ( .A(p_input[6760]), .B(p_input[16760]), .Z(o[6760]) );
  AND U3602 ( .A(p_input[675]), .B(p_input[10675]), .Z(o[675]) );
  AND U3603 ( .A(p_input[6759]), .B(p_input[16759]), .Z(o[6759]) );
  AND U3604 ( .A(p_input[6758]), .B(p_input[16758]), .Z(o[6758]) );
  AND U3605 ( .A(p_input[6757]), .B(p_input[16757]), .Z(o[6757]) );
  AND U3606 ( .A(p_input[6756]), .B(p_input[16756]), .Z(o[6756]) );
  AND U3607 ( .A(p_input[6755]), .B(p_input[16755]), .Z(o[6755]) );
  AND U3608 ( .A(p_input[6754]), .B(p_input[16754]), .Z(o[6754]) );
  AND U3609 ( .A(p_input[6753]), .B(p_input[16753]), .Z(o[6753]) );
  AND U3610 ( .A(p_input[6752]), .B(p_input[16752]), .Z(o[6752]) );
  AND U3611 ( .A(p_input[6751]), .B(p_input[16751]), .Z(o[6751]) );
  AND U3612 ( .A(p_input[6750]), .B(p_input[16750]), .Z(o[6750]) );
  AND U3613 ( .A(p_input[674]), .B(p_input[10674]), .Z(o[674]) );
  AND U3614 ( .A(p_input[6749]), .B(p_input[16749]), .Z(o[6749]) );
  AND U3615 ( .A(p_input[6748]), .B(p_input[16748]), .Z(o[6748]) );
  AND U3616 ( .A(p_input[6747]), .B(p_input[16747]), .Z(o[6747]) );
  AND U3617 ( .A(p_input[6746]), .B(p_input[16746]), .Z(o[6746]) );
  AND U3618 ( .A(p_input[6745]), .B(p_input[16745]), .Z(o[6745]) );
  AND U3619 ( .A(p_input[6744]), .B(p_input[16744]), .Z(o[6744]) );
  AND U3620 ( .A(p_input[6743]), .B(p_input[16743]), .Z(o[6743]) );
  AND U3621 ( .A(p_input[6742]), .B(p_input[16742]), .Z(o[6742]) );
  AND U3622 ( .A(p_input[6741]), .B(p_input[16741]), .Z(o[6741]) );
  AND U3623 ( .A(p_input[6740]), .B(p_input[16740]), .Z(o[6740]) );
  AND U3624 ( .A(p_input[673]), .B(p_input[10673]), .Z(o[673]) );
  AND U3625 ( .A(p_input[6739]), .B(p_input[16739]), .Z(o[6739]) );
  AND U3626 ( .A(p_input[6738]), .B(p_input[16738]), .Z(o[6738]) );
  AND U3627 ( .A(p_input[6737]), .B(p_input[16737]), .Z(o[6737]) );
  AND U3628 ( .A(p_input[6736]), .B(p_input[16736]), .Z(o[6736]) );
  AND U3629 ( .A(p_input[6735]), .B(p_input[16735]), .Z(o[6735]) );
  AND U3630 ( .A(p_input[6734]), .B(p_input[16734]), .Z(o[6734]) );
  AND U3631 ( .A(p_input[6733]), .B(p_input[16733]), .Z(o[6733]) );
  AND U3632 ( .A(p_input[6732]), .B(p_input[16732]), .Z(o[6732]) );
  AND U3633 ( .A(p_input[6731]), .B(p_input[16731]), .Z(o[6731]) );
  AND U3634 ( .A(p_input[6730]), .B(p_input[16730]), .Z(o[6730]) );
  AND U3635 ( .A(p_input[672]), .B(p_input[10672]), .Z(o[672]) );
  AND U3636 ( .A(p_input[6729]), .B(p_input[16729]), .Z(o[6729]) );
  AND U3637 ( .A(p_input[6728]), .B(p_input[16728]), .Z(o[6728]) );
  AND U3638 ( .A(p_input[6727]), .B(p_input[16727]), .Z(o[6727]) );
  AND U3639 ( .A(p_input[6726]), .B(p_input[16726]), .Z(o[6726]) );
  AND U3640 ( .A(p_input[6725]), .B(p_input[16725]), .Z(o[6725]) );
  AND U3641 ( .A(p_input[6724]), .B(p_input[16724]), .Z(o[6724]) );
  AND U3642 ( .A(p_input[6723]), .B(p_input[16723]), .Z(o[6723]) );
  AND U3643 ( .A(p_input[6722]), .B(p_input[16722]), .Z(o[6722]) );
  AND U3644 ( .A(p_input[6721]), .B(p_input[16721]), .Z(o[6721]) );
  AND U3645 ( .A(p_input[6720]), .B(p_input[16720]), .Z(o[6720]) );
  AND U3646 ( .A(p_input[671]), .B(p_input[10671]), .Z(o[671]) );
  AND U3647 ( .A(p_input[6719]), .B(p_input[16719]), .Z(o[6719]) );
  AND U3648 ( .A(p_input[6718]), .B(p_input[16718]), .Z(o[6718]) );
  AND U3649 ( .A(p_input[6717]), .B(p_input[16717]), .Z(o[6717]) );
  AND U3650 ( .A(p_input[6716]), .B(p_input[16716]), .Z(o[6716]) );
  AND U3651 ( .A(p_input[6715]), .B(p_input[16715]), .Z(o[6715]) );
  AND U3652 ( .A(p_input[6714]), .B(p_input[16714]), .Z(o[6714]) );
  AND U3653 ( .A(p_input[6713]), .B(p_input[16713]), .Z(o[6713]) );
  AND U3654 ( .A(p_input[6712]), .B(p_input[16712]), .Z(o[6712]) );
  AND U3655 ( .A(p_input[6711]), .B(p_input[16711]), .Z(o[6711]) );
  AND U3656 ( .A(p_input[6710]), .B(p_input[16710]), .Z(o[6710]) );
  AND U3657 ( .A(p_input[670]), .B(p_input[10670]), .Z(o[670]) );
  AND U3658 ( .A(p_input[6709]), .B(p_input[16709]), .Z(o[6709]) );
  AND U3659 ( .A(p_input[6708]), .B(p_input[16708]), .Z(o[6708]) );
  AND U3660 ( .A(p_input[6707]), .B(p_input[16707]), .Z(o[6707]) );
  AND U3661 ( .A(p_input[6706]), .B(p_input[16706]), .Z(o[6706]) );
  AND U3662 ( .A(p_input[6705]), .B(p_input[16705]), .Z(o[6705]) );
  AND U3663 ( .A(p_input[6704]), .B(p_input[16704]), .Z(o[6704]) );
  AND U3664 ( .A(p_input[6703]), .B(p_input[16703]), .Z(o[6703]) );
  AND U3665 ( .A(p_input[6702]), .B(p_input[16702]), .Z(o[6702]) );
  AND U3666 ( .A(p_input[6701]), .B(p_input[16701]), .Z(o[6701]) );
  AND U3667 ( .A(p_input[6700]), .B(p_input[16700]), .Z(o[6700]) );
  AND U3668 ( .A(p_input[66]), .B(p_input[10066]), .Z(o[66]) );
  AND U3669 ( .A(p_input[669]), .B(p_input[10669]), .Z(o[669]) );
  AND U3670 ( .A(p_input[6699]), .B(p_input[16699]), .Z(o[6699]) );
  AND U3671 ( .A(p_input[6698]), .B(p_input[16698]), .Z(o[6698]) );
  AND U3672 ( .A(p_input[6697]), .B(p_input[16697]), .Z(o[6697]) );
  AND U3673 ( .A(p_input[6696]), .B(p_input[16696]), .Z(o[6696]) );
  AND U3674 ( .A(p_input[6695]), .B(p_input[16695]), .Z(o[6695]) );
  AND U3675 ( .A(p_input[6694]), .B(p_input[16694]), .Z(o[6694]) );
  AND U3676 ( .A(p_input[6693]), .B(p_input[16693]), .Z(o[6693]) );
  AND U3677 ( .A(p_input[6692]), .B(p_input[16692]), .Z(o[6692]) );
  AND U3678 ( .A(p_input[6691]), .B(p_input[16691]), .Z(o[6691]) );
  AND U3679 ( .A(p_input[6690]), .B(p_input[16690]), .Z(o[6690]) );
  AND U3680 ( .A(p_input[668]), .B(p_input[10668]), .Z(o[668]) );
  AND U3681 ( .A(p_input[6689]), .B(p_input[16689]), .Z(o[6689]) );
  AND U3682 ( .A(p_input[6688]), .B(p_input[16688]), .Z(o[6688]) );
  AND U3683 ( .A(p_input[6687]), .B(p_input[16687]), .Z(o[6687]) );
  AND U3684 ( .A(p_input[6686]), .B(p_input[16686]), .Z(o[6686]) );
  AND U3685 ( .A(p_input[6685]), .B(p_input[16685]), .Z(o[6685]) );
  AND U3686 ( .A(p_input[6684]), .B(p_input[16684]), .Z(o[6684]) );
  AND U3687 ( .A(p_input[6683]), .B(p_input[16683]), .Z(o[6683]) );
  AND U3688 ( .A(p_input[6682]), .B(p_input[16682]), .Z(o[6682]) );
  AND U3689 ( .A(p_input[6681]), .B(p_input[16681]), .Z(o[6681]) );
  AND U3690 ( .A(p_input[6680]), .B(p_input[16680]), .Z(o[6680]) );
  AND U3691 ( .A(p_input[667]), .B(p_input[10667]), .Z(o[667]) );
  AND U3692 ( .A(p_input[6679]), .B(p_input[16679]), .Z(o[6679]) );
  AND U3693 ( .A(p_input[6678]), .B(p_input[16678]), .Z(o[6678]) );
  AND U3694 ( .A(p_input[6677]), .B(p_input[16677]), .Z(o[6677]) );
  AND U3695 ( .A(p_input[6676]), .B(p_input[16676]), .Z(o[6676]) );
  AND U3696 ( .A(p_input[6675]), .B(p_input[16675]), .Z(o[6675]) );
  AND U3697 ( .A(p_input[6674]), .B(p_input[16674]), .Z(o[6674]) );
  AND U3698 ( .A(p_input[6673]), .B(p_input[16673]), .Z(o[6673]) );
  AND U3699 ( .A(p_input[6672]), .B(p_input[16672]), .Z(o[6672]) );
  AND U3700 ( .A(p_input[6671]), .B(p_input[16671]), .Z(o[6671]) );
  AND U3701 ( .A(p_input[6670]), .B(p_input[16670]), .Z(o[6670]) );
  AND U3702 ( .A(p_input[666]), .B(p_input[10666]), .Z(o[666]) );
  AND U3703 ( .A(p_input[6669]), .B(p_input[16669]), .Z(o[6669]) );
  AND U3704 ( .A(p_input[6668]), .B(p_input[16668]), .Z(o[6668]) );
  AND U3705 ( .A(p_input[6667]), .B(p_input[16667]), .Z(o[6667]) );
  AND U3706 ( .A(p_input[6666]), .B(p_input[16666]), .Z(o[6666]) );
  AND U3707 ( .A(p_input[6665]), .B(p_input[16665]), .Z(o[6665]) );
  AND U3708 ( .A(p_input[6664]), .B(p_input[16664]), .Z(o[6664]) );
  AND U3709 ( .A(p_input[6663]), .B(p_input[16663]), .Z(o[6663]) );
  AND U3710 ( .A(p_input[6662]), .B(p_input[16662]), .Z(o[6662]) );
  AND U3711 ( .A(p_input[6661]), .B(p_input[16661]), .Z(o[6661]) );
  AND U3712 ( .A(p_input[6660]), .B(p_input[16660]), .Z(o[6660]) );
  AND U3713 ( .A(p_input[665]), .B(p_input[10665]), .Z(o[665]) );
  AND U3714 ( .A(p_input[6659]), .B(p_input[16659]), .Z(o[6659]) );
  AND U3715 ( .A(p_input[6658]), .B(p_input[16658]), .Z(o[6658]) );
  AND U3716 ( .A(p_input[6657]), .B(p_input[16657]), .Z(o[6657]) );
  AND U3717 ( .A(p_input[6656]), .B(p_input[16656]), .Z(o[6656]) );
  AND U3718 ( .A(p_input[6655]), .B(p_input[16655]), .Z(o[6655]) );
  AND U3719 ( .A(p_input[6654]), .B(p_input[16654]), .Z(o[6654]) );
  AND U3720 ( .A(p_input[6653]), .B(p_input[16653]), .Z(o[6653]) );
  AND U3721 ( .A(p_input[6652]), .B(p_input[16652]), .Z(o[6652]) );
  AND U3722 ( .A(p_input[6651]), .B(p_input[16651]), .Z(o[6651]) );
  AND U3723 ( .A(p_input[6650]), .B(p_input[16650]), .Z(o[6650]) );
  AND U3724 ( .A(p_input[664]), .B(p_input[10664]), .Z(o[664]) );
  AND U3725 ( .A(p_input[6649]), .B(p_input[16649]), .Z(o[6649]) );
  AND U3726 ( .A(p_input[6648]), .B(p_input[16648]), .Z(o[6648]) );
  AND U3727 ( .A(p_input[6647]), .B(p_input[16647]), .Z(o[6647]) );
  AND U3728 ( .A(p_input[6646]), .B(p_input[16646]), .Z(o[6646]) );
  AND U3729 ( .A(p_input[6645]), .B(p_input[16645]), .Z(o[6645]) );
  AND U3730 ( .A(p_input[6644]), .B(p_input[16644]), .Z(o[6644]) );
  AND U3731 ( .A(p_input[6643]), .B(p_input[16643]), .Z(o[6643]) );
  AND U3732 ( .A(p_input[6642]), .B(p_input[16642]), .Z(o[6642]) );
  AND U3733 ( .A(p_input[6641]), .B(p_input[16641]), .Z(o[6641]) );
  AND U3734 ( .A(p_input[6640]), .B(p_input[16640]), .Z(o[6640]) );
  AND U3735 ( .A(p_input[663]), .B(p_input[10663]), .Z(o[663]) );
  AND U3736 ( .A(p_input[6639]), .B(p_input[16639]), .Z(o[6639]) );
  AND U3737 ( .A(p_input[6638]), .B(p_input[16638]), .Z(o[6638]) );
  AND U3738 ( .A(p_input[6637]), .B(p_input[16637]), .Z(o[6637]) );
  AND U3739 ( .A(p_input[6636]), .B(p_input[16636]), .Z(o[6636]) );
  AND U3740 ( .A(p_input[6635]), .B(p_input[16635]), .Z(o[6635]) );
  AND U3741 ( .A(p_input[6634]), .B(p_input[16634]), .Z(o[6634]) );
  AND U3742 ( .A(p_input[6633]), .B(p_input[16633]), .Z(o[6633]) );
  AND U3743 ( .A(p_input[6632]), .B(p_input[16632]), .Z(o[6632]) );
  AND U3744 ( .A(p_input[6631]), .B(p_input[16631]), .Z(o[6631]) );
  AND U3745 ( .A(p_input[6630]), .B(p_input[16630]), .Z(o[6630]) );
  AND U3746 ( .A(p_input[662]), .B(p_input[10662]), .Z(o[662]) );
  AND U3747 ( .A(p_input[6629]), .B(p_input[16629]), .Z(o[6629]) );
  AND U3748 ( .A(p_input[6628]), .B(p_input[16628]), .Z(o[6628]) );
  AND U3749 ( .A(p_input[6627]), .B(p_input[16627]), .Z(o[6627]) );
  AND U3750 ( .A(p_input[6626]), .B(p_input[16626]), .Z(o[6626]) );
  AND U3751 ( .A(p_input[6625]), .B(p_input[16625]), .Z(o[6625]) );
  AND U3752 ( .A(p_input[6624]), .B(p_input[16624]), .Z(o[6624]) );
  AND U3753 ( .A(p_input[6623]), .B(p_input[16623]), .Z(o[6623]) );
  AND U3754 ( .A(p_input[6622]), .B(p_input[16622]), .Z(o[6622]) );
  AND U3755 ( .A(p_input[6621]), .B(p_input[16621]), .Z(o[6621]) );
  AND U3756 ( .A(p_input[6620]), .B(p_input[16620]), .Z(o[6620]) );
  AND U3757 ( .A(p_input[661]), .B(p_input[10661]), .Z(o[661]) );
  AND U3758 ( .A(p_input[6619]), .B(p_input[16619]), .Z(o[6619]) );
  AND U3759 ( .A(p_input[6618]), .B(p_input[16618]), .Z(o[6618]) );
  AND U3760 ( .A(p_input[6617]), .B(p_input[16617]), .Z(o[6617]) );
  AND U3761 ( .A(p_input[6616]), .B(p_input[16616]), .Z(o[6616]) );
  AND U3762 ( .A(p_input[6615]), .B(p_input[16615]), .Z(o[6615]) );
  AND U3763 ( .A(p_input[6614]), .B(p_input[16614]), .Z(o[6614]) );
  AND U3764 ( .A(p_input[6613]), .B(p_input[16613]), .Z(o[6613]) );
  AND U3765 ( .A(p_input[6612]), .B(p_input[16612]), .Z(o[6612]) );
  AND U3766 ( .A(p_input[6611]), .B(p_input[16611]), .Z(o[6611]) );
  AND U3767 ( .A(p_input[6610]), .B(p_input[16610]), .Z(o[6610]) );
  AND U3768 ( .A(p_input[660]), .B(p_input[10660]), .Z(o[660]) );
  AND U3769 ( .A(p_input[6609]), .B(p_input[16609]), .Z(o[6609]) );
  AND U3770 ( .A(p_input[6608]), .B(p_input[16608]), .Z(o[6608]) );
  AND U3771 ( .A(p_input[6607]), .B(p_input[16607]), .Z(o[6607]) );
  AND U3772 ( .A(p_input[6606]), .B(p_input[16606]), .Z(o[6606]) );
  AND U3773 ( .A(p_input[6605]), .B(p_input[16605]), .Z(o[6605]) );
  AND U3774 ( .A(p_input[6604]), .B(p_input[16604]), .Z(o[6604]) );
  AND U3775 ( .A(p_input[6603]), .B(p_input[16603]), .Z(o[6603]) );
  AND U3776 ( .A(p_input[6602]), .B(p_input[16602]), .Z(o[6602]) );
  AND U3777 ( .A(p_input[6601]), .B(p_input[16601]), .Z(o[6601]) );
  AND U3778 ( .A(p_input[6600]), .B(p_input[16600]), .Z(o[6600]) );
  AND U3779 ( .A(p_input[65]), .B(p_input[10065]), .Z(o[65]) );
  AND U3780 ( .A(p_input[659]), .B(p_input[10659]), .Z(o[659]) );
  AND U3781 ( .A(p_input[6599]), .B(p_input[16599]), .Z(o[6599]) );
  AND U3782 ( .A(p_input[6598]), .B(p_input[16598]), .Z(o[6598]) );
  AND U3783 ( .A(p_input[6597]), .B(p_input[16597]), .Z(o[6597]) );
  AND U3784 ( .A(p_input[6596]), .B(p_input[16596]), .Z(o[6596]) );
  AND U3785 ( .A(p_input[6595]), .B(p_input[16595]), .Z(o[6595]) );
  AND U3786 ( .A(p_input[6594]), .B(p_input[16594]), .Z(o[6594]) );
  AND U3787 ( .A(p_input[6593]), .B(p_input[16593]), .Z(o[6593]) );
  AND U3788 ( .A(p_input[6592]), .B(p_input[16592]), .Z(o[6592]) );
  AND U3789 ( .A(p_input[6591]), .B(p_input[16591]), .Z(o[6591]) );
  AND U3790 ( .A(p_input[6590]), .B(p_input[16590]), .Z(o[6590]) );
  AND U3791 ( .A(p_input[658]), .B(p_input[10658]), .Z(o[658]) );
  AND U3792 ( .A(p_input[6589]), .B(p_input[16589]), .Z(o[6589]) );
  AND U3793 ( .A(p_input[6588]), .B(p_input[16588]), .Z(o[6588]) );
  AND U3794 ( .A(p_input[6587]), .B(p_input[16587]), .Z(o[6587]) );
  AND U3795 ( .A(p_input[6586]), .B(p_input[16586]), .Z(o[6586]) );
  AND U3796 ( .A(p_input[6585]), .B(p_input[16585]), .Z(o[6585]) );
  AND U3797 ( .A(p_input[6584]), .B(p_input[16584]), .Z(o[6584]) );
  AND U3798 ( .A(p_input[6583]), .B(p_input[16583]), .Z(o[6583]) );
  AND U3799 ( .A(p_input[6582]), .B(p_input[16582]), .Z(o[6582]) );
  AND U3800 ( .A(p_input[6581]), .B(p_input[16581]), .Z(o[6581]) );
  AND U3801 ( .A(p_input[6580]), .B(p_input[16580]), .Z(o[6580]) );
  AND U3802 ( .A(p_input[657]), .B(p_input[10657]), .Z(o[657]) );
  AND U3803 ( .A(p_input[6579]), .B(p_input[16579]), .Z(o[6579]) );
  AND U3804 ( .A(p_input[6578]), .B(p_input[16578]), .Z(o[6578]) );
  AND U3805 ( .A(p_input[6577]), .B(p_input[16577]), .Z(o[6577]) );
  AND U3806 ( .A(p_input[6576]), .B(p_input[16576]), .Z(o[6576]) );
  AND U3807 ( .A(p_input[6575]), .B(p_input[16575]), .Z(o[6575]) );
  AND U3808 ( .A(p_input[6574]), .B(p_input[16574]), .Z(o[6574]) );
  AND U3809 ( .A(p_input[6573]), .B(p_input[16573]), .Z(o[6573]) );
  AND U3810 ( .A(p_input[6572]), .B(p_input[16572]), .Z(o[6572]) );
  AND U3811 ( .A(p_input[6571]), .B(p_input[16571]), .Z(o[6571]) );
  AND U3812 ( .A(p_input[6570]), .B(p_input[16570]), .Z(o[6570]) );
  AND U3813 ( .A(p_input[656]), .B(p_input[10656]), .Z(o[656]) );
  AND U3814 ( .A(p_input[6569]), .B(p_input[16569]), .Z(o[6569]) );
  AND U3815 ( .A(p_input[6568]), .B(p_input[16568]), .Z(o[6568]) );
  AND U3816 ( .A(p_input[6567]), .B(p_input[16567]), .Z(o[6567]) );
  AND U3817 ( .A(p_input[6566]), .B(p_input[16566]), .Z(o[6566]) );
  AND U3818 ( .A(p_input[6565]), .B(p_input[16565]), .Z(o[6565]) );
  AND U3819 ( .A(p_input[6564]), .B(p_input[16564]), .Z(o[6564]) );
  AND U3820 ( .A(p_input[6563]), .B(p_input[16563]), .Z(o[6563]) );
  AND U3821 ( .A(p_input[6562]), .B(p_input[16562]), .Z(o[6562]) );
  AND U3822 ( .A(p_input[6561]), .B(p_input[16561]), .Z(o[6561]) );
  AND U3823 ( .A(p_input[6560]), .B(p_input[16560]), .Z(o[6560]) );
  AND U3824 ( .A(p_input[655]), .B(p_input[10655]), .Z(o[655]) );
  AND U3825 ( .A(p_input[6559]), .B(p_input[16559]), .Z(o[6559]) );
  AND U3826 ( .A(p_input[6558]), .B(p_input[16558]), .Z(o[6558]) );
  AND U3827 ( .A(p_input[6557]), .B(p_input[16557]), .Z(o[6557]) );
  AND U3828 ( .A(p_input[6556]), .B(p_input[16556]), .Z(o[6556]) );
  AND U3829 ( .A(p_input[6555]), .B(p_input[16555]), .Z(o[6555]) );
  AND U3830 ( .A(p_input[6554]), .B(p_input[16554]), .Z(o[6554]) );
  AND U3831 ( .A(p_input[6553]), .B(p_input[16553]), .Z(o[6553]) );
  AND U3832 ( .A(p_input[6552]), .B(p_input[16552]), .Z(o[6552]) );
  AND U3833 ( .A(p_input[6551]), .B(p_input[16551]), .Z(o[6551]) );
  AND U3834 ( .A(p_input[6550]), .B(p_input[16550]), .Z(o[6550]) );
  AND U3835 ( .A(p_input[654]), .B(p_input[10654]), .Z(o[654]) );
  AND U3836 ( .A(p_input[6549]), .B(p_input[16549]), .Z(o[6549]) );
  AND U3837 ( .A(p_input[6548]), .B(p_input[16548]), .Z(o[6548]) );
  AND U3838 ( .A(p_input[6547]), .B(p_input[16547]), .Z(o[6547]) );
  AND U3839 ( .A(p_input[6546]), .B(p_input[16546]), .Z(o[6546]) );
  AND U3840 ( .A(p_input[6545]), .B(p_input[16545]), .Z(o[6545]) );
  AND U3841 ( .A(p_input[6544]), .B(p_input[16544]), .Z(o[6544]) );
  AND U3842 ( .A(p_input[6543]), .B(p_input[16543]), .Z(o[6543]) );
  AND U3843 ( .A(p_input[6542]), .B(p_input[16542]), .Z(o[6542]) );
  AND U3844 ( .A(p_input[6541]), .B(p_input[16541]), .Z(o[6541]) );
  AND U3845 ( .A(p_input[6540]), .B(p_input[16540]), .Z(o[6540]) );
  AND U3846 ( .A(p_input[653]), .B(p_input[10653]), .Z(o[653]) );
  AND U3847 ( .A(p_input[6539]), .B(p_input[16539]), .Z(o[6539]) );
  AND U3848 ( .A(p_input[6538]), .B(p_input[16538]), .Z(o[6538]) );
  AND U3849 ( .A(p_input[6537]), .B(p_input[16537]), .Z(o[6537]) );
  AND U3850 ( .A(p_input[6536]), .B(p_input[16536]), .Z(o[6536]) );
  AND U3851 ( .A(p_input[6535]), .B(p_input[16535]), .Z(o[6535]) );
  AND U3852 ( .A(p_input[6534]), .B(p_input[16534]), .Z(o[6534]) );
  AND U3853 ( .A(p_input[6533]), .B(p_input[16533]), .Z(o[6533]) );
  AND U3854 ( .A(p_input[6532]), .B(p_input[16532]), .Z(o[6532]) );
  AND U3855 ( .A(p_input[6531]), .B(p_input[16531]), .Z(o[6531]) );
  AND U3856 ( .A(p_input[6530]), .B(p_input[16530]), .Z(o[6530]) );
  AND U3857 ( .A(p_input[652]), .B(p_input[10652]), .Z(o[652]) );
  AND U3858 ( .A(p_input[6529]), .B(p_input[16529]), .Z(o[6529]) );
  AND U3859 ( .A(p_input[6528]), .B(p_input[16528]), .Z(o[6528]) );
  AND U3860 ( .A(p_input[6527]), .B(p_input[16527]), .Z(o[6527]) );
  AND U3861 ( .A(p_input[6526]), .B(p_input[16526]), .Z(o[6526]) );
  AND U3862 ( .A(p_input[6525]), .B(p_input[16525]), .Z(o[6525]) );
  AND U3863 ( .A(p_input[6524]), .B(p_input[16524]), .Z(o[6524]) );
  AND U3864 ( .A(p_input[6523]), .B(p_input[16523]), .Z(o[6523]) );
  AND U3865 ( .A(p_input[6522]), .B(p_input[16522]), .Z(o[6522]) );
  AND U3866 ( .A(p_input[6521]), .B(p_input[16521]), .Z(o[6521]) );
  AND U3867 ( .A(p_input[6520]), .B(p_input[16520]), .Z(o[6520]) );
  AND U3868 ( .A(p_input[651]), .B(p_input[10651]), .Z(o[651]) );
  AND U3869 ( .A(p_input[6519]), .B(p_input[16519]), .Z(o[6519]) );
  AND U3870 ( .A(p_input[6518]), .B(p_input[16518]), .Z(o[6518]) );
  AND U3871 ( .A(p_input[6517]), .B(p_input[16517]), .Z(o[6517]) );
  AND U3872 ( .A(p_input[6516]), .B(p_input[16516]), .Z(o[6516]) );
  AND U3873 ( .A(p_input[6515]), .B(p_input[16515]), .Z(o[6515]) );
  AND U3874 ( .A(p_input[6514]), .B(p_input[16514]), .Z(o[6514]) );
  AND U3875 ( .A(p_input[6513]), .B(p_input[16513]), .Z(o[6513]) );
  AND U3876 ( .A(p_input[6512]), .B(p_input[16512]), .Z(o[6512]) );
  AND U3877 ( .A(p_input[6511]), .B(p_input[16511]), .Z(o[6511]) );
  AND U3878 ( .A(p_input[6510]), .B(p_input[16510]), .Z(o[6510]) );
  AND U3879 ( .A(p_input[650]), .B(p_input[10650]), .Z(o[650]) );
  AND U3880 ( .A(p_input[6509]), .B(p_input[16509]), .Z(o[6509]) );
  AND U3881 ( .A(p_input[6508]), .B(p_input[16508]), .Z(o[6508]) );
  AND U3882 ( .A(p_input[6507]), .B(p_input[16507]), .Z(o[6507]) );
  AND U3883 ( .A(p_input[6506]), .B(p_input[16506]), .Z(o[6506]) );
  AND U3884 ( .A(p_input[6505]), .B(p_input[16505]), .Z(o[6505]) );
  AND U3885 ( .A(p_input[6504]), .B(p_input[16504]), .Z(o[6504]) );
  AND U3886 ( .A(p_input[6503]), .B(p_input[16503]), .Z(o[6503]) );
  AND U3887 ( .A(p_input[6502]), .B(p_input[16502]), .Z(o[6502]) );
  AND U3888 ( .A(p_input[6501]), .B(p_input[16501]), .Z(o[6501]) );
  AND U3889 ( .A(p_input[6500]), .B(p_input[16500]), .Z(o[6500]) );
  AND U3890 ( .A(p_input[64]), .B(p_input[10064]), .Z(o[64]) );
  AND U3891 ( .A(p_input[649]), .B(p_input[10649]), .Z(o[649]) );
  AND U3892 ( .A(p_input[6499]), .B(p_input[16499]), .Z(o[6499]) );
  AND U3893 ( .A(p_input[6498]), .B(p_input[16498]), .Z(o[6498]) );
  AND U3894 ( .A(p_input[6497]), .B(p_input[16497]), .Z(o[6497]) );
  AND U3895 ( .A(p_input[6496]), .B(p_input[16496]), .Z(o[6496]) );
  AND U3896 ( .A(p_input[6495]), .B(p_input[16495]), .Z(o[6495]) );
  AND U3897 ( .A(p_input[6494]), .B(p_input[16494]), .Z(o[6494]) );
  AND U3898 ( .A(p_input[6493]), .B(p_input[16493]), .Z(o[6493]) );
  AND U3899 ( .A(p_input[6492]), .B(p_input[16492]), .Z(o[6492]) );
  AND U3900 ( .A(p_input[6491]), .B(p_input[16491]), .Z(o[6491]) );
  AND U3901 ( .A(p_input[6490]), .B(p_input[16490]), .Z(o[6490]) );
  AND U3902 ( .A(p_input[648]), .B(p_input[10648]), .Z(o[648]) );
  AND U3903 ( .A(p_input[6489]), .B(p_input[16489]), .Z(o[6489]) );
  AND U3904 ( .A(p_input[6488]), .B(p_input[16488]), .Z(o[6488]) );
  AND U3905 ( .A(p_input[6487]), .B(p_input[16487]), .Z(o[6487]) );
  AND U3906 ( .A(p_input[6486]), .B(p_input[16486]), .Z(o[6486]) );
  AND U3907 ( .A(p_input[6485]), .B(p_input[16485]), .Z(o[6485]) );
  AND U3908 ( .A(p_input[6484]), .B(p_input[16484]), .Z(o[6484]) );
  AND U3909 ( .A(p_input[6483]), .B(p_input[16483]), .Z(o[6483]) );
  AND U3910 ( .A(p_input[6482]), .B(p_input[16482]), .Z(o[6482]) );
  AND U3911 ( .A(p_input[6481]), .B(p_input[16481]), .Z(o[6481]) );
  AND U3912 ( .A(p_input[6480]), .B(p_input[16480]), .Z(o[6480]) );
  AND U3913 ( .A(p_input[647]), .B(p_input[10647]), .Z(o[647]) );
  AND U3914 ( .A(p_input[6479]), .B(p_input[16479]), .Z(o[6479]) );
  AND U3915 ( .A(p_input[6478]), .B(p_input[16478]), .Z(o[6478]) );
  AND U3916 ( .A(p_input[6477]), .B(p_input[16477]), .Z(o[6477]) );
  AND U3917 ( .A(p_input[6476]), .B(p_input[16476]), .Z(o[6476]) );
  AND U3918 ( .A(p_input[6475]), .B(p_input[16475]), .Z(o[6475]) );
  AND U3919 ( .A(p_input[6474]), .B(p_input[16474]), .Z(o[6474]) );
  AND U3920 ( .A(p_input[6473]), .B(p_input[16473]), .Z(o[6473]) );
  AND U3921 ( .A(p_input[6472]), .B(p_input[16472]), .Z(o[6472]) );
  AND U3922 ( .A(p_input[6471]), .B(p_input[16471]), .Z(o[6471]) );
  AND U3923 ( .A(p_input[6470]), .B(p_input[16470]), .Z(o[6470]) );
  AND U3924 ( .A(p_input[646]), .B(p_input[10646]), .Z(o[646]) );
  AND U3925 ( .A(p_input[6469]), .B(p_input[16469]), .Z(o[6469]) );
  AND U3926 ( .A(p_input[6468]), .B(p_input[16468]), .Z(o[6468]) );
  AND U3927 ( .A(p_input[6467]), .B(p_input[16467]), .Z(o[6467]) );
  AND U3928 ( .A(p_input[6466]), .B(p_input[16466]), .Z(o[6466]) );
  AND U3929 ( .A(p_input[6465]), .B(p_input[16465]), .Z(o[6465]) );
  AND U3930 ( .A(p_input[6464]), .B(p_input[16464]), .Z(o[6464]) );
  AND U3931 ( .A(p_input[6463]), .B(p_input[16463]), .Z(o[6463]) );
  AND U3932 ( .A(p_input[6462]), .B(p_input[16462]), .Z(o[6462]) );
  AND U3933 ( .A(p_input[6461]), .B(p_input[16461]), .Z(o[6461]) );
  AND U3934 ( .A(p_input[6460]), .B(p_input[16460]), .Z(o[6460]) );
  AND U3935 ( .A(p_input[645]), .B(p_input[10645]), .Z(o[645]) );
  AND U3936 ( .A(p_input[6459]), .B(p_input[16459]), .Z(o[6459]) );
  AND U3937 ( .A(p_input[6458]), .B(p_input[16458]), .Z(o[6458]) );
  AND U3938 ( .A(p_input[6457]), .B(p_input[16457]), .Z(o[6457]) );
  AND U3939 ( .A(p_input[6456]), .B(p_input[16456]), .Z(o[6456]) );
  AND U3940 ( .A(p_input[6455]), .B(p_input[16455]), .Z(o[6455]) );
  AND U3941 ( .A(p_input[6454]), .B(p_input[16454]), .Z(o[6454]) );
  AND U3942 ( .A(p_input[6453]), .B(p_input[16453]), .Z(o[6453]) );
  AND U3943 ( .A(p_input[6452]), .B(p_input[16452]), .Z(o[6452]) );
  AND U3944 ( .A(p_input[6451]), .B(p_input[16451]), .Z(o[6451]) );
  AND U3945 ( .A(p_input[6450]), .B(p_input[16450]), .Z(o[6450]) );
  AND U3946 ( .A(p_input[644]), .B(p_input[10644]), .Z(o[644]) );
  AND U3947 ( .A(p_input[6449]), .B(p_input[16449]), .Z(o[6449]) );
  AND U3948 ( .A(p_input[6448]), .B(p_input[16448]), .Z(o[6448]) );
  AND U3949 ( .A(p_input[6447]), .B(p_input[16447]), .Z(o[6447]) );
  AND U3950 ( .A(p_input[6446]), .B(p_input[16446]), .Z(o[6446]) );
  AND U3951 ( .A(p_input[6445]), .B(p_input[16445]), .Z(o[6445]) );
  AND U3952 ( .A(p_input[6444]), .B(p_input[16444]), .Z(o[6444]) );
  AND U3953 ( .A(p_input[6443]), .B(p_input[16443]), .Z(o[6443]) );
  AND U3954 ( .A(p_input[6442]), .B(p_input[16442]), .Z(o[6442]) );
  AND U3955 ( .A(p_input[6441]), .B(p_input[16441]), .Z(o[6441]) );
  AND U3956 ( .A(p_input[6440]), .B(p_input[16440]), .Z(o[6440]) );
  AND U3957 ( .A(p_input[643]), .B(p_input[10643]), .Z(o[643]) );
  AND U3958 ( .A(p_input[6439]), .B(p_input[16439]), .Z(o[6439]) );
  AND U3959 ( .A(p_input[6438]), .B(p_input[16438]), .Z(o[6438]) );
  AND U3960 ( .A(p_input[6437]), .B(p_input[16437]), .Z(o[6437]) );
  AND U3961 ( .A(p_input[6436]), .B(p_input[16436]), .Z(o[6436]) );
  AND U3962 ( .A(p_input[6435]), .B(p_input[16435]), .Z(o[6435]) );
  AND U3963 ( .A(p_input[6434]), .B(p_input[16434]), .Z(o[6434]) );
  AND U3964 ( .A(p_input[6433]), .B(p_input[16433]), .Z(o[6433]) );
  AND U3965 ( .A(p_input[6432]), .B(p_input[16432]), .Z(o[6432]) );
  AND U3966 ( .A(p_input[6431]), .B(p_input[16431]), .Z(o[6431]) );
  AND U3967 ( .A(p_input[6430]), .B(p_input[16430]), .Z(o[6430]) );
  AND U3968 ( .A(p_input[642]), .B(p_input[10642]), .Z(o[642]) );
  AND U3969 ( .A(p_input[6429]), .B(p_input[16429]), .Z(o[6429]) );
  AND U3970 ( .A(p_input[6428]), .B(p_input[16428]), .Z(o[6428]) );
  AND U3971 ( .A(p_input[6427]), .B(p_input[16427]), .Z(o[6427]) );
  AND U3972 ( .A(p_input[6426]), .B(p_input[16426]), .Z(o[6426]) );
  AND U3973 ( .A(p_input[6425]), .B(p_input[16425]), .Z(o[6425]) );
  AND U3974 ( .A(p_input[6424]), .B(p_input[16424]), .Z(o[6424]) );
  AND U3975 ( .A(p_input[6423]), .B(p_input[16423]), .Z(o[6423]) );
  AND U3976 ( .A(p_input[6422]), .B(p_input[16422]), .Z(o[6422]) );
  AND U3977 ( .A(p_input[6421]), .B(p_input[16421]), .Z(o[6421]) );
  AND U3978 ( .A(p_input[6420]), .B(p_input[16420]), .Z(o[6420]) );
  AND U3979 ( .A(p_input[641]), .B(p_input[10641]), .Z(o[641]) );
  AND U3980 ( .A(p_input[6419]), .B(p_input[16419]), .Z(o[6419]) );
  AND U3981 ( .A(p_input[6418]), .B(p_input[16418]), .Z(o[6418]) );
  AND U3982 ( .A(p_input[6417]), .B(p_input[16417]), .Z(o[6417]) );
  AND U3983 ( .A(p_input[6416]), .B(p_input[16416]), .Z(o[6416]) );
  AND U3984 ( .A(p_input[6415]), .B(p_input[16415]), .Z(o[6415]) );
  AND U3985 ( .A(p_input[6414]), .B(p_input[16414]), .Z(o[6414]) );
  AND U3986 ( .A(p_input[6413]), .B(p_input[16413]), .Z(o[6413]) );
  AND U3987 ( .A(p_input[6412]), .B(p_input[16412]), .Z(o[6412]) );
  AND U3988 ( .A(p_input[6411]), .B(p_input[16411]), .Z(o[6411]) );
  AND U3989 ( .A(p_input[6410]), .B(p_input[16410]), .Z(o[6410]) );
  AND U3990 ( .A(p_input[640]), .B(p_input[10640]), .Z(o[640]) );
  AND U3991 ( .A(p_input[6409]), .B(p_input[16409]), .Z(o[6409]) );
  AND U3992 ( .A(p_input[6408]), .B(p_input[16408]), .Z(o[6408]) );
  AND U3993 ( .A(p_input[6407]), .B(p_input[16407]), .Z(o[6407]) );
  AND U3994 ( .A(p_input[6406]), .B(p_input[16406]), .Z(o[6406]) );
  AND U3995 ( .A(p_input[6405]), .B(p_input[16405]), .Z(o[6405]) );
  AND U3996 ( .A(p_input[6404]), .B(p_input[16404]), .Z(o[6404]) );
  AND U3997 ( .A(p_input[6403]), .B(p_input[16403]), .Z(o[6403]) );
  AND U3998 ( .A(p_input[6402]), .B(p_input[16402]), .Z(o[6402]) );
  AND U3999 ( .A(p_input[6401]), .B(p_input[16401]), .Z(o[6401]) );
  AND U4000 ( .A(p_input[6400]), .B(p_input[16400]), .Z(o[6400]) );
  AND U4001 ( .A(p_input[63]), .B(p_input[10063]), .Z(o[63]) );
  AND U4002 ( .A(p_input[639]), .B(p_input[10639]), .Z(o[639]) );
  AND U4003 ( .A(p_input[6399]), .B(p_input[16399]), .Z(o[6399]) );
  AND U4004 ( .A(p_input[6398]), .B(p_input[16398]), .Z(o[6398]) );
  AND U4005 ( .A(p_input[6397]), .B(p_input[16397]), .Z(o[6397]) );
  AND U4006 ( .A(p_input[6396]), .B(p_input[16396]), .Z(o[6396]) );
  AND U4007 ( .A(p_input[6395]), .B(p_input[16395]), .Z(o[6395]) );
  AND U4008 ( .A(p_input[6394]), .B(p_input[16394]), .Z(o[6394]) );
  AND U4009 ( .A(p_input[6393]), .B(p_input[16393]), .Z(o[6393]) );
  AND U4010 ( .A(p_input[6392]), .B(p_input[16392]), .Z(o[6392]) );
  AND U4011 ( .A(p_input[6391]), .B(p_input[16391]), .Z(o[6391]) );
  AND U4012 ( .A(p_input[6390]), .B(p_input[16390]), .Z(o[6390]) );
  AND U4013 ( .A(p_input[638]), .B(p_input[10638]), .Z(o[638]) );
  AND U4014 ( .A(p_input[6389]), .B(p_input[16389]), .Z(o[6389]) );
  AND U4015 ( .A(p_input[6388]), .B(p_input[16388]), .Z(o[6388]) );
  AND U4016 ( .A(p_input[6387]), .B(p_input[16387]), .Z(o[6387]) );
  AND U4017 ( .A(p_input[6386]), .B(p_input[16386]), .Z(o[6386]) );
  AND U4018 ( .A(p_input[6385]), .B(p_input[16385]), .Z(o[6385]) );
  AND U4019 ( .A(p_input[6384]), .B(p_input[16384]), .Z(o[6384]) );
  AND U4020 ( .A(p_input[6383]), .B(p_input[16383]), .Z(o[6383]) );
  AND U4021 ( .A(p_input[6382]), .B(p_input[16382]), .Z(o[6382]) );
  AND U4022 ( .A(p_input[6381]), .B(p_input[16381]), .Z(o[6381]) );
  AND U4023 ( .A(p_input[6380]), .B(p_input[16380]), .Z(o[6380]) );
  AND U4024 ( .A(p_input[637]), .B(p_input[10637]), .Z(o[637]) );
  AND U4025 ( .A(p_input[6379]), .B(p_input[16379]), .Z(o[6379]) );
  AND U4026 ( .A(p_input[6378]), .B(p_input[16378]), .Z(o[6378]) );
  AND U4027 ( .A(p_input[6377]), .B(p_input[16377]), .Z(o[6377]) );
  AND U4028 ( .A(p_input[6376]), .B(p_input[16376]), .Z(o[6376]) );
  AND U4029 ( .A(p_input[6375]), .B(p_input[16375]), .Z(o[6375]) );
  AND U4030 ( .A(p_input[6374]), .B(p_input[16374]), .Z(o[6374]) );
  AND U4031 ( .A(p_input[6373]), .B(p_input[16373]), .Z(o[6373]) );
  AND U4032 ( .A(p_input[6372]), .B(p_input[16372]), .Z(o[6372]) );
  AND U4033 ( .A(p_input[6371]), .B(p_input[16371]), .Z(o[6371]) );
  AND U4034 ( .A(p_input[6370]), .B(p_input[16370]), .Z(o[6370]) );
  AND U4035 ( .A(p_input[636]), .B(p_input[10636]), .Z(o[636]) );
  AND U4036 ( .A(p_input[6369]), .B(p_input[16369]), .Z(o[6369]) );
  AND U4037 ( .A(p_input[6368]), .B(p_input[16368]), .Z(o[6368]) );
  AND U4038 ( .A(p_input[6367]), .B(p_input[16367]), .Z(o[6367]) );
  AND U4039 ( .A(p_input[6366]), .B(p_input[16366]), .Z(o[6366]) );
  AND U4040 ( .A(p_input[6365]), .B(p_input[16365]), .Z(o[6365]) );
  AND U4041 ( .A(p_input[6364]), .B(p_input[16364]), .Z(o[6364]) );
  AND U4042 ( .A(p_input[6363]), .B(p_input[16363]), .Z(o[6363]) );
  AND U4043 ( .A(p_input[6362]), .B(p_input[16362]), .Z(o[6362]) );
  AND U4044 ( .A(p_input[6361]), .B(p_input[16361]), .Z(o[6361]) );
  AND U4045 ( .A(p_input[6360]), .B(p_input[16360]), .Z(o[6360]) );
  AND U4046 ( .A(p_input[635]), .B(p_input[10635]), .Z(o[635]) );
  AND U4047 ( .A(p_input[6359]), .B(p_input[16359]), .Z(o[6359]) );
  AND U4048 ( .A(p_input[6358]), .B(p_input[16358]), .Z(o[6358]) );
  AND U4049 ( .A(p_input[6357]), .B(p_input[16357]), .Z(o[6357]) );
  AND U4050 ( .A(p_input[6356]), .B(p_input[16356]), .Z(o[6356]) );
  AND U4051 ( .A(p_input[6355]), .B(p_input[16355]), .Z(o[6355]) );
  AND U4052 ( .A(p_input[6354]), .B(p_input[16354]), .Z(o[6354]) );
  AND U4053 ( .A(p_input[6353]), .B(p_input[16353]), .Z(o[6353]) );
  AND U4054 ( .A(p_input[6352]), .B(p_input[16352]), .Z(o[6352]) );
  AND U4055 ( .A(p_input[6351]), .B(p_input[16351]), .Z(o[6351]) );
  AND U4056 ( .A(p_input[6350]), .B(p_input[16350]), .Z(o[6350]) );
  AND U4057 ( .A(p_input[634]), .B(p_input[10634]), .Z(o[634]) );
  AND U4058 ( .A(p_input[6349]), .B(p_input[16349]), .Z(o[6349]) );
  AND U4059 ( .A(p_input[6348]), .B(p_input[16348]), .Z(o[6348]) );
  AND U4060 ( .A(p_input[6347]), .B(p_input[16347]), .Z(o[6347]) );
  AND U4061 ( .A(p_input[6346]), .B(p_input[16346]), .Z(o[6346]) );
  AND U4062 ( .A(p_input[6345]), .B(p_input[16345]), .Z(o[6345]) );
  AND U4063 ( .A(p_input[6344]), .B(p_input[16344]), .Z(o[6344]) );
  AND U4064 ( .A(p_input[6343]), .B(p_input[16343]), .Z(o[6343]) );
  AND U4065 ( .A(p_input[6342]), .B(p_input[16342]), .Z(o[6342]) );
  AND U4066 ( .A(p_input[6341]), .B(p_input[16341]), .Z(o[6341]) );
  AND U4067 ( .A(p_input[6340]), .B(p_input[16340]), .Z(o[6340]) );
  AND U4068 ( .A(p_input[633]), .B(p_input[10633]), .Z(o[633]) );
  AND U4069 ( .A(p_input[6339]), .B(p_input[16339]), .Z(o[6339]) );
  AND U4070 ( .A(p_input[6338]), .B(p_input[16338]), .Z(o[6338]) );
  AND U4071 ( .A(p_input[6337]), .B(p_input[16337]), .Z(o[6337]) );
  AND U4072 ( .A(p_input[6336]), .B(p_input[16336]), .Z(o[6336]) );
  AND U4073 ( .A(p_input[6335]), .B(p_input[16335]), .Z(o[6335]) );
  AND U4074 ( .A(p_input[6334]), .B(p_input[16334]), .Z(o[6334]) );
  AND U4075 ( .A(p_input[6333]), .B(p_input[16333]), .Z(o[6333]) );
  AND U4076 ( .A(p_input[6332]), .B(p_input[16332]), .Z(o[6332]) );
  AND U4077 ( .A(p_input[6331]), .B(p_input[16331]), .Z(o[6331]) );
  AND U4078 ( .A(p_input[6330]), .B(p_input[16330]), .Z(o[6330]) );
  AND U4079 ( .A(p_input[632]), .B(p_input[10632]), .Z(o[632]) );
  AND U4080 ( .A(p_input[6329]), .B(p_input[16329]), .Z(o[6329]) );
  AND U4081 ( .A(p_input[6328]), .B(p_input[16328]), .Z(o[6328]) );
  AND U4082 ( .A(p_input[6327]), .B(p_input[16327]), .Z(o[6327]) );
  AND U4083 ( .A(p_input[6326]), .B(p_input[16326]), .Z(o[6326]) );
  AND U4084 ( .A(p_input[6325]), .B(p_input[16325]), .Z(o[6325]) );
  AND U4085 ( .A(p_input[6324]), .B(p_input[16324]), .Z(o[6324]) );
  AND U4086 ( .A(p_input[6323]), .B(p_input[16323]), .Z(o[6323]) );
  AND U4087 ( .A(p_input[6322]), .B(p_input[16322]), .Z(o[6322]) );
  AND U4088 ( .A(p_input[6321]), .B(p_input[16321]), .Z(o[6321]) );
  AND U4089 ( .A(p_input[6320]), .B(p_input[16320]), .Z(o[6320]) );
  AND U4090 ( .A(p_input[631]), .B(p_input[10631]), .Z(o[631]) );
  AND U4091 ( .A(p_input[6319]), .B(p_input[16319]), .Z(o[6319]) );
  AND U4092 ( .A(p_input[6318]), .B(p_input[16318]), .Z(o[6318]) );
  AND U4093 ( .A(p_input[6317]), .B(p_input[16317]), .Z(o[6317]) );
  AND U4094 ( .A(p_input[6316]), .B(p_input[16316]), .Z(o[6316]) );
  AND U4095 ( .A(p_input[6315]), .B(p_input[16315]), .Z(o[6315]) );
  AND U4096 ( .A(p_input[6314]), .B(p_input[16314]), .Z(o[6314]) );
  AND U4097 ( .A(p_input[6313]), .B(p_input[16313]), .Z(o[6313]) );
  AND U4098 ( .A(p_input[6312]), .B(p_input[16312]), .Z(o[6312]) );
  AND U4099 ( .A(p_input[6311]), .B(p_input[16311]), .Z(o[6311]) );
  AND U4100 ( .A(p_input[6310]), .B(p_input[16310]), .Z(o[6310]) );
  AND U4101 ( .A(p_input[630]), .B(p_input[10630]), .Z(o[630]) );
  AND U4102 ( .A(p_input[6309]), .B(p_input[16309]), .Z(o[6309]) );
  AND U4103 ( .A(p_input[6308]), .B(p_input[16308]), .Z(o[6308]) );
  AND U4104 ( .A(p_input[6307]), .B(p_input[16307]), .Z(o[6307]) );
  AND U4105 ( .A(p_input[6306]), .B(p_input[16306]), .Z(o[6306]) );
  AND U4106 ( .A(p_input[6305]), .B(p_input[16305]), .Z(o[6305]) );
  AND U4107 ( .A(p_input[6304]), .B(p_input[16304]), .Z(o[6304]) );
  AND U4108 ( .A(p_input[6303]), .B(p_input[16303]), .Z(o[6303]) );
  AND U4109 ( .A(p_input[6302]), .B(p_input[16302]), .Z(o[6302]) );
  AND U4110 ( .A(p_input[6301]), .B(p_input[16301]), .Z(o[6301]) );
  AND U4111 ( .A(p_input[6300]), .B(p_input[16300]), .Z(o[6300]) );
  AND U4112 ( .A(p_input[62]), .B(p_input[10062]), .Z(o[62]) );
  AND U4113 ( .A(p_input[629]), .B(p_input[10629]), .Z(o[629]) );
  AND U4114 ( .A(p_input[6299]), .B(p_input[16299]), .Z(o[6299]) );
  AND U4115 ( .A(p_input[6298]), .B(p_input[16298]), .Z(o[6298]) );
  AND U4116 ( .A(p_input[6297]), .B(p_input[16297]), .Z(o[6297]) );
  AND U4117 ( .A(p_input[6296]), .B(p_input[16296]), .Z(o[6296]) );
  AND U4118 ( .A(p_input[6295]), .B(p_input[16295]), .Z(o[6295]) );
  AND U4119 ( .A(p_input[6294]), .B(p_input[16294]), .Z(o[6294]) );
  AND U4120 ( .A(p_input[6293]), .B(p_input[16293]), .Z(o[6293]) );
  AND U4121 ( .A(p_input[6292]), .B(p_input[16292]), .Z(o[6292]) );
  AND U4122 ( .A(p_input[6291]), .B(p_input[16291]), .Z(o[6291]) );
  AND U4123 ( .A(p_input[6290]), .B(p_input[16290]), .Z(o[6290]) );
  AND U4124 ( .A(p_input[628]), .B(p_input[10628]), .Z(o[628]) );
  AND U4125 ( .A(p_input[6289]), .B(p_input[16289]), .Z(o[6289]) );
  AND U4126 ( .A(p_input[6288]), .B(p_input[16288]), .Z(o[6288]) );
  AND U4127 ( .A(p_input[6287]), .B(p_input[16287]), .Z(o[6287]) );
  AND U4128 ( .A(p_input[6286]), .B(p_input[16286]), .Z(o[6286]) );
  AND U4129 ( .A(p_input[6285]), .B(p_input[16285]), .Z(o[6285]) );
  AND U4130 ( .A(p_input[6284]), .B(p_input[16284]), .Z(o[6284]) );
  AND U4131 ( .A(p_input[6283]), .B(p_input[16283]), .Z(o[6283]) );
  AND U4132 ( .A(p_input[6282]), .B(p_input[16282]), .Z(o[6282]) );
  AND U4133 ( .A(p_input[6281]), .B(p_input[16281]), .Z(o[6281]) );
  AND U4134 ( .A(p_input[6280]), .B(p_input[16280]), .Z(o[6280]) );
  AND U4135 ( .A(p_input[627]), .B(p_input[10627]), .Z(o[627]) );
  AND U4136 ( .A(p_input[6279]), .B(p_input[16279]), .Z(o[6279]) );
  AND U4137 ( .A(p_input[6278]), .B(p_input[16278]), .Z(o[6278]) );
  AND U4138 ( .A(p_input[6277]), .B(p_input[16277]), .Z(o[6277]) );
  AND U4139 ( .A(p_input[6276]), .B(p_input[16276]), .Z(o[6276]) );
  AND U4140 ( .A(p_input[6275]), .B(p_input[16275]), .Z(o[6275]) );
  AND U4141 ( .A(p_input[6274]), .B(p_input[16274]), .Z(o[6274]) );
  AND U4142 ( .A(p_input[6273]), .B(p_input[16273]), .Z(o[6273]) );
  AND U4143 ( .A(p_input[6272]), .B(p_input[16272]), .Z(o[6272]) );
  AND U4144 ( .A(p_input[6271]), .B(p_input[16271]), .Z(o[6271]) );
  AND U4145 ( .A(p_input[6270]), .B(p_input[16270]), .Z(o[6270]) );
  AND U4146 ( .A(p_input[626]), .B(p_input[10626]), .Z(o[626]) );
  AND U4147 ( .A(p_input[6269]), .B(p_input[16269]), .Z(o[6269]) );
  AND U4148 ( .A(p_input[6268]), .B(p_input[16268]), .Z(o[6268]) );
  AND U4149 ( .A(p_input[6267]), .B(p_input[16267]), .Z(o[6267]) );
  AND U4150 ( .A(p_input[6266]), .B(p_input[16266]), .Z(o[6266]) );
  AND U4151 ( .A(p_input[6265]), .B(p_input[16265]), .Z(o[6265]) );
  AND U4152 ( .A(p_input[6264]), .B(p_input[16264]), .Z(o[6264]) );
  AND U4153 ( .A(p_input[6263]), .B(p_input[16263]), .Z(o[6263]) );
  AND U4154 ( .A(p_input[6262]), .B(p_input[16262]), .Z(o[6262]) );
  AND U4155 ( .A(p_input[6261]), .B(p_input[16261]), .Z(o[6261]) );
  AND U4156 ( .A(p_input[6260]), .B(p_input[16260]), .Z(o[6260]) );
  AND U4157 ( .A(p_input[625]), .B(p_input[10625]), .Z(o[625]) );
  AND U4158 ( .A(p_input[6259]), .B(p_input[16259]), .Z(o[6259]) );
  AND U4159 ( .A(p_input[6258]), .B(p_input[16258]), .Z(o[6258]) );
  AND U4160 ( .A(p_input[6257]), .B(p_input[16257]), .Z(o[6257]) );
  AND U4161 ( .A(p_input[6256]), .B(p_input[16256]), .Z(o[6256]) );
  AND U4162 ( .A(p_input[6255]), .B(p_input[16255]), .Z(o[6255]) );
  AND U4163 ( .A(p_input[6254]), .B(p_input[16254]), .Z(o[6254]) );
  AND U4164 ( .A(p_input[6253]), .B(p_input[16253]), .Z(o[6253]) );
  AND U4165 ( .A(p_input[6252]), .B(p_input[16252]), .Z(o[6252]) );
  AND U4166 ( .A(p_input[6251]), .B(p_input[16251]), .Z(o[6251]) );
  AND U4167 ( .A(p_input[6250]), .B(p_input[16250]), .Z(o[6250]) );
  AND U4168 ( .A(p_input[624]), .B(p_input[10624]), .Z(o[624]) );
  AND U4169 ( .A(p_input[6249]), .B(p_input[16249]), .Z(o[6249]) );
  AND U4170 ( .A(p_input[6248]), .B(p_input[16248]), .Z(o[6248]) );
  AND U4171 ( .A(p_input[6247]), .B(p_input[16247]), .Z(o[6247]) );
  AND U4172 ( .A(p_input[6246]), .B(p_input[16246]), .Z(o[6246]) );
  AND U4173 ( .A(p_input[6245]), .B(p_input[16245]), .Z(o[6245]) );
  AND U4174 ( .A(p_input[6244]), .B(p_input[16244]), .Z(o[6244]) );
  AND U4175 ( .A(p_input[6243]), .B(p_input[16243]), .Z(o[6243]) );
  AND U4176 ( .A(p_input[6242]), .B(p_input[16242]), .Z(o[6242]) );
  AND U4177 ( .A(p_input[6241]), .B(p_input[16241]), .Z(o[6241]) );
  AND U4178 ( .A(p_input[6240]), .B(p_input[16240]), .Z(o[6240]) );
  AND U4179 ( .A(p_input[623]), .B(p_input[10623]), .Z(o[623]) );
  AND U4180 ( .A(p_input[6239]), .B(p_input[16239]), .Z(o[6239]) );
  AND U4181 ( .A(p_input[6238]), .B(p_input[16238]), .Z(o[6238]) );
  AND U4182 ( .A(p_input[6237]), .B(p_input[16237]), .Z(o[6237]) );
  AND U4183 ( .A(p_input[6236]), .B(p_input[16236]), .Z(o[6236]) );
  AND U4184 ( .A(p_input[6235]), .B(p_input[16235]), .Z(o[6235]) );
  AND U4185 ( .A(p_input[6234]), .B(p_input[16234]), .Z(o[6234]) );
  AND U4186 ( .A(p_input[6233]), .B(p_input[16233]), .Z(o[6233]) );
  AND U4187 ( .A(p_input[6232]), .B(p_input[16232]), .Z(o[6232]) );
  AND U4188 ( .A(p_input[6231]), .B(p_input[16231]), .Z(o[6231]) );
  AND U4189 ( .A(p_input[6230]), .B(p_input[16230]), .Z(o[6230]) );
  AND U4190 ( .A(p_input[622]), .B(p_input[10622]), .Z(o[622]) );
  AND U4191 ( .A(p_input[6229]), .B(p_input[16229]), .Z(o[6229]) );
  AND U4192 ( .A(p_input[6228]), .B(p_input[16228]), .Z(o[6228]) );
  AND U4193 ( .A(p_input[6227]), .B(p_input[16227]), .Z(o[6227]) );
  AND U4194 ( .A(p_input[6226]), .B(p_input[16226]), .Z(o[6226]) );
  AND U4195 ( .A(p_input[6225]), .B(p_input[16225]), .Z(o[6225]) );
  AND U4196 ( .A(p_input[6224]), .B(p_input[16224]), .Z(o[6224]) );
  AND U4197 ( .A(p_input[6223]), .B(p_input[16223]), .Z(o[6223]) );
  AND U4198 ( .A(p_input[6222]), .B(p_input[16222]), .Z(o[6222]) );
  AND U4199 ( .A(p_input[6221]), .B(p_input[16221]), .Z(o[6221]) );
  AND U4200 ( .A(p_input[6220]), .B(p_input[16220]), .Z(o[6220]) );
  AND U4201 ( .A(p_input[621]), .B(p_input[10621]), .Z(o[621]) );
  AND U4202 ( .A(p_input[6219]), .B(p_input[16219]), .Z(o[6219]) );
  AND U4203 ( .A(p_input[6218]), .B(p_input[16218]), .Z(o[6218]) );
  AND U4204 ( .A(p_input[6217]), .B(p_input[16217]), .Z(o[6217]) );
  AND U4205 ( .A(p_input[6216]), .B(p_input[16216]), .Z(o[6216]) );
  AND U4206 ( .A(p_input[6215]), .B(p_input[16215]), .Z(o[6215]) );
  AND U4207 ( .A(p_input[6214]), .B(p_input[16214]), .Z(o[6214]) );
  AND U4208 ( .A(p_input[6213]), .B(p_input[16213]), .Z(o[6213]) );
  AND U4209 ( .A(p_input[6212]), .B(p_input[16212]), .Z(o[6212]) );
  AND U4210 ( .A(p_input[6211]), .B(p_input[16211]), .Z(o[6211]) );
  AND U4211 ( .A(p_input[6210]), .B(p_input[16210]), .Z(o[6210]) );
  AND U4212 ( .A(p_input[620]), .B(p_input[10620]), .Z(o[620]) );
  AND U4213 ( .A(p_input[6209]), .B(p_input[16209]), .Z(o[6209]) );
  AND U4214 ( .A(p_input[6208]), .B(p_input[16208]), .Z(o[6208]) );
  AND U4215 ( .A(p_input[6207]), .B(p_input[16207]), .Z(o[6207]) );
  AND U4216 ( .A(p_input[6206]), .B(p_input[16206]), .Z(o[6206]) );
  AND U4217 ( .A(p_input[6205]), .B(p_input[16205]), .Z(o[6205]) );
  AND U4218 ( .A(p_input[6204]), .B(p_input[16204]), .Z(o[6204]) );
  AND U4219 ( .A(p_input[6203]), .B(p_input[16203]), .Z(o[6203]) );
  AND U4220 ( .A(p_input[6202]), .B(p_input[16202]), .Z(o[6202]) );
  AND U4221 ( .A(p_input[6201]), .B(p_input[16201]), .Z(o[6201]) );
  AND U4222 ( .A(p_input[6200]), .B(p_input[16200]), .Z(o[6200]) );
  AND U4223 ( .A(p_input[61]), .B(p_input[10061]), .Z(o[61]) );
  AND U4224 ( .A(p_input[619]), .B(p_input[10619]), .Z(o[619]) );
  AND U4225 ( .A(p_input[6199]), .B(p_input[16199]), .Z(o[6199]) );
  AND U4226 ( .A(p_input[6198]), .B(p_input[16198]), .Z(o[6198]) );
  AND U4227 ( .A(p_input[6197]), .B(p_input[16197]), .Z(o[6197]) );
  AND U4228 ( .A(p_input[6196]), .B(p_input[16196]), .Z(o[6196]) );
  AND U4229 ( .A(p_input[6195]), .B(p_input[16195]), .Z(o[6195]) );
  AND U4230 ( .A(p_input[6194]), .B(p_input[16194]), .Z(o[6194]) );
  AND U4231 ( .A(p_input[6193]), .B(p_input[16193]), .Z(o[6193]) );
  AND U4232 ( .A(p_input[6192]), .B(p_input[16192]), .Z(o[6192]) );
  AND U4233 ( .A(p_input[6191]), .B(p_input[16191]), .Z(o[6191]) );
  AND U4234 ( .A(p_input[6190]), .B(p_input[16190]), .Z(o[6190]) );
  AND U4235 ( .A(p_input[618]), .B(p_input[10618]), .Z(o[618]) );
  AND U4236 ( .A(p_input[6189]), .B(p_input[16189]), .Z(o[6189]) );
  AND U4237 ( .A(p_input[6188]), .B(p_input[16188]), .Z(o[6188]) );
  AND U4238 ( .A(p_input[6187]), .B(p_input[16187]), .Z(o[6187]) );
  AND U4239 ( .A(p_input[6186]), .B(p_input[16186]), .Z(o[6186]) );
  AND U4240 ( .A(p_input[6185]), .B(p_input[16185]), .Z(o[6185]) );
  AND U4241 ( .A(p_input[6184]), .B(p_input[16184]), .Z(o[6184]) );
  AND U4242 ( .A(p_input[6183]), .B(p_input[16183]), .Z(o[6183]) );
  AND U4243 ( .A(p_input[6182]), .B(p_input[16182]), .Z(o[6182]) );
  AND U4244 ( .A(p_input[6181]), .B(p_input[16181]), .Z(o[6181]) );
  AND U4245 ( .A(p_input[6180]), .B(p_input[16180]), .Z(o[6180]) );
  AND U4246 ( .A(p_input[617]), .B(p_input[10617]), .Z(o[617]) );
  AND U4247 ( .A(p_input[6179]), .B(p_input[16179]), .Z(o[6179]) );
  AND U4248 ( .A(p_input[6178]), .B(p_input[16178]), .Z(o[6178]) );
  AND U4249 ( .A(p_input[6177]), .B(p_input[16177]), .Z(o[6177]) );
  AND U4250 ( .A(p_input[6176]), .B(p_input[16176]), .Z(o[6176]) );
  AND U4251 ( .A(p_input[6175]), .B(p_input[16175]), .Z(o[6175]) );
  AND U4252 ( .A(p_input[6174]), .B(p_input[16174]), .Z(o[6174]) );
  AND U4253 ( .A(p_input[6173]), .B(p_input[16173]), .Z(o[6173]) );
  AND U4254 ( .A(p_input[6172]), .B(p_input[16172]), .Z(o[6172]) );
  AND U4255 ( .A(p_input[6171]), .B(p_input[16171]), .Z(o[6171]) );
  AND U4256 ( .A(p_input[6170]), .B(p_input[16170]), .Z(o[6170]) );
  AND U4257 ( .A(p_input[616]), .B(p_input[10616]), .Z(o[616]) );
  AND U4258 ( .A(p_input[6169]), .B(p_input[16169]), .Z(o[6169]) );
  AND U4259 ( .A(p_input[6168]), .B(p_input[16168]), .Z(o[6168]) );
  AND U4260 ( .A(p_input[6167]), .B(p_input[16167]), .Z(o[6167]) );
  AND U4261 ( .A(p_input[6166]), .B(p_input[16166]), .Z(o[6166]) );
  AND U4262 ( .A(p_input[6165]), .B(p_input[16165]), .Z(o[6165]) );
  AND U4263 ( .A(p_input[6164]), .B(p_input[16164]), .Z(o[6164]) );
  AND U4264 ( .A(p_input[6163]), .B(p_input[16163]), .Z(o[6163]) );
  AND U4265 ( .A(p_input[6162]), .B(p_input[16162]), .Z(o[6162]) );
  AND U4266 ( .A(p_input[6161]), .B(p_input[16161]), .Z(o[6161]) );
  AND U4267 ( .A(p_input[6160]), .B(p_input[16160]), .Z(o[6160]) );
  AND U4268 ( .A(p_input[615]), .B(p_input[10615]), .Z(o[615]) );
  AND U4269 ( .A(p_input[6159]), .B(p_input[16159]), .Z(o[6159]) );
  AND U4270 ( .A(p_input[6158]), .B(p_input[16158]), .Z(o[6158]) );
  AND U4271 ( .A(p_input[6157]), .B(p_input[16157]), .Z(o[6157]) );
  AND U4272 ( .A(p_input[6156]), .B(p_input[16156]), .Z(o[6156]) );
  AND U4273 ( .A(p_input[6155]), .B(p_input[16155]), .Z(o[6155]) );
  AND U4274 ( .A(p_input[6154]), .B(p_input[16154]), .Z(o[6154]) );
  AND U4275 ( .A(p_input[6153]), .B(p_input[16153]), .Z(o[6153]) );
  AND U4276 ( .A(p_input[6152]), .B(p_input[16152]), .Z(o[6152]) );
  AND U4277 ( .A(p_input[6151]), .B(p_input[16151]), .Z(o[6151]) );
  AND U4278 ( .A(p_input[6150]), .B(p_input[16150]), .Z(o[6150]) );
  AND U4279 ( .A(p_input[614]), .B(p_input[10614]), .Z(o[614]) );
  AND U4280 ( .A(p_input[6149]), .B(p_input[16149]), .Z(o[6149]) );
  AND U4281 ( .A(p_input[6148]), .B(p_input[16148]), .Z(o[6148]) );
  AND U4282 ( .A(p_input[6147]), .B(p_input[16147]), .Z(o[6147]) );
  AND U4283 ( .A(p_input[6146]), .B(p_input[16146]), .Z(o[6146]) );
  AND U4284 ( .A(p_input[6145]), .B(p_input[16145]), .Z(o[6145]) );
  AND U4285 ( .A(p_input[6144]), .B(p_input[16144]), .Z(o[6144]) );
  AND U4286 ( .A(p_input[6143]), .B(p_input[16143]), .Z(o[6143]) );
  AND U4287 ( .A(p_input[6142]), .B(p_input[16142]), .Z(o[6142]) );
  AND U4288 ( .A(p_input[6141]), .B(p_input[16141]), .Z(o[6141]) );
  AND U4289 ( .A(p_input[6140]), .B(p_input[16140]), .Z(o[6140]) );
  AND U4290 ( .A(p_input[613]), .B(p_input[10613]), .Z(o[613]) );
  AND U4291 ( .A(p_input[6139]), .B(p_input[16139]), .Z(o[6139]) );
  AND U4292 ( .A(p_input[6138]), .B(p_input[16138]), .Z(o[6138]) );
  AND U4293 ( .A(p_input[6137]), .B(p_input[16137]), .Z(o[6137]) );
  AND U4294 ( .A(p_input[6136]), .B(p_input[16136]), .Z(o[6136]) );
  AND U4295 ( .A(p_input[6135]), .B(p_input[16135]), .Z(o[6135]) );
  AND U4296 ( .A(p_input[6134]), .B(p_input[16134]), .Z(o[6134]) );
  AND U4297 ( .A(p_input[6133]), .B(p_input[16133]), .Z(o[6133]) );
  AND U4298 ( .A(p_input[6132]), .B(p_input[16132]), .Z(o[6132]) );
  AND U4299 ( .A(p_input[6131]), .B(p_input[16131]), .Z(o[6131]) );
  AND U4300 ( .A(p_input[6130]), .B(p_input[16130]), .Z(o[6130]) );
  AND U4301 ( .A(p_input[612]), .B(p_input[10612]), .Z(o[612]) );
  AND U4302 ( .A(p_input[6129]), .B(p_input[16129]), .Z(o[6129]) );
  AND U4303 ( .A(p_input[6128]), .B(p_input[16128]), .Z(o[6128]) );
  AND U4304 ( .A(p_input[6127]), .B(p_input[16127]), .Z(o[6127]) );
  AND U4305 ( .A(p_input[6126]), .B(p_input[16126]), .Z(o[6126]) );
  AND U4306 ( .A(p_input[6125]), .B(p_input[16125]), .Z(o[6125]) );
  AND U4307 ( .A(p_input[6124]), .B(p_input[16124]), .Z(o[6124]) );
  AND U4308 ( .A(p_input[6123]), .B(p_input[16123]), .Z(o[6123]) );
  AND U4309 ( .A(p_input[6122]), .B(p_input[16122]), .Z(o[6122]) );
  AND U4310 ( .A(p_input[6121]), .B(p_input[16121]), .Z(o[6121]) );
  AND U4311 ( .A(p_input[6120]), .B(p_input[16120]), .Z(o[6120]) );
  AND U4312 ( .A(p_input[611]), .B(p_input[10611]), .Z(o[611]) );
  AND U4313 ( .A(p_input[6119]), .B(p_input[16119]), .Z(o[6119]) );
  AND U4314 ( .A(p_input[6118]), .B(p_input[16118]), .Z(o[6118]) );
  AND U4315 ( .A(p_input[6117]), .B(p_input[16117]), .Z(o[6117]) );
  AND U4316 ( .A(p_input[6116]), .B(p_input[16116]), .Z(o[6116]) );
  AND U4317 ( .A(p_input[6115]), .B(p_input[16115]), .Z(o[6115]) );
  AND U4318 ( .A(p_input[6114]), .B(p_input[16114]), .Z(o[6114]) );
  AND U4319 ( .A(p_input[6113]), .B(p_input[16113]), .Z(o[6113]) );
  AND U4320 ( .A(p_input[6112]), .B(p_input[16112]), .Z(o[6112]) );
  AND U4321 ( .A(p_input[6111]), .B(p_input[16111]), .Z(o[6111]) );
  AND U4322 ( .A(p_input[6110]), .B(p_input[16110]), .Z(o[6110]) );
  AND U4323 ( .A(p_input[610]), .B(p_input[10610]), .Z(o[610]) );
  AND U4324 ( .A(p_input[6109]), .B(p_input[16109]), .Z(o[6109]) );
  AND U4325 ( .A(p_input[6108]), .B(p_input[16108]), .Z(o[6108]) );
  AND U4326 ( .A(p_input[6107]), .B(p_input[16107]), .Z(o[6107]) );
  AND U4327 ( .A(p_input[6106]), .B(p_input[16106]), .Z(o[6106]) );
  AND U4328 ( .A(p_input[6105]), .B(p_input[16105]), .Z(o[6105]) );
  AND U4329 ( .A(p_input[6104]), .B(p_input[16104]), .Z(o[6104]) );
  AND U4330 ( .A(p_input[6103]), .B(p_input[16103]), .Z(o[6103]) );
  AND U4331 ( .A(p_input[6102]), .B(p_input[16102]), .Z(o[6102]) );
  AND U4332 ( .A(p_input[6101]), .B(p_input[16101]), .Z(o[6101]) );
  AND U4333 ( .A(p_input[6100]), .B(p_input[16100]), .Z(o[6100]) );
  AND U4334 ( .A(p_input[60]), .B(p_input[10060]), .Z(o[60]) );
  AND U4335 ( .A(p_input[609]), .B(p_input[10609]), .Z(o[609]) );
  AND U4336 ( .A(p_input[6099]), .B(p_input[16099]), .Z(o[6099]) );
  AND U4337 ( .A(p_input[6098]), .B(p_input[16098]), .Z(o[6098]) );
  AND U4338 ( .A(p_input[6097]), .B(p_input[16097]), .Z(o[6097]) );
  AND U4339 ( .A(p_input[6096]), .B(p_input[16096]), .Z(o[6096]) );
  AND U4340 ( .A(p_input[6095]), .B(p_input[16095]), .Z(o[6095]) );
  AND U4341 ( .A(p_input[6094]), .B(p_input[16094]), .Z(o[6094]) );
  AND U4342 ( .A(p_input[6093]), .B(p_input[16093]), .Z(o[6093]) );
  AND U4343 ( .A(p_input[6092]), .B(p_input[16092]), .Z(o[6092]) );
  AND U4344 ( .A(p_input[6091]), .B(p_input[16091]), .Z(o[6091]) );
  AND U4345 ( .A(p_input[6090]), .B(p_input[16090]), .Z(o[6090]) );
  AND U4346 ( .A(p_input[608]), .B(p_input[10608]), .Z(o[608]) );
  AND U4347 ( .A(p_input[6089]), .B(p_input[16089]), .Z(o[6089]) );
  AND U4348 ( .A(p_input[6088]), .B(p_input[16088]), .Z(o[6088]) );
  AND U4349 ( .A(p_input[6087]), .B(p_input[16087]), .Z(o[6087]) );
  AND U4350 ( .A(p_input[6086]), .B(p_input[16086]), .Z(o[6086]) );
  AND U4351 ( .A(p_input[6085]), .B(p_input[16085]), .Z(o[6085]) );
  AND U4352 ( .A(p_input[6084]), .B(p_input[16084]), .Z(o[6084]) );
  AND U4353 ( .A(p_input[6083]), .B(p_input[16083]), .Z(o[6083]) );
  AND U4354 ( .A(p_input[6082]), .B(p_input[16082]), .Z(o[6082]) );
  AND U4355 ( .A(p_input[6081]), .B(p_input[16081]), .Z(o[6081]) );
  AND U4356 ( .A(p_input[6080]), .B(p_input[16080]), .Z(o[6080]) );
  AND U4357 ( .A(p_input[607]), .B(p_input[10607]), .Z(o[607]) );
  AND U4358 ( .A(p_input[6079]), .B(p_input[16079]), .Z(o[6079]) );
  AND U4359 ( .A(p_input[6078]), .B(p_input[16078]), .Z(o[6078]) );
  AND U4360 ( .A(p_input[6077]), .B(p_input[16077]), .Z(o[6077]) );
  AND U4361 ( .A(p_input[6076]), .B(p_input[16076]), .Z(o[6076]) );
  AND U4362 ( .A(p_input[6075]), .B(p_input[16075]), .Z(o[6075]) );
  AND U4363 ( .A(p_input[6074]), .B(p_input[16074]), .Z(o[6074]) );
  AND U4364 ( .A(p_input[6073]), .B(p_input[16073]), .Z(o[6073]) );
  AND U4365 ( .A(p_input[6072]), .B(p_input[16072]), .Z(o[6072]) );
  AND U4366 ( .A(p_input[6071]), .B(p_input[16071]), .Z(o[6071]) );
  AND U4367 ( .A(p_input[6070]), .B(p_input[16070]), .Z(o[6070]) );
  AND U4368 ( .A(p_input[606]), .B(p_input[10606]), .Z(o[606]) );
  AND U4369 ( .A(p_input[6069]), .B(p_input[16069]), .Z(o[6069]) );
  AND U4370 ( .A(p_input[6068]), .B(p_input[16068]), .Z(o[6068]) );
  AND U4371 ( .A(p_input[6067]), .B(p_input[16067]), .Z(o[6067]) );
  AND U4372 ( .A(p_input[6066]), .B(p_input[16066]), .Z(o[6066]) );
  AND U4373 ( .A(p_input[6065]), .B(p_input[16065]), .Z(o[6065]) );
  AND U4374 ( .A(p_input[6064]), .B(p_input[16064]), .Z(o[6064]) );
  AND U4375 ( .A(p_input[6063]), .B(p_input[16063]), .Z(o[6063]) );
  AND U4376 ( .A(p_input[6062]), .B(p_input[16062]), .Z(o[6062]) );
  AND U4377 ( .A(p_input[6061]), .B(p_input[16061]), .Z(o[6061]) );
  AND U4378 ( .A(p_input[6060]), .B(p_input[16060]), .Z(o[6060]) );
  AND U4379 ( .A(p_input[605]), .B(p_input[10605]), .Z(o[605]) );
  AND U4380 ( .A(p_input[6059]), .B(p_input[16059]), .Z(o[6059]) );
  AND U4381 ( .A(p_input[6058]), .B(p_input[16058]), .Z(o[6058]) );
  AND U4382 ( .A(p_input[6057]), .B(p_input[16057]), .Z(o[6057]) );
  AND U4383 ( .A(p_input[6056]), .B(p_input[16056]), .Z(o[6056]) );
  AND U4384 ( .A(p_input[6055]), .B(p_input[16055]), .Z(o[6055]) );
  AND U4385 ( .A(p_input[6054]), .B(p_input[16054]), .Z(o[6054]) );
  AND U4386 ( .A(p_input[6053]), .B(p_input[16053]), .Z(o[6053]) );
  AND U4387 ( .A(p_input[6052]), .B(p_input[16052]), .Z(o[6052]) );
  AND U4388 ( .A(p_input[6051]), .B(p_input[16051]), .Z(o[6051]) );
  AND U4389 ( .A(p_input[6050]), .B(p_input[16050]), .Z(o[6050]) );
  AND U4390 ( .A(p_input[604]), .B(p_input[10604]), .Z(o[604]) );
  AND U4391 ( .A(p_input[6049]), .B(p_input[16049]), .Z(o[6049]) );
  AND U4392 ( .A(p_input[6048]), .B(p_input[16048]), .Z(o[6048]) );
  AND U4393 ( .A(p_input[6047]), .B(p_input[16047]), .Z(o[6047]) );
  AND U4394 ( .A(p_input[6046]), .B(p_input[16046]), .Z(o[6046]) );
  AND U4395 ( .A(p_input[6045]), .B(p_input[16045]), .Z(o[6045]) );
  AND U4396 ( .A(p_input[6044]), .B(p_input[16044]), .Z(o[6044]) );
  AND U4397 ( .A(p_input[6043]), .B(p_input[16043]), .Z(o[6043]) );
  AND U4398 ( .A(p_input[6042]), .B(p_input[16042]), .Z(o[6042]) );
  AND U4399 ( .A(p_input[6041]), .B(p_input[16041]), .Z(o[6041]) );
  AND U4400 ( .A(p_input[6040]), .B(p_input[16040]), .Z(o[6040]) );
  AND U4401 ( .A(p_input[603]), .B(p_input[10603]), .Z(o[603]) );
  AND U4402 ( .A(p_input[6039]), .B(p_input[16039]), .Z(o[6039]) );
  AND U4403 ( .A(p_input[6038]), .B(p_input[16038]), .Z(o[6038]) );
  AND U4404 ( .A(p_input[6037]), .B(p_input[16037]), .Z(o[6037]) );
  AND U4405 ( .A(p_input[6036]), .B(p_input[16036]), .Z(o[6036]) );
  AND U4406 ( .A(p_input[6035]), .B(p_input[16035]), .Z(o[6035]) );
  AND U4407 ( .A(p_input[6034]), .B(p_input[16034]), .Z(o[6034]) );
  AND U4408 ( .A(p_input[6033]), .B(p_input[16033]), .Z(o[6033]) );
  AND U4409 ( .A(p_input[6032]), .B(p_input[16032]), .Z(o[6032]) );
  AND U4410 ( .A(p_input[6031]), .B(p_input[16031]), .Z(o[6031]) );
  AND U4411 ( .A(p_input[6030]), .B(p_input[16030]), .Z(o[6030]) );
  AND U4412 ( .A(p_input[602]), .B(p_input[10602]), .Z(o[602]) );
  AND U4413 ( .A(p_input[6029]), .B(p_input[16029]), .Z(o[6029]) );
  AND U4414 ( .A(p_input[6028]), .B(p_input[16028]), .Z(o[6028]) );
  AND U4415 ( .A(p_input[6027]), .B(p_input[16027]), .Z(o[6027]) );
  AND U4416 ( .A(p_input[6026]), .B(p_input[16026]), .Z(o[6026]) );
  AND U4417 ( .A(p_input[6025]), .B(p_input[16025]), .Z(o[6025]) );
  AND U4418 ( .A(p_input[6024]), .B(p_input[16024]), .Z(o[6024]) );
  AND U4419 ( .A(p_input[6023]), .B(p_input[16023]), .Z(o[6023]) );
  AND U4420 ( .A(p_input[6022]), .B(p_input[16022]), .Z(o[6022]) );
  AND U4421 ( .A(p_input[6021]), .B(p_input[16021]), .Z(o[6021]) );
  AND U4422 ( .A(p_input[6020]), .B(p_input[16020]), .Z(o[6020]) );
  AND U4423 ( .A(p_input[601]), .B(p_input[10601]), .Z(o[601]) );
  AND U4424 ( .A(p_input[6019]), .B(p_input[16019]), .Z(o[6019]) );
  AND U4425 ( .A(p_input[6018]), .B(p_input[16018]), .Z(o[6018]) );
  AND U4426 ( .A(p_input[6017]), .B(p_input[16017]), .Z(o[6017]) );
  AND U4427 ( .A(p_input[6016]), .B(p_input[16016]), .Z(o[6016]) );
  AND U4428 ( .A(p_input[6015]), .B(p_input[16015]), .Z(o[6015]) );
  AND U4429 ( .A(p_input[6014]), .B(p_input[16014]), .Z(o[6014]) );
  AND U4430 ( .A(p_input[6013]), .B(p_input[16013]), .Z(o[6013]) );
  AND U4431 ( .A(p_input[6012]), .B(p_input[16012]), .Z(o[6012]) );
  AND U4432 ( .A(p_input[6011]), .B(p_input[16011]), .Z(o[6011]) );
  AND U4433 ( .A(p_input[6010]), .B(p_input[16010]), .Z(o[6010]) );
  AND U4434 ( .A(p_input[600]), .B(p_input[10600]), .Z(o[600]) );
  AND U4435 ( .A(p_input[6009]), .B(p_input[16009]), .Z(o[6009]) );
  AND U4436 ( .A(p_input[6008]), .B(p_input[16008]), .Z(o[6008]) );
  AND U4437 ( .A(p_input[6007]), .B(p_input[16007]), .Z(o[6007]) );
  AND U4438 ( .A(p_input[6006]), .B(p_input[16006]), .Z(o[6006]) );
  AND U4439 ( .A(p_input[6005]), .B(p_input[16005]), .Z(o[6005]) );
  AND U4440 ( .A(p_input[6004]), .B(p_input[16004]), .Z(o[6004]) );
  AND U4441 ( .A(p_input[6003]), .B(p_input[16003]), .Z(o[6003]) );
  AND U4442 ( .A(p_input[6002]), .B(p_input[16002]), .Z(o[6002]) );
  AND U4443 ( .A(p_input[6001]), .B(p_input[16001]), .Z(o[6001]) );
  AND U4444 ( .A(p_input[6000]), .B(p_input[16000]), .Z(o[6000]) );
  AND U4445 ( .A(p_input[5]), .B(p_input[10005]), .Z(o[5]) );
  AND U4446 ( .A(p_input[59]), .B(p_input[10059]), .Z(o[59]) );
  AND U4447 ( .A(p_input[599]), .B(p_input[10599]), .Z(o[599]) );
  AND U4448 ( .A(p_input[5999]), .B(p_input[15999]), .Z(o[5999]) );
  AND U4449 ( .A(p_input[5998]), .B(p_input[15998]), .Z(o[5998]) );
  AND U4450 ( .A(p_input[5997]), .B(p_input[15997]), .Z(o[5997]) );
  AND U4451 ( .A(p_input[5996]), .B(p_input[15996]), .Z(o[5996]) );
  AND U4452 ( .A(p_input[5995]), .B(p_input[15995]), .Z(o[5995]) );
  AND U4453 ( .A(p_input[5994]), .B(p_input[15994]), .Z(o[5994]) );
  AND U4454 ( .A(p_input[5993]), .B(p_input[15993]), .Z(o[5993]) );
  AND U4455 ( .A(p_input[5992]), .B(p_input[15992]), .Z(o[5992]) );
  AND U4456 ( .A(p_input[5991]), .B(p_input[15991]), .Z(o[5991]) );
  AND U4457 ( .A(p_input[5990]), .B(p_input[15990]), .Z(o[5990]) );
  AND U4458 ( .A(p_input[598]), .B(p_input[10598]), .Z(o[598]) );
  AND U4459 ( .A(p_input[5989]), .B(p_input[15989]), .Z(o[5989]) );
  AND U4460 ( .A(p_input[5988]), .B(p_input[15988]), .Z(o[5988]) );
  AND U4461 ( .A(p_input[5987]), .B(p_input[15987]), .Z(o[5987]) );
  AND U4462 ( .A(p_input[5986]), .B(p_input[15986]), .Z(o[5986]) );
  AND U4463 ( .A(p_input[5985]), .B(p_input[15985]), .Z(o[5985]) );
  AND U4464 ( .A(p_input[5984]), .B(p_input[15984]), .Z(o[5984]) );
  AND U4465 ( .A(p_input[5983]), .B(p_input[15983]), .Z(o[5983]) );
  AND U4466 ( .A(p_input[5982]), .B(p_input[15982]), .Z(o[5982]) );
  AND U4467 ( .A(p_input[5981]), .B(p_input[15981]), .Z(o[5981]) );
  AND U4468 ( .A(p_input[5980]), .B(p_input[15980]), .Z(o[5980]) );
  AND U4469 ( .A(p_input[597]), .B(p_input[10597]), .Z(o[597]) );
  AND U4470 ( .A(p_input[5979]), .B(p_input[15979]), .Z(o[5979]) );
  AND U4471 ( .A(p_input[5978]), .B(p_input[15978]), .Z(o[5978]) );
  AND U4472 ( .A(p_input[5977]), .B(p_input[15977]), .Z(o[5977]) );
  AND U4473 ( .A(p_input[5976]), .B(p_input[15976]), .Z(o[5976]) );
  AND U4474 ( .A(p_input[5975]), .B(p_input[15975]), .Z(o[5975]) );
  AND U4475 ( .A(p_input[5974]), .B(p_input[15974]), .Z(o[5974]) );
  AND U4476 ( .A(p_input[5973]), .B(p_input[15973]), .Z(o[5973]) );
  AND U4477 ( .A(p_input[5972]), .B(p_input[15972]), .Z(o[5972]) );
  AND U4478 ( .A(p_input[5971]), .B(p_input[15971]), .Z(o[5971]) );
  AND U4479 ( .A(p_input[5970]), .B(p_input[15970]), .Z(o[5970]) );
  AND U4480 ( .A(p_input[596]), .B(p_input[10596]), .Z(o[596]) );
  AND U4481 ( .A(p_input[5969]), .B(p_input[15969]), .Z(o[5969]) );
  AND U4482 ( .A(p_input[5968]), .B(p_input[15968]), .Z(o[5968]) );
  AND U4483 ( .A(p_input[5967]), .B(p_input[15967]), .Z(o[5967]) );
  AND U4484 ( .A(p_input[5966]), .B(p_input[15966]), .Z(o[5966]) );
  AND U4485 ( .A(p_input[5965]), .B(p_input[15965]), .Z(o[5965]) );
  AND U4486 ( .A(p_input[5964]), .B(p_input[15964]), .Z(o[5964]) );
  AND U4487 ( .A(p_input[5963]), .B(p_input[15963]), .Z(o[5963]) );
  AND U4488 ( .A(p_input[5962]), .B(p_input[15962]), .Z(o[5962]) );
  AND U4489 ( .A(p_input[5961]), .B(p_input[15961]), .Z(o[5961]) );
  AND U4490 ( .A(p_input[5960]), .B(p_input[15960]), .Z(o[5960]) );
  AND U4491 ( .A(p_input[595]), .B(p_input[10595]), .Z(o[595]) );
  AND U4492 ( .A(p_input[5959]), .B(p_input[15959]), .Z(o[5959]) );
  AND U4493 ( .A(p_input[5958]), .B(p_input[15958]), .Z(o[5958]) );
  AND U4494 ( .A(p_input[5957]), .B(p_input[15957]), .Z(o[5957]) );
  AND U4495 ( .A(p_input[5956]), .B(p_input[15956]), .Z(o[5956]) );
  AND U4496 ( .A(p_input[5955]), .B(p_input[15955]), .Z(o[5955]) );
  AND U4497 ( .A(p_input[5954]), .B(p_input[15954]), .Z(o[5954]) );
  AND U4498 ( .A(p_input[5953]), .B(p_input[15953]), .Z(o[5953]) );
  AND U4499 ( .A(p_input[5952]), .B(p_input[15952]), .Z(o[5952]) );
  AND U4500 ( .A(p_input[5951]), .B(p_input[15951]), .Z(o[5951]) );
  AND U4501 ( .A(p_input[5950]), .B(p_input[15950]), .Z(o[5950]) );
  AND U4502 ( .A(p_input[594]), .B(p_input[10594]), .Z(o[594]) );
  AND U4503 ( .A(p_input[5949]), .B(p_input[15949]), .Z(o[5949]) );
  AND U4504 ( .A(p_input[5948]), .B(p_input[15948]), .Z(o[5948]) );
  AND U4505 ( .A(p_input[5947]), .B(p_input[15947]), .Z(o[5947]) );
  AND U4506 ( .A(p_input[5946]), .B(p_input[15946]), .Z(o[5946]) );
  AND U4507 ( .A(p_input[5945]), .B(p_input[15945]), .Z(o[5945]) );
  AND U4508 ( .A(p_input[5944]), .B(p_input[15944]), .Z(o[5944]) );
  AND U4509 ( .A(p_input[5943]), .B(p_input[15943]), .Z(o[5943]) );
  AND U4510 ( .A(p_input[5942]), .B(p_input[15942]), .Z(o[5942]) );
  AND U4511 ( .A(p_input[5941]), .B(p_input[15941]), .Z(o[5941]) );
  AND U4512 ( .A(p_input[5940]), .B(p_input[15940]), .Z(o[5940]) );
  AND U4513 ( .A(p_input[593]), .B(p_input[10593]), .Z(o[593]) );
  AND U4514 ( .A(p_input[5939]), .B(p_input[15939]), .Z(o[5939]) );
  AND U4515 ( .A(p_input[5938]), .B(p_input[15938]), .Z(o[5938]) );
  AND U4516 ( .A(p_input[5937]), .B(p_input[15937]), .Z(o[5937]) );
  AND U4517 ( .A(p_input[5936]), .B(p_input[15936]), .Z(o[5936]) );
  AND U4518 ( .A(p_input[5935]), .B(p_input[15935]), .Z(o[5935]) );
  AND U4519 ( .A(p_input[5934]), .B(p_input[15934]), .Z(o[5934]) );
  AND U4520 ( .A(p_input[5933]), .B(p_input[15933]), .Z(o[5933]) );
  AND U4521 ( .A(p_input[5932]), .B(p_input[15932]), .Z(o[5932]) );
  AND U4522 ( .A(p_input[5931]), .B(p_input[15931]), .Z(o[5931]) );
  AND U4523 ( .A(p_input[5930]), .B(p_input[15930]), .Z(o[5930]) );
  AND U4524 ( .A(p_input[592]), .B(p_input[10592]), .Z(o[592]) );
  AND U4525 ( .A(p_input[5929]), .B(p_input[15929]), .Z(o[5929]) );
  AND U4526 ( .A(p_input[5928]), .B(p_input[15928]), .Z(o[5928]) );
  AND U4527 ( .A(p_input[5927]), .B(p_input[15927]), .Z(o[5927]) );
  AND U4528 ( .A(p_input[5926]), .B(p_input[15926]), .Z(o[5926]) );
  AND U4529 ( .A(p_input[5925]), .B(p_input[15925]), .Z(o[5925]) );
  AND U4530 ( .A(p_input[5924]), .B(p_input[15924]), .Z(o[5924]) );
  AND U4531 ( .A(p_input[5923]), .B(p_input[15923]), .Z(o[5923]) );
  AND U4532 ( .A(p_input[5922]), .B(p_input[15922]), .Z(o[5922]) );
  AND U4533 ( .A(p_input[5921]), .B(p_input[15921]), .Z(o[5921]) );
  AND U4534 ( .A(p_input[5920]), .B(p_input[15920]), .Z(o[5920]) );
  AND U4535 ( .A(p_input[591]), .B(p_input[10591]), .Z(o[591]) );
  AND U4536 ( .A(p_input[5919]), .B(p_input[15919]), .Z(o[5919]) );
  AND U4537 ( .A(p_input[5918]), .B(p_input[15918]), .Z(o[5918]) );
  AND U4538 ( .A(p_input[5917]), .B(p_input[15917]), .Z(o[5917]) );
  AND U4539 ( .A(p_input[5916]), .B(p_input[15916]), .Z(o[5916]) );
  AND U4540 ( .A(p_input[5915]), .B(p_input[15915]), .Z(o[5915]) );
  AND U4541 ( .A(p_input[5914]), .B(p_input[15914]), .Z(o[5914]) );
  AND U4542 ( .A(p_input[5913]), .B(p_input[15913]), .Z(o[5913]) );
  AND U4543 ( .A(p_input[5912]), .B(p_input[15912]), .Z(o[5912]) );
  AND U4544 ( .A(p_input[5911]), .B(p_input[15911]), .Z(o[5911]) );
  AND U4545 ( .A(p_input[5910]), .B(p_input[15910]), .Z(o[5910]) );
  AND U4546 ( .A(p_input[590]), .B(p_input[10590]), .Z(o[590]) );
  AND U4547 ( .A(p_input[5909]), .B(p_input[15909]), .Z(o[5909]) );
  AND U4548 ( .A(p_input[5908]), .B(p_input[15908]), .Z(o[5908]) );
  AND U4549 ( .A(p_input[5907]), .B(p_input[15907]), .Z(o[5907]) );
  AND U4550 ( .A(p_input[5906]), .B(p_input[15906]), .Z(o[5906]) );
  AND U4551 ( .A(p_input[5905]), .B(p_input[15905]), .Z(o[5905]) );
  AND U4552 ( .A(p_input[5904]), .B(p_input[15904]), .Z(o[5904]) );
  AND U4553 ( .A(p_input[5903]), .B(p_input[15903]), .Z(o[5903]) );
  AND U4554 ( .A(p_input[5902]), .B(p_input[15902]), .Z(o[5902]) );
  AND U4555 ( .A(p_input[5901]), .B(p_input[15901]), .Z(o[5901]) );
  AND U4556 ( .A(p_input[5900]), .B(p_input[15900]), .Z(o[5900]) );
  AND U4557 ( .A(p_input[58]), .B(p_input[10058]), .Z(o[58]) );
  AND U4558 ( .A(p_input[589]), .B(p_input[10589]), .Z(o[589]) );
  AND U4559 ( .A(p_input[5899]), .B(p_input[15899]), .Z(o[5899]) );
  AND U4560 ( .A(p_input[5898]), .B(p_input[15898]), .Z(o[5898]) );
  AND U4561 ( .A(p_input[5897]), .B(p_input[15897]), .Z(o[5897]) );
  AND U4562 ( .A(p_input[5896]), .B(p_input[15896]), .Z(o[5896]) );
  AND U4563 ( .A(p_input[5895]), .B(p_input[15895]), .Z(o[5895]) );
  AND U4564 ( .A(p_input[5894]), .B(p_input[15894]), .Z(o[5894]) );
  AND U4565 ( .A(p_input[5893]), .B(p_input[15893]), .Z(o[5893]) );
  AND U4566 ( .A(p_input[5892]), .B(p_input[15892]), .Z(o[5892]) );
  AND U4567 ( .A(p_input[5891]), .B(p_input[15891]), .Z(o[5891]) );
  AND U4568 ( .A(p_input[5890]), .B(p_input[15890]), .Z(o[5890]) );
  AND U4569 ( .A(p_input[588]), .B(p_input[10588]), .Z(o[588]) );
  AND U4570 ( .A(p_input[5889]), .B(p_input[15889]), .Z(o[5889]) );
  AND U4571 ( .A(p_input[5888]), .B(p_input[15888]), .Z(o[5888]) );
  AND U4572 ( .A(p_input[5887]), .B(p_input[15887]), .Z(o[5887]) );
  AND U4573 ( .A(p_input[5886]), .B(p_input[15886]), .Z(o[5886]) );
  AND U4574 ( .A(p_input[5885]), .B(p_input[15885]), .Z(o[5885]) );
  AND U4575 ( .A(p_input[5884]), .B(p_input[15884]), .Z(o[5884]) );
  AND U4576 ( .A(p_input[5883]), .B(p_input[15883]), .Z(o[5883]) );
  AND U4577 ( .A(p_input[5882]), .B(p_input[15882]), .Z(o[5882]) );
  AND U4578 ( .A(p_input[5881]), .B(p_input[15881]), .Z(o[5881]) );
  AND U4579 ( .A(p_input[5880]), .B(p_input[15880]), .Z(o[5880]) );
  AND U4580 ( .A(p_input[587]), .B(p_input[10587]), .Z(o[587]) );
  AND U4581 ( .A(p_input[5879]), .B(p_input[15879]), .Z(o[5879]) );
  AND U4582 ( .A(p_input[5878]), .B(p_input[15878]), .Z(o[5878]) );
  AND U4583 ( .A(p_input[5877]), .B(p_input[15877]), .Z(o[5877]) );
  AND U4584 ( .A(p_input[5876]), .B(p_input[15876]), .Z(o[5876]) );
  AND U4585 ( .A(p_input[5875]), .B(p_input[15875]), .Z(o[5875]) );
  AND U4586 ( .A(p_input[5874]), .B(p_input[15874]), .Z(o[5874]) );
  AND U4587 ( .A(p_input[5873]), .B(p_input[15873]), .Z(o[5873]) );
  AND U4588 ( .A(p_input[5872]), .B(p_input[15872]), .Z(o[5872]) );
  AND U4589 ( .A(p_input[5871]), .B(p_input[15871]), .Z(o[5871]) );
  AND U4590 ( .A(p_input[5870]), .B(p_input[15870]), .Z(o[5870]) );
  AND U4591 ( .A(p_input[586]), .B(p_input[10586]), .Z(o[586]) );
  AND U4592 ( .A(p_input[5869]), .B(p_input[15869]), .Z(o[5869]) );
  AND U4593 ( .A(p_input[5868]), .B(p_input[15868]), .Z(o[5868]) );
  AND U4594 ( .A(p_input[5867]), .B(p_input[15867]), .Z(o[5867]) );
  AND U4595 ( .A(p_input[5866]), .B(p_input[15866]), .Z(o[5866]) );
  AND U4596 ( .A(p_input[5865]), .B(p_input[15865]), .Z(o[5865]) );
  AND U4597 ( .A(p_input[5864]), .B(p_input[15864]), .Z(o[5864]) );
  AND U4598 ( .A(p_input[5863]), .B(p_input[15863]), .Z(o[5863]) );
  AND U4599 ( .A(p_input[5862]), .B(p_input[15862]), .Z(o[5862]) );
  AND U4600 ( .A(p_input[5861]), .B(p_input[15861]), .Z(o[5861]) );
  AND U4601 ( .A(p_input[5860]), .B(p_input[15860]), .Z(o[5860]) );
  AND U4602 ( .A(p_input[585]), .B(p_input[10585]), .Z(o[585]) );
  AND U4603 ( .A(p_input[5859]), .B(p_input[15859]), .Z(o[5859]) );
  AND U4604 ( .A(p_input[5858]), .B(p_input[15858]), .Z(o[5858]) );
  AND U4605 ( .A(p_input[5857]), .B(p_input[15857]), .Z(o[5857]) );
  AND U4606 ( .A(p_input[5856]), .B(p_input[15856]), .Z(o[5856]) );
  AND U4607 ( .A(p_input[5855]), .B(p_input[15855]), .Z(o[5855]) );
  AND U4608 ( .A(p_input[5854]), .B(p_input[15854]), .Z(o[5854]) );
  AND U4609 ( .A(p_input[5853]), .B(p_input[15853]), .Z(o[5853]) );
  AND U4610 ( .A(p_input[5852]), .B(p_input[15852]), .Z(o[5852]) );
  AND U4611 ( .A(p_input[5851]), .B(p_input[15851]), .Z(o[5851]) );
  AND U4612 ( .A(p_input[5850]), .B(p_input[15850]), .Z(o[5850]) );
  AND U4613 ( .A(p_input[584]), .B(p_input[10584]), .Z(o[584]) );
  AND U4614 ( .A(p_input[5849]), .B(p_input[15849]), .Z(o[5849]) );
  AND U4615 ( .A(p_input[5848]), .B(p_input[15848]), .Z(o[5848]) );
  AND U4616 ( .A(p_input[5847]), .B(p_input[15847]), .Z(o[5847]) );
  AND U4617 ( .A(p_input[5846]), .B(p_input[15846]), .Z(o[5846]) );
  AND U4618 ( .A(p_input[5845]), .B(p_input[15845]), .Z(o[5845]) );
  AND U4619 ( .A(p_input[5844]), .B(p_input[15844]), .Z(o[5844]) );
  AND U4620 ( .A(p_input[5843]), .B(p_input[15843]), .Z(o[5843]) );
  AND U4621 ( .A(p_input[5842]), .B(p_input[15842]), .Z(o[5842]) );
  AND U4622 ( .A(p_input[5841]), .B(p_input[15841]), .Z(o[5841]) );
  AND U4623 ( .A(p_input[5840]), .B(p_input[15840]), .Z(o[5840]) );
  AND U4624 ( .A(p_input[583]), .B(p_input[10583]), .Z(o[583]) );
  AND U4625 ( .A(p_input[5839]), .B(p_input[15839]), .Z(o[5839]) );
  AND U4626 ( .A(p_input[5838]), .B(p_input[15838]), .Z(o[5838]) );
  AND U4627 ( .A(p_input[5837]), .B(p_input[15837]), .Z(o[5837]) );
  AND U4628 ( .A(p_input[5836]), .B(p_input[15836]), .Z(o[5836]) );
  AND U4629 ( .A(p_input[5835]), .B(p_input[15835]), .Z(o[5835]) );
  AND U4630 ( .A(p_input[5834]), .B(p_input[15834]), .Z(o[5834]) );
  AND U4631 ( .A(p_input[5833]), .B(p_input[15833]), .Z(o[5833]) );
  AND U4632 ( .A(p_input[5832]), .B(p_input[15832]), .Z(o[5832]) );
  AND U4633 ( .A(p_input[5831]), .B(p_input[15831]), .Z(o[5831]) );
  AND U4634 ( .A(p_input[5830]), .B(p_input[15830]), .Z(o[5830]) );
  AND U4635 ( .A(p_input[582]), .B(p_input[10582]), .Z(o[582]) );
  AND U4636 ( .A(p_input[5829]), .B(p_input[15829]), .Z(o[5829]) );
  AND U4637 ( .A(p_input[5828]), .B(p_input[15828]), .Z(o[5828]) );
  AND U4638 ( .A(p_input[5827]), .B(p_input[15827]), .Z(o[5827]) );
  AND U4639 ( .A(p_input[5826]), .B(p_input[15826]), .Z(o[5826]) );
  AND U4640 ( .A(p_input[5825]), .B(p_input[15825]), .Z(o[5825]) );
  AND U4641 ( .A(p_input[5824]), .B(p_input[15824]), .Z(o[5824]) );
  AND U4642 ( .A(p_input[5823]), .B(p_input[15823]), .Z(o[5823]) );
  AND U4643 ( .A(p_input[5822]), .B(p_input[15822]), .Z(o[5822]) );
  AND U4644 ( .A(p_input[5821]), .B(p_input[15821]), .Z(o[5821]) );
  AND U4645 ( .A(p_input[5820]), .B(p_input[15820]), .Z(o[5820]) );
  AND U4646 ( .A(p_input[581]), .B(p_input[10581]), .Z(o[581]) );
  AND U4647 ( .A(p_input[5819]), .B(p_input[15819]), .Z(o[5819]) );
  AND U4648 ( .A(p_input[5818]), .B(p_input[15818]), .Z(o[5818]) );
  AND U4649 ( .A(p_input[5817]), .B(p_input[15817]), .Z(o[5817]) );
  AND U4650 ( .A(p_input[5816]), .B(p_input[15816]), .Z(o[5816]) );
  AND U4651 ( .A(p_input[5815]), .B(p_input[15815]), .Z(o[5815]) );
  AND U4652 ( .A(p_input[5814]), .B(p_input[15814]), .Z(o[5814]) );
  AND U4653 ( .A(p_input[5813]), .B(p_input[15813]), .Z(o[5813]) );
  AND U4654 ( .A(p_input[5812]), .B(p_input[15812]), .Z(o[5812]) );
  AND U4655 ( .A(p_input[5811]), .B(p_input[15811]), .Z(o[5811]) );
  AND U4656 ( .A(p_input[5810]), .B(p_input[15810]), .Z(o[5810]) );
  AND U4657 ( .A(p_input[580]), .B(p_input[10580]), .Z(o[580]) );
  AND U4658 ( .A(p_input[5809]), .B(p_input[15809]), .Z(o[5809]) );
  AND U4659 ( .A(p_input[5808]), .B(p_input[15808]), .Z(o[5808]) );
  AND U4660 ( .A(p_input[5807]), .B(p_input[15807]), .Z(o[5807]) );
  AND U4661 ( .A(p_input[5806]), .B(p_input[15806]), .Z(o[5806]) );
  AND U4662 ( .A(p_input[5805]), .B(p_input[15805]), .Z(o[5805]) );
  AND U4663 ( .A(p_input[5804]), .B(p_input[15804]), .Z(o[5804]) );
  AND U4664 ( .A(p_input[5803]), .B(p_input[15803]), .Z(o[5803]) );
  AND U4665 ( .A(p_input[5802]), .B(p_input[15802]), .Z(o[5802]) );
  AND U4666 ( .A(p_input[5801]), .B(p_input[15801]), .Z(o[5801]) );
  AND U4667 ( .A(p_input[5800]), .B(p_input[15800]), .Z(o[5800]) );
  AND U4668 ( .A(p_input[57]), .B(p_input[10057]), .Z(o[57]) );
  AND U4669 ( .A(p_input[579]), .B(p_input[10579]), .Z(o[579]) );
  AND U4670 ( .A(p_input[5799]), .B(p_input[15799]), .Z(o[5799]) );
  AND U4671 ( .A(p_input[5798]), .B(p_input[15798]), .Z(o[5798]) );
  AND U4672 ( .A(p_input[5797]), .B(p_input[15797]), .Z(o[5797]) );
  AND U4673 ( .A(p_input[5796]), .B(p_input[15796]), .Z(o[5796]) );
  AND U4674 ( .A(p_input[5795]), .B(p_input[15795]), .Z(o[5795]) );
  AND U4675 ( .A(p_input[5794]), .B(p_input[15794]), .Z(o[5794]) );
  AND U4676 ( .A(p_input[5793]), .B(p_input[15793]), .Z(o[5793]) );
  AND U4677 ( .A(p_input[5792]), .B(p_input[15792]), .Z(o[5792]) );
  AND U4678 ( .A(p_input[5791]), .B(p_input[15791]), .Z(o[5791]) );
  AND U4679 ( .A(p_input[5790]), .B(p_input[15790]), .Z(o[5790]) );
  AND U4680 ( .A(p_input[578]), .B(p_input[10578]), .Z(o[578]) );
  AND U4681 ( .A(p_input[5789]), .B(p_input[15789]), .Z(o[5789]) );
  AND U4682 ( .A(p_input[5788]), .B(p_input[15788]), .Z(o[5788]) );
  AND U4683 ( .A(p_input[5787]), .B(p_input[15787]), .Z(o[5787]) );
  AND U4684 ( .A(p_input[5786]), .B(p_input[15786]), .Z(o[5786]) );
  AND U4685 ( .A(p_input[5785]), .B(p_input[15785]), .Z(o[5785]) );
  AND U4686 ( .A(p_input[5784]), .B(p_input[15784]), .Z(o[5784]) );
  AND U4687 ( .A(p_input[5783]), .B(p_input[15783]), .Z(o[5783]) );
  AND U4688 ( .A(p_input[5782]), .B(p_input[15782]), .Z(o[5782]) );
  AND U4689 ( .A(p_input[5781]), .B(p_input[15781]), .Z(o[5781]) );
  AND U4690 ( .A(p_input[5780]), .B(p_input[15780]), .Z(o[5780]) );
  AND U4691 ( .A(p_input[577]), .B(p_input[10577]), .Z(o[577]) );
  AND U4692 ( .A(p_input[5779]), .B(p_input[15779]), .Z(o[5779]) );
  AND U4693 ( .A(p_input[5778]), .B(p_input[15778]), .Z(o[5778]) );
  AND U4694 ( .A(p_input[5777]), .B(p_input[15777]), .Z(o[5777]) );
  AND U4695 ( .A(p_input[5776]), .B(p_input[15776]), .Z(o[5776]) );
  AND U4696 ( .A(p_input[5775]), .B(p_input[15775]), .Z(o[5775]) );
  AND U4697 ( .A(p_input[5774]), .B(p_input[15774]), .Z(o[5774]) );
  AND U4698 ( .A(p_input[5773]), .B(p_input[15773]), .Z(o[5773]) );
  AND U4699 ( .A(p_input[5772]), .B(p_input[15772]), .Z(o[5772]) );
  AND U4700 ( .A(p_input[5771]), .B(p_input[15771]), .Z(o[5771]) );
  AND U4701 ( .A(p_input[5770]), .B(p_input[15770]), .Z(o[5770]) );
  AND U4702 ( .A(p_input[576]), .B(p_input[10576]), .Z(o[576]) );
  AND U4703 ( .A(p_input[5769]), .B(p_input[15769]), .Z(o[5769]) );
  AND U4704 ( .A(p_input[5768]), .B(p_input[15768]), .Z(o[5768]) );
  AND U4705 ( .A(p_input[5767]), .B(p_input[15767]), .Z(o[5767]) );
  AND U4706 ( .A(p_input[5766]), .B(p_input[15766]), .Z(o[5766]) );
  AND U4707 ( .A(p_input[5765]), .B(p_input[15765]), .Z(o[5765]) );
  AND U4708 ( .A(p_input[5764]), .B(p_input[15764]), .Z(o[5764]) );
  AND U4709 ( .A(p_input[5763]), .B(p_input[15763]), .Z(o[5763]) );
  AND U4710 ( .A(p_input[5762]), .B(p_input[15762]), .Z(o[5762]) );
  AND U4711 ( .A(p_input[5761]), .B(p_input[15761]), .Z(o[5761]) );
  AND U4712 ( .A(p_input[5760]), .B(p_input[15760]), .Z(o[5760]) );
  AND U4713 ( .A(p_input[575]), .B(p_input[10575]), .Z(o[575]) );
  AND U4714 ( .A(p_input[5759]), .B(p_input[15759]), .Z(o[5759]) );
  AND U4715 ( .A(p_input[5758]), .B(p_input[15758]), .Z(o[5758]) );
  AND U4716 ( .A(p_input[5757]), .B(p_input[15757]), .Z(o[5757]) );
  AND U4717 ( .A(p_input[5756]), .B(p_input[15756]), .Z(o[5756]) );
  AND U4718 ( .A(p_input[5755]), .B(p_input[15755]), .Z(o[5755]) );
  AND U4719 ( .A(p_input[5754]), .B(p_input[15754]), .Z(o[5754]) );
  AND U4720 ( .A(p_input[5753]), .B(p_input[15753]), .Z(o[5753]) );
  AND U4721 ( .A(p_input[5752]), .B(p_input[15752]), .Z(o[5752]) );
  AND U4722 ( .A(p_input[5751]), .B(p_input[15751]), .Z(o[5751]) );
  AND U4723 ( .A(p_input[5750]), .B(p_input[15750]), .Z(o[5750]) );
  AND U4724 ( .A(p_input[574]), .B(p_input[10574]), .Z(o[574]) );
  AND U4725 ( .A(p_input[5749]), .B(p_input[15749]), .Z(o[5749]) );
  AND U4726 ( .A(p_input[5748]), .B(p_input[15748]), .Z(o[5748]) );
  AND U4727 ( .A(p_input[5747]), .B(p_input[15747]), .Z(o[5747]) );
  AND U4728 ( .A(p_input[5746]), .B(p_input[15746]), .Z(o[5746]) );
  AND U4729 ( .A(p_input[5745]), .B(p_input[15745]), .Z(o[5745]) );
  AND U4730 ( .A(p_input[5744]), .B(p_input[15744]), .Z(o[5744]) );
  AND U4731 ( .A(p_input[5743]), .B(p_input[15743]), .Z(o[5743]) );
  AND U4732 ( .A(p_input[5742]), .B(p_input[15742]), .Z(o[5742]) );
  AND U4733 ( .A(p_input[5741]), .B(p_input[15741]), .Z(o[5741]) );
  AND U4734 ( .A(p_input[5740]), .B(p_input[15740]), .Z(o[5740]) );
  AND U4735 ( .A(p_input[573]), .B(p_input[10573]), .Z(o[573]) );
  AND U4736 ( .A(p_input[5739]), .B(p_input[15739]), .Z(o[5739]) );
  AND U4737 ( .A(p_input[5738]), .B(p_input[15738]), .Z(o[5738]) );
  AND U4738 ( .A(p_input[5737]), .B(p_input[15737]), .Z(o[5737]) );
  AND U4739 ( .A(p_input[5736]), .B(p_input[15736]), .Z(o[5736]) );
  AND U4740 ( .A(p_input[5735]), .B(p_input[15735]), .Z(o[5735]) );
  AND U4741 ( .A(p_input[5734]), .B(p_input[15734]), .Z(o[5734]) );
  AND U4742 ( .A(p_input[5733]), .B(p_input[15733]), .Z(o[5733]) );
  AND U4743 ( .A(p_input[5732]), .B(p_input[15732]), .Z(o[5732]) );
  AND U4744 ( .A(p_input[5731]), .B(p_input[15731]), .Z(o[5731]) );
  AND U4745 ( .A(p_input[5730]), .B(p_input[15730]), .Z(o[5730]) );
  AND U4746 ( .A(p_input[572]), .B(p_input[10572]), .Z(o[572]) );
  AND U4747 ( .A(p_input[5729]), .B(p_input[15729]), .Z(o[5729]) );
  AND U4748 ( .A(p_input[5728]), .B(p_input[15728]), .Z(o[5728]) );
  AND U4749 ( .A(p_input[5727]), .B(p_input[15727]), .Z(o[5727]) );
  AND U4750 ( .A(p_input[5726]), .B(p_input[15726]), .Z(o[5726]) );
  AND U4751 ( .A(p_input[5725]), .B(p_input[15725]), .Z(o[5725]) );
  AND U4752 ( .A(p_input[5724]), .B(p_input[15724]), .Z(o[5724]) );
  AND U4753 ( .A(p_input[5723]), .B(p_input[15723]), .Z(o[5723]) );
  AND U4754 ( .A(p_input[5722]), .B(p_input[15722]), .Z(o[5722]) );
  AND U4755 ( .A(p_input[5721]), .B(p_input[15721]), .Z(o[5721]) );
  AND U4756 ( .A(p_input[5720]), .B(p_input[15720]), .Z(o[5720]) );
  AND U4757 ( .A(p_input[571]), .B(p_input[10571]), .Z(o[571]) );
  AND U4758 ( .A(p_input[5719]), .B(p_input[15719]), .Z(o[5719]) );
  AND U4759 ( .A(p_input[5718]), .B(p_input[15718]), .Z(o[5718]) );
  AND U4760 ( .A(p_input[5717]), .B(p_input[15717]), .Z(o[5717]) );
  AND U4761 ( .A(p_input[5716]), .B(p_input[15716]), .Z(o[5716]) );
  AND U4762 ( .A(p_input[5715]), .B(p_input[15715]), .Z(o[5715]) );
  AND U4763 ( .A(p_input[5714]), .B(p_input[15714]), .Z(o[5714]) );
  AND U4764 ( .A(p_input[5713]), .B(p_input[15713]), .Z(o[5713]) );
  AND U4765 ( .A(p_input[5712]), .B(p_input[15712]), .Z(o[5712]) );
  AND U4766 ( .A(p_input[5711]), .B(p_input[15711]), .Z(o[5711]) );
  AND U4767 ( .A(p_input[5710]), .B(p_input[15710]), .Z(o[5710]) );
  AND U4768 ( .A(p_input[570]), .B(p_input[10570]), .Z(o[570]) );
  AND U4769 ( .A(p_input[5709]), .B(p_input[15709]), .Z(o[5709]) );
  AND U4770 ( .A(p_input[5708]), .B(p_input[15708]), .Z(o[5708]) );
  AND U4771 ( .A(p_input[5707]), .B(p_input[15707]), .Z(o[5707]) );
  AND U4772 ( .A(p_input[5706]), .B(p_input[15706]), .Z(o[5706]) );
  AND U4773 ( .A(p_input[5705]), .B(p_input[15705]), .Z(o[5705]) );
  AND U4774 ( .A(p_input[5704]), .B(p_input[15704]), .Z(o[5704]) );
  AND U4775 ( .A(p_input[5703]), .B(p_input[15703]), .Z(o[5703]) );
  AND U4776 ( .A(p_input[5702]), .B(p_input[15702]), .Z(o[5702]) );
  AND U4777 ( .A(p_input[5701]), .B(p_input[15701]), .Z(o[5701]) );
  AND U4778 ( .A(p_input[5700]), .B(p_input[15700]), .Z(o[5700]) );
  AND U4779 ( .A(p_input[56]), .B(p_input[10056]), .Z(o[56]) );
  AND U4780 ( .A(p_input[569]), .B(p_input[10569]), .Z(o[569]) );
  AND U4781 ( .A(p_input[5699]), .B(p_input[15699]), .Z(o[5699]) );
  AND U4782 ( .A(p_input[5698]), .B(p_input[15698]), .Z(o[5698]) );
  AND U4783 ( .A(p_input[5697]), .B(p_input[15697]), .Z(o[5697]) );
  AND U4784 ( .A(p_input[5696]), .B(p_input[15696]), .Z(o[5696]) );
  AND U4785 ( .A(p_input[5695]), .B(p_input[15695]), .Z(o[5695]) );
  AND U4786 ( .A(p_input[5694]), .B(p_input[15694]), .Z(o[5694]) );
  AND U4787 ( .A(p_input[5693]), .B(p_input[15693]), .Z(o[5693]) );
  AND U4788 ( .A(p_input[5692]), .B(p_input[15692]), .Z(o[5692]) );
  AND U4789 ( .A(p_input[5691]), .B(p_input[15691]), .Z(o[5691]) );
  AND U4790 ( .A(p_input[5690]), .B(p_input[15690]), .Z(o[5690]) );
  AND U4791 ( .A(p_input[568]), .B(p_input[10568]), .Z(o[568]) );
  AND U4792 ( .A(p_input[5689]), .B(p_input[15689]), .Z(o[5689]) );
  AND U4793 ( .A(p_input[5688]), .B(p_input[15688]), .Z(o[5688]) );
  AND U4794 ( .A(p_input[5687]), .B(p_input[15687]), .Z(o[5687]) );
  AND U4795 ( .A(p_input[5686]), .B(p_input[15686]), .Z(o[5686]) );
  AND U4796 ( .A(p_input[5685]), .B(p_input[15685]), .Z(o[5685]) );
  AND U4797 ( .A(p_input[5684]), .B(p_input[15684]), .Z(o[5684]) );
  AND U4798 ( .A(p_input[5683]), .B(p_input[15683]), .Z(o[5683]) );
  AND U4799 ( .A(p_input[5682]), .B(p_input[15682]), .Z(o[5682]) );
  AND U4800 ( .A(p_input[5681]), .B(p_input[15681]), .Z(o[5681]) );
  AND U4801 ( .A(p_input[5680]), .B(p_input[15680]), .Z(o[5680]) );
  AND U4802 ( .A(p_input[567]), .B(p_input[10567]), .Z(o[567]) );
  AND U4803 ( .A(p_input[5679]), .B(p_input[15679]), .Z(o[5679]) );
  AND U4804 ( .A(p_input[5678]), .B(p_input[15678]), .Z(o[5678]) );
  AND U4805 ( .A(p_input[5677]), .B(p_input[15677]), .Z(o[5677]) );
  AND U4806 ( .A(p_input[5676]), .B(p_input[15676]), .Z(o[5676]) );
  AND U4807 ( .A(p_input[5675]), .B(p_input[15675]), .Z(o[5675]) );
  AND U4808 ( .A(p_input[5674]), .B(p_input[15674]), .Z(o[5674]) );
  AND U4809 ( .A(p_input[5673]), .B(p_input[15673]), .Z(o[5673]) );
  AND U4810 ( .A(p_input[5672]), .B(p_input[15672]), .Z(o[5672]) );
  AND U4811 ( .A(p_input[5671]), .B(p_input[15671]), .Z(o[5671]) );
  AND U4812 ( .A(p_input[5670]), .B(p_input[15670]), .Z(o[5670]) );
  AND U4813 ( .A(p_input[566]), .B(p_input[10566]), .Z(o[566]) );
  AND U4814 ( .A(p_input[5669]), .B(p_input[15669]), .Z(o[5669]) );
  AND U4815 ( .A(p_input[5668]), .B(p_input[15668]), .Z(o[5668]) );
  AND U4816 ( .A(p_input[5667]), .B(p_input[15667]), .Z(o[5667]) );
  AND U4817 ( .A(p_input[5666]), .B(p_input[15666]), .Z(o[5666]) );
  AND U4818 ( .A(p_input[5665]), .B(p_input[15665]), .Z(o[5665]) );
  AND U4819 ( .A(p_input[5664]), .B(p_input[15664]), .Z(o[5664]) );
  AND U4820 ( .A(p_input[5663]), .B(p_input[15663]), .Z(o[5663]) );
  AND U4821 ( .A(p_input[5662]), .B(p_input[15662]), .Z(o[5662]) );
  AND U4822 ( .A(p_input[5661]), .B(p_input[15661]), .Z(o[5661]) );
  AND U4823 ( .A(p_input[5660]), .B(p_input[15660]), .Z(o[5660]) );
  AND U4824 ( .A(p_input[565]), .B(p_input[10565]), .Z(o[565]) );
  AND U4825 ( .A(p_input[5659]), .B(p_input[15659]), .Z(o[5659]) );
  AND U4826 ( .A(p_input[5658]), .B(p_input[15658]), .Z(o[5658]) );
  AND U4827 ( .A(p_input[5657]), .B(p_input[15657]), .Z(o[5657]) );
  AND U4828 ( .A(p_input[5656]), .B(p_input[15656]), .Z(o[5656]) );
  AND U4829 ( .A(p_input[5655]), .B(p_input[15655]), .Z(o[5655]) );
  AND U4830 ( .A(p_input[5654]), .B(p_input[15654]), .Z(o[5654]) );
  AND U4831 ( .A(p_input[5653]), .B(p_input[15653]), .Z(o[5653]) );
  AND U4832 ( .A(p_input[5652]), .B(p_input[15652]), .Z(o[5652]) );
  AND U4833 ( .A(p_input[5651]), .B(p_input[15651]), .Z(o[5651]) );
  AND U4834 ( .A(p_input[5650]), .B(p_input[15650]), .Z(o[5650]) );
  AND U4835 ( .A(p_input[564]), .B(p_input[10564]), .Z(o[564]) );
  AND U4836 ( .A(p_input[5649]), .B(p_input[15649]), .Z(o[5649]) );
  AND U4837 ( .A(p_input[5648]), .B(p_input[15648]), .Z(o[5648]) );
  AND U4838 ( .A(p_input[5647]), .B(p_input[15647]), .Z(o[5647]) );
  AND U4839 ( .A(p_input[5646]), .B(p_input[15646]), .Z(o[5646]) );
  AND U4840 ( .A(p_input[5645]), .B(p_input[15645]), .Z(o[5645]) );
  AND U4841 ( .A(p_input[5644]), .B(p_input[15644]), .Z(o[5644]) );
  AND U4842 ( .A(p_input[5643]), .B(p_input[15643]), .Z(o[5643]) );
  AND U4843 ( .A(p_input[5642]), .B(p_input[15642]), .Z(o[5642]) );
  AND U4844 ( .A(p_input[5641]), .B(p_input[15641]), .Z(o[5641]) );
  AND U4845 ( .A(p_input[5640]), .B(p_input[15640]), .Z(o[5640]) );
  AND U4846 ( .A(p_input[563]), .B(p_input[10563]), .Z(o[563]) );
  AND U4847 ( .A(p_input[5639]), .B(p_input[15639]), .Z(o[5639]) );
  AND U4848 ( .A(p_input[5638]), .B(p_input[15638]), .Z(o[5638]) );
  AND U4849 ( .A(p_input[5637]), .B(p_input[15637]), .Z(o[5637]) );
  AND U4850 ( .A(p_input[5636]), .B(p_input[15636]), .Z(o[5636]) );
  AND U4851 ( .A(p_input[5635]), .B(p_input[15635]), .Z(o[5635]) );
  AND U4852 ( .A(p_input[5634]), .B(p_input[15634]), .Z(o[5634]) );
  AND U4853 ( .A(p_input[5633]), .B(p_input[15633]), .Z(o[5633]) );
  AND U4854 ( .A(p_input[5632]), .B(p_input[15632]), .Z(o[5632]) );
  AND U4855 ( .A(p_input[5631]), .B(p_input[15631]), .Z(o[5631]) );
  AND U4856 ( .A(p_input[5630]), .B(p_input[15630]), .Z(o[5630]) );
  AND U4857 ( .A(p_input[562]), .B(p_input[10562]), .Z(o[562]) );
  AND U4858 ( .A(p_input[5629]), .B(p_input[15629]), .Z(o[5629]) );
  AND U4859 ( .A(p_input[5628]), .B(p_input[15628]), .Z(o[5628]) );
  AND U4860 ( .A(p_input[5627]), .B(p_input[15627]), .Z(o[5627]) );
  AND U4861 ( .A(p_input[5626]), .B(p_input[15626]), .Z(o[5626]) );
  AND U4862 ( .A(p_input[5625]), .B(p_input[15625]), .Z(o[5625]) );
  AND U4863 ( .A(p_input[5624]), .B(p_input[15624]), .Z(o[5624]) );
  AND U4864 ( .A(p_input[5623]), .B(p_input[15623]), .Z(o[5623]) );
  AND U4865 ( .A(p_input[5622]), .B(p_input[15622]), .Z(o[5622]) );
  AND U4866 ( .A(p_input[5621]), .B(p_input[15621]), .Z(o[5621]) );
  AND U4867 ( .A(p_input[5620]), .B(p_input[15620]), .Z(o[5620]) );
  AND U4868 ( .A(p_input[561]), .B(p_input[10561]), .Z(o[561]) );
  AND U4869 ( .A(p_input[5619]), .B(p_input[15619]), .Z(o[5619]) );
  AND U4870 ( .A(p_input[5618]), .B(p_input[15618]), .Z(o[5618]) );
  AND U4871 ( .A(p_input[5617]), .B(p_input[15617]), .Z(o[5617]) );
  AND U4872 ( .A(p_input[5616]), .B(p_input[15616]), .Z(o[5616]) );
  AND U4873 ( .A(p_input[5615]), .B(p_input[15615]), .Z(o[5615]) );
  AND U4874 ( .A(p_input[5614]), .B(p_input[15614]), .Z(o[5614]) );
  AND U4875 ( .A(p_input[5613]), .B(p_input[15613]), .Z(o[5613]) );
  AND U4876 ( .A(p_input[5612]), .B(p_input[15612]), .Z(o[5612]) );
  AND U4877 ( .A(p_input[5611]), .B(p_input[15611]), .Z(o[5611]) );
  AND U4878 ( .A(p_input[5610]), .B(p_input[15610]), .Z(o[5610]) );
  AND U4879 ( .A(p_input[560]), .B(p_input[10560]), .Z(o[560]) );
  AND U4880 ( .A(p_input[5609]), .B(p_input[15609]), .Z(o[5609]) );
  AND U4881 ( .A(p_input[5608]), .B(p_input[15608]), .Z(o[5608]) );
  AND U4882 ( .A(p_input[5607]), .B(p_input[15607]), .Z(o[5607]) );
  AND U4883 ( .A(p_input[5606]), .B(p_input[15606]), .Z(o[5606]) );
  AND U4884 ( .A(p_input[5605]), .B(p_input[15605]), .Z(o[5605]) );
  AND U4885 ( .A(p_input[5604]), .B(p_input[15604]), .Z(o[5604]) );
  AND U4886 ( .A(p_input[5603]), .B(p_input[15603]), .Z(o[5603]) );
  AND U4887 ( .A(p_input[5602]), .B(p_input[15602]), .Z(o[5602]) );
  AND U4888 ( .A(p_input[5601]), .B(p_input[15601]), .Z(o[5601]) );
  AND U4889 ( .A(p_input[5600]), .B(p_input[15600]), .Z(o[5600]) );
  AND U4890 ( .A(p_input[55]), .B(p_input[10055]), .Z(o[55]) );
  AND U4891 ( .A(p_input[559]), .B(p_input[10559]), .Z(o[559]) );
  AND U4892 ( .A(p_input[5599]), .B(p_input[15599]), .Z(o[5599]) );
  AND U4893 ( .A(p_input[5598]), .B(p_input[15598]), .Z(o[5598]) );
  AND U4894 ( .A(p_input[5597]), .B(p_input[15597]), .Z(o[5597]) );
  AND U4895 ( .A(p_input[5596]), .B(p_input[15596]), .Z(o[5596]) );
  AND U4896 ( .A(p_input[5595]), .B(p_input[15595]), .Z(o[5595]) );
  AND U4897 ( .A(p_input[5594]), .B(p_input[15594]), .Z(o[5594]) );
  AND U4898 ( .A(p_input[5593]), .B(p_input[15593]), .Z(o[5593]) );
  AND U4899 ( .A(p_input[5592]), .B(p_input[15592]), .Z(o[5592]) );
  AND U4900 ( .A(p_input[5591]), .B(p_input[15591]), .Z(o[5591]) );
  AND U4901 ( .A(p_input[5590]), .B(p_input[15590]), .Z(o[5590]) );
  AND U4902 ( .A(p_input[558]), .B(p_input[10558]), .Z(o[558]) );
  AND U4903 ( .A(p_input[5589]), .B(p_input[15589]), .Z(o[5589]) );
  AND U4904 ( .A(p_input[5588]), .B(p_input[15588]), .Z(o[5588]) );
  AND U4905 ( .A(p_input[5587]), .B(p_input[15587]), .Z(o[5587]) );
  AND U4906 ( .A(p_input[5586]), .B(p_input[15586]), .Z(o[5586]) );
  AND U4907 ( .A(p_input[5585]), .B(p_input[15585]), .Z(o[5585]) );
  AND U4908 ( .A(p_input[5584]), .B(p_input[15584]), .Z(o[5584]) );
  AND U4909 ( .A(p_input[5583]), .B(p_input[15583]), .Z(o[5583]) );
  AND U4910 ( .A(p_input[5582]), .B(p_input[15582]), .Z(o[5582]) );
  AND U4911 ( .A(p_input[5581]), .B(p_input[15581]), .Z(o[5581]) );
  AND U4912 ( .A(p_input[5580]), .B(p_input[15580]), .Z(o[5580]) );
  AND U4913 ( .A(p_input[557]), .B(p_input[10557]), .Z(o[557]) );
  AND U4914 ( .A(p_input[5579]), .B(p_input[15579]), .Z(o[5579]) );
  AND U4915 ( .A(p_input[5578]), .B(p_input[15578]), .Z(o[5578]) );
  AND U4916 ( .A(p_input[5577]), .B(p_input[15577]), .Z(o[5577]) );
  AND U4917 ( .A(p_input[5576]), .B(p_input[15576]), .Z(o[5576]) );
  AND U4918 ( .A(p_input[5575]), .B(p_input[15575]), .Z(o[5575]) );
  AND U4919 ( .A(p_input[5574]), .B(p_input[15574]), .Z(o[5574]) );
  AND U4920 ( .A(p_input[5573]), .B(p_input[15573]), .Z(o[5573]) );
  AND U4921 ( .A(p_input[5572]), .B(p_input[15572]), .Z(o[5572]) );
  AND U4922 ( .A(p_input[5571]), .B(p_input[15571]), .Z(o[5571]) );
  AND U4923 ( .A(p_input[5570]), .B(p_input[15570]), .Z(o[5570]) );
  AND U4924 ( .A(p_input[556]), .B(p_input[10556]), .Z(o[556]) );
  AND U4925 ( .A(p_input[5569]), .B(p_input[15569]), .Z(o[5569]) );
  AND U4926 ( .A(p_input[5568]), .B(p_input[15568]), .Z(o[5568]) );
  AND U4927 ( .A(p_input[5567]), .B(p_input[15567]), .Z(o[5567]) );
  AND U4928 ( .A(p_input[5566]), .B(p_input[15566]), .Z(o[5566]) );
  AND U4929 ( .A(p_input[5565]), .B(p_input[15565]), .Z(o[5565]) );
  AND U4930 ( .A(p_input[5564]), .B(p_input[15564]), .Z(o[5564]) );
  AND U4931 ( .A(p_input[5563]), .B(p_input[15563]), .Z(o[5563]) );
  AND U4932 ( .A(p_input[5562]), .B(p_input[15562]), .Z(o[5562]) );
  AND U4933 ( .A(p_input[5561]), .B(p_input[15561]), .Z(o[5561]) );
  AND U4934 ( .A(p_input[5560]), .B(p_input[15560]), .Z(o[5560]) );
  AND U4935 ( .A(p_input[555]), .B(p_input[10555]), .Z(o[555]) );
  AND U4936 ( .A(p_input[5559]), .B(p_input[15559]), .Z(o[5559]) );
  AND U4937 ( .A(p_input[5558]), .B(p_input[15558]), .Z(o[5558]) );
  AND U4938 ( .A(p_input[5557]), .B(p_input[15557]), .Z(o[5557]) );
  AND U4939 ( .A(p_input[5556]), .B(p_input[15556]), .Z(o[5556]) );
  AND U4940 ( .A(p_input[5555]), .B(p_input[15555]), .Z(o[5555]) );
  AND U4941 ( .A(p_input[5554]), .B(p_input[15554]), .Z(o[5554]) );
  AND U4942 ( .A(p_input[5553]), .B(p_input[15553]), .Z(o[5553]) );
  AND U4943 ( .A(p_input[5552]), .B(p_input[15552]), .Z(o[5552]) );
  AND U4944 ( .A(p_input[5551]), .B(p_input[15551]), .Z(o[5551]) );
  AND U4945 ( .A(p_input[5550]), .B(p_input[15550]), .Z(o[5550]) );
  AND U4946 ( .A(p_input[554]), .B(p_input[10554]), .Z(o[554]) );
  AND U4947 ( .A(p_input[5549]), .B(p_input[15549]), .Z(o[5549]) );
  AND U4948 ( .A(p_input[5548]), .B(p_input[15548]), .Z(o[5548]) );
  AND U4949 ( .A(p_input[5547]), .B(p_input[15547]), .Z(o[5547]) );
  AND U4950 ( .A(p_input[5546]), .B(p_input[15546]), .Z(o[5546]) );
  AND U4951 ( .A(p_input[5545]), .B(p_input[15545]), .Z(o[5545]) );
  AND U4952 ( .A(p_input[5544]), .B(p_input[15544]), .Z(o[5544]) );
  AND U4953 ( .A(p_input[5543]), .B(p_input[15543]), .Z(o[5543]) );
  AND U4954 ( .A(p_input[5542]), .B(p_input[15542]), .Z(o[5542]) );
  AND U4955 ( .A(p_input[5541]), .B(p_input[15541]), .Z(o[5541]) );
  AND U4956 ( .A(p_input[5540]), .B(p_input[15540]), .Z(o[5540]) );
  AND U4957 ( .A(p_input[553]), .B(p_input[10553]), .Z(o[553]) );
  AND U4958 ( .A(p_input[5539]), .B(p_input[15539]), .Z(o[5539]) );
  AND U4959 ( .A(p_input[5538]), .B(p_input[15538]), .Z(o[5538]) );
  AND U4960 ( .A(p_input[5537]), .B(p_input[15537]), .Z(o[5537]) );
  AND U4961 ( .A(p_input[5536]), .B(p_input[15536]), .Z(o[5536]) );
  AND U4962 ( .A(p_input[5535]), .B(p_input[15535]), .Z(o[5535]) );
  AND U4963 ( .A(p_input[5534]), .B(p_input[15534]), .Z(o[5534]) );
  AND U4964 ( .A(p_input[5533]), .B(p_input[15533]), .Z(o[5533]) );
  AND U4965 ( .A(p_input[5532]), .B(p_input[15532]), .Z(o[5532]) );
  AND U4966 ( .A(p_input[5531]), .B(p_input[15531]), .Z(o[5531]) );
  AND U4967 ( .A(p_input[5530]), .B(p_input[15530]), .Z(o[5530]) );
  AND U4968 ( .A(p_input[552]), .B(p_input[10552]), .Z(o[552]) );
  AND U4969 ( .A(p_input[5529]), .B(p_input[15529]), .Z(o[5529]) );
  AND U4970 ( .A(p_input[5528]), .B(p_input[15528]), .Z(o[5528]) );
  AND U4971 ( .A(p_input[5527]), .B(p_input[15527]), .Z(o[5527]) );
  AND U4972 ( .A(p_input[5526]), .B(p_input[15526]), .Z(o[5526]) );
  AND U4973 ( .A(p_input[5525]), .B(p_input[15525]), .Z(o[5525]) );
  AND U4974 ( .A(p_input[5524]), .B(p_input[15524]), .Z(o[5524]) );
  AND U4975 ( .A(p_input[5523]), .B(p_input[15523]), .Z(o[5523]) );
  AND U4976 ( .A(p_input[5522]), .B(p_input[15522]), .Z(o[5522]) );
  AND U4977 ( .A(p_input[5521]), .B(p_input[15521]), .Z(o[5521]) );
  AND U4978 ( .A(p_input[5520]), .B(p_input[15520]), .Z(o[5520]) );
  AND U4979 ( .A(p_input[551]), .B(p_input[10551]), .Z(o[551]) );
  AND U4980 ( .A(p_input[5519]), .B(p_input[15519]), .Z(o[5519]) );
  AND U4981 ( .A(p_input[5518]), .B(p_input[15518]), .Z(o[5518]) );
  AND U4982 ( .A(p_input[5517]), .B(p_input[15517]), .Z(o[5517]) );
  AND U4983 ( .A(p_input[5516]), .B(p_input[15516]), .Z(o[5516]) );
  AND U4984 ( .A(p_input[5515]), .B(p_input[15515]), .Z(o[5515]) );
  AND U4985 ( .A(p_input[5514]), .B(p_input[15514]), .Z(o[5514]) );
  AND U4986 ( .A(p_input[5513]), .B(p_input[15513]), .Z(o[5513]) );
  AND U4987 ( .A(p_input[5512]), .B(p_input[15512]), .Z(o[5512]) );
  AND U4988 ( .A(p_input[5511]), .B(p_input[15511]), .Z(o[5511]) );
  AND U4989 ( .A(p_input[5510]), .B(p_input[15510]), .Z(o[5510]) );
  AND U4990 ( .A(p_input[550]), .B(p_input[10550]), .Z(o[550]) );
  AND U4991 ( .A(p_input[5509]), .B(p_input[15509]), .Z(o[5509]) );
  AND U4992 ( .A(p_input[5508]), .B(p_input[15508]), .Z(o[5508]) );
  AND U4993 ( .A(p_input[5507]), .B(p_input[15507]), .Z(o[5507]) );
  AND U4994 ( .A(p_input[5506]), .B(p_input[15506]), .Z(o[5506]) );
  AND U4995 ( .A(p_input[5505]), .B(p_input[15505]), .Z(o[5505]) );
  AND U4996 ( .A(p_input[5504]), .B(p_input[15504]), .Z(o[5504]) );
  AND U4997 ( .A(p_input[5503]), .B(p_input[15503]), .Z(o[5503]) );
  AND U4998 ( .A(p_input[5502]), .B(p_input[15502]), .Z(o[5502]) );
  AND U4999 ( .A(p_input[5501]), .B(p_input[15501]), .Z(o[5501]) );
  AND U5000 ( .A(p_input[5500]), .B(p_input[15500]), .Z(o[5500]) );
  AND U5001 ( .A(p_input[54]), .B(p_input[10054]), .Z(o[54]) );
  AND U5002 ( .A(p_input[549]), .B(p_input[10549]), .Z(o[549]) );
  AND U5003 ( .A(p_input[5499]), .B(p_input[15499]), .Z(o[5499]) );
  AND U5004 ( .A(p_input[5498]), .B(p_input[15498]), .Z(o[5498]) );
  AND U5005 ( .A(p_input[5497]), .B(p_input[15497]), .Z(o[5497]) );
  AND U5006 ( .A(p_input[5496]), .B(p_input[15496]), .Z(o[5496]) );
  AND U5007 ( .A(p_input[5495]), .B(p_input[15495]), .Z(o[5495]) );
  AND U5008 ( .A(p_input[5494]), .B(p_input[15494]), .Z(o[5494]) );
  AND U5009 ( .A(p_input[5493]), .B(p_input[15493]), .Z(o[5493]) );
  AND U5010 ( .A(p_input[5492]), .B(p_input[15492]), .Z(o[5492]) );
  AND U5011 ( .A(p_input[5491]), .B(p_input[15491]), .Z(o[5491]) );
  AND U5012 ( .A(p_input[5490]), .B(p_input[15490]), .Z(o[5490]) );
  AND U5013 ( .A(p_input[548]), .B(p_input[10548]), .Z(o[548]) );
  AND U5014 ( .A(p_input[5489]), .B(p_input[15489]), .Z(o[5489]) );
  AND U5015 ( .A(p_input[5488]), .B(p_input[15488]), .Z(o[5488]) );
  AND U5016 ( .A(p_input[5487]), .B(p_input[15487]), .Z(o[5487]) );
  AND U5017 ( .A(p_input[5486]), .B(p_input[15486]), .Z(o[5486]) );
  AND U5018 ( .A(p_input[5485]), .B(p_input[15485]), .Z(o[5485]) );
  AND U5019 ( .A(p_input[5484]), .B(p_input[15484]), .Z(o[5484]) );
  AND U5020 ( .A(p_input[5483]), .B(p_input[15483]), .Z(o[5483]) );
  AND U5021 ( .A(p_input[5482]), .B(p_input[15482]), .Z(o[5482]) );
  AND U5022 ( .A(p_input[5481]), .B(p_input[15481]), .Z(o[5481]) );
  AND U5023 ( .A(p_input[5480]), .B(p_input[15480]), .Z(o[5480]) );
  AND U5024 ( .A(p_input[547]), .B(p_input[10547]), .Z(o[547]) );
  AND U5025 ( .A(p_input[5479]), .B(p_input[15479]), .Z(o[5479]) );
  AND U5026 ( .A(p_input[5478]), .B(p_input[15478]), .Z(o[5478]) );
  AND U5027 ( .A(p_input[5477]), .B(p_input[15477]), .Z(o[5477]) );
  AND U5028 ( .A(p_input[5476]), .B(p_input[15476]), .Z(o[5476]) );
  AND U5029 ( .A(p_input[5475]), .B(p_input[15475]), .Z(o[5475]) );
  AND U5030 ( .A(p_input[5474]), .B(p_input[15474]), .Z(o[5474]) );
  AND U5031 ( .A(p_input[5473]), .B(p_input[15473]), .Z(o[5473]) );
  AND U5032 ( .A(p_input[5472]), .B(p_input[15472]), .Z(o[5472]) );
  AND U5033 ( .A(p_input[5471]), .B(p_input[15471]), .Z(o[5471]) );
  AND U5034 ( .A(p_input[5470]), .B(p_input[15470]), .Z(o[5470]) );
  AND U5035 ( .A(p_input[546]), .B(p_input[10546]), .Z(o[546]) );
  AND U5036 ( .A(p_input[5469]), .B(p_input[15469]), .Z(o[5469]) );
  AND U5037 ( .A(p_input[5468]), .B(p_input[15468]), .Z(o[5468]) );
  AND U5038 ( .A(p_input[5467]), .B(p_input[15467]), .Z(o[5467]) );
  AND U5039 ( .A(p_input[5466]), .B(p_input[15466]), .Z(o[5466]) );
  AND U5040 ( .A(p_input[5465]), .B(p_input[15465]), .Z(o[5465]) );
  AND U5041 ( .A(p_input[5464]), .B(p_input[15464]), .Z(o[5464]) );
  AND U5042 ( .A(p_input[5463]), .B(p_input[15463]), .Z(o[5463]) );
  AND U5043 ( .A(p_input[5462]), .B(p_input[15462]), .Z(o[5462]) );
  AND U5044 ( .A(p_input[5461]), .B(p_input[15461]), .Z(o[5461]) );
  AND U5045 ( .A(p_input[5460]), .B(p_input[15460]), .Z(o[5460]) );
  AND U5046 ( .A(p_input[545]), .B(p_input[10545]), .Z(o[545]) );
  AND U5047 ( .A(p_input[5459]), .B(p_input[15459]), .Z(o[5459]) );
  AND U5048 ( .A(p_input[5458]), .B(p_input[15458]), .Z(o[5458]) );
  AND U5049 ( .A(p_input[5457]), .B(p_input[15457]), .Z(o[5457]) );
  AND U5050 ( .A(p_input[5456]), .B(p_input[15456]), .Z(o[5456]) );
  AND U5051 ( .A(p_input[5455]), .B(p_input[15455]), .Z(o[5455]) );
  AND U5052 ( .A(p_input[5454]), .B(p_input[15454]), .Z(o[5454]) );
  AND U5053 ( .A(p_input[5453]), .B(p_input[15453]), .Z(o[5453]) );
  AND U5054 ( .A(p_input[5452]), .B(p_input[15452]), .Z(o[5452]) );
  AND U5055 ( .A(p_input[5451]), .B(p_input[15451]), .Z(o[5451]) );
  AND U5056 ( .A(p_input[5450]), .B(p_input[15450]), .Z(o[5450]) );
  AND U5057 ( .A(p_input[544]), .B(p_input[10544]), .Z(o[544]) );
  AND U5058 ( .A(p_input[5449]), .B(p_input[15449]), .Z(o[5449]) );
  AND U5059 ( .A(p_input[5448]), .B(p_input[15448]), .Z(o[5448]) );
  AND U5060 ( .A(p_input[5447]), .B(p_input[15447]), .Z(o[5447]) );
  AND U5061 ( .A(p_input[5446]), .B(p_input[15446]), .Z(o[5446]) );
  AND U5062 ( .A(p_input[5445]), .B(p_input[15445]), .Z(o[5445]) );
  AND U5063 ( .A(p_input[5444]), .B(p_input[15444]), .Z(o[5444]) );
  AND U5064 ( .A(p_input[5443]), .B(p_input[15443]), .Z(o[5443]) );
  AND U5065 ( .A(p_input[5442]), .B(p_input[15442]), .Z(o[5442]) );
  AND U5066 ( .A(p_input[5441]), .B(p_input[15441]), .Z(o[5441]) );
  AND U5067 ( .A(p_input[5440]), .B(p_input[15440]), .Z(o[5440]) );
  AND U5068 ( .A(p_input[543]), .B(p_input[10543]), .Z(o[543]) );
  AND U5069 ( .A(p_input[5439]), .B(p_input[15439]), .Z(o[5439]) );
  AND U5070 ( .A(p_input[5438]), .B(p_input[15438]), .Z(o[5438]) );
  AND U5071 ( .A(p_input[5437]), .B(p_input[15437]), .Z(o[5437]) );
  AND U5072 ( .A(p_input[5436]), .B(p_input[15436]), .Z(o[5436]) );
  AND U5073 ( .A(p_input[5435]), .B(p_input[15435]), .Z(o[5435]) );
  AND U5074 ( .A(p_input[5434]), .B(p_input[15434]), .Z(o[5434]) );
  AND U5075 ( .A(p_input[5433]), .B(p_input[15433]), .Z(o[5433]) );
  AND U5076 ( .A(p_input[5432]), .B(p_input[15432]), .Z(o[5432]) );
  AND U5077 ( .A(p_input[5431]), .B(p_input[15431]), .Z(o[5431]) );
  AND U5078 ( .A(p_input[5430]), .B(p_input[15430]), .Z(o[5430]) );
  AND U5079 ( .A(p_input[542]), .B(p_input[10542]), .Z(o[542]) );
  AND U5080 ( .A(p_input[5429]), .B(p_input[15429]), .Z(o[5429]) );
  AND U5081 ( .A(p_input[5428]), .B(p_input[15428]), .Z(o[5428]) );
  AND U5082 ( .A(p_input[5427]), .B(p_input[15427]), .Z(o[5427]) );
  AND U5083 ( .A(p_input[5426]), .B(p_input[15426]), .Z(o[5426]) );
  AND U5084 ( .A(p_input[5425]), .B(p_input[15425]), .Z(o[5425]) );
  AND U5085 ( .A(p_input[5424]), .B(p_input[15424]), .Z(o[5424]) );
  AND U5086 ( .A(p_input[5423]), .B(p_input[15423]), .Z(o[5423]) );
  AND U5087 ( .A(p_input[5422]), .B(p_input[15422]), .Z(o[5422]) );
  AND U5088 ( .A(p_input[5421]), .B(p_input[15421]), .Z(o[5421]) );
  AND U5089 ( .A(p_input[5420]), .B(p_input[15420]), .Z(o[5420]) );
  AND U5090 ( .A(p_input[541]), .B(p_input[10541]), .Z(o[541]) );
  AND U5091 ( .A(p_input[5419]), .B(p_input[15419]), .Z(o[5419]) );
  AND U5092 ( .A(p_input[5418]), .B(p_input[15418]), .Z(o[5418]) );
  AND U5093 ( .A(p_input[5417]), .B(p_input[15417]), .Z(o[5417]) );
  AND U5094 ( .A(p_input[5416]), .B(p_input[15416]), .Z(o[5416]) );
  AND U5095 ( .A(p_input[5415]), .B(p_input[15415]), .Z(o[5415]) );
  AND U5096 ( .A(p_input[5414]), .B(p_input[15414]), .Z(o[5414]) );
  AND U5097 ( .A(p_input[5413]), .B(p_input[15413]), .Z(o[5413]) );
  AND U5098 ( .A(p_input[5412]), .B(p_input[15412]), .Z(o[5412]) );
  AND U5099 ( .A(p_input[5411]), .B(p_input[15411]), .Z(o[5411]) );
  AND U5100 ( .A(p_input[5410]), .B(p_input[15410]), .Z(o[5410]) );
  AND U5101 ( .A(p_input[540]), .B(p_input[10540]), .Z(o[540]) );
  AND U5102 ( .A(p_input[5409]), .B(p_input[15409]), .Z(o[5409]) );
  AND U5103 ( .A(p_input[5408]), .B(p_input[15408]), .Z(o[5408]) );
  AND U5104 ( .A(p_input[5407]), .B(p_input[15407]), .Z(o[5407]) );
  AND U5105 ( .A(p_input[5406]), .B(p_input[15406]), .Z(o[5406]) );
  AND U5106 ( .A(p_input[5405]), .B(p_input[15405]), .Z(o[5405]) );
  AND U5107 ( .A(p_input[5404]), .B(p_input[15404]), .Z(o[5404]) );
  AND U5108 ( .A(p_input[5403]), .B(p_input[15403]), .Z(o[5403]) );
  AND U5109 ( .A(p_input[5402]), .B(p_input[15402]), .Z(o[5402]) );
  AND U5110 ( .A(p_input[5401]), .B(p_input[15401]), .Z(o[5401]) );
  AND U5111 ( .A(p_input[5400]), .B(p_input[15400]), .Z(o[5400]) );
  AND U5112 ( .A(p_input[53]), .B(p_input[10053]), .Z(o[53]) );
  AND U5113 ( .A(p_input[539]), .B(p_input[10539]), .Z(o[539]) );
  AND U5114 ( .A(p_input[5399]), .B(p_input[15399]), .Z(o[5399]) );
  AND U5115 ( .A(p_input[5398]), .B(p_input[15398]), .Z(o[5398]) );
  AND U5116 ( .A(p_input[5397]), .B(p_input[15397]), .Z(o[5397]) );
  AND U5117 ( .A(p_input[5396]), .B(p_input[15396]), .Z(o[5396]) );
  AND U5118 ( .A(p_input[5395]), .B(p_input[15395]), .Z(o[5395]) );
  AND U5119 ( .A(p_input[5394]), .B(p_input[15394]), .Z(o[5394]) );
  AND U5120 ( .A(p_input[5393]), .B(p_input[15393]), .Z(o[5393]) );
  AND U5121 ( .A(p_input[5392]), .B(p_input[15392]), .Z(o[5392]) );
  AND U5122 ( .A(p_input[5391]), .B(p_input[15391]), .Z(o[5391]) );
  AND U5123 ( .A(p_input[5390]), .B(p_input[15390]), .Z(o[5390]) );
  AND U5124 ( .A(p_input[538]), .B(p_input[10538]), .Z(o[538]) );
  AND U5125 ( .A(p_input[5389]), .B(p_input[15389]), .Z(o[5389]) );
  AND U5126 ( .A(p_input[5388]), .B(p_input[15388]), .Z(o[5388]) );
  AND U5127 ( .A(p_input[5387]), .B(p_input[15387]), .Z(o[5387]) );
  AND U5128 ( .A(p_input[5386]), .B(p_input[15386]), .Z(o[5386]) );
  AND U5129 ( .A(p_input[5385]), .B(p_input[15385]), .Z(o[5385]) );
  AND U5130 ( .A(p_input[5384]), .B(p_input[15384]), .Z(o[5384]) );
  AND U5131 ( .A(p_input[5383]), .B(p_input[15383]), .Z(o[5383]) );
  AND U5132 ( .A(p_input[5382]), .B(p_input[15382]), .Z(o[5382]) );
  AND U5133 ( .A(p_input[5381]), .B(p_input[15381]), .Z(o[5381]) );
  AND U5134 ( .A(p_input[5380]), .B(p_input[15380]), .Z(o[5380]) );
  AND U5135 ( .A(p_input[537]), .B(p_input[10537]), .Z(o[537]) );
  AND U5136 ( .A(p_input[5379]), .B(p_input[15379]), .Z(o[5379]) );
  AND U5137 ( .A(p_input[5378]), .B(p_input[15378]), .Z(o[5378]) );
  AND U5138 ( .A(p_input[5377]), .B(p_input[15377]), .Z(o[5377]) );
  AND U5139 ( .A(p_input[5376]), .B(p_input[15376]), .Z(o[5376]) );
  AND U5140 ( .A(p_input[5375]), .B(p_input[15375]), .Z(o[5375]) );
  AND U5141 ( .A(p_input[5374]), .B(p_input[15374]), .Z(o[5374]) );
  AND U5142 ( .A(p_input[5373]), .B(p_input[15373]), .Z(o[5373]) );
  AND U5143 ( .A(p_input[5372]), .B(p_input[15372]), .Z(o[5372]) );
  AND U5144 ( .A(p_input[5371]), .B(p_input[15371]), .Z(o[5371]) );
  AND U5145 ( .A(p_input[5370]), .B(p_input[15370]), .Z(o[5370]) );
  AND U5146 ( .A(p_input[536]), .B(p_input[10536]), .Z(o[536]) );
  AND U5147 ( .A(p_input[5369]), .B(p_input[15369]), .Z(o[5369]) );
  AND U5148 ( .A(p_input[5368]), .B(p_input[15368]), .Z(o[5368]) );
  AND U5149 ( .A(p_input[5367]), .B(p_input[15367]), .Z(o[5367]) );
  AND U5150 ( .A(p_input[5366]), .B(p_input[15366]), .Z(o[5366]) );
  AND U5151 ( .A(p_input[5365]), .B(p_input[15365]), .Z(o[5365]) );
  AND U5152 ( .A(p_input[5364]), .B(p_input[15364]), .Z(o[5364]) );
  AND U5153 ( .A(p_input[5363]), .B(p_input[15363]), .Z(o[5363]) );
  AND U5154 ( .A(p_input[5362]), .B(p_input[15362]), .Z(o[5362]) );
  AND U5155 ( .A(p_input[5361]), .B(p_input[15361]), .Z(o[5361]) );
  AND U5156 ( .A(p_input[5360]), .B(p_input[15360]), .Z(o[5360]) );
  AND U5157 ( .A(p_input[535]), .B(p_input[10535]), .Z(o[535]) );
  AND U5158 ( .A(p_input[5359]), .B(p_input[15359]), .Z(o[5359]) );
  AND U5159 ( .A(p_input[5358]), .B(p_input[15358]), .Z(o[5358]) );
  AND U5160 ( .A(p_input[5357]), .B(p_input[15357]), .Z(o[5357]) );
  AND U5161 ( .A(p_input[5356]), .B(p_input[15356]), .Z(o[5356]) );
  AND U5162 ( .A(p_input[5355]), .B(p_input[15355]), .Z(o[5355]) );
  AND U5163 ( .A(p_input[5354]), .B(p_input[15354]), .Z(o[5354]) );
  AND U5164 ( .A(p_input[5353]), .B(p_input[15353]), .Z(o[5353]) );
  AND U5165 ( .A(p_input[5352]), .B(p_input[15352]), .Z(o[5352]) );
  AND U5166 ( .A(p_input[5351]), .B(p_input[15351]), .Z(o[5351]) );
  AND U5167 ( .A(p_input[5350]), .B(p_input[15350]), .Z(o[5350]) );
  AND U5168 ( .A(p_input[534]), .B(p_input[10534]), .Z(o[534]) );
  AND U5169 ( .A(p_input[5349]), .B(p_input[15349]), .Z(o[5349]) );
  AND U5170 ( .A(p_input[5348]), .B(p_input[15348]), .Z(o[5348]) );
  AND U5171 ( .A(p_input[5347]), .B(p_input[15347]), .Z(o[5347]) );
  AND U5172 ( .A(p_input[5346]), .B(p_input[15346]), .Z(o[5346]) );
  AND U5173 ( .A(p_input[5345]), .B(p_input[15345]), .Z(o[5345]) );
  AND U5174 ( .A(p_input[5344]), .B(p_input[15344]), .Z(o[5344]) );
  AND U5175 ( .A(p_input[5343]), .B(p_input[15343]), .Z(o[5343]) );
  AND U5176 ( .A(p_input[5342]), .B(p_input[15342]), .Z(o[5342]) );
  AND U5177 ( .A(p_input[5341]), .B(p_input[15341]), .Z(o[5341]) );
  AND U5178 ( .A(p_input[5340]), .B(p_input[15340]), .Z(o[5340]) );
  AND U5179 ( .A(p_input[533]), .B(p_input[10533]), .Z(o[533]) );
  AND U5180 ( .A(p_input[5339]), .B(p_input[15339]), .Z(o[5339]) );
  AND U5181 ( .A(p_input[5338]), .B(p_input[15338]), .Z(o[5338]) );
  AND U5182 ( .A(p_input[5337]), .B(p_input[15337]), .Z(o[5337]) );
  AND U5183 ( .A(p_input[5336]), .B(p_input[15336]), .Z(o[5336]) );
  AND U5184 ( .A(p_input[5335]), .B(p_input[15335]), .Z(o[5335]) );
  AND U5185 ( .A(p_input[5334]), .B(p_input[15334]), .Z(o[5334]) );
  AND U5186 ( .A(p_input[5333]), .B(p_input[15333]), .Z(o[5333]) );
  AND U5187 ( .A(p_input[5332]), .B(p_input[15332]), .Z(o[5332]) );
  AND U5188 ( .A(p_input[5331]), .B(p_input[15331]), .Z(o[5331]) );
  AND U5189 ( .A(p_input[5330]), .B(p_input[15330]), .Z(o[5330]) );
  AND U5190 ( .A(p_input[532]), .B(p_input[10532]), .Z(o[532]) );
  AND U5191 ( .A(p_input[5329]), .B(p_input[15329]), .Z(o[5329]) );
  AND U5192 ( .A(p_input[5328]), .B(p_input[15328]), .Z(o[5328]) );
  AND U5193 ( .A(p_input[5327]), .B(p_input[15327]), .Z(o[5327]) );
  AND U5194 ( .A(p_input[5326]), .B(p_input[15326]), .Z(o[5326]) );
  AND U5195 ( .A(p_input[5325]), .B(p_input[15325]), .Z(o[5325]) );
  AND U5196 ( .A(p_input[5324]), .B(p_input[15324]), .Z(o[5324]) );
  AND U5197 ( .A(p_input[5323]), .B(p_input[15323]), .Z(o[5323]) );
  AND U5198 ( .A(p_input[5322]), .B(p_input[15322]), .Z(o[5322]) );
  AND U5199 ( .A(p_input[5321]), .B(p_input[15321]), .Z(o[5321]) );
  AND U5200 ( .A(p_input[5320]), .B(p_input[15320]), .Z(o[5320]) );
  AND U5201 ( .A(p_input[531]), .B(p_input[10531]), .Z(o[531]) );
  AND U5202 ( .A(p_input[5319]), .B(p_input[15319]), .Z(o[5319]) );
  AND U5203 ( .A(p_input[5318]), .B(p_input[15318]), .Z(o[5318]) );
  AND U5204 ( .A(p_input[5317]), .B(p_input[15317]), .Z(o[5317]) );
  AND U5205 ( .A(p_input[5316]), .B(p_input[15316]), .Z(o[5316]) );
  AND U5206 ( .A(p_input[5315]), .B(p_input[15315]), .Z(o[5315]) );
  AND U5207 ( .A(p_input[5314]), .B(p_input[15314]), .Z(o[5314]) );
  AND U5208 ( .A(p_input[5313]), .B(p_input[15313]), .Z(o[5313]) );
  AND U5209 ( .A(p_input[5312]), .B(p_input[15312]), .Z(o[5312]) );
  AND U5210 ( .A(p_input[5311]), .B(p_input[15311]), .Z(o[5311]) );
  AND U5211 ( .A(p_input[5310]), .B(p_input[15310]), .Z(o[5310]) );
  AND U5212 ( .A(p_input[530]), .B(p_input[10530]), .Z(o[530]) );
  AND U5213 ( .A(p_input[5309]), .B(p_input[15309]), .Z(o[5309]) );
  AND U5214 ( .A(p_input[5308]), .B(p_input[15308]), .Z(o[5308]) );
  AND U5215 ( .A(p_input[5307]), .B(p_input[15307]), .Z(o[5307]) );
  AND U5216 ( .A(p_input[5306]), .B(p_input[15306]), .Z(o[5306]) );
  AND U5217 ( .A(p_input[5305]), .B(p_input[15305]), .Z(o[5305]) );
  AND U5218 ( .A(p_input[5304]), .B(p_input[15304]), .Z(o[5304]) );
  AND U5219 ( .A(p_input[5303]), .B(p_input[15303]), .Z(o[5303]) );
  AND U5220 ( .A(p_input[5302]), .B(p_input[15302]), .Z(o[5302]) );
  AND U5221 ( .A(p_input[5301]), .B(p_input[15301]), .Z(o[5301]) );
  AND U5222 ( .A(p_input[5300]), .B(p_input[15300]), .Z(o[5300]) );
  AND U5223 ( .A(p_input[52]), .B(p_input[10052]), .Z(o[52]) );
  AND U5224 ( .A(p_input[529]), .B(p_input[10529]), .Z(o[529]) );
  AND U5225 ( .A(p_input[5299]), .B(p_input[15299]), .Z(o[5299]) );
  AND U5226 ( .A(p_input[5298]), .B(p_input[15298]), .Z(o[5298]) );
  AND U5227 ( .A(p_input[5297]), .B(p_input[15297]), .Z(o[5297]) );
  AND U5228 ( .A(p_input[5296]), .B(p_input[15296]), .Z(o[5296]) );
  AND U5229 ( .A(p_input[5295]), .B(p_input[15295]), .Z(o[5295]) );
  AND U5230 ( .A(p_input[5294]), .B(p_input[15294]), .Z(o[5294]) );
  AND U5231 ( .A(p_input[5293]), .B(p_input[15293]), .Z(o[5293]) );
  AND U5232 ( .A(p_input[5292]), .B(p_input[15292]), .Z(o[5292]) );
  AND U5233 ( .A(p_input[5291]), .B(p_input[15291]), .Z(o[5291]) );
  AND U5234 ( .A(p_input[5290]), .B(p_input[15290]), .Z(o[5290]) );
  AND U5235 ( .A(p_input[528]), .B(p_input[10528]), .Z(o[528]) );
  AND U5236 ( .A(p_input[5289]), .B(p_input[15289]), .Z(o[5289]) );
  AND U5237 ( .A(p_input[5288]), .B(p_input[15288]), .Z(o[5288]) );
  AND U5238 ( .A(p_input[5287]), .B(p_input[15287]), .Z(o[5287]) );
  AND U5239 ( .A(p_input[5286]), .B(p_input[15286]), .Z(o[5286]) );
  AND U5240 ( .A(p_input[5285]), .B(p_input[15285]), .Z(o[5285]) );
  AND U5241 ( .A(p_input[5284]), .B(p_input[15284]), .Z(o[5284]) );
  AND U5242 ( .A(p_input[5283]), .B(p_input[15283]), .Z(o[5283]) );
  AND U5243 ( .A(p_input[5282]), .B(p_input[15282]), .Z(o[5282]) );
  AND U5244 ( .A(p_input[5281]), .B(p_input[15281]), .Z(o[5281]) );
  AND U5245 ( .A(p_input[5280]), .B(p_input[15280]), .Z(o[5280]) );
  AND U5246 ( .A(p_input[527]), .B(p_input[10527]), .Z(o[527]) );
  AND U5247 ( .A(p_input[5279]), .B(p_input[15279]), .Z(o[5279]) );
  AND U5248 ( .A(p_input[5278]), .B(p_input[15278]), .Z(o[5278]) );
  AND U5249 ( .A(p_input[5277]), .B(p_input[15277]), .Z(o[5277]) );
  AND U5250 ( .A(p_input[5276]), .B(p_input[15276]), .Z(o[5276]) );
  AND U5251 ( .A(p_input[5275]), .B(p_input[15275]), .Z(o[5275]) );
  AND U5252 ( .A(p_input[5274]), .B(p_input[15274]), .Z(o[5274]) );
  AND U5253 ( .A(p_input[5273]), .B(p_input[15273]), .Z(o[5273]) );
  AND U5254 ( .A(p_input[5272]), .B(p_input[15272]), .Z(o[5272]) );
  AND U5255 ( .A(p_input[5271]), .B(p_input[15271]), .Z(o[5271]) );
  AND U5256 ( .A(p_input[5270]), .B(p_input[15270]), .Z(o[5270]) );
  AND U5257 ( .A(p_input[526]), .B(p_input[10526]), .Z(o[526]) );
  AND U5258 ( .A(p_input[5269]), .B(p_input[15269]), .Z(o[5269]) );
  AND U5259 ( .A(p_input[5268]), .B(p_input[15268]), .Z(o[5268]) );
  AND U5260 ( .A(p_input[5267]), .B(p_input[15267]), .Z(o[5267]) );
  AND U5261 ( .A(p_input[5266]), .B(p_input[15266]), .Z(o[5266]) );
  AND U5262 ( .A(p_input[5265]), .B(p_input[15265]), .Z(o[5265]) );
  AND U5263 ( .A(p_input[5264]), .B(p_input[15264]), .Z(o[5264]) );
  AND U5264 ( .A(p_input[5263]), .B(p_input[15263]), .Z(o[5263]) );
  AND U5265 ( .A(p_input[5262]), .B(p_input[15262]), .Z(o[5262]) );
  AND U5266 ( .A(p_input[5261]), .B(p_input[15261]), .Z(o[5261]) );
  AND U5267 ( .A(p_input[5260]), .B(p_input[15260]), .Z(o[5260]) );
  AND U5268 ( .A(p_input[525]), .B(p_input[10525]), .Z(o[525]) );
  AND U5269 ( .A(p_input[5259]), .B(p_input[15259]), .Z(o[5259]) );
  AND U5270 ( .A(p_input[5258]), .B(p_input[15258]), .Z(o[5258]) );
  AND U5271 ( .A(p_input[5257]), .B(p_input[15257]), .Z(o[5257]) );
  AND U5272 ( .A(p_input[5256]), .B(p_input[15256]), .Z(o[5256]) );
  AND U5273 ( .A(p_input[5255]), .B(p_input[15255]), .Z(o[5255]) );
  AND U5274 ( .A(p_input[5254]), .B(p_input[15254]), .Z(o[5254]) );
  AND U5275 ( .A(p_input[5253]), .B(p_input[15253]), .Z(o[5253]) );
  AND U5276 ( .A(p_input[5252]), .B(p_input[15252]), .Z(o[5252]) );
  AND U5277 ( .A(p_input[5251]), .B(p_input[15251]), .Z(o[5251]) );
  AND U5278 ( .A(p_input[5250]), .B(p_input[15250]), .Z(o[5250]) );
  AND U5279 ( .A(p_input[524]), .B(p_input[10524]), .Z(o[524]) );
  AND U5280 ( .A(p_input[5249]), .B(p_input[15249]), .Z(o[5249]) );
  AND U5281 ( .A(p_input[5248]), .B(p_input[15248]), .Z(o[5248]) );
  AND U5282 ( .A(p_input[5247]), .B(p_input[15247]), .Z(o[5247]) );
  AND U5283 ( .A(p_input[5246]), .B(p_input[15246]), .Z(o[5246]) );
  AND U5284 ( .A(p_input[5245]), .B(p_input[15245]), .Z(o[5245]) );
  AND U5285 ( .A(p_input[5244]), .B(p_input[15244]), .Z(o[5244]) );
  AND U5286 ( .A(p_input[5243]), .B(p_input[15243]), .Z(o[5243]) );
  AND U5287 ( .A(p_input[5242]), .B(p_input[15242]), .Z(o[5242]) );
  AND U5288 ( .A(p_input[5241]), .B(p_input[15241]), .Z(o[5241]) );
  AND U5289 ( .A(p_input[5240]), .B(p_input[15240]), .Z(o[5240]) );
  AND U5290 ( .A(p_input[523]), .B(p_input[10523]), .Z(o[523]) );
  AND U5291 ( .A(p_input[5239]), .B(p_input[15239]), .Z(o[5239]) );
  AND U5292 ( .A(p_input[5238]), .B(p_input[15238]), .Z(o[5238]) );
  AND U5293 ( .A(p_input[5237]), .B(p_input[15237]), .Z(o[5237]) );
  AND U5294 ( .A(p_input[5236]), .B(p_input[15236]), .Z(o[5236]) );
  AND U5295 ( .A(p_input[5235]), .B(p_input[15235]), .Z(o[5235]) );
  AND U5296 ( .A(p_input[5234]), .B(p_input[15234]), .Z(o[5234]) );
  AND U5297 ( .A(p_input[5233]), .B(p_input[15233]), .Z(o[5233]) );
  AND U5298 ( .A(p_input[5232]), .B(p_input[15232]), .Z(o[5232]) );
  AND U5299 ( .A(p_input[5231]), .B(p_input[15231]), .Z(o[5231]) );
  AND U5300 ( .A(p_input[5230]), .B(p_input[15230]), .Z(o[5230]) );
  AND U5301 ( .A(p_input[522]), .B(p_input[10522]), .Z(o[522]) );
  AND U5302 ( .A(p_input[5229]), .B(p_input[15229]), .Z(o[5229]) );
  AND U5303 ( .A(p_input[5228]), .B(p_input[15228]), .Z(o[5228]) );
  AND U5304 ( .A(p_input[5227]), .B(p_input[15227]), .Z(o[5227]) );
  AND U5305 ( .A(p_input[5226]), .B(p_input[15226]), .Z(o[5226]) );
  AND U5306 ( .A(p_input[5225]), .B(p_input[15225]), .Z(o[5225]) );
  AND U5307 ( .A(p_input[5224]), .B(p_input[15224]), .Z(o[5224]) );
  AND U5308 ( .A(p_input[5223]), .B(p_input[15223]), .Z(o[5223]) );
  AND U5309 ( .A(p_input[5222]), .B(p_input[15222]), .Z(o[5222]) );
  AND U5310 ( .A(p_input[5221]), .B(p_input[15221]), .Z(o[5221]) );
  AND U5311 ( .A(p_input[5220]), .B(p_input[15220]), .Z(o[5220]) );
  AND U5312 ( .A(p_input[521]), .B(p_input[10521]), .Z(o[521]) );
  AND U5313 ( .A(p_input[5219]), .B(p_input[15219]), .Z(o[5219]) );
  AND U5314 ( .A(p_input[5218]), .B(p_input[15218]), .Z(o[5218]) );
  AND U5315 ( .A(p_input[5217]), .B(p_input[15217]), .Z(o[5217]) );
  AND U5316 ( .A(p_input[5216]), .B(p_input[15216]), .Z(o[5216]) );
  AND U5317 ( .A(p_input[5215]), .B(p_input[15215]), .Z(o[5215]) );
  AND U5318 ( .A(p_input[5214]), .B(p_input[15214]), .Z(o[5214]) );
  AND U5319 ( .A(p_input[5213]), .B(p_input[15213]), .Z(o[5213]) );
  AND U5320 ( .A(p_input[5212]), .B(p_input[15212]), .Z(o[5212]) );
  AND U5321 ( .A(p_input[5211]), .B(p_input[15211]), .Z(o[5211]) );
  AND U5322 ( .A(p_input[5210]), .B(p_input[15210]), .Z(o[5210]) );
  AND U5323 ( .A(p_input[520]), .B(p_input[10520]), .Z(o[520]) );
  AND U5324 ( .A(p_input[5209]), .B(p_input[15209]), .Z(o[5209]) );
  AND U5325 ( .A(p_input[5208]), .B(p_input[15208]), .Z(o[5208]) );
  AND U5326 ( .A(p_input[5207]), .B(p_input[15207]), .Z(o[5207]) );
  AND U5327 ( .A(p_input[5206]), .B(p_input[15206]), .Z(o[5206]) );
  AND U5328 ( .A(p_input[5205]), .B(p_input[15205]), .Z(o[5205]) );
  AND U5329 ( .A(p_input[5204]), .B(p_input[15204]), .Z(o[5204]) );
  AND U5330 ( .A(p_input[5203]), .B(p_input[15203]), .Z(o[5203]) );
  AND U5331 ( .A(p_input[5202]), .B(p_input[15202]), .Z(o[5202]) );
  AND U5332 ( .A(p_input[5201]), .B(p_input[15201]), .Z(o[5201]) );
  AND U5333 ( .A(p_input[5200]), .B(p_input[15200]), .Z(o[5200]) );
  AND U5334 ( .A(p_input[51]), .B(p_input[10051]), .Z(o[51]) );
  AND U5335 ( .A(p_input[519]), .B(p_input[10519]), .Z(o[519]) );
  AND U5336 ( .A(p_input[5199]), .B(p_input[15199]), .Z(o[5199]) );
  AND U5337 ( .A(p_input[5198]), .B(p_input[15198]), .Z(o[5198]) );
  AND U5338 ( .A(p_input[5197]), .B(p_input[15197]), .Z(o[5197]) );
  AND U5339 ( .A(p_input[5196]), .B(p_input[15196]), .Z(o[5196]) );
  AND U5340 ( .A(p_input[5195]), .B(p_input[15195]), .Z(o[5195]) );
  AND U5341 ( .A(p_input[5194]), .B(p_input[15194]), .Z(o[5194]) );
  AND U5342 ( .A(p_input[5193]), .B(p_input[15193]), .Z(o[5193]) );
  AND U5343 ( .A(p_input[5192]), .B(p_input[15192]), .Z(o[5192]) );
  AND U5344 ( .A(p_input[5191]), .B(p_input[15191]), .Z(o[5191]) );
  AND U5345 ( .A(p_input[5190]), .B(p_input[15190]), .Z(o[5190]) );
  AND U5346 ( .A(p_input[518]), .B(p_input[10518]), .Z(o[518]) );
  AND U5347 ( .A(p_input[5189]), .B(p_input[15189]), .Z(o[5189]) );
  AND U5348 ( .A(p_input[5188]), .B(p_input[15188]), .Z(o[5188]) );
  AND U5349 ( .A(p_input[5187]), .B(p_input[15187]), .Z(o[5187]) );
  AND U5350 ( .A(p_input[5186]), .B(p_input[15186]), .Z(o[5186]) );
  AND U5351 ( .A(p_input[5185]), .B(p_input[15185]), .Z(o[5185]) );
  AND U5352 ( .A(p_input[5184]), .B(p_input[15184]), .Z(o[5184]) );
  AND U5353 ( .A(p_input[5183]), .B(p_input[15183]), .Z(o[5183]) );
  AND U5354 ( .A(p_input[5182]), .B(p_input[15182]), .Z(o[5182]) );
  AND U5355 ( .A(p_input[5181]), .B(p_input[15181]), .Z(o[5181]) );
  AND U5356 ( .A(p_input[5180]), .B(p_input[15180]), .Z(o[5180]) );
  AND U5357 ( .A(p_input[517]), .B(p_input[10517]), .Z(o[517]) );
  AND U5358 ( .A(p_input[5179]), .B(p_input[15179]), .Z(o[5179]) );
  AND U5359 ( .A(p_input[5178]), .B(p_input[15178]), .Z(o[5178]) );
  AND U5360 ( .A(p_input[5177]), .B(p_input[15177]), .Z(o[5177]) );
  AND U5361 ( .A(p_input[5176]), .B(p_input[15176]), .Z(o[5176]) );
  AND U5362 ( .A(p_input[5175]), .B(p_input[15175]), .Z(o[5175]) );
  AND U5363 ( .A(p_input[5174]), .B(p_input[15174]), .Z(o[5174]) );
  AND U5364 ( .A(p_input[5173]), .B(p_input[15173]), .Z(o[5173]) );
  AND U5365 ( .A(p_input[5172]), .B(p_input[15172]), .Z(o[5172]) );
  AND U5366 ( .A(p_input[5171]), .B(p_input[15171]), .Z(o[5171]) );
  AND U5367 ( .A(p_input[5170]), .B(p_input[15170]), .Z(o[5170]) );
  AND U5368 ( .A(p_input[516]), .B(p_input[10516]), .Z(o[516]) );
  AND U5369 ( .A(p_input[5169]), .B(p_input[15169]), .Z(o[5169]) );
  AND U5370 ( .A(p_input[5168]), .B(p_input[15168]), .Z(o[5168]) );
  AND U5371 ( .A(p_input[5167]), .B(p_input[15167]), .Z(o[5167]) );
  AND U5372 ( .A(p_input[5166]), .B(p_input[15166]), .Z(o[5166]) );
  AND U5373 ( .A(p_input[5165]), .B(p_input[15165]), .Z(o[5165]) );
  AND U5374 ( .A(p_input[5164]), .B(p_input[15164]), .Z(o[5164]) );
  AND U5375 ( .A(p_input[5163]), .B(p_input[15163]), .Z(o[5163]) );
  AND U5376 ( .A(p_input[5162]), .B(p_input[15162]), .Z(o[5162]) );
  AND U5377 ( .A(p_input[5161]), .B(p_input[15161]), .Z(o[5161]) );
  AND U5378 ( .A(p_input[5160]), .B(p_input[15160]), .Z(o[5160]) );
  AND U5379 ( .A(p_input[515]), .B(p_input[10515]), .Z(o[515]) );
  AND U5380 ( .A(p_input[5159]), .B(p_input[15159]), .Z(o[5159]) );
  AND U5381 ( .A(p_input[5158]), .B(p_input[15158]), .Z(o[5158]) );
  AND U5382 ( .A(p_input[5157]), .B(p_input[15157]), .Z(o[5157]) );
  AND U5383 ( .A(p_input[5156]), .B(p_input[15156]), .Z(o[5156]) );
  AND U5384 ( .A(p_input[5155]), .B(p_input[15155]), .Z(o[5155]) );
  AND U5385 ( .A(p_input[5154]), .B(p_input[15154]), .Z(o[5154]) );
  AND U5386 ( .A(p_input[5153]), .B(p_input[15153]), .Z(o[5153]) );
  AND U5387 ( .A(p_input[5152]), .B(p_input[15152]), .Z(o[5152]) );
  AND U5388 ( .A(p_input[5151]), .B(p_input[15151]), .Z(o[5151]) );
  AND U5389 ( .A(p_input[5150]), .B(p_input[15150]), .Z(o[5150]) );
  AND U5390 ( .A(p_input[514]), .B(p_input[10514]), .Z(o[514]) );
  AND U5391 ( .A(p_input[5149]), .B(p_input[15149]), .Z(o[5149]) );
  AND U5392 ( .A(p_input[5148]), .B(p_input[15148]), .Z(o[5148]) );
  AND U5393 ( .A(p_input[5147]), .B(p_input[15147]), .Z(o[5147]) );
  AND U5394 ( .A(p_input[5146]), .B(p_input[15146]), .Z(o[5146]) );
  AND U5395 ( .A(p_input[5145]), .B(p_input[15145]), .Z(o[5145]) );
  AND U5396 ( .A(p_input[5144]), .B(p_input[15144]), .Z(o[5144]) );
  AND U5397 ( .A(p_input[5143]), .B(p_input[15143]), .Z(o[5143]) );
  AND U5398 ( .A(p_input[5142]), .B(p_input[15142]), .Z(o[5142]) );
  AND U5399 ( .A(p_input[5141]), .B(p_input[15141]), .Z(o[5141]) );
  AND U5400 ( .A(p_input[5140]), .B(p_input[15140]), .Z(o[5140]) );
  AND U5401 ( .A(p_input[513]), .B(p_input[10513]), .Z(o[513]) );
  AND U5402 ( .A(p_input[5139]), .B(p_input[15139]), .Z(o[5139]) );
  AND U5403 ( .A(p_input[5138]), .B(p_input[15138]), .Z(o[5138]) );
  AND U5404 ( .A(p_input[5137]), .B(p_input[15137]), .Z(o[5137]) );
  AND U5405 ( .A(p_input[5136]), .B(p_input[15136]), .Z(o[5136]) );
  AND U5406 ( .A(p_input[5135]), .B(p_input[15135]), .Z(o[5135]) );
  AND U5407 ( .A(p_input[5134]), .B(p_input[15134]), .Z(o[5134]) );
  AND U5408 ( .A(p_input[5133]), .B(p_input[15133]), .Z(o[5133]) );
  AND U5409 ( .A(p_input[5132]), .B(p_input[15132]), .Z(o[5132]) );
  AND U5410 ( .A(p_input[5131]), .B(p_input[15131]), .Z(o[5131]) );
  AND U5411 ( .A(p_input[5130]), .B(p_input[15130]), .Z(o[5130]) );
  AND U5412 ( .A(p_input[512]), .B(p_input[10512]), .Z(o[512]) );
  AND U5413 ( .A(p_input[5129]), .B(p_input[15129]), .Z(o[5129]) );
  AND U5414 ( .A(p_input[5128]), .B(p_input[15128]), .Z(o[5128]) );
  AND U5415 ( .A(p_input[5127]), .B(p_input[15127]), .Z(o[5127]) );
  AND U5416 ( .A(p_input[5126]), .B(p_input[15126]), .Z(o[5126]) );
  AND U5417 ( .A(p_input[5125]), .B(p_input[15125]), .Z(o[5125]) );
  AND U5418 ( .A(p_input[5124]), .B(p_input[15124]), .Z(o[5124]) );
  AND U5419 ( .A(p_input[5123]), .B(p_input[15123]), .Z(o[5123]) );
  AND U5420 ( .A(p_input[5122]), .B(p_input[15122]), .Z(o[5122]) );
  AND U5421 ( .A(p_input[5121]), .B(p_input[15121]), .Z(o[5121]) );
  AND U5422 ( .A(p_input[5120]), .B(p_input[15120]), .Z(o[5120]) );
  AND U5423 ( .A(p_input[511]), .B(p_input[10511]), .Z(o[511]) );
  AND U5424 ( .A(p_input[5119]), .B(p_input[15119]), .Z(o[5119]) );
  AND U5425 ( .A(p_input[5118]), .B(p_input[15118]), .Z(o[5118]) );
  AND U5426 ( .A(p_input[5117]), .B(p_input[15117]), .Z(o[5117]) );
  AND U5427 ( .A(p_input[5116]), .B(p_input[15116]), .Z(o[5116]) );
  AND U5428 ( .A(p_input[5115]), .B(p_input[15115]), .Z(o[5115]) );
  AND U5429 ( .A(p_input[5114]), .B(p_input[15114]), .Z(o[5114]) );
  AND U5430 ( .A(p_input[5113]), .B(p_input[15113]), .Z(o[5113]) );
  AND U5431 ( .A(p_input[5112]), .B(p_input[15112]), .Z(o[5112]) );
  AND U5432 ( .A(p_input[5111]), .B(p_input[15111]), .Z(o[5111]) );
  AND U5433 ( .A(p_input[5110]), .B(p_input[15110]), .Z(o[5110]) );
  AND U5434 ( .A(p_input[510]), .B(p_input[10510]), .Z(o[510]) );
  AND U5435 ( .A(p_input[5109]), .B(p_input[15109]), .Z(o[5109]) );
  AND U5436 ( .A(p_input[5108]), .B(p_input[15108]), .Z(o[5108]) );
  AND U5437 ( .A(p_input[5107]), .B(p_input[15107]), .Z(o[5107]) );
  AND U5438 ( .A(p_input[5106]), .B(p_input[15106]), .Z(o[5106]) );
  AND U5439 ( .A(p_input[5105]), .B(p_input[15105]), .Z(o[5105]) );
  AND U5440 ( .A(p_input[5104]), .B(p_input[15104]), .Z(o[5104]) );
  AND U5441 ( .A(p_input[5103]), .B(p_input[15103]), .Z(o[5103]) );
  AND U5442 ( .A(p_input[5102]), .B(p_input[15102]), .Z(o[5102]) );
  AND U5443 ( .A(p_input[5101]), .B(p_input[15101]), .Z(o[5101]) );
  AND U5444 ( .A(p_input[5100]), .B(p_input[15100]), .Z(o[5100]) );
  AND U5445 ( .A(p_input[50]), .B(p_input[10050]), .Z(o[50]) );
  AND U5446 ( .A(p_input[509]), .B(p_input[10509]), .Z(o[509]) );
  AND U5447 ( .A(p_input[5099]), .B(p_input[15099]), .Z(o[5099]) );
  AND U5448 ( .A(p_input[5098]), .B(p_input[15098]), .Z(o[5098]) );
  AND U5449 ( .A(p_input[5097]), .B(p_input[15097]), .Z(o[5097]) );
  AND U5450 ( .A(p_input[5096]), .B(p_input[15096]), .Z(o[5096]) );
  AND U5451 ( .A(p_input[5095]), .B(p_input[15095]), .Z(o[5095]) );
  AND U5452 ( .A(p_input[5094]), .B(p_input[15094]), .Z(o[5094]) );
  AND U5453 ( .A(p_input[5093]), .B(p_input[15093]), .Z(o[5093]) );
  AND U5454 ( .A(p_input[5092]), .B(p_input[15092]), .Z(o[5092]) );
  AND U5455 ( .A(p_input[5091]), .B(p_input[15091]), .Z(o[5091]) );
  AND U5456 ( .A(p_input[5090]), .B(p_input[15090]), .Z(o[5090]) );
  AND U5457 ( .A(p_input[508]), .B(p_input[10508]), .Z(o[508]) );
  AND U5458 ( .A(p_input[5089]), .B(p_input[15089]), .Z(o[5089]) );
  AND U5459 ( .A(p_input[5088]), .B(p_input[15088]), .Z(o[5088]) );
  AND U5460 ( .A(p_input[5087]), .B(p_input[15087]), .Z(o[5087]) );
  AND U5461 ( .A(p_input[5086]), .B(p_input[15086]), .Z(o[5086]) );
  AND U5462 ( .A(p_input[5085]), .B(p_input[15085]), .Z(o[5085]) );
  AND U5463 ( .A(p_input[5084]), .B(p_input[15084]), .Z(o[5084]) );
  AND U5464 ( .A(p_input[5083]), .B(p_input[15083]), .Z(o[5083]) );
  AND U5465 ( .A(p_input[5082]), .B(p_input[15082]), .Z(o[5082]) );
  AND U5466 ( .A(p_input[5081]), .B(p_input[15081]), .Z(o[5081]) );
  AND U5467 ( .A(p_input[5080]), .B(p_input[15080]), .Z(o[5080]) );
  AND U5468 ( .A(p_input[507]), .B(p_input[10507]), .Z(o[507]) );
  AND U5469 ( .A(p_input[5079]), .B(p_input[15079]), .Z(o[5079]) );
  AND U5470 ( .A(p_input[5078]), .B(p_input[15078]), .Z(o[5078]) );
  AND U5471 ( .A(p_input[5077]), .B(p_input[15077]), .Z(o[5077]) );
  AND U5472 ( .A(p_input[5076]), .B(p_input[15076]), .Z(o[5076]) );
  AND U5473 ( .A(p_input[5075]), .B(p_input[15075]), .Z(o[5075]) );
  AND U5474 ( .A(p_input[5074]), .B(p_input[15074]), .Z(o[5074]) );
  AND U5475 ( .A(p_input[5073]), .B(p_input[15073]), .Z(o[5073]) );
  AND U5476 ( .A(p_input[5072]), .B(p_input[15072]), .Z(o[5072]) );
  AND U5477 ( .A(p_input[5071]), .B(p_input[15071]), .Z(o[5071]) );
  AND U5478 ( .A(p_input[5070]), .B(p_input[15070]), .Z(o[5070]) );
  AND U5479 ( .A(p_input[506]), .B(p_input[10506]), .Z(o[506]) );
  AND U5480 ( .A(p_input[5069]), .B(p_input[15069]), .Z(o[5069]) );
  AND U5481 ( .A(p_input[5068]), .B(p_input[15068]), .Z(o[5068]) );
  AND U5482 ( .A(p_input[5067]), .B(p_input[15067]), .Z(o[5067]) );
  AND U5483 ( .A(p_input[5066]), .B(p_input[15066]), .Z(o[5066]) );
  AND U5484 ( .A(p_input[5065]), .B(p_input[15065]), .Z(o[5065]) );
  AND U5485 ( .A(p_input[5064]), .B(p_input[15064]), .Z(o[5064]) );
  AND U5486 ( .A(p_input[5063]), .B(p_input[15063]), .Z(o[5063]) );
  AND U5487 ( .A(p_input[5062]), .B(p_input[15062]), .Z(o[5062]) );
  AND U5488 ( .A(p_input[5061]), .B(p_input[15061]), .Z(o[5061]) );
  AND U5489 ( .A(p_input[5060]), .B(p_input[15060]), .Z(o[5060]) );
  AND U5490 ( .A(p_input[505]), .B(p_input[10505]), .Z(o[505]) );
  AND U5491 ( .A(p_input[5059]), .B(p_input[15059]), .Z(o[5059]) );
  AND U5492 ( .A(p_input[5058]), .B(p_input[15058]), .Z(o[5058]) );
  AND U5493 ( .A(p_input[5057]), .B(p_input[15057]), .Z(o[5057]) );
  AND U5494 ( .A(p_input[5056]), .B(p_input[15056]), .Z(o[5056]) );
  AND U5495 ( .A(p_input[5055]), .B(p_input[15055]), .Z(o[5055]) );
  AND U5496 ( .A(p_input[5054]), .B(p_input[15054]), .Z(o[5054]) );
  AND U5497 ( .A(p_input[5053]), .B(p_input[15053]), .Z(o[5053]) );
  AND U5498 ( .A(p_input[5052]), .B(p_input[15052]), .Z(o[5052]) );
  AND U5499 ( .A(p_input[5051]), .B(p_input[15051]), .Z(o[5051]) );
  AND U5500 ( .A(p_input[5050]), .B(p_input[15050]), .Z(o[5050]) );
  AND U5501 ( .A(p_input[504]), .B(p_input[10504]), .Z(o[504]) );
  AND U5502 ( .A(p_input[5049]), .B(p_input[15049]), .Z(o[5049]) );
  AND U5503 ( .A(p_input[5048]), .B(p_input[15048]), .Z(o[5048]) );
  AND U5504 ( .A(p_input[5047]), .B(p_input[15047]), .Z(o[5047]) );
  AND U5505 ( .A(p_input[5046]), .B(p_input[15046]), .Z(o[5046]) );
  AND U5506 ( .A(p_input[5045]), .B(p_input[15045]), .Z(o[5045]) );
  AND U5507 ( .A(p_input[5044]), .B(p_input[15044]), .Z(o[5044]) );
  AND U5508 ( .A(p_input[5043]), .B(p_input[15043]), .Z(o[5043]) );
  AND U5509 ( .A(p_input[5042]), .B(p_input[15042]), .Z(o[5042]) );
  AND U5510 ( .A(p_input[5041]), .B(p_input[15041]), .Z(o[5041]) );
  AND U5511 ( .A(p_input[5040]), .B(p_input[15040]), .Z(o[5040]) );
  AND U5512 ( .A(p_input[503]), .B(p_input[10503]), .Z(o[503]) );
  AND U5513 ( .A(p_input[5039]), .B(p_input[15039]), .Z(o[5039]) );
  AND U5514 ( .A(p_input[5038]), .B(p_input[15038]), .Z(o[5038]) );
  AND U5515 ( .A(p_input[5037]), .B(p_input[15037]), .Z(o[5037]) );
  AND U5516 ( .A(p_input[5036]), .B(p_input[15036]), .Z(o[5036]) );
  AND U5517 ( .A(p_input[5035]), .B(p_input[15035]), .Z(o[5035]) );
  AND U5518 ( .A(p_input[5034]), .B(p_input[15034]), .Z(o[5034]) );
  AND U5519 ( .A(p_input[5033]), .B(p_input[15033]), .Z(o[5033]) );
  AND U5520 ( .A(p_input[5032]), .B(p_input[15032]), .Z(o[5032]) );
  AND U5521 ( .A(p_input[5031]), .B(p_input[15031]), .Z(o[5031]) );
  AND U5522 ( .A(p_input[5030]), .B(p_input[15030]), .Z(o[5030]) );
  AND U5523 ( .A(p_input[502]), .B(p_input[10502]), .Z(o[502]) );
  AND U5524 ( .A(p_input[5029]), .B(p_input[15029]), .Z(o[5029]) );
  AND U5525 ( .A(p_input[5028]), .B(p_input[15028]), .Z(o[5028]) );
  AND U5526 ( .A(p_input[5027]), .B(p_input[15027]), .Z(o[5027]) );
  AND U5527 ( .A(p_input[5026]), .B(p_input[15026]), .Z(o[5026]) );
  AND U5528 ( .A(p_input[5025]), .B(p_input[15025]), .Z(o[5025]) );
  AND U5529 ( .A(p_input[5024]), .B(p_input[15024]), .Z(o[5024]) );
  AND U5530 ( .A(p_input[5023]), .B(p_input[15023]), .Z(o[5023]) );
  AND U5531 ( .A(p_input[5022]), .B(p_input[15022]), .Z(o[5022]) );
  AND U5532 ( .A(p_input[5021]), .B(p_input[15021]), .Z(o[5021]) );
  AND U5533 ( .A(p_input[5020]), .B(p_input[15020]), .Z(o[5020]) );
  AND U5534 ( .A(p_input[501]), .B(p_input[10501]), .Z(o[501]) );
  AND U5535 ( .A(p_input[5019]), .B(p_input[15019]), .Z(o[5019]) );
  AND U5536 ( .A(p_input[5018]), .B(p_input[15018]), .Z(o[5018]) );
  AND U5537 ( .A(p_input[5017]), .B(p_input[15017]), .Z(o[5017]) );
  AND U5538 ( .A(p_input[5016]), .B(p_input[15016]), .Z(o[5016]) );
  AND U5539 ( .A(p_input[5015]), .B(p_input[15015]), .Z(o[5015]) );
  AND U5540 ( .A(p_input[5014]), .B(p_input[15014]), .Z(o[5014]) );
  AND U5541 ( .A(p_input[5013]), .B(p_input[15013]), .Z(o[5013]) );
  AND U5542 ( .A(p_input[5012]), .B(p_input[15012]), .Z(o[5012]) );
  AND U5543 ( .A(p_input[5011]), .B(p_input[15011]), .Z(o[5011]) );
  AND U5544 ( .A(p_input[5010]), .B(p_input[15010]), .Z(o[5010]) );
  AND U5545 ( .A(p_input[500]), .B(p_input[10500]), .Z(o[500]) );
  AND U5546 ( .A(p_input[5009]), .B(p_input[15009]), .Z(o[5009]) );
  AND U5547 ( .A(p_input[5008]), .B(p_input[15008]), .Z(o[5008]) );
  AND U5548 ( .A(p_input[5007]), .B(p_input[15007]), .Z(o[5007]) );
  AND U5549 ( .A(p_input[5006]), .B(p_input[15006]), .Z(o[5006]) );
  AND U5550 ( .A(p_input[5005]), .B(p_input[15005]), .Z(o[5005]) );
  AND U5551 ( .A(p_input[5004]), .B(p_input[15004]), .Z(o[5004]) );
  AND U5552 ( .A(p_input[5003]), .B(p_input[15003]), .Z(o[5003]) );
  AND U5553 ( .A(p_input[5002]), .B(p_input[15002]), .Z(o[5002]) );
  AND U5554 ( .A(p_input[5001]), .B(p_input[15001]), .Z(o[5001]) );
  AND U5555 ( .A(p_input[5000]), .B(p_input[15000]), .Z(o[5000]) );
  AND U5556 ( .A(p_input[4]), .B(p_input[10004]), .Z(o[4]) );
  AND U5557 ( .A(p_input[49]), .B(p_input[10049]), .Z(o[49]) );
  AND U5558 ( .A(p_input[499]), .B(p_input[10499]), .Z(o[499]) );
  AND U5559 ( .A(p_input[4999]), .B(p_input[14999]), .Z(o[4999]) );
  AND U5560 ( .A(p_input[4998]), .B(p_input[14998]), .Z(o[4998]) );
  AND U5561 ( .A(p_input[4997]), .B(p_input[14997]), .Z(o[4997]) );
  AND U5562 ( .A(p_input[4996]), .B(p_input[14996]), .Z(o[4996]) );
  AND U5563 ( .A(p_input[4995]), .B(p_input[14995]), .Z(o[4995]) );
  AND U5564 ( .A(p_input[4994]), .B(p_input[14994]), .Z(o[4994]) );
  AND U5565 ( .A(p_input[4993]), .B(p_input[14993]), .Z(o[4993]) );
  AND U5566 ( .A(p_input[4992]), .B(p_input[14992]), .Z(o[4992]) );
  AND U5567 ( .A(p_input[4991]), .B(p_input[14991]), .Z(o[4991]) );
  AND U5568 ( .A(p_input[4990]), .B(p_input[14990]), .Z(o[4990]) );
  AND U5569 ( .A(p_input[498]), .B(p_input[10498]), .Z(o[498]) );
  AND U5570 ( .A(p_input[4989]), .B(p_input[14989]), .Z(o[4989]) );
  AND U5571 ( .A(p_input[4988]), .B(p_input[14988]), .Z(o[4988]) );
  AND U5572 ( .A(p_input[4987]), .B(p_input[14987]), .Z(o[4987]) );
  AND U5573 ( .A(p_input[4986]), .B(p_input[14986]), .Z(o[4986]) );
  AND U5574 ( .A(p_input[4985]), .B(p_input[14985]), .Z(o[4985]) );
  AND U5575 ( .A(p_input[4984]), .B(p_input[14984]), .Z(o[4984]) );
  AND U5576 ( .A(p_input[4983]), .B(p_input[14983]), .Z(o[4983]) );
  AND U5577 ( .A(p_input[4982]), .B(p_input[14982]), .Z(o[4982]) );
  AND U5578 ( .A(p_input[4981]), .B(p_input[14981]), .Z(o[4981]) );
  AND U5579 ( .A(p_input[4980]), .B(p_input[14980]), .Z(o[4980]) );
  AND U5580 ( .A(p_input[497]), .B(p_input[10497]), .Z(o[497]) );
  AND U5581 ( .A(p_input[4979]), .B(p_input[14979]), .Z(o[4979]) );
  AND U5582 ( .A(p_input[4978]), .B(p_input[14978]), .Z(o[4978]) );
  AND U5583 ( .A(p_input[4977]), .B(p_input[14977]), .Z(o[4977]) );
  AND U5584 ( .A(p_input[4976]), .B(p_input[14976]), .Z(o[4976]) );
  AND U5585 ( .A(p_input[4975]), .B(p_input[14975]), .Z(o[4975]) );
  AND U5586 ( .A(p_input[4974]), .B(p_input[14974]), .Z(o[4974]) );
  AND U5587 ( .A(p_input[4973]), .B(p_input[14973]), .Z(o[4973]) );
  AND U5588 ( .A(p_input[4972]), .B(p_input[14972]), .Z(o[4972]) );
  AND U5589 ( .A(p_input[4971]), .B(p_input[14971]), .Z(o[4971]) );
  AND U5590 ( .A(p_input[4970]), .B(p_input[14970]), .Z(o[4970]) );
  AND U5591 ( .A(p_input[496]), .B(p_input[10496]), .Z(o[496]) );
  AND U5592 ( .A(p_input[4969]), .B(p_input[14969]), .Z(o[4969]) );
  AND U5593 ( .A(p_input[4968]), .B(p_input[14968]), .Z(o[4968]) );
  AND U5594 ( .A(p_input[4967]), .B(p_input[14967]), .Z(o[4967]) );
  AND U5595 ( .A(p_input[4966]), .B(p_input[14966]), .Z(o[4966]) );
  AND U5596 ( .A(p_input[4965]), .B(p_input[14965]), .Z(o[4965]) );
  AND U5597 ( .A(p_input[4964]), .B(p_input[14964]), .Z(o[4964]) );
  AND U5598 ( .A(p_input[4963]), .B(p_input[14963]), .Z(o[4963]) );
  AND U5599 ( .A(p_input[4962]), .B(p_input[14962]), .Z(o[4962]) );
  AND U5600 ( .A(p_input[4961]), .B(p_input[14961]), .Z(o[4961]) );
  AND U5601 ( .A(p_input[4960]), .B(p_input[14960]), .Z(o[4960]) );
  AND U5602 ( .A(p_input[495]), .B(p_input[10495]), .Z(o[495]) );
  AND U5603 ( .A(p_input[4959]), .B(p_input[14959]), .Z(o[4959]) );
  AND U5604 ( .A(p_input[4958]), .B(p_input[14958]), .Z(o[4958]) );
  AND U5605 ( .A(p_input[4957]), .B(p_input[14957]), .Z(o[4957]) );
  AND U5606 ( .A(p_input[4956]), .B(p_input[14956]), .Z(o[4956]) );
  AND U5607 ( .A(p_input[4955]), .B(p_input[14955]), .Z(o[4955]) );
  AND U5608 ( .A(p_input[4954]), .B(p_input[14954]), .Z(o[4954]) );
  AND U5609 ( .A(p_input[4953]), .B(p_input[14953]), .Z(o[4953]) );
  AND U5610 ( .A(p_input[4952]), .B(p_input[14952]), .Z(o[4952]) );
  AND U5611 ( .A(p_input[4951]), .B(p_input[14951]), .Z(o[4951]) );
  AND U5612 ( .A(p_input[4950]), .B(p_input[14950]), .Z(o[4950]) );
  AND U5613 ( .A(p_input[494]), .B(p_input[10494]), .Z(o[494]) );
  AND U5614 ( .A(p_input[4949]), .B(p_input[14949]), .Z(o[4949]) );
  AND U5615 ( .A(p_input[4948]), .B(p_input[14948]), .Z(o[4948]) );
  AND U5616 ( .A(p_input[4947]), .B(p_input[14947]), .Z(o[4947]) );
  AND U5617 ( .A(p_input[4946]), .B(p_input[14946]), .Z(o[4946]) );
  AND U5618 ( .A(p_input[4945]), .B(p_input[14945]), .Z(o[4945]) );
  AND U5619 ( .A(p_input[4944]), .B(p_input[14944]), .Z(o[4944]) );
  AND U5620 ( .A(p_input[4943]), .B(p_input[14943]), .Z(o[4943]) );
  AND U5621 ( .A(p_input[4942]), .B(p_input[14942]), .Z(o[4942]) );
  AND U5622 ( .A(p_input[4941]), .B(p_input[14941]), .Z(o[4941]) );
  AND U5623 ( .A(p_input[4940]), .B(p_input[14940]), .Z(o[4940]) );
  AND U5624 ( .A(p_input[493]), .B(p_input[10493]), .Z(o[493]) );
  AND U5625 ( .A(p_input[4939]), .B(p_input[14939]), .Z(o[4939]) );
  AND U5626 ( .A(p_input[4938]), .B(p_input[14938]), .Z(o[4938]) );
  AND U5627 ( .A(p_input[4937]), .B(p_input[14937]), .Z(o[4937]) );
  AND U5628 ( .A(p_input[4936]), .B(p_input[14936]), .Z(o[4936]) );
  AND U5629 ( .A(p_input[4935]), .B(p_input[14935]), .Z(o[4935]) );
  AND U5630 ( .A(p_input[4934]), .B(p_input[14934]), .Z(o[4934]) );
  AND U5631 ( .A(p_input[4933]), .B(p_input[14933]), .Z(o[4933]) );
  AND U5632 ( .A(p_input[4932]), .B(p_input[14932]), .Z(o[4932]) );
  AND U5633 ( .A(p_input[4931]), .B(p_input[14931]), .Z(o[4931]) );
  AND U5634 ( .A(p_input[4930]), .B(p_input[14930]), .Z(o[4930]) );
  AND U5635 ( .A(p_input[492]), .B(p_input[10492]), .Z(o[492]) );
  AND U5636 ( .A(p_input[4929]), .B(p_input[14929]), .Z(o[4929]) );
  AND U5637 ( .A(p_input[4928]), .B(p_input[14928]), .Z(o[4928]) );
  AND U5638 ( .A(p_input[4927]), .B(p_input[14927]), .Z(o[4927]) );
  AND U5639 ( .A(p_input[4926]), .B(p_input[14926]), .Z(o[4926]) );
  AND U5640 ( .A(p_input[4925]), .B(p_input[14925]), .Z(o[4925]) );
  AND U5641 ( .A(p_input[4924]), .B(p_input[14924]), .Z(o[4924]) );
  AND U5642 ( .A(p_input[4923]), .B(p_input[14923]), .Z(o[4923]) );
  AND U5643 ( .A(p_input[4922]), .B(p_input[14922]), .Z(o[4922]) );
  AND U5644 ( .A(p_input[4921]), .B(p_input[14921]), .Z(o[4921]) );
  AND U5645 ( .A(p_input[4920]), .B(p_input[14920]), .Z(o[4920]) );
  AND U5646 ( .A(p_input[491]), .B(p_input[10491]), .Z(o[491]) );
  AND U5647 ( .A(p_input[4919]), .B(p_input[14919]), .Z(o[4919]) );
  AND U5648 ( .A(p_input[4918]), .B(p_input[14918]), .Z(o[4918]) );
  AND U5649 ( .A(p_input[4917]), .B(p_input[14917]), .Z(o[4917]) );
  AND U5650 ( .A(p_input[4916]), .B(p_input[14916]), .Z(o[4916]) );
  AND U5651 ( .A(p_input[4915]), .B(p_input[14915]), .Z(o[4915]) );
  AND U5652 ( .A(p_input[4914]), .B(p_input[14914]), .Z(o[4914]) );
  AND U5653 ( .A(p_input[4913]), .B(p_input[14913]), .Z(o[4913]) );
  AND U5654 ( .A(p_input[4912]), .B(p_input[14912]), .Z(o[4912]) );
  AND U5655 ( .A(p_input[4911]), .B(p_input[14911]), .Z(o[4911]) );
  AND U5656 ( .A(p_input[4910]), .B(p_input[14910]), .Z(o[4910]) );
  AND U5657 ( .A(p_input[490]), .B(p_input[10490]), .Z(o[490]) );
  AND U5658 ( .A(p_input[4909]), .B(p_input[14909]), .Z(o[4909]) );
  AND U5659 ( .A(p_input[4908]), .B(p_input[14908]), .Z(o[4908]) );
  AND U5660 ( .A(p_input[4907]), .B(p_input[14907]), .Z(o[4907]) );
  AND U5661 ( .A(p_input[4906]), .B(p_input[14906]), .Z(o[4906]) );
  AND U5662 ( .A(p_input[4905]), .B(p_input[14905]), .Z(o[4905]) );
  AND U5663 ( .A(p_input[4904]), .B(p_input[14904]), .Z(o[4904]) );
  AND U5664 ( .A(p_input[4903]), .B(p_input[14903]), .Z(o[4903]) );
  AND U5665 ( .A(p_input[4902]), .B(p_input[14902]), .Z(o[4902]) );
  AND U5666 ( .A(p_input[4901]), .B(p_input[14901]), .Z(o[4901]) );
  AND U5667 ( .A(p_input[4900]), .B(p_input[14900]), .Z(o[4900]) );
  AND U5668 ( .A(p_input[48]), .B(p_input[10048]), .Z(o[48]) );
  AND U5669 ( .A(p_input[489]), .B(p_input[10489]), .Z(o[489]) );
  AND U5670 ( .A(p_input[4899]), .B(p_input[14899]), .Z(o[4899]) );
  AND U5671 ( .A(p_input[4898]), .B(p_input[14898]), .Z(o[4898]) );
  AND U5672 ( .A(p_input[4897]), .B(p_input[14897]), .Z(o[4897]) );
  AND U5673 ( .A(p_input[4896]), .B(p_input[14896]), .Z(o[4896]) );
  AND U5674 ( .A(p_input[4895]), .B(p_input[14895]), .Z(o[4895]) );
  AND U5675 ( .A(p_input[4894]), .B(p_input[14894]), .Z(o[4894]) );
  AND U5676 ( .A(p_input[4893]), .B(p_input[14893]), .Z(o[4893]) );
  AND U5677 ( .A(p_input[4892]), .B(p_input[14892]), .Z(o[4892]) );
  AND U5678 ( .A(p_input[4891]), .B(p_input[14891]), .Z(o[4891]) );
  AND U5679 ( .A(p_input[4890]), .B(p_input[14890]), .Z(o[4890]) );
  AND U5680 ( .A(p_input[488]), .B(p_input[10488]), .Z(o[488]) );
  AND U5681 ( .A(p_input[4889]), .B(p_input[14889]), .Z(o[4889]) );
  AND U5682 ( .A(p_input[4888]), .B(p_input[14888]), .Z(o[4888]) );
  AND U5683 ( .A(p_input[4887]), .B(p_input[14887]), .Z(o[4887]) );
  AND U5684 ( .A(p_input[4886]), .B(p_input[14886]), .Z(o[4886]) );
  AND U5685 ( .A(p_input[4885]), .B(p_input[14885]), .Z(o[4885]) );
  AND U5686 ( .A(p_input[4884]), .B(p_input[14884]), .Z(o[4884]) );
  AND U5687 ( .A(p_input[4883]), .B(p_input[14883]), .Z(o[4883]) );
  AND U5688 ( .A(p_input[4882]), .B(p_input[14882]), .Z(o[4882]) );
  AND U5689 ( .A(p_input[4881]), .B(p_input[14881]), .Z(o[4881]) );
  AND U5690 ( .A(p_input[4880]), .B(p_input[14880]), .Z(o[4880]) );
  AND U5691 ( .A(p_input[487]), .B(p_input[10487]), .Z(o[487]) );
  AND U5692 ( .A(p_input[4879]), .B(p_input[14879]), .Z(o[4879]) );
  AND U5693 ( .A(p_input[4878]), .B(p_input[14878]), .Z(o[4878]) );
  AND U5694 ( .A(p_input[4877]), .B(p_input[14877]), .Z(o[4877]) );
  AND U5695 ( .A(p_input[4876]), .B(p_input[14876]), .Z(o[4876]) );
  AND U5696 ( .A(p_input[4875]), .B(p_input[14875]), .Z(o[4875]) );
  AND U5697 ( .A(p_input[4874]), .B(p_input[14874]), .Z(o[4874]) );
  AND U5698 ( .A(p_input[4873]), .B(p_input[14873]), .Z(o[4873]) );
  AND U5699 ( .A(p_input[4872]), .B(p_input[14872]), .Z(o[4872]) );
  AND U5700 ( .A(p_input[4871]), .B(p_input[14871]), .Z(o[4871]) );
  AND U5701 ( .A(p_input[4870]), .B(p_input[14870]), .Z(o[4870]) );
  AND U5702 ( .A(p_input[486]), .B(p_input[10486]), .Z(o[486]) );
  AND U5703 ( .A(p_input[4869]), .B(p_input[14869]), .Z(o[4869]) );
  AND U5704 ( .A(p_input[4868]), .B(p_input[14868]), .Z(o[4868]) );
  AND U5705 ( .A(p_input[4867]), .B(p_input[14867]), .Z(o[4867]) );
  AND U5706 ( .A(p_input[4866]), .B(p_input[14866]), .Z(o[4866]) );
  AND U5707 ( .A(p_input[4865]), .B(p_input[14865]), .Z(o[4865]) );
  AND U5708 ( .A(p_input[4864]), .B(p_input[14864]), .Z(o[4864]) );
  AND U5709 ( .A(p_input[4863]), .B(p_input[14863]), .Z(o[4863]) );
  AND U5710 ( .A(p_input[4862]), .B(p_input[14862]), .Z(o[4862]) );
  AND U5711 ( .A(p_input[4861]), .B(p_input[14861]), .Z(o[4861]) );
  AND U5712 ( .A(p_input[4860]), .B(p_input[14860]), .Z(o[4860]) );
  AND U5713 ( .A(p_input[485]), .B(p_input[10485]), .Z(o[485]) );
  AND U5714 ( .A(p_input[4859]), .B(p_input[14859]), .Z(o[4859]) );
  AND U5715 ( .A(p_input[4858]), .B(p_input[14858]), .Z(o[4858]) );
  AND U5716 ( .A(p_input[4857]), .B(p_input[14857]), .Z(o[4857]) );
  AND U5717 ( .A(p_input[4856]), .B(p_input[14856]), .Z(o[4856]) );
  AND U5718 ( .A(p_input[4855]), .B(p_input[14855]), .Z(o[4855]) );
  AND U5719 ( .A(p_input[4854]), .B(p_input[14854]), .Z(o[4854]) );
  AND U5720 ( .A(p_input[4853]), .B(p_input[14853]), .Z(o[4853]) );
  AND U5721 ( .A(p_input[4852]), .B(p_input[14852]), .Z(o[4852]) );
  AND U5722 ( .A(p_input[4851]), .B(p_input[14851]), .Z(o[4851]) );
  AND U5723 ( .A(p_input[4850]), .B(p_input[14850]), .Z(o[4850]) );
  AND U5724 ( .A(p_input[484]), .B(p_input[10484]), .Z(o[484]) );
  AND U5725 ( .A(p_input[4849]), .B(p_input[14849]), .Z(o[4849]) );
  AND U5726 ( .A(p_input[4848]), .B(p_input[14848]), .Z(o[4848]) );
  AND U5727 ( .A(p_input[4847]), .B(p_input[14847]), .Z(o[4847]) );
  AND U5728 ( .A(p_input[4846]), .B(p_input[14846]), .Z(o[4846]) );
  AND U5729 ( .A(p_input[4845]), .B(p_input[14845]), .Z(o[4845]) );
  AND U5730 ( .A(p_input[4844]), .B(p_input[14844]), .Z(o[4844]) );
  AND U5731 ( .A(p_input[4843]), .B(p_input[14843]), .Z(o[4843]) );
  AND U5732 ( .A(p_input[4842]), .B(p_input[14842]), .Z(o[4842]) );
  AND U5733 ( .A(p_input[4841]), .B(p_input[14841]), .Z(o[4841]) );
  AND U5734 ( .A(p_input[4840]), .B(p_input[14840]), .Z(o[4840]) );
  AND U5735 ( .A(p_input[483]), .B(p_input[10483]), .Z(o[483]) );
  AND U5736 ( .A(p_input[4839]), .B(p_input[14839]), .Z(o[4839]) );
  AND U5737 ( .A(p_input[4838]), .B(p_input[14838]), .Z(o[4838]) );
  AND U5738 ( .A(p_input[4837]), .B(p_input[14837]), .Z(o[4837]) );
  AND U5739 ( .A(p_input[4836]), .B(p_input[14836]), .Z(o[4836]) );
  AND U5740 ( .A(p_input[4835]), .B(p_input[14835]), .Z(o[4835]) );
  AND U5741 ( .A(p_input[4834]), .B(p_input[14834]), .Z(o[4834]) );
  AND U5742 ( .A(p_input[4833]), .B(p_input[14833]), .Z(o[4833]) );
  AND U5743 ( .A(p_input[4832]), .B(p_input[14832]), .Z(o[4832]) );
  AND U5744 ( .A(p_input[4831]), .B(p_input[14831]), .Z(o[4831]) );
  AND U5745 ( .A(p_input[4830]), .B(p_input[14830]), .Z(o[4830]) );
  AND U5746 ( .A(p_input[482]), .B(p_input[10482]), .Z(o[482]) );
  AND U5747 ( .A(p_input[4829]), .B(p_input[14829]), .Z(o[4829]) );
  AND U5748 ( .A(p_input[4828]), .B(p_input[14828]), .Z(o[4828]) );
  AND U5749 ( .A(p_input[4827]), .B(p_input[14827]), .Z(o[4827]) );
  AND U5750 ( .A(p_input[4826]), .B(p_input[14826]), .Z(o[4826]) );
  AND U5751 ( .A(p_input[4825]), .B(p_input[14825]), .Z(o[4825]) );
  AND U5752 ( .A(p_input[4824]), .B(p_input[14824]), .Z(o[4824]) );
  AND U5753 ( .A(p_input[4823]), .B(p_input[14823]), .Z(o[4823]) );
  AND U5754 ( .A(p_input[4822]), .B(p_input[14822]), .Z(o[4822]) );
  AND U5755 ( .A(p_input[4821]), .B(p_input[14821]), .Z(o[4821]) );
  AND U5756 ( .A(p_input[4820]), .B(p_input[14820]), .Z(o[4820]) );
  AND U5757 ( .A(p_input[481]), .B(p_input[10481]), .Z(o[481]) );
  AND U5758 ( .A(p_input[4819]), .B(p_input[14819]), .Z(o[4819]) );
  AND U5759 ( .A(p_input[4818]), .B(p_input[14818]), .Z(o[4818]) );
  AND U5760 ( .A(p_input[4817]), .B(p_input[14817]), .Z(o[4817]) );
  AND U5761 ( .A(p_input[4816]), .B(p_input[14816]), .Z(o[4816]) );
  AND U5762 ( .A(p_input[4815]), .B(p_input[14815]), .Z(o[4815]) );
  AND U5763 ( .A(p_input[4814]), .B(p_input[14814]), .Z(o[4814]) );
  AND U5764 ( .A(p_input[4813]), .B(p_input[14813]), .Z(o[4813]) );
  AND U5765 ( .A(p_input[4812]), .B(p_input[14812]), .Z(o[4812]) );
  AND U5766 ( .A(p_input[4811]), .B(p_input[14811]), .Z(o[4811]) );
  AND U5767 ( .A(p_input[4810]), .B(p_input[14810]), .Z(o[4810]) );
  AND U5768 ( .A(p_input[480]), .B(p_input[10480]), .Z(o[480]) );
  AND U5769 ( .A(p_input[4809]), .B(p_input[14809]), .Z(o[4809]) );
  AND U5770 ( .A(p_input[4808]), .B(p_input[14808]), .Z(o[4808]) );
  AND U5771 ( .A(p_input[4807]), .B(p_input[14807]), .Z(o[4807]) );
  AND U5772 ( .A(p_input[4806]), .B(p_input[14806]), .Z(o[4806]) );
  AND U5773 ( .A(p_input[4805]), .B(p_input[14805]), .Z(o[4805]) );
  AND U5774 ( .A(p_input[4804]), .B(p_input[14804]), .Z(o[4804]) );
  AND U5775 ( .A(p_input[4803]), .B(p_input[14803]), .Z(o[4803]) );
  AND U5776 ( .A(p_input[4802]), .B(p_input[14802]), .Z(o[4802]) );
  AND U5777 ( .A(p_input[4801]), .B(p_input[14801]), .Z(o[4801]) );
  AND U5778 ( .A(p_input[4800]), .B(p_input[14800]), .Z(o[4800]) );
  AND U5779 ( .A(p_input[47]), .B(p_input[10047]), .Z(o[47]) );
  AND U5780 ( .A(p_input[479]), .B(p_input[10479]), .Z(o[479]) );
  AND U5781 ( .A(p_input[4799]), .B(p_input[14799]), .Z(o[4799]) );
  AND U5782 ( .A(p_input[4798]), .B(p_input[14798]), .Z(o[4798]) );
  AND U5783 ( .A(p_input[4797]), .B(p_input[14797]), .Z(o[4797]) );
  AND U5784 ( .A(p_input[4796]), .B(p_input[14796]), .Z(o[4796]) );
  AND U5785 ( .A(p_input[4795]), .B(p_input[14795]), .Z(o[4795]) );
  AND U5786 ( .A(p_input[4794]), .B(p_input[14794]), .Z(o[4794]) );
  AND U5787 ( .A(p_input[4793]), .B(p_input[14793]), .Z(o[4793]) );
  AND U5788 ( .A(p_input[4792]), .B(p_input[14792]), .Z(o[4792]) );
  AND U5789 ( .A(p_input[4791]), .B(p_input[14791]), .Z(o[4791]) );
  AND U5790 ( .A(p_input[4790]), .B(p_input[14790]), .Z(o[4790]) );
  AND U5791 ( .A(p_input[478]), .B(p_input[10478]), .Z(o[478]) );
  AND U5792 ( .A(p_input[4789]), .B(p_input[14789]), .Z(o[4789]) );
  AND U5793 ( .A(p_input[4788]), .B(p_input[14788]), .Z(o[4788]) );
  AND U5794 ( .A(p_input[4787]), .B(p_input[14787]), .Z(o[4787]) );
  AND U5795 ( .A(p_input[4786]), .B(p_input[14786]), .Z(o[4786]) );
  AND U5796 ( .A(p_input[4785]), .B(p_input[14785]), .Z(o[4785]) );
  AND U5797 ( .A(p_input[4784]), .B(p_input[14784]), .Z(o[4784]) );
  AND U5798 ( .A(p_input[4783]), .B(p_input[14783]), .Z(o[4783]) );
  AND U5799 ( .A(p_input[4782]), .B(p_input[14782]), .Z(o[4782]) );
  AND U5800 ( .A(p_input[4781]), .B(p_input[14781]), .Z(o[4781]) );
  AND U5801 ( .A(p_input[4780]), .B(p_input[14780]), .Z(o[4780]) );
  AND U5802 ( .A(p_input[477]), .B(p_input[10477]), .Z(o[477]) );
  AND U5803 ( .A(p_input[4779]), .B(p_input[14779]), .Z(o[4779]) );
  AND U5804 ( .A(p_input[4778]), .B(p_input[14778]), .Z(o[4778]) );
  AND U5805 ( .A(p_input[4777]), .B(p_input[14777]), .Z(o[4777]) );
  AND U5806 ( .A(p_input[4776]), .B(p_input[14776]), .Z(o[4776]) );
  AND U5807 ( .A(p_input[4775]), .B(p_input[14775]), .Z(o[4775]) );
  AND U5808 ( .A(p_input[4774]), .B(p_input[14774]), .Z(o[4774]) );
  AND U5809 ( .A(p_input[4773]), .B(p_input[14773]), .Z(o[4773]) );
  AND U5810 ( .A(p_input[4772]), .B(p_input[14772]), .Z(o[4772]) );
  AND U5811 ( .A(p_input[4771]), .B(p_input[14771]), .Z(o[4771]) );
  AND U5812 ( .A(p_input[4770]), .B(p_input[14770]), .Z(o[4770]) );
  AND U5813 ( .A(p_input[476]), .B(p_input[10476]), .Z(o[476]) );
  AND U5814 ( .A(p_input[4769]), .B(p_input[14769]), .Z(o[4769]) );
  AND U5815 ( .A(p_input[4768]), .B(p_input[14768]), .Z(o[4768]) );
  AND U5816 ( .A(p_input[4767]), .B(p_input[14767]), .Z(o[4767]) );
  AND U5817 ( .A(p_input[4766]), .B(p_input[14766]), .Z(o[4766]) );
  AND U5818 ( .A(p_input[4765]), .B(p_input[14765]), .Z(o[4765]) );
  AND U5819 ( .A(p_input[4764]), .B(p_input[14764]), .Z(o[4764]) );
  AND U5820 ( .A(p_input[4763]), .B(p_input[14763]), .Z(o[4763]) );
  AND U5821 ( .A(p_input[4762]), .B(p_input[14762]), .Z(o[4762]) );
  AND U5822 ( .A(p_input[4761]), .B(p_input[14761]), .Z(o[4761]) );
  AND U5823 ( .A(p_input[4760]), .B(p_input[14760]), .Z(o[4760]) );
  AND U5824 ( .A(p_input[475]), .B(p_input[10475]), .Z(o[475]) );
  AND U5825 ( .A(p_input[4759]), .B(p_input[14759]), .Z(o[4759]) );
  AND U5826 ( .A(p_input[4758]), .B(p_input[14758]), .Z(o[4758]) );
  AND U5827 ( .A(p_input[4757]), .B(p_input[14757]), .Z(o[4757]) );
  AND U5828 ( .A(p_input[4756]), .B(p_input[14756]), .Z(o[4756]) );
  AND U5829 ( .A(p_input[4755]), .B(p_input[14755]), .Z(o[4755]) );
  AND U5830 ( .A(p_input[4754]), .B(p_input[14754]), .Z(o[4754]) );
  AND U5831 ( .A(p_input[4753]), .B(p_input[14753]), .Z(o[4753]) );
  AND U5832 ( .A(p_input[4752]), .B(p_input[14752]), .Z(o[4752]) );
  AND U5833 ( .A(p_input[4751]), .B(p_input[14751]), .Z(o[4751]) );
  AND U5834 ( .A(p_input[4750]), .B(p_input[14750]), .Z(o[4750]) );
  AND U5835 ( .A(p_input[474]), .B(p_input[10474]), .Z(o[474]) );
  AND U5836 ( .A(p_input[4749]), .B(p_input[14749]), .Z(o[4749]) );
  AND U5837 ( .A(p_input[4748]), .B(p_input[14748]), .Z(o[4748]) );
  AND U5838 ( .A(p_input[4747]), .B(p_input[14747]), .Z(o[4747]) );
  AND U5839 ( .A(p_input[4746]), .B(p_input[14746]), .Z(o[4746]) );
  AND U5840 ( .A(p_input[4745]), .B(p_input[14745]), .Z(o[4745]) );
  AND U5841 ( .A(p_input[4744]), .B(p_input[14744]), .Z(o[4744]) );
  AND U5842 ( .A(p_input[4743]), .B(p_input[14743]), .Z(o[4743]) );
  AND U5843 ( .A(p_input[4742]), .B(p_input[14742]), .Z(o[4742]) );
  AND U5844 ( .A(p_input[4741]), .B(p_input[14741]), .Z(o[4741]) );
  AND U5845 ( .A(p_input[4740]), .B(p_input[14740]), .Z(o[4740]) );
  AND U5846 ( .A(p_input[473]), .B(p_input[10473]), .Z(o[473]) );
  AND U5847 ( .A(p_input[4739]), .B(p_input[14739]), .Z(o[4739]) );
  AND U5848 ( .A(p_input[4738]), .B(p_input[14738]), .Z(o[4738]) );
  AND U5849 ( .A(p_input[4737]), .B(p_input[14737]), .Z(o[4737]) );
  AND U5850 ( .A(p_input[4736]), .B(p_input[14736]), .Z(o[4736]) );
  AND U5851 ( .A(p_input[4735]), .B(p_input[14735]), .Z(o[4735]) );
  AND U5852 ( .A(p_input[4734]), .B(p_input[14734]), .Z(o[4734]) );
  AND U5853 ( .A(p_input[4733]), .B(p_input[14733]), .Z(o[4733]) );
  AND U5854 ( .A(p_input[4732]), .B(p_input[14732]), .Z(o[4732]) );
  AND U5855 ( .A(p_input[4731]), .B(p_input[14731]), .Z(o[4731]) );
  AND U5856 ( .A(p_input[4730]), .B(p_input[14730]), .Z(o[4730]) );
  AND U5857 ( .A(p_input[472]), .B(p_input[10472]), .Z(o[472]) );
  AND U5858 ( .A(p_input[4729]), .B(p_input[14729]), .Z(o[4729]) );
  AND U5859 ( .A(p_input[4728]), .B(p_input[14728]), .Z(o[4728]) );
  AND U5860 ( .A(p_input[4727]), .B(p_input[14727]), .Z(o[4727]) );
  AND U5861 ( .A(p_input[4726]), .B(p_input[14726]), .Z(o[4726]) );
  AND U5862 ( .A(p_input[4725]), .B(p_input[14725]), .Z(o[4725]) );
  AND U5863 ( .A(p_input[4724]), .B(p_input[14724]), .Z(o[4724]) );
  AND U5864 ( .A(p_input[4723]), .B(p_input[14723]), .Z(o[4723]) );
  AND U5865 ( .A(p_input[4722]), .B(p_input[14722]), .Z(o[4722]) );
  AND U5866 ( .A(p_input[4721]), .B(p_input[14721]), .Z(o[4721]) );
  AND U5867 ( .A(p_input[4720]), .B(p_input[14720]), .Z(o[4720]) );
  AND U5868 ( .A(p_input[471]), .B(p_input[10471]), .Z(o[471]) );
  AND U5869 ( .A(p_input[4719]), .B(p_input[14719]), .Z(o[4719]) );
  AND U5870 ( .A(p_input[4718]), .B(p_input[14718]), .Z(o[4718]) );
  AND U5871 ( .A(p_input[4717]), .B(p_input[14717]), .Z(o[4717]) );
  AND U5872 ( .A(p_input[4716]), .B(p_input[14716]), .Z(o[4716]) );
  AND U5873 ( .A(p_input[4715]), .B(p_input[14715]), .Z(o[4715]) );
  AND U5874 ( .A(p_input[4714]), .B(p_input[14714]), .Z(o[4714]) );
  AND U5875 ( .A(p_input[4713]), .B(p_input[14713]), .Z(o[4713]) );
  AND U5876 ( .A(p_input[4712]), .B(p_input[14712]), .Z(o[4712]) );
  AND U5877 ( .A(p_input[4711]), .B(p_input[14711]), .Z(o[4711]) );
  AND U5878 ( .A(p_input[4710]), .B(p_input[14710]), .Z(o[4710]) );
  AND U5879 ( .A(p_input[470]), .B(p_input[10470]), .Z(o[470]) );
  AND U5880 ( .A(p_input[4709]), .B(p_input[14709]), .Z(o[4709]) );
  AND U5881 ( .A(p_input[4708]), .B(p_input[14708]), .Z(o[4708]) );
  AND U5882 ( .A(p_input[4707]), .B(p_input[14707]), .Z(o[4707]) );
  AND U5883 ( .A(p_input[4706]), .B(p_input[14706]), .Z(o[4706]) );
  AND U5884 ( .A(p_input[4705]), .B(p_input[14705]), .Z(o[4705]) );
  AND U5885 ( .A(p_input[4704]), .B(p_input[14704]), .Z(o[4704]) );
  AND U5886 ( .A(p_input[4703]), .B(p_input[14703]), .Z(o[4703]) );
  AND U5887 ( .A(p_input[4702]), .B(p_input[14702]), .Z(o[4702]) );
  AND U5888 ( .A(p_input[4701]), .B(p_input[14701]), .Z(o[4701]) );
  AND U5889 ( .A(p_input[4700]), .B(p_input[14700]), .Z(o[4700]) );
  AND U5890 ( .A(p_input[46]), .B(p_input[10046]), .Z(o[46]) );
  AND U5891 ( .A(p_input[469]), .B(p_input[10469]), .Z(o[469]) );
  AND U5892 ( .A(p_input[4699]), .B(p_input[14699]), .Z(o[4699]) );
  AND U5893 ( .A(p_input[4698]), .B(p_input[14698]), .Z(o[4698]) );
  AND U5894 ( .A(p_input[4697]), .B(p_input[14697]), .Z(o[4697]) );
  AND U5895 ( .A(p_input[4696]), .B(p_input[14696]), .Z(o[4696]) );
  AND U5896 ( .A(p_input[4695]), .B(p_input[14695]), .Z(o[4695]) );
  AND U5897 ( .A(p_input[4694]), .B(p_input[14694]), .Z(o[4694]) );
  AND U5898 ( .A(p_input[4693]), .B(p_input[14693]), .Z(o[4693]) );
  AND U5899 ( .A(p_input[4692]), .B(p_input[14692]), .Z(o[4692]) );
  AND U5900 ( .A(p_input[4691]), .B(p_input[14691]), .Z(o[4691]) );
  AND U5901 ( .A(p_input[4690]), .B(p_input[14690]), .Z(o[4690]) );
  AND U5902 ( .A(p_input[468]), .B(p_input[10468]), .Z(o[468]) );
  AND U5903 ( .A(p_input[4689]), .B(p_input[14689]), .Z(o[4689]) );
  AND U5904 ( .A(p_input[4688]), .B(p_input[14688]), .Z(o[4688]) );
  AND U5905 ( .A(p_input[4687]), .B(p_input[14687]), .Z(o[4687]) );
  AND U5906 ( .A(p_input[4686]), .B(p_input[14686]), .Z(o[4686]) );
  AND U5907 ( .A(p_input[4685]), .B(p_input[14685]), .Z(o[4685]) );
  AND U5908 ( .A(p_input[4684]), .B(p_input[14684]), .Z(o[4684]) );
  AND U5909 ( .A(p_input[4683]), .B(p_input[14683]), .Z(o[4683]) );
  AND U5910 ( .A(p_input[4682]), .B(p_input[14682]), .Z(o[4682]) );
  AND U5911 ( .A(p_input[4681]), .B(p_input[14681]), .Z(o[4681]) );
  AND U5912 ( .A(p_input[4680]), .B(p_input[14680]), .Z(o[4680]) );
  AND U5913 ( .A(p_input[467]), .B(p_input[10467]), .Z(o[467]) );
  AND U5914 ( .A(p_input[4679]), .B(p_input[14679]), .Z(o[4679]) );
  AND U5915 ( .A(p_input[4678]), .B(p_input[14678]), .Z(o[4678]) );
  AND U5916 ( .A(p_input[4677]), .B(p_input[14677]), .Z(o[4677]) );
  AND U5917 ( .A(p_input[4676]), .B(p_input[14676]), .Z(o[4676]) );
  AND U5918 ( .A(p_input[4675]), .B(p_input[14675]), .Z(o[4675]) );
  AND U5919 ( .A(p_input[4674]), .B(p_input[14674]), .Z(o[4674]) );
  AND U5920 ( .A(p_input[4673]), .B(p_input[14673]), .Z(o[4673]) );
  AND U5921 ( .A(p_input[4672]), .B(p_input[14672]), .Z(o[4672]) );
  AND U5922 ( .A(p_input[4671]), .B(p_input[14671]), .Z(o[4671]) );
  AND U5923 ( .A(p_input[4670]), .B(p_input[14670]), .Z(o[4670]) );
  AND U5924 ( .A(p_input[466]), .B(p_input[10466]), .Z(o[466]) );
  AND U5925 ( .A(p_input[4669]), .B(p_input[14669]), .Z(o[4669]) );
  AND U5926 ( .A(p_input[4668]), .B(p_input[14668]), .Z(o[4668]) );
  AND U5927 ( .A(p_input[4667]), .B(p_input[14667]), .Z(o[4667]) );
  AND U5928 ( .A(p_input[4666]), .B(p_input[14666]), .Z(o[4666]) );
  AND U5929 ( .A(p_input[4665]), .B(p_input[14665]), .Z(o[4665]) );
  AND U5930 ( .A(p_input[4664]), .B(p_input[14664]), .Z(o[4664]) );
  AND U5931 ( .A(p_input[4663]), .B(p_input[14663]), .Z(o[4663]) );
  AND U5932 ( .A(p_input[4662]), .B(p_input[14662]), .Z(o[4662]) );
  AND U5933 ( .A(p_input[4661]), .B(p_input[14661]), .Z(o[4661]) );
  AND U5934 ( .A(p_input[4660]), .B(p_input[14660]), .Z(o[4660]) );
  AND U5935 ( .A(p_input[465]), .B(p_input[10465]), .Z(o[465]) );
  AND U5936 ( .A(p_input[4659]), .B(p_input[14659]), .Z(o[4659]) );
  AND U5937 ( .A(p_input[4658]), .B(p_input[14658]), .Z(o[4658]) );
  AND U5938 ( .A(p_input[4657]), .B(p_input[14657]), .Z(o[4657]) );
  AND U5939 ( .A(p_input[4656]), .B(p_input[14656]), .Z(o[4656]) );
  AND U5940 ( .A(p_input[4655]), .B(p_input[14655]), .Z(o[4655]) );
  AND U5941 ( .A(p_input[4654]), .B(p_input[14654]), .Z(o[4654]) );
  AND U5942 ( .A(p_input[4653]), .B(p_input[14653]), .Z(o[4653]) );
  AND U5943 ( .A(p_input[4652]), .B(p_input[14652]), .Z(o[4652]) );
  AND U5944 ( .A(p_input[4651]), .B(p_input[14651]), .Z(o[4651]) );
  AND U5945 ( .A(p_input[4650]), .B(p_input[14650]), .Z(o[4650]) );
  AND U5946 ( .A(p_input[464]), .B(p_input[10464]), .Z(o[464]) );
  AND U5947 ( .A(p_input[4649]), .B(p_input[14649]), .Z(o[4649]) );
  AND U5948 ( .A(p_input[4648]), .B(p_input[14648]), .Z(o[4648]) );
  AND U5949 ( .A(p_input[4647]), .B(p_input[14647]), .Z(o[4647]) );
  AND U5950 ( .A(p_input[4646]), .B(p_input[14646]), .Z(o[4646]) );
  AND U5951 ( .A(p_input[4645]), .B(p_input[14645]), .Z(o[4645]) );
  AND U5952 ( .A(p_input[4644]), .B(p_input[14644]), .Z(o[4644]) );
  AND U5953 ( .A(p_input[4643]), .B(p_input[14643]), .Z(o[4643]) );
  AND U5954 ( .A(p_input[4642]), .B(p_input[14642]), .Z(o[4642]) );
  AND U5955 ( .A(p_input[4641]), .B(p_input[14641]), .Z(o[4641]) );
  AND U5956 ( .A(p_input[4640]), .B(p_input[14640]), .Z(o[4640]) );
  AND U5957 ( .A(p_input[463]), .B(p_input[10463]), .Z(o[463]) );
  AND U5958 ( .A(p_input[4639]), .B(p_input[14639]), .Z(o[4639]) );
  AND U5959 ( .A(p_input[4638]), .B(p_input[14638]), .Z(o[4638]) );
  AND U5960 ( .A(p_input[4637]), .B(p_input[14637]), .Z(o[4637]) );
  AND U5961 ( .A(p_input[4636]), .B(p_input[14636]), .Z(o[4636]) );
  AND U5962 ( .A(p_input[4635]), .B(p_input[14635]), .Z(o[4635]) );
  AND U5963 ( .A(p_input[4634]), .B(p_input[14634]), .Z(o[4634]) );
  AND U5964 ( .A(p_input[4633]), .B(p_input[14633]), .Z(o[4633]) );
  AND U5965 ( .A(p_input[4632]), .B(p_input[14632]), .Z(o[4632]) );
  AND U5966 ( .A(p_input[4631]), .B(p_input[14631]), .Z(o[4631]) );
  AND U5967 ( .A(p_input[4630]), .B(p_input[14630]), .Z(o[4630]) );
  AND U5968 ( .A(p_input[462]), .B(p_input[10462]), .Z(o[462]) );
  AND U5969 ( .A(p_input[4629]), .B(p_input[14629]), .Z(o[4629]) );
  AND U5970 ( .A(p_input[4628]), .B(p_input[14628]), .Z(o[4628]) );
  AND U5971 ( .A(p_input[4627]), .B(p_input[14627]), .Z(o[4627]) );
  AND U5972 ( .A(p_input[4626]), .B(p_input[14626]), .Z(o[4626]) );
  AND U5973 ( .A(p_input[4625]), .B(p_input[14625]), .Z(o[4625]) );
  AND U5974 ( .A(p_input[4624]), .B(p_input[14624]), .Z(o[4624]) );
  AND U5975 ( .A(p_input[4623]), .B(p_input[14623]), .Z(o[4623]) );
  AND U5976 ( .A(p_input[4622]), .B(p_input[14622]), .Z(o[4622]) );
  AND U5977 ( .A(p_input[4621]), .B(p_input[14621]), .Z(o[4621]) );
  AND U5978 ( .A(p_input[4620]), .B(p_input[14620]), .Z(o[4620]) );
  AND U5979 ( .A(p_input[461]), .B(p_input[10461]), .Z(o[461]) );
  AND U5980 ( .A(p_input[4619]), .B(p_input[14619]), .Z(o[4619]) );
  AND U5981 ( .A(p_input[4618]), .B(p_input[14618]), .Z(o[4618]) );
  AND U5982 ( .A(p_input[4617]), .B(p_input[14617]), .Z(o[4617]) );
  AND U5983 ( .A(p_input[4616]), .B(p_input[14616]), .Z(o[4616]) );
  AND U5984 ( .A(p_input[4615]), .B(p_input[14615]), .Z(o[4615]) );
  AND U5985 ( .A(p_input[4614]), .B(p_input[14614]), .Z(o[4614]) );
  AND U5986 ( .A(p_input[4613]), .B(p_input[14613]), .Z(o[4613]) );
  AND U5987 ( .A(p_input[4612]), .B(p_input[14612]), .Z(o[4612]) );
  AND U5988 ( .A(p_input[4611]), .B(p_input[14611]), .Z(o[4611]) );
  AND U5989 ( .A(p_input[4610]), .B(p_input[14610]), .Z(o[4610]) );
  AND U5990 ( .A(p_input[460]), .B(p_input[10460]), .Z(o[460]) );
  AND U5991 ( .A(p_input[4609]), .B(p_input[14609]), .Z(o[4609]) );
  AND U5992 ( .A(p_input[4608]), .B(p_input[14608]), .Z(o[4608]) );
  AND U5993 ( .A(p_input[4607]), .B(p_input[14607]), .Z(o[4607]) );
  AND U5994 ( .A(p_input[4606]), .B(p_input[14606]), .Z(o[4606]) );
  AND U5995 ( .A(p_input[4605]), .B(p_input[14605]), .Z(o[4605]) );
  AND U5996 ( .A(p_input[4604]), .B(p_input[14604]), .Z(o[4604]) );
  AND U5997 ( .A(p_input[4603]), .B(p_input[14603]), .Z(o[4603]) );
  AND U5998 ( .A(p_input[4602]), .B(p_input[14602]), .Z(o[4602]) );
  AND U5999 ( .A(p_input[4601]), .B(p_input[14601]), .Z(o[4601]) );
  AND U6000 ( .A(p_input[4600]), .B(p_input[14600]), .Z(o[4600]) );
  AND U6001 ( .A(p_input[45]), .B(p_input[10045]), .Z(o[45]) );
  AND U6002 ( .A(p_input[459]), .B(p_input[10459]), .Z(o[459]) );
  AND U6003 ( .A(p_input[4599]), .B(p_input[14599]), .Z(o[4599]) );
  AND U6004 ( .A(p_input[4598]), .B(p_input[14598]), .Z(o[4598]) );
  AND U6005 ( .A(p_input[4597]), .B(p_input[14597]), .Z(o[4597]) );
  AND U6006 ( .A(p_input[4596]), .B(p_input[14596]), .Z(o[4596]) );
  AND U6007 ( .A(p_input[4595]), .B(p_input[14595]), .Z(o[4595]) );
  AND U6008 ( .A(p_input[4594]), .B(p_input[14594]), .Z(o[4594]) );
  AND U6009 ( .A(p_input[4593]), .B(p_input[14593]), .Z(o[4593]) );
  AND U6010 ( .A(p_input[4592]), .B(p_input[14592]), .Z(o[4592]) );
  AND U6011 ( .A(p_input[4591]), .B(p_input[14591]), .Z(o[4591]) );
  AND U6012 ( .A(p_input[4590]), .B(p_input[14590]), .Z(o[4590]) );
  AND U6013 ( .A(p_input[458]), .B(p_input[10458]), .Z(o[458]) );
  AND U6014 ( .A(p_input[4589]), .B(p_input[14589]), .Z(o[4589]) );
  AND U6015 ( .A(p_input[4588]), .B(p_input[14588]), .Z(o[4588]) );
  AND U6016 ( .A(p_input[4587]), .B(p_input[14587]), .Z(o[4587]) );
  AND U6017 ( .A(p_input[4586]), .B(p_input[14586]), .Z(o[4586]) );
  AND U6018 ( .A(p_input[4585]), .B(p_input[14585]), .Z(o[4585]) );
  AND U6019 ( .A(p_input[4584]), .B(p_input[14584]), .Z(o[4584]) );
  AND U6020 ( .A(p_input[4583]), .B(p_input[14583]), .Z(o[4583]) );
  AND U6021 ( .A(p_input[4582]), .B(p_input[14582]), .Z(o[4582]) );
  AND U6022 ( .A(p_input[4581]), .B(p_input[14581]), .Z(o[4581]) );
  AND U6023 ( .A(p_input[4580]), .B(p_input[14580]), .Z(o[4580]) );
  AND U6024 ( .A(p_input[457]), .B(p_input[10457]), .Z(o[457]) );
  AND U6025 ( .A(p_input[4579]), .B(p_input[14579]), .Z(o[4579]) );
  AND U6026 ( .A(p_input[4578]), .B(p_input[14578]), .Z(o[4578]) );
  AND U6027 ( .A(p_input[4577]), .B(p_input[14577]), .Z(o[4577]) );
  AND U6028 ( .A(p_input[4576]), .B(p_input[14576]), .Z(o[4576]) );
  AND U6029 ( .A(p_input[4575]), .B(p_input[14575]), .Z(o[4575]) );
  AND U6030 ( .A(p_input[4574]), .B(p_input[14574]), .Z(o[4574]) );
  AND U6031 ( .A(p_input[4573]), .B(p_input[14573]), .Z(o[4573]) );
  AND U6032 ( .A(p_input[4572]), .B(p_input[14572]), .Z(o[4572]) );
  AND U6033 ( .A(p_input[4571]), .B(p_input[14571]), .Z(o[4571]) );
  AND U6034 ( .A(p_input[4570]), .B(p_input[14570]), .Z(o[4570]) );
  AND U6035 ( .A(p_input[456]), .B(p_input[10456]), .Z(o[456]) );
  AND U6036 ( .A(p_input[4569]), .B(p_input[14569]), .Z(o[4569]) );
  AND U6037 ( .A(p_input[4568]), .B(p_input[14568]), .Z(o[4568]) );
  AND U6038 ( .A(p_input[4567]), .B(p_input[14567]), .Z(o[4567]) );
  AND U6039 ( .A(p_input[4566]), .B(p_input[14566]), .Z(o[4566]) );
  AND U6040 ( .A(p_input[4565]), .B(p_input[14565]), .Z(o[4565]) );
  AND U6041 ( .A(p_input[4564]), .B(p_input[14564]), .Z(o[4564]) );
  AND U6042 ( .A(p_input[4563]), .B(p_input[14563]), .Z(o[4563]) );
  AND U6043 ( .A(p_input[4562]), .B(p_input[14562]), .Z(o[4562]) );
  AND U6044 ( .A(p_input[4561]), .B(p_input[14561]), .Z(o[4561]) );
  AND U6045 ( .A(p_input[4560]), .B(p_input[14560]), .Z(o[4560]) );
  AND U6046 ( .A(p_input[455]), .B(p_input[10455]), .Z(o[455]) );
  AND U6047 ( .A(p_input[4559]), .B(p_input[14559]), .Z(o[4559]) );
  AND U6048 ( .A(p_input[4558]), .B(p_input[14558]), .Z(o[4558]) );
  AND U6049 ( .A(p_input[4557]), .B(p_input[14557]), .Z(o[4557]) );
  AND U6050 ( .A(p_input[4556]), .B(p_input[14556]), .Z(o[4556]) );
  AND U6051 ( .A(p_input[4555]), .B(p_input[14555]), .Z(o[4555]) );
  AND U6052 ( .A(p_input[4554]), .B(p_input[14554]), .Z(o[4554]) );
  AND U6053 ( .A(p_input[4553]), .B(p_input[14553]), .Z(o[4553]) );
  AND U6054 ( .A(p_input[4552]), .B(p_input[14552]), .Z(o[4552]) );
  AND U6055 ( .A(p_input[4551]), .B(p_input[14551]), .Z(o[4551]) );
  AND U6056 ( .A(p_input[4550]), .B(p_input[14550]), .Z(o[4550]) );
  AND U6057 ( .A(p_input[454]), .B(p_input[10454]), .Z(o[454]) );
  AND U6058 ( .A(p_input[4549]), .B(p_input[14549]), .Z(o[4549]) );
  AND U6059 ( .A(p_input[4548]), .B(p_input[14548]), .Z(o[4548]) );
  AND U6060 ( .A(p_input[4547]), .B(p_input[14547]), .Z(o[4547]) );
  AND U6061 ( .A(p_input[4546]), .B(p_input[14546]), .Z(o[4546]) );
  AND U6062 ( .A(p_input[4545]), .B(p_input[14545]), .Z(o[4545]) );
  AND U6063 ( .A(p_input[4544]), .B(p_input[14544]), .Z(o[4544]) );
  AND U6064 ( .A(p_input[4543]), .B(p_input[14543]), .Z(o[4543]) );
  AND U6065 ( .A(p_input[4542]), .B(p_input[14542]), .Z(o[4542]) );
  AND U6066 ( .A(p_input[4541]), .B(p_input[14541]), .Z(o[4541]) );
  AND U6067 ( .A(p_input[4540]), .B(p_input[14540]), .Z(o[4540]) );
  AND U6068 ( .A(p_input[453]), .B(p_input[10453]), .Z(o[453]) );
  AND U6069 ( .A(p_input[4539]), .B(p_input[14539]), .Z(o[4539]) );
  AND U6070 ( .A(p_input[4538]), .B(p_input[14538]), .Z(o[4538]) );
  AND U6071 ( .A(p_input[4537]), .B(p_input[14537]), .Z(o[4537]) );
  AND U6072 ( .A(p_input[4536]), .B(p_input[14536]), .Z(o[4536]) );
  AND U6073 ( .A(p_input[4535]), .B(p_input[14535]), .Z(o[4535]) );
  AND U6074 ( .A(p_input[4534]), .B(p_input[14534]), .Z(o[4534]) );
  AND U6075 ( .A(p_input[4533]), .B(p_input[14533]), .Z(o[4533]) );
  AND U6076 ( .A(p_input[4532]), .B(p_input[14532]), .Z(o[4532]) );
  AND U6077 ( .A(p_input[4531]), .B(p_input[14531]), .Z(o[4531]) );
  AND U6078 ( .A(p_input[4530]), .B(p_input[14530]), .Z(o[4530]) );
  AND U6079 ( .A(p_input[452]), .B(p_input[10452]), .Z(o[452]) );
  AND U6080 ( .A(p_input[4529]), .B(p_input[14529]), .Z(o[4529]) );
  AND U6081 ( .A(p_input[4528]), .B(p_input[14528]), .Z(o[4528]) );
  AND U6082 ( .A(p_input[4527]), .B(p_input[14527]), .Z(o[4527]) );
  AND U6083 ( .A(p_input[4526]), .B(p_input[14526]), .Z(o[4526]) );
  AND U6084 ( .A(p_input[4525]), .B(p_input[14525]), .Z(o[4525]) );
  AND U6085 ( .A(p_input[4524]), .B(p_input[14524]), .Z(o[4524]) );
  AND U6086 ( .A(p_input[4523]), .B(p_input[14523]), .Z(o[4523]) );
  AND U6087 ( .A(p_input[4522]), .B(p_input[14522]), .Z(o[4522]) );
  AND U6088 ( .A(p_input[4521]), .B(p_input[14521]), .Z(o[4521]) );
  AND U6089 ( .A(p_input[4520]), .B(p_input[14520]), .Z(o[4520]) );
  AND U6090 ( .A(p_input[451]), .B(p_input[10451]), .Z(o[451]) );
  AND U6091 ( .A(p_input[4519]), .B(p_input[14519]), .Z(o[4519]) );
  AND U6092 ( .A(p_input[4518]), .B(p_input[14518]), .Z(o[4518]) );
  AND U6093 ( .A(p_input[4517]), .B(p_input[14517]), .Z(o[4517]) );
  AND U6094 ( .A(p_input[4516]), .B(p_input[14516]), .Z(o[4516]) );
  AND U6095 ( .A(p_input[4515]), .B(p_input[14515]), .Z(o[4515]) );
  AND U6096 ( .A(p_input[4514]), .B(p_input[14514]), .Z(o[4514]) );
  AND U6097 ( .A(p_input[4513]), .B(p_input[14513]), .Z(o[4513]) );
  AND U6098 ( .A(p_input[4512]), .B(p_input[14512]), .Z(o[4512]) );
  AND U6099 ( .A(p_input[4511]), .B(p_input[14511]), .Z(o[4511]) );
  AND U6100 ( .A(p_input[4510]), .B(p_input[14510]), .Z(o[4510]) );
  AND U6101 ( .A(p_input[450]), .B(p_input[10450]), .Z(o[450]) );
  AND U6102 ( .A(p_input[4509]), .B(p_input[14509]), .Z(o[4509]) );
  AND U6103 ( .A(p_input[4508]), .B(p_input[14508]), .Z(o[4508]) );
  AND U6104 ( .A(p_input[4507]), .B(p_input[14507]), .Z(o[4507]) );
  AND U6105 ( .A(p_input[4506]), .B(p_input[14506]), .Z(o[4506]) );
  AND U6106 ( .A(p_input[4505]), .B(p_input[14505]), .Z(o[4505]) );
  AND U6107 ( .A(p_input[4504]), .B(p_input[14504]), .Z(o[4504]) );
  AND U6108 ( .A(p_input[4503]), .B(p_input[14503]), .Z(o[4503]) );
  AND U6109 ( .A(p_input[4502]), .B(p_input[14502]), .Z(o[4502]) );
  AND U6110 ( .A(p_input[4501]), .B(p_input[14501]), .Z(o[4501]) );
  AND U6111 ( .A(p_input[4500]), .B(p_input[14500]), .Z(o[4500]) );
  AND U6112 ( .A(p_input[44]), .B(p_input[10044]), .Z(o[44]) );
  AND U6113 ( .A(p_input[449]), .B(p_input[10449]), .Z(o[449]) );
  AND U6114 ( .A(p_input[4499]), .B(p_input[14499]), .Z(o[4499]) );
  AND U6115 ( .A(p_input[4498]), .B(p_input[14498]), .Z(o[4498]) );
  AND U6116 ( .A(p_input[4497]), .B(p_input[14497]), .Z(o[4497]) );
  AND U6117 ( .A(p_input[4496]), .B(p_input[14496]), .Z(o[4496]) );
  AND U6118 ( .A(p_input[4495]), .B(p_input[14495]), .Z(o[4495]) );
  AND U6119 ( .A(p_input[4494]), .B(p_input[14494]), .Z(o[4494]) );
  AND U6120 ( .A(p_input[4493]), .B(p_input[14493]), .Z(o[4493]) );
  AND U6121 ( .A(p_input[4492]), .B(p_input[14492]), .Z(o[4492]) );
  AND U6122 ( .A(p_input[4491]), .B(p_input[14491]), .Z(o[4491]) );
  AND U6123 ( .A(p_input[4490]), .B(p_input[14490]), .Z(o[4490]) );
  AND U6124 ( .A(p_input[448]), .B(p_input[10448]), .Z(o[448]) );
  AND U6125 ( .A(p_input[4489]), .B(p_input[14489]), .Z(o[4489]) );
  AND U6126 ( .A(p_input[4488]), .B(p_input[14488]), .Z(o[4488]) );
  AND U6127 ( .A(p_input[4487]), .B(p_input[14487]), .Z(o[4487]) );
  AND U6128 ( .A(p_input[4486]), .B(p_input[14486]), .Z(o[4486]) );
  AND U6129 ( .A(p_input[4485]), .B(p_input[14485]), .Z(o[4485]) );
  AND U6130 ( .A(p_input[4484]), .B(p_input[14484]), .Z(o[4484]) );
  AND U6131 ( .A(p_input[4483]), .B(p_input[14483]), .Z(o[4483]) );
  AND U6132 ( .A(p_input[4482]), .B(p_input[14482]), .Z(o[4482]) );
  AND U6133 ( .A(p_input[4481]), .B(p_input[14481]), .Z(o[4481]) );
  AND U6134 ( .A(p_input[4480]), .B(p_input[14480]), .Z(o[4480]) );
  AND U6135 ( .A(p_input[447]), .B(p_input[10447]), .Z(o[447]) );
  AND U6136 ( .A(p_input[4479]), .B(p_input[14479]), .Z(o[4479]) );
  AND U6137 ( .A(p_input[4478]), .B(p_input[14478]), .Z(o[4478]) );
  AND U6138 ( .A(p_input[4477]), .B(p_input[14477]), .Z(o[4477]) );
  AND U6139 ( .A(p_input[4476]), .B(p_input[14476]), .Z(o[4476]) );
  AND U6140 ( .A(p_input[4475]), .B(p_input[14475]), .Z(o[4475]) );
  AND U6141 ( .A(p_input[4474]), .B(p_input[14474]), .Z(o[4474]) );
  AND U6142 ( .A(p_input[4473]), .B(p_input[14473]), .Z(o[4473]) );
  AND U6143 ( .A(p_input[4472]), .B(p_input[14472]), .Z(o[4472]) );
  AND U6144 ( .A(p_input[4471]), .B(p_input[14471]), .Z(o[4471]) );
  AND U6145 ( .A(p_input[4470]), .B(p_input[14470]), .Z(o[4470]) );
  AND U6146 ( .A(p_input[446]), .B(p_input[10446]), .Z(o[446]) );
  AND U6147 ( .A(p_input[4469]), .B(p_input[14469]), .Z(o[4469]) );
  AND U6148 ( .A(p_input[4468]), .B(p_input[14468]), .Z(o[4468]) );
  AND U6149 ( .A(p_input[4467]), .B(p_input[14467]), .Z(o[4467]) );
  AND U6150 ( .A(p_input[4466]), .B(p_input[14466]), .Z(o[4466]) );
  AND U6151 ( .A(p_input[4465]), .B(p_input[14465]), .Z(o[4465]) );
  AND U6152 ( .A(p_input[4464]), .B(p_input[14464]), .Z(o[4464]) );
  AND U6153 ( .A(p_input[4463]), .B(p_input[14463]), .Z(o[4463]) );
  AND U6154 ( .A(p_input[4462]), .B(p_input[14462]), .Z(o[4462]) );
  AND U6155 ( .A(p_input[4461]), .B(p_input[14461]), .Z(o[4461]) );
  AND U6156 ( .A(p_input[4460]), .B(p_input[14460]), .Z(o[4460]) );
  AND U6157 ( .A(p_input[445]), .B(p_input[10445]), .Z(o[445]) );
  AND U6158 ( .A(p_input[4459]), .B(p_input[14459]), .Z(o[4459]) );
  AND U6159 ( .A(p_input[4458]), .B(p_input[14458]), .Z(o[4458]) );
  AND U6160 ( .A(p_input[4457]), .B(p_input[14457]), .Z(o[4457]) );
  AND U6161 ( .A(p_input[4456]), .B(p_input[14456]), .Z(o[4456]) );
  AND U6162 ( .A(p_input[4455]), .B(p_input[14455]), .Z(o[4455]) );
  AND U6163 ( .A(p_input[4454]), .B(p_input[14454]), .Z(o[4454]) );
  AND U6164 ( .A(p_input[4453]), .B(p_input[14453]), .Z(o[4453]) );
  AND U6165 ( .A(p_input[4452]), .B(p_input[14452]), .Z(o[4452]) );
  AND U6166 ( .A(p_input[4451]), .B(p_input[14451]), .Z(o[4451]) );
  AND U6167 ( .A(p_input[4450]), .B(p_input[14450]), .Z(o[4450]) );
  AND U6168 ( .A(p_input[444]), .B(p_input[10444]), .Z(o[444]) );
  AND U6169 ( .A(p_input[4449]), .B(p_input[14449]), .Z(o[4449]) );
  AND U6170 ( .A(p_input[4448]), .B(p_input[14448]), .Z(o[4448]) );
  AND U6171 ( .A(p_input[4447]), .B(p_input[14447]), .Z(o[4447]) );
  AND U6172 ( .A(p_input[4446]), .B(p_input[14446]), .Z(o[4446]) );
  AND U6173 ( .A(p_input[4445]), .B(p_input[14445]), .Z(o[4445]) );
  AND U6174 ( .A(p_input[4444]), .B(p_input[14444]), .Z(o[4444]) );
  AND U6175 ( .A(p_input[4443]), .B(p_input[14443]), .Z(o[4443]) );
  AND U6176 ( .A(p_input[4442]), .B(p_input[14442]), .Z(o[4442]) );
  AND U6177 ( .A(p_input[4441]), .B(p_input[14441]), .Z(o[4441]) );
  AND U6178 ( .A(p_input[4440]), .B(p_input[14440]), .Z(o[4440]) );
  AND U6179 ( .A(p_input[443]), .B(p_input[10443]), .Z(o[443]) );
  AND U6180 ( .A(p_input[4439]), .B(p_input[14439]), .Z(o[4439]) );
  AND U6181 ( .A(p_input[4438]), .B(p_input[14438]), .Z(o[4438]) );
  AND U6182 ( .A(p_input[4437]), .B(p_input[14437]), .Z(o[4437]) );
  AND U6183 ( .A(p_input[4436]), .B(p_input[14436]), .Z(o[4436]) );
  AND U6184 ( .A(p_input[4435]), .B(p_input[14435]), .Z(o[4435]) );
  AND U6185 ( .A(p_input[4434]), .B(p_input[14434]), .Z(o[4434]) );
  AND U6186 ( .A(p_input[4433]), .B(p_input[14433]), .Z(o[4433]) );
  AND U6187 ( .A(p_input[4432]), .B(p_input[14432]), .Z(o[4432]) );
  AND U6188 ( .A(p_input[4431]), .B(p_input[14431]), .Z(o[4431]) );
  AND U6189 ( .A(p_input[4430]), .B(p_input[14430]), .Z(o[4430]) );
  AND U6190 ( .A(p_input[442]), .B(p_input[10442]), .Z(o[442]) );
  AND U6191 ( .A(p_input[4429]), .B(p_input[14429]), .Z(o[4429]) );
  AND U6192 ( .A(p_input[4428]), .B(p_input[14428]), .Z(o[4428]) );
  AND U6193 ( .A(p_input[4427]), .B(p_input[14427]), .Z(o[4427]) );
  AND U6194 ( .A(p_input[4426]), .B(p_input[14426]), .Z(o[4426]) );
  AND U6195 ( .A(p_input[4425]), .B(p_input[14425]), .Z(o[4425]) );
  AND U6196 ( .A(p_input[4424]), .B(p_input[14424]), .Z(o[4424]) );
  AND U6197 ( .A(p_input[4423]), .B(p_input[14423]), .Z(o[4423]) );
  AND U6198 ( .A(p_input[4422]), .B(p_input[14422]), .Z(o[4422]) );
  AND U6199 ( .A(p_input[4421]), .B(p_input[14421]), .Z(o[4421]) );
  AND U6200 ( .A(p_input[4420]), .B(p_input[14420]), .Z(o[4420]) );
  AND U6201 ( .A(p_input[441]), .B(p_input[10441]), .Z(o[441]) );
  AND U6202 ( .A(p_input[4419]), .B(p_input[14419]), .Z(o[4419]) );
  AND U6203 ( .A(p_input[4418]), .B(p_input[14418]), .Z(o[4418]) );
  AND U6204 ( .A(p_input[4417]), .B(p_input[14417]), .Z(o[4417]) );
  AND U6205 ( .A(p_input[4416]), .B(p_input[14416]), .Z(o[4416]) );
  AND U6206 ( .A(p_input[4415]), .B(p_input[14415]), .Z(o[4415]) );
  AND U6207 ( .A(p_input[4414]), .B(p_input[14414]), .Z(o[4414]) );
  AND U6208 ( .A(p_input[4413]), .B(p_input[14413]), .Z(o[4413]) );
  AND U6209 ( .A(p_input[4412]), .B(p_input[14412]), .Z(o[4412]) );
  AND U6210 ( .A(p_input[4411]), .B(p_input[14411]), .Z(o[4411]) );
  AND U6211 ( .A(p_input[4410]), .B(p_input[14410]), .Z(o[4410]) );
  AND U6212 ( .A(p_input[440]), .B(p_input[10440]), .Z(o[440]) );
  AND U6213 ( .A(p_input[4409]), .B(p_input[14409]), .Z(o[4409]) );
  AND U6214 ( .A(p_input[4408]), .B(p_input[14408]), .Z(o[4408]) );
  AND U6215 ( .A(p_input[4407]), .B(p_input[14407]), .Z(o[4407]) );
  AND U6216 ( .A(p_input[4406]), .B(p_input[14406]), .Z(o[4406]) );
  AND U6217 ( .A(p_input[4405]), .B(p_input[14405]), .Z(o[4405]) );
  AND U6218 ( .A(p_input[4404]), .B(p_input[14404]), .Z(o[4404]) );
  AND U6219 ( .A(p_input[4403]), .B(p_input[14403]), .Z(o[4403]) );
  AND U6220 ( .A(p_input[4402]), .B(p_input[14402]), .Z(o[4402]) );
  AND U6221 ( .A(p_input[4401]), .B(p_input[14401]), .Z(o[4401]) );
  AND U6222 ( .A(p_input[4400]), .B(p_input[14400]), .Z(o[4400]) );
  AND U6223 ( .A(p_input[43]), .B(p_input[10043]), .Z(o[43]) );
  AND U6224 ( .A(p_input[439]), .B(p_input[10439]), .Z(o[439]) );
  AND U6225 ( .A(p_input[4399]), .B(p_input[14399]), .Z(o[4399]) );
  AND U6226 ( .A(p_input[4398]), .B(p_input[14398]), .Z(o[4398]) );
  AND U6227 ( .A(p_input[4397]), .B(p_input[14397]), .Z(o[4397]) );
  AND U6228 ( .A(p_input[4396]), .B(p_input[14396]), .Z(o[4396]) );
  AND U6229 ( .A(p_input[4395]), .B(p_input[14395]), .Z(o[4395]) );
  AND U6230 ( .A(p_input[4394]), .B(p_input[14394]), .Z(o[4394]) );
  AND U6231 ( .A(p_input[4393]), .B(p_input[14393]), .Z(o[4393]) );
  AND U6232 ( .A(p_input[4392]), .B(p_input[14392]), .Z(o[4392]) );
  AND U6233 ( .A(p_input[4391]), .B(p_input[14391]), .Z(o[4391]) );
  AND U6234 ( .A(p_input[4390]), .B(p_input[14390]), .Z(o[4390]) );
  AND U6235 ( .A(p_input[438]), .B(p_input[10438]), .Z(o[438]) );
  AND U6236 ( .A(p_input[4389]), .B(p_input[14389]), .Z(o[4389]) );
  AND U6237 ( .A(p_input[4388]), .B(p_input[14388]), .Z(o[4388]) );
  AND U6238 ( .A(p_input[4387]), .B(p_input[14387]), .Z(o[4387]) );
  AND U6239 ( .A(p_input[4386]), .B(p_input[14386]), .Z(o[4386]) );
  AND U6240 ( .A(p_input[4385]), .B(p_input[14385]), .Z(o[4385]) );
  AND U6241 ( .A(p_input[4384]), .B(p_input[14384]), .Z(o[4384]) );
  AND U6242 ( .A(p_input[4383]), .B(p_input[14383]), .Z(o[4383]) );
  AND U6243 ( .A(p_input[4382]), .B(p_input[14382]), .Z(o[4382]) );
  AND U6244 ( .A(p_input[4381]), .B(p_input[14381]), .Z(o[4381]) );
  AND U6245 ( .A(p_input[4380]), .B(p_input[14380]), .Z(o[4380]) );
  AND U6246 ( .A(p_input[437]), .B(p_input[10437]), .Z(o[437]) );
  AND U6247 ( .A(p_input[4379]), .B(p_input[14379]), .Z(o[4379]) );
  AND U6248 ( .A(p_input[4378]), .B(p_input[14378]), .Z(o[4378]) );
  AND U6249 ( .A(p_input[4377]), .B(p_input[14377]), .Z(o[4377]) );
  AND U6250 ( .A(p_input[4376]), .B(p_input[14376]), .Z(o[4376]) );
  AND U6251 ( .A(p_input[4375]), .B(p_input[14375]), .Z(o[4375]) );
  AND U6252 ( .A(p_input[4374]), .B(p_input[14374]), .Z(o[4374]) );
  AND U6253 ( .A(p_input[4373]), .B(p_input[14373]), .Z(o[4373]) );
  AND U6254 ( .A(p_input[4372]), .B(p_input[14372]), .Z(o[4372]) );
  AND U6255 ( .A(p_input[4371]), .B(p_input[14371]), .Z(o[4371]) );
  AND U6256 ( .A(p_input[4370]), .B(p_input[14370]), .Z(o[4370]) );
  AND U6257 ( .A(p_input[436]), .B(p_input[10436]), .Z(o[436]) );
  AND U6258 ( .A(p_input[4369]), .B(p_input[14369]), .Z(o[4369]) );
  AND U6259 ( .A(p_input[4368]), .B(p_input[14368]), .Z(o[4368]) );
  AND U6260 ( .A(p_input[4367]), .B(p_input[14367]), .Z(o[4367]) );
  AND U6261 ( .A(p_input[4366]), .B(p_input[14366]), .Z(o[4366]) );
  AND U6262 ( .A(p_input[4365]), .B(p_input[14365]), .Z(o[4365]) );
  AND U6263 ( .A(p_input[4364]), .B(p_input[14364]), .Z(o[4364]) );
  AND U6264 ( .A(p_input[4363]), .B(p_input[14363]), .Z(o[4363]) );
  AND U6265 ( .A(p_input[4362]), .B(p_input[14362]), .Z(o[4362]) );
  AND U6266 ( .A(p_input[4361]), .B(p_input[14361]), .Z(o[4361]) );
  AND U6267 ( .A(p_input[4360]), .B(p_input[14360]), .Z(o[4360]) );
  AND U6268 ( .A(p_input[435]), .B(p_input[10435]), .Z(o[435]) );
  AND U6269 ( .A(p_input[4359]), .B(p_input[14359]), .Z(o[4359]) );
  AND U6270 ( .A(p_input[4358]), .B(p_input[14358]), .Z(o[4358]) );
  AND U6271 ( .A(p_input[4357]), .B(p_input[14357]), .Z(o[4357]) );
  AND U6272 ( .A(p_input[4356]), .B(p_input[14356]), .Z(o[4356]) );
  AND U6273 ( .A(p_input[4355]), .B(p_input[14355]), .Z(o[4355]) );
  AND U6274 ( .A(p_input[4354]), .B(p_input[14354]), .Z(o[4354]) );
  AND U6275 ( .A(p_input[4353]), .B(p_input[14353]), .Z(o[4353]) );
  AND U6276 ( .A(p_input[4352]), .B(p_input[14352]), .Z(o[4352]) );
  AND U6277 ( .A(p_input[4351]), .B(p_input[14351]), .Z(o[4351]) );
  AND U6278 ( .A(p_input[4350]), .B(p_input[14350]), .Z(o[4350]) );
  AND U6279 ( .A(p_input[434]), .B(p_input[10434]), .Z(o[434]) );
  AND U6280 ( .A(p_input[4349]), .B(p_input[14349]), .Z(o[4349]) );
  AND U6281 ( .A(p_input[4348]), .B(p_input[14348]), .Z(o[4348]) );
  AND U6282 ( .A(p_input[4347]), .B(p_input[14347]), .Z(o[4347]) );
  AND U6283 ( .A(p_input[4346]), .B(p_input[14346]), .Z(o[4346]) );
  AND U6284 ( .A(p_input[4345]), .B(p_input[14345]), .Z(o[4345]) );
  AND U6285 ( .A(p_input[4344]), .B(p_input[14344]), .Z(o[4344]) );
  AND U6286 ( .A(p_input[4343]), .B(p_input[14343]), .Z(o[4343]) );
  AND U6287 ( .A(p_input[4342]), .B(p_input[14342]), .Z(o[4342]) );
  AND U6288 ( .A(p_input[4341]), .B(p_input[14341]), .Z(o[4341]) );
  AND U6289 ( .A(p_input[4340]), .B(p_input[14340]), .Z(o[4340]) );
  AND U6290 ( .A(p_input[433]), .B(p_input[10433]), .Z(o[433]) );
  AND U6291 ( .A(p_input[4339]), .B(p_input[14339]), .Z(o[4339]) );
  AND U6292 ( .A(p_input[4338]), .B(p_input[14338]), .Z(o[4338]) );
  AND U6293 ( .A(p_input[4337]), .B(p_input[14337]), .Z(o[4337]) );
  AND U6294 ( .A(p_input[4336]), .B(p_input[14336]), .Z(o[4336]) );
  AND U6295 ( .A(p_input[4335]), .B(p_input[14335]), .Z(o[4335]) );
  AND U6296 ( .A(p_input[4334]), .B(p_input[14334]), .Z(o[4334]) );
  AND U6297 ( .A(p_input[4333]), .B(p_input[14333]), .Z(o[4333]) );
  AND U6298 ( .A(p_input[4332]), .B(p_input[14332]), .Z(o[4332]) );
  AND U6299 ( .A(p_input[4331]), .B(p_input[14331]), .Z(o[4331]) );
  AND U6300 ( .A(p_input[4330]), .B(p_input[14330]), .Z(o[4330]) );
  AND U6301 ( .A(p_input[432]), .B(p_input[10432]), .Z(o[432]) );
  AND U6302 ( .A(p_input[4329]), .B(p_input[14329]), .Z(o[4329]) );
  AND U6303 ( .A(p_input[4328]), .B(p_input[14328]), .Z(o[4328]) );
  AND U6304 ( .A(p_input[4327]), .B(p_input[14327]), .Z(o[4327]) );
  AND U6305 ( .A(p_input[4326]), .B(p_input[14326]), .Z(o[4326]) );
  AND U6306 ( .A(p_input[4325]), .B(p_input[14325]), .Z(o[4325]) );
  AND U6307 ( .A(p_input[4324]), .B(p_input[14324]), .Z(o[4324]) );
  AND U6308 ( .A(p_input[4323]), .B(p_input[14323]), .Z(o[4323]) );
  AND U6309 ( .A(p_input[4322]), .B(p_input[14322]), .Z(o[4322]) );
  AND U6310 ( .A(p_input[4321]), .B(p_input[14321]), .Z(o[4321]) );
  AND U6311 ( .A(p_input[4320]), .B(p_input[14320]), .Z(o[4320]) );
  AND U6312 ( .A(p_input[431]), .B(p_input[10431]), .Z(o[431]) );
  AND U6313 ( .A(p_input[4319]), .B(p_input[14319]), .Z(o[4319]) );
  AND U6314 ( .A(p_input[4318]), .B(p_input[14318]), .Z(o[4318]) );
  AND U6315 ( .A(p_input[4317]), .B(p_input[14317]), .Z(o[4317]) );
  AND U6316 ( .A(p_input[4316]), .B(p_input[14316]), .Z(o[4316]) );
  AND U6317 ( .A(p_input[4315]), .B(p_input[14315]), .Z(o[4315]) );
  AND U6318 ( .A(p_input[4314]), .B(p_input[14314]), .Z(o[4314]) );
  AND U6319 ( .A(p_input[4313]), .B(p_input[14313]), .Z(o[4313]) );
  AND U6320 ( .A(p_input[4312]), .B(p_input[14312]), .Z(o[4312]) );
  AND U6321 ( .A(p_input[4311]), .B(p_input[14311]), .Z(o[4311]) );
  AND U6322 ( .A(p_input[4310]), .B(p_input[14310]), .Z(o[4310]) );
  AND U6323 ( .A(p_input[430]), .B(p_input[10430]), .Z(o[430]) );
  AND U6324 ( .A(p_input[4309]), .B(p_input[14309]), .Z(o[4309]) );
  AND U6325 ( .A(p_input[4308]), .B(p_input[14308]), .Z(o[4308]) );
  AND U6326 ( .A(p_input[4307]), .B(p_input[14307]), .Z(o[4307]) );
  AND U6327 ( .A(p_input[4306]), .B(p_input[14306]), .Z(o[4306]) );
  AND U6328 ( .A(p_input[4305]), .B(p_input[14305]), .Z(o[4305]) );
  AND U6329 ( .A(p_input[4304]), .B(p_input[14304]), .Z(o[4304]) );
  AND U6330 ( .A(p_input[4303]), .B(p_input[14303]), .Z(o[4303]) );
  AND U6331 ( .A(p_input[4302]), .B(p_input[14302]), .Z(o[4302]) );
  AND U6332 ( .A(p_input[4301]), .B(p_input[14301]), .Z(o[4301]) );
  AND U6333 ( .A(p_input[4300]), .B(p_input[14300]), .Z(o[4300]) );
  AND U6334 ( .A(p_input[42]), .B(p_input[10042]), .Z(o[42]) );
  AND U6335 ( .A(p_input[429]), .B(p_input[10429]), .Z(o[429]) );
  AND U6336 ( .A(p_input[4299]), .B(p_input[14299]), .Z(o[4299]) );
  AND U6337 ( .A(p_input[4298]), .B(p_input[14298]), .Z(o[4298]) );
  AND U6338 ( .A(p_input[4297]), .B(p_input[14297]), .Z(o[4297]) );
  AND U6339 ( .A(p_input[4296]), .B(p_input[14296]), .Z(o[4296]) );
  AND U6340 ( .A(p_input[4295]), .B(p_input[14295]), .Z(o[4295]) );
  AND U6341 ( .A(p_input[4294]), .B(p_input[14294]), .Z(o[4294]) );
  AND U6342 ( .A(p_input[4293]), .B(p_input[14293]), .Z(o[4293]) );
  AND U6343 ( .A(p_input[4292]), .B(p_input[14292]), .Z(o[4292]) );
  AND U6344 ( .A(p_input[4291]), .B(p_input[14291]), .Z(o[4291]) );
  AND U6345 ( .A(p_input[4290]), .B(p_input[14290]), .Z(o[4290]) );
  AND U6346 ( .A(p_input[428]), .B(p_input[10428]), .Z(o[428]) );
  AND U6347 ( .A(p_input[4289]), .B(p_input[14289]), .Z(o[4289]) );
  AND U6348 ( .A(p_input[4288]), .B(p_input[14288]), .Z(o[4288]) );
  AND U6349 ( .A(p_input[4287]), .B(p_input[14287]), .Z(o[4287]) );
  AND U6350 ( .A(p_input[4286]), .B(p_input[14286]), .Z(o[4286]) );
  AND U6351 ( .A(p_input[4285]), .B(p_input[14285]), .Z(o[4285]) );
  AND U6352 ( .A(p_input[4284]), .B(p_input[14284]), .Z(o[4284]) );
  AND U6353 ( .A(p_input[4283]), .B(p_input[14283]), .Z(o[4283]) );
  AND U6354 ( .A(p_input[4282]), .B(p_input[14282]), .Z(o[4282]) );
  AND U6355 ( .A(p_input[4281]), .B(p_input[14281]), .Z(o[4281]) );
  AND U6356 ( .A(p_input[4280]), .B(p_input[14280]), .Z(o[4280]) );
  AND U6357 ( .A(p_input[427]), .B(p_input[10427]), .Z(o[427]) );
  AND U6358 ( .A(p_input[4279]), .B(p_input[14279]), .Z(o[4279]) );
  AND U6359 ( .A(p_input[4278]), .B(p_input[14278]), .Z(o[4278]) );
  AND U6360 ( .A(p_input[4277]), .B(p_input[14277]), .Z(o[4277]) );
  AND U6361 ( .A(p_input[4276]), .B(p_input[14276]), .Z(o[4276]) );
  AND U6362 ( .A(p_input[4275]), .B(p_input[14275]), .Z(o[4275]) );
  AND U6363 ( .A(p_input[4274]), .B(p_input[14274]), .Z(o[4274]) );
  AND U6364 ( .A(p_input[4273]), .B(p_input[14273]), .Z(o[4273]) );
  AND U6365 ( .A(p_input[4272]), .B(p_input[14272]), .Z(o[4272]) );
  AND U6366 ( .A(p_input[4271]), .B(p_input[14271]), .Z(o[4271]) );
  AND U6367 ( .A(p_input[4270]), .B(p_input[14270]), .Z(o[4270]) );
  AND U6368 ( .A(p_input[426]), .B(p_input[10426]), .Z(o[426]) );
  AND U6369 ( .A(p_input[4269]), .B(p_input[14269]), .Z(o[4269]) );
  AND U6370 ( .A(p_input[4268]), .B(p_input[14268]), .Z(o[4268]) );
  AND U6371 ( .A(p_input[4267]), .B(p_input[14267]), .Z(o[4267]) );
  AND U6372 ( .A(p_input[4266]), .B(p_input[14266]), .Z(o[4266]) );
  AND U6373 ( .A(p_input[4265]), .B(p_input[14265]), .Z(o[4265]) );
  AND U6374 ( .A(p_input[4264]), .B(p_input[14264]), .Z(o[4264]) );
  AND U6375 ( .A(p_input[4263]), .B(p_input[14263]), .Z(o[4263]) );
  AND U6376 ( .A(p_input[4262]), .B(p_input[14262]), .Z(o[4262]) );
  AND U6377 ( .A(p_input[4261]), .B(p_input[14261]), .Z(o[4261]) );
  AND U6378 ( .A(p_input[4260]), .B(p_input[14260]), .Z(o[4260]) );
  AND U6379 ( .A(p_input[425]), .B(p_input[10425]), .Z(o[425]) );
  AND U6380 ( .A(p_input[4259]), .B(p_input[14259]), .Z(o[4259]) );
  AND U6381 ( .A(p_input[4258]), .B(p_input[14258]), .Z(o[4258]) );
  AND U6382 ( .A(p_input[4257]), .B(p_input[14257]), .Z(o[4257]) );
  AND U6383 ( .A(p_input[4256]), .B(p_input[14256]), .Z(o[4256]) );
  AND U6384 ( .A(p_input[4255]), .B(p_input[14255]), .Z(o[4255]) );
  AND U6385 ( .A(p_input[4254]), .B(p_input[14254]), .Z(o[4254]) );
  AND U6386 ( .A(p_input[4253]), .B(p_input[14253]), .Z(o[4253]) );
  AND U6387 ( .A(p_input[4252]), .B(p_input[14252]), .Z(o[4252]) );
  AND U6388 ( .A(p_input[4251]), .B(p_input[14251]), .Z(o[4251]) );
  AND U6389 ( .A(p_input[4250]), .B(p_input[14250]), .Z(o[4250]) );
  AND U6390 ( .A(p_input[424]), .B(p_input[10424]), .Z(o[424]) );
  AND U6391 ( .A(p_input[4249]), .B(p_input[14249]), .Z(o[4249]) );
  AND U6392 ( .A(p_input[4248]), .B(p_input[14248]), .Z(o[4248]) );
  AND U6393 ( .A(p_input[4247]), .B(p_input[14247]), .Z(o[4247]) );
  AND U6394 ( .A(p_input[4246]), .B(p_input[14246]), .Z(o[4246]) );
  AND U6395 ( .A(p_input[4245]), .B(p_input[14245]), .Z(o[4245]) );
  AND U6396 ( .A(p_input[4244]), .B(p_input[14244]), .Z(o[4244]) );
  AND U6397 ( .A(p_input[4243]), .B(p_input[14243]), .Z(o[4243]) );
  AND U6398 ( .A(p_input[4242]), .B(p_input[14242]), .Z(o[4242]) );
  AND U6399 ( .A(p_input[4241]), .B(p_input[14241]), .Z(o[4241]) );
  AND U6400 ( .A(p_input[4240]), .B(p_input[14240]), .Z(o[4240]) );
  AND U6401 ( .A(p_input[423]), .B(p_input[10423]), .Z(o[423]) );
  AND U6402 ( .A(p_input[4239]), .B(p_input[14239]), .Z(o[4239]) );
  AND U6403 ( .A(p_input[4238]), .B(p_input[14238]), .Z(o[4238]) );
  AND U6404 ( .A(p_input[4237]), .B(p_input[14237]), .Z(o[4237]) );
  AND U6405 ( .A(p_input[4236]), .B(p_input[14236]), .Z(o[4236]) );
  AND U6406 ( .A(p_input[4235]), .B(p_input[14235]), .Z(o[4235]) );
  AND U6407 ( .A(p_input[4234]), .B(p_input[14234]), .Z(o[4234]) );
  AND U6408 ( .A(p_input[4233]), .B(p_input[14233]), .Z(o[4233]) );
  AND U6409 ( .A(p_input[4232]), .B(p_input[14232]), .Z(o[4232]) );
  AND U6410 ( .A(p_input[4231]), .B(p_input[14231]), .Z(o[4231]) );
  AND U6411 ( .A(p_input[4230]), .B(p_input[14230]), .Z(o[4230]) );
  AND U6412 ( .A(p_input[422]), .B(p_input[10422]), .Z(o[422]) );
  AND U6413 ( .A(p_input[4229]), .B(p_input[14229]), .Z(o[4229]) );
  AND U6414 ( .A(p_input[4228]), .B(p_input[14228]), .Z(o[4228]) );
  AND U6415 ( .A(p_input[4227]), .B(p_input[14227]), .Z(o[4227]) );
  AND U6416 ( .A(p_input[4226]), .B(p_input[14226]), .Z(o[4226]) );
  AND U6417 ( .A(p_input[4225]), .B(p_input[14225]), .Z(o[4225]) );
  AND U6418 ( .A(p_input[4224]), .B(p_input[14224]), .Z(o[4224]) );
  AND U6419 ( .A(p_input[4223]), .B(p_input[14223]), .Z(o[4223]) );
  AND U6420 ( .A(p_input[4222]), .B(p_input[14222]), .Z(o[4222]) );
  AND U6421 ( .A(p_input[4221]), .B(p_input[14221]), .Z(o[4221]) );
  AND U6422 ( .A(p_input[4220]), .B(p_input[14220]), .Z(o[4220]) );
  AND U6423 ( .A(p_input[421]), .B(p_input[10421]), .Z(o[421]) );
  AND U6424 ( .A(p_input[4219]), .B(p_input[14219]), .Z(o[4219]) );
  AND U6425 ( .A(p_input[4218]), .B(p_input[14218]), .Z(o[4218]) );
  AND U6426 ( .A(p_input[4217]), .B(p_input[14217]), .Z(o[4217]) );
  AND U6427 ( .A(p_input[4216]), .B(p_input[14216]), .Z(o[4216]) );
  AND U6428 ( .A(p_input[4215]), .B(p_input[14215]), .Z(o[4215]) );
  AND U6429 ( .A(p_input[4214]), .B(p_input[14214]), .Z(o[4214]) );
  AND U6430 ( .A(p_input[4213]), .B(p_input[14213]), .Z(o[4213]) );
  AND U6431 ( .A(p_input[4212]), .B(p_input[14212]), .Z(o[4212]) );
  AND U6432 ( .A(p_input[4211]), .B(p_input[14211]), .Z(o[4211]) );
  AND U6433 ( .A(p_input[4210]), .B(p_input[14210]), .Z(o[4210]) );
  AND U6434 ( .A(p_input[420]), .B(p_input[10420]), .Z(o[420]) );
  AND U6435 ( .A(p_input[4209]), .B(p_input[14209]), .Z(o[4209]) );
  AND U6436 ( .A(p_input[4208]), .B(p_input[14208]), .Z(o[4208]) );
  AND U6437 ( .A(p_input[4207]), .B(p_input[14207]), .Z(o[4207]) );
  AND U6438 ( .A(p_input[4206]), .B(p_input[14206]), .Z(o[4206]) );
  AND U6439 ( .A(p_input[4205]), .B(p_input[14205]), .Z(o[4205]) );
  AND U6440 ( .A(p_input[4204]), .B(p_input[14204]), .Z(o[4204]) );
  AND U6441 ( .A(p_input[4203]), .B(p_input[14203]), .Z(o[4203]) );
  AND U6442 ( .A(p_input[4202]), .B(p_input[14202]), .Z(o[4202]) );
  AND U6443 ( .A(p_input[4201]), .B(p_input[14201]), .Z(o[4201]) );
  AND U6444 ( .A(p_input[4200]), .B(p_input[14200]), .Z(o[4200]) );
  AND U6445 ( .A(p_input[41]), .B(p_input[10041]), .Z(o[41]) );
  AND U6446 ( .A(p_input[419]), .B(p_input[10419]), .Z(o[419]) );
  AND U6447 ( .A(p_input[4199]), .B(p_input[14199]), .Z(o[4199]) );
  AND U6448 ( .A(p_input[4198]), .B(p_input[14198]), .Z(o[4198]) );
  AND U6449 ( .A(p_input[4197]), .B(p_input[14197]), .Z(o[4197]) );
  AND U6450 ( .A(p_input[4196]), .B(p_input[14196]), .Z(o[4196]) );
  AND U6451 ( .A(p_input[4195]), .B(p_input[14195]), .Z(o[4195]) );
  AND U6452 ( .A(p_input[4194]), .B(p_input[14194]), .Z(o[4194]) );
  AND U6453 ( .A(p_input[4193]), .B(p_input[14193]), .Z(o[4193]) );
  AND U6454 ( .A(p_input[4192]), .B(p_input[14192]), .Z(o[4192]) );
  AND U6455 ( .A(p_input[4191]), .B(p_input[14191]), .Z(o[4191]) );
  AND U6456 ( .A(p_input[4190]), .B(p_input[14190]), .Z(o[4190]) );
  AND U6457 ( .A(p_input[418]), .B(p_input[10418]), .Z(o[418]) );
  AND U6458 ( .A(p_input[4189]), .B(p_input[14189]), .Z(o[4189]) );
  AND U6459 ( .A(p_input[4188]), .B(p_input[14188]), .Z(o[4188]) );
  AND U6460 ( .A(p_input[4187]), .B(p_input[14187]), .Z(o[4187]) );
  AND U6461 ( .A(p_input[4186]), .B(p_input[14186]), .Z(o[4186]) );
  AND U6462 ( .A(p_input[4185]), .B(p_input[14185]), .Z(o[4185]) );
  AND U6463 ( .A(p_input[4184]), .B(p_input[14184]), .Z(o[4184]) );
  AND U6464 ( .A(p_input[4183]), .B(p_input[14183]), .Z(o[4183]) );
  AND U6465 ( .A(p_input[4182]), .B(p_input[14182]), .Z(o[4182]) );
  AND U6466 ( .A(p_input[4181]), .B(p_input[14181]), .Z(o[4181]) );
  AND U6467 ( .A(p_input[4180]), .B(p_input[14180]), .Z(o[4180]) );
  AND U6468 ( .A(p_input[417]), .B(p_input[10417]), .Z(o[417]) );
  AND U6469 ( .A(p_input[4179]), .B(p_input[14179]), .Z(o[4179]) );
  AND U6470 ( .A(p_input[4178]), .B(p_input[14178]), .Z(o[4178]) );
  AND U6471 ( .A(p_input[4177]), .B(p_input[14177]), .Z(o[4177]) );
  AND U6472 ( .A(p_input[4176]), .B(p_input[14176]), .Z(o[4176]) );
  AND U6473 ( .A(p_input[4175]), .B(p_input[14175]), .Z(o[4175]) );
  AND U6474 ( .A(p_input[4174]), .B(p_input[14174]), .Z(o[4174]) );
  AND U6475 ( .A(p_input[4173]), .B(p_input[14173]), .Z(o[4173]) );
  AND U6476 ( .A(p_input[4172]), .B(p_input[14172]), .Z(o[4172]) );
  AND U6477 ( .A(p_input[4171]), .B(p_input[14171]), .Z(o[4171]) );
  AND U6478 ( .A(p_input[4170]), .B(p_input[14170]), .Z(o[4170]) );
  AND U6479 ( .A(p_input[416]), .B(p_input[10416]), .Z(o[416]) );
  AND U6480 ( .A(p_input[4169]), .B(p_input[14169]), .Z(o[4169]) );
  AND U6481 ( .A(p_input[4168]), .B(p_input[14168]), .Z(o[4168]) );
  AND U6482 ( .A(p_input[4167]), .B(p_input[14167]), .Z(o[4167]) );
  AND U6483 ( .A(p_input[4166]), .B(p_input[14166]), .Z(o[4166]) );
  AND U6484 ( .A(p_input[4165]), .B(p_input[14165]), .Z(o[4165]) );
  AND U6485 ( .A(p_input[4164]), .B(p_input[14164]), .Z(o[4164]) );
  AND U6486 ( .A(p_input[4163]), .B(p_input[14163]), .Z(o[4163]) );
  AND U6487 ( .A(p_input[4162]), .B(p_input[14162]), .Z(o[4162]) );
  AND U6488 ( .A(p_input[4161]), .B(p_input[14161]), .Z(o[4161]) );
  AND U6489 ( .A(p_input[4160]), .B(p_input[14160]), .Z(o[4160]) );
  AND U6490 ( .A(p_input[415]), .B(p_input[10415]), .Z(o[415]) );
  AND U6491 ( .A(p_input[4159]), .B(p_input[14159]), .Z(o[4159]) );
  AND U6492 ( .A(p_input[4158]), .B(p_input[14158]), .Z(o[4158]) );
  AND U6493 ( .A(p_input[4157]), .B(p_input[14157]), .Z(o[4157]) );
  AND U6494 ( .A(p_input[4156]), .B(p_input[14156]), .Z(o[4156]) );
  AND U6495 ( .A(p_input[4155]), .B(p_input[14155]), .Z(o[4155]) );
  AND U6496 ( .A(p_input[4154]), .B(p_input[14154]), .Z(o[4154]) );
  AND U6497 ( .A(p_input[4153]), .B(p_input[14153]), .Z(o[4153]) );
  AND U6498 ( .A(p_input[4152]), .B(p_input[14152]), .Z(o[4152]) );
  AND U6499 ( .A(p_input[4151]), .B(p_input[14151]), .Z(o[4151]) );
  AND U6500 ( .A(p_input[4150]), .B(p_input[14150]), .Z(o[4150]) );
  AND U6501 ( .A(p_input[414]), .B(p_input[10414]), .Z(o[414]) );
  AND U6502 ( .A(p_input[4149]), .B(p_input[14149]), .Z(o[4149]) );
  AND U6503 ( .A(p_input[4148]), .B(p_input[14148]), .Z(o[4148]) );
  AND U6504 ( .A(p_input[4147]), .B(p_input[14147]), .Z(o[4147]) );
  AND U6505 ( .A(p_input[4146]), .B(p_input[14146]), .Z(o[4146]) );
  AND U6506 ( .A(p_input[4145]), .B(p_input[14145]), .Z(o[4145]) );
  AND U6507 ( .A(p_input[4144]), .B(p_input[14144]), .Z(o[4144]) );
  AND U6508 ( .A(p_input[4143]), .B(p_input[14143]), .Z(o[4143]) );
  AND U6509 ( .A(p_input[4142]), .B(p_input[14142]), .Z(o[4142]) );
  AND U6510 ( .A(p_input[4141]), .B(p_input[14141]), .Z(o[4141]) );
  AND U6511 ( .A(p_input[4140]), .B(p_input[14140]), .Z(o[4140]) );
  AND U6512 ( .A(p_input[413]), .B(p_input[10413]), .Z(o[413]) );
  AND U6513 ( .A(p_input[4139]), .B(p_input[14139]), .Z(o[4139]) );
  AND U6514 ( .A(p_input[4138]), .B(p_input[14138]), .Z(o[4138]) );
  AND U6515 ( .A(p_input[4137]), .B(p_input[14137]), .Z(o[4137]) );
  AND U6516 ( .A(p_input[4136]), .B(p_input[14136]), .Z(o[4136]) );
  AND U6517 ( .A(p_input[4135]), .B(p_input[14135]), .Z(o[4135]) );
  AND U6518 ( .A(p_input[4134]), .B(p_input[14134]), .Z(o[4134]) );
  AND U6519 ( .A(p_input[4133]), .B(p_input[14133]), .Z(o[4133]) );
  AND U6520 ( .A(p_input[4132]), .B(p_input[14132]), .Z(o[4132]) );
  AND U6521 ( .A(p_input[4131]), .B(p_input[14131]), .Z(o[4131]) );
  AND U6522 ( .A(p_input[4130]), .B(p_input[14130]), .Z(o[4130]) );
  AND U6523 ( .A(p_input[412]), .B(p_input[10412]), .Z(o[412]) );
  AND U6524 ( .A(p_input[4129]), .B(p_input[14129]), .Z(o[4129]) );
  AND U6525 ( .A(p_input[4128]), .B(p_input[14128]), .Z(o[4128]) );
  AND U6526 ( .A(p_input[4127]), .B(p_input[14127]), .Z(o[4127]) );
  AND U6527 ( .A(p_input[4126]), .B(p_input[14126]), .Z(o[4126]) );
  AND U6528 ( .A(p_input[4125]), .B(p_input[14125]), .Z(o[4125]) );
  AND U6529 ( .A(p_input[4124]), .B(p_input[14124]), .Z(o[4124]) );
  AND U6530 ( .A(p_input[4123]), .B(p_input[14123]), .Z(o[4123]) );
  AND U6531 ( .A(p_input[4122]), .B(p_input[14122]), .Z(o[4122]) );
  AND U6532 ( .A(p_input[4121]), .B(p_input[14121]), .Z(o[4121]) );
  AND U6533 ( .A(p_input[4120]), .B(p_input[14120]), .Z(o[4120]) );
  AND U6534 ( .A(p_input[411]), .B(p_input[10411]), .Z(o[411]) );
  AND U6535 ( .A(p_input[4119]), .B(p_input[14119]), .Z(o[4119]) );
  AND U6536 ( .A(p_input[4118]), .B(p_input[14118]), .Z(o[4118]) );
  AND U6537 ( .A(p_input[4117]), .B(p_input[14117]), .Z(o[4117]) );
  AND U6538 ( .A(p_input[4116]), .B(p_input[14116]), .Z(o[4116]) );
  AND U6539 ( .A(p_input[4115]), .B(p_input[14115]), .Z(o[4115]) );
  AND U6540 ( .A(p_input[4114]), .B(p_input[14114]), .Z(o[4114]) );
  AND U6541 ( .A(p_input[4113]), .B(p_input[14113]), .Z(o[4113]) );
  AND U6542 ( .A(p_input[4112]), .B(p_input[14112]), .Z(o[4112]) );
  AND U6543 ( .A(p_input[4111]), .B(p_input[14111]), .Z(o[4111]) );
  AND U6544 ( .A(p_input[4110]), .B(p_input[14110]), .Z(o[4110]) );
  AND U6545 ( .A(p_input[410]), .B(p_input[10410]), .Z(o[410]) );
  AND U6546 ( .A(p_input[4109]), .B(p_input[14109]), .Z(o[4109]) );
  AND U6547 ( .A(p_input[4108]), .B(p_input[14108]), .Z(o[4108]) );
  AND U6548 ( .A(p_input[4107]), .B(p_input[14107]), .Z(o[4107]) );
  AND U6549 ( .A(p_input[4106]), .B(p_input[14106]), .Z(o[4106]) );
  AND U6550 ( .A(p_input[4105]), .B(p_input[14105]), .Z(o[4105]) );
  AND U6551 ( .A(p_input[4104]), .B(p_input[14104]), .Z(o[4104]) );
  AND U6552 ( .A(p_input[4103]), .B(p_input[14103]), .Z(o[4103]) );
  AND U6553 ( .A(p_input[4102]), .B(p_input[14102]), .Z(o[4102]) );
  AND U6554 ( .A(p_input[4101]), .B(p_input[14101]), .Z(o[4101]) );
  AND U6555 ( .A(p_input[4100]), .B(p_input[14100]), .Z(o[4100]) );
  AND U6556 ( .A(p_input[40]), .B(p_input[10040]), .Z(o[40]) );
  AND U6557 ( .A(p_input[409]), .B(p_input[10409]), .Z(o[409]) );
  AND U6558 ( .A(p_input[4099]), .B(p_input[14099]), .Z(o[4099]) );
  AND U6559 ( .A(p_input[4098]), .B(p_input[14098]), .Z(o[4098]) );
  AND U6560 ( .A(p_input[4097]), .B(p_input[14097]), .Z(o[4097]) );
  AND U6561 ( .A(p_input[4096]), .B(p_input[14096]), .Z(o[4096]) );
  AND U6562 ( .A(p_input[4095]), .B(p_input[14095]), .Z(o[4095]) );
  AND U6563 ( .A(p_input[4094]), .B(p_input[14094]), .Z(o[4094]) );
  AND U6564 ( .A(p_input[4093]), .B(p_input[14093]), .Z(o[4093]) );
  AND U6565 ( .A(p_input[4092]), .B(p_input[14092]), .Z(o[4092]) );
  AND U6566 ( .A(p_input[4091]), .B(p_input[14091]), .Z(o[4091]) );
  AND U6567 ( .A(p_input[4090]), .B(p_input[14090]), .Z(o[4090]) );
  AND U6568 ( .A(p_input[408]), .B(p_input[10408]), .Z(o[408]) );
  AND U6569 ( .A(p_input[4089]), .B(p_input[14089]), .Z(o[4089]) );
  AND U6570 ( .A(p_input[4088]), .B(p_input[14088]), .Z(o[4088]) );
  AND U6571 ( .A(p_input[4087]), .B(p_input[14087]), .Z(o[4087]) );
  AND U6572 ( .A(p_input[4086]), .B(p_input[14086]), .Z(o[4086]) );
  AND U6573 ( .A(p_input[4085]), .B(p_input[14085]), .Z(o[4085]) );
  AND U6574 ( .A(p_input[4084]), .B(p_input[14084]), .Z(o[4084]) );
  AND U6575 ( .A(p_input[4083]), .B(p_input[14083]), .Z(o[4083]) );
  AND U6576 ( .A(p_input[4082]), .B(p_input[14082]), .Z(o[4082]) );
  AND U6577 ( .A(p_input[4081]), .B(p_input[14081]), .Z(o[4081]) );
  AND U6578 ( .A(p_input[4080]), .B(p_input[14080]), .Z(o[4080]) );
  AND U6579 ( .A(p_input[407]), .B(p_input[10407]), .Z(o[407]) );
  AND U6580 ( .A(p_input[4079]), .B(p_input[14079]), .Z(o[4079]) );
  AND U6581 ( .A(p_input[4078]), .B(p_input[14078]), .Z(o[4078]) );
  AND U6582 ( .A(p_input[4077]), .B(p_input[14077]), .Z(o[4077]) );
  AND U6583 ( .A(p_input[4076]), .B(p_input[14076]), .Z(o[4076]) );
  AND U6584 ( .A(p_input[4075]), .B(p_input[14075]), .Z(o[4075]) );
  AND U6585 ( .A(p_input[4074]), .B(p_input[14074]), .Z(o[4074]) );
  AND U6586 ( .A(p_input[4073]), .B(p_input[14073]), .Z(o[4073]) );
  AND U6587 ( .A(p_input[4072]), .B(p_input[14072]), .Z(o[4072]) );
  AND U6588 ( .A(p_input[4071]), .B(p_input[14071]), .Z(o[4071]) );
  AND U6589 ( .A(p_input[4070]), .B(p_input[14070]), .Z(o[4070]) );
  AND U6590 ( .A(p_input[406]), .B(p_input[10406]), .Z(o[406]) );
  AND U6591 ( .A(p_input[4069]), .B(p_input[14069]), .Z(o[4069]) );
  AND U6592 ( .A(p_input[4068]), .B(p_input[14068]), .Z(o[4068]) );
  AND U6593 ( .A(p_input[4067]), .B(p_input[14067]), .Z(o[4067]) );
  AND U6594 ( .A(p_input[4066]), .B(p_input[14066]), .Z(o[4066]) );
  AND U6595 ( .A(p_input[4065]), .B(p_input[14065]), .Z(o[4065]) );
  AND U6596 ( .A(p_input[4064]), .B(p_input[14064]), .Z(o[4064]) );
  AND U6597 ( .A(p_input[4063]), .B(p_input[14063]), .Z(o[4063]) );
  AND U6598 ( .A(p_input[4062]), .B(p_input[14062]), .Z(o[4062]) );
  AND U6599 ( .A(p_input[4061]), .B(p_input[14061]), .Z(o[4061]) );
  AND U6600 ( .A(p_input[4060]), .B(p_input[14060]), .Z(o[4060]) );
  AND U6601 ( .A(p_input[405]), .B(p_input[10405]), .Z(o[405]) );
  AND U6602 ( .A(p_input[4059]), .B(p_input[14059]), .Z(o[4059]) );
  AND U6603 ( .A(p_input[4058]), .B(p_input[14058]), .Z(o[4058]) );
  AND U6604 ( .A(p_input[4057]), .B(p_input[14057]), .Z(o[4057]) );
  AND U6605 ( .A(p_input[4056]), .B(p_input[14056]), .Z(o[4056]) );
  AND U6606 ( .A(p_input[4055]), .B(p_input[14055]), .Z(o[4055]) );
  AND U6607 ( .A(p_input[4054]), .B(p_input[14054]), .Z(o[4054]) );
  AND U6608 ( .A(p_input[4053]), .B(p_input[14053]), .Z(o[4053]) );
  AND U6609 ( .A(p_input[4052]), .B(p_input[14052]), .Z(o[4052]) );
  AND U6610 ( .A(p_input[4051]), .B(p_input[14051]), .Z(o[4051]) );
  AND U6611 ( .A(p_input[4050]), .B(p_input[14050]), .Z(o[4050]) );
  AND U6612 ( .A(p_input[404]), .B(p_input[10404]), .Z(o[404]) );
  AND U6613 ( .A(p_input[4049]), .B(p_input[14049]), .Z(o[4049]) );
  AND U6614 ( .A(p_input[4048]), .B(p_input[14048]), .Z(o[4048]) );
  AND U6615 ( .A(p_input[4047]), .B(p_input[14047]), .Z(o[4047]) );
  AND U6616 ( .A(p_input[4046]), .B(p_input[14046]), .Z(o[4046]) );
  AND U6617 ( .A(p_input[4045]), .B(p_input[14045]), .Z(o[4045]) );
  AND U6618 ( .A(p_input[4044]), .B(p_input[14044]), .Z(o[4044]) );
  AND U6619 ( .A(p_input[4043]), .B(p_input[14043]), .Z(o[4043]) );
  AND U6620 ( .A(p_input[4042]), .B(p_input[14042]), .Z(o[4042]) );
  AND U6621 ( .A(p_input[4041]), .B(p_input[14041]), .Z(o[4041]) );
  AND U6622 ( .A(p_input[4040]), .B(p_input[14040]), .Z(o[4040]) );
  AND U6623 ( .A(p_input[403]), .B(p_input[10403]), .Z(o[403]) );
  AND U6624 ( .A(p_input[4039]), .B(p_input[14039]), .Z(o[4039]) );
  AND U6625 ( .A(p_input[4038]), .B(p_input[14038]), .Z(o[4038]) );
  AND U6626 ( .A(p_input[4037]), .B(p_input[14037]), .Z(o[4037]) );
  AND U6627 ( .A(p_input[4036]), .B(p_input[14036]), .Z(o[4036]) );
  AND U6628 ( .A(p_input[4035]), .B(p_input[14035]), .Z(o[4035]) );
  AND U6629 ( .A(p_input[4034]), .B(p_input[14034]), .Z(o[4034]) );
  AND U6630 ( .A(p_input[4033]), .B(p_input[14033]), .Z(o[4033]) );
  AND U6631 ( .A(p_input[4032]), .B(p_input[14032]), .Z(o[4032]) );
  AND U6632 ( .A(p_input[4031]), .B(p_input[14031]), .Z(o[4031]) );
  AND U6633 ( .A(p_input[4030]), .B(p_input[14030]), .Z(o[4030]) );
  AND U6634 ( .A(p_input[402]), .B(p_input[10402]), .Z(o[402]) );
  AND U6635 ( .A(p_input[4029]), .B(p_input[14029]), .Z(o[4029]) );
  AND U6636 ( .A(p_input[4028]), .B(p_input[14028]), .Z(o[4028]) );
  AND U6637 ( .A(p_input[4027]), .B(p_input[14027]), .Z(o[4027]) );
  AND U6638 ( .A(p_input[4026]), .B(p_input[14026]), .Z(o[4026]) );
  AND U6639 ( .A(p_input[4025]), .B(p_input[14025]), .Z(o[4025]) );
  AND U6640 ( .A(p_input[4024]), .B(p_input[14024]), .Z(o[4024]) );
  AND U6641 ( .A(p_input[4023]), .B(p_input[14023]), .Z(o[4023]) );
  AND U6642 ( .A(p_input[4022]), .B(p_input[14022]), .Z(o[4022]) );
  AND U6643 ( .A(p_input[4021]), .B(p_input[14021]), .Z(o[4021]) );
  AND U6644 ( .A(p_input[4020]), .B(p_input[14020]), .Z(o[4020]) );
  AND U6645 ( .A(p_input[401]), .B(p_input[10401]), .Z(o[401]) );
  AND U6646 ( .A(p_input[4019]), .B(p_input[14019]), .Z(o[4019]) );
  AND U6647 ( .A(p_input[4018]), .B(p_input[14018]), .Z(o[4018]) );
  AND U6648 ( .A(p_input[4017]), .B(p_input[14017]), .Z(o[4017]) );
  AND U6649 ( .A(p_input[4016]), .B(p_input[14016]), .Z(o[4016]) );
  AND U6650 ( .A(p_input[4015]), .B(p_input[14015]), .Z(o[4015]) );
  AND U6651 ( .A(p_input[4014]), .B(p_input[14014]), .Z(o[4014]) );
  AND U6652 ( .A(p_input[4013]), .B(p_input[14013]), .Z(o[4013]) );
  AND U6653 ( .A(p_input[4012]), .B(p_input[14012]), .Z(o[4012]) );
  AND U6654 ( .A(p_input[4011]), .B(p_input[14011]), .Z(o[4011]) );
  AND U6655 ( .A(p_input[4010]), .B(p_input[14010]), .Z(o[4010]) );
  AND U6656 ( .A(p_input[400]), .B(p_input[10400]), .Z(o[400]) );
  AND U6657 ( .A(p_input[4009]), .B(p_input[14009]), .Z(o[4009]) );
  AND U6658 ( .A(p_input[4008]), .B(p_input[14008]), .Z(o[4008]) );
  AND U6659 ( .A(p_input[4007]), .B(p_input[14007]), .Z(o[4007]) );
  AND U6660 ( .A(p_input[4006]), .B(p_input[14006]), .Z(o[4006]) );
  AND U6661 ( .A(p_input[4005]), .B(p_input[14005]), .Z(o[4005]) );
  AND U6662 ( .A(p_input[4004]), .B(p_input[14004]), .Z(o[4004]) );
  AND U6663 ( .A(p_input[4003]), .B(p_input[14003]), .Z(o[4003]) );
  AND U6664 ( .A(p_input[4002]), .B(p_input[14002]), .Z(o[4002]) );
  AND U6665 ( .A(p_input[4001]), .B(p_input[14001]), .Z(o[4001]) );
  AND U6666 ( .A(p_input[4000]), .B(p_input[14000]), .Z(o[4000]) );
  AND U6667 ( .A(p_input[3]), .B(p_input[10003]), .Z(o[3]) );
  AND U6668 ( .A(p_input[39]), .B(p_input[10039]), .Z(o[39]) );
  AND U6669 ( .A(p_input[399]), .B(p_input[10399]), .Z(o[399]) );
  AND U6670 ( .A(p_input[3999]), .B(p_input[13999]), .Z(o[3999]) );
  AND U6671 ( .A(p_input[3998]), .B(p_input[13998]), .Z(o[3998]) );
  AND U6672 ( .A(p_input[3997]), .B(p_input[13997]), .Z(o[3997]) );
  AND U6673 ( .A(p_input[3996]), .B(p_input[13996]), .Z(o[3996]) );
  AND U6674 ( .A(p_input[3995]), .B(p_input[13995]), .Z(o[3995]) );
  AND U6675 ( .A(p_input[3994]), .B(p_input[13994]), .Z(o[3994]) );
  AND U6676 ( .A(p_input[3993]), .B(p_input[13993]), .Z(o[3993]) );
  AND U6677 ( .A(p_input[3992]), .B(p_input[13992]), .Z(o[3992]) );
  AND U6678 ( .A(p_input[3991]), .B(p_input[13991]), .Z(o[3991]) );
  AND U6679 ( .A(p_input[3990]), .B(p_input[13990]), .Z(o[3990]) );
  AND U6680 ( .A(p_input[398]), .B(p_input[10398]), .Z(o[398]) );
  AND U6681 ( .A(p_input[3989]), .B(p_input[13989]), .Z(o[3989]) );
  AND U6682 ( .A(p_input[3988]), .B(p_input[13988]), .Z(o[3988]) );
  AND U6683 ( .A(p_input[3987]), .B(p_input[13987]), .Z(o[3987]) );
  AND U6684 ( .A(p_input[3986]), .B(p_input[13986]), .Z(o[3986]) );
  AND U6685 ( .A(p_input[3985]), .B(p_input[13985]), .Z(o[3985]) );
  AND U6686 ( .A(p_input[3984]), .B(p_input[13984]), .Z(o[3984]) );
  AND U6687 ( .A(p_input[3983]), .B(p_input[13983]), .Z(o[3983]) );
  AND U6688 ( .A(p_input[3982]), .B(p_input[13982]), .Z(o[3982]) );
  AND U6689 ( .A(p_input[3981]), .B(p_input[13981]), .Z(o[3981]) );
  AND U6690 ( .A(p_input[3980]), .B(p_input[13980]), .Z(o[3980]) );
  AND U6691 ( .A(p_input[397]), .B(p_input[10397]), .Z(o[397]) );
  AND U6692 ( .A(p_input[3979]), .B(p_input[13979]), .Z(o[3979]) );
  AND U6693 ( .A(p_input[3978]), .B(p_input[13978]), .Z(o[3978]) );
  AND U6694 ( .A(p_input[3977]), .B(p_input[13977]), .Z(o[3977]) );
  AND U6695 ( .A(p_input[3976]), .B(p_input[13976]), .Z(o[3976]) );
  AND U6696 ( .A(p_input[3975]), .B(p_input[13975]), .Z(o[3975]) );
  AND U6697 ( .A(p_input[3974]), .B(p_input[13974]), .Z(o[3974]) );
  AND U6698 ( .A(p_input[3973]), .B(p_input[13973]), .Z(o[3973]) );
  AND U6699 ( .A(p_input[3972]), .B(p_input[13972]), .Z(o[3972]) );
  AND U6700 ( .A(p_input[3971]), .B(p_input[13971]), .Z(o[3971]) );
  AND U6701 ( .A(p_input[3970]), .B(p_input[13970]), .Z(o[3970]) );
  AND U6702 ( .A(p_input[396]), .B(p_input[10396]), .Z(o[396]) );
  AND U6703 ( .A(p_input[3969]), .B(p_input[13969]), .Z(o[3969]) );
  AND U6704 ( .A(p_input[3968]), .B(p_input[13968]), .Z(o[3968]) );
  AND U6705 ( .A(p_input[3967]), .B(p_input[13967]), .Z(o[3967]) );
  AND U6706 ( .A(p_input[3966]), .B(p_input[13966]), .Z(o[3966]) );
  AND U6707 ( .A(p_input[3965]), .B(p_input[13965]), .Z(o[3965]) );
  AND U6708 ( .A(p_input[3964]), .B(p_input[13964]), .Z(o[3964]) );
  AND U6709 ( .A(p_input[3963]), .B(p_input[13963]), .Z(o[3963]) );
  AND U6710 ( .A(p_input[3962]), .B(p_input[13962]), .Z(o[3962]) );
  AND U6711 ( .A(p_input[3961]), .B(p_input[13961]), .Z(o[3961]) );
  AND U6712 ( .A(p_input[3960]), .B(p_input[13960]), .Z(o[3960]) );
  AND U6713 ( .A(p_input[395]), .B(p_input[10395]), .Z(o[395]) );
  AND U6714 ( .A(p_input[3959]), .B(p_input[13959]), .Z(o[3959]) );
  AND U6715 ( .A(p_input[3958]), .B(p_input[13958]), .Z(o[3958]) );
  AND U6716 ( .A(p_input[3957]), .B(p_input[13957]), .Z(o[3957]) );
  AND U6717 ( .A(p_input[3956]), .B(p_input[13956]), .Z(o[3956]) );
  AND U6718 ( .A(p_input[3955]), .B(p_input[13955]), .Z(o[3955]) );
  AND U6719 ( .A(p_input[3954]), .B(p_input[13954]), .Z(o[3954]) );
  AND U6720 ( .A(p_input[3953]), .B(p_input[13953]), .Z(o[3953]) );
  AND U6721 ( .A(p_input[3952]), .B(p_input[13952]), .Z(o[3952]) );
  AND U6722 ( .A(p_input[3951]), .B(p_input[13951]), .Z(o[3951]) );
  AND U6723 ( .A(p_input[3950]), .B(p_input[13950]), .Z(o[3950]) );
  AND U6724 ( .A(p_input[394]), .B(p_input[10394]), .Z(o[394]) );
  AND U6725 ( .A(p_input[3949]), .B(p_input[13949]), .Z(o[3949]) );
  AND U6726 ( .A(p_input[3948]), .B(p_input[13948]), .Z(o[3948]) );
  AND U6727 ( .A(p_input[3947]), .B(p_input[13947]), .Z(o[3947]) );
  AND U6728 ( .A(p_input[3946]), .B(p_input[13946]), .Z(o[3946]) );
  AND U6729 ( .A(p_input[3945]), .B(p_input[13945]), .Z(o[3945]) );
  AND U6730 ( .A(p_input[3944]), .B(p_input[13944]), .Z(o[3944]) );
  AND U6731 ( .A(p_input[3943]), .B(p_input[13943]), .Z(o[3943]) );
  AND U6732 ( .A(p_input[3942]), .B(p_input[13942]), .Z(o[3942]) );
  AND U6733 ( .A(p_input[3941]), .B(p_input[13941]), .Z(o[3941]) );
  AND U6734 ( .A(p_input[3940]), .B(p_input[13940]), .Z(o[3940]) );
  AND U6735 ( .A(p_input[393]), .B(p_input[10393]), .Z(o[393]) );
  AND U6736 ( .A(p_input[3939]), .B(p_input[13939]), .Z(o[3939]) );
  AND U6737 ( .A(p_input[3938]), .B(p_input[13938]), .Z(o[3938]) );
  AND U6738 ( .A(p_input[3937]), .B(p_input[13937]), .Z(o[3937]) );
  AND U6739 ( .A(p_input[3936]), .B(p_input[13936]), .Z(o[3936]) );
  AND U6740 ( .A(p_input[3935]), .B(p_input[13935]), .Z(o[3935]) );
  AND U6741 ( .A(p_input[3934]), .B(p_input[13934]), .Z(o[3934]) );
  AND U6742 ( .A(p_input[3933]), .B(p_input[13933]), .Z(o[3933]) );
  AND U6743 ( .A(p_input[3932]), .B(p_input[13932]), .Z(o[3932]) );
  AND U6744 ( .A(p_input[3931]), .B(p_input[13931]), .Z(o[3931]) );
  AND U6745 ( .A(p_input[3930]), .B(p_input[13930]), .Z(o[3930]) );
  AND U6746 ( .A(p_input[392]), .B(p_input[10392]), .Z(o[392]) );
  AND U6747 ( .A(p_input[3929]), .B(p_input[13929]), .Z(o[3929]) );
  AND U6748 ( .A(p_input[3928]), .B(p_input[13928]), .Z(o[3928]) );
  AND U6749 ( .A(p_input[3927]), .B(p_input[13927]), .Z(o[3927]) );
  AND U6750 ( .A(p_input[3926]), .B(p_input[13926]), .Z(o[3926]) );
  AND U6751 ( .A(p_input[3925]), .B(p_input[13925]), .Z(o[3925]) );
  AND U6752 ( .A(p_input[3924]), .B(p_input[13924]), .Z(o[3924]) );
  AND U6753 ( .A(p_input[3923]), .B(p_input[13923]), .Z(o[3923]) );
  AND U6754 ( .A(p_input[3922]), .B(p_input[13922]), .Z(o[3922]) );
  AND U6755 ( .A(p_input[3921]), .B(p_input[13921]), .Z(o[3921]) );
  AND U6756 ( .A(p_input[3920]), .B(p_input[13920]), .Z(o[3920]) );
  AND U6757 ( .A(p_input[391]), .B(p_input[10391]), .Z(o[391]) );
  AND U6758 ( .A(p_input[3919]), .B(p_input[13919]), .Z(o[3919]) );
  AND U6759 ( .A(p_input[3918]), .B(p_input[13918]), .Z(o[3918]) );
  AND U6760 ( .A(p_input[3917]), .B(p_input[13917]), .Z(o[3917]) );
  AND U6761 ( .A(p_input[3916]), .B(p_input[13916]), .Z(o[3916]) );
  AND U6762 ( .A(p_input[3915]), .B(p_input[13915]), .Z(o[3915]) );
  AND U6763 ( .A(p_input[3914]), .B(p_input[13914]), .Z(o[3914]) );
  AND U6764 ( .A(p_input[3913]), .B(p_input[13913]), .Z(o[3913]) );
  AND U6765 ( .A(p_input[3912]), .B(p_input[13912]), .Z(o[3912]) );
  AND U6766 ( .A(p_input[3911]), .B(p_input[13911]), .Z(o[3911]) );
  AND U6767 ( .A(p_input[3910]), .B(p_input[13910]), .Z(o[3910]) );
  AND U6768 ( .A(p_input[390]), .B(p_input[10390]), .Z(o[390]) );
  AND U6769 ( .A(p_input[3909]), .B(p_input[13909]), .Z(o[3909]) );
  AND U6770 ( .A(p_input[3908]), .B(p_input[13908]), .Z(o[3908]) );
  AND U6771 ( .A(p_input[3907]), .B(p_input[13907]), .Z(o[3907]) );
  AND U6772 ( .A(p_input[3906]), .B(p_input[13906]), .Z(o[3906]) );
  AND U6773 ( .A(p_input[3905]), .B(p_input[13905]), .Z(o[3905]) );
  AND U6774 ( .A(p_input[3904]), .B(p_input[13904]), .Z(o[3904]) );
  AND U6775 ( .A(p_input[3903]), .B(p_input[13903]), .Z(o[3903]) );
  AND U6776 ( .A(p_input[3902]), .B(p_input[13902]), .Z(o[3902]) );
  AND U6777 ( .A(p_input[3901]), .B(p_input[13901]), .Z(o[3901]) );
  AND U6778 ( .A(p_input[3900]), .B(p_input[13900]), .Z(o[3900]) );
  AND U6779 ( .A(p_input[38]), .B(p_input[10038]), .Z(o[38]) );
  AND U6780 ( .A(p_input[389]), .B(p_input[10389]), .Z(o[389]) );
  AND U6781 ( .A(p_input[3899]), .B(p_input[13899]), .Z(o[3899]) );
  AND U6782 ( .A(p_input[3898]), .B(p_input[13898]), .Z(o[3898]) );
  AND U6783 ( .A(p_input[3897]), .B(p_input[13897]), .Z(o[3897]) );
  AND U6784 ( .A(p_input[3896]), .B(p_input[13896]), .Z(o[3896]) );
  AND U6785 ( .A(p_input[3895]), .B(p_input[13895]), .Z(o[3895]) );
  AND U6786 ( .A(p_input[3894]), .B(p_input[13894]), .Z(o[3894]) );
  AND U6787 ( .A(p_input[3893]), .B(p_input[13893]), .Z(o[3893]) );
  AND U6788 ( .A(p_input[3892]), .B(p_input[13892]), .Z(o[3892]) );
  AND U6789 ( .A(p_input[3891]), .B(p_input[13891]), .Z(o[3891]) );
  AND U6790 ( .A(p_input[3890]), .B(p_input[13890]), .Z(o[3890]) );
  AND U6791 ( .A(p_input[388]), .B(p_input[10388]), .Z(o[388]) );
  AND U6792 ( .A(p_input[3889]), .B(p_input[13889]), .Z(o[3889]) );
  AND U6793 ( .A(p_input[3888]), .B(p_input[13888]), .Z(o[3888]) );
  AND U6794 ( .A(p_input[3887]), .B(p_input[13887]), .Z(o[3887]) );
  AND U6795 ( .A(p_input[3886]), .B(p_input[13886]), .Z(o[3886]) );
  AND U6796 ( .A(p_input[3885]), .B(p_input[13885]), .Z(o[3885]) );
  AND U6797 ( .A(p_input[3884]), .B(p_input[13884]), .Z(o[3884]) );
  AND U6798 ( .A(p_input[3883]), .B(p_input[13883]), .Z(o[3883]) );
  AND U6799 ( .A(p_input[3882]), .B(p_input[13882]), .Z(o[3882]) );
  AND U6800 ( .A(p_input[3881]), .B(p_input[13881]), .Z(o[3881]) );
  AND U6801 ( .A(p_input[3880]), .B(p_input[13880]), .Z(o[3880]) );
  AND U6802 ( .A(p_input[387]), .B(p_input[10387]), .Z(o[387]) );
  AND U6803 ( .A(p_input[3879]), .B(p_input[13879]), .Z(o[3879]) );
  AND U6804 ( .A(p_input[3878]), .B(p_input[13878]), .Z(o[3878]) );
  AND U6805 ( .A(p_input[3877]), .B(p_input[13877]), .Z(o[3877]) );
  AND U6806 ( .A(p_input[3876]), .B(p_input[13876]), .Z(o[3876]) );
  AND U6807 ( .A(p_input[3875]), .B(p_input[13875]), .Z(o[3875]) );
  AND U6808 ( .A(p_input[3874]), .B(p_input[13874]), .Z(o[3874]) );
  AND U6809 ( .A(p_input[3873]), .B(p_input[13873]), .Z(o[3873]) );
  AND U6810 ( .A(p_input[3872]), .B(p_input[13872]), .Z(o[3872]) );
  AND U6811 ( .A(p_input[3871]), .B(p_input[13871]), .Z(o[3871]) );
  AND U6812 ( .A(p_input[3870]), .B(p_input[13870]), .Z(o[3870]) );
  AND U6813 ( .A(p_input[386]), .B(p_input[10386]), .Z(o[386]) );
  AND U6814 ( .A(p_input[3869]), .B(p_input[13869]), .Z(o[3869]) );
  AND U6815 ( .A(p_input[3868]), .B(p_input[13868]), .Z(o[3868]) );
  AND U6816 ( .A(p_input[3867]), .B(p_input[13867]), .Z(o[3867]) );
  AND U6817 ( .A(p_input[3866]), .B(p_input[13866]), .Z(o[3866]) );
  AND U6818 ( .A(p_input[3865]), .B(p_input[13865]), .Z(o[3865]) );
  AND U6819 ( .A(p_input[3864]), .B(p_input[13864]), .Z(o[3864]) );
  AND U6820 ( .A(p_input[3863]), .B(p_input[13863]), .Z(o[3863]) );
  AND U6821 ( .A(p_input[3862]), .B(p_input[13862]), .Z(o[3862]) );
  AND U6822 ( .A(p_input[3861]), .B(p_input[13861]), .Z(o[3861]) );
  AND U6823 ( .A(p_input[3860]), .B(p_input[13860]), .Z(o[3860]) );
  AND U6824 ( .A(p_input[385]), .B(p_input[10385]), .Z(o[385]) );
  AND U6825 ( .A(p_input[3859]), .B(p_input[13859]), .Z(o[3859]) );
  AND U6826 ( .A(p_input[3858]), .B(p_input[13858]), .Z(o[3858]) );
  AND U6827 ( .A(p_input[3857]), .B(p_input[13857]), .Z(o[3857]) );
  AND U6828 ( .A(p_input[3856]), .B(p_input[13856]), .Z(o[3856]) );
  AND U6829 ( .A(p_input[3855]), .B(p_input[13855]), .Z(o[3855]) );
  AND U6830 ( .A(p_input[3854]), .B(p_input[13854]), .Z(o[3854]) );
  AND U6831 ( .A(p_input[3853]), .B(p_input[13853]), .Z(o[3853]) );
  AND U6832 ( .A(p_input[3852]), .B(p_input[13852]), .Z(o[3852]) );
  AND U6833 ( .A(p_input[3851]), .B(p_input[13851]), .Z(o[3851]) );
  AND U6834 ( .A(p_input[3850]), .B(p_input[13850]), .Z(o[3850]) );
  AND U6835 ( .A(p_input[384]), .B(p_input[10384]), .Z(o[384]) );
  AND U6836 ( .A(p_input[3849]), .B(p_input[13849]), .Z(o[3849]) );
  AND U6837 ( .A(p_input[3848]), .B(p_input[13848]), .Z(o[3848]) );
  AND U6838 ( .A(p_input[3847]), .B(p_input[13847]), .Z(o[3847]) );
  AND U6839 ( .A(p_input[3846]), .B(p_input[13846]), .Z(o[3846]) );
  AND U6840 ( .A(p_input[3845]), .B(p_input[13845]), .Z(o[3845]) );
  AND U6841 ( .A(p_input[3844]), .B(p_input[13844]), .Z(o[3844]) );
  AND U6842 ( .A(p_input[3843]), .B(p_input[13843]), .Z(o[3843]) );
  AND U6843 ( .A(p_input[3842]), .B(p_input[13842]), .Z(o[3842]) );
  AND U6844 ( .A(p_input[3841]), .B(p_input[13841]), .Z(o[3841]) );
  AND U6845 ( .A(p_input[3840]), .B(p_input[13840]), .Z(o[3840]) );
  AND U6846 ( .A(p_input[383]), .B(p_input[10383]), .Z(o[383]) );
  AND U6847 ( .A(p_input[3839]), .B(p_input[13839]), .Z(o[3839]) );
  AND U6848 ( .A(p_input[3838]), .B(p_input[13838]), .Z(o[3838]) );
  AND U6849 ( .A(p_input[3837]), .B(p_input[13837]), .Z(o[3837]) );
  AND U6850 ( .A(p_input[3836]), .B(p_input[13836]), .Z(o[3836]) );
  AND U6851 ( .A(p_input[3835]), .B(p_input[13835]), .Z(o[3835]) );
  AND U6852 ( .A(p_input[3834]), .B(p_input[13834]), .Z(o[3834]) );
  AND U6853 ( .A(p_input[3833]), .B(p_input[13833]), .Z(o[3833]) );
  AND U6854 ( .A(p_input[3832]), .B(p_input[13832]), .Z(o[3832]) );
  AND U6855 ( .A(p_input[3831]), .B(p_input[13831]), .Z(o[3831]) );
  AND U6856 ( .A(p_input[3830]), .B(p_input[13830]), .Z(o[3830]) );
  AND U6857 ( .A(p_input[382]), .B(p_input[10382]), .Z(o[382]) );
  AND U6858 ( .A(p_input[3829]), .B(p_input[13829]), .Z(o[3829]) );
  AND U6859 ( .A(p_input[3828]), .B(p_input[13828]), .Z(o[3828]) );
  AND U6860 ( .A(p_input[3827]), .B(p_input[13827]), .Z(o[3827]) );
  AND U6861 ( .A(p_input[3826]), .B(p_input[13826]), .Z(o[3826]) );
  AND U6862 ( .A(p_input[3825]), .B(p_input[13825]), .Z(o[3825]) );
  AND U6863 ( .A(p_input[3824]), .B(p_input[13824]), .Z(o[3824]) );
  AND U6864 ( .A(p_input[3823]), .B(p_input[13823]), .Z(o[3823]) );
  AND U6865 ( .A(p_input[3822]), .B(p_input[13822]), .Z(o[3822]) );
  AND U6866 ( .A(p_input[3821]), .B(p_input[13821]), .Z(o[3821]) );
  AND U6867 ( .A(p_input[3820]), .B(p_input[13820]), .Z(o[3820]) );
  AND U6868 ( .A(p_input[381]), .B(p_input[10381]), .Z(o[381]) );
  AND U6869 ( .A(p_input[3819]), .B(p_input[13819]), .Z(o[3819]) );
  AND U6870 ( .A(p_input[3818]), .B(p_input[13818]), .Z(o[3818]) );
  AND U6871 ( .A(p_input[3817]), .B(p_input[13817]), .Z(o[3817]) );
  AND U6872 ( .A(p_input[3816]), .B(p_input[13816]), .Z(o[3816]) );
  AND U6873 ( .A(p_input[3815]), .B(p_input[13815]), .Z(o[3815]) );
  AND U6874 ( .A(p_input[3814]), .B(p_input[13814]), .Z(o[3814]) );
  AND U6875 ( .A(p_input[3813]), .B(p_input[13813]), .Z(o[3813]) );
  AND U6876 ( .A(p_input[3812]), .B(p_input[13812]), .Z(o[3812]) );
  AND U6877 ( .A(p_input[3811]), .B(p_input[13811]), .Z(o[3811]) );
  AND U6878 ( .A(p_input[3810]), .B(p_input[13810]), .Z(o[3810]) );
  AND U6879 ( .A(p_input[380]), .B(p_input[10380]), .Z(o[380]) );
  AND U6880 ( .A(p_input[3809]), .B(p_input[13809]), .Z(o[3809]) );
  AND U6881 ( .A(p_input[3808]), .B(p_input[13808]), .Z(o[3808]) );
  AND U6882 ( .A(p_input[3807]), .B(p_input[13807]), .Z(o[3807]) );
  AND U6883 ( .A(p_input[3806]), .B(p_input[13806]), .Z(o[3806]) );
  AND U6884 ( .A(p_input[3805]), .B(p_input[13805]), .Z(o[3805]) );
  AND U6885 ( .A(p_input[3804]), .B(p_input[13804]), .Z(o[3804]) );
  AND U6886 ( .A(p_input[3803]), .B(p_input[13803]), .Z(o[3803]) );
  AND U6887 ( .A(p_input[3802]), .B(p_input[13802]), .Z(o[3802]) );
  AND U6888 ( .A(p_input[3801]), .B(p_input[13801]), .Z(o[3801]) );
  AND U6889 ( .A(p_input[3800]), .B(p_input[13800]), .Z(o[3800]) );
  AND U6890 ( .A(p_input[37]), .B(p_input[10037]), .Z(o[37]) );
  AND U6891 ( .A(p_input[379]), .B(p_input[10379]), .Z(o[379]) );
  AND U6892 ( .A(p_input[3799]), .B(p_input[13799]), .Z(o[3799]) );
  AND U6893 ( .A(p_input[3798]), .B(p_input[13798]), .Z(o[3798]) );
  AND U6894 ( .A(p_input[3797]), .B(p_input[13797]), .Z(o[3797]) );
  AND U6895 ( .A(p_input[3796]), .B(p_input[13796]), .Z(o[3796]) );
  AND U6896 ( .A(p_input[3795]), .B(p_input[13795]), .Z(o[3795]) );
  AND U6897 ( .A(p_input[3794]), .B(p_input[13794]), .Z(o[3794]) );
  AND U6898 ( .A(p_input[3793]), .B(p_input[13793]), .Z(o[3793]) );
  AND U6899 ( .A(p_input[3792]), .B(p_input[13792]), .Z(o[3792]) );
  AND U6900 ( .A(p_input[3791]), .B(p_input[13791]), .Z(o[3791]) );
  AND U6901 ( .A(p_input[3790]), .B(p_input[13790]), .Z(o[3790]) );
  AND U6902 ( .A(p_input[378]), .B(p_input[10378]), .Z(o[378]) );
  AND U6903 ( .A(p_input[3789]), .B(p_input[13789]), .Z(o[3789]) );
  AND U6904 ( .A(p_input[3788]), .B(p_input[13788]), .Z(o[3788]) );
  AND U6905 ( .A(p_input[3787]), .B(p_input[13787]), .Z(o[3787]) );
  AND U6906 ( .A(p_input[3786]), .B(p_input[13786]), .Z(o[3786]) );
  AND U6907 ( .A(p_input[3785]), .B(p_input[13785]), .Z(o[3785]) );
  AND U6908 ( .A(p_input[3784]), .B(p_input[13784]), .Z(o[3784]) );
  AND U6909 ( .A(p_input[3783]), .B(p_input[13783]), .Z(o[3783]) );
  AND U6910 ( .A(p_input[3782]), .B(p_input[13782]), .Z(o[3782]) );
  AND U6911 ( .A(p_input[3781]), .B(p_input[13781]), .Z(o[3781]) );
  AND U6912 ( .A(p_input[3780]), .B(p_input[13780]), .Z(o[3780]) );
  AND U6913 ( .A(p_input[377]), .B(p_input[10377]), .Z(o[377]) );
  AND U6914 ( .A(p_input[3779]), .B(p_input[13779]), .Z(o[3779]) );
  AND U6915 ( .A(p_input[3778]), .B(p_input[13778]), .Z(o[3778]) );
  AND U6916 ( .A(p_input[3777]), .B(p_input[13777]), .Z(o[3777]) );
  AND U6917 ( .A(p_input[3776]), .B(p_input[13776]), .Z(o[3776]) );
  AND U6918 ( .A(p_input[3775]), .B(p_input[13775]), .Z(o[3775]) );
  AND U6919 ( .A(p_input[3774]), .B(p_input[13774]), .Z(o[3774]) );
  AND U6920 ( .A(p_input[3773]), .B(p_input[13773]), .Z(o[3773]) );
  AND U6921 ( .A(p_input[3772]), .B(p_input[13772]), .Z(o[3772]) );
  AND U6922 ( .A(p_input[3771]), .B(p_input[13771]), .Z(o[3771]) );
  AND U6923 ( .A(p_input[3770]), .B(p_input[13770]), .Z(o[3770]) );
  AND U6924 ( .A(p_input[376]), .B(p_input[10376]), .Z(o[376]) );
  AND U6925 ( .A(p_input[3769]), .B(p_input[13769]), .Z(o[3769]) );
  AND U6926 ( .A(p_input[3768]), .B(p_input[13768]), .Z(o[3768]) );
  AND U6927 ( .A(p_input[3767]), .B(p_input[13767]), .Z(o[3767]) );
  AND U6928 ( .A(p_input[3766]), .B(p_input[13766]), .Z(o[3766]) );
  AND U6929 ( .A(p_input[3765]), .B(p_input[13765]), .Z(o[3765]) );
  AND U6930 ( .A(p_input[3764]), .B(p_input[13764]), .Z(o[3764]) );
  AND U6931 ( .A(p_input[3763]), .B(p_input[13763]), .Z(o[3763]) );
  AND U6932 ( .A(p_input[3762]), .B(p_input[13762]), .Z(o[3762]) );
  AND U6933 ( .A(p_input[3761]), .B(p_input[13761]), .Z(o[3761]) );
  AND U6934 ( .A(p_input[3760]), .B(p_input[13760]), .Z(o[3760]) );
  AND U6935 ( .A(p_input[375]), .B(p_input[10375]), .Z(o[375]) );
  AND U6936 ( .A(p_input[3759]), .B(p_input[13759]), .Z(o[3759]) );
  AND U6937 ( .A(p_input[3758]), .B(p_input[13758]), .Z(o[3758]) );
  AND U6938 ( .A(p_input[3757]), .B(p_input[13757]), .Z(o[3757]) );
  AND U6939 ( .A(p_input[3756]), .B(p_input[13756]), .Z(o[3756]) );
  AND U6940 ( .A(p_input[3755]), .B(p_input[13755]), .Z(o[3755]) );
  AND U6941 ( .A(p_input[3754]), .B(p_input[13754]), .Z(o[3754]) );
  AND U6942 ( .A(p_input[3753]), .B(p_input[13753]), .Z(o[3753]) );
  AND U6943 ( .A(p_input[3752]), .B(p_input[13752]), .Z(o[3752]) );
  AND U6944 ( .A(p_input[3751]), .B(p_input[13751]), .Z(o[3751]) );
  AND U6945 ( .A(p_input[3750]), .B(p_input[13750]), .Z(o[3750]) );
  AND U6946 ( .A(p_input[374]), .B(p_input[10374]), .Z(o[374]) );
  AND U6947 ( .A(p_input[3749]), .B(p_input[13749]), .Z(o[3749]) );
  AND U6948 ( .A(p_input[3748]), .B(p_input[13748]), .Z(o[3748]) );
  AND U6949 ( .A(p_input[3747]), .B(p_input[13747]), .Z(o[3747]) );
  AND U6950 ( .A(p_input[3746]), .B(p_input[13746]), .Z(o[3746]) );
  AND U6951 ( .A(p_input[3745]), .B(p_input[13745]), .Z(o[3745]) );
  AND U6952 ( .A(p_input[3744]), .B(p_input[13744]), .Z(o[3744]) );
  AND U6953 ( .A(p_input[3743]), .B(p_input[13743]), .Z(o[3743]) );
  AND U6954 ( .A(p_input[3742]), .B(p_input[13742]), .Z(o[3742]) );
  AND U6955 ( .A(p_input[3741]), .B(p_input[13741]), .Z(o[3741]) );
  AND U6956 ( .A(p_input[3740]), .B(p_input[13740]), .Z(o[3740]) );
  AND U6957 ( .A(p_input[373]), .B(p_input[10373]), .Z(o[373]) );
  AND U6958 ( .A(p_input[3739]), .B(p_input[13739]), .Z(o[3739]) );
  AND U6959 ( .A(p_input[3738]), .B(p_input[13738]), .Z(o[3738]) );
  AND U6960 ( .A(p_input[3737]), .B(p_input[13737]), .Z(o[3737]) );
  AND U6961 ( .A(p_input[3736]), .B(p_input[13736]), .Z(o[3736]) );
  AND U6962 ( .A(p_input[3735]), .B(p_input[13735]), .Z(o[3735]) );
  AND U6963 ( .A(p_input[3734]), .B(p_input[13734]), .Z(o[3734]) );
  AND U6964 ( .A(p_input[3733]), .B(p_input[13733]), .Z(o[3733]) );
  AND U6965 ( .A(p_input[3732]), .B(p_input[13732]), .Z(o[3732]) );
  AND U6966 ( .A(p_input[3731]), .B(p_input[13731]), .Z(o[3731]) );
  AND U6967 ( .A(p_input[3730]), .B(p_input[13730]), .Z(o[3730]) );
  AND U6968 ( .A(p_input[372]), .B(p_input[10372]), .Z(o[372]) );
  AND U6969 ( .A(p_input[3729]), .B(p_input[13729]), .Z(o[3729]) );
  AND U6970 ( .A(p_input[3728]), .B(p_input[13728]), .Z(o[3728]) );
  AND U6971 ( .A(p_input[3727]), .B(p_input[13727]), .Z(o[3727]) );
  AND U6972 ( .A(p_input[3726]), .B(p_input[13726]), .Z(o[3726]) );
  AND U6973 ( .A(p_input[3725]), .B(p_input[13725]), .Z(o[3725]) );
  AND U6974 ( .A(p_input[3724]), .B(p_input[13724]), .Z(o[3724]) );
  AND U6975 ( .A(p_input[3723]), .B(p_input[13723]), .Z(o[3723]) );
  AND U6976 ( .A(p_input[3722]), .B(p_input[13722]), .Z(o[3722]) );
  AND U6977 ( .A(p_input[3721]), .B(p_input[13721]), .Z(o[3721]) );
  AND U6978 ( .A(p_input[3720]), .B(p_input[13720]), .Z(o[3720]) );
  AND U6979 ( .A(p_input[371]), .B(p_input[10371]), .Z(o[371]) );
  AND U6980 ( .A(p_input[3719]), .B(p_input[13719]), .Z(o[3719]) );
  AND U6981 ( .A(p_input[3718]), .B(p_input[13718]), .Z(o[3718]) );
  AND U6982 ( .A(p_input[3717]), .B(p_input[13717]), .Z(o[3717]) );
  AND U6983 ( .A(p_input[3716]), .B(p_input[13716]), .Z(o[3716]) );
  AND U6984 ( .A(p_input[3715]), .B(p_input[13715]), .Z(o[3715]) );
  AND U6985 ( .A(p_input[3714]), .B(p_input[13714]), .Z(o[3714]) );
  AND U6986 ( .A(p_input[3713]), .B(p_input[13713]), .Z(o[3713]) );
  AND U6987 ( .A(p_input[3712]), .B(p_input[13712]), .Z(o[3712]) );
  AND U6988 ( .A(p_input[3711]), .B(p_input[13711]), .Z(o[3711]) );
  AND U6989 ( .A(p_input[3710]), .B(p_input[13710]), .Z(o[3710]) );
  AND U6990 ( .A(p_input[370]), .B(p_input[10370]), .Z(o[370]) );
  AND U6991 ( .A(p_input[3709]), .B(p_input[13709]), .Z(o[3709]) );
  AND U6992 ( .A(p_input[3708]), .B(p_input[13708]), .Z(o[3708]) );
  AND U6993 ( .A(p_input[3707]), .B(p_input[13707]), .Z(o[3707]) );
  AND U6994 ( .A(p_input[3706]), .B(p_input[13706]), .Z(o[3706]) );
  AND U6995 ( .A(p_input[3705]), .B(p_input[13705]), .Z(o[3705]) );
  AND U6996 ( .A(p_input[3704]), .B(p_input[13704]), .Z(o[3704]) );
  AND U6997 ( .A(p_input[3703]), .B(p_input[13703]), .Z(o[3703]) );
  AND U6998 ( .A(p_input[3702]), .B(p_input[13702]), .Z(o[3702]) );
  AND U6999 ( .A(p_input[3701]), .B(p_input[13701]), .Z(o[3701]) );
  AND U7000 ( .A(p_input[3700]), .B(p_input[13700]), .Z(o[3700]) );
  AND U7001 ( .A(p_input[36]), .B(p_input[10036]), .Z(o[36]) );
  AND U7002 ( .A(p_input[369]), .B(p_input[10369]), .Z(o[369]) );
  AND U7003 ( .A(p_input[3699]), .B(p_input[13699]), .Z(o[3699]) );
  AND U7004 ( .A(p_input[3698]), .B(p_input[13698]), .Z(o[3698]) );
  AND U7005 ( .A(p_input[3697]), .B(p_input[13697]), .Z(o[3697]) );
  AND U7006 ( .A(p_input[3696]), .B(p_input[13696]), .Z(o[3696]) );
  AND U7007 ( .A(p_input[3695]), .B(p_input[13695]), .Z(o[3695]) );
  AND U7008 ( .A(p_input[3694]), .B(p_input[13694]), .Z(o[3694]) );
  AND U7009 ( .A(p_input[3693]), .B(p_input[13693]), .Z(o[3693]) );
  AND U7010 ( .A(p_input[3692]), .B(p_input[13692]), .Z(o[3692]) );
  AND U7011 ( .A(p_input[3691]), .B(p_input[13691]), .Z(o[3691]) );
  AND U7012 ( .A(p_input[3690]), .B(p_input[13690]), .Z(o[3690]) );
  AND U7013 ( .A(p_input[368]), .B(p_input[10368]), .Z(o[368]) );
  AND U7014 ( .A(p_input[3689]), .B(p_input[13689]), .Z(o[3689]) );
  AND U7015 ( .A(p_input[3688]), .B(p_input[13688]), .Z(o[3688]) );
  AND U7016 ( .A(p_input[3687]), .B(p_input[13687]), .Z(o[3687]) );
  AND U7017 ( .A(p_input[3686]), .B(p_input[13686]), .Z(o[3686]) );
  AND U7018 ( .A(p_input[3685]), .B(p_input[13685]), .Z(o[3685]) );
  AND U7019 ( .A(p_input[3684]), .B(p_input[13684]), .Z(o[3684]) );
  AND U7020 ( .A(p_input[3683]), .B(p_input[13683]), .Z(o[3683]) );
  AND U7021 ( .A(p_input[3682]), .B(p_input[13682]), .Z(o[3682]) );
  AND U7022 ( .A(p_input[3681]), .B(p_input[13681]), .Z(o[3681]) );
  AND U7023 ( .A(p_input[3680]), .B(p_input[13680]), .Z(o[3680]) );
  AND U7024 ( .A(p_input[367]), .B(p_input[10367]), .Z(o[367]) );
  AND U7025 ( .A(p_input[3679]), .B(p_input[13679]), .Z(o[3679]) );
  AND U7026 ( .A(p_input[3678]), .B(p_input[13678]), .Z(o[3678]) );
  AND U7027 ( .A(p_input[3677]), .B(p_input[13677]), .Z(o[3677]) );
  AND U7028 ( .A(p_input[3676]), .B(p_input[13676]), .Z(o[3676]) );
  AND U7029 ( .A(p_input[3675]), .B(p_input[13675]), .Z(o[3675]) );
  AND U7030 ( .A(p_input[3674]), .B(p_input[13674]), .Z(o[3674]) );
  AND U7031 ( .A(p_input[3673]), .B(p_input[13673]), .Z(o[3673]) );
  AND U7032 ( .A(p_input[3672]), .B(p_input[13672]), .Z(o[3672]) );
  AND U7033 ( .A(p_input[3671]), .B(p_input[13671]), .Z(o[3671]) );
  AND U7034 ( .A(p_input[3670]), .B(p_input[13670]), .Z(o[3670]) );
  AND U7035 ( .A(p_input[366]), .B(p_input[10366]), .Z(o[366]) );
  AND U7036 ( .A(p_input[3669]), .B(p_input[13669]), .Z(o[3669]) );
  AND U7037 ( .A(p_input[3668]), .B(p_input[13668]), .Z(o[3668]) );
  AND U7038 ( .A(p_input[3667]), .B(p_input[13667]), .Z(o[3667]) );
  AND U7039 ( .A(p_input[3666]), .B(p_input[13666]), .Z(o[3666]) );
  AND U7040 ( .A(p_input[3665]), .B(p_input[13665]), .Z(o[3665]) );
  AND U7041 ( .A(p_input[3664]), .B(p_input[13664]), .Z(o[3664]) );
  AND U7042 ( .A(p_input[3663]), .B(p_input[13663]), .Z(o[3663]) );
  AND U7043 ( .A(p_input[3662]), .B(p_input[13662]), .Z(o[3662]) );
  AND U7044 ( .A(p_input[3661]), .B(p_input[13661]), .Z(o[3661]) );
  AND U7045 ( .A(p_input[3660]), .B(p_input[13660]), .Z(o[3660]) );
  AND U7046 ( .A(p_input[365]), .B(p_input[10365]), .Z(o[365]) );
  AND U7047 ( .A(p_input[3659]), .B(p_input[13659]), .Z(o[3659]) );
  AND U7048 ( .A(p_input[3658]), .B(p_input[13658]), .Z(o[3658]) );
  AND U7049 ( .A(p_input[3657]), .B(p_input[13657]), .Z(o[3657]) );
  AND U7050 ( .A(p_input[3656]), .B(p_input[13656]), .Z(o[3656]) );
  AND U7051 ( .A(p_input[3655]), .B(p_input[13655]), .Z(o[3655]) );
  AND U7052 ( .A(p_input[3654]), .B(p_input[13654]), .Z(o[3654]) );
  AND U7053 ( .A(p_input[3653]), .B(p_input[13653]), .Z(o[3653]) );
  AND U7054 ( .A(p_input[3652]), .B(p_input[13652]), .Z(o[3652]) );
  AND U7055 ( .A(p_input[3651]), .B(p_input[13651]), .Z(o[3651]) );
  AND U7056 ( .A(p_input[3650]), .B(p_input[13650]), .Z(o[3650]) );
  AND U7057 ( .A(p_input[364]), .B(p_input[10364]), .Z(o[364]) );
  AND U7058 ( .A(p_input[3649]), .B(p_input[13649]), .Z(o[3649]) );
  AND U7059 ( .A(p_input[3648]), .B(p_input[13648]), .Z(o[3648]) );
  AND U7060 ( .A(p_input[3647]), .B(p_input[13647]), .Z(o[3647]) );
  AND U7061 ( .A(p_input[3646]), .B(p_input[13646]), .Z(o[3646]) );
  AND U7062 ( .A(p_input[3645]), .B(p_input[13645]), .Z(o[3645]) );
  AND U7063 ( .A(p_input[3644]), .B(p_input[13644]), .Z(o[3644]) );
  AND U7064 ( .A(p_input[3643]), .B(p_input[13643]), .Z(o[3643]) );
  AND U7065 ( .A(p_input[3642]), .B(p_input[13642]), .Z(o[3642]) );
  AND U7066 ( .A(p_input[3641]), .B(p_input[13641]), .Z(o[3641]) );
  AND U7067 ( .A(p_input[3640]), .B(p_input[13640]), .Z(o[3640]) );
  AND U7068 ( .A(p_input[363]), .B(p_input[10363]), .Z(o[363]) );
  AND U7069 ( .A(p_input[3639]), .B(p_input[13639]), .Z(o[3639]) );
  AND U7070 ( .A(p_input[3638]), .B(p_input[13638]), .Z(o[3638]) );
  AND U7071 ( .A(p_input[3637]), .B(p_input[13637]), .Z(o[3637]) );
  AND U7072 ( .A(p_input[3636]), .B(p_input[13636]), .Z(o[3636]) );
  AND U7073 ( .A(p_input[3635]), .B(p_input[13635]), .Z(o[3635]) );
  AND U7074 ( .A(p_input[3634]), .B(p_input[13634]), .Z(o[3634]) );
  AND U7075 ( .A(p_input[3633]), .B(p_input[13633]), .Z(o[3633]) );
  AND U7076 ( .A(p_input[3632]), .B(p_input[13632]), .Z(o[3632]) );
  AND U7077 ( .A(p_input[3631]), .B(p_input[13631]), .Z(o[3631]) );
  AND U7078 ( .A(p_input[3630]), .B(p_input[13630]), .Z(o[3630]) );
  AND U7079 ( .A(p_input[362]), .B(p_input[10362]), .Z(o[362]) );
  AND U7080 ( .A(p_input[3629]), .B(p_input[13629]), .Z(o[3629]) );
  AND U7081 ( .A(p_input[3628]), .B(p_input[13628]), .Z(o[3628]) );
  AND U7082 ( .A(p_input[3627]), .B(p_input[13627]), .Z(o[3627]) );
  AND U7083 ( .A(p_input[3626]), .B(p_input[13626]), .Z(o[3626]) );
  AND U7084 ( .A(p_input[3625]), .B(p_input[13625]), .Z(o[3625]) );
  AND U7085 ( .A(p_input[3624]), .B(p_input[13624]), .Z(o[3624]) );
  AND U7086 ( .A(p_input[3623]), .B(p_input[13623]), .Z(o[3623]) );
  AND U7087 ( .A(p_input[3622]), .B(p_input[13622]), .Z(o[3622]) );
  AND U7088 ( .A(p_input[3621]), .B(p_input[13621]), .Z(o[3621]) );
  AND U7089 ( .A(p_input[3620]), .B(p_input[13620]), .Z(o[3620]) );
  AND U7090 ( .A(p_input[361]), .B(p_input[10361]), .Z(o[361]) );
  AND U7091 ( .A(p_input[3619]), .B(p_input[13619]), .Z(o[3619]) );
  AND U7092 ( .A(p_input[3618]), .B(p_input[13618]), .Z(o[3618]) );
  AND U7093 ( .A(p_input[3617]), .B(p_input[13617]), .Z(o[3617]) );
  AND U7094 ( .A(p_input[3616]), .B(p_input[13616]), .Z(o[3616]) );
  AND U7095 ( .A(p_input[3615]), .B(p_input[13615]), .Z(o[3615]) );
  AND U7096 ( .A(p_input[3614]), .B(p_input[13614]), .Z(o[3614]) );
  AND U7097 ( .A(p_input[3613]), .B(p_input[13613]), .Z(o[3613]) );
  AND U7098 ( .A(p_input[3612]), .B(p_input[13612]), .Z(o[3612]) );
  AND U7099 ( .A(p_input[3611]), .B(p_input[13611]), .Z(o[3611]) );
  AND U7100 ( .A(p_input[3610]), .B(p_input[13610]), .Z(o[3610]) );
  AND U7101 ( .A(p_input[360]), .B(p_input[10360]), .Z(o[360]) );
  AND U7102 ( .A(p_input[3609]), .B(p_input[13609]), .Z(o[3609]) );
  AND U7103 ( .A(p_input[3608]), .B(p_input[13608]), .Z(o[3608]) );
  AND U7104 ( .A(p_input[3607]), .B(p_input[13607]), .Z(o[3607]) );
  AND U7105 ( .A(p_input[3606]), .B(p_input[13606]), .Z(o[3606]) );
  AND U7106 ( .A(p_input[3605]), .B(p_input[13605]), .Z(o[3605]) );
  AND U7107 ( .A(p_input[3604]), .B(p_input[13604]), .Z(o[3604]) );
  AND U7108 ( .A(p_input[3603]), .B(p_input[13603]), .Z(o[3603]) );
  AND U7109 ( .A(p_input[3602]), .B(p_input[13602]), .Z(o[3602]) );
  AND U7110 ( .A(p_input[3601]), .B(p_input[13601]), .Z(o[3601]) );
  AND U7111 ( .A(p_input[3600]), .B(p_input[13600]), .Z(o[3600]) );
  AND U7112 ( .A(p_input[35]), .B(p_input[10035]), .Z(o[35]) );
  AND U7113 ( .A(p_input[359]), .B(p_input[10359]), .Z(o[359]) );
  AND U7114 ( .A(p_input[3599]), .B(p_input[13599]), .Z(o[3599]) );
  AND U7115 ( .A(p_input[3598]), .B(p_input[13598]), .Z(o[3598]) );
  AND U7116 ( .A(p_input[3597]), .B(p_input[13597]), .Z(o[3597]) );
  AND U7117 ( .A(p_input[3596]), .B(p_input[13596]), .Z(o[3596]) );
  AND U7118 ( .A(p_input[3595]), .B(p_input[13595]), .Z(o[3595]) );
  AND U7119 ( .A(p_input[3594]), .B(p_input[13594]), .Z(o[3594]) );
  AND U7120 ( .A(p_input[3593]), .B(p_input[13593]), .Z(o[3593]) );
  AND U7121 ( .A(p_input[3592]), .B(p_input[13592]), .Z(o[3592]) );
  AND U7122 ( .A(p_input[3591]), .B(p_input[13591]), .Z(o[3591]) );
  AND U7123 ( .A(p_input[3590]), .B(p_input[13590]), .Z(o[3590]) );
  AND U7124 ( .A(p_input[358]), .B(p_input[10358]), .Z(o[358]) );
  AND U7125 ( .A(p_input[3589]), .B(p_input[13589]), .Z(o[3589]) );
  AND U7126 ( .A(p_input[3588]), .B(p_input[13588]), .Z(o[3588]) );
  AND U7127 ( .A(p_input[3587]), .B(p_input[13587]), .Z(o[3587]) );
  AND U7128 ( .A(p_input[3586]), .B(p_input[13586]), .Z(o[3586]) );
  AND U7129 ( .A(p_input[3585]), .B(p_input[13585]), .Z(o[3585]) );
  AND U7130 ( .A(p_input[3584]), .B(p_input[13584]), .Z(o[3584]) );
  AND U7131 ( .A(p_input[3583]), .B(p_input[13583]), .Z(o[3583]) );
  AND U7132 ( .A(p_input[3582]), .B(p_input[13582]), .Z(o[3582]) );
  AND U7133 ( .A(p_input[3581]), .B(p_input[13581]), .Z(o[3581]) );
  AND U7134 ( .A(p_input[3580]), .B(p_input[13580]), .Z(o[3580]) );
  AND U7135 ( .A(p_input[357]), .B(p_input[10357]), .Z(o[357]) );
  AND U7136 ( .A(p_input[3579]), .B(p_input[13579]), .Z(o[3579]) );
  AND U7137 ( .A(p_input[3578]), .B(p_input[13578]), .Z(o[3578]) );
  AND U7138 ( .A(p_input[3577]), .B(p_input[13577]), .Z(o[3577]) );
  AND U7139 ( .A(p_input[3576]), .B(p_input[13576]), .Z(o[3576]) );
  AND U7140 ( .A(p_input[3575]), .B(p_input[13575]), .Z(o[3575]) );
  AND U7141 ( .A(p_input[3574]), .B(p_input[13574]), .Z(o[3574]) );
  AND U7142 ( .A(p_input[3573]), .B(p_input[13573]), .Z(o[3573]) );
  AND U7143 ( .A(p_input[3572]), .B(p_input[13572]), .Z(o[3572]) );
  AND U7144 ( .A(p_input[3571]), .B(p_input[13571]), .Z(o[3571]) );
  AND U7145 ( .A(p_input[3570]), .B(p_input[13570]), .Z(o[3570]) );
  AND U7146 ( .A(p_input[356]), .B(p_input[10356]), .Z(o[356]) );
  AND U7147 ( .A(p_input[3569]), .B(p_input[13569]), .Z(o[3569]) );
  AND U7148 ( .A(p_input[3568]), .B(p_input[13568]), .Z(o[3568]) );
  AND U7149 ( .A(p_input[3567]), .B(p_input[13567]), .Z(o[3567]) );
  AND U7150 ( .A(p_input[3566]), .B(p_input[13566]), .Z(o[3566]) );
  AND U7151 ( .A(p_input[3565]), .B(p_input[13565]), .Z(o[3565]) );
  AND U7152 ( .A(p_input[3564]), .B(p_input[13564]), .Z(o[3564]) );
  AND U7153 ( .A(p_input[3563]), .B(p_input[13563]), .Z(o[3563]) );
  AND U7154 ( .A(p_input[3562]), .B(p_input[13562]), .Z(o[3562]) );
  AND U7155 ( .A(p_input[3561]), .B(p_input[13561]), .Z(o[3561]) );
  AND U7156 ( .A(p_input[3560]), .B(p_input[13560]), .Z(o[3560]) );
  AND U7157 ( .A(p_input[355]), .B(p_input[10355]), .Z(o[355]) );
  AND U7158 ( .A(p_input[3559]), .B(p_input[13559]), .Z(o[3559]) );
  AND U7159 ( .A(p_input[3558]), .B(p_input[13558]), .Z(o[3558]) );
  AND U7160 ( .A(p_input[3557]), .B(p_input[13557]), .Z(o[3557]) );
  AND U7161 ( .A(p_input[3556]), .B(p_input[13556]), .Z(o[3556]) );
  AND U7162 ( .A(p_input[3555]), .B(p_input[13555]), .Z(o[3555]) );
  AND U7163 ( .A(p_input[3554]), .B(p_input[13554]), .Z(o[3554]) );
  AND U7164 ( .A(p_input[3553]), .B(p_input[13553]), .Z(o[3553]) );
  AND U7165 ( .A(p_input[3552]), .B(p_input[13552]), .Z(o[3552]) );
  AND U7166 ( .A(p_input[3551]), .B(p_input[13551]), .Z(o[3551]) );
  AND U7167 ( .A(p_input[3550]), .B(p_input[13550]), .Z(o[3550]) );
  AND U7168 ( .A(p_input[354]), .B(p_input[10354]), .Z(o[354]) );
  AND U7169 ( .A(p_input[3549]), .B(p_input[13549]), .Z(o[3549]) );
  AND U7170 ( .A(p_input[3548]), .B(p_input[13548]), .Z(o[3548]) );
  AND U7171 ( .A(p_input[3547]), .B(p_input[13547]), .Z(o[3547]) );
  AND U7172 ( .A(p_input[3546]), .B(p_input[13546]), .Z(o[3546]) );
  AND U7173 ( .A(p_input[3545]), .B(p_input[13545]), .Z(o[3545]) );
  AND U7174 ( .A(p_input[3544]), .B(p_input[13544]), .Z(o[3544]) );
  AND U7175 ( .A(p_input[3543]), .B(p_input[13543]), .Z(o[3543]) );
  AND U7176 ( .A(p_input[3542]), .B(p_input[13542]), .Z(o[3542]) );
  AND U7177 ( .A(p_input[3541]), .B(p_input[13541]), .Z(o[3541]) );
  AND U7178 ( .A(p_input[3540]), .B(p_input[13540]), .Z(o[3540]) );
  AND U7179 ( .A(p_input[353]), .B(p_input[10353]), .Z(o[353]) );
  AND U7180 ( .A(p_input[3539]), .B(p_input[13539]), .Z(o[3539]) );
  AND U7181 ( .A(p_input[3538]), .B(p_input[13538]), .Z(o[3538]) );
  AND U7182 ( .A(p_input[3537]), .B(p_input[13537]), .Z(o[3537]) );
  AND U7183 ( .A(p_input[3536]), .B(p_input[13536]), .Z(o[3536]) );
  AND U7184 ( .A(p_input[3535]), .B(p_input[13535]), .Z(o[3535]) );
  AND U7185 ( .A(p_input[3534]), .B(p_input[13534]), .Z(o[3534]) );
  AND U7186 ( .A(p_input[3533]), .B(p_input[13533]), .Z(o[3533]) );
  AND U7187 ( .A(p_input[3532]), .B(p_input[13532]), .Z(o[3532]) );
  AND U7188 ( .A(p_input[3531]), .B(p_input[13531]), .Z(o[3531]) );
  AND U7189 ( .A(p_input[3530]), .B(p_input[13530]), .Z(o[3530]) );
  AND U7190 ( .A(p_input[352]), .B(p_input[10352]), .Z(o[352]) );
  AND U7191 ( .A(p_input[3529]), .B(p_input[13529]), .Z(o[3529]) );
  AND U7192 ( .A(p_input[3528]), .B(p_input[13528]), .Z(o[3528]) );
  AND U7193 ( .A(p_input[3527]), .B(p_input[13527]), .Z(o[3527]) );
  AND U7194 ( .A(p_input[3526]), .B(p_input[13526]), .Z(o[3526]) );
  AND U7195 ( .A(p_input[3525]), .B(p_input[13525]), .Z(o[3525]) );
  AND U7196 ( .A(p_input[3524]), .B(p_input[13524]), .Z(o[3524]) );
  AND U7197 ( .A(p_input[3523]), .B(p_input[13523]), .Z(o[3523]) );
  AND U7198 ( .A(p_input[3522]), .B(p_input[13522]), .Z(o[3522]) );
  AND U7199 ( .A(p_input[3521]), .B(p_input[13521]), .Z(o[3521]) );
  AND U7200 ( .A(p_input[3520]), .B(p_input[13520]), .Z(o[3520]) );
  AND U7201 ( .A(p_input[351]), .B(p_input[10351]), .Z(o[351]) );
  AND U7202 ( .A(p_input[3519]), .B(p_input[13519]), .Z(o[3519]) );
  AND U7203 ( .A(p_input[3518]), .B(p_input[13518]), .Z(o[3518]) );
  AND U7204 ( .A(p_input[3517]), .B(p_input[13517]), .Z(o[3517]) );
  AND U7205 ( .A(p_input[3516]), .B(p_input[13516]), .Z(o[3516]) );
  AND U7206 ( .A(p_input[3515]), .B(p_input[13515]), .Z(o[3515]) );
  AND U7207 ( .A(p_input[3514]), .B(p_input[13514]), .Z(o[3514]) );
  AND U7208 ( .A(p_input[3513]), .B(p_input[13513]), .Z(o[3513]) );
  AND U7209 ( .A(p_input[3512]), .B(p_input[13512]), .Z(o[3512]) );
  AND U7210 ( .A(p_input[3511]), .B(p_input[13511]), .Z(o[3511]) );
  AND U7211 ( .A(p_input[3510]), .B(p_input[13510]), .Z(o[3510]) );
  AND U7212 ( .A(p_input[350]), .B(p_input[10350]), .Z(o[350]) );
  AND U7213 ( .A(p_input[3509]), .B(p_input[13509]), .Z(o[3509]) );
  AND U7214 ( .A(p_input[3508]), .B(p_input[13508]), .Z(o[3508]) );
  AND U7215 ( .A(p_input[3507]), .B(p_input[13507]), .Z(o[3507]) );
  AND U7216 ( .A(p_input[3506]), .B(p_input[13506]), .Z(o[3506]) );
  AND U7217 ( .A(p_input[3505]), .B(p_input[13505]), .Z(o[3505]) );
  AND U7218 ( .A(p_input[3504]), .B(p_input[13504]), .Z(o[3504]) );
  AND U7219 ( .A(p_input[3503]), .B(p_input[13503]), .Z(o[3503]) );
  AND U7220 ( .A(p_input[3502]), .B(p_input[13502]), .Z(o[3502]) );
  AND U7221 ( .A(p_input[3501]), .B(p_input[13501]), .Z(o[3501]) );
  AND U7222 ( .A(p_input[3500]), .B(p_input[13500]), .Z(o[3500]) );
  AND U7223 ( .A(p_input[34]), .B(p_input[10034]), .Z(o[34]) );
  AND U7224 ( .A(p_input[349]), .B(p_input[10349]), .Z(o[349]) );
  AND U7225 ( .A(p_input[3499]), .B(p_input[13499]), .Z(o[3499]) );
  AND U7226 ( .A(p_input[3498]), .B(p_input[13498]), .Z(o[3498]) );
  AND U7227 ( .A(p_input[3497]), .B(p_input[13497]), .Z(o[3497]) );
  AND U7228 ( .A(p_input[3496]), .B(p_input[13496]), .Z(o[3496]) );
  AND U7229 ( .A(p_input[3495]), .B(p_input[13495]), .Z(o[3495]) );
  AND U7230 ( .A(p_input[3494]), .B(p_input[13494]), .Z(o[3494]) );
  AND U7231 ( .A(p_input[3493]), .B(p_input[13493]), .Z(o[3493]) );
  AND U7232 ( .A(p_input[3492]), .B(p_input[13492]), .Z(o[3492]) );
  AND U7233 ( .A(p_input[3491]), .B(p_input[13491]), .Z(o[3491]) );
  AND U7234 ( .A(p_input[3490]), .B(p_input[13490]), .Z(o[3490]) );
  AND U7235 ( .A(p_input[348]), .B(p_input[10348]), .Z(o[348]) );
  AND U7236 ( .A(p_input[3489]), .B(p_input[13489]), .Z(o[3489]) );
  AND U7237 ( .A(p_input[3488]), .B(p_input[13488]), .Z(o[3488]) );
  AND U7238 ( .A(p_input[3487]), .B(p_input[13487]), .Z(o[3487]) );
  AND U7239 ( .A(p_input[3486]), .B(p_input[13486]), .Z(o[3486]) );
  AND U7240 ( .A(p_input[3485]), .B(p_input[13485]), .Z(o[3485]) );
  AND U7241 ( .A(p_input[3484]), .B(p_input[13484]), .Z(o[3484]) );
  AND U7242 ( .A(p_input[3483]), .B(p_input[13483]), .Z(o[3483]) );
  AND U7243 ( .A(p_input[3482]), .B(p_input[13482]), .Z(o[3482]) );
  AND U7244 ( .A(p_input[3481]), .B(p_input[13481]), .Z(o[3481]) );
  AND U7245 ( .A(p_input[3480]), .B(p_input[13480]), .Z(o[3480]) );
  AND U7246 ( .A(p_input[347]), .B(p_input[10347]), .Z(o[347]) );
  AND U7247 ( .A(p_input[3479]), .B(p_input[13479]), .Z(o[3479]) );
  AND U7248 ( .A(p_input[3478]), .B(p_input[13478]), .Z(o[3478]) );
  AND U7249 ( .A(p_input[3477]), .B(p_input[13477]), .Z(o[3477]) );
  AND U7250 ( .A(p_input[3476]), .B(p_input[13476]), .Z(o[3476]) );
  AND U7251 ( .A(p_input[3475]), .B(p_input[13475]), .Z(o[3475]) );
  AND U7252 ( .A(p_input[3474]), .B(p_input[13474]), .Z(o[3474]) );
  AND U7253 ( .A(p_input[3473]), .B(p_input[13473]), .Z(o[3473]) );
  AND U7254 ( .A(p_input[3472]), .B(p_input[13472]), .Z(o[3472]) );
  AND U7255 ( .A(p_input[3471]), .B(p_input[13471]), .Z(o[3471]) );
  AND U7256 ( .A(p_input[3470]), .B(p_input[13470]), .Z(o[3470]) );
  AND U7257 ( .A(p_input[346]), .B(p_input[10346]), .Z(o[346]) );
  AND U7258 ( .A(p_input[3469]), .B(p_input[13469]), .Z(o[3469]) );
  AND U7259 ( .A(p_input[3468]), .B(p_input[13468]), .Z(o[3468]) );
  AND U7260 ( .A(p_input[3467]), .B(p_input[13467]), .Z(o[3467]) );
  AND U7261 ( .A(p_input[3466]), .B(p_input[13466]), .Z(o[3466]) );
  AND U7262 ( .A(p_input[3465]), .B(p_input[13465]), .Z(o[3465]) );
  AND U7263 ( .A(p_input[3464]), .B(p_input[13464]), .Z(o[3464]) );
  AND U7264 ( .A(p_input[3463]), .B(p_input[13463]), .Z(o[3463]) );
  AND U7265 ( .A(p_input[3462]), .B(p_input[13462]), .Z(o[3462]) );
  AND U7266 ( .A(p_input[3461]), .B(p_input[13461]), .Z(o[3461]) );
  AND U7267 ( .A(p_input[3460]), .B(p_input[13460]), .Z(o[3460]) );
  AND U7268 ( .A(p_input[345]), .B(p_input[10345]), .Z(o[345]) );
  AND U7269 ( .A(p_input[3459]), .B(p_input[13459]), .Z(o[3459]) );
  AND U7270 ( .A(p_input[3458]), .B(p_input[13458]), .Z(o[3458]) );
  AND U7271 ( .A(p_input[3457]), .B(p_input[13457]), .Z(o[3457]) );
  AND U7272 ( .A(p_input[3456]), .B(p_input[13456]), .Z(o[3456]) );
  AND U7273 ( .A(p_input[3455]), .B(p_input[13455]), .Z(o[3455]) );
  AND U7274 ( .A(p_input[3454]), .B(p_input[13454]), .Z(o[3454]) );
  AND U7275 ( .A(p_input[3453]), .B(p_input[13453]), .Z(o[3453]) );
  AND U7276 ( .A(p_input[3452]), .B(p_input[13452]), .Z(o[3452]) );
  AND U7277 ( .A(p_input[3451]), .B(p_input[13451]), .Z(o[3451]) );
  AND U7278 ( .A(p_input[3450]), .B(p_input[13450]), .Z(o[3450]) );
  AND U7279 ( .A(p_input[344]), .B(p_input[10344]), .Z(o[344]) );
  AND U7280 ( .A(p_input[3449]), .B(p_input[13449]), .Z(o[3449]) );
  AND U7281 ( .A(p_input[3448]), .B(p_input[13448]), .Z(o[3448]) );
  AND U7282 ( .A(p_input[3447]), .B(p_input[13447]), .Z(o[3447]) );
  AND U7283 ( .A(p_input[3446]), .B(p_input[13446]), .Z(o[3446]) );
  AND U7284 ( .A(p_input[3445]), .B(p_input[13445]), .Z(o[3445]) );
  AND U7285 ( .A(p_input[3444]), .B(p_input[13444]), .Z(o[3444]) );
  AND U7286 ( .A(p_input[3443]), .B(p_input[13443]), .Z(o[3443]) );
  AND U7287 ( .A(p_input[3442]), .B(p_input[13442]), .Z(o[3442]) );
  AND U7288 ( .A(p_input[3441]), .B(p_input[13441]), .Z(o[3441]) );
  AND U7289 ( .A(p_input[3440]), .B(p_input[13440]), .Z(o[3440]) );
  AND U7290 ( .A(p_input[343]), .B(p_input[10343]), .Z(o[343]) );
  AND U7291 ( .A(p_input[3439]), .B(p_input[13439]), .Z(o[3439]) );
  AND U7292 ( .A(p_input[3438]), .B(p_input[13438]), .Z(o[3438]) );
  AND U7293 ( .A(p_input[3437]), .B(p_input[13437]), .Z(o[3437]) );
  AND U7294 ( .A(p_input[3436]), .B(p_input[13436]), .Z(o[3436]) );
  AND U7295 ( .A(p_input[3435]), .B(p_input[13435]), .Z(o[3435]) );
  AND U7296 ( .A(p_input[3434]), .B(p_input[13434]), .Z(o[3434]) );
  AND U7297 ( .A(p_input[3433]), .B(p_input[13433]), .Z(o[3433]) );
  AND U7298 ( .A(p_input[3432]), .B(p_input[13432]), .Z(o[3432]) );
  AND U7299 ( .A(p_input[3431]), .B(p_input[13431]), .Z(o[3431]) );
  AND U7300 ( .A(p_input[3430]), .B(p_input[13430]), .Z(o[3430]) );
  AND U7301 ( .A(p_input[342]), .B(p_input[10342]), .Z(o[342]) );
  AND U7302 ( .A(p_input[3429]), .B(p_input[13429]), .Z(o[3429]) );
  AND U7303 ( .A(p_input[3428]), .B(p_input[13428]), .Z(o[3428]) );
  AND U7304 ( .A(p_input[3427]), .B(p_input[13427]), .Z(o[3427]) );
  AND U7305 ( .A(p_input[3426]), .B(p_input[13426]), .Z(o[3426]) );
  AND U7306 ( .A(p_input[3425]), .B(p_input[13425]), .Z(o[3425]) );
  AND U7307 ( .A(p_input[3424]), .B(p_input[13424]), .Z(o[3424]) );
  AND U7308 ( .A(p_input[3423]), .B(p_input[13423]), .Z(o[3423]) );
  AND U7309 ( .A(p_input[3422]), .B(p_input[13422]), .Z(o[3422]) );
  AND U7310 ( .A(p_input[3421]), .B(p_input[13421]), .Z(o[3421]) );
  AND U7311 ( .A(p_input[3420]), .B(p_input[13420]), .Z(o[3420]) );
  AND U7312 ( .A(p_input[341]), .B(p_input[10341]), .Z(o[341]) );
  AND U7313 ( .A(p_input[3419]), .B(p_input[13419]), .Z(o[3419]) );
  AND U7314 ( .A(p_input[3418]), .B(p_input[13418]), .Z(o[3418]) );
  AND U7315 ( .A(p_input[3417]), .B(p_input[13417]), .Z(o[3417]) );
  AND U7316 ( .A(p_input[3416]), .B(p_input[13416]), .Z(o[3416]) );
  AND U7317 ( .A(p_input[3415]), .B(p_input[13415]), .Z(o[3415]) );
  AND U7318 ( .A(p_input[3414]), .B(p_input[13414]), .Z(o[3414]) );
  AND U7319 ( .A(p_input[3413]), .B(p_input[13413]), .Z(o[3413]) );
  AND U7320 ( .A(p_input[3412]), .B(p_input[13412]), .Z(o[3412]) );
  AND U7321 ( .A(p_input[3411]), .B(p_input[13411]), .Z(o[3411]) );
  AND U7322 ( .A(p_input[3410]), .B(p_input[13410]), .Z(o[3410]) );
  AND U7323 ( .A(p_input[340]), .B(p_input[10340]), .Z(o[340]) );
  AND U7324 ( .A(p_input[3409]), .B(p_input[13409]), .Z(o[3409]) );
  AND U7325 ( .A(p_input[3408]), .B(p_input[13408]), .Z(o[3408]) );
  AND U7326 ( .A(p_input[3407]), .B(p_input[13407]), .Z(o[3407]) );
  AND U7327 ( .A(p_input[3406]), .B(p_input[13406]), .Z(o[3406]) );
  AND U7328 ( .A(p_input[3405]), .B(p_input[13405]), .Z(o[3405]) );
  AND U7329 ( .A(p_input[3404]), .B(p_input[13404]), .Z(o[3404]) );
  AND U7330 ( .A(p_input[3403]), .B(p_input[13403]), .Z(o[3403]) );
  AND U7331 ( .A(p_input[3402]), .B(p_input[13402]), .Z(o[3402]) );
  AND U7332 ( .A(p_input[3401]), .B(p_input[13401]), .Z(o[3401]) );
  AND U7333 ( .A(p_input[3400]), .B(p_input[13400]), .Z(o[3400]) );
  AND U7334 ( .A(p_input[33]), .B(p_input[10033]), .Z(o[33]) );
  AND U7335 ( .A(p_input[339]), .B(p_input[10339]), .Z(o[339]) );
  AND U7336 ( .A(p_input[3399]), .B(p_input[13399]), .Z(o[3399]) );
  AND U7337 ( .A(p_input[3398]), .B(p_input[13398]), .Z(o[3398]) );
  AND U7338 ( .A(p_input[3397]), .B(p_input[13397]), .Z(o[3397]) );
  AND U7339 ( .A(p_input[3396]), .B(p_input[13396]), .Z(o[3396]) );
  AND U7340 ( .A(p_input[3395]), .B(p_input[13395]), .Z(o[3395]) );
  AND U7341 ( .A(p_input[3394]), .B(p_input[13394]), .Z(o[3394]) );
  AND U7342 ( .A(p_input[3393]), .B(p_input[13393]), .Z(o[3393]) );
  AND U7343 ( .A(p_input[3392]), .B(p_input[13392]), .Z(o[3392]) );
  AND U7344 ( .A(p_input[3391]), .B(p_input[13391]), .Z(o[3391]) );
  AND U7345 ( .A(p_input[3390]), .B(p_input[13390]), .Z(o[3390]) );
  AND U7346 ( .A(p_input[338]), .B(p_input[10338]), .Z(o[338]) );
  AND U7347 ( .A(p_input[3389]), .B(p_input[13389]), .Z(o[3389]) );
  AND U7348 ( .A(p_input[3388]), .B(p_input[13388]), .Z(o[3388]) );
  AND U7349 ( .A(p_input[3387]), .B(p_input[13387]), .Z(o[3387]) );
  AND U7350 ( .A(p_input[3386]), .B(p_input[13386]), .Z(o[3386]) );
  AND U7351 ( .A(p_input[3385]), .B(p_input[13385]), .Z(o[3385]) );
  AND U7352 ( .A(p_input[3384]), .B(p_input[13384]), .Z(o[3384]) );
  AND U7353 ( .A(p_input[3383]), .B(p_input[13383]), .Z(o[3383]) );
  AND U7354 ( .A(p_input[3382]), .B(p_input[13382]), .Z(o[3382]) );
  AND U7355 ( .A(p_input[3381]), .B(p_input[13381]), .Z(o[3381]) );
  AND U7356 ( .A(p_input[3380]), .B(p_input[13380]), .Z(o[3380]) );
  AND U7357 ( .A(p_input[337]), .B(p_input[10337]), .Z(o[337]) );
  AND U7358 ( .A(p_input[3379]), .B(p_input[13379]), .Z(o[3379]) );
  AND U7359 ( .A(p_input[3378]), .B(p_input[13378]), .Z(o[3378]) );
  AND U7360 ( .A(p_input[3377]), .B(p_input[13377]), .Z(o[3377]) );
  AND U7361 ( .A(p_input[3376]), .B(p_input[13376]), .Z(o[3376]) );
  AND U7362 ( .A(p_input[3375]), .B(p_input[13375]), .Z(o[3375]) );
  AND U7363 ( .A(p_input[3374]), .B(p_input[13374]), .Z(o[3374]) );
  AND U7364 ( .A(p_input[3373]), .B(p_input[13373]), .Z(o[3373]) );
  AND U7365 ( .A(p_input[3372]), .B(p_input[13372]), .Z(o[3372]) );
  AND U7366 ( .A(p_input[3371]), .B(p_input[13371]), .Z(o[3371]) );
  AND U7367 ( .A(p_input[3370]), .B(p_input[13370]), .Z(o[3370]) );
  AND U7368 ( .A(p_input[336]), .B(p_input[10336]), .Z(o[336]) );
  AND U7369 ( .A(p_input[3369]), .B(p_input[13369]), .Z(o[3369]) );
  AND U7370 ( .A(p_input[3368]), .B(p_input[13368]), .Z(o[3368]) );
  AND U7371 ( .A(p_input[3367]), .B(p_input[13367]), .Z(o[3367]) );
  AND U7372 ( .A(p_input[3366]), .B(p_input[13366]), .Z(o[3366]) );
  AND U7373 ( .A(p_input[3365]), .B(p_input[13365]), .Z(o[3365]) );
  AND U7374 ( .A(p_input[3364]), .B(p_input[13364]), .Z(o[3364]) );
  AND U7375 ( .A(p_input[3363]), .B(p_input[13363]), .Z(o[3363]) );
  AND U7376 ( .A(p_input[3362]), .B(p_input[13362]), .Z(o[3362]) );
  AND U7377 ( .A(p_input[3361]), .B(p_input[13361]), .Z(o[3361]) );
  AND U7378 ( .A(p_input[3360]), .B(p_input[13360]), .Z(o[3360]) );
  AND U7379 ( .A(p_input[335]), .B(p_input[10335]), .Z(o[335]) );
  AND U7380 ( .A(p_input[3359]), .B(p_input[13359]), .Z(o[3359]) );
  AND U7381 ( .A(p_input[3358]), .B(p_input[13358]), .Z(o[3358]) );
  AND U7382 ( .A(p_input[3357]), .B(p_input[13357]), .Z(o[3357]) );
  AND U7383 ( .A(p_input[3356]), .B(p_input[13356]), .Z(o[3356]) );
  AND U7384 ( .A(p_input[3355]), .B(p_input[13355]), .Z(o[3355]) );
  AND U7385 ( .A(p_input[3354]), .B(p_input[13354]), .Z(o[3354]) );
  AND U7386 ( .A(p_input[3353]), .B(p_input[13353]), .Z(o[3353]) );
  AND U7387 ( .A(p_input[3352]), .B(p_input[13352]), .Z(o[3352]) );
  AND U7388 ( .A(p_input[3351]), .B(p_input[13351]), .Z(o[3351]) );
  AND U7389 ( .A(p_input[3350]), .B(p_input[13350]), .Z(o[3350]) );
  AND U7390 ( .A(p_input[334]), .B(p_input[10334]), .Z(o[334]) );
  AND U7391 ( .A(p_input[3349]), .B(p_input[13349]), .Z(o[3349]) );
  AND U7392 ( .A(p_input[3348]), .B(p_input[13348]), .Z(o[3348]) );
  AND U7393 ( .A(p_input[3347]), .B(p_input[13347]), .Z(o[3347]) );
  AND U7394 ( .A(p_input[3346]), .B(p_input[13346]), .Z(o[3346]) );
  AND U7395 ( .A(p_input[3345]), .B(p_input[13345]), .Z(o[3345]) );
  AND U7396 ( .A(p_input[3344]), .B(p_input[13344]), .Z(o[3344]) );
  AND U7397 ( .A(p_input[3343]), .B(p_input[13343]), .Z(o[3343]) );
  AND U7398 ( .A(p_input[3342]), .B(p_input[13342]), .Z(o[3342]) );
  AND U7399 ( .A(p_input[3341]), .B(p_input[13341]), .Z(o[3341]) );
  AND U7400 ( .A(p_input[3340]), .B(p_input[13340]), .Z(o[3340]) );
  AND U7401 ( .A(p_input[333]), .B(p_input[10333]), .Z(o[333]) );
  AND U7402 ( .A(p_input[3339]), .B(p_input[13339]), .Z(o[3339]) );
  AND U7403 ( .A(p_input[3338]), .B(p_input[13338]), .Z(o[3338]) );
  AND U7404 ( .A(p_input[3337]), .B(p_input[13337]), .Z(o[3337]) );
  AND U7405 ( .A(p_input[3336]), .B(p_input[13336]), .Z(o[3336]) );
  AND U7406 ( .A(p_input[3335]), .B(p_input[13335]), .Z(o[3335]) );
  AND U7407 ( .A(p_input[3334]), .B(p_input[13334]), .Z(o[3334]) );
  AND U7408 ( .A(p_input[3333]), .B(p_input[13333]), .Z(o[3333]) );
  AND U7409 ( .A(p_input[3332]), .B(p_input[13332]), .Z(o[3332]) );
  AND U7410 ( .A(p_input[3331]), .B(p_input[13331]), .Z(o[3331]) );
  AND U7411 ( .A(p_input[3330]), .B(p_input[13330]), .Z(o[3330]) );
  AND U7412 ( .A(p_input[332]), .B(p_input[10332]), .Z(o[332]) );
  AND U7413 ( .A(p_input[3329]), .B(p_input[13329]), .Z(o[3329]) );
  AND U7414 ( .A(p_input[3328]), .B(p_input[13328]), .Z(o[3328]) );
  AND U7415 ( .A(p_input[3327]), .B(p_input[13327]), .Z(o[3327]) );
  AND U7416 ( .A(p_input[3326]), .B(p_input[13326]), .Z(o[3326]) );
  AND U7417 ( .A(p_input[3325]), .B(p_input[13325]), .Z(o[3325]) );
  AND U7418 ( .A(p_input[3324]), .B(p_input[13324]), .Z(o[3324]) );
  AND U7419 ( .A(p_input[3323]), .B(p_input[13323]), .Z(o[3323]) );
  AND U7420 ( .A(p_input[3322]), .B(p_input[13322]), .Z(o[3322]) );
  AND U7421 ( .A(p_input[3321]), .B(p_input[13321]), .Z(o[3321]) );
  AND U7422 ( .A(p_input[3320]), .B(p_input[13320]), .Z(o[3320]) );
  AND U7423 ( .A(p_input[331]), .B(p_input[10331]), .Z(o[331]) );
  AND U7424 ( .A(p_input[3319]), .B(p_input[13319]), .Z(o[3319]) );
  AND U7425 ( .A(p_input[3318]), .B(p_input[13318]), .Z(o[3318]) );
  AND U7426 ( .A(p_input[3317]), .B(p_input[13317]), .Z(o[3317]) );
  AND U7427 ( .A(p_input[3316]), .B(p_input[13316]), .Z(o[3316]) );
  AND U7428 ( .A(p_input[3315]), .B(p_input[13315]), .Z(o[3315]) );
  AND U7429 ( .A(p_input[3314]), .B(p_input[13314]), .Z(o[3314]) );
  AND U7430 ( .A(p_input[3313]), .B(p_input[13313]), .Z(o[3313]) );
  AND U7431 ( .A(p_input[3312]), .B(p_input[13312]), .Z(o[3312]) );
  AND U7432 ( .A(p_input[3311]), .B(p_input[13311]), .Z(o[3311]) );
  AND U7433 ( .A(p_input[3310]), .B(p_input[13310]), .Z(o[3310]) );
  AND U7434 ( .A(p_input[330]), .B(p_input[10330]), .Z(o[330]) );
  AND U7435 ( .A(p_input[3309]), .B(p_input[13309]), .Z(o[3309]) );
  AND U7436 ( .A(p_input[3308]), .B(p_input[13308]), .Z(o[3308]) );
  AND U7437 ( .A(p_input[3307]), .B(p_input[13307]), .Z(o[3307]) );
  AND U7438 ( .A(p_input[3306]), .B(p_input[13306]), .Z(o[3306]) );
  AND U7439 ( .A(p_input[3305]), .B(p_input[13305]), .Z(o[3305]) );
  AND U7440 ( .A(p_input[3304]), .B(p_input[13304]), .Z(o[3304]) );
  AND U7441 ( .A(p_input[3303]), .B(p_input[13303]), .Z(o[3303]) );
  AND U7442 ( .A(p_input[3302]), .B(p_input[13302]), .Z(o[3302]) );
  AND U7443 ( .A(p_input[3301]), .B(p_input[13301]), .Z(o[3301]) );
  AND U7444 ( .A(p_input[3300]), .B(p_input[13300]), .Z(o[3300]) );
  AND U7445 ( .A(p_input[32]), .B(p_input[10032]), .Z(o[32]) );
  AND U7446 ( .A(p_input[329]), .B(p_input[10329]), .Z(o[329]) );
  AND U7447 ( .A(p_input[3299]), .B(p_input[13299]), .Z(o[3299]) );
  AND U7448 ( .A(p_input[3298]), .B(p_input[13298]), .Z(o[3298]) );
  AND U7449 ( .A(p_input[3297]), .B(p_input[13297]), .Z(o[3297]) );
  AND U7450 ( .A(p_input[3296]), .B(p_input[13296]), .Z(o[3296]) );
  AND U7451 ( .A(p_input[3295]), .B(p_input[13295]), .Z(o[3295]) );
  AND U7452 ( .A(p_input[3294]), .B(p_input[13294]), .Z(o[3294]) );
  AND U7453 ( .A(p_input[3293]), .B(p_input[13293]), .Z(o[3293]) );
  AND U7454 ( .A(p_input[3292]), .B(p_input[13292]), .Z(o[3292]) );
  AND U7455 ( .A(p_input[3291]), .B(p_input[13291]), .Z(o[3291]) );
  AND U7456 ( .A(p_input[3290]), .B(p_input[13290]), .Z(o[3290]) );
  AND U7457 ( .A(p_input[328]), .B(p_input[10328]), .Z(o[328]) );
  AND U7458 ( .A(p_input[3289]), .B(p_input[13289]), .Z(o[3289]) );
  AND U7459 ( .A(p_input[3288]), .B(p_input[13288]), .Z(o[3288]) );
  AND U7460 ( .A(p_input[3287]), .B(p_input[13287]), .Z(o[3287]) );
  AND U7461 ( .A(p_input[3286]), .B(p_input[13286]), .Z(o[3286]) );
  AND U7462 ( .A(p_input[3285]), .B(p_input[13285]), .Z(o[3285]) );
  AND U7463 ( .A(p_input[3284]), .B(p_input[13284]), .Z(o[3284]) );
  AND U7464 ( .A(p_input[3283]), .B(p_input[13283]), .Z(o[3283]) );
  AND U7465 ( .A(p_input[3282]), .B(p_input[13282]), .Z(o[3282]) );
  AND U7466 ( .A(p_input[3281]), .B(p_input[13281]), .Z(o[3281]) );
  AND U7467 ( .A(p_input[3280]), .B(p_input[13280]), .Z(o[3280]) );
  AND U7468 ( .A(p_input[327]), .B(p_input[10327]), .Z(o[327]) );
  AND U7469 ( .A(p_input[3279]), .B(p_input[13279]), .Z(o[3279]) );
  AND U7470 ( .A(p_input[3278]), .B(p_input[13278]), .Z(o[3278]) );
  AND U7471 ( .A(p_input[3277]), .B(p_input[13277]), .Z(o[3277]) );
  AND U7472 ( .A(p_input[3276]), .B(p_input[13276]), .Z(o[3276]) );
  AND U7473 ( .A(p_input[3275]), .B(p_input[13275]), .Z(o[3275]) );
  AND U7474 ( .A(p_input[3274]), .B(p_input[13274]), .Z(o[3274]) );
  AND U7475 ( .A(p_input[3273]), .B(p_input[13273]), .Z(o[3273]) );
  AND U7476 ( .A(p_input[3272]), .B(p_input[13272]), .Z(o[3272]) );
  AND U7477 ( .A(p_input[3271]), .B(p_input[13271]), .Z(o[3271]) );
  AND U7478 ( .A(p_input[3270]), .B(p_input[13270]), .Z(o[3270]) );
  AND U7479 ( .A(p_input[326]), .B(p_input[10326]), .Z(o[326]) );
  AND U7480 ( .A(p_input[3269]), .B(p_input[13269]), .Z(o[3269]) );
  AND U7481 ( .A(p_input[3268]), .B(p_input[13268]), .Z(o[3268]) );
  AND U7482 ( .A(p_input[3267]), .B(p_input[13267]), .Z(o[3267]) );
  AND U7483 ( .A(p_input[3266]), .B(p_input[13266]), .Z(o[3266]) );
  AND U7484 ( .A(p_input[3265]), .B(p_input[13265]), .Z(o[3265]) );
  AND U7485 ( .A(p_input[3264]), .B(p_input[13264]), .Z(o[3264]) );
  AND U7486 ( .A(p_input[3263]), .B(p_input[13263]), .Z(o[3263]) );
  AND U7487 ( .A(p_input[3262]), .B(p_input[13262]), .Z(o[3262]) );
  AND U7488 ( .A(p_input[3261]), .B(p_input[13261]), .Z(o[3261]) );
  AND U7489 ( .A(p_input[3260]), .B(p_input[13260]), .Z(o[3260]) );
  AND U7490 ( .A(p_input[325]), .B(p_input[10325]), .Z(o[325]) );
  AND U7491 ( .A(p_input[3259]), .B(p_input[13259]), .Z(o[3259]) );
  AND U7492 ( .A(p_input[3258]), .B(p_input[13258]), .Z(o[3258]) );
  AND U7493 ( .A(p_input[3257]), .B(p_input[13257]), .Z(o[3257]) );
  AND U7494 ( .A(p_input[3256]), .B(p_input[13256]), .Z(o[3256]) );
  AND U7495 ( .A(p_input[3255]), .B(p_input[13255]), .Z(o[3255]) );
  AND U7496 ( .A(p_input[3254]), .B(p_input[13254]), .Z(o[3254]) );
  AND U7497 ( .A(p_input[3253]), .B(p_input[13253]), .Z(o[3253]) );
  AND U7498 ( .A(p_input[3252]), .B(p_input[13252]), .Z(o[3252]) );
  AND U7499 ( .A(p_input[3251]), .B(p_input[13251]), .Z(o[3251]) );
  AND U7500 ( .A(p_input[3250]), .B(p_input[13250]), .Z(o[3250]) );
  AND U7501 ( .A(p_input[324]), .B(p_input[10324]), .Z(o[324]) );
  AND U7502 ( .A(p_input[3249]), .B(p_input[13249]), .Z(o[3249]) );
  AND U7503 ( .A(p_input[3248]), .B(p_input[13248]), .Z(o[3248]) );
  AND U7504 ( .A(p_input[3247]), .B(p_input[13247]), .Z(o[3247]) );
  AND U7505 ( .A(p_input[3246]), .B(p_input[13246]), .Z(o[3246]) );
  AND U7506 ( .A(p_input[3245]), .B(p_input[13245]), .Z(o[3245]) );
  AND U7507 ( .A(p_input[3244]), .B(p_input[13244]), .Z(o[3244]) );
  AND U7508 ( .A(p_input[3243]), .B(p_input[13243]), .Z(o[3243]) );
  AND U7509 ( .A(p_input[3242]), .B(p_input[13242]), .Z(o[3242]) );
  AND U7510 ( .A(p_input[3241]), .B(p_input[13241]), .Z(o[3241]) );
  AND U7511 ( .A(p_input[3240]), .B(p_input[13240]), .Z(o[3240]) );
  AND U7512 ( .A(p_input[323]), .B(p_input[10323]), .Z(o[323]) );
  AND U7513 ( .A(p_input[3239]), .B(p_input[13239]), .Z(o[3239]) );
  AND U7514 ( .A(p_input[3238]), .B(p_input[13238]), .Z(o[3238]) );
  AND U7515 ( .A(p_input[3237]), .B(p_input[13237]), .Z(o[3237]) );
  AND U7516 ( .A(p_input[3236]), .B(p_input[13236]), .Z(o[3236]) );
  AND U7517 ( .A(p_input[3235]), .B(p_input[13235]), .Z(o[3235]) );
  AND U7518 ( .A(p_input[3234]), .B(p_input[13234]), .Z(o[3234]) );
  AND U7519 ( .A(p_input[3233]), .B(p_input[13233]), .Z(o[3233]) );
  AND U7520 ( .A(p_input[3232]), .B(p_input[13232]), .Z(o[3232]) );
  AND U7521 ( .A(p_input[3231]), .B(p_input[13231]), .Z(o[3231]) );
  AND U7522 ( .A(p_input[3230]), .B(p_input[13230]), .Z(o[3230]) );
  AND U7523 ( .A(p_input[322]), .B(p_input[10322]), .Z(o[322]) );
  AND U7524 ( .A(p_input[3229]), .B(p_input[13229]), .Z(o[3229]) );
  AND U7525 ( .A(p_input[3228]), .B(p_input[13228]), .Z(o[3228]) );
  AND U7526 ( .A(p_input[3227]), .B(p_input[13227]), .Z(o[3227]) );
  AND U7527 ( .A(p_input[3226]), .B(p_input[13226]), .Z(o[3226]) );
  AND U7528 ( .A(p_input[3225]), .B(p_input[13225]), .Z(o[3225]) );
  AND U7529 ( .A(p_input[3224]), .B(p_input[13224]), .Z(o[3224]) );
  AND U7530 ( .A(p_input[3223]), .B(p_input[13223]), .Z(o[3223]) );
  AND U7531 ( .A(p_input[3222]), .B(p_input[13222]), .Z(o[3222]) );
  AND U7532 ( .A(p_input[3221]), .B(p_input[13221]), .Z(o[3221]) );
  AND U7533 ( .A(p_input[3220]), .B(p_input[13220]), .Z(o[3220]) );
  AND U7534 ( .A(p_input[321]), .B(p_input[10321]), .Z(o[321]) );
  AND U7535 ( .A(p_input[3219]), .B(p_input[13219]), .Z(o[3219]) );
  AND U7536 ( .A(p_input[3218]), .B(p_input[13218]), .Z(o[3218]) );
  AND U7537 ( .A(p_input[3217]), .B(p_input[13217]), .Z(o[3217]) );
  AND U7538 ( .A(p_input[3216]), .B(p_input[13216]), .Z(o[3216]) );
  AND U7539 ( .A(p_input[3215]), .B(p_input[13215]), .Z(o[3215]) );
  AND U7540 ( .A(p_input[3214]), .B(p_input[13214]), .Z(o[3214]) );
  AND U7541 ( .A(p_input[3213]), .B(p_input[13213]), .Z(o[3213]) );
  AND U7542 ( .A(p_input[3212]), .B(p_input[13212]), .Z(o[3212]) );
  AND U7543 ( .A(p_input[3211]), .B(p_input[13211]), .Z(o[3211]) );
  AND U7544 ( .A(p_input[3210]), .B(p_input[13210]), .Z(o[3210]) );
  AND U7545 ( .A(p_input[320]), .B(p_input[10320]), .Z(o[320]) );
  AND U7546 ( .A(p_input[3209]), .B(p_input[13209]), .Z(o[3209]) );
  AND U7547 ( .A(p_input[3208]), .B(p_input[13208]), .Z(o[3208]) );
  AND U7548 ( .A(p_input[3207]), .B(p_input[13207]), .Z(o[3207]) );
  AND U7549 ( .A(p_input[3206]), .B(p_input[13206]), .Z(o[3206]) );
  AND U7550 ( .A(p_input[3205]), .B(p_input[13205]), .Z(o[3205]) );
  AND U7551 ( .A(p_input[3204]), .B(p_input[13204]), .Z(o[3204]) );
  AND U7552 ( .A(p_input[3203]), .B(p_input[13203]), .Z(o[3203]) );
  AND U7553 ( .A(p_input[3202]), .B(p_input[13202]), .Z(o[3202]) );
  AND U7554 ( .A(p_input[3201]), .B(p_input[13201]), .Z(o[3201]) );
  AND U7555 ( .A(p_input[3200]), .B(p_input[13200]), .Z(o[3200]) );
  AND U7556 ( .A(p_input[31]), .B(p_input[10031]), .Z(o[31]) );
  AND U7557 ( .A(p_input[319]), .B(p_input[10319]), .Z(o[319]) );
  AND U7558 ( .A(p_input[3199]), .B(p_input[13199]), .Z(o[3199]) );
  AND U7559 ( .A(p_input[3198]), .B(p_input[13198]), .Z(o[3198]) );
  AND U7560 ( .A(p_input[3197]), .B(p_input[13197]), .Z(o[3197]) );
  AND U7561 ( .A(p_input[3196]), .B(p_input[13196]), .Z(o[3196]) );
  AND U7562 ( .A(p_input[3195]), .B(p_input[13195]), .Z(o[3195]) );
  AND U7563 ( .A(p_input[3194]), .B(p_input[13194]), .Z(o[3194]) );
  AND U7564 ( .A(p_input[3193]), .B(p_input[13193]), .Z(o[3193]) );
  AND U7565 ( .A(p_input[3192]), .B(p_input[13192]), .Z(o[3192]) );
  AND U7566 ( .A(p_input[3191]), .B(p_input[13191]), .Z(o[3191]) );
  AND U7567 ( .A(p_input[3190]), .B(p_input[13190]), .Z(o[3190]) );
  AND U7568 ( .A(p_input[318]), .B(p_input[10318]), .Z(o[318]) );
  AND U7569 ( .A(p_input[3189]), .B(p_input[13189]), .Z(o[3189]) );
  AND U7570 ( .A(p_input[3188]), .B(p_input[13188]), .Z(o[3188]) );
  AND U7571 ( .A(p_input[3187]), .B(p_input[13187]), .Z(o[3187]) );
  AND U7572 ( .A(p_input[3186]), .B(p_input[13186]), .Z(o[3186]) );
  AND U7573 ( .A(p_input[3185]), .B(p_input[13185]), .Z(o[3185]) );
  AND U7574 ( .A(p_input[3184]), .B(p_input[13184]), .Z(o[3184]) );
  AND U7575 ( .A(p_input[3183]), .B(p_input[13183]), .Z(o[3183]) );
  AND U7576 ( .A(p_input[3182]), .B(p_input[13182]), .Z(o[3182]) );
  AND U7577 ( .A(p_input[3181]), .B(p_input[13181]), .Z(o[3181]) );
  AND U7578 ( .A(p_input[3180]), .B(p_input[13180]), .Z(o[3180]) );
  AND U7579 ( .A(p_input[317]), .B(p_input[10317]), .Z(o[317]) );
  AND U7580 ( .A(p_input[3179]), .B(p_input[13179]), .Z(o[3179]) );
  AND U7581 ( .A(p_input[3178]), .B(p_input[13178]), .Z(o[3178]) );
  AND U7582 ( .A(p_input[3177]), .B(p_input[13177]), .Z(o[3177]) );
  AND U7583 ( .A(p_input[3176]), .B(p_input[13176]), .Z(o[3176]) );
  AND U7584 ( .A(p_input[3175]), .B(p_input[13175]), .Z(o[3175]) );
  AND U7585 ( .A(p_input[3174]), .B(p_input[13174]), .Z(o[3174]) );
  AND U7586 ( .A(p_input[3173]), .B(p_input[13173]), .Z(o[3173]) );
  AND U7587 ( .A(p_input[3172]), .B(p_input[13172]), .Z(o[3172]) );
  AND U7588 ( .A(p_input[3171]), .B(p_input[13171]), .Z(o[3171]) );
  AND U7589 ( .A(p_input[3170]), .B(p_input[13170]), .Z(o[3170]) );
  AND U7590 ( .A(p_input[316]), .B(p_input[10316]), .Z(o[316]) );
  AND U7591 ( .A(p_input[3169]), .B(p_input[13169]), .Z(o[3169]) );
  AND U7592 ( .A(p_input[3168]), .B(p_input[13168]), .Z(o[3168]) );
  AND U7593 ( .A(p_input[3167]), .B(p_input[13167]), .Z(o[3167]) );
  AND U7594 ( .A(p_input[3166]), .B(p_input[13166]), .Z(o[3166]) );
  AND U7595 ( .A(p_input[3165]), .B(p_input[13165]), .Z(o[3165]) );
  AND U7596 ( .A(p_input[3164]), .B(p_input[13164]), .Z(o[3164]) );
  AND U7597 ( .A(p_input[3163]), .B(p_input[13163]), .Z(o[3163]) );
  AND U7598 ( .A(p_input[3162]), .B(p_input[13162]), .Z(o[3162]) );
  AND U7599 ( .A(p_input[3161]), .B(p_input[13161]), .Z(o[3161]) );
  AND U7600 ( .A(p_input[3160]), .B(p_input[13160]), .Z(o[3160]) );
  AND U7601 ( .A(p_input[315]), .B(p_input[10315]), .Z(o[315]) );
  AND U7602 ( .A(p_input[3159]), .B(p_input[13159]), .Z(o[3159]) );
  AND U7603 ( .A(p_input[3158]), .B(p_input[13158]), .Z(o[3158]) );
  AND U7604 ( .A(p_input[3157]), .B(p_input[13157]), .Z(o[3157]) );
  AND U7605 ( .A(p_input[3156]), .B(p_input[13156]), .Z(o[3156]) );
  AND U7606 ( .A(p_input[3155]), .B(p_input[13155]), .Z(o[3155]) );
  AND U7607 ( .A(p_input[3154]), .B(p_input[13154]), .Z(o[3154]) );
  AND U7608 ( .A(p_input[3153]), .B(p_input[13153]), .Z(o[3153]) );
  AND U7609 ( .A(p_input[3152]), .B(p_input[13152]), .Z(o[3152]) );
  AND U7610 ( .A(p_input[3151]), .B(p_input[13151]), .Z(o[3151]) );
  AND U7611 ( .A(p_input[3150]), .B(p_input[13150]), .Z(o[3150]) );
  AND U7612 ( .A(p_input[314]), .B(p_input[10314]), .Z(o[314]) );
  AND U7613 ( .A(p_input[3149]), .B(p_input[13149]), .Z(o[3149]) );
  AND U7614 ( .A(p_input[3148]), .B(p_input[13148]), .Z(o[3148]) );
  AND U7615 ( .A(p_input[3147]), .B(p_input[13147]), .Z(o[3147]) );
  AND U7616 ( .A(p_input[3146]), .B(p_input[13146]), .Z(o[3146]) );
  AND U7617 ( .A(p_input[3145]), .B(p_input[13145]), .Z(o[3145]) );
  AND U7618 ( .A(p_input[3144]), .B(p_input[13144]), .Z(o[3144]) );
  AND U7619 ( .A(p_input[3143]), .B(p_input[13143]), .Z(o[3143]) );
  AND U7620 ( .A(p_input[3142]), .B(p_input[13142]), .Z(o[3142]) );
  AND U7621 ( .A(p_input[3141]), .B(p_input[13141]), .Z(o[3141]) );
  AND U7622 ( .A(p_input[3140]), .B(p_input[13140]), .Z(o[3140]) );
  AND U7623 ( .A(p_input[313]), .B(p_input[10313]), .Z(o[313]) );
  AND U7624 ( .A(p_input[3139]), .B(p_input[13139]), .Z(o[3139]) );
  AND U7625 ( .A(p_input[3138]), .B(p_input[13138]), .Z(o[3138]) );
  AND U7626 ( .A(p_input[3137]), .B(p_input[13137]), .Z(o[3137]) );
  AND U7627 ( .A(p_input[3136]), .B(p_input[13136]), .Z(o[3136]) );
  AND U7628 ( .A(p_input[3135]), .B(p_input[13135]), .Z(o[3135]) );
  AND U7629 ( .A(p_input[3134]), .B(p_input[13134]), .Z(o[3134]) );
  AND U7630 ( .A(p_input[3133]), .B(p_input[13133]), .Z(o[3133]) );
  AND U7631 ( .A(p_input[3132]), .B(p_input[13132]), .Z(o[3132]) );
  AND U7632 ( .A(p_input[3131]), .B(p_input[13131]), .Z(o[3131]) );
  AND U7633 ( .A(p_input[3130]), .B(p_input[13130]), .Z(o[3130]) );
  AND U7634 ( .A(p_input[312]), .B(p_input[10312]), .Z(o[312]) );
  AND U7635 ( .A(p_input[3129]), .B(p_input[13129]), .Z(o[3129]) );
  AND U7636 ( .A(p_input[3128]), .B(p_input[13128]), .Z(o[3128]) );
  AND U7637 ( .A(p_input[3127]), .B(p_input[13127]), .Z(o[3127]) );
  AND U7638 ( .A(p_input[3126]), .B(p_input[13126]), .Z(o[3126]) );
  AND U7639 ( .A(p_input[3125]), .B(p_input[13125]), .Z(o[3125]) );
  AND U7640 ( .A(p_input[3124]), .B(p_input[13124]), .Z(o[3124]) );
  AND U7641 ( .A(p_input[3123]), .B(p_input[13123]), .Z(o[3123]) );
  AND U7642 ( .A(p_input[3122]), .B(p_input[13122]), .Z(o[3122]) );
  AND U7643 ( .A(p_input[3121]), .B(p_input[13121]), .Z(o[3121]) );
  AND U7644 ( .A(p_input[3120]), .B(p_input[13120]), .Z(o[3120]) );
  AND U7645 ( .A(p_input[311]), .B(p_input[10311]), .Z(o[311]) );
  AND U7646 ( .A(p_input[3119]), .B(p_input[13119]), .Z(o[3119]) );
  AND U7647 ( .A(p_input[3118]), .B(p_input[13118]), .Z(o[3118]) );
  AND U7648 ( .A(p_input[3117]), .B(p_input[13117]), .Z(o[3117]) );
  AND U7649 ( .A(p_input[3116]), .B(p_input[13116]), .Z(o[3116]) );
  AND U7650 ( .A(p_input[3115]), .B(p_input[13115]), .Z(o[3115]) );
  AND U7651 ( .A(p_input[3114]), .B(p_input[13114]), .Z(o[3114]) );
  AND U7652 ( .A(p_input[3113]), .B(p_input[13113]), .Z(o[3113]) );
  AND U7653 ( .A(p_input[3112]), .B(p_input[13112]), .Z(o[3112]) );
  AND U7654 ( .A(p_input[3111]), .B(p_input[13111]), .Z(o[3111]) );
  AND U7655 ( .A(p_input[3110]), .B(p_input[13110]), .Z(o[3110]) );
  AND U7656 ( .A(p_input[310]), .B(p_input[10310]), .Z(o[310]) );
  AND U7657 ( .A(p_input[3109]), .B(p_input[13109]), .Z(o[3109]) );
  AND U7658 ( .A(p_input[3108]), .B(p_input[13108]), .Z(o[3108]) );
  AND U7659 ( .A(p_input[3107]), .B(p_input[13107]), .Z(o[3107]) );
  AND U7660 ( .A(p_input[3106]), .B(p_input[13106]), .Z(o[3106]) );
  AND U7661 ( .A(p_input[3105]), .B(p_input[13105]), .Z(o[3105]) );
  AND U7662 ( .A(p_input[3104]), .B(p_input[13104]), .Z(o[3104]) );
  AND U7663 ( .A(p_input[3103]), .B(p_input[13103]), .Z(o[3103]) );
  AND U7664 ( .A(p_input[3102]), .B(p_input[13102]), .Z(o[3102]) );
  AND U7665 ( .A(p_input[3101]), .B(p_input[13101]), .Z(o[3101]) );
  AND U7666 ( .A(p_input[3100]), .B(p_input[13100]), .Z(o[3100]) );
  AND U7667 ( .A(p_input[30]), .B(p_input[10030]), .Z(o[30]) );
  AND U7668 ( .A(p_input[309]), .B(p_input[10309]), .Z(o[309]) );
  AND U7669 ( .A(p_input[3099]), .B(p_input[13099]), .Z(o[3099]) );
  AND U7670 ( .A(p_input[3098]), .B(p_input[13098]), .Z(o[3098]) );
  AND U7671 ( .A(p_input[3097]), .B(p_input[13097]), .Z(o[3097]) );
  AND U7672 ( .A(p_input[3096]), .B(p_input[13096]), .Z(o[3096]) );
  AND U7673 ( .A(p_input[3095]), .B(p_input[13095]), .Z(o[3095]) );
  AND U7674 ( .A(p_input[3094]), .B(p_input[13094]), .Z(o[3094]) );
  AND U7675 ( .A(p_input[3093]), .B(p_input[13093]), .Z(o[3093]) );
  AND U7676 ( .A(p_input[3092]), .B(p_input[13092]), .Z(o[3092]) );
  AND U7677 ( .A(p_input[3091]), .B(p_input[13091]), .Z(o[3091]) );
  AND U7678 ( .A(p_input[3090]), .B(p_input[13090]), .Z(o[3090]) );
  AND U7679 ( .A(p_input[308]), .B(p_input[10308]), .Z(o[308]) );
  AND U7680 ( .A(p_input[3089]), .B(p_input[13089]), .Z(o[3089]) );
  AND U7681 ( .A(p_input[3088]), .B(p_input[13088]), .Z(o[3088]) );
  AND U7682 ( .A(p_input[3087]), .B(p_input[13087]), .Z(o[3087]) );
  AND U7683 ( .A(p_input[3086]), .B(p_input[13086]), .Z(o[3086]) );
  AND U7684 ( .A(p_input[3085]), .B(p_input[13085]), .Z(o[3085]) );
  AND U7685 ( .A(p_input[3084]), .B(p_input[13084]), .Z(o[3084]) );
  AND U7686 ( .A(p_input[3083]), .B(p_input[13083]), .Z(o[3083]) );
  AND U7687 ( .A(p_input[3082]), .B(p_input[13082]), .Z(o[3082]) );
  AND U7688 ( .A(p_input[3081]), .B(p_input[13081]), .Z(o[3081]) );
  AND U7689 ( .A(p_input[3080]), .B(p_input[13080]), .Z(o[3080]) );
  AND U7690 ( .A(p_input[307]), .B(p_input[10307]), .Z(o[307]) );
  AND U7691 ( .A(p_input[3079]), .B(p_input[13079]), .Z(o[3079]) );
  AND U7692 ( .A(p_input[3078]), .B(p_input[13078]), .Z(o[3078]) );
  AND U7693 ( .A(p_input[3077]), .B(p_input[13077]), .Z(o[3077]) );
  AND U7694 ( .A(p_input[3076]), .B(p_input[13076]), .Z(o[3076]) );
  AND U7695 ( .A(p_input[3075]), .B(p_input[13075]), .Z(o[3075]) );
  AND U7696 ( .A(p_input[3074]), .B(p_input[13074]), .Z(o[3074]) );
  AND U7697 ( .A(p_input[3073]), .B(p_input[13073]), .Z(o[3073]) );
  AND U7698 ( .A(p_input[3072]), .B(p_input[13072]), .Z(o[3072]) );
  AND U7699 ( .A(p_input[3071]), .B(p_input[13071]), .Z(o[3071]) );
  AND U7700 ( .A(p_input[3070]), .B(p_input[13070]), .Z(o[3070]) );
  AND U7701 ( .A(p_input[306]), .B(p_input[10306]), .Z(o[306]) );
  AND U7702 ( .A(p_input[3069]), .B(p_input[13069]), .Z(o[3069]) );
  AND U7703 ( .A(p_input[3068]), .B(p_input[13068]), .Z(o[3068]) );
  AND U7704 ( .A(p_input[3067]), .B(p_input[13067]), .Z(o[3067]) );
  AND U7705 ( .A(p_input[3066]), .B(p_input[13066]), .Z(o[3066]) );
  AND U7706 ( .A(p_input[3065]), .B(p_input[13065]), .Z(o[3065]) );
  AND U7707 ( .A(p_input[3064]), .B(p_input[13064]), .Z(o[3064]) );
  AND U7708 ( .A(p_input[3063]), .B(p_input[13063]), .Z(o[3063]) );
  AND U7709 ( .A(p_input[3062]), .B(p_input[13062]), .Z(o[3062]) );
  AND U7710 ( .A(p_input[3061]), .B(p_input[13061]), .Z(o[3061]) );
  AND U7711 ( .A(p_input[3060]), .B(p_input[13060]), .Z(o[3060]) );
  AND U7712 ( .A(p_input[305]), .B(p_input[10305]), .Z(o[305]) );
  AND U7713 ( .A(p_input[3059]), .B(p_input[13059]), .Z(o[3059]) );
  AND U7714 ( .A(p_input[3058]), .B(p_input[13058]), .Z(o[3058]) );
  AND U7715 ( .A(p_input[3057]), .B(p_input[13057]), .Z(o[3057]) );
  AND U7716 ( .A(p_input[3056]), .B(p_input[13056]), .Z(o[3056]) );
  AND U7717 ( .A(p_input[3055]), .B(p_input[13055]), .Z(o[3055]) );
  AND U7718 ( .A(p_input[3054]), .B(p_input[13054]), .Z(o[3054]) );
  AND U7719 ( .A(p_input[3053]), .B(p_input[13053]), .Z(o[3053]) );
  AND U7720 ( .A(p_input[3052]), .B(p_input[13052]), .Z(o[3052]) );
  AND U7721 ( .A(p_input[3051]), .B(p_input[13051]), .Z(o[3051]) );
  AND U7722 ( .A(p_input[3050]), .B(p_input[13050]), .Z(o[3050]) );
  AND U7723 ( .A(p_input[304]), .B(p_input[10304]), .Z(o[304]) );
  AND U7724 ( .A(p_input[3049]), .B(p_input[13049]), .Z(o[3049]) );
  AND U7725 ( .A(p_input[3048]), .B(p_input[13048]), .Z(o[3048]) );
  AND U7726 ( .A(p_input[3047]), .B(p_input[13047]), .Z(o[3047]) );
  AND U7727 ( .A(p_input[3046]), .B(p_input[13046]), .Z(o[3046]) );
  AND U7728 ( .A(p_input[3045]), .B(p_input[13045]), .Z(o[3045]) );
  AND U7729 ( .A(p_input[3044]), .B(p_input[13044]), .Z(o[3044]) );
  AND U7730 ( .A(p_input[3043]), .B(p_input[13043]), .Z(o[3043]) );
  AND U7731 ( .A(p_input[3042]), .B(p_input[13042]), .Z(o[3042]) );
  AND U7732 ( .A(p_input[3041]), .B(p_input[13041]), .Z(o[3041]) );
  AND U7733 ( .A(p_input[3040]), .B(p_input[13040]), .Z(o[3040]) );
  AND U7734 ( .A(p_input[303]), .B(p_input[10303]), .Z(o[303]) );
  AND U7735 ( .A(p_input[3039]), .B(p_input[13039]), .Z(o[3039]) );
  AND U7736 ( .A(p_input[3038]), .B(p_input[13038]), .Z(o[3038]) );
  AND U7737 ( .A(p_input[3037]), .B(p_input[13037]), .Z(o[3037]) );
  AND U7738 ( .A(p_input[3036]), .B(p_input[13036]), .Z(o[3036]) );
  AND U7739 ( .A(p_input[3035]), .B(p_input[13035]), .Z(o[3035]) );
  AND U7740 ( .A(p_input[3034]), .B(p_input[13034]), .Z(o[3034]) );
  AND U7741 ( .A(p_input[3033]), .B(p_input[13033]), .Z(o[3033]) );
  AND U7742 ( .A(p_input[3032]), .B(p_input[13032]), .Z(o[3032]) );
  AND U7743 ( .A(p_input[3031]), .B(p_input[13031]), .Z(o[3031]) );
  AND U7744 ( .A(p_input[3030]), .B(p_input[13030]), .Z(o[3030]) );
  AND U7745 ( .A(p_input[302]), .B(p_input[10302]), .Z(o[302]) );
  AND U7746 ( .A(p_input[3029]), .B(p_input[13029]), .Z(o[3029]) );
  AND U7747 ( .A(p_input[3028]), .B(p_input[13028]), .Z(o[3028]) );
  AND U7748 ( .A(p_input[3027]), .B(p_input[13027]), .Z(o[3027]) );
  AND U7749 ( .A(p_input[3026]), .B(p_input[13026]), .Z(o[3026]) );
  AND U7750 ( .A(p_input[3025]), .B(p_input[13025]), .Z(o[3025]) );
  AND U7751 ( .A(p_input[3024]), .B(p_input[13024]), .Z(o[3024]) );
  AND U7752 ( .A(p_input[3023]), .B(p_input[13023]), .Z(o[3023]) );
  AND U7753 ( .A(p_input[3022]), .B(p_input[13022]), .Z(o[3022]) );
  AND U7754 ( .A(p_input[3021]), .B(p_input[13021]), .Z(o[3021]) );
  AND U7755 ( .A(p_input[3020]), .B(p_input[13020]), .Z(o[3020]) );
  AND U7756 ( .A(p_input[301]), .B(p_input[10301]), .Z(o[301]) );
  AND U7757 ( .A(p_input[3019]), .B(p_input[13019]), .Z(o[3019]) );
  AND U7758 ( .A(p_input[3018]), .B(p_input[13018]), .Z(o[3018]) );
  AND U7759 ( .A(p_input[3017]), .B(p_input[13017]), .Z(o[3017]) );
  AND U7760 ( .A(p_input[3016]), .B(p_input[13016]), .Z(o[3016]) );
  AND U7761 ( .A(p_input[3015]), .B(p_input[13015]), .Z(o[3015]) );
  AND U7762 ( .A(p_input[3014]), .B(p_input[13014]), .Z(o[3014]) );
  AND U7763 ( .A(p_input[3013]), .B(p_input[13013]), .Z(o[3013]) );
  AND U7764 ( .A(p_input[3012]), .B(p_input[13012]), .Z(o[3012]) );
  AND U7765 ( .A(p_input[3011]), .B(p_input[13011]), .Z(o[3011]) );
  AND U7766 ( .A(p_input[3010]), .B(p_input[13010]), .Z(o[3010]) );
  AND U7767 ( .A(p_input[300]), .B(p_input[10300]), .Z(o[300]) );
  AND U7768 ( .A(p_input[3009]), .B(p_input[13009]), .Z(o[3009]) );
  AND U7769 ( .A(p_input[3008]), .B(p_input[13008]), .Z(o[3008]) );
  AND U7770 ( .A(p_input[3007]), .B(p_input[13007]), .Z(o[3007]) );
  AND U7771 ( .A(p_input[3006]), .B(p_input[13006]), .Z(o[3006]) );
  AND U7772 ( .A(p_input[3005]), .B(p_input[13005]), .Z(o[3005]) );
  AND U7773 ( .A(p_input[3004]), .B(p_input[13004]), .Z(o[3004]) );
  AND U7774 ( .A(p_input[3003]), .B(p_input[13003]), .Z(o[3003]) );
  AND U7775 ( .A(p_input[3002]), .B(p_input[13002]), .Z(o[3002]) );
  AND U7776 ( .A(p_input[3001]), .B(p_input[13001]), .Z(o[3001]) );
  AND U7777 ( .A(p_input[3000]), .B(p_input[13000]), .Z(o[3000]) );
  AND U7778 ( .A(p_input[2]), .B(p_input[10002]), .Z(o[2]) );
  AND U7779 ( .A(p_input[29]), .B(p_input[10029]), .Z(o[29]) );
  AND U7780 ( .A(p_input[299]), .B(p_input[10299]), .Z(o[299]) );
  AND U7781 ( .A(p_input[2999]), .B(p_input[12999]), .Z(o[2999]) );
  AND U7782 ( .A(p_input[2998]), .B(p_input[12998]), .Z(o[2998]) );
  AND U7783 ( .A(p_input[2997]), .B(p_input[12997]), .Z(o[2997]) );
  AND U7784 ( .A(p_input[2996]), .B(p_input[12996]), .Z(o[2996]) );
  AND U7785 ( .A(p_input[2995]), .B(p_input[12995]), .Z(o[2995]) );
  AND U7786 ( .A(p_input[2994]), .B(p_input[12994]), .Z(o[2994]) );
  AND U7787 ( .A(p_input[2993]), .B(p_input[12993]), .Z(o[2993]) );
  AND U7788 ( .A(p_input[2992]), .B(p_input[12992]), .Z(o[2992]) );
  AND U7789 ( .A(p_input[2991]), .B(p_input[12991]), .Z(o[2991]) );
  AND U7790 ( .A(p_input[2990]), .B(p_input[12990]), .Z(o[2990]) );
  AND U7791 ( .A(p_input[298]), .B(p_input[10298]), .Z(o[298]) );
  AND U7792 ( .A(p_input[2989]), .B(p_input[12989]), .Z(o[2989]) );
  AND U7793 ( .A(p_input[2988]), .B(p_input[12988]), .Z(o[2988]) );
  AND U7794 ( .A(p_input[2987]), .B(p_input[12987]), .Z(o[2987]) );
  AND U7795 ( .A(p_input[2986]), .B(p_input[12986]), .Z(o[2986]) );
  AND U7796 ( .A(p_input[2985]), .B(p_input[12985]), .Z(o[2985]) );
  AND U7797 ( .A(p_input[2984]), .B(p_input[12984]), .Z(o[2984]) );
  AND U7798 ( .A(p_input[2983]), .B(p_input[12983]), .Z(o[2983]) );
  AND U7799 ( .A(p_input[2982]), .B(p_input[12982]), .Z(o[2982]) );
  AND U7800 ( .A(p_input[2981]), .B(p_input[12981]), .Z(o[2981]) );
  AND U7801 ( .A(p_input[2980]), .B(p_input[12980]), .Z(o[2980]) );
  AND U7802 ( .A(p_input[297]), .B(p_input[10297]), .Z(o[297]) );
  AND U7803 ( .A(p_input[2979]), .B(p_input[12979]), .Z(o[2979]) );
  AND U7804 ( .A(p_input[2978]), .B(p_input[12978]), .Z(o[2978]) );
  AND U7805 ( .A(p_input[2977]), .B(p_input[12977]), .Z(o[2977]) );
  AND U7806 ( .A(p_input[2976]), .B(p_input[12976]), .Z(o[2976]) );
  AND U7807 ( .A(p_input[2975]), .B(p_input[12975]), .Z(o[2975]) );
  AND U7808 ( .A(p_input[2974]), .B(p_input[12974]), .Z(o[2974]) );
  AND U7809 ( .A(p_input[2973]), .B(p_input[12973]), .Z(o[2973]) );
  AND U7810 ( .A(p_input[2972]), .B(p_input[12972]), .Z(o[2972]) );
  AND U7811 ( .A(p_input[2971]), .B(p_input[12971]), .Z(o[2971]) );
  AND U7812 ( .A(p_input[2970]), .B(p_input[12970]), .Z(o[2970]) );
  AND U7813 ( .A(p_input[296]), .B(p_input[10296]), .Z(o[296]) );
  AND U7814 ( .A(p_input[2969]), .B(p_input[12969]), .Z(o[2969]) );
  AND U7815 ( .A(p_input[2968]), .B(p_input[12968]), .Z(o[2968]) );
  AND U7816 ( .A(p_input[2967]), .B(p_input[12967]), .Z(o[2967]) );
  AND U7817 ( .A(p_input[2966]), .B(p_input[12966]), .Z(o[2966]) );
  AND U7818 ( .A(p_input[2965]), .B(p_input[12965]), .Z(o[2965]) );
  AND U7819 ( .A(p_input[2964]), .B(p_input[12964]), .Z(o[2964]) );
  AND U7820 ( .A(p_input[2963]), .B(p_input[12963]), .Z(o[2963]) );
  AND U7821 ( .A(p_input[2962]), .B(p_input[12962]), .Z(o[2962]) );
  AND U7822 ( .A(p_input[2961]), .B(p_input[12961]), .Z(o[2961]) );
  AND U7823 ( .A(p_input[2960]), .B(p_input[12960]), .Z(o[2960]) );
  AND U7824 ( .A(p_input[295]), .B(p_input[10295]), .Z(o[295]) );
  AND U7825 ( .A(p_input[2959]), .B(p_input[12959]), .Z(o[2959]) );
  AND U7826 ( .A(p_input[2958]), .B(p_input[12958]), .Z(o[2958]) );
  AND U7827 ( .A(p_input[2957]), .B(p_input[12957]), .Z(o[2957]) );
  AND U7828 ( .A(p_input[2956]), .B(p_input[12956]), .Z(o[2956]) );
  AND U7829 ( .A(p_input[2955]), .B(p_input[12955]), .Z(o[2955]) );
  AND U7830 ( .A(p_input[2954]), .B(p_input[12954]), .Z(o[2954]) );
  AND U7831 ( .A(p_input[2953]), .B(p_input[12953]), .Z(o[2953]) );
  AND U7832 ( .A(p_input[2952]), .B(p_input[12952]), .Z(o[2952]) );
  AND U7833 ( .A(p_input[2951]), .B(p_input[12951]), .Z(o[2951]) );
  AND U7834 ( .A(p_input[2950]), .B(p_input[12950]), .Z(o[2950]) );
  AND U7835 ( .A(p_input[294]), .B(p_input[10294]), .Z(o[294]) );
  AND U7836 ( .A(p_input[2949]), .B(p_input[12949]), .Z(o[2949]) );
  AND U7837 ( .A(p_input[2948]), .B(p_input[12948]), .Z(o[2948]) );
  AND U7838 ( .A(p_input[2947]), .B(p_input[12947]), .Z(o[2947]) );
  AND U7839 ( .A(p_input[2946]), .B(p_input[12946]), .Z(o[2946]) );
  AND U7840 ( .A(p_input[2945]), .B(p_input[12945]), .Z(o[2945]) );
  AND U7841 ( .A(p_input[2944]), .B(p_input[12944]), .Z(o[2944]) );
  AND U7842 ( .A(p_input[2943]), .B(p_input[12943]), .Z(o[2943]) );
  AND U7843 ( .A(p_input[2942]), .B(p_input[12942]), .Z(o[2942]) );
  AND U7844 ( .A(p_input[2941]), .B(p_input[12941]), .Z(o[2941]) );
  AND U7845 ( .A(p_input[2940]), .B(p_input[12940]), .Z(o[2940]) );
  AND U7846 ( .A(p_input[293]), .B(p_input[10293]), .Z(o[293]) );
  AND U7847 ( .A(p_input[2939]), .B(p_input[12939]), .Z(o[2939]) );
  AND U7848 ( .A(p_input[2938]), .B(p_input[12938]), .Z(o[2938]) );
  AND U7849 ( .A(p_input[2937]), .B(p_input[12937]), .Z(o[2937]) );
  AND U7850 ( .A(p_input[2936]), .B(p_input[12936]), .Z(o[2936]) );
  AND U7851 ( .A(p_input[2935]), .B(p_input[12935]), .Z(o[2935]) );
  AND U7852 ( .A(p_input[2934]), .B(p_input[12934]), .Z(o[2934]) );
  AND U7853 ( .A(p_input[2933]), .B(p_input[12933]), .Z(o[2933]) );
  AND U7854 ( .A(p_input[2932]), .B(p_input[12932]), .Z(o[2932]) );
  AND U7855 ( .A(p_input[2931]), .B(p_input[12931]), .Z(o[2931]) );
  AND U7856 ( .A(p_input[2930]), .B(p_input[12930]), .Z(o[2930]) );
  AND U7857 ( .A(p_input[292]), .B(p_input[10292]), .Z(o[292]) );
  AND U7858 ( .A(p_input[2929]), .B(p_input[12929]), .Z(o[2929]) );
  AND U7859 ( .A(p_input[2928]), .B(p_input[12928]), .Z(o[2928]) );
  AND U7860 ( .A(p_input[2927]), .B(p_input[12927]), .Z(o[2927]) );
  AND U7861 ( .A(p_input[2926]), .B(p_input[12926]), .Z(o[2926]) );
  AND U7862 ( .A(p_input[2925]), .B(p_input[12925]), .Z(o[2925]) );
  AND U7863 ( .A(p_input[2924]), .B(p_input[12924]), .Z(o[2924]) );
  AND U7864 ( .A(p_input[2923]), .B(p_input[12923]), .Z(o[2923]) );
  AND U7865 ( .A(p_input[2922]), .B(p_input[12922]), .Z(o[2922]) );
  AND U7866 ( .A(p_input[2921]), .B(p_input[12921]), .Z(o[2921]) );
  AND U7867 ( .A(p_input[2920]), .B(p_input[12920]), .Z(o[2920]) );
  AND U7868 ( .A(p_input[291]), .B(p_input[10291]), .Z(o[291]) );
  AND U7869 ( .A(p_input[2919]), .B(p_input[12919]), .Z(o[2919]) );
  AND U7870 ( .A(p_input[2918]), .B(p_input[12918]), .Z(o[2918]) );
  AND U7871 ( .A(p_input[2917]), .B(p_input[12917]), .Z(o[2917]) );
  AND U7872 ( .A(p_input[2916]), .B(p_input[12916]), .Z(o[2916]) );
  AND U7873 ( .A(p_input[2915]), .B(p_input[12915]), .Z(o[2915]) );
  AND U7874 ( .A(p_input[2914]), .B(p_input[12914]), .Z(o[2914]) );
  AND U7875 ( .A(p_input[2913]), .B(p_input[12913]), .Z(o[2913]) );
  AND U7876 ( .A(p_input[2912]), .B(p_input[12912]), .Z(o[2912]) );
  AND U7877 ( .A(p_input[2911]), .B(p_input[12911]), .Z(o[2911]) );
  AND U7878 ( .A(p_input[2910]), .B(p_input[12910]), .Z(o[2910]) );
  AND U7879 ( .A(p_input[290]), .B(p_input[10290]), .Z(o[290]) );
  AND U7880 ( .A(p_input[2909]), .B(p_input[12909]), .Z(o[2909]) );
  AND U7881 ( .A(p_input[2908]), .B(p_input[12908]), .Z(o[2908]) );
  AND U7882 ( .A(p_input[2907]), .B(p_input[12907]), .Z(o[2907]) );
  AND U7883 ( .A(p_input[2906]), .B(p_input[12906]), .Z(o[2906]) );
  AND U7884 ( .A(p_input[2905]), .B(p_input[12905]), .Z(o[2905]) );
  AND U7885 ( .A(p_input[2904]), .B(p_input[12904]), .Z(o[2904]) );
  AND U7886 ( .A(p_input[2903]), .B(p_input[12903]), .Z(o[2903]) );
  AND U7887 ( .A(p_input[2902]), .B(p_input[12902]), .Z(o[2902]) );
  AND U7888 ( .A(p_input[2901]), .B(p_input[12901]), .Z(o[2901]) );
  AND U7889 ( .A(p_input[2900]), .B(p_input[12900]), .Z(o[2900]) );
  AND U7890 ( .A(p_input[28]), .B(p_input[10028]), .Z(o[28]) );
  AND U7891 ( .A(p_input[289]), .B(p_input[10289]), .Z(o[289]) );
  AND U7892 ( .A(p_input[2899]), .B(p_input[12899]), .Z(o[2899]) );
  AND U7893 ( .A(p_input[2898]), .B(p_input[12898]), .Z(o[2898]) );
  AND U7894 ( .A(p_input[2897]), .B(p_input[12897]), .Z(o[2897]) );
  AND U7895 ( .A(p_input[2896]), .B(p_input[12896]), .Z(o[2896]) );
  AND U7896 ( .A(p_input[2895]), .B(p_input[12895]), .Z(o[2895]) );
  AND U7897 ( .A(p_input[2894]), .B(p_input[12894]), .Z(o[2894]) );
  AND U7898 ( .A(p_input[2893]), .B(p_input[12893]), .Z(o[2893]) );
  AND U7899 ( .A(p_input[2892]), .B(p_input[12892]), .Z(o[2892]) );
  AND U7900 ( .A(p_input[2891]), .B(p_input[12891]), .Z(o[2891]) );
  AND U7901 ( .A(p_input[2890]), .B(p_input[12890]), .Z(o[2890]) );
  AND U7902 ( .A(p_input[288]), .B(p_input[10288]), .Z(o[288]) );
  AND U7903 ( .A(p_input[2889]), .B(p_input[12889]), .Z(o[2889]) );
  AND U7904 ( .A(p_input[2888]), .B(p_input[12888]), .Z(o[2888]) );
  AND U7905 ( .A(p_input[2887]), .B(p_input[12887]), .Z(o[2887]) );
  AND U7906 ( .A(p_input[2886]), .B(p_input[12886]), .Z(o[2886]) );
  AND U7907 ( .A(p_input[2885]), .B(p_input[12885]), .Z(o[2885]) );
  AND U7908 ( .A(p_input[2884]), .B(p_input[12884]), .Z(o[2884]) );
  AND U7909 ( .A(p_input[2883]), .B(p_input[12883]), .Z(o[2883]) );
  AND U7910 ( .A(p_input[2882]), .B(p_input[12882]), .Z(o[2882]) );
  AND U7911 ( .A(p_input[2881]), .B(p_input[12881]), .Z(o[2881]) );
  AND U7912 ( .A(p_input[2880]), .B(p_input[12880]), .Z(o[2880]) );
  AND U7913 ( .A(p_input[287]), .B(p_input[10287]), .Z(o[287]) );
  AND U7914 ( .A(p_input[2879]), .B(p_input[12879]), .Z(o[2879]) );
  AND U7915 ( .A(p_input[2878]), .B(p_input[12878]), .Z(o[2878]) );
  AND U7916 ( .A(p_input[2877]), .B(p_input[12877]), .Z(o[2877]) );
  AND U7917 ( .A(p_input[2876]), .B(p_input[12876]), .Z(o[2876]) );
  AND U7918 ( .A(p_input[2875]), .B(p_input[12875]), .Z(o[2875]) );
  AND U7919 ( .A(p_input[2874]), .B(p_input[12874]), .Z(o[2874]) );
  AND U7920 ( .A(p_input[2873]), .B(p_input[12873]), .Z(o[2873]) );
  AND U7921 ( .A(p_input[2872]), .B(p_input[12872]), .Z(o[2872]) );
  AND U7922 ( .A(p_input[2871]), .B(p_input[12871]), .Z(o[2871]) );
  AND U7923 ( .A(p_input[2870]), .B(p_input[12870]), .Z(o[2870]) );
  AND U7924 ( .A(p_input[286]), .B(p_input[10286]), .Z(o[286]) );
  AND U7925 ( .A(p_input[2869]), .B(p_input[12869]), .Z(o[2869]) );
  AND U7926 ( .A(p_input[2868]), .B(p_input[12868]), .Z(o[2868]) );
  AND U7927 ( .A(p_input[2867]), .B(p_input[12867]), .Z(o[2867]) );
  AND U7928 ( .A(p_input[2866]), .B(p_input[12866]), .Z(o[2866]) );
  AND U7929 ( .A(p_input[2865]), .B(p_input[12865]), .Z(o[2865]) );
  AND U7930 ( .A(p_input[2864]), .B(p_input[12864]), .Z(o[2864]) );
  AND U7931 ( .A(p_input[2863]), .B(p_input[12863]), .Z(o[2863]) );
  AND U7932 ( .A(p_input[2862]), .B(p_input[12862]), .Z(o[2862]) );
  AND U7933 ( .A(p_input[2861]), .B(p_input[12861]), .Z(o[2861]) );
  AND U7934 ( .A(p_input[2860]), .B(p_input[12860]), .Z(o[2860]) );
  AND U7935 ( .A(p_input[285]), .B(p_input[10285]), .Z(o[285]) );
  AND U7936 ( .A(p_input[2859]), .B(p_input[12859]), .Z(o[2859]) );
  AND U7937 ( .A(p_input[2858]), .B(p_input[12858]), .Z(o[2858]) );
  AND U7938 ( .A(p_input[2857]), .B(p_input[12857]), .Z(o[2857]) );
  AND U7939 ( .A(p_input[2856]), .B(p_input[12856]), .Z(o[2856]) );
  AND U7940 ( .A(p_input[2855]), .B(p_input[12855]), .Z(o[2855]) );
  AND U7941 ( .A(p_input[2854]), .B(p_input[12854]), .Z(o[2854]) );
  AND U7942 ( .A(p_input[2853]), .B(p_input[12853]), .Z(o[2853]) );
  AND U7943 ( .A(p_input[2852]), .B(p_input[12852]), .Z(o[2852]) );
  AND U7944 ( .A(p_input[2851]), .B(p_input[12851]), .Z(o[2851]) );
  AND U7945 ( .A(p_input[2850]), .B(p_input[12850]), .Z(o[2850]) );
  AND U7946 ( .A(p_input[284]), .B(p_input[10284]), .Z(o[284]) );
  AND U7947 ( .A(p_input[2849]), .B(p_input[12849]), .Z(o[2849]) );
  AND U7948 ( .A(p_input[2848]), .B(p_input[12848]), .Z(o[2848]) );
  AND U7949 ( .A(p_input[2847]), .B(p_input[12847]), .Z(o[2847]) );
  AND U7950 ( .A(p_input[2846]), .B(p_input[12846]), .Z(o[2846]) );
  AND U7951 ( .A(p_input[2845]), .B(p_input[12845]), .Z(o[2845]) );
  AND U7952 ( .A(p_input[2844]), .B(p_input[12844]), .Z(o[2844]) );
  AND U7953 ( .A(p_input[2843]), .B(p_input[12843]), .Z(o[2843]) );
  AND U7954 ( .A(p_input[2842]), .B(p_input[12842]), .Z(o[2842]) );
  AND U7955 ( .A(p_input[2841]), .B(p_input[12841]), .Z(o[2841]) );
  AND U7956 ( .A(p_input[2840]), .B(p_input[12840]), .Z(o[2840]) );
  AND U7957 ( .A(p_input[283]), .B(p_input[10283]), .Z(o[283]) );
  AND U7958 ( .A(p_input[2839]), .B(p_input[12839]), .Z(o[2839]) );
  AND U7959 ( .A(p_input[2838]), .B(p_input[12838]), .Z(o[2838]) );
  AND U7960 ( .A(p_input[2837]), .B(p_input[12837]), .Z(o[2837]) );
  AND U7961 ( .A(p_input[2836]), .B(p_input[12836]), .Z(o[2836]) );
  AND U7962 ( .A(p_input[2835]), .B(p_input[12835]), .Z(o[2835]) );
  AND U7963 ( .A(p_input[2834]), .B(p_input[12834]), .Z(o[2834]) );
  AND U7964 ( .A(p_input[2833]), .B(p_input[12833]), .Z(o[2833]) );
  AND U7965 ( .A(p_input[2832]), .B(p_input[12832]), .Z(o[2832]) );
  AND U7966 ( .A(p_input[2831]), .B(p_input[12831]), .Z(o[2831]) );
  AND U7967 ( .A(p_input[2830]), .B(p_input[12830]), .Z(o[2830]) );
  AND U7968 ( .A(p_input[282]), .B(p_input[10282]), .Z(o[282]) );
  AND U7969 ( .A(p_input[2829]), .B(p_input[12829]), .Z(o[2829]) );
  AND U7970 ( .A(p_input[2828]), .B(p_input[12828]), .Z(o[2828]) );
  AND U7971 ( .A(p_input[2827]), .B(p_input[12827]), .Z(o[2827]) );
  AND U7972 ( .A(p_input[2826]), .B(p_input[12826]), .Z(o[2826]) );
  AND U7973 ( .A(p_input[2825]), .B(p_input[12825]), .Z(o[2825]) );
  AND U7974 ( .A(p_input[2824]), .B(p_input[12824]), .Z(o[2824]) );
  AND U7975 ( .A(p_input[2823]), .B(p_input[12823]), .Z(o[2823]) );
  AND U7976 ( .A(p_input[2822]), .B(p_input[12822]), .Z(o[2822]) );
  AND U7977 ( .A(p_input[2821]), .B(p_input[12821]), .Z(o[2821]) );
  AND U7978 ( .A(p_input[2820]), .B(p_input[12820]), .Z(o[2820]) );
  AND U7979 ( .A(p_input[281]), .B(p_input[10281]), .Z(o[281]) );
  AND U7980 ( .A(p_input[2819]), .B(p_input[12819]), .Z(o[2819]) );
  AND U7981 ( .A(p_input[2818]), .B(p_input[12818]), .Z(o[2818]) );
  AND U7982 ( .A(p_input[2817]), .B(p_input[12817]), .Z(o[2817]) );
  AND U7983 ( .A(p_input[2816]), .B(p_input[12816]), .Z(o[2816]) );
  AND U7984 ( .A(p_input[2815]), .B(p_input[12815]), .Z(o[2815]) );
  AND U7985 ( .A(p_input[2814]), .B(p_input[12814]), .Z(o[2814]) );
  AND U7986 ( .A(p_input[2813]), .B(p_input[12813]), .Z(o[2813]) );
  AND U7987 ( .A(p_input[2812]), .B(p_input[12812]), .Z(o[2812]) );
  AND U7988 ( .A(p_input[2811]), .B(p_input[12811]), .Z(o[2811]) );
  AND U7989 ( .A(p_input[2810]), .B(p_input[12810]), .Z(o[2810]) );
  AND U7990 ( .A(p_input[280]), .B(p_input[10280]), .Z(o[280]) );
  AND U7991 ( .A(p_input[2809]), .B(p_input[12809]), .Z(o[2809]) );
  AND U7992 ( .A(p_input[2808]), .B(p_input[12808]), .Z(o[2808]) );
  AND U7993 ( .A(p_input[2807]), .B(p_input[12807]), .Z(o[2807]) );
  AND U7994 ( .A(p_input[2806]), .B(p_input[12806]), .Z(o[2806]) );
  AND U7995 ( .A(p_input[2805]), .B(p_input[12805]), .Z(o[2805]) );
  AND U7996 ( .A(p_input[2804]), .B(p_input[12804]), .Z(o[2804]) );
  AND U7997 ( .A(p_input[2803]), .B(p_input[12803]), .Z(o[2803]) );
  AND U7998 ( .A(p_input[2802]), .B(p_input[12802]), .Z(o[2802]) );
  AND U7999 ( .A(p_input[2801]), .B(p_input[12801]), .Z(o[2801]) );
  AND U8000 ( .A(p_input[2800]), .B(p_input[12800]), .Z(o[2800]) );
  AND U8001 ( .A(p_input[27]), .B(p_input[10027]), .Z(o[27]) );
  AND U8002 ( .A(p_input[279]), .B(p_input[10279]), .Z(o[279]) );
  AND U8003 ( .A(p_input[2799]), .B(p_input[12799]), .Z(o[2799]) );
  AND U8004 ( .A(p_input[2798]), .B(p_input[12798]), .Z(o[2798]) );
  AND U8005 ( .A(p_input[2797]), .B(p_input[12797]), .Z(o[2797]) );
  AND U8006 ( .A(p_input[2796]), .B(p_input[12796]), .Z(o[2796]) );
  AND U8007 ( .A(p_input[2795]), .B(p_input[12795]), .Z(o[2795]) );
  AND U8008 ( .A(p_input[2794]), .B(p_input[12794]), .Z(o[2794]) );
  AND U8009 ( .A(p_input[2793]), .B(p_input[12793]), .Z(o[2793]) );
  AND U8010 ( .A(p_input[2792]), .B(p_input[12792]), .Z(o[2792]) );
  AND U8011 ( .A(p_input[2791]), .B(p_input[12791]), .Z(o[2791]) );
  AND U8012 ( .A(p_input[2790]), .B(p_input[12790]), .Z(o[2790]) );
  AND U8013 ( .A(p_input[278]), .B(p_input[10278]), .Z(o[278]) );
  AND U8014 ( .A(p_input[2789]), .B(p_input[12789]), .Z(o[2789]) );
  AND U8015 ( .A(p_input[2788]), .B(p_input[12788]), .Z(o[2788]) );
  AND U8016 ( .A(p_input[2787]), .B(p_input[12787]), .Z(o[2787]) );
  AND U8017 ( .A(p_input[2786]), .B(p_input[12786]), .Z(o[2786]) );
  AND U8018 ( .A(p_input[2785]), .B(p_input[12785]), .Z(o[2785]) );
  AND U8019 ( .A(p_input[2784]), .B(p_input[12784]), .Z(o[2784]) );
  AND U8020 ( .A(p_input[2783]), .B(p_input[12783]), .Z(o[2783]) );
  AND U8021 ( .A(p_input[2782]), .B(p_input[12782]), .Z(o[2782]) );
  AND U8022 ( .A(p_input[2781]), .B(p_input[12781]), .Z(o[2781]) );
  AND U8023 ( .A(p_input[2780]), .B(p_input[12780]), .Z(o[2780]) );
  AND U8024 ( .A(p_input[277]), .B(p_input[10277]), .Z(o[277]) );
  AND U8025 ( .A(p_input[2779]), .B(p_input[12779]), .Z(o[2779]) );
  AND U8026 ( .A(p_input[2778]), .B(p_input[12778]), .Z(o[2778]) );
  AND U8027 ( .A(p_input[2777]), .B(p_input[12777]), .Z(o[2777]) );
  AND U8028 ( .A(p_input[2776]), .B(p_input[12776]), .Z(o[2776]) );
  AND U8029 ( .A(p_input[2775]), .B(p_input[12775]), .Z(o[2775]) );
  AND U8030 ( .A(p_input[2774]), .B(p_input[12774]), .Z(o[2774]) );
  AND U8031 ( .A(p_input[2773]), .B(p_input[12773]), .Z(o[2773]) );
  AND U8032 ( .A(p_input[2772]), .B(p_input[12772]), .Z(o[2772]) );
  AND U8033 ( .A(p_input[2771]), .B(p_input[12771]), .Z(o[2771]) );
  AND U8034 ( .A(p_input[2770]), .B(p_input[12770]), .Z(o[2770]) );
  AND U8035 ( .A(p_input[276]), .B(p_input[10276]), .Z(o[276]) );
  AND U8036 ( .A(p_input[2769]), .B(p_input[12769]), .Z(o[2769]) );
  AND U8037 ( .A(p_input[2768]), .B(p_input[12768]), .Z(o[2768]) );
  AND U8038 ( .A(p_input[2767]), .B(p_input[12767]), .Z(o[2767]) );
  AND U8039 ( .A(p_input[2766]), .B(p_input[12766]), .Z(o[2766]) );
  AND U8040 ( .A(p_input[2765]), .B(p_input[12765]), .Z(o[2765]) );
  AND U8041 ( .A(p_input[2764]), .B(p_input[12764]), .Z(o[2764]) );
  AND U8042 ( .A(p_input[2763]), .B(p_input[12763]), .Z(o[2763]) );
  AND U8043 ( .A(p_input[2762]), .B(p_input[12762]), .Z(o[2762]) );
  AND U8044 ( .A(p_input[2761]), .B(p_input[12761]), .Z(o[2761]) );
  AND U8045 ( .A(p_input[2760]), .B(p_input[12760]), .Z(o[2760]) );
  AND U8046 ( .A(p_input[275]), .B(p_input[10275]), .Z(o[275]) );
  AND U8047 ( .A(p_input[2759]), .B(p_input[12759]), .Z(o[2759]) );
  AND U8048 ( .A(p_input[2758]), .B(p_input[12758]), .Z(o[2758]) );
  AND U8049 ( .A(p_input[2757]), .B(p_input[12757]), .Z(o[2757]) );
  AND U8050 ( .A(p_input[2756]), .B(p_input[12756]), .Z(o[2756]) );
  AND U8051 ( .A(p_input[2755]), .B(p_input[12755]), .Z(o[2755]) );
  AND U8052 ( .A(p_input[2754]), .B(p_input[12754]), .Z(o[2754]) );
  AND U8053 ( .A(p_input[2753]), .B(p_input[12753]), .Z(o[2753]) );
  AND U8054 ( .A(p_input[2752]), .B(p_input[12752]), .Z(o[2752]) );
  AND U8055 ( .A(p_input[2751]), .B(p_input[12751]), .Z(o[2751]) );
  AND U8056 ( .A(p_input[2750]), .B(p_input[12750]), .Z(o[2750]) );
  AND U8057 ( .A(p_input[274]), .B(p_input[10274]), .Z(o[274]) );
  AND U8058 ( .A(p_input[2749]), .B(p_input[12749]), .Z(o[2749]) );
  AND U8059 ( .A(p_input[2748]), .B(p_input[12748]), .Z(o[2748]) );
  AND U8060 ( .A(p_input[2747]), .B(p_input[12747]), .Z(o[2747]) );
  AND U8061 ( .A(p_input[2746]), .B(p_input[12746]), .Z(o[2746]) );
  AND U8062 ( .A(p_input[2745]), .B(p_input[12745]), .Z(o[2745]) );
  AND U8063 ( .A(p_input[2744]), .B(p_input[12744]), .Z(o[2744]) );
  AND U8064 ( .A(p_input[2743]), .B(p_input[12743]), .Z(o[2743]) );
  AND U8065 ( .A(p_input[2742]), .B(p_input[12742]), .Z(o[2742]) );
  AND U8066 ( .A(p_input[2741]), .B(p_input[12741]), .Z(o[2741]) );
  AND U8067 ( .A(p_input[2740]), .B(p_input[12740]), .Z(o[2740]) );
  AND U8068 ( .A(p_input[273]), .B(p_input[10273]), .Z(o[273]) );
  AND U8069 ( .A(p_input[2739]), .B(p_input[12739]), .Z(o[2739]) );
  AND U8070 ( .A(p_input[2738]), .B(p_input[12738]), .Z(o[2738]) );
  AND U8071 ( .A(p_input[2737]), .B(p_input[12737]), .Z(o[2737]) );
  AND U8072 ( .A(p_input[2736]), .B(p_input[12736]), .Z(o[2736]) );
  AND U8073 ( .A(p_input[2735]), .B(p_input[12735]), .Z(o[2735]) );
  AND U8074 ( .A(p_input[2734]), .B(p_input[12734]), .Z(o[2734]) );
  AND U8075 ( .A(p_input[2733]), .B(p_input[12733]), .Z(o[2733]) );
  AND U8076 ( .A(p_input[2732]), .B(p_input[12732]), .Z(o[2732]) );
  AND U8077 ( .A(p_input[2731]), .B(p_input[12731]), .Z(o[2731]) );
  AND U8078 ( .A(p_input[2730]), .B(p_input[12730]), .Z(o[2730]) );
  AND U8079 ( .A(p_input[272]), .B(p_input[10272]), .Z(o[272]) );
  AND U8080 ( .A(p_input[2729]), .B(p_input[12729]), .Z(o[2729]) );
  AND U8081 ( .A(p_input[2728]), .B(p_input[12728]), .Z(o[2728]) );
  AND U8082 ( .A(p_input[2727]), .B(p_input[12727]), .Z(o[2727]) );
  AND U8083 ( .A(p_input[2726]), .B(p_input[12726]), .Z(o[2726]) );
  AND U8084 ( .A(p_input[2725]), .B(p_input[12725]), .Z(o[2725]) );
  AND U8085 ( .A(p_input[2724]), .B(p_input[12724]), .Z(o[2724]) );
  AND U8086 ( .A(p_input[2723]), .B(p_input[12723]), .Z(o[2723]) );
  AND U8087 ( .A(p_input[2722]), .B(p_input[12722]), .Z(o[2722]) );
  AND U8088 ( .A(p_input[2721]), .B(p_input[12721]), .Z(o[2721]) );
  AND U8089 ( .A(p_input[2720]), .B(p_input[12720]), .Z(o[2720]) );
  AND U8090 ( .A(p_input[271]), .B(p_input[10271]), .Z(o[271]) );
  AND U8091 ( .A(p_input[2719]), .B(p_input[12719]), .Z(o[2719]) );
  AND U8092 ( .A(p_input[2718]), .B(p_input[12718]), .Z(o[2718]) );
  AND U8093 ( .A(p_input[2717]), .B(p_input[12717]), .Z(o[2717]) );
  AND U8094 ( .A(p_input[2716]), .B(p_input[12716]), .Z(o[2716]) );
  AND U8095 ( .A(p_input[2715]), .B(p_input[12715]), .Z(o[2715]) );
  AND U8096 ( .A(p_input[2714]), .B(p_input[12714]), .Z(o[2714]) );
  AND U8097 ( .A(p_input[2713]), .B(p_input[12713]), .Z(o[2713]) );
  AND U8098 ( .A(p_input[2712]), .B(p_input[12712]), .Z(o[2712]) );
  AND U8099 ( .A(p_input[2711]), .B(p_input[12711]), .Z(o[2711]) );
  AND U8100 ( .A(p_input[2710]), .B(p_input[12710]), .Z(o[2710]) );
  AND U8101 ( .A(p_input[270]), .B(p_input[10270]), .Z(o[270]) );
  AND U8102 ( .A(p_input[2709]), .B(p_input[12709]), .Z(o[2709]) );
  AND U8103 ( .A(p_input[2708]), .B(p_input[12708]), .Z(o[2708]) );
  AND U8104 ( .A(p_input[2707]), .B(p_input[12707]), .Z(o[2707]) );
  AND U8105 ( .A(p_input[2706]), .B(p_input[12706]), .Z(o[2706]) );
  AND U8106 ( .A(p_input[2705]), .B(p_input[12705]), .Z(o[2705]) );
  AND U8107 ( .A(p_input[2704]), .B(p_input[12704]), .Z(o[2704]) );
  AND U8108 ( .A(p_input[2703]), .B(p_input[12703]), .Z(o[2703]) );
  AND U8109 ( .A(p_input[2702]), .B(p_input[12702]), .Z(o[2702]) );
  AND U8110 ( .A(p_input[2701]), .B(p_input[12701]), .Z(o[2701]) );
  AND U8111 ( .A(p_input[2700]), .B(p_input[12700]), .Z(o[2700]) );
  AND U8112 ( .A(p_input[26]), .B(p_input[10026]), .Z(o[26]) );
  AND U8113 ( .A(p_input[269]), .B(p_input[10269]), .Z(o[269]) );
  AND U8114 ( .A(p_input[2699]), .B(p_input[12699]), .Z(o[2699]) );
  AND U8115 ( .A(p_input[2698]), .B(p_input[12698]), .Z(o[2698]) );
  AND U8116 ( .A(p_input[2697]), .B(p_input[12697]), .Z(o[2697]) );
  AND U8117 ( .A(p_input[2696]), .B(p_input[12696]), .Z(o[2696]) );
  AND U8118 ( .A(p_input[2695]), .B(p_input[12695]), .Z(o[2695]) );
  AND U8119 ( .A(p_input[2694]), .B(p_input[12694]), .Z(o[2694]) );
  AND U8120 ( .A(p_input[2693]), .B(p_input[12693]), .Z(o[2693]) );
  AND U8121 ( .A(p_input[2692]), .B(p_input[12692]), .Z(o[2692]) );
  AND U8122 ( .A(p_input[2691]), .B(p_input[12691]), .Z(o[2691]) );
  AND U8123 ( .A(p_input[2690]), .B(p_input[12690]), .Z(o[2690]) );
  AND U8124 ( .A(p_input[268]), .B(p_input[10268]), .Z(o[268]) );
  AND U8125 ( .A(p_input[2689]), .B(p_input[12689]), .Z(o[2689]) );
  AND U8126 ( .A(p_input[2688]), .B(p_input[12688]), .Z(o[2688]) );
  AND U8127 ( .A(p_input[2687]), .B(p_input[12687]), .Z(o[2687]) );
  AND U8128 ( .A(p_input[2686]), .B(p_input[12686]), .Z(o[2686]) );
  AND U8129 ( .A(p_input[2685]), .B(p_input[12685]), .Z(o[2685]) );
  AND U8130 ( .A(p_input[2684]), .B(p_input[12684]), .Z(o[2684]) );
  AND U8131 ( .A(p_input[2683]), .B(p_input[12683]), .Z(o[2683]) );
  AND U8132 ( .A(p_input[2682]), .B(p_input[12682]), .Z(o[2682]) );
  AND U8133 ( .A(p_input[2681]), .B(p_input[12681]), .Z(o[2681]) );
  AND U8134 ( .A(p_input[2680]), .B(p_input[12680]), .Z(o[2680]) );
  AND U8135 ( .A(p_input[267]), .B(p_input[10267]), .Z(o[267]) );
  AND U8136 ( .A(p_input[2679]), .B(p_input[12679]), .Z(o[2679]) );
  AND U8137 ( .A(p_input[2678]), .B(p_input[12678]), .Z(o[2678]) );
  AND U8138 ( .A(p_input[2677]), .B(p_input[12677]), .Z(o[2677]) );
  AND U8139 ( .A(p_input[2676]), .B(p_input[12676]), .Z(o[2676]) );
  AND U8140 ( .A(p_input[2675]), .B(p_input[12675]), .Z(o[2675]) );
  AND U8141 ( .A(p_input[2674]), .B(p_input[12674]), .Z(o[2674]) );
  AND U8142 ( .A(p_input[2673]), .B(p_input[12673]), .Z(o[2673]) );
  AND U8143 ( .A(p_input[2672]), .B(p_input[12672]), .Z(o[2672]) );
  AND U8144 ( .A(p_input[2671]), .B(p_input[12671]), .Z(o[2671]) );
  AND U8145 ( .A(p_input[2670]), .B(p_input[12670]), .Z(o[2670]) );
  AND U8146 ( .A(p_input[266]), .B(p_input[10266]), .Z(o[266]) );
  AND U8147 ( .A(p_input[2669]), .B(p_input[12669]), .Z(o[2669]) );
  AND U8148 ( .A(p_input[2668]), .B(p_input[12668]), .Z(o[2668]) );
  AND U8149 ( .A(p_input[2667]), .B(p_input[12667]), .Z(o[2667]) );
  AND U8150 ( .A(p_input[2666]), .B(p_input[12666]), .Z(o[2666]) );
  AND U8151 ( .A(p_input[2665]), .B(p_input[12665]), .Z(o[2665]) );
  AND U8152 ( .A(p_input[2664]), .B(p_input[12664]), .Z(o[2664]) );
  AND U8153 ( .A(p_input[2663]), .B(p_input[12663]), .Z(o[2663]) );
  AND U8154 ( .A(p_input[2662]), .B(p_input[12662]), .Z(o[2662]) );
  AND U8155 ( .A(p_input[2661]), .B(p_input[12661]), .Z(o[2661]) );
  AND U8156 ( .A(p_input[2660]), .B(p_input[12660]), .Z(o[2660]) );
  AND U8157 ( .A(p_input[265]), .B(p_input[10265]), .Z(o[265]) );
  AND U8158 ( .A(p_input[2659]), .B(p_input[12659]), .Z(o[2659]) );
  AND U8159 ( .A(p_input[2658]), .B(p_input[12658]), .Z(o[2658]) );
  AND U8160 ( .A(p_input[2657]), .B(p_input[12657]), .Z(o[2657]) );
  AND U8161 ( .A(p_input[2656]), .B(p_input[12656]), .Z(o[2656]) );
  AND U8162 ( .A(p_input[2655]), .B(p_input[12655]), .Z(o[2655]) );
  AND U8163 ( .A(p_input[2654]), .B(p_input[12654]), .Z(o[2654]) );
  AND U8164 ( .A(p_input[2653]), .B(p_input[12653]), .Z(o[2653]) );
  AND U8165 ( .A(p_input[2652]), .B(p_input[12652]), .Z(o[2652]) );
  AND U8166 ( .A(p_input[2651]), .B(p_input[12651]), .Z(o[2651]) );
  AND U8167 ( .A(p_input[2650]), .B(p_input[12650]), .Z(o[2650]) );
  AND U8168 ( .A(p_input[264]), .B(p_input[10264]), .Z(o[264]) );
  AND U8169 ( .A(p_input[2649]), .B(p_input[12649]), .Z(o[2649]) );
  AND U8170 ( .A(p_input[2648]), .B(p_input[12648]), .Z(o[2648]) );
  AND U8171 ( .A(p_input[2647]), .B(p_input[12647]), .Z(o[2647]) );
  AND U8172 ( .A(p_input[2646]), .B(p_input[12646]), .Z(o[2646]) );
  AND U8173 ( .A(p_input[2645]), .B(p_input[12645]), .Z(o[2645]) );
  AND U8174 ( .A(p_input[2644]), .B(p_input[12644]), .Z(o[2644]) );
  AND U8175 ( .A(p_input[2643]), .B(p_input[12643]), .Z(o[2643]) );
  AND U8176 ( .A(p_input[2642]), .B(p_input[12642]), .Z(o[2642]) );
  AND U8177 ( .A(p_input[2641]), .B(p_input[12641]), .Z(o[2641]) );
  AND U8178 ( .A(p_input[2640]), .B(p_input[12640]), .Z(o[2640]) );
  AND U8179 ( .A(p_input[263]), .B(p_input[10263]), .Z(o[263]) );
  AND U8180 ( .A(p_input[2639]), .B(p_input[12639]), .Z(o[2639]) );
  AND U8181 ( .A(p_input[2638]), .B(p_input[12638]), .Z(o[2638]) );
  AND U8182 ( .A(p_input[2637]), .B(p_input[12637]), .Z(o[2637]) );
  AND U8183 ( .A(p_input[2636]), .B(p_input[12636]), .Z(o[2636]) );
  AND U8184 ( .A(p_input[2635]), .B(p_input[12635]), .Z(o[2635]) );
  AND U8185 ( .A(p_input[2634]), .B(p_input[12634]), .Z(o[2634]) );
  AND U8186 ( .A(p_input[2633]), .B(p_input[12633]), .Z(o[2633]) );
  AND U8187 ( .A(p_input[2632]), .B(p_input[12632]), .Z(o[2632]) );
  AND U8188 ( .A(p_input[2631]), .B(p_input[12631]), .Z(o[2631]) );
  AND U8189 ( .A(p_input[2630]), .B(p_input[12630]), .Z(o[2630]) );
  AND U8190 ( .A(p_input[262]), .B(p_input[10262]), .Z(o[262]) );
  AND U8191 ( .A(p_input[2629]), .B(p_input[12629]), .Z(o[2629]) );
  AND U8192 ( .A(p_input[2628]), .B(p_input[12628]), .Z(o[2628]) );
  AND U8193 ( .A(p_input[2627]), .B(p_input[12627]), .Z(o[2627]) );
  AND U8194 ( .A(p_input[2626]), .B(p_input[12626]), .Z(o[2626]) );
  AND U8195 ( .A(p_input[2625]), .B(p_input[12625]), .Z(o[2625]) );
  AND U8196 ( .A(p_input[2624]), .B(p_input[12624]), .Z(o[2624]) );
  AND U8197 ( .A(p_input[2623]), .B(p_input[12623]), .Z(o[2623]) );
  AND U8198 ( .A(p_input[2622]), .B(p_input[12622]), .Z(o[2622]) );
  AND U8199 ( .A(p_input[2621]), .B(p_input[12621]), .Z(o[2621]) );
  AND U8200 ( .A(p_input[2620]), .B(p_input[12620]), .Z(o[2620]) );
  AND U8201 ( .A(p_input[261]), .B(p_input[10261]), .Z(o[261]) );
  AND U8202 ( .A(p_input[2619]), .B(p_input[12619]), .Z(o[2619]) );
  AND U8203 ( .A(p_input[2618]), .B(p_input[12618]), .Z(o[2618]) );
  AND U8204 ( .A(p_input[2617]), .B(p_input[12617]), .Z(o[2617]) );
  AND U8205 ( .A(p_input[2616]), .B(p_input[12616]), .Z(o[2616]) );
  AND U8206 ( .A(p_input[2615]), .B(p_input[12615]), .Z(o[2615]) );
  AND U8207 ( .A(p_input[2614]), .B(p_input[12614]), .Z(o[2614]) );
  AND U8208 ( .A(p_input[2613]), .B(p_input[12613]), .Z(o[2613]) );
  AND U8209 ( .A(p_input[2612]), .B(p_input[12612]), .Z(o[2612]) );
  AND U8210 ( .A(p_input[2611]), .B(p_input[12611]), .Z(o[2611]) );
  AND U8211 ( .A(p_input[2610]), .B(p_input[12610]), .Z(o[2610]) );
  AND U8212 ( .A(p_input[260]), .B(p_input[10260]), .Z(o[260]) );
  AND U8213 ( .A(p_input[2609]), .B(p_input[12609]), .Z(o[2609]) );
  AND U8214 ( .A(p_input[2608]), .B(p_input[12608]), .Z(o[2608]) );
  AND U8215 ( .A(p_input[2607]), .B(p_input[12607]), .Z(o[2607]) );
  AND U8216 ( .A(p_input[2606]), .B(p_input[12606]), .Z(o[2606]) );
  AND U8217 ( .A(p_input[2605]), .B(p_input[12605]), .Z(o[2605]) );
  AND U8218 ( .A(p_input[2604]), .B(p_input[12604]), .Z(o[2604]) );
  AND U8219 ( .A(p_input[2603]), .B(p_input[12603]), .Z(o[2603]) );
  AND U8220 ( .A(p_input[2602]), .B(p_input[12602]), .Z(o[2602]) );
  AND U8221 ( .A(p_input[2601]), .B(p_input[12601]), .Z(o[2601]) );
  AND U8222 ( .A(p_input[2600]), .B(p_input[12600]), .Z(o[2600]) );
  AND U8223 ( .A(p_input[25]), .B(p_input[10025]), .Z(o[25]) );
  AND U8224 ( .A(p_input[259]), .B(p_input[10259]), .Z(o[259]) );
  AND U8225 ( .A(p_input[2599]), .B(p_input[12599]), .Z(o[2599]) );
  AND U8226 ( .A(p_input[2598]), .B(p_input[12598]), .Z(o[2598]) );
  AND U8227 ( .A(p_input[2597]), .B(p_input[12597]), .Z(o[2597]) );
  AND U8228 ( .A(p_input[2596]), .B(p_input[12596]), .Z(o[2596]) );
  AND U8229 ( .A(p_input[2595]), .B(p_input[12595]), .Z(o[2595]) );
  AND U8230 ( .A(p_input[2594]), .B(p_input[12594]), .Z(o[2594]) );
  AND U8231 ( .A(p_input[2593]), .B(p_input[12593]), .Z(o[2593]) );
  AND U8232 ( .A(p_input[2592]), .B(p_input[12592]), .Z(o[2592]) );
  AND U8233 ( .A(p_input[2591]), .B(p_input[12591]), .Z(o[2591]) );
  AND U8234 ( .A(p_input[2590]), .B(p_input[12590]), .Z(o[2590]) );
  AND U8235 ( .A(p_input[258]), .B(p_input[10258]), .Z(o[258]) );
  AND U8236 ( .A(p_input[2589]), .B(p_input[12589]), .Z(o[2589]) );
  AND U8237 ( .A(p_input[2588]), .B(p_input[12588]), .Z(o[2588]) );
  AND U8238 ( .A(p_input[2587]), .B(p_input[12587]), .Z(o[2587]) );
  AND U8239 ( .A(p_input[2586]), .B(p_input[12586]), .Z(o[2586]) );
  AND U8240 ( .A(p_input[2585]), .B(p_input[12585]), .Z(o[2585]) );
  AND U8241 ( .A(p_input[2584]), .B(p_input[12584]), .Z(o[2584]) );
  AND U8242 ( .A(p_input[2583]), .B(p_input[12583]), .Z(o[2583]) );
  AND U8243 ( .A(p_input[2582]), .B(p_input[12582]), .Z(o[2582]) );
  AND U8244 ( .A(p_input[2581]), .B(p_input[12581]), .Z(o[2581]) );
  AND U8245 ( .A(p_input[2580]), .B(p_input[12580]), .Z(o[2580]) );
  AND U8246 ( .A(p_input[257]), .B(p_input[10257]), .Z(o[257]) );
  AND U8247 ( .A(p_input[2579]), .B(p_input[12579]), .Z(o[2579]) );
  AND U8248 ( .A(p_input[2578]), .B(p_input[12578]), .Z(o[2578]) );
  AND U8249 ( .A(p_input[2577]), .B(p_input[12577]), .Z(o[2577]) );
  AND U8250 ( .A(p_input[2576]), .B(p_input[12576]), .Z(o[2576]) );
  AND U8251 ( .A(p_input[2575]), .B(p_input[12575]), .Z(o[2575]) );
  AND U8252 ( .A(p_input[2574]), .B(p_input[12574]), .Z(o[2574]) );
  AND U8253 ( .A(p_input[2573]), .B(p_input[12573]), .Z(o[2573]) );
  AND U8254 ( .A(p_input[2572]), .B(p_input[12572]), .Z(o[2572]) );
  AND U8255 ( .A(p_input[2571]), .B(p_input[12571]), .Z(o[2571]) );
  AND U8256 ( .A(p_input[2570]), .B(p_input[12570]), .Z(o[2570]) );
  AND U8257 ( .A(p_input[256]), .B(p_input[10256]), .Z(o[256]) );
  AND U8258 ( .A(p_input[2569]), .B(p_input[12569]), .Z(o[2569]) );
  AND U8259 ( .A(p_input[2568]), .B(p_input[12568]), .Z(o[2568]) );
  AND U8260 ( .A(p_input[2567]), .B(p_input[12567]), .Z(o[2567]) );
  AND U8261 ( .A(p_input[2566]), .B(p_input[12566]), .Z(o[2566]) );
  AND U8262 ( .A(p_input[2565]), .B(p_input[12565]), .Z(o[2565]) );
  AND U8263 ( .A(p_input[2564]), .B(p_input[12564]), .Z(o[2564]) );
  AND U8264 ( .A(p_input[2563]), .B(p_input[12563]), .Z(o[2563]) );
  AND U8265 ( .A(p_input[2562]), .B(p_input[12562]), .Z(o[2562]) );
  AND U8266 ( .A(p_input[2561]), .B(p_input[12561]), .Z(o[2561]) );
  AND U8267 ( .A(p_input[2560]), .B(p_input[12560]), .Z(o[2560]) );
  AND U8268 ( .A(p_input[255]), .B(p_input[10255]), .Z(o[255]) );
  AND U8269 ( .A(p_input[2559]), .B(p_input[12559]), .Z(o[2559]) );
  AND U8270 ( .A(p_input[2558]), .B(p_input[12558]), .Z(o[2558]) );
  AND U8271 ( .A(p_input[2557]), .B(p_input[12557]), .Z(o[2557]) );
  AND U8272 ( .A(p_input[2556]), .B(p_input[12556]), .Z(o[2556]) );
  AND U8273 ( .A(p_input[2555]), .B(p_input[12555]), .Z(o[2555]) );
  AND U8274 ( .A(p_input[2554]), .B(p_input[12554]), .Z(o[2554]) );
  AND U8275 ( .A(p_input[2553]), .B(p_input[12553]), .Z(o[2553]) );
  AND U8276 ( .A(p_input[2552]), .B(p_input[12552]), .Z(o[2552]) );
  AND U8277 ( .A(p_input[2551]), .B(p_input[12551]), .Z(o[2551]) );
  AND U8278 ( .A(p_input[2550]), .B(p_input[12550]), .Z(o[2550]) );
  AND U8279 ( .A(p_input[254]), .B(p_input[10254]), .Z(o[254]) );
  AND U8280 ( .A(p_input[2549]), .B(p_input[12549]), .Z(o[2549]) );
  AND U8281 ( .A(p_input[2548]), .B(p_input[12548]), .Z(o[2548]) );
  AND U8282 ( .A(p_input[2547]), .B(p_input[12547]), .Z(o[2547]) );
  AND U8283 ( .A(p_input[2546]), .B(p_input[12546]), .Z(o[2546]) );
  AND U8284 ( .A(p_input[2545]), .B(p_input[12545]), .Z(o[2545]) );
  AND U8285 ( .A(p_input[2544]), .B(p_input[12544]), .Z(o[2544]) );
  AND U8286 ( .A(p_input[2543]), .B(p_input[12543]), .Z(o[2543]) );
  AND U8287 ( .A(p_input[2542]), .B(p_input[12542]), .Z(o[2542]) );
  AND U8288 ( .A(p_input[2541]), .B(p_input[12541]), .Z(o[2541]) );
  AND U8289 ( .A(p_input[2540]), .B(p_input[12540]), .Z(o[2540]) );
  AND U8290 ( .A(p_input[253]), .B(p_input[10253]), .Z(o[253]) );
  AND U8291 ( .A(p_input[2539]), .B(p_input[12539]), .Z(o[2539]) );
  AND U8292 ( .A(p_input[2538]), .B(p_input[12538]), .Z(o[2538]) );
  AND U8293 ( .A(p_input[2537]), .B(p_input[12537]), .Z(o[2537]) );
  AND U8294 ( .A(p_input[2536]), .B(p_input[12536]), .Z(o[2536]) );
  AND U8295 ( .A(p_input[2535]), .B(p_input[12535]), .Z(o[2535]) );
  AND U8296 ( .A(p_input[2534]), .B(p_input[12534]), .Z(o[2534]) );
  AND U8297 ( .A(p_input[2533]), .B(p_input[12533]), .Z(o[2533]) );
  AND U8298 ( .A(p_input[2532]), .B(p_input[12532]), .Z(o[2532]) );
  AND U8299 ( .A(p_input[2531]), .B(p_input[12531]), .Z(o[2531]) );
  AND U8300 ( .A(p_input[2530]), .B(p_input[12530]), .Z(o[2530]) );
  AND U8301 ( .A(p_input[252]), .B(p_input[10252]), .Z(o[252]) );
  AND U8302 ( .A(p_input[2529]), .B(p_input[12529]), .Z(o[2529]) );
  AND U8303 ( .A(p_input[2528]), .B(p_input[12528]), .Z(o[2528]) );
  AND U8304 ( .A(p_input[2527]), .B(p_input[12527]), .Z(o[2527]) );
  AND U8305 ( .A(p_input[2526]), .B(p_input[12526]), .Z(o[2526]) );
  AND U8306 ( .A(p_input[2525]), .B(p_input[12525]), .Z(o[2525]) );
  AND U8307 ( .A(p_input[2524]), .B(p_input[12524]), .Z(o[2524]) );
  AND U8308 ( .A(p_input[2523]), .B(p_input[12523]), .Z(o[2523]) );
  AND U8309 ( .A(p_input[2522]), .B(p_input[12522]), .Z(o[2522]) );
  AND U8310 ( .A(p_input[2521]), .B(p_input[12521]), .Z(o[2521]) );
  AND U8311 ( .A(p_input[2520]), .B(p_input[12520]), .Z(o[2520]) );
  AND U8312 ( .A(p_input[251]), .B(p_input[10251]), .Z(o[251]) );
  AND U8313 ( .A(p_input[2519]), .B(p_input[12519]), .Z(o[2519]) );
  AND U8314 ( .A(p_input[2518]), .B(p_input[12518]), .Z(o[2518]) );
  AND U8315 ( .A(p_input[2517]), .B(p_input[12517]), .Z(o[2517]) );
  AND U8316 ( .A(p_input[2516]), .B(p_input[12516]), .Z(o[2516]) );
  AND U8317 ( .A(p_input[2515]), .B(p_input[12515]), .Z(o[2515]) );
  AND U8318 ( .A(p_input[2514]), .B(p_input[12514]), .Z(o[2514]) );
  AND U8319 ( .A(p_input[2513]), .B(p_input[12513]), .Z(o[2513]) );
  AND U8320 ( .A(p_input[2512]), .B(p_input[12512]), .Z(o[2512]) );
  AND U8321 ( .A(p_input[2511]), .B(p_input[12511]), .Z(o[2511]) );
  AND U8322 ( .A(p_input[2510]), .B(p_input[12510]), .Z(o[2510]) );
  AND U8323 ( .A(p_input[250]), .B(p_input[10250]), .Z(o[250]) );
  AND U8324 ( .A(p_input[2509]), .B(p_input[12509]), .Z(o[2509]) );
  AND U8325 ( .A(p_input[2508]), .B(p_input[12508]), .Z(o[2508]) );
  AND U8326 ( .A(p_input[2507]), .B(p_input[12507]), .Z(o[2507]) );
  AND U8327 ( .A(p_input[2506]), .B(p_input[12506]), .Z(o[2506]) );
  AND U8328 ( .A(p_input[2505]), .B(p_input[12505]), .Z(o[2505]) );
  AND U8329 ( .A(p_input[2504]), .B(p_input[12504]), .Z(o[2504]) );
  AND U8330 ( .A(p_input[2503]), .B(p_input[12503]), .Z(o[2503]) );
  AND U8331 ( .A(p_input[2502]), .B(p_input[12502]), .Z(o[2502]) );
  AND U8332 ( .A(p_input[2501]), .B(p_input[12501]), .Z(o[2501]) );
  AND U8333 ( .A(p_input[2500]), .B(p_input[12500]), .Z(o[2500]) );
  AND U8334 ( .A(p_input[24]), .B(p_input[10024]), .Z(o[24]) );
  AND U8335 ( .A(p_input[249]), .B(p_input[10249]), .Z(o[249]) );
  AND U8336 ( .A(p_input[2499]), .B(p_input[12499]), .Z(o[2499]) );
  AND U8337 ( .A(p_input[2498]), .B(p_input[12498]), .Z(o[2498]) );
  AND U8338 ( .A(p_input[2497]), .B(p_input[12497]), .Z(o[2497]) );
  AND U8339 ( .A(p_input[2496]), .B(p_input[12496]), .Z(o[2496]) );
  AND U8340 ( .A(p_input[2495]), .B(p_input[12495]), .Z(o[2495]) );
  AND U8341 ( .A(p_input[2494]), .B(p_input[12494]), .Z(o[2494]) );
  AND U8342 ( .A(p_input[2493]), .B(p_input[12493]), .Z(o[2493]) );
  AND U8343 ( .A(p_input[2492]), .B(p_input[12492]), .Z(o[2492]) );
  AND U8344 ( .A(p_input[2491]), .B(p_input[12491]), .Z(o[2491]) );
  AND U8345 ( .A(p_input[2490]), .B(p_input[12490]), .Z(o[2490]) );
  AND U8346 ( .A(p_input[248]), .B(p_input[10248]), .Z(o[248]) );
  AND U8347 ( .A(p_input[2489]), .B(p_input[12489]), .Z(o[2489]) );
  AND U8348 ( .A(p_input[2488]), .B(p_input[12488]), .Z(o[2488]) );
  AND U8349 ( .A(p_input[2487]), .B(p_input[12487]), .Z(o[2487]) );
  AND U8350 ( .A(p_input[2486]), .B(p_input[12486]), .Z(o[2486]) );
  AND U8351 ( .A(p_input[2485]), .B(p_input[12485]), .Z(o[2485]) );
  AND U8352 ( .A(p_input[2484]), .B(p_input[12484]), .Z(o[2484]) );
  AND U8353 ( .A(p_input[2483]), .B(p_input[12483]), .Z(o[2483]) );
  AND U8354 ( .A(p_input[2482]), .B(p_input[12482]), .Z(o[2482]) );
  AND U8355 ( .A(p_input[2481]), .B(p_input[12481]), .Z(o[2481]) );
  AND U8356 ( .A(p_input[2480]), .B(p_input[12480]), .Z(o[2480]) );
  AND U8357 ( .A(p_input[247]), .B(p_input[10247]), .Z(o[247]) );
  AND U8358 ( .A(p_input[2479]), .B(p_input[12479]), .Z(o[2479]) );
  AND U8359 ( .A(p_input[2478]), .B(p_input[12478]), .Z(o[2478]) );
  AND U8360 ( .A(p_input[2477]), .B(p_input[12477]), .Z(o[2477]) );
  AND U8361 ( .A(p_input[2476]), .B(p_input[12476]), .Z(o[2476]) );
  AND U8362 ( .A(p_input[2475]), .B(p_input[12475]), .Z(o[2475]) );
  AND U8363 ( .A(p_input[2474]), .B(p_input[12474]), .Z(o[2474]) );
  AND U8364 ( .A(p_input[2473]), .B(p_input[12473]), .Z(o[2473]) );
  AND U8365 ( .A(p_input[2472]), .B(p_input[12472]), .Z(o[2472]) );
  AND U8366 ( .A(p_input[2471]), .B(p_input[12471]), .Z(o[2471]) );
  AND U8367 ( .A(p_input[2470]), .B(p_input[12470]), .Z(o[2470]) );
  AND U8368 ( .A(p_input[246]), .B(p_input[10246]), .Z(o[246]) );
  AND U8369 ( .A(p_input[2469]), .B(p_input[12469]), .Z(o[2469]) );
  AND U8370 ( .A(p_input[2468]), .B(p_input[12468]), .Z(o[2468]) );
  AND U8371 ( .A(p_input[2467]), .B(p_input[12467]), .Z(o[2467]) );
  AND U8372 ( .A(p_input[2466]), .B(p_input[12466]), .Z(o[2466]) );
  AND U8373 ( .A(p_input[2465]), .B(p_input[12465]), .Z(o[2465]) );
  AND U8374 ( .A(p_input[2464]), .B(p_input[12464]), .Z(o[2464]) );
  AND U8375 ( .A(p_input[2463]), .B(p_input[12463]), .Z(o[2463]) );
  AND U8376 ( .A(p_input[2462]), .B(p_input[12462]), .Z(o[2462]) );
  AND U8377 ( .A(p_input[2461]), .B(p_input[12461]), .Z(o[2461]) );
  AND U8378 ( .A(p_input[2460]), .B(p_input[12460]), .Z(o[2460]) );
  AND U8379 ( .A(p_input[245]), .B(p_input[10245]), .Z(o[245]) );
  AND U8380 ( .A(p_input[2459]), .B(p_input[12459]), .Z(o[2459]) );
  AND U8381 ( .A(p_input[2458]), .B(p_input[12458]), .Z(o[2458]) );
  AND U8382 ( .A(p_input[2457]), .B(p_input[12457]), .Z(o[2457]) );
  AND U8383 ( .A(p_input[2456]), .B(p_input[12456]), .Z(o[2456]) );
  AND U8384 ( .A(p_input[2455]), .B(p_input[12455]), .Z(o[2455]) );
  AND U8385 ( .A(p_input[2454]), .B(p_input[12454]), .Z(o[2454]) );
  AND U8386 ( .A(p_input[2453]), .B(p_input[12453]), .Z(o[2453]) );
  AND U8387 ( .A(p_input[2452]), .B(p_input[12452]), .Z(o[2452]) );
  AND U8388 ( .A(p_input[2451]), .B(p_input[12451]), .Z(o[2451]) );
  AND U8389 ( .A(p_input[2450]), .B(p_input[12450]), .Z(o[2450]) );
  AND U8390 ( .A(p_input[244]), .B(p_input[10244]), .Z(o[244]) );
  AND U8391 ( .A(p_input[2449]), .B(p_input[12449]), .Z(o[2449]) );
  AND U8392 ( .A(p_input[2448]), .B(p_input[12448]), .Z(o[2448]) );
  AND U8393 ( .A(p_input[2447]), .B(p_input[12447]), .Z(o[2447]) );
  AND U8394 ( .A(p_input[2446]), .B(p_input[12446]), .Z(o[2446]) );
  AND U8395 ( .A(p_input[2445]), .B(p_input[12445]), .Z(o[2445]) );
  AND U8396 ( .A(p_input[2444]), .B(p_input[12444]), .Z(o[2444]) );
  AND U8397 ( .A(p_input[2443]), .B(p_input[12443]), .Z(o[2443]) );
  AND U8398 ( .A(p_input[2442]), .B(p_input[12442]), .Z(o[2442]) );
  AND U8399 ( .A(p_input[2441]), .B(p_input[12441]), .Z(o[2441]) );
  AND U8400 ( .A(p_input[2440]), .B(p_input[12440]), .Z(o[2440]) );
  AND U8401 ( .A(p_input[243]), .B(p_input[10243]), .Z(o[243]) );
  AND U8402 ( .A(p_input[2439]), .B(p_input[12439]), .Z(o[2439]) );
  AND U8403 ( .A(p_input[2438]), .B(p_input[12438]), .Z(o[2438]) );
  AND U8404 ( .A(p_input[2437]), .B(p_input[12437]), .Z(o[2437]) );
  AND U8405 ( .A(p_input[2436]), .B(p_input[12436]), .Z(o[2436]) );
  AND U8406 ( .A(p_input[2435]), .B(p_input[12435]), .Z(o[2435]) );
  AND U8407 ( .A(p_input[2434]), .B(p_input[12434]), .Z(o[2434]) );
  AND U8408 ( .A(p_input[2433]), .B(p_input[12433]), .Z(o[2433]) );
  AND U8409 ( .A(p_input[2432]), .B(p_input[12432]), .Z(o[2432]) );
  AND U8410 ( .A(p_input[2431]), .B(p_input[12431]), .Z(o[2431]) );
  AND U8411 ( .A(p_input[2430]), .B(p_input[12430]), .Z(o[2430]) );
  AND U8412 ( .A(p_input[242]), .B(p_input[10242]), .Z(o[242]) );
  AND U8413 ( .A(p_input[2429]), .B(p_input[12429]), .Z(o[2429]) );
  AND U8414 ( .A(p_input[2428]), .B(p_input[12428]), .Z(o[2428]) );
  AND U8415 ( .A(p_input[2427]), .B(p_input[12427]), .Z(o[2427]) );
  AND U8416 ( .A(p_input[2426]), .B(p_input[12426]), .Z(o[2426]) );
  AND U8417 ( .A(p_input[2425]), .B(p_input[12425]), .Z(o[2425]) );
  AND U8418 ( .A(p_input[2424]), .B(p_input[12424]), .Z(o[2424]) );
  AND U8419 ( .A(p_input[2423]), .B(p_input[12423]), .Z(o[2423]) );
  AND U8420 ( .A(p_input[2422]), .B(p_input[12422]), .Z(o[2422]) );
  AND U8421 ( .A(p_input[2421]), .B(p_input[12421]), .Z(o[2421]) );
  AND U8422 ( .A(p_input[2420]), .B(p_input[12420]), .Z(o[2420]) );
  AND U8423 ( .A(p_input[241]), .B(p_input[10241]), .Z(o[241]) );
  AND U8424 ( .A(p_input[2419]), .B(p_input[12419]), .Z(o[2419]) );
  AND U8425 ( .A(p_input[2418]), .B(p_input[12418]), .Z(o[2418]) );
  AND U8426 ( .A(p_input[2417]), .B(p_input[12417]), .Z(o[2417]) );
  AND U8427 ( .A(p_input[2416]), .B(p_input[12416]), .Z(o[2416]) );
  AND U8428 ( .A(p_input[2415]), .B(p_input[12415]), .Z(o[2415]) );
  AND U8429 ( .A(p_input[2414]), .B(p_input[12414]), .Z(o[2414]) );
  AND U8430 ( .A(p_input[2413]), .B(p_input[12413]), .Z(o[2413]) );
  AND U8431 ( .A(p_input[2412]), .B(p_input[12412]), .Z(o[2412]) );
  AND U8432 ( .A(p_input[2411]), .B(p_input[12411]), .Z(o[2411]) );
  AND U8433 ( .A(p_input[2410]), .B(p_input[12410]), .Z(o[2410]) );
  AND U8434 ( .A(p_input[240]), .B(p_input[10240]), .Z(o[240]) );
  AND U8435 ( .A(p_input[2409]), .B(p_input[12409]), .Z(o[2409]) );
  AND U8436 ( .A(p_input[2408]), .B(p_input[12408]), .Z(o[2408]) );
  AND U8437 ( .A(p_input[2407]), .B(p_input[12407]), .Z(o[2407]) );
  AND U8438 ( .A(p_input[2406]), .B(p_input[12406]), .Z(o[2406]) );
  AND U8439 ( .A(p_input[2405]), .B(p_input[12405]), .Z(o[2405]) );
  AND U8440 ( .A(p_input[2404]), .B(p_input[12404]), .Z(o[2404]) );
  AND U8441 ( .A(p_input[2403]), .B(p_input[12403]), .Z(o[2403]) );
  AND U8442 ( .A(p_input[2402]), .B(p_input[12402]), .Z(o[2402]) );
  AND U8443 ( .A(p_input[2401]), .B(p_input[12401]), .Z(o[2401]) );
  AND U8444 ( .A(p_input[2400]), .B(p_input[12400]), .Z(o[2400]) );
  AND U8445 ( .A(p_input[23]), .B(p_input[10023]), .Z(o[23]) );
  AND U8446 ( .A(p_input[239]), .B(p_input[10239]), .Z(o[239]) );
  AND U8447 ( .A(p_input[2399]), .B(p_input[12399]), .Z(o[2399]) );
  AND U8448 ( .A(p_input[2398]), .B(p_input[12398]), .Z(o[2398]) );
  AND U8449 ( .A(p_input[2397]), .B(p_input[12397]), .Z(o[2397]) );
  AND U8450 ( .A(p_input[2396]), .B(p_input[12396]), .Z(o[2396]) );
  AND U8451 ( .A(p_input[2395]), .B(p_input[12395]), .Z(o[2395]) );
  AND U8452 ( .A(p_input[2394]), .B(p_input[12394]), .Z(o[2394]) );
  AND U8453 ( .A(p_input[2393]), .B(p_input[12393]), .Z(o[2393]) );
  AND U8454 ( .A(p_input[2392]), .B(p_input[12392]), .Z(o[2392]) );
  AND U8455 ( .A(p_input[2391]), .B(p_input[12391]), .Z(o[2391]) );
  AND U8456 ( .A(p_input[2390]), .B(p_input[12390]), .Z(o[2390]) );
  AND U8457 ( .A(p_input[238]), .B(p_input[10238]), .Z(o[238]) );
  AND U8458 ( .A(p_input[2389]), .B(p_input[12389]), .Z(o[2389]) );
  AND U8459 ( .A(p_input[2388]), .B(p_input[12388]), .Z(o[2388]) );
  AND U8460 ( .A(p_input[2387]), .B(p_input[12387]), .Z(o[2387]) );
  AND U8461 ( .A(p_input[2386]), .B(p_input[12386]), .Z(o[2386]) );
  AND U8462 ( .A(p_input[2385]), .B(p_input[12385]), .Z(o[2385]) );
  AND U8463 ( .A(p_input[2384]), .B(p_input[12384]), .Z(o[2384]) );
  AND U8464 ( .A(p_input[2383]), .B(p_input[12383]), .Z(o[2383]) );
  AND U8465 ( .A(p_input[2382]), .B(p_input[12382]), .Z(o[2382]) );
  AND U8466 ( .A(p_input[2381]), .B(p_input[12381]), .Z(o[2381]) );
  AND U8467 ( .A(p_input[2380]), .B(p_input[12380]), .Z(o[2380]) );
  AND U8468 ( .A(p_input[237]), .B(p_input[10237]), .Z(o[237]) );
  AND U8469 ( .A(p_input[2379]), .B(p_input[12379]), .Z(o[2379]) );
  AND U8470 ( .A(p_input[2378]), .B(p_input[12378]), .Z(o[2378]) );
  AND U8471 ( .A(p_input[2377]), .B(p_input[12377]), .Z(o[2377]) );
  AND U8472 ( .A(p_input[2376]), .B(p_input[12376]), .Z(o[2376]) );
  AND U8473 ( .A(p_input[2375]), .B(p_input[12375]), .Z(o[2375]) );
  AND U8474 ( .A(p_input[2374]), .B(p_input[12374]), .Z(o[2374]) );
  AND U8475 ( .A(p_input[2373]), .B(p_input[12373]), .Z(o[2373]) );
  AND U8476 ( .A(p_input[2372]), .B(p_input[12372]), .Z(o[2372]) );
  AND U8477 ( .A(p_input[2371]), .B(p_input[12371]), .Z(o[2371]) );
  AND U8478 ( .A(p_input[2370]), .B(p_input[12370]), .Z(o[2370]) );
  AND U8479 ( .A(p_input[236]), .B(p_input[10236]), .Z(o[236]) );
  AND U8480 ( .A(p_input[2369]), .B(p_input[12369]), .Z(o[2369]) );
  AND U8481 ( .A(p_input[2368]), .B(p_input[12368]), .Z(o[2368]) );
  AND U8482 ( .A(p_input[2367]), .B(p_input[12367]), .Z(o[2367]) );
  AND U8483 ( .A(p_input[2366]), .B(p_input[12366]), .Z(o[2366]) );
  AND U8484 ( .A(p_input[2365]), .B(p_input[12365]), .Z(o[2365]) );
  AND U8485 ( .A(p_input[2364]), .B(p_input[12364]), .Z(o[2364]) );
  AND U8486 ( .A(p_input[2363]), .B(p_input[12363]), .Z(o[2363]) );
  AND U8487 ( .A(p_input[2362]), .B(p_input[12362]), .Z(o[2362]) );
  AND U8488 ( .A(p_input[2361]), .B(p_input[12361]), .Z(o[2361]) );
  AND U8489 ( .A(p_input[2360]), .B(p_input[12360]), .Z(o[2360]) );
  AND U8490 ( .A(p_input[235]), .B(p_input[10235]), .Z(o[235]) );
  AND U8491 ( .A(p_input[2359]), .B(p_input[12359]), .Z(o[2359]) );
  AND U8492 ( .A(p_input[2358]), .B(p_input[12358]), .Z(o[2358]) );
  AND U8493 ( .A(p_input[2357]), .B(p_input[12357]), .Z(o[2357]) );
  AND U8494 ( .A(p_input[2356]), .B(p_input[12356]), .Z(o[2356]) );
  AND U8495 ( .A(p_input[2355]), .B(p_input[12355]), .Z(o[2355]) );
  AND U8496 ( .A(p_input[2354]), .B(p_input[12354]), .Z(o[2354]) );
  AND U8497 ( .A(p_input[2353]), .B(p_input[12353]), .Z(o[2353]) );
  AND U8498 ( .A(p_input[2352]), .B(p_input[12352]), .Z(o[2352]) );
  AND U8499 ( .A(p_input[2351]), .B(p_input[12351]), .Z(o[2351]) );
  AND U8500 ( .A(p_input[2350]), .B(p_input[12350]), .Z(o[2350]) );
  AND U8501 ( .A(p_input[234]), .B(p_input[10234]), .Z(o[234]) );
  AND U8502 ( .A(p_input[2349]), .B(p_input[12349]), .Z(o[2349]) );
  AND U8503 ( .A(p_input[2348]), .B(p_input[12348]), .Z(o[2348]) );
  AND U8504 ( .A(p_input[2347]), .B(p_input[12347]), .Z(o[2347]) );
  AND U8505 ( .A(p_input[2346]), .B(p_input[12346]), .Z(o[2346]) );
  AND U8506 ( .A(p_input[2345]), .B(p_input[12345]), .Z(o[2345]) );
  AND U8507 ( .A(p_input[2344]), .B(p_input[12344]), .Z(o[2344]) );
  AND U8508 ( .A(p_input[2343]), .B(p_input[12343]), .Z(o[2343]) );
  AND U8509 ( .A(p_input[2342]), .B(p_input[12342]), .Z(o[2342]) );
  AND U8510 ( .A(p_input[2341]), .B(p_input[12341]), .Z(o[2341]) );
  AND U8511 ( .A(p_input[2340]), .B(p_input[12340]), .Z(o[2340]) );
  AND U8512 ( .A(p_input[233]), .B(p_input[10233]), .Z(o[233]) );
  AND U8513 ( .A(p_input[2339]), .B(p_input[12339]), .Z(o[2339]) );
  AND U8514 ( .A(p_input[2338]), .B(p_input[12338]), .Z(o[2338]) );
  AND U8515 ( .A(p_input[2337]), .B(p_input[12337]), .Z(o[2337]) );
  AND U8516 ( .A(p_input[2336]), .B(p_input[12336]), .Z(o[2336]) );
  AND U8517 ( .A(p_input[2335]), .B(p_input[12335]), .Z(o[2335]) );
  AND U8518 ( .A(p_input[2334]), .B(p_input[12334]), .Z(o[2334]) );
  AND U8519 ( .A(p_input[2333]), .B(p_input[12333]), .Z(o[2333]) );
  AND U8520 ( .A(p_input[2332]), .B(p_input[12332]), .Z(o[2332]) );
  AND U8521 ( .A(p_input[2331]), .B(p_input[12331]), .Z(o[2331]) );
  AND U8522 ( .A(p_input[2330]), .B(p_input[12330]), .Z(o[2330]) );
  AND U8523 ( .A(p_input[232]), .B(p_input[10232]), .Z(o[232]) );
  AND U8524 ( .A(p_input[2329]), .B(p_input[12329]), .Z(o[2329]) );
  AND U8525 ( .A(p_input[2328]), .B(p_input[12328]), .Z(o[2328]) );
  AND U8526 ( .A(p_input[2327]), .B(p_input[12327]), .Z(o[2327]) );
  AND U8527 ( .A(p_input[2326]), .B(p_input[12326]), .Z(o[2326]) );
  AND U8528 ( .A(p_input[2325]), .B(p_input[12325]), .Z(o[2325]) );
  AND U8529 ( .A(p_input[2324]), .B(p_input[12324]), .Z(o[2324]) );
  AND U8530 ( .A(p_input[2323]), .B(p_input[12323]), .Z(o[2323]) );
  AND U8531 ( .A(p_input[2322]), .B(p_input[12322]), .Z(o[2322]) );
  AND U8532 ( .A(p_input[2321]), .B(p_input[12321]), .Z(o[2321]) );
  AND U8533 ( .A(p_input[2320]), .B(p_input[12320]), .Z(o[2320]) );
  AND U8534 ( .A(p_input[231]), .B(p_input[10231]), .Z(o[231]) );
  AND U8535 ( .A(p_input[2319]), .B(p_input[12319]), .Z(o[2319]) );
  AND U8536 ( .A(p_input[2318]), .B(p_input[12318]), .Z(o[2318]) );
  AND U8537 ( .A(p_input[2317]), .B(p_input[12317]), .Z(o[2317]) );
  AND U8538 ( .A(p_input[2316]), .B(p_input[12316]), .Z(o[2316]) );
  AND U8539 ( .A(p_input[2315]), .B(p_input[12315]), .Z(o[2315]) );
  AND U8540 ( .A(p_input[2314]), .B(p_input[12314]), .Z(o[2314]) );
  AND U8541 ( .A(p_input[2313]), .B(p_input[12313]), .Z(o[2313]) );
  AND U8542 ( .A(p_input[2312]), .B(p_input[12312]), .Z(o[2312]) );
  AND U8543 ( .A(p_input[2311]), .B(p_input[12311]), .Z(o[2311]) );
  AND U8544 ( .A(p_input[2310]), .B(p_input[12310]), .Z(o[2310]) );
  AND U8545 ( .A(p_input[230]), .B(p_input[10230]), .Z(o[230]) );
  AND U8546 ( .A(p_input[2309]), .B(p_input[12309]), .Z(o[2309]) );
  AND U8547 ( .A(p_input[2308]), .B(p_input[12308]), .Z(o[2308]) );
  AND U8548 ( .A(p_input[2307]), .B(p_input[12307]), .Z(o[2307]) );
  AND U8549 ( .A(p_input[2306]), .B(p_input[12306]), .Z(o[2306]) );
  AND U8550 ( .A(p_input[2305]), .B(p_input[12305]), .Z(o[2305]) );
  AND U8551 ( .A(p_input[2304]), .B(p_input[12304]), .Z(o[2304]) );
  AND U8552 ( .A(p_input[2303]), .B(p_input[12303]), .Z(o[2303]) );
  AND U8553 ( .A(p_input[2302]), .B(p_input[12302]), .Z(o[2302]) );
  AND U8554 ( .A(p_input[2301]), .B(p_input[12301]), .Z(o[2301]) );
  AND U8555 ( .A(p_input[2300]), .B(p_input[12300]), .Z(o[2300]) );
  AND U8556 ( .A(p_input[22]), .B(p_input[10022]), .Z(o[22]) );
  AND U8557 ( .A(p_input[229]), .B(p_input[10229]), .Z(o[229]) );
  AND U8558 ( .A(p_input[2299]), .B(p_input[12299]), .Z(o[2299]) );
  AND U8559 ( .A(p_input[2298]), .B(p_input[12298]), .Z(o[2298]) );
  AND U8560 ( .A(p_input[2297]), .B(p_input[12297]), .Z(o[2297]) );
  AND U8561 ( .A(p_input[2296]), .B(p_input[12296]), .Z(o[2296]) );
  AND U8562 ( .A(p_input[2295]), .B(p_input[12295]), .Z(o[2295]) );
  AND U8563 ( .A(p_input[2294]), .B(p_input[12294]), .Z(o[2294]) );
  AND U8564 ( .A(p_input[2293]), .B(p_input[12293]), .Z(o[2293]) );
  AND U8565 ( .A(p_input[2292]), .B(p_input[12292]), .Z(o[2292]) );
  AND U8566 ( .A(p_input[2291]), .B(p_input[12291]), .Z(o[2291]) );
  AND U8567 ( .A(p_input[2290]), .B(p_input[12290]), .Z(o[2290]) );
  AND U8568 ( .A(p_input[228]), .B(p_input[10228]), .Z(o[228]) );
  AND U8569 ( .A(p_input[2289]), .B(p_input[12289]), .Z(o[2289]) );
  AND U8570 ( .A(p_input[2288]), .B(p_input[12288]), .Z(o[2288]) );
  AND U8571 ( .A(p_input[2287]), .B(p_input[12287]), .Z(o[2287]) );
  AND U8572 ( .A(p_input[2286]), .B(p_input[12286]), .Z(o[2286]) );
  AND U8573 ( .A(p_input[2285]), .B(p_input[12285]), .Z(o[2285]) );
  AND U8574 ( .A(p_input[2284]), .B(p_input[12284]), .Z(o[2284]) );
  AND U8575 ( .A(p_input[2283]), .B(p_input[12283]), .Z(o[2283]) );
  AND U8576 ( .A(p_input[2282]), .B(p_input[12282]), .Z(o[2282]) );
  AND U8577 ( .A(p_input[2281]), .B(p_input[12281]), .Z(o[2281]) );
  AND U8578 ( .A(p_input[2280]), .B(p_input[12280]), .Z(o[2280]) );
  AND U8579 ( .A(p_input[227]), .B(p_input[10227]), .Z(o[227]) );
  AND U8580 ( .A(p_input[2279]), .B(p_input[12279]), .Z(o[2279]) );
  AND U8581 ( .A(p_input[2278]), .B(p_input[12278]), .Z(o[2278]) );
  AND U8582 ( .A(p_input[2277]), .B(p_input[12277]), .Z(o[2277]) );
  AND U8583 ( .A(p_input[2276]), .B(p_input[12276]), .Z(o[2276]) );
  AND U8584 ( .A(p_input[2275]), .B(p_input[12275]), .Z(o[2275]) );
  AND U8585 ( .A(p_input[2274]), .B(p_input[12274]), .Z(o[2274]) );
  AND U8586 ( .A(p_input[2273]), .B(p_input[12273]), .Z(o[2273]) );
  AND U8587 ( .A(p_input[2272]), .B(p_input[12272]), .Z(o[2272]) );
  AND U8588 ( .A(p_input[2271]), .B(p_input[12271]), .Z(o[2271]) );
  AND U8589 ( .A(p_input[2270]), .B(p_input[12270]), .Z(o[2270]) );
  AND U8590 ( .A(p_input[226]), .B(p_input[10226]), .Z(o[226]) );
  AND U8591 ( .A(p_input[2269]), .B(p_input[12269]), .Z(o[2269]) );
  AND U8592 ( .A(p_input[2268]), .B(p_input[12268]), .Z(o[2268]) );
  AND U8593 ( .A(p_input[2267]), .B(p_input[12267]), .Z(o[2267]) );
  AND U8594 ( .A(p_input[2266]), .B(p_input[12266]), .Z(o[2266]) );
  AND U8595 ( .A(p_input[2265]), .B(p_input[12265]), .Z(o[2265]) );
  AND U8596 ( .A(p_input[2264]), .B(p_input[12264]), .Z(o[2264]) );
  AND U8597 ( .A(p_input[2263]), .B(p_input[12263]), .Z(o[2263]) );
  AND U8598 ( .A(p_input[2262]), .B(p_input[12262]), .Z(o[2262]) );
  AND U8599 ( .A(p_input[2261]), .B(p_input[12261]), .Z(o[2261]) );
  AND U8600 ( .A(p_input[2260]), .B(p_input[12260]), .Z(o[2260]) );
  AND U8601 ( .A(p_input[225]), .B(p_input[10225]), .Z(o[225]) );
  AND U8602 ( .A(p_input[2259]), .B(p_input[12259]), .Z(o[2259]) );
  AND U8603 ( .A(p_input[2258]), .B(p_input[12258]), .Z(o[2258]) );
  AND U8604 ( .A(p_input[2257]), .B(p_input[12257]), .Z(o[2257]) );
  AND U8605 ( .A(p_input[2256]), .B(p_input[12256]), .Z(o[2256]) );
  AND U8606 ( .A(p_input[2255]), .B(p_input[12255]), .Z(o[2255]) );
  AND U8607 ( .A(p_input[2254]), .B(p_input[12254]), .Z(o[2254]) );
  AND U8608 ( .A(p_input[2253]), .B(p_input[12253]), .Z(o[2253]) );
  AND U8609 ( .A(p_input[2252]), .B(p_input[12252]), .Z(o[2252]) );
  AND U8610 ( .A(p_input[2251]), .B(p_input[12251]), .Z(o[2251]) );
  AND U8611 ( .A(p_input[2250]), .B(p_input[12250]), .Z(o[2250]) );
  AND U8612 ( .A(p_input[224]), .B(p_input[10224]), .Z(o[224]) );
  AND U8613 ( .A(p_input[2249]), .B(p_input[12249]), .Z(o[2249]) );
  AND U8614 ( .A(p_input[2248]), .B(p_input[12248]), .Z(o[2248]) );
  AND U8615 ( .A(p_input[2247]), .B(p_input[12247]), .Z(o[2247]) );
  AND U8616 ( .A(p_input[2246]), .B(p_input[12246]), .Z(o[2246]) );
  AND U8617 ( .A(p_input[2245]), .B(p_input[12245]), .Z(o[2245]) );
  AND U8618 ( .A(p_input[2244]), .B(p_input[12244]), .Z(o[2244]) );
  AND U8619 ( .A(p_input[2243]), .B(p_input[12243]), .Z(o[2243]) );
  AND U8620 ( .A(p_input[2242]), .B(p_input[12242]), .Z(o[2242]) );
  AND U8621 ( .A(p_input[2241]), .B(p_input[12241]), .Z(o[2241]) );
  AND U8622 ( .A(p_input[2240]), .B(p_input[12240]), .Z(o[2240]) );
  AND U8623 ( .A(p_input[223]), .B(p_input[10223]), .Z(o[223]) );
  AND U8624 ( .A(p_input[2239]), .B(p_input[12239]), .Z(o[2239]) );
  AND U8625 ( .A(p_input[2238]), .B(p_input[12238]), .Z(o[2238]) );
  AND U8626 ( .A(p_input[2237]), .B(p_input[12237]), .Z(o[2237]) );
  AND U8627 ( .A(p_input[2236]), .B(p_input[12236]), .Z(o[2236]) );
  AND U8628 ( .A(p_input[2235]), .B(p_input[12235]), .Z(o[2235]) );
  AND U8629 ( .A(p_input[2234]), .B(p_input[12234]), .Z(o[2234]) );
  AND U8630 ( .A(p_input[2233]), .B(p_input[12233]), .Z(o[2233]) );
  AND U8631 ( .A(p_input[2232]), .B(p_input[12232]), .Z(o[2232]) );
  AND U8632 ( .A(p_input[2231]), .B(p_input[12231]), .Z(o[2231]) );
  AND U8633 ( .A(p_input[2230]), .B(p_input[12230]), .Z(o[2230]) );
  AND U8634 ( .A(p_input[222]), .B(p_input[10222]), .Z(o[222]) );
  AND U8635 ( .A(p_input[2229]), .B(p_input[12229]), .Z(o[2229]) );
  AND U8636 ( .A(p_input[2228]), .B(p_input[12228]), .Z(o[2228]) );
  AND U8637 ( .A(p_input[2227]), .B(p_input[12227]), .Z(o[2227]) );
  AND U8638 ( .A(p_input[2226]), .B(p_input[12226]), .Z(o[2226]) );
  AND U8639 ( .A(p_input[2225]), .B(p_input[12225]), .Z(o[2225]) );
  AND U8640 ( .A(p_input[2224]), .B(p_input[12224]), .Z(o[2224]) );
  AND U8641 ( .A(p_input[2223]), .B(p_input[12223]), .Z(o[2223]) );
  AND U8642 ( .A(p_input[2222]), .B(p_input[12222]), .Z(o[2222]) );
  AND U8643 ( .A(p_input[2221]), .B(p_input[12221]), .Z(o[2221]) );
  AND U8644 ( .A(p_input[2220]), .B(p_input[12220]), .Z(o[2220]) );
  AND U8645 ( .A(p_input[221]), .B(p_input[10221]), .Z(o[221]) );
  AND U8646 ( .A(p_input[2219]), .B(p_input[12219]), .Z(o[2219]) );
  AND U8647 ( .A(p_input[2218]), .B(p_input[12218]), .Z(o[2218]) );
  AND U8648 ( .A(p_input[2217]), .B(p_input[12217]), .Z(o[2217]) );
  AND U8649 ( .A(p_input[2216]), .B(p_input[12216]), .Z(o[2216]) );
  AND U8650 ( .A(p_input[2215]), .B(p_input[12215]), .Z(o[2215]) );
  AND U8651 ( .A(p_input[2214]), .B(p_input[12214]), .Z(o[2214]) );
  AND U8652 ( .A(p_input[2213]), .B(p_input[12213]), .Z(o[2213]) );
  AND U8653 ( .A(p_input[2212]), .B(p_input[12212]), .Z(o[2212]) );
  AND U8654 ( .A(p_input[2211]), .B(p_input[12211]), .Z(o[2211]) );
  AND U8655 ( .A(p_input[2210]), .B(p_input[12210]), .Z(o[2210]) );
  AND U8656 ( .A(p_input[220]), .B(p_input[10220]), .Z(o[220]) );
  AND U8657 ( .A(p_input[2209]), .B(p_input[12209]), .Z(o[2209]) );
  AND U8658 ( .A(p_input[2208]), .B(p_input[12208]), .Z(o[2208]) );
  AND U8659 ( .A(p_input[2207]), .B(p_input[12207]), .Z(o[2207]) );
  AND U8660 ( .A(p_input[2206]), .B(p_input[12206]), .Z(o[2206]) );
  AND U8661 ( .A(p_input[2205]), .B(p_input[12205]), .Z(o[2205]) );
  AND U8662 ( .A(p_input[2204]), .B(p_input[12204]), .Z(o[2204]) );
  AND U8663 ( .A(p_input[2203]), .B(p_input[12203]), .Z(o[2203]) );
  AND U8664 ( .A(p_input[2202]), .B(p_input[12202]), .Z(o[2202]) );
  AND U8665 ( .A(p_input[2201]), .B(p_input[12201]), .Z(o[2201]) );
  AND U8666 ( .A(p_input[2200]), .B(p_input[12200]), .Z(o[2200]) );
  AND U8667 ( .A(p_input[21]), .B(p_input[10021]), .Z(o[21]) );
  AND U8668 ( .A(p_input[219]), .B(p_input[10219]), .Z(o[219]) );
  AND U8669 ( .A(p_input[2199]), .B(p_input[12199]), .Z(o[2199]) );
  AND U8670 ( .A(p_input[2198]), .B(p_input[12198]), .Z(o[2198]) );
  AND U8671 ( .A(p_input[2197]), .B(p_input[12197]), .Z(o[2197]) );
  AND U8672 ( .A(p_input[2196]), .B(p_input[12196]), .Z(o[2196]) );
  AND U8673 ( .A(p_input[2195]), .B(p_input[12195]), .Z(o[2195]) );
  AND U8674 ( .A(p_input[2194]), .B(p_input[12194]), .Z(o[2194]) );
  AND U8675 ( .A(p_input[2193]), .B(p_input[12193]), .Z(o[2193]) );
  AND U8676 ( .A(p_input[2192]), .B(p_input[12192]), .Z(o[2192]) );
  AND U8677 ( .A(p_input[2191]), .B(p_input[12191]), .Z(o[2191]) );
  AND U8678 ( .A(p_input[2190]), .B(p_input[12190]), .Z(o[2190]) );
  AND U8679 ( .A(p_input[218]), .B(p_input[10218]), .Z(o[218]) );
  AND U8680 ( .A(p_input[2189]), .B(p_input[12189]), .Z(o[2189]) );
  AND U8681 ( .A(p_input[2188]), .B(p_input[12188]), .Z(o[2188]) );
  AND U8682 ( .A(p_input[2187]), .B(p_input[12187]), .Z(o[2187]) );
  AND U8683 ( .A(p_input[2186]), .B(p_input[12186]), .Z(o[2186]) );
  AND U8684 ( .A(p_input[2185]), .B(p_input[12185]), .Z(o[2185]) );
  AND U8685 ( .A(p_input[2184]), .B(p_input[12184]), .Z(o[2184]) );
  AND U8686 ( .A(p_input[2183]), .B(p_input[12183]), .Z(o[2183]) );
  AND U8687 ( .A(p_input[2182]), .B(p_input[12182]), .Z(o[2182]) );
  AND U8688 ( .A(p_input[2181]), .B(p_input[12181]), .Z(o[2181]) );
  AND U8689 ( .A(p_input[2180]), .B(p_input[12180]), .Z(o[2180]) );
  AND U8690 ( .A(p_input[217]), .B(p_input[10217]), .Z(o[217]) );
  AND U8691 ( .A(p_input[2179]), .B(p_input[12179]), .Z(o[2179]) );
  AND U8692 ( .A(p_input[2178]), .B(p_input[12178]), .Z(o[2178]) );
  AND U8693 ( .A(p_input[2177]), .B(p_input[12177]), .Z(o[2177]) );
  AND U8694 ( .A(p_input[2176]), .B(p_input[12176]), .Z(o[2176]) );
  AND U8695 ( .A(p_input[2175]), .B(p_input[12175]), .Z(o[2175]) );
  AND U8696 ( .A(p_input[2174]), .B(p_input[12174]), .Z(o[2174]) );
  AND U8697 ( .A(p_input[2173]), .B(p_input[12173]), .Z(o[2173]) );
  AND U8698 ( .A(p_input[2172]), .B(p_input[12172]), .Z(o[2172]) );
  AND U8699 ( .A(p_input[2171]), .B(p_input[12171]), .Z(o[2171]) );
  AND U8700 ( .A(p_input[2170]), .B(p_input[12170]), .Z(o[2170]) );
  AND U8701 ( .A(p_input[216]), .B(p_input[10216]), .Z(o[216]) );
  AND U8702 ( .A(p_input[2169]), .B(p_input[12169]), .Z(o[2169]) );
  AND U8703 ( .A(p_input[2168]), .B(p_input[12168]), .Z(o[2168]) );
  AND U8704 ( .A(p_input[2167]), .B(p_input[12167]), .Z(o[2167]) );
  AND U8705 ( .A(p_input[2166]), .B(p_input[12166]), .Z(o[2166]) );
  AND U8706 ( .A(p_input[2165]), .B(p_input[12165]), .Z(o[2165]) );
  AND U8707 ( .A(p_input[2164]), .B(p_input[12164]), .Z(o[2164]) );
  AND U8708 ( .A(p_input[2163]), .B(p_input[12163]), .Z(o[2163]) );
  AND U8709 ( .A(p_input[2162]), .B(p_input[12162]), .Z(o[2162]) );
  AND U8710 ( .A(p_input[2161]), .B(p_input[12161]), .Z(o[2161]) );
  AND U8711 ( .A(p_input[2160]), .B(p_input[12160]), .Z(o[2160]) );
  AND U8712 ( .A(p_input[215]), .B(p_input[10215]), .Z(o[215]) );
  AND U8713 ( .A(p_input[2159]), .B(p_input[12159]), .Z(o[2159]) );
  AND U8714 ( .A(p_input[2158]), .B(p_input[12158]), .Z(o[2158]) );
  AND U8715 ( .A(p_input[2157]), .B(p_input[12157]), .Z(o[2157]) );
  AND U8716 ( .A(p_input[2156]), .B(p_input[12156]), .Z(o[2156]) );
  AND U8717 ( .A(p_input[2155]), .B(p_input[12155]), .Z(o[2155]) );
  AND U8718 ( .A(p_input[2154]), .B(p_input[12154]), .Z(o[2154]) );
  AND U8719 ( .A(p_input[2153]), .B(p_input[12153]), .Z(o[2153]) );
  AND U8720 ( .A(p_input[2152]), .B(p_input[12152]), .Z(o[2152]) );
  AND U8721 ( .A(p_input[2151]), .B(p_input[12151]), .Z(o[2151]) );
  AND U8722 ( .A(p_input[2150]), .B(p_input[12150]), .Z(o[2150]) );
  AND U8723 ( .A(p_input[214]), .B(p_input[10214]), .Z(o[214]) );
  AND U8724 ( .A(p_input[2149]), .B(p_input[12149]), .Z(o[2149]) );
  AND U8725 ( .A(p_input[2148]), .B(p_input[12148]), .Z(o[2148]) );
  AND U8726 ( .A(p_input[2147]), .B(p_input[12147]), .Z(o[2147]) );
  AND U8727 ( .A(p_input[2146]), .B(p_input[12146]), .Z(o[2146]) );
  AND U8728 ( .A(p_input[2145]), .B(p_input[12145]), .Z(o[2145]) );
  AND U8729 ( .A(p_input[2144]), .B(p_input[12144]), .Z(o[2144]) );
  AND U8730 ( .A(p_input[2143]), .B(p_input[12143]), .Z(o[2143]) );
  AND U8731 ( .A(p_input[2142]), .B(p_input[12142]), .Z(o[2142]) );
  AND U8732 ( .A(p_input[2141]), .B(p_input[12141]), .Z(o[2141]) );
  AND U8733 ( .A(p_input[2140]), .B(p_input[12140]), .Z(o[2140]) );
  AND U8734 ( .A(p_input[213]), .B(p_input[10213]), .Z(o[213]) );
  AND U8735 ( .A(p_input[2139]), .B(p_input[12139]), .Z(o[2139]) );
  AND U8736 ( .A(p_input[2138]), .B(p_input[12138]), .Z(o[2138]) );
  AND U8737 ( .A(p_input[2137]), .B(p_input[12137]), .Z(o[2137]) );
  AND U8738 ( .A(p_input[2136]), .B(p_input[12136]), .Z(o[2136]) );
  AND U8739 ( .A(p_input[2135]), .B(p_input[12135]), .Z(o[2135]) );
  AND U8740 ( .A(p_input[2134]), .B(p_input[12134]), .Z(o[2134]) );
  AND U8741 ( .A(p_input[2133]), .B(p_input[12133]), .Z(o[2133]) );
  AND U8742 ( .A(p_input[2132]), .B(p_input[12132]), .Z(o[2132]) );
  AND U8743 ( .A(p_input[2131]), .B(p_input[12131]), .Z(o[2131]) );
  AND U8744 ( .A(p_input[2130]), .B(p_input[12130]), .Z(o[2130]) );
  AND U8745 ( .A(p_input[212]), .B(p_input[10212]), .Z(o[212]) );
  AND U8746 ( .A(p_input[2129]), .B(p_input[12129]), .Z(o[2129]) );
  AND U8747 ( .A(p_input[2128]), .B(p_input[12128]), .Z(o[2128]) );
  AND U8748 ( .A(p_input[2127]), .B(p_input[12127]), .Z(o[2127]) );
  AND U8749 ( .A(p_input[2126]), .B(p_input[12126]), .Z(o[2126]) );
  AND U8750 ( .A(p_input[2125]), .B(p_input[12125]), .Z(o[2125]) );
  AND U8751 ( .A(p_input[2124]), .B(p_input[12124]), .Z(o[2124]) );
  AND U8752 ( .A(p_input[2123]), .B(p_input[12123]), .Z(o[2123]) );
  AND U8753 ( .A(p_input[2122]), .B(p_input[12122]), .Z(o[2122]) );
  AND U8754 ( .A(p_input[2121]), .B(p_input[12121]), .Z(o[2121]) );
  AND U8755 ( .A(p_input[2120]), .B(p_input[12120]), .Z(o[2120]) );
  AND U8756 ( .A(p_input[211]), .B(p_input[10211]), .Z(o[211]) );
  AND U8757 ( .A(p_input[2119]), .B(p_input[12119]), .Z(o[2119]) );
  AND U8758 ( .A(p_input[2118]), .B(p_input[12118]), .Z(o[2118]) );
  AND U8759 ( .A(p_input[2117]), .B(p_input[12117]), .Z(o[2117]) );
  AND U8760 ( .A(p_input[2116]), .B(p_input[12116]), .Z(o[2116]) );
  AND U8761 ( .A(p_input[2115]), .B(p_input[12115]), .Z(o[2115]) );
  AND U8762 ( .A(p_input[2114]), .B(p_input[12114]), .Z(o[2114]) );
  AND U8763 ( .A(p_input[2113]), .B(p_input[12113]), .Z(o[2113]) );
  AND U8764 ( .A(p_input[2112]), .B(p_input[12112]), .Z(o[2112]) );
  AND U8765 ( .A(p_input[2111]), .B(p_input[12111]), .Z(o[2111]) );
  AND U8766 ( .A(p_input[2110]), .B(p_input[12110]), .Z(o[2110]) );
  AND U8767 ( .A(p_input[210]), .B(p_input[10210]), .Z(o[210]) );
  AND U8768 ( .A(p_input[2109]), .B(p_input[12109]), .Z(o[2109]) );
  AND U8769 ( .A(p_input[2108]), .B(p_input[12108]), .Z(o[2108]) );
  AND U8770 ( .A(p_input[2107]), .B(p_input[12107]), .Z(o[2107]) );
  AND U8771 ( .A(p_input[2106]), .B(p_input[12106]), .Z(o[2106]) );
  AND U8772 ( .A(p_input[2105]), .B(p_input[12105]), .Z(o[2105]) );
  AND U8773 ( .A(p_input[2104]), .B(p_input[12104]), .Z(o[2104]) );
  AND U8774 ( .A(p_input[2103]), .B(p_input[12103]), .Z(o[2103]) );
  AND U8775 ( .A(p_input[2102]), .B(p_input[12102]), .Z(o[2102]) );
  AND U8776 ( .A(p_input[2101]), .B(p_input[12101]), .Z(o[2101]) );
  AND U8777 ( .A(p_input[2100]), .B(p_input[12100]), .Z(o[2100]) );
  AND U8778 ( .A(p_input[20]), .B(p_input[10020]), .Z(o[20]) );
  AND U8779 ( .A(p_input[209]), .B(p_input[10209]), .Z(o[209]) );
  AND U8780 ( .A(p_input[2099]), .B(p_input[12099]), .Z(o[2099]) );
  AND U8781 ( .A(p_input[2098]), .B(p_input[12098]), .Z(o[2098]) );
  AND U8782 ( .A(p_input[2097]), .B(p_input[12097]), .Z(o[2097]) );
  AND U8783 ( .A(p_input[2096]), .B(p_input[12096]), .Z(o[2096]) );
  AND U8784 ( .A(p_input[2095]), .B(p_input[12095]), .Z(o[2095]) );
  AND U8785 ( .A(p_input[2094]), .B(p_input[12094]), .Z(o[2094]) );
  AND U8786 ( .A(p_input[2093]), .B(p_input[12093]), .Z(o[2093]) );
  AND U8787 ( .A(p_input[2092]), .B(p_input[12092]), .Z(o[2092]) );
  AND U8788 ( .A(p_input[2091]), .B(p_input[12091]), .Z(o[2091]) );
  AND U8789 ( .A(p_input[2090]), .B(p_input[12090]), .Z(o[2090]) );
  AND U8790 ( .A(p_input[208]), .B(p_input[10208]), .Z(o[208]) );
  AND U8791 ( .A(p_input[2089]), .B(p_input[12089]), .Z(o[2089]) );
  AND U8792 ( .A(p_input[2088]), .B(p_input[12088]), .Z(o[2088]) );
  AND U8793 ( .A(p_input[2087]), .B(p_input[12087]), .Z(o[2087]) );
  AND U8794 ( .A(p_input[2086]), .B(p_input[12086]), .Z(o[2086]) );
  AND U8795 ( .A(p_input[2085]), .B(p_input[12085]), .Z(o[2085]) );
  AND U8796 ( .A(p_input[2084]), .B(p_input[12084]), .Z(o[2084]) );
  AND U8797 ( .A(p_input[2083]), .B(p_input[12083]), .Z(o[2083]) );
  AND U8798 ( .A(p_input[2082]), .B(p_input[12082]), .Z(o[2082]) );
  AND U8799 ( .A(p_input[2081]), .B(p_input[12081]), .Z(o[2081]) );
  AND U8800 ( .A(p_input[2080]), .B(p_input[12080]), .Z(o[2080]) );
  AND U8801 ( .A(p_input[207]), .B(p_input[10207]), .Z(o[207]) );
  AND U8802 ( .A(p_input[2079]), .B(p_input[12079]), .Z(o[2079]) );
  AND U8803 ( .A(p_input[2078]), .B(p_input[12078]), .Z(o[2078]) );
  AND U8804 ( .A(p_input[2077]), .B(p_input[12077]), .Z(o[2077]) );
  AND U8805 ( .A(p_input[2076]), .B(p_input[12076]), .Z(o[2076]) );
  AND U8806 ( .A(p_input[2075]), .B(p_input[12075]), .Z(o[2075]) );
  AND U8807 ( .A(p_input[2074]), .B(p_input[12074]), .Z(o[2074]) );
  AND U8808 ( .A(p_input[2073]), .B(p_input[12073]), .Z(o[2073]) );
  AND U8809 ( .A(p_input[2072]), .B(p_input[12072]), .Z(o[2072]) );
  AND U8810 ( .A(p_input[2071]), .B(p_input[12071]), .Z(o[2071]) );
  AND U8811 ( .A(p_input[2070]), .B(p_input[12070]), .Z(o[2070]) );
  AND U8812 ( .A(p_input[206]), .B(p_input[10206]), .Z(o[206]) );
  AND U8813 ( .A(p_input[2069]), .B(p_input[12069]), .Z(o[2069]) );
  AND U8814 ( .A(p_input[2068]), .B(p_input[12068]), .Z(o[2068]) );
  AND U8815 ( .A(p_input[2067]), .B(p_input[12067]), .Z(o[2067]) );
  AND U8816 ( .A(p_input[2066]), .B(p_input[12066]), .Z(o[2066]) );
  AND U8817 ( .A(p_input[2065]), .B(p_input[12065]), .Z(o[2065]) );
  AND U8818 ( .A(p_input[2064]), .B(p_input[12064]), .Z(o[2064]) );
  AND U8819 ( .A(p_input[2063]), .B(p_input[12063]), .Z(o[2063]) );
  AND U8820 ( .A(p_input[2062]), .B(p_input[12062]), .Z(o[2062]) );
  AND U8821 ( .A(p_input[2061]), .B(p_input[12061]), .Z(o[2061]) );
  AND U8822 ( .A(p_input[2060]), .B(p_input[12060]), .Z(o[2060]) );
  AND U8823 ( .A(p_input[205]), .B(p_input[10205]), .Z(o[205]) );
  AND U8824 ( .A(p_input[2059]), .B(p_input[12059]), .Z(o[2059]) );
  AND U8825 ( .A(p_input[2058]), .B(p_input[12058]), .Z(o[2058]) );
  AND U8826 ( .A(p_input[2057]), .B(p_input[12057]), .Z(o[2057]) );
  AND U8827 ( .A(p_input[2056]), .B(p_input[12056]), .Z(o[2056]) );
  AND U8828 ( .A(p_input[2055]), .B(p_input[12055]), .Z(o[2055]) );
  AND U8829 ( .A(p_input[2054]), .B(p_input[12054]), .Z(o[2054]) );
  AND U8830 ( .A(p_input[2053]), .B(p_input[12053]), .Z(o[2053]) );
  AND U8831 ( .A(p_input[2052]), .B(p_input[12052]), .Z(o[2052]) );
  AND U8832 ( .A(p_input[2051]), .B(p_input[12051]), .Z(o[2051]) );
  AND U8833 ( .A(p_input[2050]), .B(p_input[12050]), .Z(o[2050]) );
  AND U8834 ( .A(p_input[204]), .B(p_input[10204]), .Z(o[204]) );
  AND U8835 ( .A(p_input[2049]), .B(p_input[12049]), .Z(o[2049]) );
  AND U8836 ( .A(p_input[2048]), .B(p_input[12048]), .Z(o[2048]) );
  AND U8837 ( .A(p_input[2047]), .B(p_input[12047]), .Z(o[2047]) );
  AND U8838 ( .A(p_input[2046]), .B(p_input[12046]), .Z(o[2046]) );
  AND U8839 ( .A(p_input[2045]), .B(p_input[12045]), .Z(o[2045]) );
  AND U8840 ( .A(p_input[2044]), .B(p_input[12044]), .Z(o[2044]) );
  AND U8841 ( .A(p_input[2043]), .B(p_input[12043]), .Z(o[2043]) );
  AND U8842 ( .A(p_input[2042]), .B(p_input[12042]), .Z(o[2042]) );
  AND U8843 ( .A(p_input[2041]), .B(p_input[12041]), .Z(o[2041]) );
  AND U8844 ( .A(p_input[2040]), .B(p_input[12040]), .Z(o[2040]) );
  AND U8845 ( .A(p_input[203]), .B(p_input[10203]), .Z(o[203]) );
  AND U8846 ( .A(p_input[2039]), .B(p_input[12039]), .Z(o[2039]) );
  AND U8847 ( .A(p_input[2038]), .B(p_input[12038]), .Z(o[2038]) );
  AND U8848 ( .A(p_input[2037]), .B(p_input[12037]), .Z(o[2037]) );
  AND U8849 ( .A(p_input[2036]), .B(p_input[12036]), .Z(o[2036]) );
  AND U8850 ( .A(p_input[2035]), .B(p_input[12035]), .Z(o[2035]) );
  AND U8851 ( .A(p_input[2034]), .B(p_input[12034]), .Z(o[2034]) );
  AND U8852 ( .A(p_input[2033]), .B(p_input[12033]), .Z(o[2033]) );
  AND U8853 ( .A(p_input[2032]), .B(p_input[12032]), .Z(o[2032]) );
  AND U8854 ( .A(p_input[2031]), .B(p_input[12031]), .Z(o[2031]) );
  AND U8855 ( .A(p_input[2030]), .B(p_input[12030]), .Z(o[2030]) );
  AND U8856 ( .A(p_input[202]), .B(p_input[10202]), .Z(o[202]) );
  AND U8857 ( .A(p_input[2029]), .B(p_input[12029]), .Z(o[2029]) );
  AND U8858 ( .A(p_input[2028]), .B(p_input[12028]), .Z(o[2028]) );
  AND U8859 ( .A(p_input[2027]), .B(p_input[12027]), .Z(o[2027]) );
  AND U8860 ( .A(p_input[2026]), .B(p_input[12026]), .Z(o[2026]) );
  AND U8861 ( .A(p_input[2025]), .B(p_input[12025]), .Z(o[2025]) );
  AND U8862 ( .A(p_input[2024]), .B(p_input[12024]), .Z(o[2024]) );
  AND U8863 ( .A(p_input[2023]), .B(p_input[12023]), .Z(o[2023]) );
  AND U8864 ( .A(p_input[2022]), .B(p_input[12022]), .Z(o[2022]) );
  AND U8865 ( .A(p_input[2021]), .B(p_input[12021]), .Z(o[2021]) );
  AND U8866 ( .A(p_input[2020]), .B(p_input[12020]), .Z(o[2020]) );
  AND U8867 ( .A(p_input[201]), .B(p_input[10201]), .Z(o[201]) );
  AND U8868 ( .A(p_input[2019]), .B(p_input[12019]), .Z(o[2019]) );
  AND U8869 ( .A(p_input[2018]), .B(p_input[12018]), .Z(o[2018]) );
  AND U8870 ( .A(p_input[2017]), .B(p_input[12017]), .Z(o[2017]) );
  AND U8871 ( .A(p_input[2016]), .B(p_input[12016]), .Z(o[2016]) );
  AND U8872 ( .A(p_input[2015]), .B(p_input[12015]), .Z(o[2015]) );
  AND U8873 ( .A(p_input[2014]), .B(p_input[12014]), .Z(o[2014]) );
  AND U8874 ( .A(p_input[2013]), .B(p_input[12013]), .Z(o[2013]) );
  AND U8875 ( .A(p_input[2012]), .B(p_input[12012]), .Z(o[2012]) );
  AND U8876 ( .A(p_input[2011]), .B(p_input[12011]), .Z(o[2011]) );
  AND U8877 ( .A(p_input[2010]), .B(p_input[12010]), .Z(o[2010]) );
  AND U8878 ( .A(p_input[200]), .B(p_input[10200]), .Z(o[200]) );
  AND U8879 ( .A(p_input[2009]), .B(p_input[12009]), .Z(o[2009]) );
  AND U8880 ( .A(p_input[2008]), .B(p_input[12008]), .Z(o[2008]) );
  AND U8881 ( .A(p_input[2007]), .B(p_input[12007]), .Z(o[2007]) );
  AND U8882 ( .A(p_input[2006]), .B(p_input[12006]), .Z(o[2006]) );
  AND U8883 ( .A(p_input[2005]), .B(p_input[12005]), .Z(o[2005]) );
  AND U8884 ( .A(p_input[2004]), .B(p_input[12004]), .Z(o[2004]) );
  AND U8885 ( .A(p_input[2003]), .B(p_input[12003]), .Z(o[2003]) );
  AND U8886 ( .A(p_input[2002]), .B(p_input[12002]), .Z(o[2002]) );
  AND U8887 ( .A(p_input[2001]), .B(p_input[12001]), .Z(o[2001]) );
  AND U8888 ( .A(p_input[2000]), .B(p_input[12000]), .Z(o[2000]) );
  AND U8889 ( .A(p_input[1]), .B(p_input[10001]), .Z(o[1]) );
  AND U8890 ( .A(p_input[19]), .B(p_input[10019]), .Z(o[19]) );
  AND U8891 ( .A(p_input[199]), .B(p_input[10199]), .Z(o[199]) );
  AND U8892 ( .A(p_input[1999]), .B(p_input[11999]), .Z(o[1999]) );
  AND U8893 ( .A(p_input[1998]), .B(p_input[11998]), .Z(o[1998]) );
  AND U8894 ( .A(p_input[1997]), .B(p_input[11997]), .Z(o[1997]) );
  AND U8895 ( .A(p_input[1996]), .B(p_input[11996]), .Z(o[1996]) );
  AND U8896 ( .A(p_input[1995]), .B(p_input[11995]), .Z(o[1995]) );
  AND U8897 ( .A(p_input[1994]), .B(p_input[11994]), .Z(o[1994]) );
  AND U8898 ( .A(p_input[1993]), .B(p_input[11993]), .Z(o[1993]) );
  AND U8899 ( .A(p_input[1992]), .B(p_input[11992]), .Z(o[1992]) );
  AND U8900 ( .A(p_input[1991]), .B(p_input[11991]), .Z(o[1991]) );
  AND U8901 ( .A(p_input[1990]), .B(p_input[11990]), .Z(o[1990]) );
  AND U8902 ( .A(p_input[198]), .B(p_input[10198]), .Z(o[198]) );
  AND U8903 ( .A(p_input[1989]), .B(p_input[11989]), .Z(o[1989]) );
  AND U8904 ( .A(p_input[1988]), .B(p_input[11988]), .Z(o[1988]) );
  AND U8905 ( .A(p_input[1987]), .B(p_input[11987]), .Z(o[1987]) );
  AND U8906 ( .A(p_input[1986]), .B(p_input[11986]), .Z(o[1986]) );
  AND U8907 ( .A(p_input[1985]), .B(p_input[11985]), .Z(o[1985]) );
  AND U8908 ( .A(p_input[1984]), .B(p_input[11984]), .Z(o[1984]) );
  AND U8909 ( .A(p_input[1983]), .B(p_input[11983]), .Z(o[1983]) );
  AND U8910 ( .A(p_input[1982]), .B(p_input[11982]), .Z(o[1982]) );
  AND U8911 ( .A(p_input[1981]), .B(p_input[11981]), .Z(o[1981]) );
  AND U8912 ( .A(p_input[1980]), .B(p_input[11980]), .Z(o[1980]) );
  AND U8913 ( .A(p_input[197]), .B(p_input[10197]), .Z(o[197]) );
  AND U8914 ( .A(p_input[1979]), .B(p_input[11979]), .Z(o[1979]) );
  AND U8915 ( .A(p_input[1978]), .B(p_input[11978]), .Z(o[1978]) );
  AND U8916 ( .A(p_input[1977]), .B(p_input[11977]), .Z(o[1977]) );
  AND U8917 ( .A(p_input[1976]), .B(p_input[11976]), .Z(o[1976]) );
  AND U8918 ( .A(p_input[1975]), .B(p_input[11975]), .Z(o[1975]) );
  AND U8919 ( .A(p_input[1974]), .B(p_input[11974]), .Z(o[1974]) );
  AND U8920 ( .A(p_input[1973]), .B(p_input[11973]), .Z(o[1973]) );
  AND U8921 ( .A(p_input[1972]), .B(p_input[11972]), .Z(o[1972]) );
  AND U8922 ( .A(p_input[1971]), .B(p_input[11971]), .Z(o[1971]) );
  AND U8923 ( .A(p_input[1970]), .B(p_input[11970]), .Z(o[1970]) );
  AND U8924 ( .A(p_input[196]), .B(p_input[10196]), .Z(o[196]) );
  AND U8925 ( .A(p_input[1969]), .B(p_input[11969]), .Z(o[1969]) );
  AND U8926 ( .A(p_input[1968]), .B(p_input[11968]), .Z(o[1968]) );
  AND U8927 ( .A(p_input[1967]), .B(p_input[11967]), .Z(o[1967]) );
  AND U8928 ( .A(p_input[1966]), .B(p_input[11966]), .Z(o[1966]) );
  AND U8929 ( .A(p_input[1965]), .B(p_input[11965]), .Z(o[1965]) );
  AND U8930 ( .A(p_input[1964]), .B(p_input[11964]), .Z(o[1964]) );
  AND U8931 ( .A(p_input[1963]), .B(p_input[11963]), .Z(o[1963]) );
  AND U8932 ( .A(p_input[1962]), .B(p_input[11962]), .Z(o[1962]) );
  AND U8933 ( .A(p_input[1961]), .B(p_input[11961]), .Z(o[1961]) );
  AND U8934 ( .A(p_input[1960]), .B(p_input[11960]), .Z(o[1960]) );
  AND U8935 ( .A(p_input[195]), .B(p_input[10195]), .Z(o[195]) );
  AND U8936 ( .A(p_input[1959]), .B(p_input[11959]), .Z(o[1959]) );
  AND U8937 ( .A(p_input[1958]), .B(p_input[11958]), .Z(o[1958]) );
  AND U8938 ( .A(p_input[1957]), .B(p_input[11957]), .Z(o[1957]) );
  AND U8939 ( .A(p_input[1956]), .B(p_input[11956]), .Z(o[1956]) );
  AND U8940 ( .A(p_input[1955]), .B(p_input[11955]), .Z(o[1955]) );
  AND U8941 ( .A(p_input[1954]), .B(p_input[11954]), .Z(o[1954]) );
  AND U8942 ( .A(p_input[1953]), .B(p_input[11953]), .Z(o[1953]) );
  AND U8943 ( .A(p_input[1952]), .B(p_input[11952]), .Z(o[1952]) );
  AND U8944 ( .A(p_input[1951]), .B(p_input[11951]), .Z(o[1951]) );
  AND U8945 ( .A(p_input[1950]), .B(p_input[11950]), .Z(o[1950]) );
  AND U8946 ( .A(p_input[194]), .B(p_input[10194]), .Z(o[194]) );
  AND U8947 ( .A(p_input[1949]), .B(p_input[11949]), .Z(o[1949]) );
  AND U8948 ( .A(p_input[1948]), .B(p_input[11948]), .Z(o[1948]) );
  AND U8949 ( .A(p_input[1947]), .B(p_input[11947]), .Z(o[1947]) );
  AND U8950 ( .A(p_input[1946]), .B(p_input[11946]), .Z(o[1946]) );
  AND U8951 ( .A(p_input[1945]), .B(p_input[11945]), .Z(o[1945]) );
  AND U8952 ( .A(p_input[1944]), .B(p_input[11944]), .Z(o[1944]) );
  AND U8953 ( .A(p_input[1943]), .B(p_input[11943]), .Z(o[1943]) );
  AND U8954 ( .A(p_input[1942]), .B(p_input[11942]), .Z(o[1942]) );
  AND U8955 ( .A(p_input[1941]), .B(p_input[11941]), .Z(o[1941]) );
  AND U8956 ( .A(p_input[1940]), .B(p_input[11940]), .Z(o[1940]) );
  AND U8957 ( .A(p_input[193]), .B(p_input[10193]), .Z(o[193]) );
  AND U8958 ( .A(p_input[1939]), .B(p_input[11939]), .Z(o[1939]) );
  AND U8959 ( .A(p_input[1938]), .B(p_input[11938]), .Z(o[1938]) );
  AND U8960 ( .A(p_input[1937]), .B(p_input[11937]), .Z(o[1937]) );
  AND U8961 ( .A(p_input[1936]), .B(p_input[11936]), .Z(o[1936]) );
  AND U8962 ( .A(p_input[1935]), .B(p_input[11935]), .Z(o[1935]) );
  AND U8963 ( .A(p_input[1934]), .B(p_input[11934]), .Z(o[1934]) );
  AND U8964 ( .A(p_input[1933]), .B(p_input[11933]), .Z(o[1933]) );
  AND U8965 ( .A(p_input[1932]), .B(p_input[11932]), .Z(o[1932]) );
  AND U8966 ( .A(p_input[1931]), .B(p_input[11931]), .Z(o[1931]) );
  AND U8967 ( .A(p_input[1930]), .B(p_input[11930]), .Z(o[1930]) );
  AND U8968 ( .A(p_input[192]), .B(p_input[10192]), .Z(o[192]) );
  AND U8969 ( .A(p_input[1929]), .B(p_input[11929]), .Z(o[1929]) );
  AND U8970 ( .A(p_input[1928]), .B(p_input[11928]), .Z(o[1928]) );
  AND U8971 ( .A(p_input[1927]), .B(p_input[11927]), .Z(o[1927]) );
  AND U8972 ( .A(p_input[1926]), .B(p_input[11926]), .Z(o[1926]) );
  AND U8973 ( .A(p_input[1925]), .B(p_input[11925]), .Z(o[1925]) );
  AND U8974 ( .A(p_input[1924]), .B(p_input[11924]), .Z(o[1924]) );
  AND U8975 ( .A(p_input[1923]), .B(p_input[11923]), .Z(o[1923]) );
  AND U8976 ( .A(p_input[1922]), .B(p_input[11922]), .Z(o[1922]) );
  AND U8977 ( .A(p_input[1921]), .B(p_input[11921]), .Z(o[1921]) );
  AND U8978 ( .A(p_input[1920]), .B(p_input[11920]), .Z(o[1920]) );
  AND U8979 ( .A(p_input[191]), .B(p_input[10191]), .Z(o[191]) );
  AND U8980 ( .A(p_input[1919]), .B(p_input[11919]), .Z(o[1919]) );
  AND U8981 ( .A(p_input[1918]), .B(p_input[11918]), .Z(o[1918]) );
  AND U8982 ( .A(p_input[1917]), .B(p_input[11917]), .Z(o[1917]) );
  AND U8983 ( .A(p_input[1916]), .B(p_input[11916]), .Z(o[1916]) );
  AND U8984 ( .A(p_input[1915]), .B(p_input[11915]), .Z(o[1915]) );
  AND U8985 ( .A(p_input[1914]), .B(p_input[11914]), .Z(o[1914]) );
  AND U8986 ( .A(p_input[1913]), .B(p_input[11913]), .Z(o[1913]) );
  AND U8987 ( .A(p_input[1912]), .B(p_input[11912]), .Z(o[1912]) );
  AND U8988 ( .A(p_input[1911]), .B(p_input[11911]), .Z(o[1911]) );
  AND U8989 ( .A(p_input[1910]), .B(p_input[11910]), .Z(o[1910]) );
  AND U8990 ( .A(p_input[190]), .B(p_input[10190]), .Z(o[190]) );
  AND U8991 ( .A(p_input[1909]), .B(p_input[11909]), .Z(o[1909]) );
  AND U8992 ( .A(p_input[1908]), .B(p_input[11908]), .Z(o[1908]) );
  AND U8993 ( .A(p_input[1907]), .B(p_input[11907]), .Z(o[1907]) );
  AND U8994 ( .A(p_input[1906]), .B(p_input[11906]), .Z(o[1906]) );
  AND U8995 ( .A(p_input[1905]), .B(p_input[11905]), .Z(o[1905]) );
  AND U8996 ( .A(p_input[1904]), .B(p_input[11904]), .Z(o[1904]) );
  AND U8997 ( .A(p_input[1903]), .B(p_input[11903]), .Z(o[1903]) );
  AND U8998 ( .A(p_input[1902]), .B(p_input[11902]), .Z(o[1902]) );
  AND U8999 ( .A(p_input[1901]), .B(p_input[11901]), .Z(o[1901]) );
  AND U9000 ( .A(p_input[1900]), .B(p_input[11900]), .Z(o[1900]) );
  AND U9001 ( .A(p_input[18]), .B(p_input[10018]), .Z(o[18]) );
  AND U9002 ( .A(p_input[189]), .B(p_input[10189]), .Z(o[189]) );
  AND U9003 ( .A(p_input[1899]), .B(p_input[11899]), .Z(o[1899]) );
  AND U9004 ( .A(p_input[1898]), .B(p_input[11898]), .Z(o[1898]) );
  AND U9005 ( .A(p_input[1897]), .B(p_input[11897]), .Z(o[1897]) );
  AND U9006 ( .A(p_input[1896]), .B(p_input[11896]), .Z(o[1896]) );
  AND U9007 ( .A(p_input[1895]), .B(p_input[11895]), .Z(o[1895]) );
  AND U9008 ( .A(p_input[1894]), .B(p_input[11894]), .Z(o[1894]) );
  AND U9009 ( .A(p_input[1893]), .B(p_input[11893]), .Z(o[1893]) );
  AND U9010 ( .A(p_input[1892]), .B(p_input[11892]), .Z(o[1892]) );
  AND U9011 ( .A(p_input[1891]), .B(p_input[11891]), .Z(o[1891]) );
  AND U9012 ( .A(p_input[1890]), .B(p_input[11890]), .Z(o[1890]) );
  AND U9013 ( .A(p_input[188]), .B(p_input[10188]), .Z(o[188]) );
  AND U9014 ( .A(p_input[1889]), .B(p_input[11889]), .Z(o[1889]) );
  AND U9015 ( .A(p_input[1888]), .B(p_input[11888]), .Z(o[1888]) );
  AND U9016 ( .A(p_input[1887]), .B(p_input[11887]), .Z(o[1887]) );
  AND U9017 ( .A(p_input[1886]), .B(p_input[11886]), .Z(o[1886]) );
  AND U9018 ( .A(p_input[1885]), .B(p_input[11885]), .Z(o[1885]) );
  AND U9019 ( .A(p_input[1884]), .B(p_input[11884]), .Z(o[1884]) );
  AND U9020 ( .A(p_input[1883]), .B(p_input[11883]), .Z(o[1883]) );
  AND U9021 ( .A(p_input[1882]), .B(p_input[11882]), .Z(o[1882]) );
  AND U9022 ( .A(p_input[1881]), .B(p_input[11881]), .Z(o[1881]) );
  AND U9023 ( .A(p_input[1880]), .B(p_input[11880]), .Z(o[1880]) );
  AND U9024 ( .A(p_input[187]), .B(p_input[10187]), .Z(o[187]) );
  AND U9025 ( .A(p_input[1879]), .B(p_input[11879]), .Z(o[1879]) );
  AND U9026 ( .A(p_input[1878]), .B(p_input[11878]), .Z(o[1878]) );
  AND U9027 ( .A(p_input[1877]), .B(p_input[11877]), .Z(o[1877]) );
  AND U9028 ( .A(p_input[1876]), .B(p_input[11876]), .Z(o[1876]) );
  AND U9029 ( .A(p_input[1875]), .B(p_input[11875]), .Z(o[1875]) );
  AND U9030 ( .A(p_input[1874]), .B(p_input[11874]), .Z(o[1874]) );
  AND U9031 ( .A(p_input[1873]), .B(p_input[11873]), .Z(o[1873]) );
  AND U9032 ( .A(p_input[1872]), .B(p_input[11872]), .Z(o[1872]) );
  AND U9033 ( .A(p_input[1871]), .B(p_input[11871]), .Z(o[1871]) );
  AND U9034 ( .A(p_input[1870]), .B(p_input[11870]), .Z(o[1870]) );
  AND U9035 ( .A(p_input[186]), .B(p_input[10186]), .Z(o[186]) );
  AND U9036 ( .A(p_input[1869]), .B(p_input[11869]), .Z(o[1869]) );
  AND U9037 ( .A(p_input[1868]), .B(p_input[11868]), .Z(o[1868]) );
  AND U9038 ( .A(p_input[1867]), .B(p_input[11867]), .Z(o[1867]) );
  AND U9039 ( .A(p_input[1866]), .B(p_input[11866]), .Z(o[1866]) );
  AND U9040 ( .A(p_input[1865]), .B(p_input[11865]), .Z(o[1865]) );
  AND U9041 ( .A(p_input[1864]), .B(p_input[11864]), .Z(o[1864]) );
  AND U9042 ( .A(p_input[1863]), .B(p_input[11863]), .Z(o[1863]) );
  AND U9043 ( .A(p_input[1862]), .B(p_input[11862]), .Z(o[1862]) );
  AND U9044 ( .A(p_input[1861]), .B(p_input[11861]), .Z(o[1861]) );
  AND U9045 ( .A(p_input[1860]), .B(p_input[11860]), .Z(o[1860]) );
  AND U9046 ( .A(p_input[185]), .B(p_input[10185]), .Z(o[185]) );
  AND U9047 ( .A(p_input[1859]), .B(p_input[11859]), .Z(o[1859]) );
  AND U9048 ( .A(p_input[1858]), .B(p_input[11858]), .Z(o[1858]) );
  AND U9049 ( .A(p_input[1857]), .B(p_input[11857]), .Z(o[1857]) );
  AND U9050 ( .A(p_input[1856]), .B(p_input[11856]), .Z(o[1856]) );
  AND U9051 ( .A(p_input[1855]), .B(p_input[11855]), .Z(o[1855]) );
  AND U9052 ( .A(p_input[1854]), .B(p_input[11854]), .Z(o[1854]) );
  AND U9053 ( .A(p_input[1853]), .B(p_input[11853]), .Z(o[1853]) );
  AND U9054 ( .A(p_input[1852]), .B(p_input[11852]), .Z(o[1852]) );
  AND U9055 ( .A(p_input[1851]), .B(p_input[11851]), .Z(o[1851]) );
  AND U9056 ( .A(p_input[1850]), .B(p_input[11850]), .Z(o[1850]) );
  AND U9057 ( .A(p_input[184]), .B(p_input[10184]), .Z(o[184]) );
  AND U9058 ( .A(p_input[1849]), .B(p_input[11849]), .Z(o[1849]) );
  AND U9059 ( .A(p_input[1848]), .B(p_input[11848]), .Z(o[1848]) );
  AND U9060 ( .A(p_input[1847]), .B(p_input[11847]), .Z(o[1847]) );
  AND U9061 ( .A(p_input[1846]), .B(p_input[11846]), .Z(o[1846]) );
  AND U9062 ( .A(p_input[1845]), .B(p_input[11845]), .Z(o[1845]) );
  AND U9063 ( .A(p_input[1844]), .B(p_input[11844]), .Z(o[1844]) );
  AND U9064 ( .A(p_input[1843]), .B(p_input[11843]), .Z(o[1843]) );
  AND U9065 ( .A(p_input[1842]), .B(p_input[11842]), .Z(o[1842]) );
  AND U9066 ( .A(p_input[1841]), .B(p_input[11841]), .Z(o[1841]) );
  AND U9067 ( .A(p_input[1840]), .B(p_input[11840]), .Z(o[1840]) );
  AND U9068 ( .A(p_input[183]), .B(p_input[10183]), .Z(o[183]) );
  AND U9069 ( .A(p_input[1839]), .B(p_input[11839]), .Z(o[1839]) );
  AND U9070 ( .A(p_input[1838]), .B(p_input[11838]), .Z(o[1838]) );
  AND U9071 ( .A(p_input[1837]), .B(p_input[11837]), .Z(o[1837]) );
  AND U9072 ( .A(p_input[1836]), .B(p_input[11836]), .Z(o[1836]) );
  AND U9073 ( .A(p_input[1835]), .B(p_input[11835]), .Z(o[1835]) );
  AND U9074 ( .A(p_input[1834]), .B(p_input[11834]), .Z(o[1834]) );
  AND U9075 ( .A(p_input[1833]), .B(p_input[11833]), .Z(o[1833]) );
  AND U9076 ( .A(p_input[1832]), .B(p_input[11832]), .Z(o[1832]) );
  AND U9077 ( .A(p_input[1831]), .B(p_input[11831]), .Z(o[1831]) );
  AND U9078 ( .A(p_input[1830]), .B(p_input[11830]), .Z(o[1830]) );
  AND U9079 ( .A(p_input[182]), .B(p_input[10182]), .Z(o[182]) );
  AND U9080 ( .A(p_input[1829]), .B(p_input[11829]), .Z(o[1829]) );
  AND U9081 ( .A(p_input[1828]), .B(p_input[11828]), .Z(o[1828]) );
  AND U9082 ( .A(p_input[1827]), .B(p_input[11827]), .Z(o[1827]) );
  AND U9083 ( .A(p_input[1826]), .B(p_input[11826]), .Z(o[1826]) );
  AND U9084 ( .A(p_input[1825]), .B(p_input[11825]), .Z(o[1825]) );
  AND U9085 ( .A(p_input[1824]), .B(p_input[11824]), .Z(o[1824]) );
  AND U9086 ( .A(p_input[1823]), .B(p_input[11823]), .Z(o[1823]) );
  AND U9087 ( .A(p_input[1822]), .B(p_input[11822]), .Z(o[1822]) );
  AND U9088 ( .A(p_input[1821]), .B(p_input[11821]), .Z(o[1821]) );
  AND U9089 ( .A(p_input[1820]), .B(p_input[11820]), .Z(o[1820]) );
  AND U9090 ( .A(p_input[181]), .B(p_input[10181]), .Z(o[181]) );
  AND U9091 ( .A(p_input[1819]), .B(p_input[11819]), .Z(o[1819]) );
  AND U9092 ( .A(p_input[1818]), .B(p_input[11818]), .Z(o[1818]) );
  AND U9093 ( .A(p_input[1817]), .B(p_input[11817]), .Z(o[1817]) );
  AND U9094 ( .A(p_input[1816]), .B(p_input[11816]), .Z(o[1816]) );
  AND U9095 ( .A(p_input[1815]), .B(p_input[11815]), .Z(o[1815]) );
  AND U9096 ( .A(p_input[1814]), .B(p_input[11814]), .Z(o[1814]) );
  AND U9097 ( .A(p_input[1813]), .B(p_input[11813]), .Z(o[1813]) );
  AND U9098 ( .A(p_input[1812]), .B(p_input[11812]), .Z(o[1812]) );
  AND U9099 ( .A(p_input[1811]), .B(p_input[11811]), .Z(o[1811]) );
  AND U9100 ( .A(p_input[1810]), .B(p_input[11810]), .Z(o[1810]) );
  AND U9101 ( .A(p_input[180]), .B(p_input[10180]), .Z(o[180]) );
  AND U9102 ( .A(p_input[1809]), .B(p_input[11809]), .Z(o[1809]) );
  AND U9103 ( .A(p_input[1808]), .B(p_input[11808]), .Z(o[1808]) );
  AND U9104 ( .A(p_input[1807]), .B(p_input[11807]), .Z(o[1807]) );
  AND U9105 ( .A(p_input[1806]), .B(p_input[11806]), .Z(o[1806]) );
  AND U9106 ( .A(p_input[1805]), .B(p_input[11805]), .Z(o[1805]) );
  AND U9107 ( .A(p_input[1804]), .B(p_input[11804]), .Z(o[1804]) );
  AND U9108 ( .A(p_input[1803]), .B(p_input[11803]), .Z(o[1803]) );
  AND U9109 ( .A(p_input[1802]), .B(p_input[11802]), .Z(o[1802]) );
  AND U9110 ( .A(p_input[1801]), .B(p_input[11801]), .Z(o[1801]) );
  AND U9111 ( .A(p_input[1800]), .B(p_input[11800]), .Z(o[1800]) );
  AND U9112 ( .A(p_input[17]), .B(p_input[10017]), .Z(o[17]) );
  AND U9113 ( .A(p_input[179]), .B(p_input[10179]), .Z(o[179]) );
  AND U9114 ( .A(p_input[1799]), .B(p_input[11799]), .Z(o[1799]) );
  AND U9115 ( .A(p_input[1798]), .B(p_input[11798]), .Z(o[1798]) );
  AND U9116 ( .A(p_input[1797]), .B(p_input[11797]), .Z(o[1797]) );
  AND U9117 ( .A(p_input[1796]), .B(p_input[11796]), .Z(o[1796]) );
  AND U9118 ( .A(p_input[1795]), .B(p_input[11795]), .Z(o[1795]) );
  AND U9119 ( .A(p_input[1794]), .B(p_input[11794]), .Z(o[1794]) );
  AND U9120 ( .A(p_input[1793]), .B(p_input[11793]), .Z(o[1793]) );
  AND U9121 ( .A(p_input[1792]), .B(p_input[11792]), .Z(o[1792]) );
  AND U9122 ( .A(p_input[1791]), .B(p_input[11791]), .Z(o[1791]) );
  AND U9123 ( .A(p_input[1790]), .B(p_input[11790]), .Z(o[1790]) );
  AND U9124 ( .A(p_input[178]), .B(p_input[10178]), .Z(o[178]) );
  AND U9125 ( .A(p_input[1789]), .B(p_input[11789]), .Z(o[1789]) );
  AND U9126 ( .A(p_input[1788]), .B(p_input[11788]), .Z(o[1788]) );
  AND U9127 ( .A(p_input[1787]), .B(p_input[11787]), .Z(o[1787]) );
  AND U9128 ( .A(p_input[1786]), .B(p_input[11786]), .Z(o[1786]) );
  AND U9129 ( .A(p_input[1785]), .B(p_input[11785]), .Z(o[1785]) );
  AND U9130 ( .A(p_input[1784]), .B(p_input[11784]), .Z(o[1784]) );
  AND U9131 ( .A(p_input[1783]), .B(p_input[11783]), .Z(o[1783]) );
  AND U9132 ( .A(p_input[1782]), .B(p_input[11782]), .Z(o[1782]) );
  AND U9133 ( .A(p_input[1781]), .B(p_input[11781]), .Z(o[1781]) );
  AND U9134 ( .A(p_input[1780]), .B(p_input[11780]), .Z(o[1780]) );
  AND U9135 ( .A(p_input[177]), .B(p_input[10177]), .Z(o[177]) );
  AND U9136 ( .A(p_input[1779]), .B(p_input[11779]), .Z(o[1779]) );
  AND U9137 ( .A(p_input[1778]), .B(p_input[11778]), .Z(o[1778]) );
  AND U9138 ( .A(p_input[1777]), .B(p_input[11777]), .Z(o[1777]) );
  AND U9139 ( .A(p_input[1776]), .B(p_input[11776]), .Z(o[1776]) );
  AND U9140 ( .A(p_input[1775]), .B(p_input[11775]), .Z(o[1775]) );
  AND U9141 ( .A(p_input[1774]), .B(p_input[11774]), .Z(o[1774]) );
  AND U9142 ( .A(p_input[1773]), .B(p_input[11773]), .Z(o[1773]) );
  AND U9143 ( .A(p_input[1772]), .B(p_input[11772]), .Z(o[1772]) );
  AND U9144 ( .A(p_input[1771]), .B(p_input[11771]), .Z(o[1771]) );
  AND U9145 ( .A(p_input[1770]), .B(p_input[11770]), .Z(o[1770]) );
  AND U9146 ( .A(p_input[176]), .B(p_input[10176]), .Z(o[176]) );
  AND U9147 ( .A(p_input[1769]), .B(p_input[11769]), .Z(o[1769]) );
  AND U9148 ( .A(p_input[1768]), .B(p_input[11768]), .Z(o[1768]) );
  AND U9149 ( .A(p_input[1767]), .B(p_input[11767]), .Z(o[1767]) );
  AND U9150 ( .A(p_input[1766]), .B(p_input[11766]), .Z(o[1766]) );
  AND U9151 ( .A(p_input[1765]), .B(p_input[11765]), .Z(o[1765]) );
  AND U9152 ( .A(p_input[1764]), .B(p_input[11764]), .Z(o[1764]) );
  AND U9153 ( .A(p_input[1763]), .B(p_input[11763]), .Z(o[1763]) );
  AND U9154 ( .A(p_input[1762]), .B(p_input[11762]), .Z(o[1762]) );
  AND U9155 ( .A(p_input[1761]), .B(p_input[11761]), .Z(o[1761]) );
  AND U9156 ( .A(p_input[1760]), .B(p_input[11760]), .Z(o[1760]) );
  AND U9157 ( .A(p_input[175]), .B(p_input[10175]), .Z(o[175]) );
  AND U9158 ( .A(p_input[1759]), .B(p_input[11759]), .Z(o[1759]) );
  AND U9159 ( .A(p_input[1758]), .B(p_input[11758]), .Z(o[1758]) );
  AND U9160 ( .A(p_input[1757]), .B(p_input[11757]), .Z(o[1757]) );
  AND U9161 ( .A(p_input[1756]), .B(p_input[11756]), .Z(o[1756]) );
  AND U9162 ( .A(p_input[1755]), .B(p_input[11755]), .Z(o[1755]) );
  AND U9163 ( .A(p_input[1754]), .B(p_input[11754]), .Z(o[1754]) );
  AND U9164 ( .A(p_input[1753]), .B(p_input[11753]), .Z(o[1753]) );
  AND U9165 ( .A(p_input[1752]), .B(p_input[11752]), .Z(o[1752]) );
  AND U9166 ( .A(p_input[1751]), .B(p_input[11751]), .Z(o[1751]) );
  AND U9167 ( .A(p_input[1750]), .B(p_input[11750]), .Z(o[1750]) );
  AND U9168 ( .A(p_input[174]), .B(p_input[10174]), .Z(o[174]) );
  AND U9169 ( .A(p_input[1749]), .B(p_input[11749]), .Z(o[1749]) );
  AND U9170 ( .A(p_input[1748]), .B(p_input[11748]), .Z(o[1748]) );
  AND U9171 ( .A(p_input[1747]), .B(p_input[11747]), .Z(o[1747]) );
  AND U9172 ( .A(p_input[1746]), .B(p_input[11746]), .Z(o[1746]) );
  AND U9173 ( .A(p_input[1745]), .B(p_input[11745]), .Z(o[1745]) );
  AND U9174 ( .A(p_input[1744]), .B(p_input[11744]), .Z(o[1744]) );
  AND U9175 ( .A(p_input[1743]), .B(p_input[11743]), .Z(o[1743]) );
  AND U9176 ( .A(p_input[1742]), .B(p_input[11742]), .Z(o[1742]) );
  AND U9177 ( .A(p_input[1741]), .B(p_input[11741]), .Z(o[1741]) );
  AND U9178 ( .A(p_input[1740]), .B(p_input[11740]), .Z(o[1740]) );
  AND U9179 ( .A(p_input[173]), .B(p_input[10173]), .Z(o[173]) );
  AND U9180 ( .A(p_input[1739]), .B(p_input[11739]), .Z(o[1739]) );
  AND U9181 ( .A(p_input[1738]), .B(p_input[11738]), .Z(o[1738]) );
  AND U9182 ( .A(p_input[1737]), .B(p_input[11737]), .Z(o[1737]) );
  AND U9183 ( .A(p_input[1736]), .B(p_input[11736]), .Z(o[1736]) );
  AND U9184 ( .A(p_input[1735]), .B(p_input[11735]), .Z(o[1735]) );
  AND U9185 ( .A(p_input[1734]), .B(p_input[11734]), .Z(o[1734]) );
  AND U9186 ( .A(p_input[1733]), .B(p_input[11733]), .Z(o[1733]) );
  AND U9187 ( .A(p_input[1732]), .B(p_input[11732]), .Z(o[1732]) );
  AND U9188 ( .A(p_input[1731]), .B(p_input[11731]), .Z(o[1731]) );
  AND U9189 ( .A(p_input[1730]), .B(p_input[11730]), .Z(o[1730]) );
  AND U9190 ( .A(p_input[172]), .B(p_input[10172]), .Z(o[172]) );
  AND U9191 ( .A(p_input[1729]), .B(p_input[11729]), .Z(o[1729]) );
  AND U9192 ( .A(p_input[1728]), .B(p_input[11728]), .Z(o[1728]) );
  AND U9193 ( .A(p_input[1727]), .B(p_input[11727]), .Z(o[1727]) );
  AND U9194 ( .A(p_input[1726]), .B(p_input[11726]), .Z(o[1726]) );
  AND U9195 ( .A(p_input[1725]), .B(p_input[11725]), .Z(o[1725]) );
  AND U9196 ( .A(p_input[1724]), .B(p_input[11724]), .Z(o[1724]) );
  AND U9197 ( .A(p_input[1723]), .B(p_input[11723]), .Z(o[1723]) );
  AND U9198 ( .A(p_input[1722]), .B(p_input[11722]), .Z(o[1722]) );
  AND U9199 ( .A(p_input[1721]), .B(p_input[11721]), .Z(o[1721]) );
  AND U9200 ( .A(p_input[1720]), .B(p_input[11720]), .Z(o[1720]) );
  AND U9201 ( .A(p_input[171]), .B(p_input[10171]), .Z(o[171]) );
  AND U9202 ( .A(p_input[1719]), .B(p_input[11719]), .Z(o[1719]) );
  AND U9203 ( .A(p_input[1718]), .B(p_input[11718]), .Z(o[1718]) );
  AND U9204 ( .A(p_input[1717]), .B(p_input[11717]), .Z(o[1717]) );
  AND U9205 ( .A(p_input[1716]), .B(p_input[11716]), .Z(o[1716]) );
  AND U9206 ( .A(p_input[1715]), .B(p_input[11715]), .Z(o[1715]) );
  AND U9207 ( .A(p_input[1714]), .B(p_input[11714]), .Z(o[1714]) );
  AND U9208 ( .A(p_input[1713]), .B(p_input[11713]), .Z(o[1713]) );
  AND U9209 ( .A(p_input[1712]), .B(p_input[11712]), .Z(o[1712]) );
  AND U9210 ( .A(p_input[1711]), .B(p_input[11711]), .Z(o[1711]) );
  AND U9211 ( .A(p_input[1710]), .B(p_input[11710]), .Z(o[1710]) );
  AND U9212 ( .A(p_input[170]), .B(p_input[10170]), .Z(o[170]) );
  AND U9213 ( .A(p_input[1709]), .B(p_input[11709]), .Z(o[1709]) );
  AND U9214 ( .A(p_input[1708]), .B(p_input[11708]), .Z(o[1708]) );
  AND U9215 ( .A(p_input[1707]), .B(p_input[11707]), .Z(o[1707]) );
  AND U9216 ( .A(p_input[1706]), .B(p_input[11706]), .Z(o[1706]) );
  AND U9217 ( .A(p_input[1705]), .B(p_input[11705]), .Z(o[1705]) );
  AND U9218 ( .A(p_input[1704]), .B(p_input[11704]), .Z(o[1704]) );
  AND U9219 ( .A(p_input[1703]), .B(p_input[11703]), .Z(o[1703]) );
  AND U9220 ( .A(p_input[1702]), .B(p_input[11702]), .Z(o[1702]) );
  AND U9221 ( .A(p_input[1701]), .B(p_input[11701]), .Z(o[1701]) );
  AND U9222 ( .A(p_input[1700]), .B(p_input[11700]), .Z(o[1700]) );
  AND U9223 ( .A(p_input[16]), .B(p_input[10016]), .Z(o[16]) );
  AND U9224 ( .A(p_input[169]), .B(p_input[10169]), .Z(o[169]) );
  AND U9225 ( .A(p_input[1699]), .B(p_input[11699]), .Z(o[1699]) );
  AND U9226 ( .A(p_input[1698]), .B(p_input[11698]), .Z(o[1698]) );
  AND U9227 ( .A(p_input[1697]), .B(p_input[11697]), .Z(o[1697]) );
  AND U9228 ( .A(p_input[1696]), .B(p_input[11696]), .Z(o[1696]) );
  AND U9229 ( .A(p_input[1695]), .B(p_input[11695]), .Z(o[1695]) );
  AND U9230 ( .A(p_input[1694]), .B(p_input[11694]), .Z(o[1694]) );
  AND U9231 ( .A(p_input[1693]), .B(p_input[11693]), .Z(o[1693]) );
  AND U9232 ( .A(p_input[1692]), .B(p_input[11692]), .Z(o[1692]) );
  AND U9233 ( .A(p_input[1691]), .B(p_input[11691]), .Z(o[1691]) );
  AND U9234 ( .A(p_input[1690]), .B(p_input[11690]), .Z(o[1690]) );
  AND U9235 ( .A(p_input[168]), .B(p_input[10168]), .Z(o[168]) );
  AND U9236 ( .A(p_input[1689]), .B(p_input[11689]), .Z(o[1689]) );
  AND U9237 ( .A(p_input[1688]), .B(p_input[11688]), .Z(o[1688]) );
  AND U9238 ( .A(p_input[1687]), .B(p_input[11687]), .Z(o[1687]) );
  AND U9239 ( .A(p_input[1686]), .B(p_input[11686]), .Z(o[1686]) );
  AND U9240 ( .A(p_input[1685]), .B(p_input[11685]), .Z(o[1685]) );
  AND U9241 ( .A(p_input[1684]), .B(p_input[11684]), .Z(o[1684]) );
  AND U9242 ( .A(p_input[1683]), .B(p_input[11683]), .Z(o[1683]) );
  AND U9243 ( .A(p_input[1682]), .B(p_input[11682]), .Z(o[1682]) );
  AND U9244 ( .A(p_input[1681]), .B(p_input[11681]), .Z(o[1681]) );
  AND U9245 ( .A(p_input[1680]), .B(p_input[11680]), .Z(o[1680]) );
  AND U9246 ( .A(p_input[167]), .B(p_input[10167]), .Z(o[167]) );
  AND U9247 ( .A(p_input[1679]), .B(p_input[11679]), .Z(o[1679]) );
  AND U9248 ( .A(p_input[1678]), .B(p_input[11678]), .Z(o[1678]) );
  AND U9249 ( .A(p_input[1677]), .B(p_input[11677]), .Z(o[1677]) );
  AND U9250 ( .A(p_input[1676]), .B(p_input[11676]), .Z(o[1676]) );
  AND U9251 ( .A(p_input[1675]), .B(p_input[11675]), .Z(o[1675]) );
  AND U9252 ( .A(p_input[1674]), .B(p_input[11674]), .Z(o[1674]) );
  AND U9253 ( .A(p_input[1673]), .B(p_input[11673]), .Z(o[1673]) );
  AND U9254 ( .A(p_input[1672]), .B(p_input[11672]), .Z(o[1672]) );
  AND U9255 ( .A(p_input[1671]), .B(p_input[11671]), .Z(o[1671]) );
  AND U9256 ( .A(p_input[1670]), .B(p_input[11670]), .Z(o[1670]) );
  AND U9257 ( .A(p_input[166]), .B(p_input[10166]), .Z(o[166]) );
  AND U9258 ( .A(p_input[1669]), .B(p_input[11669]), .Z(o[1669]) );
  AND U9259 ( .A(p_input[1668]), .B(p_input[11668]), .Z(o[1668]) );
  AND U9260 ( .A(p_input[1667]), .B(p_input[11667]), .Z(o[1667]) );
  AND U9261 ( .A(p_input[1666]), .B(p_input[11666]), .Z(o[1666]) );
  AND U9262 ( .A(p_input[1665]), .B(p_input[11665]), .Z(o[1665]) );
  AND U9263 ( .A(p_input[1664]), .B(p_input[11664]), .Z(o[1664]) );
  AND U9264 ( .A(p_input[1663]), .B(p_input[11663]), .Z(o[1663]) );
  AND U9265 ( .A(p_input[1662]), .B(p_input[11662]), .Z(o[1662]) );
  AND U9266 ( .A(p_input[1661]), .B(p_input[11661]), .Z(o[1661]) );
  AND U9267 ( .A(p_input[1660]), .B(p_input[11660]), .Z(o[1660]) );
  AND U9268 ( .A(p_input[165]), .B(p_input[10165]), .Z(o[165]) );
  AND U9269 ( .A(p_input[1659]), .B(p_input[11659]), .Z(o[1659]) );
  AND U9270 ( .A(p_input[1658]), .B(p_input[11658]), .Z(o[1658]) );
  AND U9271 ( .A(p_input[1657]), .B(p_input[11657]), .Z(o[1657]) );
  AND U9272 ( .A(p_input[1656]), .B(p_input[11656]), .Z(o[1656]) );
  AND U9273 ( .A(p_input[1655]), .B(p_input[11655]), .Z(o[1655]) );
  AND U9274 ( .A(p_input[1654]), .B(p_input[11654]), .Z(o[1654]) );
  AND U9275 ( .A(p_input[1653]), .B(p_input[11653]), .Z(o[1653]) );
  AND U9276 ( .A(p_input[1652]), .B(p_input[11652]), .Z(o[1652]) );
  AND U9277 ( .A(p_input[1651]), .B(p_input[11651]), .Z(o[1651]) );
  AND U9278 ( .A(p_input[1650]), .B(p_input[11650]), .Z(o[1650]) );
  AND U9279 ( .A(p_input[164]), .B(p_input[10164]), .Z(o[164]) );
  AND U9280 ( .A(p_input[1649]), .B(p_input[11649]), .Z(o[1649]) );
  AND U9281 ( .A(p_input[1648]), .B(p_input[11648]), .Z(o[1648]) );
  AND U9282 ( .A(p_input[1647]), .B(p_input[11647]), .Z(o[1647]) );
  AND U9283 ( .A(p_input[1646]), .B(p_input[11646]), .Z(o[1646]) );
  AND U9284 ( .A(p_input[1645]), .B(p_input[11645]), .Z(o[1645]) );
  AND U9285 ( .A(p_input[1644]), .B(p_input[11644]), .Z(o[1644]) );
  AND U9286 ( .A(p_input[1643]), .B(p_input[11643]), .Z(o[1643]) );
  AND U9287 ( .A(p_input[1642]), .B(p_input[11642]), .Z(o[1642]) );
  AND U9288 ( .A(p_input[1641]), .B(p_input[11641]), .Z(o[1641]) );
  AND U9289 ( .A(p_input[1640]), .B(p_input[11640]), .Z(o[1640]) );
  AND U9290 ( .A(p_input[163]), .B(p_input[10163]), .Z(o[163]) );
  AND U9291 ( .A(p_input[1639]), .B(p_input[11639]), .Z(o[1639]) );
  AND U9292 ( .A(p_input[1638]), .B(p_input[11638]), .Z(o[1638]) );
  AND U9293 ( .A(p_input[1637]), .B(p_input[11637]), .Z(o[1637]) );
  AND U9294 ( .A(p_input[1636]), .B(p_input[11636]), .Z(o[1636]) );
  AND U9295 ( .A(p_input[1635]), .B(p_input[11635]), .Z(o[1635]) );
  AND U9296 ( .A(p_input[1634]), .B(p_input[11634]), .Z(o[1634]) );
  AND U9297 ( .A(p_input[1633]), .B(p_input[11633]), .Z(o[1633]) );
  AND U9298 ( .A(p_input[1632]), .B(p_input[11632]), .Z(o[1632]) );
  AND U9299 ( .A(p_input[1631]), .B(p_input[11631]), .Z(o[1631]) );
  AND U9300 ( .A(p_input[1630]), .B(p_input[11630]), .Z(o[1630]) );
  AND U9301 ( .A(p_input[162]), .B(p_input[10162]), .Z(o[162]) );
  AND U9302 ( .A(p_input[1629]), .B(p_input[11629]), .Z(o[1629]) );
  AND U9303 ( .A(p_input[1628]), .B(p_input[11628]), .Z(o[1628]) );
  AND U9304 ( .A(p_input[1627]), .B(p_input[11627]), .Z(o[1627]) );
  AND U9305 ( .A(p_input[1626]), .B(p_input[11626]), .Z(o[1626]) );
  AND U9306 ( .A(p_input[1625]), .B(p_input[11625]), .Z(o[1625]) );
  AND U9307 ( .A(p_input[1624]), .B(p_input[11624]), .Z(o[1624]) );
  AND U9308 ( .A(p_input[1623]), .B(p_input[11623]), .Z(o[1623]) );
  AND U9309 ( .A(p_input[1622]), .B(p_input[11622]), .Z(o[1622]) );
  AND U9310 ( .A(p_input[1621]), .B(p_input[11621]), .Z(o[1621]) );
  AND U9311 ( .A(p_input[1620]), .B(p_input[11620]), .Z(o[1620]) );
  AND U9312 ( .A(p_input[161]), .B(p_input[10161]), .Z(o[161]) );
  AND U9313 ( .A(p_input[1619]), .B(p_input[11619]), .Z(o[1619]) );
  AND U9314 ( .A(p_input[1618]), .B(p_input[11618]), .Z(o[1618]) );
  AND U9315 ( .A(p_input[1617]), .B(p_input[11617]), .Z(o[1617]) );
  AND U9316 ( .A(p_input[1616]), .B(p_input[11616]), .Z(o[1616]) );
  AND U9317 ( .A(p_input[1615]), .B(p_input[11615]), .Z(o[1615]) );
  AND U9318 ( .A(p_input[1614]), .B(p_input[11614]), .Z(o[1614]) );
  AND U9319 ( .A(p_input[1613]), .B(p_input[11613]), .Z(o[1613]) );
  AND U9320 ( .A(p_input[1612]), .B(p_input[11612]), .Z(o[1612]) );
  AND U9321 ( .A(p_input[1611]), .B(p_input[11611]), .Z(o[1611]) );
  AND U9322 ( .A(p_input[1610]), .B(p_input[11610]), .Z(o[1610]) );
  AND U9323 ( .A(p_input[160]), .B(p_input[10160]), .Z(o[160]) );
  AND U9324 ( .A(p_input[1609]), .B(p_input[11609]), .Z(o[1609]) );
  AND U9325 ( .A(p_input[1608]), .B(p_input[11608]), .Z(o[1608]) );
  AND U9326 ( .A(p_input[1607]), .B(p_input[11607]), .Z(o[1607]) );
  AND U9327 ( .A(p_input[1606]), .B(p_input[11606]), .Z(o[1606]) );
  AND U9328 ( .A(p_input[1605]), .B(p_input[11605]), .Z(o[1605]) );
  AND U9329 ( .A(p_input[1604]), .B(p_input[11604]), .Z(o[1604]) );
  AND U9330 ( .A(p_input[1603]), .B(p_input[11603]), .Z(o[1603]) );
  AND U9331 ( .A(p_input[1602]), .B(p_input[11602]), .Z(o[1602]) );
  AND U9332 ( .A(p_input[1601]), .B(p_input[11601]), .Z(o[1601]) );
  AND U9333 ( .A(p_input[1600]), .B(p_input[11600]), .Z(o[1600]) );
  AND U9334 ( .A(p_input[15]), .B(p_input[10015]), .Z(o[15]) );
  AND U9335 ( .A(p_input[159]), .B(p_input[10159]), .Z(o[159]) );
  AND U9336 ( .A(p_input[1599]), .B(p_input[11599]), .Z(o[1599]) );
  AND U9337 ( .A(p_input[1598]), .B(p_input[11598]), .Z(o[1598]) );
  AND U9338 ( .A(p_input[1597]), .B(p_input[11597]), .Z(o[1597]) );
  AND U9339 ( .A(p_input[1596]), .B(p_input[11596]), .Z(o[1596]) );
  AND U9340 ( .A(p_input[1595]), .B(p_input[11595]), .Z(o[1595]) );
  AND U9341 ( .A(p_input[1594]), .B(p_input[11594]), .Z(o[1594]) );
  AND U9342 ( .A(p_input[1593]), .B(p_input[11593]), .Z(o[1593]) );
  AND U9343 ( .A(p_input[1592]), .B(p_input[11592]), .Z(o[1592]) );
  AND U9344 ( .A(p_input[1591]), .B(p_input[11591]), .Z(o[1591]) );
  AND U9345 ( .A(p_input[1590]), .B(p_input[11590]), .Z(o[1590]) );
  AND U9346 ( .A(p_input[158]), .B(p_input[10158]), .Z(o[158]) );
  AND U9347 ( .A(p_input[1589]), .B(p_input[11589]), .Z(o[1589]) );
  AND U9348 ( .A(p_input[1588]), .B(p_input[11588]), .Z(o[1588]) );
  AND U9349 ( .A(p_input[1587]), .B(p_input[11587]), .Z(o[1587]) );
  AND U9350 ( .A(p_input[1586]), .B(p_input[11586]), .Z(o[1586]) );
  AND U9351 ( .A(p_input[1585]), .B(p_input[11585]), .Z(o[1585]) );
  AND U9352 ( .A(p_input[1584]), .B(p_input[11584]), .Z(o[1584]) );
  AND U9353 ( .A(p_input[1583]), .B(p_input[11583]), .Z(o[1583]) );
  AND U9354 ( .A(p_input[1582]), .B(p_input[11582]), .Z(o[1582]) );
  AND U9355 ( .A(p_input[1581]), .B(p_input[11581]), .Z(o[1581]) );
  AND U9356 ( .A(p_input[1580]), .B(p_input[11580]), .Z(o[1580]) );
  AND U9357 ( .A(p_input[157]), .B(p_input[10157]), .Z(o[157]) );
  AND U9358 ( .A(p_input[1579]), .B(p_input[11579]), .Z(o[1579]) );
  AND U9359 ( .A(p_input[1578]), .B(p_input[11578]), .Z(o[1578]) );
  AND U9360 ( .A(p_input[1577]), .B(p_input[11577]), .Z(o[1577]) );
  AND U9361 ( .A(p_input[1576]), .B(p_input[11576]), .Z(o[1576]) );
  AND U9362 ( .A(p_input[1575]), .B(p_input[11575]), .Z(o[1575]) );
  AND U9363 ( .A(p_input[1574]), .B(p_input[11574]), .Z(o[1574]) );
  AND U9364 ( .A(p_input[1573]), .B(p_input[11573]), .Z(o[1573]) );
  AND U9365 ( .A(p_input[1572]), .B(p_input[11572]), .Z(o[1572]) );
  AND U9366 ( .A(p_input[1571]), .B(p_input[11571]), .Z(o[1571]) );
  AND U9367 ( .A(p_input[1570]), .B(p_input[11570]), .Z(o[1570]) );
  AND U9368 ( .A(p_input[156]), .B(p_input[10156]), .Z(o[156]) );
  AND U9369 ( .A(p_input[1569]), .B(p_input[11569]), .Z(o[1569]) );
  AND U9370 ( .A(p_input[1568]), .B(p_input[11568]), .Z(o[1568]) );
  AND U9371 ( .A(p_input[1567]), .B(p_input[11567]), .Z(o[1567]) );
  AND U9372 ( .A(p_input[1566]), .B(p_input[11566]), .Z(o[1566]) );
  AND U9373 ( .A(p_input[1565]), .B(p_input[11565]), .Z(o[1565]) );
  AND U9374 ( .A(p_input[1564]), .B(p_input[11564]), .Z(o[1564]) );
  AND U9375 ( .A(p_input[1563]), .B(p_input[11563]), .Z(o[1563]) );
  AND U9376 ( .A(p_input[1562]), .B(p_input[11562]), .Z(o[1562]) );
  AND U9377 ( .A(p_input[1561]), .B(p_input[11561]), .Z(o[1561]) );
  AND U9378 ( .A(p_input[1560]), .B(p_input[11560]), .Z(o[1560]) );
  AND U9379 ( .A(p_input[155]), .B(p_input[10155]), .Z(o[155]) );
  AND U9380 ( .A(p_input[1559]), .B(p_input[11559]), .Z(o[1559]) );
  AND U9381 ( .A(p_input[1558]), .B(p_input[11558]), .Z(o[1558]) );
  AND U9382 ( .A(p_input[1557]), .B(p_input[11557]), .Z(o[1557]) );
  AND U9383 ( .A(p_input[1556]), .B(p_input[11556]), .Z(o[1556]) );
  AND U9384 ( .A(p_input[1555]), .B(p_input[11555]), .Z(o[1555]) );
  AND U9385 ( .A(p_input[1554]), .B(p_input[11554]), .Z(o[1554]) );
  AND U9386 ( .A(p_input[1553]), .B(p_input[11553]), .Z(o[1553]) );
  AND U9387 ( .A(p_input[1552]), .B(p_input[11552]), .Z(o[1552]) );
  AND U9388 ( .A(p_input[1551]), .B(p_input[11551]), .Z(o[1551]) );
  AND U9389 ( .A(p_input[1550]), .B(p_input[11550]), .Z(o[1550]) );
  AND U9390 ( .A(p_input[154]), .B(p_input[10154]), .Z(o[154]) );
  AND U9391 ( .A(p_input[1549]), .B(p_input[11549]), .Z(o[1549]) );
  AND U9392 ( .A(p_input[1548]), .B(p_input[11548]), .Z(o[1548]) );
  AND U9393 ( .A(p_input[1547]), .B(p_input[11547]), .Z(o[1547]) );
  AND U9394 ( .A(p_input[1546]), .B(p_input[11546]), .Z(o[1546]) );
  AND U9395 ( .A(p_input[1545]), .B(p_input[11545]), .Z(o[1545]) );
  AND U9396 ( .A(p_input[1544]), .B(p_input[11544]), .Z(o[1544]) );
  AND U9397 ( .A(p_input[1543]), .B(p_input[11543]), .Z(o[1543]) );
  AND U9398 ( .A(p_input[1542]), .B(p_input[11542]), .Z(o[1542]) );
  AND U9399 ( .A(p_input[1541]), .B(p_input[11541]), .Z(o[1541]) );
  AND U9400 ( .A(p_input[1540]), .B(p_input[11540]), .Z(o[1540]) );
  AND U9401 ( .A(p_input[153]), .B(p_input[10153]), .Z(o[153]) );
  AND U9402 ( .A(p_input[1539]), .B(p_input[11539]), .Z(o[1539]) );
  AND U9403 ( .A(p_input[1538]), .B(p_input[11538]), .Z(o[1538]) );
  AND U9404 ( .A(p_input[1537]), .B(p_input[11537]), .Z(o[1537]) );
  AND U9405 ( .A(p_input[1536]), .B(p_input[11536]), .Z(o[1536]) );
  AND U9406 ( .A(p_input[1535]), .B(p_input[11535]), .Z(o[1535]) );
  AND U9407 ( .A(p_input[1534]), .B(p_input[11534]), .Z(o[1534]) );
  AND U9408 ( .A(p_input[1533]), .B(p_input[11533]), .Z(o[1533]) );
  AND U9409 ( .A(p_input[1532]), .B(p_input[11532]), .Z(o[1532]) );
  AND U9410 ( .A(p_input[1531]), .B(p_input[11531]), .Z(o[1531]) );
  AND U9411 ( .A(p_input[1530]), .B(p_input[11530]), .Z(o[1530]) );
  AND U9412 ( .A(p_input[152]), .B(p_input[10152]), .Z(o[152]) );
  AND U9413 ( .A(p_input[1529]), .B(p_input[11529]), .Z(o[1529]) );
  AND U9414 ( .A(p_input[1528]), .B(p_input[11528]), .Z(o[1528]) );
  AND U9415 ( .A(p_input[1527]), .B(p_input[11527]), .Z(o[1527]) );
  AND U9416 ( .A(p_input[1526]), .B(p_input[11526]), .Z(o[1526]) );
  AND U9417 ( .A(p_input[1525]), .B(p_input[11525]), .Z(o[1525]) );
  AND U9418 ( .A(p_input[1524]), .B(p_input[11524]), .Z(o[1524]) );
  AND U9419 ( .A(p_input[1523]), .B(p_input[11523]), .Z(o[1523]) );
  AND U9420 ( .A(p_input[1522]), .B(p_input[11522]), .Z(o[1522]) );
  AND U9421 ( .A(p_input[1521]), .B(p_input[11521]), .Z(o[1521]) );
  AND U9422 ( .A(p_input[1520]), .B(p_input[11520]), .Z(o[1520]) );
  AND U9423 ( .A(p_input[151]), .B(p_input[10151]), .Z(o[151]) );
  AND U9424 ( .A(p_input[1519]), .B(p_input[11519]), .Z(o[1519]) );
  AND U9425 ( .A(p_input[1518]), .B(p_input[11518]), .Z(o[1518]) );
  AND U9426 ( .A(p_input[1517]), .B(p_input[11517]), .Z(o[1517]) );
  AND U9427 ( .A(p_input[1516]), .B(p_input[11516]), .Z(o[1516]) );
  AND U9428 ( .A(p_input[1515]), .B(p_input[11515]), .Z(o[1515]) );
  AND U9429 ( .A(p_input[1514]), .B(p_input[11514]), .Z(o[1514]) );
  AND U9430 ( .A(p_input[1513]), .B(p_input[11513]), .Z(o[1513]) );
  AND U9431 ( .A(p_input[1512]), .B(p_input[11512]), .Z(o[1512]) );
  AND U9432 ( .A(p_input[1511]), .B(p_input[11511]), .Z(o[1511]) );
  AND U9433 ( .A(p_input[1510]), .B(p_input[11510]), .Z(o[1510]) );
  AND U9434 ( .A(p_input[150]), .B(p_input[10150]), .Z(o[150]) );
  AND U9435 ( .A(p_input[1509]), .B(p_input[11509]), .Z(o[1509]) );
  AND U9436 ( .A(p_input[1508]), .B(p_input[11508]), .Z(o[1508]) );
  AND U9437 ( .A(p_input[1507]), .B(p_input[11507]), .Z(o[1507]) );
  AND U9438 ( .A(p_input[1506]), .B(p_input[11506]), .Z(o[1506]) );
  AND U9439 ( .A(p_input[1505]), .B(p_input[11505]), .Z(o[1505]) );
  AND U9440 ( .A(p_input[1504]), .B(p_input[11504]), .Z(o[1504]) );
  AND U9441 ( .A(p_input[1503]), .B(p_input[11503]), .Z(o[1503]) );
  AND U9442 ( .A(p_input[1502]), .B(p_input[11502]), .Z(o[1502]) );
  AND U9443 ( .A(p_input[1501]), .B(p_input[11501]), .Z(o[1501]) );
  AND U9444 ( .A(p_input[1500]), .B(p_input[11500]), .Z(o[1500]) );
  AND U9445 ( .A(p_input[14]), .B(p_input[10014]), .Z(o[14]) );
  AND U9446 ( .A(p_input[149]), .B(p_input[10149]), .Z(o[149]) );
  AND U9447 ( .A(p_input[1499]), .B(p_input[11499]), .Z(o[1499]) );
  AND U9448 ( .A(p_input[1498]), .B(p_input[11498]), .Z(o[1498]) );
  AND U9449 ( .A(p_input[1497]), .B(p_input[11497]), .Z(o[1497]) );
  AND U9450 ( .A(p_input[1496]), .B(p_input[11496]), .Z(o[1496]) );
  AND U9451 ( .A(p_input[1495]), .B(p_input[11495]), .Z(o[1495]) );
  AND U9452 ( .A(p_input[1494]), .B(p_input[11494]), .Z(o[1494]) );
  AND U9453 ( .A(p_input[1493]), .B(p_input[11493]), .Z(o[1493]) );
  AND U9454 ( .A(p_input[1492]), .B(p_input[11492]), .Z(o[1492]) );
  AND U9455 ( .A(p_input[1491]), .B(p_input[11491]), .Z(o[1491]) );
  AND U9456 ( .A(p_input[1490]), .B(p_input[11490]), .Z(o[1490]) );
  AND U9457 ( .A(p_input[148]), .B(p_input[10148]), .Z(o[148]) );
  AND U9458 ( .A(p_input[1489]), .B(p_input[11489]), .Z(o[1489]) );
  AND U9459 ( .A(p_input[1488]), .B(p_input[11488]), .Z(o[1488]) );
  AND U9460 ( .A(p_input[1487]), .B(p_input[11487]), .Z(o[1487]) );
  AND U9461 ( .A(p_input[1486]), .B(p_input[11486]), .Z(o[1486]) );
  AND U9462 ( .A(p_input[1485]), .B(p_input[11485]), .Z(o[1485]) );
  AND U9463 ( .A(p_input[1484]), .B(p_input[11484]), .Z(o[1484]) );
  AND U9464 ( .A(p_input[1483]), .B(p_input[11483]), .Z(o[1483]) );
  AND U9465 ( .A(p_input[1482]), .B(p_input[11482]), .Z(o[1482]) );
  AND U9466 ( .A(p_input[1481]), .B(p_input[11481]), .Z(o[1481]) );
  AND U9467 ( .A(p_input[1480]), .B(p_input[11480]), .Z(o[1480]) );
  AND U9468 ( .A(p_input[147]), .B(p_input[10147]), .Z(o[147]) );
  AND U9469 ( .A(p_input[1479]), .B(p_input[11479]), .Z(o[1479]) );
  AND U9470 ( .A(p_input[1478]), .B(p_input[11478]), .Z(o[1478]) );
  AND U9471 ( .A(p_input[1477]), .B(p_input[11477]), .Z(o[1477]) );
  AND U9472 ( .A(p_input[1476]), .B(p_input[11476]), .Z(o[1476]) );
  AND U9473 ( .A(p_input[1475]), .B(p_input[11475]), .Z(o[1475]) );
  AND U9474 ( .A(p_input[1474]), .B(p_input[11474]), .Z(o[1474]) );
  AND U9475 ( .A(p_input[1473]), .B(p_input[11473]), .Z(o[1473]) );
  AND U9476 ( .A(p_input[1472]), .B(p_input[11472]), .Z(o[1472]) );
  AND U9477 ( .A(p_input[1471]), .B(p_input[11471]), .Z(o[1471]) );
  AND U9478 ( .A(p_input[1470]), .B(p_input[11470]), .Z(o[1470]) );
  AND U9479 ( .A(p_input[146]), .B(p_input[10146]), .Z(o[146]) );
  AND U9480 ( .A(p_input[1469]), .B(p_input[11469]), .Z(o[1469]) );
  AND U9481 ( .A(p_input[1468]), .B(p_input[11468]), .Z(o[1468]) );
  AND U9482 ( .A(p_input[1467]), .B(p_input[11467]), .Z(o[1467]) );
  AND U9483 ( .A(p_input[1466]), .B(p_input[11466]), .Z(o[1466]) );
  AND U9484 ( .A(p_input[1465]), .B(p_input[11465]), .Z(o[1465]) );
  AND U9485 ( .A(p_input[1464]), .B(p_input[11464]), .Z(o[1464]) );
  AND U9486 ( .A(p_input[1463]), .B(p_input[11463]), .Z(o[1463]) );
  AND U9487 ( .A(p_input[1462]), .B(p_input[11462]), .Z(o[1462]) );
  AND U9488 ( .A(p_input[1461]), .B(p_input[11461]), .Z(o[1461]) );
  AND U9489 ( .A(p_input[1460]), .B(p_input[11460]), .Z(o[1460]) );
  AND U9490 ( .A(p_input[145]), .B(p_input[10145]), .Z(o[145]) );
  AND U9491 ( .A(p_input[1459]), .B(p_input[11459]), .Z(o[1459]) );
  AND U9492 ( .A(p_input[1458]), .B(p_input[11458]), .Z(o[1458]) );
  AND U9493 ( .A(p_input[1457]), .B(p_input[11457]), .Z(o[1457]) );
  AND U9494 ( .A(p_input[1456]), .B(p_input[11456]), .Z(o[1456]) );
  AND U9495 ( .A(p_input[1455]), .B(p_input[11455]), .Z(o[1455]) );
  AND U9496 ( .A(p_input[1454]), .B(p_input[11454]), .Z(o[1454]) );
  AND U9497 ( .A(p_input[1453]), .B(p_input[11453]), .Z(o[1453]) );
  AND U9498 ( .A(p_input[1452]), .B(p_input[11452]), .Z(o[1452]) );
  AND U9499 ( .A(p_input[1451]), .B(p_input[11451]), .Z(o[1451]) );
  AND U9500 ( .A(p_input[1450]), .B(p_input[11450]), .Z(o[1450]) );
  AND U9501 ( .A(p_input[144]), .B(p_input[10144]), .Z(o[144]) );
  AND U9502 ( .A(p_input[1449]), .B(p_input[11449]), .Z(o[1449]) );
  AND U9503 ( .A(p_input[1448]), .B(p_input[11448]), .Z(o[1448]) );
  AND U9504 ( .A(p_input[1447]), .B(p_input[11447]), .Z(o[1447]) );
  AND U9505 ( .A(p_input[1446]), .B(p_input[11446]), .Z(o[1446]) );
  AND U9506 ( .A(p_input[1445]), .B(p_input[11445]), .Z(o[1445]) );
  AND U9507 ( .A(p_input[1444]), .B(p_input[11444]), .Z(o[1444]) );
  AND U9508 ( .A(p_input[1443]), .B(p_input[11443]), .Z(o[1443]) );
  AND U9509 ( .A(p_input[1442]), .B(p_input[11442]), .Z(o[1442]) );
  AND U9510 ( .A(p_input[1441]), .B(p_input[11441]), .Z(o[1441]) );
  AND U9511 ( .A(p_input[1440]), .B(p_input[11440]), .Z(o[1440]) );
  AND U9512 ( .A(p_input[143]), .B(p_input[10143]), .Z(o[143]) );
  AND U9513 ( .A(p_input[1439]), .B(p_input[11439]), .Z(o[1439]) );
  AND U9514 ( .A(p_input[1438]), .B(p_input[11438]), .Z(o[1438]) );
  AND U9515 ( .A(p_input[1437]), .B(p_input[11437]), .Z(o[1437]) );
  AND U9516 ( .A(p_input[1436]), .B(p_input[11436]), .Z(o[1436]) );
  AND U9517 ( .A(p_input[1435]), .B(p_input[11435]), .Z(o[1435]) );
  AND U9518 ( .A(p_input[1434]), .B(p_input[11434]), .Z(o[1434]) );
  AND U9519 ( .A(p_input[1433]), .B(p_input[11433]), .Z(o[1433]) );
  AND U9520 ( .A(p_input[1432]), .B(p_input[11432]), .Z(o[1432]) );
  AND U9521 ( .A(p_input[1431]), .B(p_input[11431]), .Z(o[1431]) );
  AND U9522 ( .A(p_input[1430]), .B(p_input[11430]), .Z(o[1430]) );
  AND U9523 ( .A(p_input[142]), .B(p_input[10142]), .Z(o[142]) );
  AND U9524 ( .A(p_input[1429]), .B(p_input[11429]), .Z(o[1429]) );
  AND U9525 ( .A(p_input[1428]), .B(p_input[11428]), .Z(o[1428]) );
  AND U9526 ( .A(p_input[1427]), .B(p_input[11427]), .Z(o[1427]) );
  AND U9527 ( .A(p_input[1426]), .B(p_input[11426]), .Z(o[1426]) );
  AND U9528 ( .A(p_input[1425]), .B(p_input[11425]), .Z(o[1425]) );
  AND U9529 ( .A(p_input[1424]), .B(p_input[11424]), .Z(o[1424]) );
  AND U9530 ( .A(p_input[1423]), .B(p_input[11423]), .Z(o[1423]) );
  AND U9531 ( .A(p_input[1422]), .B(p_input[11422]), .Z(o[1422]) );
  AND U9532 ( .A(p_input[1421]), .B(p_input[11421]), .Z(o[1421]) );
  AND U9533 ( .A(p_input[1420]), .B(p_input[11420]), .Z(o[1420]) );
  AND U9534 ( .A(p_input[141]), .B(p_input[10141]), .Z(o[141]) );
  AND U9535 ( .A(p_input[1419]), .B(p_input[11419]), .Z(o[1419]) );
  AND U9536 ( .A(p_input[1418]), .B(p_input[11418]), .Z(o[1418]) );
  AND U9537 ( .A(p_input[1417]), .B(p_input[11417]), .Z(o[1417]) );
  AND U9538 ( .A(p_input[1416]), .B(p_input[11416]), .Z(o[1416]) );
  AND U9539 ( .A(p_input[1415]), .B(p_input[11415]), .Z(o[1415]) );
  AND U9540 ( .A(p_input[1414]), .B(p_input[11414]), .Z(o[1414]) );
  AND U9541 ( .A(p_input[1413]), .B(p_input[11413]), .Z(o[1413]) );
  AND U9542 ( .A(p_input[1412]), .B(p_input[11412]), .Z(o[1412]) );
  AND U9543 ( .A(p_input[1411]), .B(p_input[11411]), .Z(o[1411]) );
  AND U9544 ( .A(p_input[1410]), .B(p_input[11410]), .Z(o[1410]) );
  AND U9545 ( .A(p_input[140]), .B(p_input[10140]), .Z(o[140]) );
  AND U9546 ( .A(p_input[1409]), .B(p_input[11409]), .Z(o[1409]) );
  AND U9547 ( .A(p_input[1408]), .B(p_input[11408]), .Z(o[1408]) );
  AND U9548 ( .A(p_input[1407]), .B(p_input[11407]), .Z(o[1407]) );
  AND U9549 ( .A(p_input[1406]), .B(p_input[11406]), .Z(o[1406]) );
  AND U9550 ( .A(p_input[1405]), .B(p_input[11405]), .Z(o[1405]) );
  AND U9551 ( .A(p_input[1404]), .B(p_input[11404]), .Z(o[1404]) );
  AND U9552 ( .A(p_input[1403]), .B(p_input[11403]), .Z(o[1403]) );
  AND U9553 ( .A(p_input[1402]), .B(p_input[11402]), .Z(o[1402]) );
  AND U9554 ( .A(p_input[1401]), .B(p_input[11401]), .Z(o[1401]) );
  AND U9555 ( .A(p_input[1400]), .B(p_input[11400]), .Z(o[1400]) );
  AND U9556 ( .A(p_input[13]), .B(p_input[10013]), .Z(o[13]) );
  AND U9557 ( .A(p_input[139]), .B(p_input[10139]), .Z(o[139]) );
  AND U9558 ( .A(p_input[1399]), .B(p_input[11399]), .Z(o[1399]) );
  AND U9559 ( .A(p_input[1398]), .B(p_input[11398]), .Z(o[1398]) );
  AND U9560 ( .A(p_input[1397]), .B(p_input[11397]), .Z(o[1397]) );
  AND U9561 ( .A(p_input[1396]), .B(p_input[11396]), .Z(o[1396]) );
  AND U9562 ( .A(p_input[1395]), .B(p_input[11395]), .Z(o[1395]) );
  AND U9563 ( .A(p_input[1394]), .B(p_input[11394]), .Z(o[1394]) );
  AND U9564 ( .A(p_input[1393]), .B(p_input[11393]), .Z(o[1393]) );
  AND U9565 ( .A(p_input[1392]), .B(p_input[11392]), .Z(o[1392]) );
  AND U9566 ( .A(p_input[1391]), .B(p_input[11391]), .Z(o[1391]) );
  AND U9567 ( .A(p_input[1390]), .B(p_input[11390]), .Z(o[1390]) );
  AND U9568 ( .A(p_input[138]), .B(p_input[10138]), .Z(o[138]) );
  AND U9569 ( .A(p_input[1389]), .B(p_input[11389]), .Z(o[1389]) );
  AND U9570 ( .A(p_input[1388]), .B(p_input[11388]), .Z(o[1388]) );
  AND U9571 ( .A(p_input[1387]), .B(p_input[11387]), .Z(o[1387]) );
  AND U9572 ( .A(p_input[1386]), .B(p_input[11386]), .Z(o[1386]) );
  AND U9573 ( .A(p_input[1385]), .B(p_input[11385]), .Z(o[1385]) );
  AND U9574 ( .A(p_input[1384]), .B(p_input[11384]), .Z(o[1384]) );
  AND U9575 ( .A(p_input[1383]), .B(p_input[11383]), .Z(o[1383]) );
  AND U9576 ( .A(p_input[1382]), .B(p_input[11382]), .Z(o[1382]) );
  AND U9577 ( .A(p_input[1381]), .B(p_input[11381]), .Z(o[1381]) );
  AND U9578 ( .A(p_input[1380]), .B(p_input[11380]), .Z(o[1380]) );
  AND U9579 ( .A(p_input[137]), .B(p_input[10137]), .Z(o[137]) );
  AND U9580 ( .A(p_input[1379]), .B(p_input[11379]), .Z(o[1379]) );
  AND U9581 ( .A(p_input[1378]), .B(p_input[11378]), .Z(o[1378]) );
  AND U9582 ( .A(p_input[1377]), .B(p_input[11377]), .Z(o[1377]) );
  AND U9583 ( .A(p_input[1376]), .B(p_input[11376]), .Z(o[1376]) );
  AND U9584 ( .A(p_input[1375]), .B(p_input[11375]), .Z(o[1375]) );
  AND U9585 ( .A(p_input[1374]), .B(p_input[11374]), .Z(o[1374]) );
  AND U9586 ( .A(p_input[1373]), .B(p_input[11373]), .Z(o[1373]) );
  AND U9587 ( .A(p_input[1372]), .B(p_input[11372]), .Z(o[1372]) );
  AND U9588 ( .A(p_input[1371]), .B(p_input[11371]), .Z(o[1371]) );
  AND U9589 ( .A(p_input[1370]), .B(p_input[11370]), .Z(o[1370]) );
  AND U9590 ( .A(p_input[136]), .B(p_input[10136]), .Z(o[136]) );
  AND U9591 ( .A(p_input[1369]), .B(p_input[11369]), .Z(o[1369]) );
  AND U9592 ( .A(p_input[1368]), .B(p_input[11368]), .Z(o[1368]) );
  AND U9593 ( .A(p_input[1367]), .B(p_input[11367]), .Z(o[1367]) );
  AND U9594 ( .A(p_input[1366]), .B(p_input[11366]), .Z(o[1366]) );
  AND U9595 ( .A(p_input[1365]), .B(p_input[11365]), .Z(o[1365]) );
  AND U9596 ( .A(p_input[1364]), .B(p_input[11364]), .Z(o[1364]) );
  AND U9597 ( .A(p_input[1363]), .B(p_input[11363]), .Z(o[1363]) );
  AND U9598 ( .A(p_input[1362]), .B(p_input[11362]), .Z(o[1362]) );
  AND U9599 ( .A(p_input[1361]), .B(p_input[11361]), .Z(o[1361]) );
  AND U9600 ( .A(p_input[1360]), .B(p_input[11360]), .Z(o[1360]) );
  AND U9601 ( .A(p_input[135]), .B(p_input[10135]), .Z(o[135]) );
  AND U9602 ( .A(p_input[1359]), .B(p_input[11359]), .Z(o[1359]) );
  AND U9603 ( .A(p_input[1358]), .B(p_input[11358]), .Z(o[1358]) );
  AND U9604 ( .A(p_input[1357]), .B(p_input[11357]), .Z(o[1357]) );
  AND U9605 ( .A(p_input[1356]), .B(p_input[11356]), .Z(o[1356]) );
  AND U9606 ( .A(p_input[1355]), .B(p_input[11355]), .Z(o[1355]) );
  AND U9607 ( .A(p_input[1354]), .B(p_input[11354]), .Z(o[1354]) );
  AND U9608 ( .A(p_input[1353]), .B(p_input[11353]), .Z(o[1353]) );
  AND U9609 ( .A(p_input[1352]), .B(p_input[11352]), .Z(o[1352]) );
  AND U9610 ( .A(p_input[1351]), .B(p_input[11351]), .Z(o[1351]) );
  AND U9611 ( .A(p_input[1350]), .B(p_input[11350]), .Z(o[1350]) );
  AND U9612 ( .A(p_input[134]), .B(p_input[10134]), .Z(o[134]) );
  AND U9613 ( .A(p_input[1349]), .B(p_input[11349]), .Z(o[1349]) );
  AND U9614 ( .A(p_input[1348]), .B(p_input[11348]), .Z(o[1348]) );
  AND U9615 ( .A(p_input[1347]), .B(p_input[11347]), .Z(o[1347]) );
  AND U9616 ( .A(p_input[1346]), .B(p_input[11346]), .Z(o[1346]) );
  AND U9617 ( .A(p_input[1345]), .B(p_input[11345]), .Z(o[1345]) );
  AND U9618 ( .A(p_input[1344]), .B(p_input[11344]), .Z(o[1344]) );
  AND U9619 ( .A(p_input[1343]), .B(p_input[11343]), .Z(o[1343]) );
  AND U9620 ( .A(p_input[1342]), .B(p_input[11342]), .Z(o[1342]) );
  AND U9621 ( .A(p_input[1341]), .B(p_input[11341]), .Z(o[1341]) );
  AND U9622 ( .A(p_input[1340]), .B(p_input[11340]), .Z(o[1340]) );
  AND U9623 ( .A(p_input[133]), .B(p_input[10133]), .Z(o[133]) );
  AND U9624 ( .A(p_input[1339]), .B(p_input[11339]), .Z(o[1339]) );
  AND U9625 ( .A(p_input[1338]), .B(p_input[11338]), .Z(o[1338]) );
  AND U9626 ( .A(p_input[1337]), .B(p_input[11337]), .Z(o[1337]) );
  AND U9627 ( .A(p_input[1336]), .B(p_input[11336]), .Z(o[1336]) );
  AND U9628 ( .A(p_input[1335]), .B(p_input[11335]), .Z(o[1335]) );
  AND U9629 ( .A(p_input[1334]), .B(p_input[11334]), .Z(o[1334]) );
  AND U9630 ( .A(p_input[1333]), .B(p_input[11333]), .Z(o[1333]) );
  AND U9631 ( .A(p_input[1332]), .B(p_input[11332]), .Z(o[1332]) );
  AND U9632 ( .A(p_input[1331]), .B(p_input[11331]), .Z(o[1331]) );
  AND U9633 ( .A(p_input[1330]), .B(p_input[11330]), .Z(o[1330]) );
  AND U9634 ( .A(p_input[132]), .B(p_input[10132]), .Z(o[132]) );
  AND U9635 ( .A(p_input[1329]), .B(p_input[11329]), .Z(o[1329]) );
  AND U9636 ( .A(p_input[1328]), .B(p_input[11328]), .Z(o[1328]) );
  AND U9637 ( .A(p_input[1327]), .B(p_input[11327]), .Z(o[1327]) );
  AND U9638 ( .A(p_input[1326]), .B(p_input[11326]), .Z(o[1326]) );
  AND U9639 ( .A(p_input[1325]), .B(p_input[11325]), .Z(o[1325]) );
  AND U9640 ( .A(p_input[1324]), .B(p_input[11324]), .Z(o[1324]) );
  AND U9641 ( .A(p_input[1323]), .B(p_input[11323]), .Z(o[1323]) );
  AND U9642 ( .A(p_input[1322]), .B(p_input[11322]), .Z(o[1322]) );
  AND U9643 ( .A(p_input[1321]), .B(p_input[11321]), .Z(o[1321]) );
  AND U9644 ( .A(p_input[1320]), .B(p_input[11320]), .Z(o[1320]) );
  AND U9645 ( .A(p_input[131]), .B(p_input[10131]), .Z(o[131]) );
  AND U9646 ( .A(p_input[1319]), .B(p_input[11319]), .Z(o[1319]) );
  AND U9647 ( .A(p_input[1318]), .B(p_input[11318]), .Z(o[1318]) );
  AND U9648 ( .A(p_input[1317]), .B(p_input[11317]), .Z(o[1317]) );
  AND U9649 ( .A(p_input[1316]), .B(p_input[11316]), .Z(o[1316]) );
  AND U9650 ( .A(p_input[1315]), .B(p_input[11315]), .Z(o[1315]) );
  AND U9651 ( .A(p_input[1314]), .B(p_input[11314]), .Z(o[1314]) );
  AND U9652 ( .A(p_input[1313]), .B(p_input[11313]), .Z(o[1313]) );
  AND U9653 ( .A(p_input[1312]), .B(p_input[11312]), .Z(o[1312]) );
  AND U9654 ( .A(p_input[1311]), .B(p_input[11311]), .Z(o[1311]) );
  AND U9655 ( .A(p_input[1310]), .B(p_input[11310]), .Z(o[1310]) );
  AND U9656 ( .A(p_input[130]), .B(p_input[10130]), .Z(o[130]) );
  AND U9657 ( .A(p_input[1309]), .B(p_input[11309]), .Z(o[1309]) );
  AND U9658 ( .A(p_input[1308]), .B(p_input[11308]), .Z(o[1308]) );
  AND U9659 ( .A(p_input[1307]), .B(p_input[11307]), .Z(o[1307]) );
  AND U9660 ( .A(p_input[1306]), .B(p_input[11306]), .Z(o[1306]) );
  AND U9661 ( .A(p_input[1305]), .B(p_input[11305]), .Z(o[1305]) );
  AND U9662 ( .A(p_input[1304]), .B(p_input[11304]), .Z(o[1304]) );
  AND U9663 ( .A(p_input[1303]), .B(p_input[11303]), .Z(o[1303]) );
  AND U9664 ( .A(p_input[1302]), .B(p_input[11302]), .Z(o[1302]) );
  AND U9665 ( .A(p_input[1301]), .B(p_input[11301]), .Z(o[1301]) );
  AND U9666 ( .A(p_input[1300]), .B(p_input[11300]), .Z(o[1300]) );
  AND U9667 ( .A(p_input[12]), .B(p_input[10012]), .Z(o[12]) );
  AND U9668 ( .A(p_input[129]), .B(p_input[10129]), .Z(o[129]) );
  AND U9669 ( .A(p_input[1299]), .B(p_input[11299]), .Z(o[1299]) );
  AND U9670 ( .A(p_input[1298]), .B(p_input[11298]), .Z(o[1298]) );
  AND U9671 ( .A(p_input[1297]), .B(p_input[11297]), .Z(o[1297]) );
  AND U9672 ( .A(p_input[1296]), .B(p_input[11296]), .Z(o[1296]) );
  AND U9673 ( .A(p_input[1295]), .B(p_input[11295]), .Z(o[1295]) );
  AND U9674 ( .A(p_input[1294]), .B(p_input[11294]), .Z(o[1294]) );
  AND U9675 ( .A(p_input[1293]), .B(p_input[11293]), .Z(o[1293]) );
  AND U9676 ( .A(p_input[1292]), .B(p_input[11292]), .Z(o[1292]) );
  AND U9677 ( .A(p_input[1291]), .B(p_input[11291]), .Z(o[1291]) );
  AND U9678 ( .A(p_input[1290]), .B(p_input[11290]), .Z(o[1290]) );
  AND U9679 ( .A(p_input[128]), .B(p_input[10128]), .Z(o[128]) );
  AND U9680 ( .A(p_input[1289]), .B(p_input[11289]), .Z(o[1289]) );
  AND U9681 ( .A(p_input[1288]), .B(p_input[11288]), .Z(o[1288]) );
  AND U9682 ( .A(p_input[1287]), .B(p_input[11287]), .Z(o[1287]) );
  AND U9683 ( .A(p_input[1286]), .B(p_input[11286]), .Z(o[1286]) );
  AND U9684 ( .A(p_input[1285]), .B(p_input[11285]), .Z(o[1285]) );
  AND U9685 ( .A(p_input[1284]), .B(p_input[11284]), .Z(o[1284]) );
  AND U9686 ( .A(p_input[1283]), .B(p_input[11283]), .Z(o[1283]) );
  AND U9687 ( .A(p_input[1282]), .B(p_input[11282]), .Z(o[1282]) );
  AND U9688 ( .A(p_input[1281]), .B(p_input[11281]), .Z(o[1281]) );
  AND U9689 ( .A(p_input[1280]), .B(p_input[11280]), .Z(o[1280]) );
  AND U9690 ( .A(p_input[127]), .B(p_input[10127]), .Z(o[127]) );
  AND U9691 ( .A(p_input[1279]), .B(p_input[11279]), .Z(o[1279]) );
  AND U9692 ( .A(p_input[1278]), .B(p_input[11278]), .Z(o[1278]) );
  AND U9693 ( .A(p_input[1277]), .B(p_input[11277]), .Z(o[1277]) );
  AND U9694 ( .A(p_input[1276]), .B(p_input[11276]), .Z(o[1276]) );
  AND U9695 ( .A(p_input[1275]), .B(p_input[11275]), .Z(o[1275]) );
  AND U9696 ( .A(p_input[1274]), .B(p_input[11274]), .Z(o[1274]) );
  AND U9697 ( .A(p_input[1273]), .B(p_input[11273]), .Z(o[1273]) );
  AND U9698 ( .A(p_input[1272]), .B(p_input[11272]), .Z(o[1272]) );
  AND U9699 ( .A(p_input[1271]), .B(p_input[11271]), .Z(o[1271]) );
  AND U9700 ( .A(p_input[1270]), .B(p_input[11270]), .Z(o[1270]) );
  AND U9701 ( .A(p_input[126]), .B(p_input[10126]), .Z(o[126]) );
  AND U9702 ( .A(p_input[1269]), .B(p_input[11269]), .Z(o[1269]) );
  AND U9703 ( .A(p_input[1268]), .B(p_input[11268]), .Z(o[1268]) );
  AND U9704 ( .A(p_input[1267]), .B(p_input[11267]), .Z(o[1267]) );
  AND U9705 ( .A(p_input[1266]), .B(p_input[11266]), .Z(o[1266]) );
  AND U9706 ( .A(p_input[1265]), .B(p_input[11265]), .Z(o[1265]) );
  AND U9707 ( .A(p_input[1264]), .B(p_input[11264]), .Z(o[1264]) );
  AND U9708 ( .A(p_input[1263]), .B(p_input[11263]), .Z(o[1263]) );
  AND U9709 ( .A(p_input[1262]), .B(p_input[11262]), .Z(o[1262]) );
  AND U9710 ( .A(p_input[1261]), .B(p_input[11261]), .Z(o[1261]) );
  AND U9711 ( .A(p_input[1260]), .B(p_input[11260]), .Z(o[1260]) );
  AND U9712 ( .A(p_input[125]), .B(p_input[10125]), .Z(o[125]) );
  AND U9713 ( .A(p_input[1259]), .B(p_input[11259]), .Z(o[1259]) );
  AND U9714 ( .A(p_input[1258]), .B(p_input[11258]), .Z(o[1258]) );
  AND U9715 ( .A(p_input[1257]), .B(p_input[11257]), .Z(o[1257]) );
  AND U9716 ( .A(p_input[1256]), .B(p_input[11256]), .Z(o[1256]) );
  AND U9717 ( .A(p_input[1255]), .B(p_input[11255]), .Z(o[1255]) );
  AND U9718 ( .A(p_input[1254]), .B(p_input[11254]), .Z(o[1254]) );
  AND U9719 ( .A(p_input[1253]), .B(p_input[11253]), .Z(o[1253]) );
  AND U9720 ( .A(p_input[1252]), .B(p_input[11252]), .Z(o[1252]) );
  AND U9721 ( .A(p_input[1251]), .B(p_input[11251]), .Z(o[1251]) );
  AND U9722 ( .A(p_input[1250]), .B(p_input[11250]), .Z(o[1250]) );
  AND U9723 ( .A(p_input[124]), .B(p_input[10124]), .Z(o[124]) );
  AND U9724 ( .A(p_input[1249]), .B(p_input[11249]), .Z(o[1249]) );
  AND U9725 ( .A(p_input[1248]), .B(p_input[11248]), .Z(o[1248]) );
  AND U9726 ( .A(p_input[1247]), .B(p_input[11247]), .Z(o[1247]) );
  AND U9727 ( .A(p_input[1246]), .B(p_input[11246]), .Z(o[1246]) );
  AND U9728 ( .A(p_input[1245]), .B(p_input[11245]), .Z(o[1245]) );
  AND U9729 ( .A(p_input[1244]), .B(p_input[11244]), .Z(o[1244]) );
  AND U9730 ( .A(p_input[1243]), .B(p_input[11243]), .Z(o[1243]) );
  AND U9731 ( .A(p_input[1242]), .B(p_input[11242]), .Z(o[1242]) );
  AND U9732 ( .A(p_input[1241]), .B(p_input[11241]), .Z(o[1241]) );
  AND U9733 ( .A(p_input[1240]), .B(p_input[11240]), .Z(o[1240]) );
  AND U9734 ( .A(p_input[123]), .B(p_input[10123]), .Z(o[123]) );
  AND U9735 ( .A(p_input[1239]), .B(p_input[11239]), .Z(o[1239]) );
  AND U9736 ( .A(p_input[1238]), .B(p_input[11238]), .Z(o[1238]) );
  AND U9737 ( .A(p_input[1237]), .B(p_input[11237]), .Z(o[1237]) );
  AND U9738 ( .A(p_input[1236]), .B(p_input[11236]), .Z(o[1236]) );
  AND U9739 ( .A(p_input[1235]), .B(p_input[11235]), .Z(o[1235]) );
  AND U9740 ( .A(p_input[1234]), .B(p_input[11234]), .Z(o[1234]) );
  AND U9741 ( .A(p_input[1233]), .B(p_input[11233]), .Z(o[1233]) );
  AND U9742 ( .A(p_input[1232]), .B(p_input[11232]), .Z(o[1232]) );
  AND U9743 ( .A(p_input[1231]), .B(p_input[11231]), .Z(o[1231]) );
  AND U9744 ( .A(p_input[1230]), .B(p_input[11230]), .Z(o[1230]) );
  AND U9745 ( .A(p_input[122]), .B(p_input[10122]), .Z(o[122]) );
  AND U9746 ( .A(p_input[1229]), .B(p_input[11229]), .Z(o[1229]) );
  AND U9747 ( .A(p_input[1228]), .B(p_input[11228]), .Z(o[1228]) );
  AND U9748 ( .A(p_input[1227]), .B(p_input[11227]), .Z(o[1227]) );
  AND U9749 ( .A(p_input[1226]), .B(p_input[11226]), .Z(o[1226]) );
  AND U9750 ( .A(p_input[1225]), .B(p_input[11225]), .Z(o[1225]) );
  AND U9751 ( .A(p_input[1224]), .B(p_input[11224]), .Z(o[1224]) );
  AND U9752 ( .A(p_input[1223]), .B(p_input[11223]), .Z(o[1223]) );
  AND U9753 ( .A(p_input[1222]), .B(p_input[11222]), .Z(o[1222]) );
  AND U9754 ( .A(p_input[1221]), .B(p_input[11221]), .Z(o[1221]) );
  AND U9755 ( .A(p_input[1220]), .B(p_input[11220]), .Z(o[1220]) );
  AND U9756 ( .A(p_input[121]), .B(p_input[10121]), .Z(o[121]) );
  AND U9757 ( .A(p_input[1219]), .B(p_input[11219]), .Z(o[1219]) );
  AND U9758 ( .A(p_input[1218]), .B(p_input[11218]), .Z(o[1218]) );
  AND U9759 ( .A(p_input[1217]), .B(p_input[11217]), .Z(o[1217]) );
  AND U9760 ( .A(p_input[1216]), .B(p_input[11216]), .Z(o[1216]) );
  AND U9761 ( .A(p_input[1215]), .B(p_input[11215]), .Z(o[1215]) );
  AND U9762 ( .A(p_input[1214]), .B(p_input[11214]), .Z(o[1214]) );
  AND U9763 ( .A(p_input[1213]), .B(p_input[11213]), .Z(o[1213]) );
  AND U9764 ( .A(p_input[1212]), .B(p_input[11212]), .Z(o[1212]) );
  AND U9765 ( .A(p_input[1211]), .B(p_input[11211]), .Z(o[1211]) );
  AND U9766 ( .A(p_input[1210]), .B(p_input[11210]), .Z(o[1210]) );
  AND U9767 ( .A(p_input[120]), .B(p_input[10120]), .Z(o[120]) );
  AND U9768 ( .A(p_input[1209]), .B(p_input[11209]), .Z(o[1209]) );
  AND U9769 ( .A(p_input[1208]), .B(p_input[11208]), .Z(o[1208]) );
  AND U9770 ( .A(p_input[1207]), .B(p_input[11207]), .Z(o[1207]) );
  AND U9771 ( .A(p_input[1206]), .B(p_input[11206]), .Z(o[1206]) );
  AND U9772 ( .A(p_input[1205]), .B(p_input[11205]), .Z(o[1205]) );
  AND U9773 ( .A(p_input[1204]), .B(p_input[11204]), .Z(o[1204]) );
  AND U9774 ( .A(p_input[1203]), .B(p_input[11203]), .Z(o[1203]) );
  AND U9775 ( .A(p_input[1202]), .B(p_input[11202]), .Z(o[1202]) );
  AND U9776 ( .A(p_input[1201]), .B(p_input[11201]), .Z(o[1201]) );
  AND U9777 ( .A(p_input[1200]), .B(p_input[11200]), .Z(o[1200]) );
  AND U9778 ( .A(p_input[11]), .B(p_input[10011]), .Z(o[11]) );
  AND U9779 ( .A(p_input[119]), .B(p_input[10119]), .Z(o[119]) );
  AND U9780 ( .A(p_input[1199]), .B(p_input[11199]), .Z(o[1199]) );
  AND U9781 ( .A(p_input[1198]), .B(p_input[11198]), .Z(o[1198]) );
  AND U9782 ( .A(p_input[1197]), .B(p_input[11197]), .Z(o[1197]) );
  AND U9783 ( .A(p_input[1196]), .B(p_input[11196]), .Z(o[1196]) );
  AND U9784 ( .A(p_input[1195]), .B(p_input[11195]), .Z(o[1195]) );
  AND U9785 ( .A(p_input[1194]), .B(p_input[11194]), .Z(o[1194]) );
  AND U9786 ( .A(p_input[1193]), .B(p_input[11193]), .Z(o[1193]) );
  AND U9787 ( .A(p_input[1192]), .B(p_input[11192]), .Z(o[1192]) );
  AND U9788 ( .A(p_input[1191]), .B(p_input[11191]), .Z(o[1191]) );
  AND U9789 ( .A(p_input[1190]), .B(p_input[11190]), .Z(o[1190]) );
  AND U9790 ( .A(p_input[118]), .B(p_input[10118]), .Z(o[118]) );
  AND U9791 ( .A(p_input[1189]), .B(p_input[11189]), .Z(o[1189]) );
  AND U9792 ( .A(p_input[1188]), .B(p_input[11188]), .Z(o[1188]) );
  AND U9793 ( .A(p_input[1187]), .B(p_input[11187]), .Z(o[1187]) );
  AND U9794 ( .A(p_input[1186]), .B(p_input[11186]), .Z(o[1186]) );
  AND U9795 ( .A(p_input[1185]), .B(p_input[11185]), .Z(o[1185]) );
  AND U9796 ( .A(p_input[1184]), .B(p_input[11184]), .Z(o[1184]) );
  AND U9797 ( .A(p_input[1183]), .B(p_input[11183]), .Z(o[1183]) );
  AND U9798 ( .A(p_input[1182]), .B(p_input[11182]), .Z(o[1182]) );
  AND U9799 ( .A(p_input[1181]), .B(p_input[11181]), .Z(o[1181]) );
  AND U9800 ( .A(p_input[1180]), .B(p_input[11180]), .Z(o[1180]) );
  AND U9801 ( .A(p_input[117]), .B(p_input[10117]), .Z(o[117]) );
  AND U9802 ( .A(p_input[1179]), .B(p_input[11179]), .Z(o[1179]) );
  AND U9803 ( .A(p_input[1178]), .B(p_input[11178]), .Z(o[1178]) );
  AND U9804 ( .A(p_input[1177]), .B(p_input[11177]), .Z(o[1177]) );
  AND U9805 ( .A(p_input[1176]), .B(p_input[11176]), .Z(o[1176]) );
  AND U9806 ( .A(p_input[1175]), .B(p_input[11175]), .Z(o[1175]) );
  AND U9807 ( .A(p_input[1174]), .B(p_input[11174]), .Z(o[1174]) );
  AND U9808 ( .A(p_input[1173]), .B(p_input[11173]), .Z(o[1173]) );
  AND U9809 ( .A(p_input[1172]), .B(p_input[11172]), .Z(o[1172]) );
  AND U9810 ( .A(p_input[1171]), .B(p_input[11171]), .Z(o[1171]) );
  AND U9811 ( .A(p_input[1170]), .B(p_input[11170]), .Z(o[1170]) );
  AND U9812 ( .A(p_input[116]), .B(p_input[10116]), .Z(o[116]) );
  AND U9813 ( .A(p_input[1169]), .B(p_input[11169]), .Z(o[1169]) );
  AND U9814 ( .A(p_input[1168]), .B(p_input[11168]), .Z(o[1168]) );
  AND U9815 ( .A(p_input[1167]), .B(p_input[11167]), .Z(o[1167]) );
  AND U9816 ( .A(p_input[1166]), .B(p_input[11166]), .Z(o[1166]) );
  AND U9817 ( .A(p_input[1165]), .B(p_input[11165]), .Z(o[1165]) );
  AND U9818 ( .A(p_input[1164]), .B(p_input[11164]), .Z(o[1164]) );
  AND U9819 ( .A(p_input[1163]), .B(p_input[11163]), .Z(o[1163]) );
  AND U9820 ( .A(p_input[1162]), .B(p_input[11162]), .Z(o[1162]) );
  AND U9821 ( .A(p_input[1161]), .B(p_input[11161]), .Z(o[1161]) );
  AND U9822 ( .A(p_input[1160]), .B(p_input[11160]), .Z(o[1160]) );
  AND U9823 ( .A(p_input[115]), .B(p_input[10115]), .Z(o[115]) );
  AND U9824 ( .A(p_input[1159]), .B(p_input[11159]), .Z(o[1159]) );
  AND U9825 ( .A(p_input[1158]), .B(p_input[11158]), .Z(o[1158]) );
  AND U9826 ( .A(p_input[1157]), .B(p_input[11157]), .Z(o[1157]) );
  AND U9827 ( .A(p_input[1156]), .B(p_input[11156]), .Z(o[1156]) );
  AND U9828 ( .A(p_input[1155]), .B(p_input[11155]), .Z(o[1155]) );
  AND U9829 ( .A(p_input[1154]), .B(p_input[11154]), .Z(o[1154]) );
  AND U9830 ( .A(p_input[1153]), .B(p_input[11153]), .Z(o[1153]) );
  AND U9831 ( .A(p_input[1152]), .B(p_input[11152]), .Z(o[1152]) );
  AND U9832 ( .A(p_input[1151]), .B(p_input[11151]), .Z(o[1151]) );
  AND U9833 ( .A(p_input[1150]), .B(p_input[11150]), .Z(o[1150]) );
  AND U9834 ( .A(p_input[114]), .B(p_input[10114]), .Z(o[114]) );
  AND U9835 ( .A(p_input[1149]), .B(p_input[11149]), .Z(o[1149]) );
  AND U9836 ( .A(p_input[1148]), .B(p_input[11148]), .Z(o[1148]) );
  AND U9837 ( .A(p_input[1147]), .B(p_input[11147]), .Z(o[1147]) );
  AND U9838 ( .A(p_input[1146]), .B(p_input[11146]), .Z(o[1146]) );
  AND U9839 ( .A(p_input[1145]), .B(p_input[11145]), .Z(o[1145]) );
  AND U9840 ( .A(p_input[1144]), .B(p_input[11144]), .Z(o[1144]) );
  AND U9841 ( .A(p_input[1143]), .B(p_input[11143]), .Z(o[1143]) );
  AND U9842 ( .A(p_input[1142]), .B(p_input[11142]), .Z(o[1142]) );
  AND U9843 ( .A(p_input[1141]), .B(p_input[11141]), .Z(o[1141]) );
  AND U9844 ( .A(p_input[1140]), .B(p_input[11140]), .Z(o[1140]) );
  AND U9845 ( .A(p_input[113]), .B(p_input[10113]), .Z(o[113]) );
  AND U9846 ( .A(p_input[1139]), .B(p_input[11139]), .Z(o[1139]) );
  AND U9847 ( .A(p_input[1138]), .B(p_input[11138]), .Z(o[1138]) );
  AND U9848 ( .A(p_input[1137]), .B(p_input[11137]), .Z(o[1137]) );
  AND U9849 ( .A(p_input[1136]), .B(p_input[11136]), .Z(o[1136]) );
  AND U9850 ( .A(p_input[1135]), .B(p_input[11135]), .Z(o[1135]) );
  AND U9851 ( .A(p_input[1134]), .B(p_input[11134]), .Z(o[1134]) );
  AND U9852 ( .A(p_input[1133]), .B(p_input[11133]), .Z(o[1133]) );
  AND U9853 ( .A(p_input[1132]), .B(p_input[11132]), .Z(o[1132]) );
  AND U9854 ( .A(p_input[1131]), .B(p_input[11131]), .Z(o[1131]) );
  AND U9855 ( .A(p_input[1130]), .B(p_input[11130]), .Z(o[1130]) );
  AND U9856 ( .A(p_input[112]), .B(p_input[10112]), .Z(o[112]) );
  AND U9857 ( .A(p_input[1129]), .B(p_input[11129]), .Z(o[1129]) );
  AND U9858 ( .A(p_input[1128]), .B(p_input[11128]), .Z(o[1128]) );
  AND U9859 ( .A(p_input[1127]), .B(p_input[11127]), .Z(o[1127]) );
  AND U9860 ( .A(p_input[1126]), .B(p_input[11126]), .Z(o[1126]) );
  AND U9861 ( .A(p_input[1125]), .B(p_input[11125]), .Z(o[1125]) );
  AND U9862 ( .A(p_input[1124]), .B(p_input[11124]), .Z(o[1124]) );
  AND U9863 ( .A(p_input[1123]), .B(p_input[11123]), .Z(o[1123]) );
  AND U9864 ( .A(p_input[1122]), .B(p_input[11122]), .Z(o[1122]) );
  AND U9865 ( .A(p_input[1121]), .B(p_input[11121]), .Z(o[1121]) );
  AND U9866 ( .A(p_input[1120]), .B(p_input[11120]), .Z(o[1120]) );
  AND U9867 ( .A(p_input[111]), .B(p_input[10111]), .Z(o[111]) );
  AND U9868 ( .A(p_input[1119]), .B(p_input[11119]), .Z(o[1119]) );
  AND U9869 ( .A(p_input[1118]), .B(p_input[11118]), .Z(o[1118]) );
  AND U9870 ( .A(p_input[1117]), .B(p_input[11117]), .Z(o[1117]) );
  AND U9871 ( .A(p_input[1116]), .B(p_input[11116]), .Z(o[1116]) );
  AND U9872 ( .A(p_input[1115]), .B(p_input[11115]), .Z(o[1115]) );
  AND U9873 ( .A(p_input[1114]), .B(p_input[11114]), .Z(o[1114]) );
  AND U9874 ( .A(p_input[1113]), .B(p_input[11113]), .Z(o[1113]) );
  AND U9875 ( .A(p_input[1112]), .B(p_input[11112]), .Z(o[1112]) );
  AND U9876 ( .A(p_input[1111]), .B(p_input[11111]), .Z(o[1111]) );
  AND U9877 ( .A(p_input[11110]), .B(p_input[1110]), .Z(o[1110]) );
  AND U9878 ( .A(p_input[110]), .B(p_input[10110]), .Z(o[110]) );
  AND U9879 ( .A(p_input[11109]), .B(p_input[1109]), .Z(o[1109]) );
  AND U9880 ( .A(p_input[11108]), .B(p_input[1108]), .Z(o[1108]) );
  AND U9881 ( .A(p_input[11107]), .B(p_input[1107]), .Z(o[1107]) );
  AND U9882 ( .A(p_input[11106]), .B(p_input[1106]), .Z(o[1106]) );
  AND U9883 ( .A(p_input[11105]), .B(p_input[1105]), .Z(o[1105]) );
  AND U9884 ( .A(p_input[11104]), .B(p_input[1104]), .Z(o[1104]) );
  AND U9885 ( .A(p_input[11103]), .B(p_input[1103]), .Z(o[1103]) );
  AND U9886 ( .A(p_input[11102]), .B(p_input[1102]), .Z(o[1102]) );
  AND U9887 ( .A(p_input[11101]), .B(p_input[1101]), .Z(o[1101]) );
  AND U9888 ( .A(p_input[11100]), .B(p_input[1100]), .Z(o[1100]) );
  AND U9889 ( .A(p_input[10]), .B(p_input[10010]), .Z(o[10]) );
  AND U9890 ( .A(p_input[109]), .B(p_input[10109]), .Z(o[109]) );
  AND U9891 ( .A(p_input[11099]), .B(p_input[1099]), .Z(o[1099]) );
  AND U9892 ( .A(p_input[11098]), .B(p_input[1098]), .Z(o[1098]) );
  AND U9893 ( .A(p_input[11097]), .B(p_input[1097]), .Z(o[1097]) );
  AND U9894 ( .A(p_input[11096]), .B(p_input[1096]), .Z(o[1096]) );
  AND U9895 ( .A(p_input[11095]), .B(p_input[1095]), .Z(o[1095]) );
  AND U9896 ( .A(p_input[11094]), .B(p_input[1094]), .Z(o[1094]) );
  AND U9897 ( .A(p_input[11093]), .B(p_input[1093]), .Z(o[1093]) );
  AND U9898 ( .A(p_input[11092]), .B(p_input[1092]), .Z(o[1092]) );
  AND U9899 ( .A(p_input[11091]), .B(p_input[1091]), .Z(o[1091]) );
  AND U9900 ( .A(p_input[11090]), .B(p_input[1090]), .Z(o[1090]) );
  AND U9901 ( .A(p_input[108]), .B(p_input[10108]), .Z(o[108]) );
  AND U9902 ( .A(p_input[11089]), .B(p_input[1089]), .Z(o[1089]) );
  AND U9903 ( .A(p_input[11088]), .B(p_input[1088]), .Z(o[1088]) );
  AND U9904 ( .A(p_input[11087]), .B(p_input[1087]), .Z(o[1087]) );
  AND U9905 ( .A(p_input[11086]), .B(p_input[1086]), .Z(o[1086]) );
  AND U9906 ( .A(p_input[11085]), .B(p_input[1085]), .Z(o[1085]) );
  AND U9907 ( .A(p_input[11084]), .B(p_input[1084]), .Z(o[1084]) );
  AND U9908 ( .A(p_input[11083]), .B(p_input[1083]), .Z(o[1083]) );
  AND U9909 ( .A(p_input[11082]), .B(p_input[1082]), .Z(o[1082]) );
  AND U9910 ( .A(p_input[11081]), .B(p_input[1081]), .Z(o[1081]) );
  AND U9911 ( .A(p_input[11080]), .B(p_input[1080]), .Z(o[1080]) );
  AND U9912 ( .A(p_input[107]), .B(p_input[10107]), .Z(o[107]) );
  AND U9913 ( .A(p_input[11079]), .B(p_input[1079]), .Z(o[1079]) );
  AND U9914 ( .A(p_input[11078]), .B(p_input[1078]), .Z(o[1078]) );
  AND U9915 ( .A(p_input[11077]), .B(p_input[1077]), .Z(o[1077]) );
  AND U9916 ( .A(p_input[11076]), .B(p_input[1076]), .Z(o[1076]) );
  AND U9917 ( .A(p_input[11075]), .B(p_input[1075]), .Z(o[1075]) );
  AND U9918 ( .A(p_input[11074]), .B(p_input[1074]), .Z(o[1074]) );
  AND U9919 ( .A(p_input[11073]), .B(p_input[1073]), .Z(o[1073]) );
  AND U9920 ( .A(p_input[11072]), .B(p_input[1072]), .Z(o[1072]) );
  AND U9921 ( .A(p_input[11071]), .B(p_input[1071]), .Z(o[1071]) );
  AND U9922 ( .A(p_input[11070]), .B(p_input[1070]), .Z(o[1070]) );
  AND U9923 ( .A(p_input[106]), .B(p_input[10106]), .Z(o[106]) );
  AND U9924 ( .A(p_input[11069]), .B(p_input[1069]), .Z(o[1069]) );
  AND U9925 ( .A(p_input[11068]), .B(p_input[1068]), .Z(o[1068]) );
  AND U9926 ( .A(p_input[11067]), .B(p_input[1067]), .Z(o[1067]) );
  AND U9927 ( .A(p_input[11066]), .B(p_input[1066]), .Z(o[1066]) );
  AND U9928 ( .A(p_input[11065]), .B(p_input[1065]), .Z(o[1065]) );
  AND U9929 ( .A(p_input[11064]), .B(p_input[1064]), .Z(o[1064]) );
  AND U9930 ( .A(p_input[11063]), .B(p_input[1063]), .Z(o[1063]) );
  AND U9931 ( .A(p_input[11062]), .B(p_input[1062]), .Z(o[1062]) );
  AND U9932 ( .A(p_input[11061]), .B(p_input[1061]), .Z(o[1061]) );
  AND U9933 ( .A(p_input[11060]), .B(p_input[1060]), .Z(o[1060]) );
  AND U9934 ( .A(p_input[105]), .B(p_input[10105]), .Z(o[105]) );
  AND U9935 ( .A(p_input[11059]), .B(p_input[1059]), .Z(o[1059]) );
  AND U9936 ( .A(p_input[11058]), .B(p_input[1058]), .Z(o[1058]) );
  AND U9937 ( .A(p_input[11057]), .B(p_input[1057]), .Z(o[1057]) );
  AND U9938 ( .A(p_input[11056]), .B(p_input[1056]), .Z(o[1056]) );
  AND U9939 ( .A(p_input[11055]), .B(p_input[1055]), .Z(o[1055]) );
  AND U9940 ( .A(p_input[11054]), .B(p_input[1054]), .Z(o[1054]) );
  AND U9941 ( .A(p_input[11053]), .B(p_input[1053]), .Z(o[1053]) );
  AND U9942 ( .A(p_input[11052]), .B(p_input[1052]), .Z(o[1052]) );
  AND U9943 ( .A(p_input[11051]), .B(p_input[1051]), .Z(o[1051]) );
  AND U9944 ( .A(p_input[11050]), .B(p_input[1050]), .Z(o[1050]) );
  AND U9945 ( .A(p_input[104]), .B(p_input[10104]), .Z(o[104]) );
  AND U9946 ( .A(p_input[11049]), .B(p_input[1049]), .Z(o[1049]) );
  AND U9947 ( .A(p_input[11048]), .B(p_input[1048]), .Z(o[1048]) );
  AND U9948 ( .A(p_input[11047]), .B(p_input[1047]), .Z(o[1047]) );
  AND U9949 ( .A(p_input[11046]), .B(p_input[1046]), .Z(o[1046]) );
  AND U9950 ( .A(p_input[11045]), .B(p_input[1045]), .Z(o[1045]) );
  AND U9951 ( .A(p_input[11044]), .B(p_input[1044]), .Z(o[1044]) );
  AND U9952 ( .A(p_input[11043]), .B(p_input[1043]), .Z(o[1043]) );
  AND U9953 ( .A(p_input[11042]), .B(p_input[1042]), .Z(o[1042]) );
  AND U9954 ( .A(p_input[11041]), .B(p_input[1041]), .Z(o[1041]) );
  AND U9955 ( .A(p_input[11040]), .B(p_input[1040]), .Z(o[1040]) );
  AND U9956 ( .A(p_input[103]), .B(p_input[10103]), .Z(o[103]) );
  AND U9957 ( .A(p_input[11039]), .B(p_input[1039]), .Z(o[1039]) );
  AND U9958 ( .A(p_input[11038]), .B(p_input[1038]), .Z(o[1038]) );
  AND U9959 ( .A(p_input[11037]), .B(p_input[1037]), .Z(o[1037]) );
  AND U9960 ( .A(p_input[11036]), .B(p_input[1036]), .Z(o[1036]) );
  AND U9961 ( .A(p_input[11035]), .B(p_input[1035]), .Z(o[1035]) );
  AND U9962 ( .A(p_input[11034]), .B(p_input[1034]), .Z(o[1034]) );
  AND U9963 ( .A(p_input[11033]), .B(p_input[1033]), .Z(o[1033]) );
  AND U9964 ( .A(p_input[11032]), .B(p_input[1032]), .Z(o[1032]) );
  AND U9965 ( .A(p_input[11031]), .B(p_input[1031]), .Z(o[1031]) );
  AND U9966 ( .A(p_input[11030]), .B(p_input[1030]), .Z(o[1030]) );
  AND U9967 ( .A(p_input[102]), .B(p_input[10102]), .Z(o[102]) );
  AND U9968 ( .A(p_input[11029]), .B(p_input[1029]), .Z(o[1029]) );
  AND U9969 ( .A(p_input[11028]), .B(p_input[1028]), .Z(o[1028]) );
  AND U9970 ( .A(p_input[11027]), .B(p_input[1027]), .Z(o[1027]) );
  AND U9971 ( .A(p_input[11026]), .B(p_input[1026]), .Z(o[1026]) );
  AND U9972 ( .A(p_input[11025]), .B(p_input[1025]), .Z(o[1025]) );
  AND U9973 ( .A(p_input[11024]), .B(p_input[1024]), .Z(o[1024]) );
  AND U9974 ( .A(p_input[11023]), .B(p_input[1023]), .Z(o[1023]) );
  AND U9975 ( .A(p_input[11022]), .B(p_input[1022]), .Z(o[1022]) );
  AND U9976 ( .A(p_input[11021]), .B(p_input[1021]), .Z(o[1021]) );
  AND U9977 ( .A(p_input[11020]), .B(p_input[1020]), .Z(o[1020]) );
  AND U9978 ( .A(p_input[101]), .B(p_input[10101]), .Z(o[101]) );
  AND U9979 ( .A(p_input[11019]), .B(p_input[1019]), .Z(o[1019]) );
  AND U9980 ( .A(p_input[11018]), .B(p_input[1018]), .Z(o[1018]) );
  AND U9981 ( .A(p_input[11017]), .B(p_input[1017]), .Z(o[1017]) );
  AND U9982 ( .A(p_input[11016]), .B(p_input[1016]), .Z(o[1016]) );
  AND U9983 ( .A(p_input[11015]), .B(p_input[1015]), .Z(o[1015]) );
  AND U9984 ( .A(p_input[11014]), .B(p_input[1014]), .Z(o[1014]) );
  AND U9985 ( .A(p_input[11013]), .B(p_input[1013]), .Z(o[1013]) );
  AND U9986 ( .A(p_input[11012]), .B(p_input[1012]), .Z(o[1012]) );
  AND U9987 ( .A(p_input[11011]), .B(p_input[1011]), .Z(o[1011]) );
  AND U9988 ( .A(p_input[11010]), .B(p_input[1010]), .Z(o[1010]) );
  AND U9989 ( .A(p_input[10100]), .B(p_input[100]), .Z(o[100]) );
  AND U9990 ( .A(p_input[11009]), .B(p_input[1009]), .Z(o[1009]) );
  AND U9991 ( .A(p_input[11008]), .B(p_input[1008]), .Z(o[1008]) );
  AND U9992 ( .A(p_input[11007]), .B(p_input[1007]), .Z(o[1007]) );
  AND U9993 ( .A(p_input[11006]), .B(p_input[1006]), .Z(o[1006]) );
  AND U9994 ( .A(p_input[11005]), .B(p_input[1005]), .Z(o[1005]) );
  AND U9995 ( .A(p_input[11004]), .B(p_input[1004]), .Z(o[1004]) );
  AND U9996 ( .A(p_input[11003]), .B(p_input[1003]), .Z(o[1003]) );
  AND U9997 ( .A(p_input[11002]), .B(p_input[1002]), .Z(o[1002]) );
  AND U9998 ( .A(p_input[11001]), .B(p_input[1001]), .Z(o[1001]) );
  AND U9999 ( .A(p_input[11000]), .B(p_input[1000]), .Z(o[1000]) );
  AND U10000 ( .A(p_input[10000]), .B(p_input[0]), .Z(o[0]) );
endmodule

