
module knn_comb_BMR_W32_K1_N8 ( p_input, o );
  input [287:0] p_input;
  output [31:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/min_val_out[0][16] , \knn_comb_/min_val_out[0][17] ,
         \knn_comb_/min_val_out[0][18] , \knn_comb_/min_val_out[0][19] ,
         \knn_comb_/min_val_out[0][20] , \knn_comb_/min_val_out[0][21] ,
         \knn_comb_/min_val_out[0][22] , \knn_comb_/min_val_out[0][23] ,
         \knn_comb_/min_val_out[0][24] , \knn_comb_/min_val_out[0][25] ,
         \knn_comb_/min_val_out[0][26] , \knn_comb_/min_val_out[0][27] ,
         \knn_comb_/min_val_out[0][28] , \knn_comb_/min_val_out[0][29] ,
         \knn_comb_/min_val_out[0][30] , \knn_comb_/min_val_out[0][31] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313;
  assign \knn_comb_/min_val_out[0][0]  = p_input[224];
  assign \knn_comb_/min_val_out[0][1]  = p_input[225];
  assign \knn_comb_/min_val_out[0][2]  = p_input[226];
  assign \knn_comb_/min_val_out[0][3]  = p_input[227];
  assign \knn_comb_/min_val_out[0][4]  = p_input[228];
  assign \knn_comb_/min_val_out[0][5]  = p_input[229];
  assign \knn_comb_/min_val_out[0][6]  = p_input[230];
  assign \knn_comb_/min_val_out[0][7]  = p_input[231];
  assign \knn_comb_/min_val_out[0][8]  = p_input[232];
  assign \knn_comb_/min_val_out[0][9]  = p_input[233];
  assign \knn_comb_/min_val_out[0][10]  = p_input[234];
  assign \knn_comb_/min_val_out[0][11]  = p_input[235];
  assign \knn_comb_/min_val_out[0][12]  = p_input[236];
  assign \knn_comb_/min_val_out[0][13]  = p_input[237];
  assign \knn_comb_/min_val_out[0][14]  = p_input[238];
  assign \knn_comb_/min_val_out[0][15]  = p_input[239];
  assign \knn_comb_/min_val_out[0][16]  = p_input[240];
  assign \knn_comb_/min_val_out[0][17]  = p_input[241];
  assign \knn_comb_/min_val_out[0][18]  = p_input[242];
  assign \knn_comb_/min_val_out[0][19]  = p_input[243];
  assign \knn_comb_/min_val_out[0][20]  = p_input[244];
  assign \knn_comb_/min_val_out[0][21]  = p_input[245];
  assign \knn_comb_/min_val_out[0][22]  = p_input[246];
  assign \knn_comb_/min_val_out[0][23]  = p_input[247];
  assign \knn_comb_/min_val_out[0][24]  = p_input[248];
  assign \knn_comb_/min_val_out[0][25]  = p_input[249];
  assign \knn_comb_/min_val_out[0][26]  = p_input[250];
  assign \knn_comb_/min_val_out[0][27]  = p_input[251];
  assign \knn_comb_/min_val_out[0][28]  = p_input[252];
  assign \knn_comb_/min_val_out[0][29]  = p_input[253];
  assign \knn_comb_/min_val_out[0][30]  = p_input[254];
  assign \knn_comb_/min_val_out[0][31]  = p_input[255];

  XNOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(n3), .B(n4), .Z(n1) );
  XNOR U3 ( .A(p_input[9]), .B(n2), .Z(n4) );
  XOR U4 ( .A(n5), .B(n6), .Z(n2) );
  AND U5 ( .A(n7), .B(n8), .Z(n6) );
  XNOR U6 ( .A(p_input[41]), .B(n5), .Z(n8) );
  XOR U7 ( .A(n9), .B(n10), .Z(n5) );
  AND U8 ( .A(n11), .B(n12), .Z(n10) );
  XNOR U9 ( .A(p_input[73]), .B(n9), .Z(n12) );
  XOR U10 ( .A(n13), .B(n14), .Z(n9) );
  AND U11 ( .A(n15), .B(n16), .Z(n14) );
  XNOR U12 ( .A(p_input[105]), .B(n13), .Z(n16) );
  XOR U13 ( .A(n17), .B(n18), .Z(n13) );
  AND U14 ( .A(n19), .B(n20), .Z(n18) );
  XNOR U15 ( .A(p_input[137]), .B(n17), .Z(n20) );
  XNOR U16 ( .A(n21), .B(n22), .Z(n17) );
  AND U17 ( .A(n23), .B(n24), .Z(n22) );
  XOR U18 ( .A(p_input[169]), .B(n21), .Z(n24) );
  XOR U19 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n25), .Z(n21) );
  AND U20 ( .A(n26), .B(n27), .Z(n25) );
  XOR U21 ( .A(p_input[201]), .B(\knn_comb_/min_val_out[0][9] ), .Z(n27) );
  XNOR U22 ( .A(n28), .B(n29), .Z(o[8]) );
  AND U23 ( .A(n3), .B(n30), .Z(n28) );
  XNOR U24 ( .A(p_input[8]), .B(n29), .Z(n30) );
  XOR U25 ( .A(n31), .B(n32), .Z(n29) );
  AND U26 ( .A(n7), .B(n33), .Z(n32) );
  XNOR U27 ( .A(p_input[40]), .B(n31), .Z(n33) );
  XOR U28 ( .A(n34), .B(n35), .Z(n31) );
  AND U29 ( .A(n11), .B(n36), .Z(n35) );
  XNOR U30 ( .A(p_input[72]), .B(n34), .Z(n36) );
  XOR U31 ( .A(n37), .B(n38), .Z(n34) );
  AND U32 ( .A(n15), .B(n39), .Z(n38) );
  XNOR U33 ( .A(p_input[104]), .B(n37), .Z(n39) );
  XOR U34 ( .A(n40), .B(n41), .Z(n37) );
  AND U35 ( .A(n19), .B(n42), .Z(n41) );
  XNOR U36 ( .A(p_input[136]), .B(n40), .Z(n42) );
  XNOR U37 ( .A(n43), .B(n44), .Z(n40) );
  AND U38 ( .A(n23), .B(n45), .Z(n44) );
  XOR U39 ( .A(p_input[168]), .B(n43), .Z(n45) );
  XOR U40 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n46), .Z(n43) );
  AND U41 ( .A(n26), .B(n47), .Z(n46) );
  XOR U42 ( .A(p_input[200]), .B(\knn_comb_/min_val_out[0][8] ), .Z(n47) );
  XNOR U43 ( .A(n48), .B(n49), .Z(o[7]) );
  AND U44 ( .A(n3), .B(n50), .Z(n48) );
  XNOR U45 ( .A(p_input[7]), .B(n49), .Z(n50) );
  XOR U46 ( .A(n51), .B(n52), .Z(n49) );
  AND U47 ( .A(n7), .B(n53), .Z(n52) );
  XNOR U48 ( .A(p_input[39]), .B(n51), .Z(n53) );
  XOR U49 ( .A(n54), .B(n55), .Z(n51) );
  AND U50 ( .A(n11), .B(n56), .Z(n55) );
  XNOR U51 ( .A(p_input[71]), .B(n54), .Z(n56) );
  XOR U52 ( .A(n57), .B(n58), .Z(n54) );
  AND U53 ( .A(n15), .B(n59), .Z(n58) );
  XNOR U54 ( .A(p_input[103]), .B(n57), .Z(n59) );
  XOR U55 ( .A(n60), .B(n61), .Z(n57) );
  AND U56 ( .A(n19), .B(n62), .Z(n61) );
  XNOR U57 ( .A(p_input[135]), .B(n60), .Z(n62) );
  XNOR U58 ( .A(n63), .B(n64), .Z(n60) );
  AND U59 ( .A(n23), .B(n65), .Z(n64) );
  XOR U60 ( .A(p_input[167]), .B(n63), .Z(n65) );
  XOR U61 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n66), .Z(n63) );
  AND U62 ( .A(n26), .B(n67), .Z(n66) );
  XOR U63 ( .A(p_input[199]), .B(\knn_comb_/min_val_out[0][7] ), .Z(n67) );
  XNOR U64 ( .A(n68), .B(n69), .Z(o[6]) );
  AND U65 ( .A(n3), .B(n70), .Z(n68) );
  XNOR U66 ( .A(p_input[6]), .B(n69), .Z(n70) );
  XOR U67 ( .A(n71), .B(n72), .Z(n69) );
  AND U68 ( .A(n7), .B(n73), .Z(n72) );
  XNOR U69 ( .A(p_input[38]), .B(n71), .Z(n73) );
  XOR U70 ( .A(n74), .B(n75), .Z(n71) );
  AND U71 ( .A(n11), .B(n76), .Z(n75) );
  XNOR U72 ( .A(p_input[70]), .B(n74), .Z(n76) );
  XOR U73 ( .A(n77), .B(n78), .Z(n74) );
  AND U74 ( .A(n15), .B(n79), .Z(n78) );
  XNOR U75 ( .A(p_input[102]), .B(n77), .Z(n79) );
  XOR U76 ( .A(n80), .B(n81), .Z(n77) );
  AND U77 ( .A(n19), .B(n82), .Z(n81) );
  XNOR U78 ( .A(p_input[134]), .B(n80), .Z(n82) );
  XNOR U79 ( .A(n83), .B(n84), .Z(n80) );
  AND U80 ( .A(n23), .B(n85), .Z(n84) );
  XOR U81 ( .A(p_input[166]), .B(n83), .Z(n85) );
  XOR U82 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n86), .Z(n83) );
  AND U83 ( .A(n26), .B(n87), .Z(n86) );
  XOR U84 ( .A(p_input[198]), .B(\knn_comb_/min_val_out[0][6] ), .Z(n87) );
  XNOR U85 ( .A(n88), .B(n89), .Z(o[5]) );
  AND U86 ( .A(n3), .B(n90), .Z(n88) );
  XNOR U87 ( .A(p_input[5]), .B(n89), .Z(n90) );
  XOR U88 ( .A(n91), .B(n92), .Z(n89) );
  AND U89 ( .A(n7), .B(n93), .Z(n92) );
  XNOR U90 ( .A(p_input[37]), .B(n91), .Z(n93) );
  XOR U91 ( .A(n94), .B(n95), .Z(n91) );
  AND U92 ( .A(n11), .B(n96), .Z(n95) );
  XNOR U93 ( .A(p_input[69]), .B(n94), .Z(n96) );
  XOR U94 ( .A(n97), .B(n98), .Z(n94) );
  AND U95 ( .A(n15), .B(n99), .Z(n98) );
  XNOR U96 ( .A(p_input[101]), .B(n97), .Z(n99) );
  XOR U97 ( .A(n100), .B(n101), .Z(n97) );
  AND U98 ( .A(n19), .B(n102), .Z(n101) );
  XNOR U99 ( .A(p_input[133]), .B(n100), .Z(n102) );
  XNOR U100 ( .A(n103), .B(n104), .Z(n100) );
  AND U101 ( .A(n23), .B(n105), .Z(n104) );
  XOR U102 ( .A(p_input[165]), .B(n103), .Z(n105) );
  XOR U103 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n106), .Z(n103) );
  AND U104 ( .A(n26), .B(n107), .Z(n106) );
  XOR U105 ( .A(p_input[197]), .B(\knn_comb_/min_val_out[0][5] ), .Z(n107) );
  XNOR U106 ( .A(n108), .B(n109), .Z(o[4]) );
  AND U107 ( .A(n3), .B(n110), .Z(n108) );
  XNOR U108 ( .A(p_input[4]), .B(n109), .Z(n110) );
  XOR U109 ( .A(n111), .B(n112), .Z(n109) );
  AND U110 ( .A(n7), .B(n113), .Z(n112) );
  XNOR U111 ( .A(p_input[36]), .B(n111), .Z(n113) );
  XOR U112 ( .A(n114), .B(n115), .Z(n111) );
  AND U113 ( .A(n11), .B(n116), .Z(n115) );
  XNOR U114 ( .A(p_input[68]), .B(n114), .Z(n116) );
  XOR U115 ( .A(n117), .B(n118), .Z(n114) );
  AND U116 ( .A(n15), .B(n119), .Z(n118) );
  XNOR U117 ( .A(p_input[100]), .B(n117), .Z(n119) );
  XOR U118 ( .A(n120), .B(n121), .Z(n117) );
  AND U119 ( .A(n19), .B(n122), .Z(n121) );
  XNOR U120 ( .A(p_input[132]), .B(n120), .Z(n122) );
  XNOR U121 ( .A(n123), .B(n124), .Z(n120) );
  AND U122 ( .A(n23), .B(n125), .Z(n124) );
  XOR U123 ( .A(p_input[164]), .B(n123), .Z(n125) );
  XOR U124 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n126), .Z(n123) );
  AND U125 ( .A(n26), .B(n127), .Z(n126) );
  XOR U126 ( .A(p_input[196]), .B(\knn_comb_/min_val_out[0][4] ), .Z(n127) );
  XNOR U127 ( .A(n128), .B(n129), .Z(o[3]) );
  AND U128 ( .A(n3), .B(n130), .Z(n128) );
  XNOR U129 ( .A(p_input[3]), .B(n129), .Z(n130) );
  XOR U130 ( .A(n131), .B(n132), .Z(n129) );
  AND U131 ( .A(n7), .B(n133), .Z(n132) );
  XNOR U132 ( .A(p_input[35]), .B(n131), .Z(n133) );
  XOR U133 ( .A(n134), .B(n135), .Z(n131) );
  AND U134 ( .A(n11), .B(n136), .Z(n135) );
  XNOR U135 ( .A(p_input[67]), .B(n134), .Z(n136) );
  XOR U136 ( .A(n137), .B(n138), .Z(n134) );
  AND U137 ( .A(n15), .B(n139), .Z(n138) );
  XNOR U138 ( .A(p_input[99]), .B(n137), .Z(n139) );
  XOR U139 ( .A(n140), .B(n141), .Z(n137) );
  AND U140 ( .A(n19), .B(n142), .Z(n141) );
  XNOR U141 ( .A(p_input[131]), .B(n140), .Z(n142) );
  XNOR U142 ( .A(n143), .B(n144), .Z(n140) );
  AND U143 ( .A(n23), .B(n145), .Z(n144) );
  XOR U144 ( .A(p_input[163]), .B(n143), .Z(n145) );
  XOR U145 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n146), .Z(n143) );
  AND U146 ( .A(n26), .B(n147), .Z(n146) );
  XOR U147 ( .A(p_input[195]), .B(\knn_comb_/min_val_out[0][3] ), .Z(n147) );
  XNOR U148 ( .A(n148), .B(n149), .Z(o[31]) );
  AND U149 ( .A(n3), .B(n150), .Z(n148) );
  XNOR U150 ( .A(p_input[31]), .B(n149), .Z(n150) );
  XOR U151 ( .A(n151), .B(n152), .Z(n149) );
  AND U152 ( .A(n7), .B(n153), .Z(n152) );
  XNOR U153 ( .A(p_input[63]), .B(n151), .Z(n153) );
  XOR U154 ( .A(n154), .B(n155), .Z(n151) );
  AND U155 ( .A(n11), .B(n156), .Z(n155) );
  XNOR U156 ( .A(p_input[95]), .B(n154), .Z(n156) );
  XOR U157 ( .A(n157), .B(n158), .Z(n154) );
  AND U158 ( .A(n15), .B(n159), .Z(n158) );
  XNOR U159 ( .A(p_input[127]), .B(n157), .Z(n159) );
  XOR U160 ( .A(n160), .B(n161), .Z(n157) );
  AND U161 ( .A(n19), .B(n162), .Z(n161) );
  XNOR U162 ( .A(p_input[159]), .B(n160), .Z(n162) );
  XNOR U163 ( .A(n163), .B(n164), .Z(n160) );
  AND U164 ( .A(n23), .B(n165), .Z(n164) );
  XOR U165 ( .A(p_input[191]), .B(n163), .Z(n165) );
  XOR U166 ( .A(\knn_comb_/min_val_out[0][31] ), .B(n166), .Z(n163) );
  AND U167 ( .A(n26), .B(n167), .Z(n166) );
  XOR U168 ( .A(p_input[223]), .B(\knn_comb_/min_val_out[0][31] ), .Z(n167) );
  XNOR U169 ( .A(n168), .B(n169), .Z(o[30]) );
  AND U170 ( .A(n3), .B(n170), .Z(n168) );
  XNOR U171 ( .A(p_input[30]), .B(n169), .Z(n170) );
  XOR U172 ( .A(n171), .B(n172), .Z(n169) );
  AND U173 ( .A(n7), .B(n173), .Z(n172) );
  XNOR U174 ( .A(p_input[62]), .B(n171), .Z(n173) );
  XOR U175 ( .A(n174), .B(n175), .Z(n171) );
  AND U176 ( .A(n11), .B(n176), .Z(n175) );
  XNOR U177 ( .A(p_input[94]), .B(n174), .Z(n176) );
  XOR U178 ( .A(n177), .B(n178), .Z(n174) );
  AND U179 ( .A(n15), .B(n179), .Z(n178) );
  XNOR U180 ( .A(p_input[126]), .B(n177), .Z(n179) );
  XOR U181 ( .A(n180), .B(n181), .Z(n177) );
  AND U182 ( .A(n19), .B(n182), .Z(n181) );
  XNOR U183 ( .A(p_input[158]), .B(n180), .Z(n182) );
  XNOR U184 ( .A(n183), .B(n184), .Z(n180) );
  AND U185 ( .A(n23), .B(n185), .Z(n184) );
  XOR U186 ( .A(p_input[190]), .B(n183), .Z(n185) );
  XOR U187 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n186), .Z(n183) );
  AND U188 ( .A(n26), .B(n187), .Z(n186) );
  XOR U189 ( .A(p_input[222]), .B(\knn_comb_/min_val_out[0][30] ), .Z(n187) );
  XNOR U190 ( .A(n188), .B(n189), .Z(o[2]) );
  AND U191 ( .A(n3), .B(n190), .Z(n188) );
  XNOR U192 ( .A(p_input[2]), .B(n189), .Z(n190) );
  XOR U193 ( .A(n191), .B(n192), .Z(n189) );
  AND U194 ( .A(n7), .B(n193), .Z(n192) );
  XNOR U195 ( .A(p_input[34]), .B(n191), .Z(n193) );
  XOR U196 ( .A(n194), .B(n195), .Z(n191) );
  AND U197 ( .A(n11), .B(n196), .Z(n195) );
  XNOR U198 ( .A(p_input[66]), .B(n194), .Z(n196) );
  XOR U199 ( .A(n197), .B(n198), .Z(n194) );
  AND U200 ( .A(n15), .B(n199), .Z(n198) );
  XNOR U201 ( .A(p_input[98]), .B(n197), .Z(n199) );
  XOR U202 ( .A(n200), .B(n201), .Z(n197) );
  AND U203 ( .A(n19), .B(n202), .Z(n201) );
  XNOR U204 ( .A(p_input[130]), .B(n200), .Z(n202) );
  XNOR U205 ( .A(n203), .B(n204), .Z(n200) );
  AND U206 ( .A(n23), .B(n205), .Z(n204) );
  XOR U207 ( .A(p_input[162]), .B(n203), .Z(n205) );
  XOR U208 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n206), .Z(n203) );
  AND U209 ( .A(n26), .B(n207), .Z(n206) );
  XOR U210 ( .A(p_input[194]), .B(\knn_comb_/min_val_out[0][2] ), .Z(n207) );
  XNOR U211 ( .A(n208), .B(n209), .Z(o[29]) );
  AND U212 ( .A(n3), .B(n210), .Z(n208) );
  XNOR U213 ( .A(p_input[29]), .B(n209), .Z(n210) );
  XOR U214 ( .A(n211), .B(n212), .Z(n209) );
  AND U215 ( .A(n7), .B(n213), .Z(n212) );
  XNOR U216 ( .A(p_input[61]), .B(n211), .Z(n213) );
  XOR U217 ( .A(n214), .B(n215), .Z(n211) );
  AND U218 ( .A(n11), .B(n216), .Z(n215) );
  XNOR U219 ( .A(p_input[93]), .B(n214), .Z(n216) );
  XOR U220 ( .A(n217), .B(n218), .Z(n214) );
  AND U221 ( .A(n15), .B(n219), .Z(n218) );
  XNOR U222 ( .A(p_input[125]), .B(n217), .Z(n219) );
  XOR U223 ( .A(n220), .B(n221), .Z(n217) );
  AND U224 ( .A(n19), .B(n222), .Z(n221) );
  XNOR U225 ( .A(p_input[157]), .B(n220), .Z(n222) );
  XNOR U226 ( .A(n223), .B(n224), .Z(n220) );
  AND U227 ( .A(n23), .B(n225), .Z(n224) );
  XOR U228 ( .A(p_input[189]), .B(n223), .Z(n225) );
  XOR U229 ( .A(\knn_comb_/min_val_out[0][29] ), .B(n226), .Z(n223) );
  AND U230 ( .A(n26), .B(n227), .Z(n226) );
  XOR U231 ( .A(p_input[221]), .B(\knn_comb_/min_val_out[0][29] ), .Z(n227) );
  XNOR U232 ( .A(n228), .B(n229), .Z(o[28]) );
  AND U233 ( .A(n3), .B(n230), .Z(n228) );
  XNOR U234 ( .A(p_input[28]), .B(n229), .Z(n230) );
  XOR U235 ( .A(n231), .B(n232), .Z(n229) );
  AND U236 ( .A(n7), .B(n233), .Z(n232) );
  XNOR U237 ( .A(p_input[60]), .B(n231), .Z(n233) );
  XOR U238 ( .A(n234), .B(n235), .Z(n231) );
  AND U239 ( .A(n11), .B(n236), .Z(n235) );
  XNOR U240 ( .A(p_input[92]), .B(n234), .Z(n236) );
  XOR U241 ( .A(n237), .B(n238), .Z(n234) );
  AND U242 ( .A(n15), .B(n239), .Z(n238) );
  XNOR U243 ( .A(p_input[124]), .B(n237), .Z(n239) );
  XOR U244 ( .A(n240), .B(n241), .Z(n237) );
  AND U245 ( .A(n19), .B(n242), .Z(n241) );
  XNOR U246 ( .A(p_input[156]), .B(n240), .Z(n242) );
  XNOR U247 ( .A(n243), .B(n244), .Z(n240) );
  AND U248 ( .A(n23), .B(n245), .Z(n244) );
  XOR U249 ( .A(p_input[188]), .B(n243), .Z(n245) );
  XOR U250 ( .A(\knn_comb_/min_val_out[0][28] ), .B(n246), .Z(n243) );
  AND U251 ( .A(n26), .B(n247), .Z(n246) );
  XOR U252 ( .A(p_input[220]), .B(\knn_comb_/min_val_out[0][28] ), .Z(n247) );
  XNOR U253 ( .A(n248), .B(n249), .Z(o[27]) );
  AND U254 ( .A(n3), .B(n250), .Z(n248) );
  XNOR U255 ( .A(p_input[27]), .B(n249), .Z(n250) );
  XOR U256 ( .A(n251), .B(n252), .Z(n249) );
  AND U257 ( .A(n7), .B(n253), .Z(n252) );
  XNOR U258 ( .A(p_input[59]), .B(n251), .Z(n253) );
  XOR U259 ( .A(n254), .B(n255), .Z(n251) );
  AND U260 ( .A(n11), .B(n256), .Z(n255) );
  XNOR U261 ( .A(p_input[91]), .B(n254), .Z(n256) );
  XOR U262 ( .A(n257), .B(n258), .Z(n254) );
  AND U263 ( .A(n15), .B(n259), .Z(n258) );
  XNOR U264 ( .A(p_input[123]), .B(n257), .Z(n259) );
  XOR U265 ( .A(n260), .B(n261), .Z(n257) );
  AND U266 ( .A(n19), .B(n262), .Z(n261) );
  XNOR U267 ( .A(p_input[155]), .B(n260), .Z(n262) );
  XNOR U268 ( .A(n263), .B(n264), .Z(n260) );
  AND U269 ( .A(n23), .B(n265), .Z(n264) );
  XOR U270 ( .A(p_input[187]), .B(n263), .Z(n265) );
  XOR U271 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n266), .Z(n263) );
  AND U272 ( .A(n26), .B(n267), .Z(n266) );
  XOR U273 ( .A(p_input[219]), .B(\knn_comb_/min_val_out[0][27] ), .Z(n267) );
  XNOR U274 ( .A(n268), .B(n269), .Z(o[26]) );
  AND U275 ( .A(n3), .B(n270), .Z(n268) );
  XNOR U276 ( .A(p_input[26]), .B(n269), .Z(n270) );
  XOR U277 ( .A(n271), .B(n272), .Z(n269) );
  AND U278 ( .A(n7), .B(n273), .Z(n272) );
  XNOR U279 ( .A(p_input[58]), .B(n271), .Z(n273) );
  XOR U280 ( .A(n274), .B(n275), .Z(n271) );
  AND U281 ( .A(n11), .B(n276), .Z(n275) );
  XNOR U282 ( .A(p_input[90]), .B(n274), .Z(n276) );
  XOR U283 ( .A(n277), .B(n278), .Z(n274) );
  AND U284 ( .A(n15), .B(n279), .Z(n278) );
  XNOR U285 ( .A(p_input[122]), .B(n277), .Z(n279) );
  XOR U286 ( .A(n280), .B(n281), .Z(n277) );
  AND U287 ( .A(n19), .B(n282), .Z(n281) );
  XNOR U288 ( .A(p_input[154]), .B(n280), .Z(n282) );
  XNOR U289 ( .A(n283), .B(n284), .Z(n280) );
  AND U290 ( .A(n23), .B(n285), .Z(n284) );
  XOR U291 ( .A(p_input[186]), .B(n283), .Z(n285) );
  XOR U292 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n286), .Z(n283) );
  AND U293 ( .A(n26), .B(n287), .Z(n286) );
  XOR U294 ( .A(p_input[218]), .B(\knn_comb_/min_val_out[0][26] ), .Z(n287) );
  XNOR U295 ( .A(n288), .B(n289), .Z(o[25]) );
  AND U296 ( .A(n3), .B(n290), .Z(n288) );
  XNOR U297 ( .A(p_input[25]), .B(n289), .Z(n290) );
  XOR U298 ( .A(n291), .B(n292), .Z(n289) );
  AND U299 ( .A(n7), .B(n293), .Z(n292) );
  XNOR U300 ( .A(p_input[57]), .B(n291), .Z(n293) );
  XOR U301 ( .A(n294), .B(n295), .Z(n291) );
  AND U302 ( .A(n11), .B(n296), .Z(n295) );
  XNOR U303 ( .A(p_input[89]), .B(n294), .Z(n296) );
  XOR U304 ( .A(n297), .B(n298), .Z(n294) );
  AND U305 ( .A(n15), .B(n299), .Z(n298) );
  XNOR U306 ( .A(p_input[121]), .B(n297), .Z(n299) );
  XOR U307 ( .A(n300), .B(n301), .Z(n297) );
  AND U308 ( .A(n19), .B(n302), .Z(n301) );
  XNOR U309 ( .A(p_input[153]), .B(n300), .Z(n302) );
  XNOR U310 ( .A(n303), .B(n304), .Z(n300) );
  AND U311 ( .A(n23), .B(n305), .Z(n304) );
  XOR U312 ( .A(p_input[185]), .B(n303), .Z(n305) );
  XOR U313 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n306), .Z(n303) );
  AND U314 ( .A(n26), .B(n307), .Z(n306) );
  XOR U315 ( .A(p_input[217]), .B(\knn_comb_/min_val_out[0][25] ), .Z(n307) );
  XNOR U316 ( .A(n308), .B(n309), .Z(o[24]) );
  AND U317 ( .A(n3), .B(n310), .Z(n308) );
  XNOR U318 ( .A(p_input[24]), .B(n309), .Z(n310) );
  XOR U319 ( .A(n311), .B(n312), .Z(n309) );
  AND U320 ( .A(n7), .B(n313), .Z(n312) );
  XNOR U321 ( .A(p_input[56]), .B(n311), .Z(n313) );
  XOR U322 ( .A(n314), .B(n315), .Z(n311) );
  AND U323 ( .A(n11), .B(n316), .Z(n315) );
  XNOR U324 ( .A(p_input[88]), .B(n314), .Z(n316) );
  XOR U325 ( .A(n317), .B(n318), .Z(n314) );
  AND U326 ( .A(n15), .B(n319), .Z(n318) );
  XNOR U327 ( .A(p_input[120]), .B(n317), .Z(n319) );
  XOR U328 ( .A(n320), .B(n321), .Z(n317) );
  AND U329 ( .A(n19), .B(n322), .Z(n321) );
  XNOR U330 ( .A(p_input[152]), .B(n320), .Z(n322) );
  XNOR U331 ( .A(n323), .B(n324), .Z(n320) );
  AND U332 ( .A(n23), .B(n325), .Z(n324) );
  XOR U333 ( .A(p_input[184]), .B(n323), .Z(n325) );
  XOR U334 ( .A(\knn_comb_/min_val_out[0][24] ), .B(n326), .Z(n323) );
  AND U335 ( .A(n26), .B(n327), .Z(n326) );
  XOR U336 ( .A(p_input[216]), .B(\knn_comb_/min_val_out[0][24] ), .Z(n327) );
  XNOR U337 ( .A(n328), .B(n329), .Z(o[23]) );
  AND U338 ( .A(n3), .B(n330), .Z(n328) );
  XNOR U339 ( .A(p_input[23]), .B(n329), .Z(n330) );
  XOR U340 ( .A(n331), .B(n332), .Z(n329) );
  AND U341 ( .A(n7), .B(n333), .Z(n332) );
  XNOR U342 ( .A(p_input[55]), .B(n331), .Z(n333) );
  XOR U343 ( .A(n334), .B(n335), .Z(n331) );
  AND U344 ( .A(n11), .B(n336), .Z(n335) );
  XNOR U345 ( .A(p_input[87]), .B(n334), .Z(n336) );
  XOR U346 ( .A(n337), .B(n338), .Z(n334) );
  AND U347 ( .A(n15), .B(n339), .Z(n338) );
  XNOR U348 ( .A(p_input[119]), .B(n337), .Z(n339) );
  XOR U349 ( .A(n340), .B(n341), .Z(n337) );
  AND U350 ( .A(n19), .B(n342), .Z(n341) );
  XNOR U351 ( .A(p_input[151]), .B(n340), .Z(n342) );
  XNOR U352 ( .A(n343), .B(n344), .Z(n340) );
  AND U353 ( .A(n23), .B(n345), .Z(n344) );
  XOR U354 ( .A(p_input[183]), .B(n343), .Z(n345) );
  XOR U355 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n346), .Z(n343) );
  AND U356 ( .A(n26), .B(n347), .Z(n346) );
  XOR U357 ( .A(p_input[215]), .B(\knn_comb_/min_val_out[0][23] ), .Z(n347) );
  XNOR U358 ( .A(n348), .B(n349), .Z(o[22]) );
  AND U359 ( .A(n3), .B(n350), .Z(n348) );
  XNOR U360 ( .A(p_input[22]), .B(n349), .Z(n350) );
  XOR U361 ( .A(n351), .B(n352), .Z(n349) );
  AND U362 ( .A(n7), .B(n353), .Z(n352) );
  XNOR U363 ( .A(p_input[54]), .B(n351), .Z(n353) );
  XOR U364 ( .A(n354), .B(n355), .Z(n351) );
  AND U365 ( .A(n11), .B(n356), .Z(n355) );
  XNOR U366 ( .A(p_input[86]), .B(n354), .Z(n356) );
  XOR U367 ( .A(n357), .B(n358), .Z(n354) );
  AND U368 ( .A(n15), .B(n359), .Z(n358) );
  XNOR U369 ( .A(p_input[118]), .B(n357), .Z(n359) );
  XOR U370 ( .A(n360), .B(n361), .Z(n357) );
  AND U371 ( .A(n19), .B(n362), .Z(n361) );
  XNOR U372 ( .A(p_input[150]), .B(n360), .Z(n362) );
  XNOR U373 ( .A(n363), .B(n364), .Z(n360) );
  AND U374 ( .A(n23), .B(n365), .Z(n364) );
  XOR U375 ( .A(p_input[182]), .B(n363), .Z(n365) );
  XOR U376 ( .A(\knn_comb_/min_val_out[0][22] ), .B(n366), .Z(n363) );
  AND U377 ( .A(n26), .B(n367), .Z(n366) );
  XOR U378 ( .A(p_input[214]), .B(\knn_comb_/min_val_out[0][22] ), .Z(n367) );
  XNOR U379 ( .A(n368), .B(n369), .Z(o[21]) );
  AND U380 ( .A(n3), .B(n370), .Z(n368) );
  XNOR U381 ( .A(p_input[21]), .B(n369), .Z(n370) );
  XOR U382 ( .A(n371), .B(n372), .Z(n369) );
  AND U383 ( .A(n7), .B(n373), .Z(n372) );
  XNOR U384 ( .A(p_input[53]), .B(n371), .Z(n373) );
  XOR U385 ( .A(n374), .B(n375), .Z(n371) );
  AND U386 ( .A(n11), .B(n376), .Z(n375) );
  XNOR U387 ( .A(p_input[85]), .B(n374), .Z(n376) );
  XOR U388 ( .A(n377), .B(n378), .Z(n374) );
  AND U389 ( .A(n15), .B(n379), .Z(n378) );
  XNOR U390 ( .A(p_input[117]), .B(n377), .Z(n379) );
  XOR U391 ( .A(n380), .B(n381), .Z(n377) );
  AND U392 ( .A(n19), .B(n382), .Z(n381) );
  XNOR U393 ( .A(p_input[149]), .B(n380), .Z(n382) );
  XNOR U394 ( .A(n383), .B(n384), .Z(n380) );
  AND U395 ( .A(n23), .B(n385), .Z(n384) );
  XOR U396 ( .A(p_input[181]), .B(n383), .Z(n385) );
  XOR U397 ( .A(\knn_comb_/min_val_out[0][21] ), .B(n386), .Z(n383) );
  AND U398 ( .A(n26), .B(n387), .Z(n386) );
  XOR U399 ( .A(p_input[213]), .B(\knn_comb_/min_val_out[0][21] ), .Z(n387) );
  XNOR U400 ( .A(n388), .B(n389), .Z(o[20]) );
  AND U401 ( .A(n3), .B(n390), .Z(n388) );
  XNOR U402 ( .A(p_input[20]), .B(n389), .Z(n390) );
  XOR U403 ( .A(n391), .B(n392), .Z(n389) );
  AND U404 ( .A(n7), .B(n393), .Z(n392) );
  XNOR U405 ( .A(p_input[52]), .B(n391), .Z(n393) );
  XOR U406 ( .A(n394), .B(n395), .Z(n391) );
  AND U407 ( .A(n11), .B(n396), .Z(n395) );
  XNOR U408 ( .A(p_input[84]), .B(n394), .Z(n396) );
  XOR U409 ( .A(n397), .B(n398), .Z(n394) );
  AND U410 ( .A(n15), .B(n399), .Z(n398) );
  XNOR U411 ( .A(p_input[116]), .B(n397), .Z(n399) );
  XOR U412 ( .A(n400), .B(n401), .Z(n397) );
  AND U413 ( .A(n19), .B(n402), .Z(n401) );
  XNOR U414 ( .A(p_input[148]), .B(n400), .Z(n402) );
  XNOR U415 ( .A(n403), .B(n404), .Z(n400) );
  AND U416 ( .A(n23), .B(n405), .Z(n404) );
  XOR U417 ( .A(p_input[180]), .B(n403), .Z(n405) );
  XOR U418 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n406), .Z(n403) );
  AND U419 ( .A(n26), .B(n407), .Z(n406) );
  XOR U420 ( .A(p_input[212]), .B(\knn_comb_/min_val_out[0][20] ), .Z(n407) );
  XNOR U421 ( .A(n408), .B(n409), .Z(o[1]) );
  AND U422 ( .A(n3), .B(n410), .Z(n408) );
  XNOR U423 ( .A(p_input[1]), .B(n409), .Z(n410) );
  XOR U424 ( .A(n411), .B(n412), .Z(n409) );
  AND U425 ( .A(n7), .B(n413), .Z(n412) );
  XNOR U426 ( .A(p_input[33]), .B(n411), .Z(n413) );
  XOR U427 ( .A(n414), .B(n415), .Z(n411) );
  AND U428 ( .A(n11), .B(n416), .Z(n415) );
  XNOR U429 ( .A(p_input[65]), .B(n414), .Z(n416) );
  XOR U430 ( .A(n417), .B(n418), .Z(n414) );
  AND U431 ( .A(n15), .B(n419), .Z(n418) );
  XNOR U432 ( .A(p_input[97]), .B(n417), .Z(n419) );
  XOR U433 ( .A(n420), .B(n421), .Z(n417) );
  AND U434 ( .A(n19), .B(n422), .Z(n421) );
  XNOR U435 ( .A(p_input[129]), .B(n420), .Z(n422) );
  XNOR U436 ( .A(n423), .B(n424), .Z(n420) );
  AND U437 ( .A(n23), .B(n425), .Z(n424) );
  XOR U438 ( .A(p_input[161]), .B(n423), .Z(n425) );
  XOR U439 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n426), .Z(n423) );
  AND U440 ( .A(n26), .B(n427), .Z(n426) );
  XOR U441 ( .A(p_input[193]), .B(\knn_comb_/min_val_out[0][1] ), .Z(n427) );
  XNOR U442 ( .A(n428), .B(n429), .Z(o[19]) );
  AND U443 ( .A(n3), .B(n430), .Z(n428) );
  XNOR U444 ( .A(p_input[19]), .B(n429), .Z(n430) );
  XOR U445 ( .A(n431), .B(n432), .Z(n429) );
  AND U446 ( .A(n7), .B(n433), .Z(n432) );
  XNOR U447 ( .A(p_input[51]), .B(n431), .Z(n433) );
  XOR U448 ( .A(n434), .B(n435), .Z(n431) );
  AND U449 ( .A(n11), .B(n436), .Z(n435) );
  XNOR U450 ( .A(p_input[83]), .B(n434), .Z(n436) );
  XOR U451 ( .A(n437), .B(n438), .Z(n434) );
  AND U452 ( .A(n15), .B(n439), .Z(n438) );
  XNOR U453 ( .A(p_input[115]), .B(n437), .Z(n439) );
  XOR U454 ( .A(n440), .B(n441), .Z(n437) );
  AND U455 ( .A(n19), .B(n442), .Z(n441) );
  XNOR U456 ( .A(p_input[147]), .B(n440), .Z(n442) );
  XNOR U457 ( .A(n443), .B(n444), .Z(n440) );
  AND U458 ( .A(n23), .B(n445), .Z(n444) );
  XOR U459 ( .A(p_input[179]), .B(n443), .Z(n445) );
  XOR U460 ( .A(\knn_comb_/min_val_out[0][19] ), .B(n446), .Z(n443) );
  AND U461 ( .A(n26), .B(n447), .Z(n446) );
  XOR U462 ( .A(p_input[211]), .B(\knn_comb_/min_val_out[0][19] ), .Z(n447) );
  XNOR U463 ( .A(n448), .B(n449), .Z(o[18]) );
  AND U464 ( .A(n3), .B(n450), .Z(n448) );
  XNOR U465 ( .A(p_input[18]), .B(n449), .Z(n450) );
  XOR U466 ( .A(n451), .B(n452), .Z(n449) );
  AND U467 ( .A(n7), .B(n453), .Z(n452) );
  XNOR U468 ( .A(p_input[50]), .B(n451), .Z(n453) );
  XOR U469 ( .A(n454), .B(n455), .Z(n451) );
  AND U470 ( .A(n11), .B(n456), .Z(n455) );
  XNOR U471 ( .A(p_input[82]), .B(n454), .Z(n456) );
  XOR U472 ( .A(n457), .B(n458), .Z(n454) );
  AND U473 ( .A(n15), .B(n459), .Z(n458) );
  XNOR U474 ( .A(p_input[114]), .B(n457), .Z(n459) );
  XOR U475 ( .A(n460), .B(n461), .Z(n457) );
  AND U476 ( .A(n19), .B(n462), .Z(n461) );
  XNOR U477 ( .A(p_input[146]), .B(n460), .Z(n462) );
  XNOR U478 ( .A(n463), .B(n464), .Z(n460) );
  AND U479 ( .A(n23), .B(n465), .Z(n464) );
  XOR U480 ( .A(p_input[178]), .B(n463), .Z(n465) );
  XOR U481 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n466), .Z(n463) );
  AND U482 ( .A(n26), .B(n467), .Z(n466) );
  XOR U483 ( .A(p_input[210]), .B(\knn_comb_/min_val_out[0][18] ), .Z(n467) );
  XNOR U484 ( .A(n468), .B(n469), .Z(o[17]) );
  AND U485 ( .A(n3), .B(n470), .Z(n468) );
  XNOR U486 ( .A(p_input[17]), .B(n469), .Z(n470) );
  XOR U487 ( .A(n471), .B(n472), .Z(n469) );
  AND U488 ( .A(n7), .B(n473), .Z(n472) );
  XNOR U489 ( .A(p_input[49]), .B(n471), .Z(n473) );
  XOR U490 ( .A(n474), .B(n475), .Z(n471) );
  AND U491 ( .A(n11), .B(n476), .Z(n475) );
  XNOR U492 ( .A(p_input[81]), .B(n474), .Z(n476) );
  XOR U493 ( .A(n477), .B(n478), .Z(n474) );
  AND U494 ( .A(n15), .B(n479), .Z(n478) );
  XNOR U495 ( .A(p_input[113]), .B(n477), .Z(n479) );
  XOR U496 ( .A(n480), .B(n481), .Z(n477) );
  AND U497 ( .A(n19), .B(n482), .Z(n481) );
  XNOR U498 ( .A(p_input[145]), .B(n480), .Z(n482) );
  XNOR U499 ( .A(n483), .B(n484), .Z(n480) );
  AND U500 ( .A(n23), .B(n485), .Z(n484) );
  XOR U501 ( .A(p_input[177]), .B(n483), .Z(n485) );
  XOR U502 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n486), .Z(n483) );
  AND U503 ( .A(n26), .B(n487), .Z(n486) );
  XOR U504 ( .A(p_input[209]), .B(\knn_comb_/min_val_out[0][17] ), .Z(n487) );
  XNOR U505 ( .A(n488), .B(n489), .Z(o[16]) );
  AND U506 ( .A(n3), .B(n490), .Z(n488) );
  XNOR U507 ( .A(p_input[16]), .B(n489), .Z(n490) );
  XOR U508 ( .A(n491), .B(n492), .Z(n489) );
  AND U509 ( .A(n7), .B(n493), .Z(n492) );
  XNOR U510 ( .A(p_input[48]), .B(n491), .Z(n493) );
  XOR U511 ( .A(n494), .B(n495), .Z(n491) );
  AND U512 ( .A(n11), .B(n496), .Z(n495) );
  XNOR U513 ( .A(p_input[80]), .B(n494), .Z(n496) );
  XOR U514 ( .A(n497), .B(n498), .Z(n494) );
  AND U515 ( .A(n15), .B(n499), .Z(n498) );
  XNOR U516 ( .A(p_input[112]), .B(n497), .Z(n499) );
  XOR U517 ( .A(n500), .B(n501), .Z(n497) );
  AND U518 ( .A(n19), .B(n502), .Z(n501) );
  XNOR U519 ( .A(p_input[144]), .B(n500), .Z(n502) );
  XNOR U520 ( .A(n503), .B(n504), .Z(n500) );
  AND U521 ( .A(n23), .B(n505), .Z(n504) );
  XOR U522 ( .A(p_input[176]), .B(n503), .Z(n505) );
  XOR U523 ( .A(\knn_comb_/min_val_out[0][16] ), .B(n506), .Z(n503) );
  AND U524 ( .A(n26), .B(n507), .Z(n506) );
  XOR U525 ( .A(p_input[208]), .B(\knn_comb_/min_val_out[0][16] ), .Z(n507) );
  XNOR U526 ( .A(n508), .B(n509), .Z(o[15]) );
  AND U527 ( .A(n3), .B(n510), .Z(n508) );
  XNOR U528 ( .A(p_input[15]), .B(n509), .Z(n510) );
  XOR U529 ( .A(n511), .B(n512), .Z(n509) );
  AND U530 ( .A(n7), .B(n513), .Z(n512) );
  XNOR U531 ( .A(p_input[47]), .B(n511), .Z(n513) );
  XOR U532 ( .A(n514), .B(n515), .Z(n511) );
  AND U533 ( .A(n11), .B(n516), .Z(n515) );
  XNOR U534 ( .A(p_input[79]), .B(n514), .Z(n516) );
  XOR U535 ( .A(n517), .B(n518), .Z(n514) );
  AND U536 ( .A(n15), .B(n519), .Z(n518) );
  XNOR U537 ( .A(p_input[111]), .B(n517), .Z(n519) );
  XOR U538 ( .A(n520), .B(n521), .Z(n517) );
  AND U539 ( .A(n19), .B(n522), .Z(n521) );
  XNOR U540 ( .A(p_input[143]), .B(n520), .Z(n522) );
  XNOR U541 ( .A(n523), .B(n524), .Z(n520) );
  AND U542 ( .A(n23), .B(n525), .Z(n524) );
  XOR U543 ( .A(p_input[175]), .B(n523), .Z(n525) );
  XOR U544 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n526), .Z(n523) );
  AND U545 ( .A(n26), .B(n527), .Z(n526) );
  XOR U546 ( .A(p_input[207]), .B(\knn_comb_/min_val_out[0][15] ), .Z(n527) );
  XNOR U547 ( .A(n528), .B(n529), .Z(o[14]) );
  AND U548 ( .A(n3), .B(n530), .Z(n528) );
  XNOR U549 ( .A(p_input[14]), .B(n529), .Z(n530) );
  XOR U550 ( .A(n531), .B(n532), .Z(n529) );
  AND U551 ( .A(n7), .B(n533), .Z(n532) );
  XNOR U552 ( .A(p_input[46]), .B(n531), .Z(n533) );
  XOR U553 ( .A(n534), .B(n535), .Z(n531) );
  AND U554 ( .A(n11), .B(n536), .Z(n535) );
  XNOR U555 ( .A(p_input[78]), .B(n534), .Z(n536) );
  XOR U556 ( .A(n537), .B(n538), .Z(n534) );
  AND U557 ( .A(n15), .B(n539), .Z(n538) );
  XNOR U558 ( .A(p_input[110]), .B(n537), .Z(n539) );
  XOR U559 ( .A(n540), .B(n541), .Z(n537) );
  AND U560 ( .A(n19), .B(n542), .Z(n541) );
  XNOR U561 ( .A(p_input[142]), .B(n540), .Z(n542) );
  XNOR U562 ( .A(n543), .B(n544), .Z(n540) );
  AND U563 ( .A(n23), .B(n545), .Z(n544) );
  XOR U564 ( .A(p_input[174]), .B(n543), .Z(n545) );
  XOR U565 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n546), .Z(n543) );
  AND U566 ( .A(n26), .B(n547), .Z(n546) );
  XOR U567 ( .A(p_input[206]), .B(\knn_comb_/min_val_out[0][14] ), .Z(n547) );
  XNOR U568 ( .A(n548), .B(n549), .Z(o[13]) );
  AND U569 ( .A(n3), .B(n550), .Z(n548) );
  XNOR U570 ( .A(p_input[13]), .B(n549), .Z(n550) );
  XOR U571 ( .A(n551), .B(n552), .Z(n549) );
  AND U572 ( .A(n7), .B(n553), .Z(n552) );
  XNOR U573 ( .A(p_input[45]), .B(n551), .Z(n553) );
  XOR U574 ( .A(n554), .B(n555), .Z(n551) );
  AND U575 ( .A(n11), .B(n556), .Z(n555) );
  XNOR U576 ( .A(p_input[77]), .B(n554), .Z(n556) );
  XOR U577 ( .A(n557), .B(n558), .Z(n554) );
  AND U578 ( .A(n15), .B(n559), .Z(n558) );
  XNOR U579 ( .A(p_input[109]), .B(n557), .Z(n559) );
  XOR U580 ( .A(n560), .B(n561), .Z(n557) );
  AND U581 ( .A(n19), .B(n562), .Z(n561) );
  XNOR U582 ( .A(p_input[141]), .B(n560), .Z(n562) );
  XNOR U583 ( .A(n563), .B(n564), .Z(n560) );
  AND U584 ( .A(n23), .B(n565), .Z(n564) );
  XOR U585 ( .A(p_input[173]), .B(n563), .Z(n565) );
  XOR U586 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n566), .Z(n563) );
  AND U587 ( .A(n26), .B(n567), .Z(n566) );
  XOR U588 ( .A(p_input[205]), .B(\knn_comb_/min_val_out[0][13] ), .Z(n567) );
  XNOR U589 ( .A(n568), .B(n569), .Z(o[12]) );
  AND U590 ( .A(n3), .B(n570), .Z(n568) );
  XNOR U591 ( .A(p_input[12]), .B(n569), .Z(n570) );
  XOR U592 ( .A(n571), .B(n572), .Z(n569) );
  AND U593 ( .A(n7), .B(n573), .Z(n572) );
  XNOR U594 ( .A(p_input[44]), .B(n571), .Z(n573) );
  XOR U595 ( .A(n574), .B(n575), .Z(n571) );
  AND U596 ( .A(n11), .B(n576), .Z(n575) );
  XNOR U597 ( .A(p_input[76]), .B(n574), .Z(n576) );
  XOR U598 ( .A(n577), .B(n578), .Z(n574) );
  AND U599 ( .A(n15), .B(n579), .Z(n578) );
  XNOR U600 ( .A(p_input[108]), .B(n577), .Z(n579) );
  XOR U601 ( .A(n580), .B(n581), .Z(n577) );
  AND U602 ( .A(n19), .B(n582), .Z(n581) );
  XNOR U603 ( .A(p_input[140]), .B(n580), .Z(n582) );
  XNOR U604 ( .A(n583), .B(n584), .Z(n580) );
  AND U605 ( .A(n23), .B(n585), .Z(n584) );
  XOR U606 ( .A(p_input[172]), .B(n583), .Z(n585) );
  XOR U607 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n586), .Z(n583) );
  AND U608 ( .A(n26), .B(n587), .Z(n586) );
  XOR U609 ( .A(p_input[204]), .B(\knn_comb_/min_val_out[0][12] ), .Z(n587) );
  XNOR U610 ( .A(n588), .B(n589), .Z(o[11]) );
  AND U611 ( .A(n3), .B(n590), .Z(n588) );
  XNOR U612 ( .A(p_input[11]), .B(n589), .Z(n590) );
  XOR U613 ( .A(n591), .B(n592), .Z(n589) );
  AND U614 ( .A(n7), .B(n593), .Z(n592) );
  XNOR U615 ( .A(p_input[43]), .B(n591), .Z(n593) );
  XOR U616 ( .A(n594), .B(n595), .Z(n591) );
  AND U617 ( .A(n11), .B(n596), .Z(n595) );
  XNOR U618 ( .A(p_input[75]), .B(n594), .Z(n596) );
  XOR U619 ( .A(n597), .B(n598), .Z(n594) );
  AND U620 ( .A(n15), .B(n599), .Z(n598) );
  XNOR U621 ( .A(p_input[107]), .B(n597), .Z(n599) );
  XOR U622 ( .A(n600), .B(n601), .Z(n597) );
  AND U623 ( .A(n19), .B(n602), .Z(n601) );
  XNOR U624 ( .A(p_input[139]), .B(n600), .Z(n602) );
  XNOR U625 ( .A(n603), .B(n604), .Z(n600) );
  AND U626 ( .A(n23), .B(n605), .Z(n604) );
  XOR U627 ( .A(p_input[171]), .B(n603), .Z(n605) );
  XOR U628 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n606), .Z(n603) );
  AND U629 ( .A(n26), .B(n607), .Z(n606) );
  XOR U630 ( .A(p_input[203]), .B(\knn_comb_/min_val_out[0][11] ), .Z(n607) );
  XNOR U631 ( .A(n608), .B(n609), .Z(o[10]) );
  AND U632 ( .A(n3), .B(n610), .Z(n608) );
  XNOR U633 ( .A(p_input[10]), .B(n609), .Z(n610) );
  XOR U634 ( .A(n611), .B(n612), .Z(n609) );
  AND U635 ( .A(n7), .B(n613), .Z(n612) );
  XNOR U636 ( .A(p_input[42]), .B(n611), .Z(n613) );
  XOR U637 ( .A(n614), .B(n615), .Z(n611) );
  AND U638 ( .A(n11), .B(n616), .Z(n615) );
  XNOR U639 ( .A(p_input[74]), .B(n614), .Z(n616) );
  XOR U640 ( .A(n617), .B(n618), .Z(n614) );
  AND U641 ( .A(n15), .B(n619), .Z(n618) );
  XNOR U642 ( .A(p_input[106]), .B(n617), .Z(n619) );
  XOR U643 ( .A(n620), .B(n621), .Z(n617) );
  AND U644 ( .A(n19), .B(n622), .Z(n621) );
  XNOR U645 ( .A(p_input[138]), .B(n620), .Z(n622) );
  XNOR U646 ( .A(n623), .B(n624), .Z(n620) );
  AND U647 ( .A(n23), .B(n625), .Z(n624) );
  XOR U648 ( .A(p_input[170]), .B(n623), .Z(n625) );
  XOR U649 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n626), .Z(n623) );
  AND U650 ( .A(n26), .B(n627), .Z(n626) );
  XOR U651 ( .A(p_input[202]), .B(\knn_comb_/min_val_out[0][10] ), .Z(n627) );
  XNOR U652 ( .A(n628), .B(n629), .Z(o[0]) );
  AND U653 ( .A(n3), .B(n630), .Z(n628) );
  XNOR U654 ( .A(p_input[0]), .B(n629), .Z(n630) );
  XOR U655 ( .A(n631), .B(n632), .Z(n629) );
  AND U656 ( .A(n7), .B(n633), .Z(n632) );
  XNOR U657 ( .A(p_input[32]), .B(n631), .Z(n633) );
  XOR U658 ( .A(n634), .B(n635), .Z(n631) );
  AND U659 ( .A(n11), .B(n636), .Z(n635) );
  XNOR U660 ( .A(p_input[64]), .B(n634), .Z(n636) );
  XOR U661 ( .A(n637), .B(n638), .Z(n634) );
  AND U662 ( .A(n15), .B(n639), .Z(n638) );
  XNOR U663 ( .A(p_input[96]), .B(n637), .Z(n639) );
  XOR U664 ( .A(n640), .B(n641), .Z(n637) );
  AND U665 ( .A(n19), .B(n642), .Z(n641) );
  XNOR U666 ( .A(p_input[128]), .B(n640), .Z(n642) );
  XNOR U667 ( .A(n643), .B(n644), .Z(n640) );
  AND U668 ( .A(n23), .B(n645), .Z(n644) );
  XOR U669 ( .A(p_input[160]), .B(n643), .Z(n645) );
  XOR U670 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n646), .Z(n643) );
  AND U671 ( .A(n26), .B(n647), .Z(n646) );
  XOR U672 ( .A(p_input[192]), .B(\knn_comb_/min_val_out[0][0] ), .Z(n647) );
  XNOR U673 ( .A(n648), .B(n649), .Z(n3) );
  NOR U674 ( .A(n650), .B(n651), .Z(n649) );
  XOR U675 ( .A(n652), .B(n648), .Z(n651) );
  AND U676 ( .A(n653), .B(n654), .Z(n652) );
  NOR U677 ( .A(n655), .B(n648), .Z(n650) );
  AND U678 ( .A(n656), .B(n657), .Z(n655) );
  XOR U679 ( .A(n658), .B(n659), .Z(n648) );
  AND U680 ( .A(n660), .B(n661), .Z(n659) );
  XNOR U681 ( .A(n658), .B(n656), .Z(n661) );
  XNOR U682 ( .A(n662), .B(n663), .Z(n656) );
  XOR U683 ( .A(n664), .B(n657), .Z(n663) );
  AND U684 ( .A(n665), .B(n666), .Z(n657) );
  AND U685 ( .A(n667), .B(n668), .Z(n664) );
  XOR U686 ( .A(n669), .B(n662), .Z(n667) );
  XOR U687 ( .A(n670), .B(n658), .Z(n660) );
  XNOR U688 ( .A(n671), .B(n672), .Z(n670) );
  AND U689 ( .A(n7), .B(n673), .Z(n672) );
  XOR U690 ( .A(n674), .B(n671), .Z(n673) );
  XOR U691 ( .A(n675), .B(n676), .Z(n658) );
  AND U692 ( .A(n677), .B(n678), .Z(n676) );
  XNOR U693 ( .A(n675), .B(n665), .Z(n678) );
  XOR U694 ( .A(n679), .B(n668), .Z(n665) );
  XNOR U695 ( .A(n680), .B(n662), .Z(n668) );
  XOR U696 ( .A(n681), .B(n682), .Z(n662) );
  AND U697 ( .A(n683), .B(n684), .Z(n682) );
  XOR U698 ( .A(n685), .B(n681), .Z(n683) );
  XNOR U699 ( .A(n686), .B(n687), .Z(n680) );
  AND U700 ( .A(n688), .B(n689), .Z(n687) );
  XOR U701 ( .A(n686), .B(n690), .Z(n688) );
  XNOR U702 ( .A(n669), .B(n666), .Z(n679) );
  AND U703 ( .A(n691), .B(n692), .Z(n666) );
  XOR U704 ( .A(n693), .B(n694), .Z(n669) );
  AND U705 ( .A(n695), .B(n696), .Z(n694) );
  XOR U706 ( .A(n693), .B(n697), .Z(n695) );
  XOR U707 ( .A(n698), .B(n675), .Z(n677) );
  XNOR U708 ( .A(n699), .B(n700), .Z(n698) );
  AND U709 ( .A(n7), .B(n701), .Z(n700) );
  XNOR U710 ( .A(n702), .B(n699), .Z(n701) );
  XOR U711 ( .A(n703), .B(n704), .Z(n675) );
  AND U712 ( .A(n705), .B(n706), .Z(n704) );
  XNOR U713 ( .A(n703), .B(n691), .Z(n706) );
  XOR U714 ( .A(n707), .B(n684), .Z(n691) );
  XNOR U715 ( .A(n708), .B(n690), .Z(n684) );
  XOR U716 ( .A(n709), .B(n710), .Z(n690) );
  AND U717 ( .A(n711), .B(n712), .Z(n710) );
  XOR U718 ( .A(n709), .B(n713), .Z(n711) );
  XNOR U719 ( .A(n689), .B(n681), .Z(n708) );
  XOR U720 ( .A(n714), .B(n715), .Z(n681) );
  AND U721 ( .A(n716), .B(n717), .Z(n715) );
  XNOR U722 ( .A(n718), .B(n714), .Z(n716) );
  XNOR U723 ( .A(n719), .B(n686), .Z(n689) );
  XOR U724 ( .A(n720), .B(n721), .Z(n686) );
  AND U725 ( .A(n722), .B(n723), .Z(n721) );
  XOR U726 ( .A(n720), .B(n724), .Z(n722) );
  XNOR U727 ( .A(n725), .B(n726), .Z(n719) );
  AND U728 ( .A(n727), .B(n728), .Z(n726) );
  XNOR U729 ( .A(n725), .B(n729), .Z(n727) );
  XNOR U730 ( .A(n685), .B(n692), .Z(n707) );
  AND U731 ( .A(n730), .B(n731), .Z(n692) );
  XOR U732 ( .A(n697), .B(n696), .Z(n685) );
  XNOR U733 ( .A(n732), .B(n693), .Z(n696) );
  XOR U734 ( .A(n733), .B(n734), .Z(n693) );
  AND U735 ( .A(n735), .B(n736), .Z(n734) );
  XOR U736 ( .A(n733), .B(n737), .Z(n735) );
  XNOR U737 ( .A(n738), .B(n739), .Z(n732) );
  AND U738 ( .A(n740), .B(n741), .Z(n739) );
  XOR U739 ( .A(n738), .B(n742), .Z(n740) );
  XOR U740 ( .A(n743), .B(n744), .Z(n697) );
  AND U741 ( .A(n745), .B(n746), .Z(n744) );
  XOR U742 ( .A(n743), .B(n747), .Z(n745) );
  XOR U743 ( .A(n748), .B(n703), .Z(n705) );
  XNOR U744 ( .A(n749), .B(n750), .Z(n748) );
  AND U745 ( .A(n7), .B(n751), .Z(n750) );
  XOR U746 ( .A(n752), .B(n749), .Z(n751) );
  XOR U747 ( .A(n753), .B(n754), .Z(n703) );
  AND U748 ( .A(n755), .B(n756), .Z(n754) );
  XNOR U749 ( .A(n753), .B(n730), .Z(n756) );
  XOR U750 ( .A(n757), .B(n717), .Z(n730) );
  XNOR U751 ( .A(n758), .B(n724), .Z(n717) );
  XOR U752 ( .A(n713), .B(n712), .Z(n724) );
  XNOR U753 ( .A(n759), .B(n709), .Z(n712) );
  XOR U754 ( .A(n760), .B(n761), .Z(n709) );
  AND U755 ( .A(n762), .B(n763), .Z(n761) );
  XNOR U756 ( .A(n764), .B(n765), .Z(n762) );
  IV U757 ( .A(n760), .Z(n764) );
  XNOR U758 ( .A(n766), .B(n767), .Z(n759) );
  NOR U759 ( .A(n768), .B(n769), .Z(n767) );
  XNOR U760 ( .A(n766), .B(n770), .Z(n768) );
  XOR U761 ( .A(n771), .B(n772), .Z(n713) );
  NOR U762 ( .A(n773), .B(n774), .Z(n772) );
  XNOR U763 ( .A(n771), .B(n775), .Z(n773) );
  XNOR U764 ( .A(n723), .B(n714), .Z(n758) );
  XOR U765 ( .A(n776), .B(n777), .Z(n714) );
  AND U766 ( .A(n778), .B(n779), .Z(n777) );
  XOR U767 ( .A(n776), .B(n780), .Z(n778) );
  XOR U768 ( .A(n781), .B(n729), .Z(n723) );
  XOR U769 ( .A(n782), .B(n783), .Z(n729) );
  NOR U770 ( .A(n784), .B(n785), .Z(n783) );
  XOR U771 ( .A(n782), .B(n786), .Z(n784) );
  XNOR U772 ( .A(n728), .B(n720), .Z(n781) );
  XOR U773 ( .A(n787), .B(n788), .Z(n720) );
  AND U774 ( .A(n789), .B(n790), .Z(n788) );
  XOR U775 ( .A(n787), .B(n791), .Z(n789) );
  XNOR U776 ( .A(n792), .B(n725), .Z(n728) );
  XOR U777 ( .A(n793), .B(n794), .Z(n725) );
  AND U778 ( .A(n795), .B(n796), .Z(n794) );
  XNOR U779 ( .A(n797), .B(n798), .Z(n795) );
  IV U780 ( .A(n793), .Z(n797) );
  XNOR U781 ( .A(n799), .B(n800), .Z(n792) );
  NOR U782 ( .A(n801), .B(n802), .Z(n800) );
  XOR U783 ( .A(n799), .B(n803), .Z(n801) );
  XOR U784 ( .A(n718), .B(n731), .Z(n757) );
  NOR U785 ( .A(n804), .B(n805), .Z(n731) );
  XNOR U786 ( .A(n737), .B(n736), .Z(n718) );
  XNOR U787 ( .A(n806), .B(n742), .Z(n736) );
  XNOR U788 ( .A(n807), .B(n808), .Z(n742) );
  NOR U789 ( .A(n809), .B(n810), .Z(n808) );
  XOR U790 ( .A(n807), .B(n811), .Z(n809) );
  XNOR U791 ( .A(n741), .B(n733), .Z(n806) );
  XOR U792 ( .A(n812), .B(n813), .Z(n733) );
  AND U793 ( .A(n814), .B(n815), .Z(n813) );
  XNOR U794 ( .A(n812), .B(n816), .Z(n814) );
  XNOR U795 ( .A(n817), .B(n738), .Z(n741) );
  XOR U796 ( .A(n818), .B(n819), .Z(n738) );
  AND U797 ( .A(n820), .B(n821), .Z(n819) );
  XNOR U798 ( .A(n822), .B(n823), .Z(n820) );
  IV U799 ( .A(n818), .Z(n822) );
  XNOR U800 ( .A(n824), .B(n825), .Z(n817) );
  NOR U801 ( .A(n826), .B(n827), .Z(n825) );
  XNOR U802 ( .A(n824), .B(n828), .Z(n826) );
  XOR U803 ( .A(n747), .B(n746), .Z(n737) );
  XNOR U804 ( .A(n829), .B(n743), .Z(n746) );
  XOR U805 ( .A(n830), .B(n831), .Z(n743) );
  AND U806 ( .A(n832), .B(n833), .Z(n831) );
  XOR U807 ( .A(n830), .B(n834), .Z(n832) );
  XNOR U808 ( .A(n835), .B(n836), .Z(n829) );
  NOR U809 ( .A(n837), .B(n838), .Z(n836) );
  XNOR U810 ( .A(n835), .B(n839), .Z(n837) );
  XOR U811 ( .A(n840), .B(n841), .Z(n747) );
  NOR U812 ( .A(n842), .B(n843), .Z(n841) );
  XNOR U813 ( .A(n840), .B(n844), .Z(n842) );
  XNOR U814 ( .A(n845), .B(n846), .Z(n755) );
  XOR U815 ( .A(n753), .B(n847), .Z(n846) );
  AND U816 ( .A(n7), .B(n848), .Z(n847) );
  XNOR U817 ( .A(n849), .B(n845), .Z(n848) );
  AND U818 ( .A(n850), .B(n804), .Z(n753) );
  XOR U819 ( .A(n851), .B(n805), .Z(n804) );
  XNOR U820 ( .A(p_input[0]), .B(p_input[256]), .Z(n805) );
  XNOR U821 ( .A(n780), .B(n779), .Z(n851) );
  XNOR U822 ( .A(n852), .B(n791), .Z(n779) );
  XOR U823 ( .A(n765), .B(n763), .Z(n791) );
  XNOR U824 ( .A(n853), .B(n770), .Z(n763) );
  XOR U825 ( .A(p_input[24]), .B(p_input[280]), .Z(n770) );
  XOR U826 ( .A(n760), .B(n769), .Z(n853) );
  XOR U827 ( .A(n854), .B(n766), .Z(n769) );
  XOR U828 ( .A(p_input[22]), .B(p_input[278]), .Z(n766) );
  XOR U829 ( .A(p_input[23]), .B(n855), .Z(n854) );
  XOR U830 ( .A(p_input[18]), .B(p_input[274]), .Z(n760) );
  XNOR U831 ( .A(n775), .B(n774), .Z(n765) );
  XOR U832 ( .A(n856), .B(n771), .Z(n774) );
  XOR U833 ( .A(p_input[19]), .B(p_input[275]), .Z(n771) );
  XOR U834 ( .A(p_input[20]), .B(n857), .Z(n856) );
  XOR U835 ( .A(p_input[21]), .B(p_input[277]), .Z(n775) );
  XOR U836 ( .A(n790), .B(n858), .Z(n852) );
  IV U837 ( .A(n776), .Z(n858) );
  XOR U838 ( .A(p_input[1]), .B(p_input[257]), .Z(n776) );
  XNOR U839 ( .A(n859), .B(n798), .Z(n790) );
  XNOR U840 ( .A(n786), .B(n785), .Z(n798) );
  XNOR U841 ( .A(n860), .B(n782), .Z(n785) );
  XNOR U842 ( .A(p_input[26]), .B(p_input[282]), .Z(n782) );
  XOR U843 ( .A(p_input[27]), .B(n861), .Z(n860) );
  XOR U844 ( .A(p_input[284]), .B(p_input[28]), .Z(n786) );
  XOR U845 ( .A(n796), .B(n862), .Z(n859) );
  IV U846 ( .A(n787), .Z(n862) );
  XOR U847 ( .A(p_input[17]), .B(p_input[273]), .Z(n787) );
  XOR U848 ( .A(n863), .B(n803), .Z(n796) );
  XNOR U849 ( .A(p_input[287]), .B(p_input[31]), .Z(n803) );
  XOR U850 ( .A(n793), .B(n802), .Z(n863) );
  XOR U851 ( .A(n864), .B(n799), .Z(n802) );
  XOR U852 ( .A(p_input[285]), .B(p_input[29]), .Z(n799) );
  XNOR U853 ( .A(p_input[286]), .B(p_input[30]), .Z(n864) );
  XOR U854 ( .A(p_input[25]), .B(p_input[281]), .Z(n793) );
  XNOR U855 ( .A(n816), .B(n815), .Z(n780) );
  XNOR U856 ( .A(n865), .B(n823), .Z(n815) );
  XNOR U857 ( .A(n811), .B(n810), .Z(n823) );
  XNOR U858 ( .A(n866), .B(n807), .Z(n810) );
  XNOR U859 ( .A(p_input[11]), .B(p_input[267]), .Z(n807) );
  XOR U860 ( .A(p_input[12]), .B(n867), .Z(n866) );
  XOR U861 ( .A(p_input[13]), .B(p_input[269]), .Z(n811) );
  XNOR U862 ( .A(n821), .B(n812), .Z(n865) );
  XOR U863 ( .A(p_input[258]), .B(p_input[2]), .Z(n812) );
  XNOR U864 ( .A(n868), .B(n828), .Z(n821) );
  XNOR U865 ( .A(p_input[16]), .B(n869), .Z(n828) );
  XOR U866 ( .A(n818), .B(n827), .Z(n868) );
  XOR U867 ( .A(n870), .B(n824), .Z(n827) );
  XOR U868 ( .A(p_input[14]), .B(p_input[270]), .Z(n824) );
  XOR U869 ( .A(p_input[15]), .B(n871), .Z(n870) );
  XOR U870 ( .A(p_input[10]), .B(p_input[266]), .Z(n818) );
  XNOR U871 ( .A(n834), .B(n833), .Z(n816) );
  XNOR U872 ( .A(n872), .B(n839), .Z(n833) );
  XOR U873 ( .A(p_input[265]), .B(p_input[9]), .Z(n839) );
  XOR U874 ( .A(n830), .B(n838), .Z(n872) );
  XOR U875 ( .A(n873), .B(n835), .Z(n838) );
  XOR U876 ( .A(p_input[263]), .B(p_input[7]), .Z(n835) );
  XNOR U877 ( .A(p_input[264]), .B(p_input[8]), .Z(n873) );
  XOR U878 ( .A(p_input[259]), .B(p_input[3]), .Z(n830) );
  XNOR U879 ( .A(n844), .B(n843), .Z(n834) );
  XOR U880 ( .A(n874), .B(n840), .Z(n843) );
  XOR U881 ( .A(p_input[260]), .B(p_input[4]), .Z(n840) );
  XNOR U882 ( .A(p_input[261]), .B(p_input[5]), .Z(n874) );
  XOR U883 ( .A(p_input[262]), .B(p_input[6]), .Z(n844) );
  XNOR U884 ( .A(n875), .B(n876), .Z(n850) );
  AND U885 ( .A(n7), .B(n877), .Z(n876) );
  XNOR U886 ( .A(n878), .B(n879), .Z(n877) );
  XNOR U887 ( .A(n880), .B(n881), .Z(n7) );
  NOR U888 ( .A(n882), .B(n883), .Z(n881) );
  XOR U889 ( .A(n654), .B(n880), .Z(n883) );
  AND U890 ( .A(n884), .B(n885), .Z(n654) );
  NOR U891 ( .A(n880), .B(n653), .Z(n882) );
  AND U892 ( .A(n886), .B(n887), .Z(n653) );
  XOR U893 ( .A(n888), .B(n889), .Z(n880) );
  AND U894 ( .A(n890), .B(n891), .Z(n889) );
  XNOR U895 ( .A(n888), .B(n886), .Z(n891) );
  IV U896 ( .A(n674), .Z(n886) );
  XOR U897 ( .A(n892), .B(n893), .Z(n674) );
  XOR U898 ( .A(n894), .B(n887), .Z(n893) );
  AND U899 ( .A(n702), .B(n895), .Z(n887) );
  AND U900 ( .A(n896), .B(n897), .Z(n894) );
  XOR U901 ( .A(n898), .B(n892), .Z(n896) );
  XNOR U902 ( .A(n671), .B(n888), .Z(n890) );
  XOR U903 ( .A(n899), .B(n900), .Z(n671) );
  AND U904 ( .A(n11), .B(n901), .Z(n900) );
  XOR U905 ( .A(n902), .B(n899), .Z(n901) );
  XOR U906 ( .A(n903), .B(n904), .Z(n888) );
  AND U907 ( .A(n905), .B(n906), .Z(n904) );
  XNOR U908 ( .A(n903), .B(n702), .Z(n906) );
  XOR U909 ( .A(n907), .B(n897), .Z(n702) );
  XNOR U910 ( .A(n908), .B(n892), .Z(n897) );
  XOR U911 ( .A(n909), .B(n910), .Z(n892) );
  AND U912 ( .A(n911), .B(n912), .Z(n910) );
  XOR U913 ( .A(n913), .B(n909), .Z(n911) );
  XNOR U914 ( .A(n914), .B(n915), .Z(n908) );
  AND U915 ( .A(n916), .B(n917), .Z(n915) );
  XOR U916 ( .A(n914), .B(n918), .Z(n916) );
  XNOR U917 ( .A(n898), .B(n895), .Z(n907) );
  AND U918 ( .A(n919), .B(n920), .Z(n895) );
  XOR U919 ( .A(n921), .B(n922), .Z(n898) );
  AND U920 ( .A(n923), .B(n924), .Z(n922) );
  XOR U921 ( .A(n921), .B(n925), .Z(n923) );
  XNOR U922 ( .A(n699), .B(n903), .Z(n905) );
  XOR U923 ( .A(n926), .B(n927), .Z(n699) );
  AND U924 ( .A(n11), .B(n928), .Z(n927) );
  XNOR U925 ( .A(n929), .B(n926), .Z(n928) );
  XOR U926 ( .A(n930), .B(n931), .Z(n903) );
  AND U927 ( .A(n932), .B(n933), .Z(n931) );
  XNOR U928 ( .A(n930), .B(n919), .Z(n933) );
  IV U929 ( .A(n752), .Z(n919) );
  XNOR U930 ( .A(n934), .B(n912), .Z(n752) );
  XNOR U931 ( .A(n935), .B(n918), .Z(n912) );
  XOR U932 ( .A(n936), .B(n937), .Z(n918) );
  AND U933 ( .A(n938), .B(n939), .Z(n937) );
  XOR U934 ( .A(n936), .B(n940), .Z(n938) );
  XNOR U935 ( .A(n917), .B(n909), .Z(n935) );
  XOR U936 ( .A(n941), .B(n942), .Z(n909) );
  AND U937 ( .A(n943), .B(n944), .Z(n942) );
  XNOR U938 ( .A(n945), .B(n941), .Z(n943) );
  XNOR U939 ( .A(n946), .B(n914), .Z(n917) );
  XOR U940 ( .A(n947), .B(n948), .Z(n914) );
  AND U941 ( .A(n949), .B(n950), .Z(n948) );
  XOR U942 ( .A(n947), .B(n951), .Z(n949) );
  XNOR U943 ( .A(n952), .B(n953), .Z(n946) );
  AND U944 ( .A(n954), .B(n955), .Z(n953) );
  XNOR U945 ( .A(n952), .B(n956), .Z(n954) );
  XNOR U946 ( .A(n913), .B(n920), .Z(n934) );
  AND U947 ( .A(n849), .B(n957), .Z(n920) );
  XOR U948 ( .A(n925), .B(n924), .Z(n913) );
  XNOR U949 ( .A(n958), .B(n921), .Z(n924) );
  XOR U950 ( .A(n959), .B(n960), .Z(n921) );
  AND U951 ( .A(n961), .B(n962), .Z(n960) );
  XOR U952 ( .A(n959), .B(n963), .Z(n961) );
  XNOR U953 ( .A(n964), .B(n965), .Z(n958) );
  AND U954 ( .A(n966), .B(n967), .Z(n965) );
  XOR U955 ( .A(n964), .B(n968), .Z(n966) );
  XOR U956 ( .A(n969), .B(n970), .Z(n925) );
  AND U957 ( .A(n971), .B(n972), .Z(n970) );
  XOR U958 ( .A(n969), .B(n973), .Z(n971) );
  XNOR U959 ( .A(n749), .B(n930), .Z(n932) );
  XOR U960 ( .A(n974), .B(n975), .Z(n749) );
  AND U961 ( .A(n11), .B(n976), .Z(n975) );
  XOR U962 ( .A(n977), .B(n974), .Z(n976) );
  XOR U963 ( .A(n978), .B(n979), .Z(n930) );
  AND U964 ( .A(n980), .B(n981), .Z(n979) );
  XNOR U965 ( .A(n978), .B(n849), .Z(n981) );
  XOR U966 ( .A(n982), .B(n944), .Z(n849) );
  XNOR U967 ( .A(n983), .B(n951), .Z(n944) );
  XOR U968 ( .A(n940), .B(n939), .Z(n951) );
  XNOR U969 ( .A(n984), .B(n936), .Z(n939) );
  XOR U970 ( .A(n985), .B(n986), .Z(n936) );
  AND U971 ( .A(n987), .B(n988), .Z(n986) );
  XOR U972 ( .A(n985), .B(n989), .Z(n987) );
  XNOR U973 ( .A(n990), .B(n991), .Z(n984) );
  NOR U974 ( .A(n992), .B(n993), .Z(n991) );
  XNOR U975 ( .A(n990), .B(n994), .Z(n992) );
  XOR U976 ( .A(n995), .B(n996), .Z(n940) );
  NOR U977 ( .A(n997), .B(n998), .Z(n996) );
  XNOR U978 ( .A(n995), .B(n999), .Z(n997) );
  XNOR U979 ( .A(n950), .B(n941), .Z(n983) );
  XOR U980 ( .A(n1000), .B(n1001), .Z(n941) );
  NOR U981 ( .A(n1002), .B(n1003), .Z(n1001) );
  XNOR U982 ( .A(n1000), .B(n1004), .Z(n1002) );
  XOR U983 ( .A(n1005), .B(n956), .Z(n950) );
  XNOR U984 ( .A(n1006), .B(n1007), .Z(n956) );
  NOR U985 ( .A(n1008), .B(n1009), .Z(n1007) );
  XNOR U986 ( .A(n1006), .B(n1010), .Z(n1008) );
  XNOR U987 ( .A(n955), .B(n947), .Z(n1005) );
  XOR U988 ( .A(n1011), .B(n1012), .Z(n947) );
  AND U989 ( .A(n1013), .B(n1014), .Z(n1012) );
  XOR U990 ( .A(n1011), .B(n1015), .Z(n1013) );
  XNOR U991 ( .A(n1016), .B(n952), .Z(n955) );
  XOR U992 ( .A(n1017), .B(n1018), .Z(n952) );
  AND U993 ( .A(n1019), .B(n1020), .Z(n1018) );
  XOR U994 ( .A(n1017), .B(n1021), .Z(n1019) );
  XNOR U995 ( .A(n1022), .B(n1023), .Z(n1016) );
  NOR U996 ( .A(n1024), .B(n1025), .Z(n1023) );
  XOR U997 ( .A(n1022), .B(n1026), .Z(n1024) );
  XOR U998 ( .A(n945), .B(n957), .Z(n982) );
  NOR U999 ( .A(n878), .B(n1027), .Z(n957) );
  XNOR U1000 ( .A(n963), .B(n962), .Z(n945) );
  XNOR U1001 ( .A(n1028), .B(n968), .Z(n962) );
  XOR U1002 ( .A(n1029), .B(n1030), .Z(n968) );
  NOR U1003 ( .A(n1031), .B(n1032), .Z(n1030) );
  XNOR U1004 ( .A(n1029), .B(n1033), .Z(n1031) );
  XNOR U1005 ( .A(n967), .B(n959), .Z(n1028) );
  XOR U1006 ( .A(n1034), .B(n1035), .Z(n959) );
  AND U1007 ( .A(n1036), .B(n1037), .Z(n1035) );
  XNOR U1008 ( .A(n1034), .B(n1038), .Z(n1036) );
  XNOR U1009 ( .A(n1039), .B(n964), .Z(n967) );
  XOR U1010 ( .A(n1040), .B(n1041), .Z(n964) );
  AND U1011 ( .A(n1042), .B(n1043), .Z(n1041) );
  XOR U1012 ( .A(n1040), .B(n1044), .Z(n1042) );
  XNOR U1013 ( .A(n1045), .B(n1046), .Z(n1039) );
  NOR U1014 ( .A(n1047), .B(n1048), .Z(n1046) );
  XOR U1015 ( .A(n1045), .B(n1049), .Z(n1047) );
  XOR U1016 ( .A(n973), .B(n972), .Z(n963) );
  XNOR U1017 ( .A(n1050), .B(n969), .Z(n972) );
  XOR U1018 ( .A(n1051), .B(n1052), .Z(n969) );
  AND U1019 ( .A(n1053), .B(n1054), .Z(n1052) );
  XOR U1020 ( .A(n1051), .B(n1055), .Z(n1053) );
  XNOR U1021 ( .A(n1056), .B(n1057), .Z(n1050) );
  NOR U1022 ( .A(n1058), .B(n1059), .Z(n1057) );
  XNOR U1023 ( .A(n1056), .B(n1060), .Z(n1058) );
  XOR U1024 ( .A(n1061), .B(n1062), .Z(n973) );
  NOR U1025 ( .A(n1063), .B(n1064), .Z(n1062) );
  XNOR U1026 ( .A(n1061), .B(n1065), .Z(n1063) );
  XNOR U1027 ( .A(n845), .B(n978), .Z(n980) );
  XOR U1028 ( .A(n1066), .B(n1067), .Z(n845) );
  AND U1029 ( .A(n11), .B(n1068), .Z(n1067) );
  XNOR U1030 ( .A(n1069), .B(n1066), .Z(n1068) );
  AND U1031 ( .A(n879), .B(n878), .Z(n978) );
  XOR U1032 ( .A(n1070), .B(n1027), .Z(n878) );
  XNOR U1033 ( .A(p_input[256]), .B(p_input[32]), .Z(n1027) );
  XOR U1034 ( .A(n1004), .B(n1003), .Z(n1070) );
  XOR U1035 ( .A(n1071), .B(n1015), .Z(n1003) );
  XOR U1036 ( .A(n989), .B(n988), .Z(n1015) );
  XNOR U1037 ( .A(n1072), .B(n994), .Z(n988) );
  XOR U1038 ( .A(p_input[280]), .B(p_input[56]), .Z(n994) );
  XOR U1039 ( .A(n985), .B(n993), .Z(n1072) );
  XOR U1040 ( .A(n1073), .B(n990), .Z(n993) );
  XOR U1041 ( .A(p_input[278]), .B(p_input[54]), .Z(n990) );
  XNOR U1042 ( .A(p_input[279]), .B(p_input[55]), .Z(n1073) );
  XNOR U1043 ( .A(n1074), .B(p_input[50]), .Z(n985) );
  XNOR U1044 ( .A(n999), .B(n998), .Z(n989) );
  XOR U1045 ( .A(n1075), .B(n995), .Z(n998) );
  XOR U1046 ( .A(p_input[275]), .B(p_input[51]), .Z(n995) );
  XNOR U1047 ( .A(p_input[276]), .B(p_input[52]), .Z(n1075) );
  XOR U1048 ( .A(p_input[277]), .B(p_input[53]), .Z(n999) );
  XNOR U1049 ( .A(n1014), .B(n1000), .Z(n1071) );
  XNOR U1050 ( .A(n1076), .B(p_input[33]), .Z(n1000) );
  XNOR U1051 ( .A(n1077), .B(n1021), .Z(n1014) );
  XNOR U1052 ( .A(n1010), .B(n1009), .Z(n1021) );
  XOR U1053 ( .A(n1078), .B(n1006), .Z(n1009) );
  XNOR U1054 ( .A(n1079), .B(p_input[58]), .Z(n1006) );
  XNOR U1055 ( .A(p_input[283]), .B(p_input[59]), .Z(n1078) );
  XOR U1056 ( .A(p_input[284]), .B(p_input[60]), .Z(n1010) );
  XNOR U1057 ( .A(n1020), .B(n1011), .Z(n1077) );
  XNOR U1058 ( .A(n1080), .B(p_input[49]), .Z(n1011) );
  XOR U1059 ( .A(n1081), .B(n1026), .Z(n1020) );
  XNOR U1060 ( .A(p_input[287]), .B(p_input[63]), .Z(n1026) );
  XOR U1061 ( .A(n1017), .B(n1025), .Z(n1081) );
  XOR U1062 ( .A(n1082), .B(n1022), .Z(n1025) );
  XOR U1063 ( .A(p_input[285]), .B(p_input[61]), .Z(n1022) );
  XNOR U1064 ( .A(p_input[286]), .B(p_input[62]), .Z(n1082) );
  XNOR U1065 ( .A(n1083), .B(p_input[57]), .Z(n1017) );
  XNOR U1066 ( .A(n1038), .B(n1037), .Z(n1004) );
  XNOR U1067 ( .A(n1084), .B(n1044), .Z(n1037) );
  XNOR U1068 ( .A(n1033), .B(n1032), .Z(n1044) );
  XOR U1069 ( .A(n1085), .B(n1029), .Z(n1032) );
  XNOR U1070 ( .A(n1086), .B(p_input[43]), .Z(n1029) );
  XNOR U1071 ( .A(p_input[268]), .B(p_input[44]), .Z(n1085) );
  XOR U1072 ( .A(p_input[269]), .B(p_input[45]), .Z(n1033) );
  XNOR U1073 ( .A(n1043), .B(n1034), .Z(n1084) );
  XOR U1074 ( .A(p_input[258]), .B(p_input[34]), .Z(n1034) );
  XOR U1075 ( .A(n1087), .B(n1049), .Z(n1043) );
  XNOR U1076 ( .A(p_input[272]), .B(p_input[48]), .Z(n1049) );
  XOR U1077 ( .A(n1040), .B(n1048), .Z(n1087) );
  XOR U1078 ( .A(n1088), .B(n1045), .Z(n1048) );
  XOR U1079 ( .A(p_input[270]), .B(p_input[46]), .Z(n1045) );
  XNOR U1080 ( .A(p_input[271]), .B(p_input[47]), .Z(n1088) );
  XNOR U1081 ( .A(n1089), .B(p_input[42]), .Z(n1040) );
  XNOR U1082 ( .A(n1055), .B(n1054), .Z(n1038) );
  XNOR U1083 ( .A(n1090), .B(n1060), .Z(n1054) );
  XOR U1084 ( .A(p_input[265]), .B(p_input[41]), .Z(n1060) );
  XOR U1085 ( .A(n1051), .B(n1059), .Z(n1090) );
  XOR U1086 ( .A(n1091), .B(n1056), .Z(n1059) );
  XOR U1087 ( .A(p_input[263]), .B(p_input[39]), .Z(n1056) );
  XNOR U1088 ( .A(p_input[264]), .B(p_input[40]), .Z(n1091) );
  XOR U1089 ( .A(p_input[259]), .B(p_input[35]), .Z(n1051) );
  XNOR U1090 ( .A(n1065), .B(n1064), .Z(n1055) );
  XOR U1091 ( .A(n1092), .B(n1061), .Z(n1064) );
  XOR U1092 ( .A(p_input[260]), .B(p_input[36]), .Z(n1061) );
  XNOR U1093 ( .A(p_input[261]), .B(p_input[37]), .Z(n1092) );
  XOR U1094 ( .A(p_input[262]), .B(p_input[38]), .Z(n1065) );
  IV U1095 ( .A(n875), .Z(n879) );
  XNOR U1096 ( .A(n1093), .B(n1094), .Z(n875) );
  AND U1097 ( .A(n11), .B(n1095), .Z(n1094) );
  XNOR U1098 ( .A(n1096), .B(n1093), .Z(n1095) );
  XNOR U1099 ( .A(n1097), .B(n1098), .Z(n11) );
  NOR U1100 ( .A(n1099), .B(n1100), .Z(n1098) );
  XOR U1101 ( .A(n885), .B(n1097), .Z(n1100) );
  AND U1102 ( .A(n1101), .B(n1102), .Z(n885) );
  NOR U1103 ( .A(n1097), .B(n884), .Z(n1099) );
  AND U1104 ( .A(n1103), .B(n1104), .Z(n884) );
  XOR U1105 ( .A(n1105), .B(n1106), .Z(n1097) );
  AND U1106 ( .A(n1107), .B(n1108), .Z(n1106) );
  XNOR U1107 ( .A(n1105), .B(n1103), .Z(n1108) );
  IV U1108 ( .A(n902), .Z(n1103) );
  XOR U1109 ( .A(n1109), .B(n1110), .Z(n902) );
  XOR U1110 ( .A(n1111), .B(n1104), .Z(n1110) );
  AND U1111 ( .A(n929), .B(n1112), .Z(n1104) );
  AND U1112 ( .A(n1113), .B(n1114), .Z(n1111) );
  XOR U1113 ( .A(n1115), .B(n1109), .Z(n1113) );
  XNOR U1114 ( .A(n899), .B(n1105), .Z(n1107) );
  XOR U1115 ( .A(n1116), .B(n1117), .Z(n899) );
  AND U1116 ( .A(n15), .B(n1118), .Z(n1117) );
  XOR U1117 ( .A(n1119), .B(n1116), .Z(n1118) );
  XOR U1118 ( .A(n1120), .B(n1121), .Z(n1105) );
  AND U1119 ( .A(n1122), .B(n1123), .Z(n1121) );
  XNOR U1120 ( .A(n1120), .B(n929), .Z(n1123) );
  XOR U1121 ( .A(n1124), .B(n1114), .Z(n929) );
  XNOR U1122 ( .A(n1125), .B(n1109), .Z(n1114) );
  XOR U1123 ( .A(n1126), .B(n1127), .Z(n1109) );
  AND U1124 ( .A(n1128), .B(n1129), .Z(n1127) );
  XOR U1125 ( .A(n1130), .B(n1126), .Z(n1128) );
  XNOR U1126 ( .A(n1131), .B(n1132), .Z(n1125) );
  AND U1127 ( .A(n1133), .B(n1134), .Z(n1132) );
  XOR U1128 ( .A(n1131), .B(n1135), .Z(n1133) );
  XNOR U1129 ( .A(n1115), .B(n1112), .Z(n1124) );
  AND U1130 ( .A(n1136), .B(n1137), .Z(n1112) );
  XOR U1131 ( .A(n1138), .B(n1139), .Z(n1115) );
  AND U1132 ( .A(n1140), .B(n1141), .Z(n1139) );
  XOR U1133 ( .A(n1138), .B(n1142), .Z(n1140) );
  XNOR U1134 ( .A(n926), .B(n1120), .Z(n1122) );
  XOR U1135 ( .A(n1143), .B(n1144), .Z(n926) );
  AND U1136 ( .A(n15), .B(n1145), .Z(n1144) );
  XNOR U1137 ( .A(n1146), .B(n1143), .Z(n1145) );
  XOR U1138 ( .A(n1147), .B(n1148), .Z(n1120) );
  AND U1139 ( .A(n1149), .B(n1150), .Z(n1148) );
  XNOR U1140 ( .A(n1147), .B(n1136), .Z(n1150) );
  IV U1141 ( .A(n977), .Z(n1136) );
  XNOR U1142 ( .A(n1151), .B(n1129), .Z(n977) );
  XNOR U1143 ( .A(n1152), .B(n1135), .Z(n1129) );
  XOR U1144 ( .A(n1153), .B(n1154), .Z(n1135) );
  AND U1145 ( .A(n1155), .B(n1156), .Z(n1154) );
  XOR U1146 ( .A(n1153), .B(n1157), .Z(n1155) );
  XNOR U1147 ( .A(n1134), .B(n1126), .Z(n1152) );
  XOR U1148 ( .A(n1158), .B(n1159), .Z(n1126) );
  AND U1149 ( .A(n1160), .B(n1161), .Z(n1159) );
  XNOR U1150 ( .A(n1162), .B(n1158), .Z(n1160) );
  XNOR U1151 ( .A(n1163), .B(n1131), .Z(n1134) );
  XOR U1152 ( .A(n1164), .B(n1165), .Z(n1131) );
  AND U1153 ( .A(n1166), .B(n1167), .Z(n1165) );
  XOR U1154 ( .A(n1164), .B(n1168), .Z(n1166) );
  XNOR U1155 ( .A(n1169), .B(n1170), .Z(n1163) );
  AND U1156 ( .A(n1171), .B(n1172), .Z(n1170) );
  XNOR U1157 ( .A(n1169), .B(n1173), .Z(n1171) );
  XNOR U1158 ( .A(n1130), .B(n1137), .Z(n1151) );
  AND U1159 ( .A(n1069), .B(n1174), .Z(n1137) );
  XOR U1160 ( .A(n1142), .B(n1141), .Z(n1130) );
  XNOR U1161 ( .A(n1175), .B(n1138), .Z(n1141) );
  XOR U1162 ( .A(n1176), .B(n1177), .Z(n1138) );
  AND U1163 ( .A(n1178), .B(n1179), .Z(n1177) );
  XOR U1164 ( .A(n1176), .B(n1180), .Z(n1178) );
  XNOR U1165 ( .A(n1181), .B(n1182), .Z(n1175) );
  AND U1166 ( .A(n1183), .B(n1184), .Z(n1182) );
  XOR U1167 ( .A(n1181), .B(n1185), .Z(n1183) );
  XOR U1168 ( .A(n1186), .B(n1187), .Z(n1142) );
  AND U1169 ( .A(n1188), .B(n1189), .Z(n1187) );
  XOR U1170 ( .A(n1186), .B(n1190), .Z(n1188) );
  XNOR U1171 ( .A(n974), .B(n1147), .Z(n1149) );
  XOR U1172 ( .A(n1191), .B(n1192), .Z(n974) );
  AND U1173 ( .A(n15), .B(n1193), .Z(n1192) );
  XOR U1174 ( .A(n1194), .B(n1191), .Z(n1193) );
  XOR U1175 ( .A(n1195), .B(n1196), .Z(n1147) );
  AND U1176 ( .A(n1197), .B(n1198), .Z(n1196) );
  XNOR U1177 ( .A(n1195), .B(n1069), .Z(n1198) );
  XOR U1178 ( .A(n1199), .B(n1161), .Z(n1069) );
  XNOR U1179 ( .A(n1200), .B(n1168), .Z(n1161) );
  XOR U1180 ( .A(n1157), .B(n1156), .Z(n1168) );
  XNOR U1181 ( .A(n1201), .B(n1153), .Z(n1156) );
  XOR U1182 ( .A(n1202), .B(n1203), .Z(n1153) );
  AND U1183 ( .A(n1204), .B(n1205), .Z(n1203) );
  XOR U1184 ( .A(n1202), .B(n1206), .Z(n1204) );
  XNOR U1185 ( .A(n1207), .B(n1208), .Z(n1201) );
  NOR U1186 ( .A(n1209), .B(n1210), .Z(n1208) );
  XNOR U1187 ( .A(n1207), .B(n1211), .Z(n1209) );
  XOR U1188 ( .A(n1212), .B(n1213), .Z(n1157) );
  NOR U1189 ( .A(n1214), .B(n1215), .Z(n1213) );
  XNOR U1190 ( .A(n1212), .B(n1216), .Z(n1214) );
  XNOR U1191 ( .A(n1167), .B(n1158), .Z(n1200) );
  XOR U1192 ( .A(n1217), .B(n1218), .Z(n1158) );
  NOR U1193 ( .A(n1219), .B(n1220), .Z(n1218) );
  XNOR U1194 ( .A(n1217), .B(n1221), .Z(n1219) );
  XOR U1195 ( .A(n1222), .B(n1173), .Z(n1167) );
  XNOR U1196 ( .A(n1223), .B(n1224), .Z(n1173) );
  NOR U1197 ( .A(n1225), .B(n1226), .Z(n1224) );
  XNOR U1198 ( .A(n1223), .B(n1227), .Z(n1225) );
  XNOR U1199 ( .A(n1172), .B(n1164), .Z(n1222) );
  XOR U1200 ( .A(n1228), .B(n1229), .Z(n1164) );
  AND U1201 ( .A(n1230), .B(n1231), .Z(n1229) );
  XOR U1202 ( .A(n1228), .B(n1232), .Z(n1230) );
  XNOR U1203 ( .A(n1233), .B(n1169), .Z(n1172) );
  XOR U1204 ( .A(n1234), .B(n1235), .Z(n1169) );
  AND U1205 ( .A(n1236), .B(n1237), .Z(n1235) );
  XOR U1206 ( .A(n1234), .B(n1238), .Z(n1236) );
  XNOR U1207 ( .A(n1239), .B(n1240), .Z(n1233) );
  NOR U1208 ( .A(n1241), .B(n1242), .Z(n1240) );
  XOR U1209 ( .A(n1239), .B(n1243), .Z(n1241) );
  XOR U1210 ( .A(n1162), .B(n1174), .Z(n1199) );
  NOR U1211 ( .A(n1096), .B(n1244), .Z(n1174) );
  XNOR U1212 ( .A(n1180), .B(n1179), .Z(n1162) );
  XNOR U1213 ( .A(n1245), .B(n1185), .Z(n1179) );
  XOR U1214 ( .A(n1246), .B(n1247), .Z(n1185) );
  NOR U1215 ( .A(n1248), .B(n1249), .Z(n1247) );
  XNOR U1216 ( .A(n1246), .B(n1250), .Z(n1248) );
  XNOR U1217 ( .A(n1184), .B(n1176), .Z(n1245) );
  XOR U1218 ( .A(n1251), .B(n1252), .Z(n1176) );
  AND U1219 ( .A(n1253), .B(n1254), .Z(n1252) );
  XNOR U1220 ( .A(n1251), .B(n1255), .Z(n1253) );
  XNOR U1221 ( .A(n1256), .B(n1181), .Z(n1184) );
  XOR U1222 ( .A(n1257), .B(n1258), .Z(n1181) );
  AND U1223 ( .A(n1259), .B(n1260), .Z(n1258) );
  XOR U1224 ( .A(n1257), .B(n1261), .Z(n1259) );
  XNOR U1225 ( .A(n1262), .B(n1263), .Z(n1256) );
  NOR U1226 ( .A(n1264), .B(n1265), .Z(n1263) );
  XOR U1227 ( .A(n1262), .B(n1266), .Z(n1264) );
  XOR U1228 ( .A(n1190), .B(n1189), .Z(n1180) );
  XNOR U1229 ( .A(n1267), .B(n1186), .Z(n1189) );
  XOR U1230 ( .A(n1268), .B(n1269), .Z(n1186) );
  AND U1231 ( .A(n1270), .B(n1271), .Z(n1269) );
  XOR U1232 ( .A(n1268), .B(n1272), .Z(n1270) );
  XNOR U1233 ( .A(n1273), .B(n1274), .Z(n1267) );
  NOR U1234 ( .A(n1275), .B(n1276), .Z(n1274) );
  XNOR U1235 ( .A(n1273), .B(n1277), .Z(n1275) );
  XOR U1236 ( .A(n1278), .B(n1279), .Z(n1190) );
  NOR U1237 ( .A(n1280), .B(n1281), .Z(n1279) );
  XNOR U1238 ( .A(n1278), .B(n1282), .Z(n1280) );
  XNOR U1239 ( .A(n1066), .B(n1195), .Z(n1197) );
  XOR U1240 ( .A(n1283), .B(n1284), .Z(n1066) );
  AND U1241 ( .A(n15), .B(n1285), .Z(n1284) );
  XNOR U1242 ( .A(n1286), .B(n1283), .Z(n1285) );
  AND U1243 ( .A(n1093), .B(n1096), .Z(n1195) );
  XOR U1244 ( .A(n1287), .B(n1244), .Z(n1096) );
  XNOR U1245 ( .A(p_input[256]), .B(p_input[64]), .Z(n1244) );
  XOR U1246 ( .A(n1221), .B(n1220), .Z(n1287) );
  XOR U1247 ( .A(n1288), .B(n1232), .Z(n1220) );
  XOR U1248 ( .A(n1206), .B(n1205), .Z(n1232) );
  XNOR U1249 ( .A(n1289), .B(n1211), .Z(n1205) );
  XOR U1250 ( .A(p_input[280]), .B(p_input[88]), .Z(n1211) );
  XOR U1251 ( .A(n1202), .B(n1210), .Z(n1289) );
  XOR U1252 ( .A(n1290), .B(n1207), .Z(n1210) );
  XOR U1253 ( .A(p_input[278]), .B(p_input[86]), .Z(n1207) );
  XNOR U1254 ( .A(p_input[279]), .B(p_input[87]), .Z(n1290) );
  XNOR U1255 ( .A(n1074), .B(p_input[82]), .Z(n1202) );
  XNOR U1256 ( .A(n1216), .B(n1215), .Z(n1206) );
  XOR U1257 ( .A(n1291), .B(n1212), .Z(n1215) );
  XOR U1258 ( .A(p_input[275]), .B(p_input[83]), .Z(n1212) );
  XNOR U1259 ( .A(p_input[276]), .B(p_input[84]), .Z(n1291) );
  XOR U1260 ( .A(p_input[277]), .B(p_input[85]), .Z(n1216) );
  XNOR U1261 ( .A(n1231), .B(n1217), .Z(n1288) );
  XNOR U1262 ( .A(n1076), .B(p_input[65]), .Z(n1217) );
  XNOR U1263 ( .A(n1292), .B(n1238), .Z(n1231) );
  XNOR U1264 ( .A(n1227), .B(n1226), .Z(n1238) );
  XOR U1265 ( .A(n1293), .B(n1223), .Z(n1226) );
  XNOR U1266 ( .A(n1079), .B(p_input[90]), .Z(n1223) );
  XNOR U1267 ( .A(p_input[283]), .B(p_input[91]), .Z(n1293) );
  XOR U1268 ( .A(p_input[284]), .B(p_input[92]), .Z(n1227) );
  XNOR U1269 ( .A(n1237), .B(n1228), .Z(n1292) );
  XNOR U1270 ( .A(n1080), .B(p_input[81]), .Z(n1228) );
  XOR U1271 ( .A(n1294), .B(n1243), .Z(n1237) );
  XNOR U1272 ( .A(p_input[287]), .B(p_input[95]), .Z(n1243) );
  XOR U1273 ( .A(n1234), .B(n1242), .Z(n1294) );
  XOR U1274 ( .A(n1295), .B(n1239), .Z(n1242) );
  XOR U1275 ( .A(p_input[285]), .B(p_input[93]), .Z(n1239) );
  XNOR U1276 ( .A(p_input[286]), .B(p_input[94]), .Z(n1295) );
  XNOR U1277 ( .A(n1083), .B(p_input[89]), .Z(n1234) );
  XNOR U1278 ( .A(n1255), .B(n1254), .Z(n1221) );
  XNOR U1279 ( .A(n1296), .B(n1261), .Z(n1254) );
  XNOR U1280 ( .A(n1250), .B(n1249), .Z(n1261) );
  XOR U1281 ( .A(n1297), .B(n1246), .Z(n1249) );
  XNOR U1282 ( .A(n1086), .B(p_input[75]), .Z(n1246) );
  XNOR U1283 ( .A(p_input[268]), .B(p_input[76]), .Z(n1297) );
  XOR U1284 ( .A(p_input[269]), .B(p_input[77]), .Z(n1250) );
  XNOR U1285 ( .A(n1260), .B(n1251), .Z(n1296) );
  XOR U1286 ( .A(p_input[258]), .B(p_input[66]), .Z(n1251) );
  XOR U1287 ( .A(n1298), .B(n1266), .Z(n1260) );
  XNOR U1288 ( .A(p_input[272]), .B(p_input[80]), .Z(n1266) );
  XOR U1289 ( .A(n1257), .B(n1265), .Z(n1298) );
  XOR U1290 ( .A(n1299), .B(n1262), .Z(n1265) );
  XOR U1291 ( .A(p_input[270]), .B(p_input[78]), .Z(n1262) );
  XNOR U1292 ( .A(p_input[271]), .B(p_input[79]), .Z(n1299) );
  XNOR U1293 ( .A(n1089), .B(p_input[74]), .Z(n1257) );
  XNOR U1294 ( .A(n1272), .B(n1271), .Z(n1255) );
  XNOR U1295 ( .A(n1300), .B(n1277), .Z(n1271) );
  XOR U1296 ( .A(p_input[265]), .B(p_input[73]), .Z(n1277) );
  XOR U1297 ( .A(n1268), .B(n1276), .Z(n1300) );
  XOR U1298 ( .A(n1301), .B(n1273), .Z(n1276) );
  XOR U1299 ( .A(p_input[263]), .B(p_input[71]), .Z(n1273) );
  XNOR U1300 ( .A(p_input[264]), .B(p_input[72]), .Z(n1301) );
  XOR U1301 ( .A(p_input[259]), .B(p_input[67]), .Z(n1268) );
  XNOR U1302 ( .A(n1282), .B(n1281), .Z(n1272) );
  XOR U1303 ( .A(n1302), .B(n1278), .Z(n1281) );
  XOR U1304 ( .A(p_input[260]), .B(p_input[68]), .Z(n1278) );
  XNOR U1305 ( .A(p_input[261]), .B(p_input[69]), .Z(n1302) );
  XOR U1306 ( .A(p_input[262]), .B(p_input[70]), .Z(n1282) );
  XOR U1307 ( .A(n1303), .B(n1304), .Z(n1093) );
  AND U1308 ( .A(n15), .B(n1305), .Z(n1304) );
  XNOR U1309 ( .A(n1306), .B(n1303), .Z(n1305) );
  XNOR U1310 ( .A(n1307), .B(n1308), .Z(n15) );
  NOR U1311 ( .A(n1309), .B(n1310), .Z(n1308) );
  XOR U1312 ( .A(n1102), .B(n1307), .Z(n1310) );
  AND U1313 ( .A(n1311), .B(n1312), .Z(n1102) );
  NOR U1314 ( .A(n1307), .B(n1101), .Z(n1309) );
  AND U1315 ( .A(n1313), .B(n1314), .Z(n1101) );
  XOR U1316 ( .A(n1315), .B(n1316), .Z(n1307) );
  AND U1317 ( .A(n1317), .B(n1318), .Z(n1316) );
  XNOR U1318 ( .A(n1315), .B(n1313), .Z(n1318) );
  IV U1319 ( .A(n1119), .Z(n1313) );
  XOR U1320 ( .A(n1319), .B(n1320), .Z(n1119) );
  XOR U1321 ( .A(n1321), .B(n1314), .Z(n1320) );
  AND U1322 ( .A(n1146), .B(n1322), .Z(n1314) );
  AND U1323 ( .A(n1323), .B(n1324), .Z(n1321) );
  XOR U1324 ( .A(n1325), .B(n1319), .Z(n1323) );
  XNOR U1325 ( .A(n1116), .B(n1315), .Z(n1317) );
  XOR U1326 ( .A(n1326), .B(n1327), .Z(n1116) );
  AND U1327 ( .A(n19), .B(n1328), .Z(n1327) );
  XOR U1328 ( .A(n1329), .B(n1326), .Z(n1328) );
  XOR U1329 ( .A(n1330), .B(n1331), .Z(n1315) );
  AND U1330 ( .A(n1332), .B(n1333), .Z(n1331) );
  XNOR U1331 ( .A(n1330), .B(n1146), .Z(n1333) );
  XOR U1332 ( .A(n1334), .B(n1324), .Z(n1146) );
  XNOR U1333 ( .A(n1335), .B(n1319), .Z(n1324) );
  XOR U1334 ( .A(n1336), .B(n1337), .Z(n1319) );
  AND U1335 ( .A(n1338), .B(n1339), .Z(n1337) );
  XOR U1336 ( .A(n1340), .B(n1336), .Z(n1338) );
  XNOR U1337 ( .A(n1341), .B(n1342), .Z(n1335) );
  AND U1338 ( .A(n1343), .B(n1344), .Z(n1342) );
  XOR U1339 ( .A(n1341), .B(n1345), .Z(n1343) );
  XNOR U1340 ( .A(n1325), .B(n1322), .Z(n1334) );
  AND U1341 ( .A(n1346), .B(n1347), .Z(n1322) );
  XOR U1342 ( .A(n1348), .B(n1349), .Z(n1325) );
  AND U1343 ( .A(n1350), .B(n1351), .Z(n1349) );
  XOR U1344 ( .A(n1348), .B(n1352), .Z(n1350) );
  XNOR U1345 ( .A(n1143), .B(n1330), .Z(n1332) );
  XOR U1346 ( .A(n1353), .B(n1354), .Z(n1143) );
  AND U1347 ( .A(n19), .B(n1355), .Z(n1354) );
  XNOR U1348 ( .A(n1356), .B(n1353), .Z(n1355) );
  XOR U1349 ( .A(n1357), .B(n1358), .Z(n1330) );
  AND U1350 ( .A(n1359), .B(n1360), .Z(n1358) );
  XNOR U1351 ( .A(n1357), .B(n1346), .Z(n1360) );
  IV U1352 ( .A(n1194), .Z(n1346) );
  XNOR U1353 ( .A(n1361), .B(n1339), .Z(n1194) );
  XNOR U1354 ( .A(n1362), .B(n1345), .Z(n1339) );
  XOR U1355 ( .A(n1363), .B(n1364), .Z(n1345) );
  AND U1356 ( .A(n1365), .B(n1366), .Z(n1364) );
  XOR U1357 ( .A(n1363), .B(n1367), .Z(n1365) );
  XNOR U1358 ( .A(n1344), .B(n1336), .Z(n1362) );
  XOR U1359 ( .A(n1368), .B(n1369), .Z(n1336) );
  AND U1360 ( .A(n1370), .B(n1371), .Z(n1369) );
  XNOR U1361 ( .A(n1372), .B(n1368), .Z(n1370) );
  XNOR U1362 ( .A(n1373), .B(n1341), .Z(n1344) );
  XOR U1363 ( .A(n1374), .B(n1375), .Z(n1341) );
  AND U1364 ( .A(n1376), .B(n1377), .Z(n1375) );
  XOR U1365 ( .A(n1374), .B(n1378), .Z(n1376) );
  XNOR U1366 ( .A(n1379), .B(n1380), .Z(n1373) );
  AND U1367 ( .A(n1381), .B(n1382), .Z(n1380) );
  XNOR U1368 ( .A(n1379), .B(n1383), .Z(n1381) );
  XNOR U1369 ( .A(n1340), .B(n1347), .Z(n1361) );
  AND U1370 ( .A(n1286), .B(n1384), .Z(n1347) );
  XOR U1371 ( .A(n1352), .B(n1351), .Z(n1340) );
  XNOR U1372 ( .A(n1385), .B(n1348), .Z(n1351) );
  XOR U1373 ( .A(n1386), .B(n1387), .Z(n1348) );
  AND U1374 ( .A(n1388), .B(n1389), .Z(n1387) );
  XOR U1375 ( .A(n1386), .B(n1390), .Z(n1388) );
  XNOR U1376 ( .A(n1391), .B(n1392), .Z(n1385) );
  AND U1377 ( .A(n1393), .B(n1394), .Z(n1392) );
  XOR U1378 ( .A(n1391), .B(n1395), .Z(n1393) );
  XOR U1379 ( .A(n1396), .B(n1397), .Z(n1352) );
  AND U1380 ( .A(n1398), .B(n1399), .Z(n1397) );
  XOR U1381 ( .A(n1396), .B(n1400), .Z(n1398) );
  XNOR U1382 ( .A(n1191), .B(n1357), .Z(n1359) );
  XOR U1383 ( .A(n1401), .B(n1402), .Z(n1191) );
  AND U1384 ( .A(n19), .B(n1403), .Z(n1402) );
  XOR U1385 ( .A(n1404), .B(n1401), .Z(n1403) );
  XOR U1386 ( .A(n1405), .B(n1406), .Z(n1357) );
  AND U1387 ( .A(n1407), .B(n1408), .Z(n1406) );
  XNOR U1388 ( .A(n1405), .B(n1286), .Z(n1408) );
  XOR U1389 ( .A(n1409), .B(n1371), .Z(n1286) );
  XNOR U1390 ( .A(n1410), .B(n1378), .Z(n1371) );
  XOR U1391 ( .A(n1367), .B(n1366), .Z(n1378) );
  XNOR U1392 ( .A(n1411), .B(n1363), .Z(n1366) );
  XOR U1393 ( .A(n1412), .B(n1413), .Z(n1363) );
  AND U1394 ( .A(n1414), .B(n1415), .Z(n1413) );
  XNOR U1395 ( .A(n1416), .B(n1417), .Z(n1414) );
  IV U1396 ( .A(n1412), .Z(n1416) );
  XNOR U1397 ( .A(n1418), .B(n1419), .Z(n1411) );
  NOR U1398 ( .A(n1420), .B(n1421), .Z(n1419) );
  XNOR U1399 ( .A(n1418), .B(n1422), .Z(n1420) );
  XOR U1400 ( .A(n1423), .B(n1424), .Z(n1367) );
  NOR U1401 ( .A(n1425), .B(n1426), .Z(n1424) );
  XNOR U1402 ( .A(n1423), .B(n1427), .Z(n1425) );
  XNOR U1403 ( .A(n1377), .B(n1368), .Z(n1410) );
  XOR U1404 ( .A(n1428), .B(n1429), .Z(n1368) );
  AND U1405 ( .A(n1430), .B(n1431), .Z(n1429) );
  XOR U1406 ( .A(n1428), .B(n1432), .Z(n1430) );
  XOR U1407 ( .A(n1433), .B(n1383), .Z(n1377) );
  XOR U1408 ( .A(n1434), .B(n1435), .Z(n1383) );
  NOR U1409 ( .A(n1436), .B(n1437), .Z(n1435) );
  XOR U1410 ( .A(n1434), .B(n1438), .Z(n1436) );
  XNOR U1411 ( .A(n1382), .B(n1374), .Z(n1433) );
  XOR U1412 ( .A(n1439), .B(n1440), .Z(n1374) );
  AND U1413 ( .A(n1441), .B(n1442), .Z(n1440) );
  XOR U1414 ( .A(n1439), .B(n1443), .Z(n1441) );
  XNOR U1415 ( .A(n1444), .B(n1379), .Z(n1382) );
  XNOR U1416 ( .A(n1445), .B(n1446), .Z(n1379) );
  NOR U1417 ( .A(n1447), .B(n1448), .Z(n1446) );
  XOR U1418 ( .A(n1445), .B(n1449), .Z(n1447) );
  XNOR U1419 ( .A(n1450), .B(n1451), .Z(n1444) );
  NOR U1420 ( .A(n1452), .B(n1453), .Z(n1451) );
  XNOR U1421 ( .A(n1450), .B(n1454), .Z(n1452) );
  XOR U1422 ( .A(n1372), .B(n1384), .Z(n1409) );
  NOR U1423 ( .A(n1306), .B(n1455), .Z(n1384) );
  XNOR U1424 ( .A(n1390), .B(n1389), .Z(n1372) );
  XNOR U1425 ( .A(n1456), .B(n1395), .Z(n1389) );
  XNOR U1426 ( .A(n1457), .B(n1458), .Z(n1395) );
  NOR U1427 ( .A(n1459), .B(n1460), .Z(n1458) );
  XOR U1428 ( .A(n1457), .B(n1461), .Z(n1459) );
  XNOR U1429 ( .A(n1394), .B(n1386), .Z(n1456) );
  XOR U1430 ( .A(n1462), .B(n1463), .Z(n1386) );
  AND U1431 ( .A(n1464), .B(n1465), .Z(n1463) );
  XOR U1432 ( .A(n1462), .B(n1466), .Z(n1464) );
  XNOR U1433 ( .A(n1467), .B(n1391), .Z(n1394) );
  XOR U1434 ( .A(n1468), .B(n1469), .Z(n1391) );
  AND U1435 ( .A(n1470), .B(n1471), .Z(n1469) );
  XNOR U1436 ( .A(n1472), .B(n1473), .Z(n1470) );
  IV U1437 ( .A(n1468), .Z(n1472) );
  XNOR U1438 ( .A(n1474), .B(n1475), .Z(n1467) );
  NOR U1439 ( .A(n1476), .B(n1477), .Z(n1475) );
  XNOR U1440 ( .A(n1474), .B(n1478), .Z(n1476) );
  XOR U1441 ( .A(n1400), .B(n1399), .Z(n1390) );
  XNOR U1442 ( .A(n1479), .B(n1396), .Z(n1399) );
  XOR U1443 ( .A(n1480), .B(n1481), .Z(n1396) );
  NOR U1444 ( .A(n1482), .B(n1483), .Z(n1481) );
  XNOR U1445 ( .A(n1480), .B(n1484), .Z(n1482) );
  XNOR U1446 ( .A(n1485), .B(n1486), .Z(n1479) );
  NOR U1447 ( .A(n1487), .B(n1488), .Z(n1486) );
  XNOR U1448 ( .A(n1485), .B(n1489), .Z(n1487) );
  XOR U1449 ( .A(n1490), .B(n1491), .Z(n1400) );
  NOR U1450 ( .A(n1492), .B(n1493), .Z(n1491) );
  XNOR U1451 ( .A(n1490), .B(n1494), .Z(n1492) );
  XNOR U1452 ( .A(n1283), .B(n1405), .Z(n1407) );
  XOR U1453 ( .A(n1495), .B(n1496), .Z(n1283) );
  AND U1454 ( .A(n19), .B(n1497), .Z(n1496) );
  XNOR U1455 ( .A(n1498), .B(n1495), .Z(n1497) );
  AND U1456 ( .A(n1303), .B(n1306), .Z(n1405) );
  XOR U1457 ( .A(n1499), .B(n1455), .Z(n1306) );
  XNOR U1458 ( .A(p_input[256]), .B(p_input[96]), .Z(n1455) );
  XNOR U1459 ( .A(n1432), .B(n1431), .Z(n1499) );
  XNOR U1460 ( .A(n1500), .B(n1443), .Z(n1431) );
  XOR U1461 ( .A(n1417), .B(n1415), .Z(n1443) );
  XNOR U1462 ( .A(n1501), .B(n1422), .Z(n1415) );
  XOR U1463 ( .A(p_input[120]), .B(p_input[280]), .Z(n1422) );
  XOR U1464 ( .A(n1412), .B(n1421), .Z(n1501) );
  XOR U1465 ( .A(n1502), .B(n1418), .Z(n1421) );
  XOR U1466 ( .A(p_input[118]), .B(p_input[278]), .Z(n1418) );
  XOR U1467 ( .A(p_input[119]), .B(n855), .Z(n1502) );
  XOR U1468 ( .A(p_input[114]), .B(p_input[274]), .Z(n1412) );
  XNOR U1469 ( .A(n1427), .B(n1426), .Z(n1417) );
  XOR U1470 ( .A(n1503), .B(n1423), .Z(n1426) );
  XOR U1471 ( .A(p_input[115]), .B(p_input[275]), .Z(n1423) );
  XOR U1472 ( .A(p_input[116]), .B(n857), .Z(n1503) );
  XOR U1473 ( .A(p_input[117]), .B(p_input[277]), .Z(n1427) );
  XNOR U1474 ( .A(n1442), .B(n1428), .Z(n1500) );
  XNOR U1475 ( .A(n1076), .B(p_input[97]), .Z(n1428) );
  XNOR U1476 ( .A(n1504), .B(n1449), .Z(n1442) );
  XNOR U1477 ( .A(n1438), .B(n1437), .Z(n1449) );
  XNOR U1478 ( .A(n1505), .B(n1434), .Z(n1437) );
  XNOR U1479 ( .A(p_input[122]), .B(p_input[282]), .Z(n1434) );
  XOR U1480 ( .A(p_input[123]), .B(n861), .Z(n1505) );
  XOR U1481 ( .A(p_input[124]), .B(p_input[284]), .Z(n1438) );
  XNOR U1482 ( .A(n1448), .B(n1506), .Z(n1504) );
  IV U1483 ( .A(n1439), .Z(n1506) );
  XOR U1484 ( .A(p_input[113]), .B(p_input[273]), .Z(n1439) );
  XOR U1485 ( .A(n1507), .B(n1454), .Z(n1448) );
  XNOR U1486 ( .A(p_input[127]), .B(n1508), .Z(n1454) );
  XNOR U1487 ( .A(n1445), .B(n1453), .Z(n1507) );
  XOR U1488 ( .A(n1509), .B(n1450), .Z(n1453) );
  XOR U1489 ( .A(p_input[125]), .B(p_input[285]), .Z(n1450) );
  XNOR U1490 ( .A(p_input[126]), .B(p_input[286]), .Z(n1509) );
  XNOR U1491 ( .A(p_input[121]), .B(p_input[281]), .Z(n1445) );
  XOR U1492 ( .A(n1466), .B(n1465), .Z(n1432) );
  XNOR U1493 ( .A(n1510), .B(n1473), .Z(n1465) );
  XNOR U1494 ( .A(n1461), .B(n1460), .Z(n1473) );
  XNOR U1495 ( .A(n1511), .B(n1457), .Z(n1460) );
  XNOR U1496 ( .A(p_input[107]), .B(p_input[267]), .Z(n1457) );
  XOR U1497 ( .A(p_input[108]), .B(n867), .Z(n1511) );
  XOR U1498 ( .A(p_input[109]), .B(p_input[269]), .Z(n1461) );
  XNOR U1499 ( .A(n1471), .B(n1462), .Z(n1510) );
  XOR U1500 ( .A(p_input[258]), .B(p_input[98]), .Z(n1462) );
  XNOR U1501 ( .A(n1512), .B(n1478), .Z(n1471) );
  XNOR U1502 ( .A(p_input[112]), .B(n869), .Z(n1478) );
  XOR U1503 ( .A(n1468), .B(n1477), .Z(n1512) );
  XOR U1504 ( .A(n1513), .B(n1474), .Z(n1477) );
  XOR U1505 ( .A(p_input[110]), .B(p_input[270]), .Z(n1474) );
  XOR U1506 ( .A(p_input[111]), .B(n871), .Z(n1513) );
  XOR U1507 ( .A(p_input[106]), .B(p_input[266]), .Z(n1468) );
  XNOR U1508 ( .A(n1484), .B(n1483), .Z(n1466) );
  XOR U1509 ( .A(n1514), .B(n1489), .Z(n1483) );
  XOR U1510 ( .A(p_input[105]), .B(p_input[265]), .Z(n1489) );
  XOR U1511 ( .A(n1480), .B(n1488), .Z(n1514) );
  XOR U1512 ( .A(n1515), .B(n1485), .Z(n1488) );
  XOR U1513 ( .A(p_input[103]), .B(p_input[263]), .Z(n1485) );
  XNOR U1514 ( .A(p_input[104]), .B(p_input[264]), .Z(n1515) );
  XOR U1515 ( .A(p_input[259]), .B(p_input[99]), .Z(n1480) );
  XNOR U1516 ( .A(n1494), .B(n1493), .Z(n1484) );
  XOR U1517 ( .A(n1516), .B(n1490), .Z(n1493) );
  XOR U1518 ( .A(p_input[100]), .B(p_input[260]), .Z(n1490) );
  XNOR U1519 ( .A(p_input[101]), .B(p_input[261]), .Z(n1516) );
  XOR U1520 ( .A(p_input[102]), .B(p_input[262]), .Z(n1494) );
  XOR U1521 ( .A(n1517), .B(n1518), .Z(n1303) );
  AND U1522 ( .A(n19), .B(n1519), .Z(n1518) );
  XNOR U1523 ( .A(n1520), .B(n1517), .Z(n1519) );
  XNOR U1524 ( .A(n1521), .B(n1522), .Z(n19) );
  NOR U1525 ( .A(n1523), .B(n1524), .Z(n1522) );
  XOR U1526 ( .A(n1312), .B(n1521), .Z(n1524) );
  AND U1527 ( .A(n1525), .B(n1526), .Z(n1312) );
  NOR U1528 ( .A(n1521), .B(n1311), .Z(n1523) );
  AND U1529 ( .A(n1527), .B(n1528), .Z(n1311) );
  XOR U1530 ( .A(n1529), .B(n1530), .Z(n1521) );
  AND U1531 ( .A(n1531), .B(n1532), .Z(n1530) );
  XNOR U1532 ( .A(n1529), .B(n1527), .Z(n1532) );
  IV U1533 ( .A(n1329), .Z(n1527) );
  XOR U1534 ( .A(n1533), .B(n1534), .Z(n1329) );
  XOR U1535 ( .A(n1535), .B(n1528), .Z(n1534) );
  AND U1536 ( .A(n1356), .B(n1536), .Z(n1528) );
  AND U1537 ( .A(n1537), .B(n1538), .Z(n1535) );
  XOR U1538 ( .A(n1539), .B(n1533), .Z(n1537) );
  XNOR U1539 ( .A(n1326), .B(n1529), .Z(n1531) );
  XOR U1540 ( .A(n1540), .B(n1541), .Z(n1326) );
  AND U1541 ( .A(n23), .B(n1542), .Z(n1541) );
  XOR U1542 ( .A(n1543), .B(n1540), .Z(n1542) );
  XOR U1543 ( .A(n1544), .B(n1545), .Z(n1529) );
  AND U1544 ( .A(n1546), .B(n1547), .Z(n1545) );
  XNOR U1545 ( .A(n1544), .B(n1356), .Z(n1547) );
  XOR U1546 ( .A(n1548), .B(n1538), .Z(n1356) );
  XNOR U1547 ( .A(n1549), .B(n1533), .Z(n1538) );
  XOR U1548 ( .A(n1550), .B(n1551), .Z(n1533) );
  AND U1549 ( .A(n1552), .B(n1553), .Z(n1551) );
  XOR U1550 ( .A(n1554), .B(n1550), .Z(n1552) );
  XNOR U1551 ( .A(n1555), .B(n1556), .Z(n1549) );
  AND U1552 ( .A(n1557), .B(n1558), .Z(n1556) );
  XOR U1553 ( .A(n1555), .B(n1559), .Z(n1557) );
  XNOR U1554 ( .A(n1539), .B(n1536), .Z(n1548) );
  AND U1555 ( .A(n1560), .B(n1561), .Z(n1536) );
  XOR U1556 ( .A(n1562), .B(n1563), .Z(n1539) );
  AND U1557 ( .A(n1564), .B(n1565), .Z(n1563) );
  XOR U1558 ( .A(n1562), .B(n1566), .Z(n1564) );
  XNOR U1559 ( .A(n1353), .B(n1544), .Z(n1546) );
  XOR U1560 ( .A(n1567), .B(n1568), .Z(n1353) );
  AND U1561 ( .A(n23), .B(n1569), .Z(n1568) );
  XNOR U1562 ( .A(n1570), .B(n1567), .Z(n1569) );
  XOR U1563 ( .A(n1571), .B(n1572), .Z(n1544) );
  AND U1564 ( .A(n1573), .B(n1574), .Z(n1572) );
  XNOR U1565 ( .A(n1571), .B(n1560), .Z(n1574) );
  IV U1566 ( .A(n1404), .Z(n1560) );
  XNOR U1567 ( .A(n1575), .B(n1553), .Z(n1404) );
  XNOR U1568 ( .A(n1576), .B(n1559), .Z(n1553) );
  XOR U1569 ( .A(n1577), .B(n1578), .Z(n1559) );
  AND U1570 ( .A(n1579), .B(n1580), .Z(n1578) );
  XOR U1571 ( .A(n1577), .B(n1581), .Z(n1579) );
  XNOR U1572 ( .A(n1558), .B(n1550), .Z(n1576) );
  XOR U1573 ( .A(n1582), .B(n1583), .Z(n1550) );
  AND U1574 ( .A(n1584), .B(n1585), .Z(n1583) );
  XNOR U1575 ( .A(n1586), .B(n1582), .Z(n1584) );
  XNOR U1576 ( .A(n1587), .B(n1555), .Z(n1558) );
  XOR U1577 ( .A(n1588), .B(n1589), .Z(n1555) );
  AND U1578 ( .A(n1590), .B(n1591), .Z(n1589) );
  XOR U1579 ( .A(n1588), .B(n1592), .Z(n1590) );
  XNOR U1580 ( .A(n1593), .B(n1594), .Z(n1587) );
  AND U1581 ( .A(n1595), .B(n1596), .Z(n1594) );
  XNOR U1582 ( .A(n1593), .B(n1597), .Z(n1595) );
  XNOR U1583 ( .A(n1554), .B(n1561), .Z(n1575) );
  AND U1584 ( .A(n1498), .B(n1598), .Z(n1561) );
  XOR U1585 ( .A(n1566), .B(n1565), .Z(n1554) );
  XNOR U1586 ( .A(n1599), .B(n1562), .Z(n1565) );
  XOR U1587 ( .A(n1600), .B(n1601), .Z(n1562) );
  AND U1588 ( .A(n1602), .B(n1603), .Z(n1601) );
  XOR U1589 ( .A(n1600), .B(n1604), .Z(n1602) );
  XNOR U1590 ( .A(n1605), .B(n1606), .Z(n1599) );
  AND U1591 ( .A(n1607), .B(n1608), .Z(n1606) );
  XOR U1592 ( .A(n1605), .B(n1609), .Z(n1607) );
  XOR U1593 ( .A(n1610), .B(n1611), .Z(n1566) );
  AND U1594 ( .A(n1612), .B(n1613), .Z(n1611) );
  XOR U1595 ( .A(n1610), .B(n1614), .Z(n1612) );
  XNOR U1596 ( .A(n1401), .B(n1571), .Z(n1573) );
  XOR U1597 ( .A(n1615), .B(n1616), .Z(n1401) );
  AND U1598 ( .A(n23), .B(n1617), .Z(n1616) );
  XOR U1599 ( .A(n1618), .B(n1615), .Z(n1617) );
  XOR U1600 ( .A(n1619), .B(n1620), .Z(n1571) );
  AND U1601 ( .A(n1621), .B(n1622), .Z(n1620) );
  XNOR U1602 ( .A(n1619), .B(n1498), .Z(n1622) );
  XOR U1603 ( .A(n1623), .B(n1585), .Z(n1498) );
  XNOR U1604 ( .A(n1624), .B(n1592), .Z(n1585) );
  XOR U1605 ( .A(n1581), .B(n1580), .Z(n1592) );
  XNOR U1606 ( .A(n1625), .B(n1577), .Z(n1580) );
  XOR U1607 ( .A(n1626), .B(n1627), .Z(n1577) );
  AND U1608 ( .A(n1628), .B(n1629), .Z(n1627) );
  XNOR U1609 ( .A(n1630), .B(n1631), .Z(n1628) );
  IV U1610 ( .A(n1626), .Z(n1630) );
  XNOR U1611 ( .A(n1632), .B(n1633), .Z(n1625) );
  NOR U1612 ( .A(n1634), .B(n1635), .Z(n1633) );
  XNOR U1613 ( .A(n1632), .B(n1636), .Z(n1634) );
  XOR U1614 ( .A(n1637), .B(n1638), .Z(n1581) );
  NOR U1615 ( .A(n1639), .B(n1640), .Z(n1638) );
  XNOR U1616 ( .A(n1637), .B(n1641), .Z(n1639) );
  XNOR U1617 ( .A(n1591), .B(n1582), .Z(n1624) );
  XOR U1618 ( .A(n1642), .B(n1643), .Z(n1582) );
  AND U1619 ( .A(n1644), .B(n1645), .Z(n1643) );
  XOR U1620 ( .A(n1642), .B(n1646), .Z(n1644) );
  XOR U1621 ( .A(n1647), .B(n1597), .Z(n1591) );
  XOR U1622 ( .A(n1648), .B(n1649), .Z(n1597) );
  NOR U1623 ( .A(n1650), .B(n1651), .Z(n1649) );
  XOR U1624 ( .A(n1648), .B(n1652), .Z(n1650) );
  XNOR U1625 ( .A(n1596), .B(n1588), .Z(n1647) );
  XOR U1626 ( .A(n1653), .B(n1654), .Z(n1588) );
  AND U1627 ( .A(n1655), .B(n1656), .Z(n1654) );
  XOR U1628 ( .A(n1653), .B(n1657), .Z(n1655) );
  XNOR U1629 ( .A(n1658), .B(n1593), .Z(n1596) );
  XOR U1630 ( .A(n1659), .B(n1660), .Z(n1593) );
  AND U1631 ( .A(n1661), .B(n1662), .Z(n1660) );
  XNOR U1632 ( .A(n1663), .B(n1664), .Z(n1661) );
  IV U1633 ( .A(n1659), .Z(n1663) );
  XNOR U1634 ( .A(n1665), .B(n1666), .Z(n1658) );
  NOR U1635 ( .A(n1667), .B(n1668), .Z(n1666) );
  XNOR U1636 ( .A(n1665), .B(n1669), .Z(n1667) );
  XOR U1637 ( .A(n1586), .B(n1598), .Z(n1623) );
  NOR U1638 ( .A(n1520), .B(n1670), .Z(n1598) );
  XNOR U1639 ( .A(n1604), .B(n1603), .Z(n1586) );
  XNOR U1640 ( .A(n1671), .B(n1609), .Z(n1603) );
  XNOR U1641 ( .A(n1672), .B(n1673), .Z(n1609) );
  NOR U1642 ( .A(n1674), .B(n1675), .Z(n1673) );
  XOR U1643 ( .A(n1672), .B(n1676), .Z(n1674) );
  XNOR U1644 ( .A(n1608), .B(n1600), .Z(n1671) );
  XOR U1645 ( .A(n1677), .B(n1678), .Z(n1600) );
  AND U1646 ( .A(n1679), .B(n1680), .Z(n1678) );
  XNOR U1647 ( .A(n1681), .B(n1682), .Z(n1679) );
  XNOR U1648 ( .A(n1683), .B(n1605), .Z(n1608) );
  XOR U1649 ( .A(n1684), .B(n1685), .Z(n1605) );
  AND U1650 ( .A(n1686), .B(n1687), .Z(n1685) );
  XNOR U1651 ( .A(n1688), .B(n1689), .Z(n1686) );
  IV U1652 ( .A(n1684), .Z(n1688) );
  XNOR U1653 ( .A(n1690), .B(n1691), .Z(n1683) );
  NOR U1654 ( .A(n1692), .B(n1693), .Z(n1691) );
  XNOR U1655 ( .A(n1690), .B(n1694), .Z(n1692) );
  XOR U1656 ( .A(n1614), .B(n1613), .Z(n1604) );
  XNOR U1657 ( .A(n1695), .B(n1610), .Z(n1613) );
  XOR U1658 ( .A(n1696), .B(n1697), .Z(n1610) );
  AND U1659 ( .A(n1698), .B(n1699), .Z(n1697) );
  XOR U1660 ( .A(n1696), .B(n1700), .Z(n1698) );
  XNOR U1661 ( .A(n1701), .B(n1702), .Z(n1695) );
  NOR U1662 ( .A(n1703), .B(n1704), .Z(n1702) );
  XNOR U1663 ( .A(n1701), .B(n1705), .Z(n1703) );
  XOR U1664 ( .A(n1706), .B(n1707), .Z(n1614) );
  NOR U1665 ( .A(n1708), .B(n1709), .Z(n1707) );
  XNOR U1666 ( .A(n1706), .B(n1710), .Z(n1708) );
  XNOR U1667 ( .A(n1495), .B(n1619), .Z(n1621) );
  XOR U1668 ( .A(n1711), .B(n1712), .Z(n1495) );
  AND U1669 ( .A(n23), .B(n1713), .Z(n1712) );
  XNOR U1670 ( .A(n1714), .B(n1711), .Z(n1713) );
  AND U1671 ( .A(n1517), .B(n1520), .Z(n1619) );
  XOR U1672 ( .A(n1715), .B(n1670), .Z(n1520) );
  XNOR U1673 ( .A(p_input[128]), .B(p_input[256]), .Z(n1670) );
  XNOR U1674 ( .A(n1646), .B(n1645), .Z(n1715) );
  XNOR U1675 ( .A(n1716), .B(n1657), .Z(n1645) );
  XOR U1676 ( .A(n1631), .B(n1629), .Z(n1657) );
  XNOR U1677 ( .A(n1717), .B(n1636), .Z(n1629) );
  XOR U1678 ( .A(p_input[152]), .B(p_input[280]), .Z(n1636) );
  XOR U1679 ( .A(n1626), .B(n1635), .Z(n1717) );
  XOR U1680 ( .A(n1718), .B(n1632), .Z(n1635) );
  XOR U1681 ( .A(p_input[150]), .B(p_input[278]), .Z(n1632) );
  XOR U1682 ( .A(p_input[151]), .B(n855), .Z(n1718) );
  XOR U1683 ( .A(p_input[146]), .B(p_input[274]), .Z(n1626) );
  XNOR U1684 ( .A(n1641), .B(n1640), .Z(n1631) );
  XOR U1685 ( .A(n1719), .B(n1637), .Z(n1640) );
  XOR U1686 ( .A(p_input[147]), .B(p_input[275]), .Z(n1637) );
  XOR U1687 ( .A(p_input[148]), .B(n857), .Z(n1719) );
  XOR U1688 ( .A(p_input[149]), .B(p_input[277]), .Z(n1641) );
  XOR U1689 ( .A(n1656), .B(n1720), .Z(n1716) );
  IV U1690 ( .A(n1642), .Z(n1720) );
  XOR U1691 ( .A(p_input[129]), .B(p_input[257]), .Z(n1642) );
  XNOR U1692 ( .A(n1721), .B(n1664), .Z(n1656) );
  XNOR U1693 ( .A(n1652), .B(n1651), .Z(n1664) );
  XNOR U1694 ( .A(n1722), .B(n1648), .Z(n1651) );
  XNOR U1695 ( .A(p_input[154]), .B(p_input[282]), .Z(n1648) );
  XOR U1696 ( .A(p_input[155]), .B(n861), .Z(n1722) );
  XOR U1697 ( .A(p_input[156]), .B(p_input[284]), .Z(n1652) );
  XOR U1698 ( .A(n1662), .B(n1723), .Z(n1721) );
  IV U1699 ( .A(n1653), .Z(n1723) );
  XOR U1700 ( .A(p_input[145]), .B(p_input[273]), .Z(n1653) );
  XNOR U1701 ( .A(n1724), .B(n1669), .Z(n1662) );
  XNOR U1702 ( .A(p_input[159]), .B(n1508), .Z(n1669) );
  XOR U1703 ( .A(n1659), .B(n1668), .Z(n1724) );
  XOR U1704 ( .A(n1725), .B(n1665), .Z(n1668) );
  XOR U1705 ( .A(p_input[157]), .B(p_input[285]), .Z(n1665) );
  XNOR U1706 ( .A(p_input[158]), .B(p_input[286]), .Z(n1725) );
  XOR U1707 ( .A(p_input[153]), .B(p_input[281]), .Z(n1659) );
  XOR U1708 ( .A(n1682), .B(n1680), .Z(n1646) );
  XNOR U1709 ( .A(n1726), .B(n1689), .Z(n1680) );
  XNOR U1710 ( .A(n1676), .B(n1675), .Z(n1689) );
  XNOR U1711 ( .A(n1727), .B(n1672), .Z(n1675) );
  XNOR U1712 ( .A(p_input[139]), .B(p_input[267]), .Z(n1672) );
  XOR U1713 ( .A(p_input[140]), .B(n867), .Z(n1727) );
  XOR U1714 ( .A(p_input[141]), .B(p_input[269]), .Z(n1676) );
  XOR U1715 ( .A(n1687), .B(n1681), .Z(n1726) );
  IV U1716 ( .A(n1677), .Z(n1681) );
  XOR U1717 ( .A(p_input[130]), .B(p_input[258]), .Z(n1677) );
  XNOR U1718 ( .A(n1728), .B(n1694), .Z(n1687) );
  XNOR U1719 ( .A(p_input[144]), .B(n869), .Z(n1694) );
  XOR U1720 ( .A(n1684), .B(n1693), .Z(n1728) );
  XOR U1721 ( .A(n1729), .B(n1690), .Z(n1693) );
  XOR U1722 ( .A(p_input[142]), .B(p_input[270]), .Z(n1690) );
  XOR U1723 ( .A(p_input[143]), .B(n871), .Z(n1729) );
  XOR U1724 ( .A(p_input[138]), .B(p_input[266]), .Z(n1684) );
  XOR U1725 ( .A(n1700), .B(n1699), .Z(n1682) );
  XNOR U1726 ( .A(n1730), .B(n1705), .Z(n1699) );
  XOR U1727 ( .A(p_input[137]), .B(p_input[265]), .Z(n1705) );
  XOR U1728 ( .A(n1696), .B(n1704), .Z(n1730) );
  XOR U1729 ( .A(n1731), .B(n1701), .Z(n1704) );
  XOR U1730 ( .A(p_input[135]), .B(p_input[263]), .Z(n1701) );
  XNOR U1731 ( .A(p_input[136]), .B(p_input[264]), .Z(n1731) );
  XOR U1732 ( .A(p_input[131]), .B(p_input[259]), .Z(n1696) );
  XNOR U1733 ( .A(n1710), .B(n1709), .Z(n1700) );
  XOR U1734 ( .A(n1732), .B(n1706), .Z(n1709) );
  XOR U1735 ( .A(p_input[132]), .B(p_input[260]), .Z(n1706) );
  XNOR U1736 ( .A(p_input[133]), .B(p_input[261]), .Z(n1732) );
  XOR U1737 ( .A(p_input[134]), .B(p_input[262]), .Z(n1710) );
  XOR U1738 ( .A(n1733), .B(n1734), .Z(n1517) );
  AND U1739 ( .A(n23), .B(n1735), .Z(n1734) );
  XNOR U1740 ( .A(n1736), .B(n1733), .Z(n1735) );
  XNOR U1741 ( .A(n1737), .B(n1738), .Z(n23) );
  NOR U1742 ( .A(n1739), .B(n1740), .Z(n1738) );
  XOR U1743 ( .A(n1526), .B(n1737), .Z(n1740) );
  AND U1744 ( .A(n1741), .B(n1742), .Z(n1526) );
  NOR U1745 ( .A(n1737), .B(n1525), .Z(n1739) );
  AND U1746 ( .A(n1743), .B(n1744), .Z(n1525) );
  XOR U1747 ( .A(n1745), .B(n1746), .Z(n1737) );
  AND U1748 ( .A(n1747), .B(n1748), .Z(n1746) );
  XNOR U1749 ( .A(n1745), .B(n1743), .Z(n1748) );
  IV U1750 ( .A(n1543), .Z(n1743) );
  XOR U1751 ( .A(n1749), .B(n1750), .Z(n1543) );
  XOR U1752 ( .A(n1751), .B(n1744), .Z(n1750) );
  AND U1753 ( .A(n1570), .B(n1752), .Z(n1744) );
  AND U1754 ( .A(n1753), .B(n1754), .Z(n1751) );
  XOR U1755 ( .A(n1755), .B(n1749), .Z(n1753) );
  XNOR U1756 ( .A(n1540), .B(n1745), .Z(n1747) );
  XNOR U1757 ( .A(n1756), .B(n1757), .Z(n1540) );
  AND U1758 ( .A(n26), .B(n1758), .Z(n1757) );
  XNOR U1759 ( .A(n1759), .B(n1756), .Z(n1758) );
  XOR U1760 ( .A(n1760), .B(n1761), .Z(n1745) );
  AND U1761 ( .A(n1762), .B(n1763), .Z(n1761) );
  XNOR U1762 ( .A(n1760), .B(n1570), .Z(n1763) );
  XOR U1763 ( .A(n1764), .B(n1754), .Z(n1570) );
  XNOR U1764 ( .A(n1765), .B(n1749), .Z(n1754) );
  XOR U1765 ( .A(n1766), .B(n1767), .Z(n1749) );
  AND U1766 ( .A(n1768), .B(n1769), .Z(n1767) );
  XOR U1767 ( .A(n1770), .B(n1766), .Z(n1768) );
  XNOR U1768 ( .A(n1771), .B(n1772), .Z(n1765) );
  AND U1769 ( .A(n1773), .B(n1774), .Z(n1772) );
  XOR U1770 ( .A(n1771), .B(n1775), .Z(n1773) );
  XNOR U1771 ( .A(n1755), .B(n1752), .Z(n1764) );
  AND U1772 ( .A(n1776), .B(n1777), .Z(n1752) );
  XOR U1773 ( .A(n1778), .B(n1779), .Z(n1755) );
  AND U1774 ( .A(n1780), .B(n1781), .Z(n1779) );
  XOR U1775 ( .A(n1778), .B(n1782), .Z(n1780) );
  XNOR U1776 ( .A(n1567), .B(n1760), .Z(n1762) );
  XNOR U1777 ( .A(n1783), .B(n1784), .Z(n1567) );
  AND U1778 ( .A(n26), .B(n1785), .Z(n1784) );
  XOR U1779 ( .A(n1786), .B(n1783), .Z(n1785) );
  XOR U1780 ( .A(n1787), .B(n1788), .Z(n1760) );
  AND U1781 ( .A(n1789), .B(n1790), .Z(n1788) );
  XNOR U1782 ( .A(n1787), .B(n1776), .Z(n1790) );
  IV U1783 ( .A(n1618), .Z(n1776) );
  XNOR U1784 ( .A(n1791), .B(n1769), .Z(n1618) );
  XNOR U1785 ( .A(n1792), .B(n1775), .Z(n1769) );
  XOR U1786 ( .A(n1793), .B(n1794), .Z(n1775) );
  AND U1787 ( .A(n1795), .B(n1796), .Z(n1794) );
  XOR U1788 ( .A(n1793), .B(n1797), .Z(n1795) );
  XNOR U1789 ( .A(n1774), .B(n1766), .Z(n1792) );
  XOR U1790 ( .A(n1798), .B(n1799), .Z(n1766) );
  AND U1791 ( .A(n1800), .B(n1801), .Z(n1799) );
  XNOR U1792 ( .A(n1802), .B(n1798), .Z(n1800) );
  XNOR U1793 ( .A(n1803), .B(n1771), .Z(n1774) );
  XOR U1794 ( .A(n1804), .B(n1805), .Z(n1771) );
  AND U1795 ( .A(n1806), .B(n1807), .Z(n1805) );
  XOR U1796 ( .A(n1804), .B(n1808), .Z(n1806) );
  XNOR U1797 ( .A(n1809), .B(n1810), .Z(n1803) );
  AND U1798 ( .A(n1811), .B(n1812), .Z(n1810) );
  XNOR U1799 ( .A(n1809), .B(n1813), .Z(n1811) );
  XNOR U1800 ( .A(n1770), .B(n1777), .Z(n1791) );
  AND U1801 ( .A(n1714), .B(n1814), .Z(n1777) );
  XOR U1802 ( .A(n1782), .B(n1781), .Z(n1770) );
  XNOR U1803 ( .A(n1815), .B(n1778), .Z(n1781) );
  XOR U1804 ( .A(n1816), .B(n1817), .Z(n1778) );
  AND U1805 ( .A(n1818), .B(n1819), .Z(n1817) );
  XOR U1806 ( .A(n1816), .B(n1820), .Z(n1818) );
  XNOR U1807 ( .A(n1821), .B(n1822), .Z(n1815) );
  AND U1808 ( .A(n1823), .B(n1824), .Z(n1822) );
  XOR U1809 ( .A(n1821), .B(n1825), .Z(n1823) );
  XOR U1810 ( .A(n1826), .B(n1827), .Z(n1782) );
  AND U1811 ( .A(n1828), .B(n1829), .Z(n1827) );
  XOR U1812 ( .A(n1826), .B(n1830), .Z(n1828) );
  XNOR U1813 ( .A(n1615), .B(n1787), .Z(n1789) );
  XNOR U1814 ( .A(n1831), .B(n1832), .Z(n1615) );
  AND U1815 ( .A(n26), .B(n1833), .Z(n1832) );
  XNOR U1816 ( .A(n1834), .B(n1831), .Z(n1833) );
  XOR U1817 ( .A(n1835), .B(n1836), .Z(n1787) );
  AND U1818 ( .A(n1837), .B(n1838), .Z(n1836) );
  XNOR U1819 ( .A(n1835), .B(n1714), .Z(n1838) );
  XOR U1820 ( .A(n1839), .B(n1801), .Z(n1714) );
  XNOR U1821 ( .A(n1840), .B(n1808), .Z(n1801) );
  XOR U1822 ( .A(n1797), .B(n1796), .Z(n1808) );
  XNOR U1823 ( .A(n1841), .B(n1793), .Z(n1796) );
  XOR U1824 ( .A(n1842), .B(n1843), .Z(n1793) );
  AND U1825 ( .A(n1844), .B(n1845), .Z(n1843) );
  XNOR U1826 ( .A(n1846), .B(n1847), .Z(n1844) );
  IV U1827 ( .A(n1842), .Z(n1846) );
  XNOR U1828 ( .A(n1848), .B(n1849), .Z(n1841) );
  NOR U1829 ( .A(n1850), .B(n1851), .Z(n1849) );
  XNOR U1830 ( .A(n1848), .B(n1852), .Z(n1850) );
  XOR U1831 ( .A(n1853), .B(n1854), .Z(n1797) );
  NOR U1832 ( .A(n1855), .B(n1856), .Z(n1854) );
  XNOR U1833 ( .A(n1853), .B(n1857), .Z(n1855) );
  XNOR U1834 ( .A(n1807), .B(n1798), .Z(n1840) );
  XOR U1835 ( .A(n1858), .B(n1859), .Z(n1798) );
  AND U1836 ( .A(n1860), .B(n1861), .Z(n1859) );
  XOR U1837 ( .A(n1858), .B(n1862), .Z(n1860) );
  XOR U1838 ( .A(n1863), .B(n1813), .Z(n1807) );
  XOR U1839 ( .A(n1864), .B(n1865), .Z(n1813) );
  NOR U1840 ( .A(n1866), .B(n1867), .Z(n1865) );
  XOR U1841 ( .A(n1864), .B(n1868), .Z(n1866) );
  XNOR U1842 ( .A(n1812), .B(n1804), .Z(n1863) );
  XOR U1843 ( .A(n1869), .B(n1870), .Z(n1804) );
  AND U1844 ( .A(n1871), .B(n1872), .Z(n1870) );
  XOR U1845 ( .A(n1869), .B(n1873), .Z(n1871) );
  XNOR U1846 ( .A(n1874), .B(n1809), .Z(n1812) );
  XOR U1847 ( .A(n1875), .B(n1876), .Z(n1809) );
  AND U1848 ( .A(n1877), .B(n1878), .Z(n1876) );
  XNOR U1849 ( .A(n1879), .B(n1880), .Z(n1877) );
  IV U1850 ( .A(n1875), .Z(n1879) );
  XNOR U1851 ( .A(n1881), .B(n1882), .Z(n1874) );
  NOR U1852 ( .A(n1883), .B(n1884), .Z(n1882) );
  XNOR U1853 ( .A(n1881), .B(n1885), .Z(n1883) );
  XOR U1854 ( .A(n1802), .B(n1814), .Z(n1839) );
  NOR U1855 ( .A(n1736), .B(n1886), .Z(n1814) );
  XNOR U1856 ( .A(n1820), .B(n1819), .Z(n1802) );
  XNOR U1857 ( .A(n1887), .B(n1825), .Z(n1819) );
  XNOR U1858 ( .A(n1888), .B(n1889), .Z(n1825) );
  NOR U1859 ( .A(n1890), .B(n1891), .Z(n1889) );
  XOR U1860 ( .A(n1888), .B(n1892), .Z(n1890) );
  XNOR U1861 ( .A(n1824), .B(n1816), .Z(n1887) );
  XOR U1862 ( .A(n1893), .B(n1894), .Z(n1816) );
  AND U1863 ( .A(n1895), .B(n1896), .Z(n1894) );
  XOR U1864 ( .A(n1893), .B(n1897), .Z(n1895) );
  XNOR U1865 ( .A(n1898), .B(n1821), .Z(n1824) );
  XOR U1866 ( .A(n1899), .B(n1900), .Z(n1821) );
  AND U1867 ( .A(n1901), .B(n1902), .Z(n1900) );
  XNOR U1868 ( .A(n1903), .B(n1904), .Z(n1901) );
  IV U1869 ( .A(n1899), .Z(n1903) );
  XNOR U1870 ( .A(n1905), .B(n1906), .Z(n1898) );
  NOR U1871 ( .A(n1907), .B(n1908), .Z(n1906) );
  XNOR U1872 ( .A(n1905), .B(n1909), .Z(n1907) );
  XOR U1873 ( .A(n1830), .B(n1829), .Z(n1820) );
  XNOR U1874 ( .A(n1910), .B(n1826), .Z(n1829) );
  XOR U1875 ( .A(n1911), .B(n1912), .Z(n1826) );
  AND U1876 ( .A(n1913), .B(n1914), .Z(n1912) );
  XNOR U1877 ( .A(n1915), .B(n1916), .Z(n1913) );
  XNOR U1878 ( .A(n1917), .B(n1918), .Z(n1910) );
  NOR U1879 ( .A(n1919), .B(n1920), .Z(n1918) );
  XNOR U1880 ( .A(n1917), .B(n1921), .Z(n1919) );
  XOR U1881 ( .A(n1922), .B(n1923), .Z(n1830) );
  NOR U1882 ( .A(n1924), .B(n1925), .Z(n1923) );
  XNOR U1883 ( .A(n1922), .B(n1926), .Z(n1924) );
  XNOR U1884 ( .A(n1711), .B(n1835), .Z(n1837) );
  XNOR U1885 ( .A(n1927), .B(n1928), .Z(n1711) );
  AND U1886 ( .A(n26), .B(n1929), .Z(n1928) );
  XOR U1887 ( .A(n1930), .B(n1927), .Z(n1929) );
  AND U1888 ( .A(n1733), .B(n1736), .Z(n1835) );
  XOR U1889 ( .A(n1931), .B(n1886), .Z(n1736) );
  XNOR U1890 ( .A(p_input[160]), .B(p_input[256]), .Z(n1886) );
  XNOR U1891 ( .A(n1862), .B(n1861), .Z(n1931) );
  XNOR U1892 ( .A(n1932), .B(n1873), .Z(n1861) );
  XOR U1893 ( .A(n1847), .B(n1845), .Z(n1873) );
  XNOR U1894 ( .A(n1933), .B(n1852), .Z(n1845) );
  XOR U1895 ( .A(p_input[184]), .B(p_input[280]), .Z(n1852) );
  XOR U1896 ( .A(n1842), .B(n1851), .Z(n1933) );
  XOR U1897 ( .A(n1934), .B(n1848), .Z(n1851) );
  XOR U1898 ( .A(p_input[182]), .B(p_input[278]), .Z(n1848) );
  XOR U1899 ( .A(p_input[183]), .B(n855), .Z(n1934) );
  XOR U1900 ( .A(p_input[178]), .B(p_input[274]), .Z(n1842) );
  XNOR U1901 ( .A(n1857), .B(n1856), .Z(n1847) );
  XOR U1902 ( .A(n1935), .B(n1853), .Z(n1856) );
  XOR U1903 ( .A(p_input[179]), .B(p_input[275]), .Z(n1853) );
  XOR U1904 ( .A(p_input[180]), .B(n857), .Z(n1935) );
  XOR U1905 ( .A(p_input[181]), .B(p_input[277]), .Z(n1857) );
  XOR U1906 ( .A(n1872), .B(n1936), .Z(n1932) );
  IV U1907 ( .A(n1858), .Z(n1936) );
  XOR U1908 ( .A(p_input[161]), .B(p_input[257]), .Z(n1858) );
  XNOR U1909 ( .A(n1937), .B(n1880), .Z(n1872) );
  XNOR U1910 ( .A(n1868), .B(n1867), .Z(n1880) );
  XNOR U1911 ( .A(n1938), .B(n1864), .Z(n1867) );
  XNOR U1912 ( .A(p_input[186]), .B(p_input[282]), .Z(n1864) );
  XOR U1913 ( .A(p_input[187]), .B(n861), .Z(n1938) );
  XOR U1914 ( .A(p_input[188]), .B(p_input[284]), .Z(n1868) );
  XOR U1915 ( .A(n1878), .B(n1939), .Z(n1937) );
  IV U1916 ( .A(n1869), .Z(n1939) );
  XOR U1917 ( .A(p_input[177]), .B(p_input[273]), .Z(n1869) );
  XNOR U1918 ( .A(n1940), .B(n1885), .Z(n1878) );
  XNOR U1919 ( .A(p_input[191]), .B(n1508), .Z(n1885) );
  XOR U1920 ( .A(n1875), .B(n1884), .Z(n1940) );
  XOR U1921 ( .A(n1941), .B(n1881), .Z(n1884) );
  XOR U1922 ( .A(p_input[189]), .B(p_input[285]), .Z(n1881) );
  XNOR U1923 ( .A(p_input[190]), .B(p_input[286]), .Z(n1941) );
  XOR U1924 ( .A(p_input[185]), .B(p_input[281]), .Z(n1875) );
  XOR U1925 ( .A(n1897), .B(n1896), .Z(n1862) );
  XNOR U1926 ( .A(n1942), .B(n1904), .Z(n1896) );
  XNOR U1927 ( .A(n1892), .B(n1891), .Z(n1904) );
  XNOR U1928 ( .A(n1943), .B(n1888), .Z(n1891) );
  XNOR U1929 ( .A(p_input[171]), .B(p_input[267]), .Z(n1888) );
  XOR U1930 ( .A(p_input[172]), .B(n867), .Z(n1943) );
  XOR U1931 ( .A(p_input[173]), .B(p_input[269]), .Z(n1892) );
  XNOR U1932 ( .A(n1902), .B(n1893), .Z(n1942) );
  XOR U1933 ( .A(p_input[162]), .B(p_input[258]), .Z(n1893) );
  XNOR U1934 ( .A(n1944), .B(n1909), .Z(n1902) );
  XNOR U1935 ( .A(p_input[176]), .B(n869), .Z(n1909) );
  XOR U1936 ( .A(n1899), .B(n1908), .Z(n1944) );
  XOR U1937 ( .A(n1945), .B(n1905), .Z(n1908) );
  XOR U1938 ( .A(p_input[174]), .B(p_input[270]), .Z(n1905) );
  XOR U1939 ( .A(p_input[175]), .B(n871), .Z(n1945) );
  XOR U1940 ( .A(p_input[170]), .B(p_input[266]), .Z(n1899) );
  XOR U1941 ( .A(n1916), .B(n1914), .Z(n1897) );
  XNOR U1942 ( .A(n1946), .B(n1921), .Z(n1914) );
  XOR U1943 ( .A(p_input[169]), .B(p_input[265]), .Z(n1921) );
  XOR U1944 ( .A(n1911), .B(n1920), .Z(n1946) );
  XOR U1945 ( .A(n1947), .B(n1917), .Z(n1920) );
  XOR U1946 ( .A(p_input[167]), .B(p_input[263]), .Z(n1917) );
  XNOR U1947 ( .A(p_input[168]), .B(p_input[264]), .Z(n1947) );
  IV U1948 ( .A(n1915), .Z(n1911) );
  XNOR U1949 ( .A(p_input[163]), .B(p_input[259]), .Z(n1915) );
  XNOR U1950 ( .A(n1926), .B(n1925), .Z(n1916) );
  XOR U1951 ( .A(n1948), .B(n1922), .Z(n1925) );
  XOR U1952 ( .A(p_input[164]), .B(p_input[260]), .Z(n1922) );
  XNOR U1953 ( .A(p_input[165]), .B(p_input[261]), .Z(n1948) );
  XOR U1954 ( .A(p_input[166]), .B(p_input[262]), .Z(n1926) );
  XOR U1955 ( .A(n1949), .B(n1950), .Z(n1733) );
  AND U1956 ( .A(n26), .B(n1951), .Z(n1950) );
  XNOR U1957 ( .A(n1952), .B(n1949), .Z(n1951) );
  XNOR U1958 ( .A(n1953), .B(n1954), .Z(n26) );
  MUX U1959 ( .IN0(n1741), .IN1(n1742), .SEL(n1953), .F(n1954) );
  AND U1960 ( .A(n1756), .B(n1955), .Z(n1742) );
  AND U1961 ( .A(n1956), .B(n1957), .Z(n1741) );
  XOR U1962 ( .A(n1958), .B(n1959), .Z(n1953) );
  AND U1963 ( .A(n1960), .B(n1961), .Z(n1959) );
  XNOR U1964 ( .A(n1958), .B(n1956), .Z(n1961) );
  IV U1965 ( .A(n1759), .Z(n1956) );
  XOR U1966 ( .A(n1962), .B(n1963), .Z(n1759) );
  XOR U1967 ( .A(n1964), .B(n1957), .Z(n1963) );
  AND U1968 ( .A(n1786), .B(n1965), .Z(n1957) );
  AND U1969 ( .A(n1966), .B(n1967), .Z(n1964) );
  XOR U1970 ( .A(n1968), .B(n1962), .Z(n1966) );
  XNOR U1971 ( .A(n1969), .B(n1958), .Z(n1960) );
  IV U1972 ( .A(n1756), .Z(n1969) );
  XNOR U1973 ( .A(n1970), .B(n1971), .Z(n1756) );
  XOR U1974 ( .A(n1972), .B(n1955), .Z(n1971) );
  AND U1975 ( .A(n1783), .B(n1973), .Z(n1955) );
  AND U1976 ( .A(n1974), .B(n1975), .Z(n1972) );
  XNOR U1977 ( .A(n1970), .B(n1976), .Z(n1974) );
  XOR U1978 ( .A(n1977), .B(n1978), .Z(n1958) );
  AND U1979 ( .A(n1979), .B(n1980), .Z(n1978) );
  XNOR U1980 ( .A(n1977), .B(n1786), .Z(n1980) );
  XOR U1981 ( .A(n1981), .B(n1967), .Z(n1786) );
  XNOR U1982 ( .A(n1982), .B(n1962), .Z(n1967) );
  XOR U1983 ( .A(n1983), .B(n1984), .Z(n1962) );
  AND U1984 ( .A(n1985), .B(n1986), .Z(n1984) );
  XOR U1985 ( .A(n1987), .B(n1983), .Z(n1985) );
  XNOR U1986 ( .A(n1988), .B(n1989), .Z(n1982) );
  AND U1987 ( .A(n1990), .B(n1991), .Z(n1989) );
  XOR U1988 ( .A(n1988), .B(n1992), .Z(n1990) );
  XNOR U1989 ( .A(n1968), .B(n1965), .Z(n1981) );
  AND U1990 ( .A(n1993), .B(n1994), .Z(n1965) );
  XOR U1991 ( .A(n1995), .B(n1996), .Z(n1968) );
  AND U1992 ( .A(n1997), .B(n1998), .Z(n1996) );
  XOR U1993 ( .A(n1995), .B(n1999), .Z(n1997) );
  XOR U1994 ( .A(n1783), .B(n1977), .Z(n1979) );
  XNOR U1995 ( .A(n2000), .B(n1976), .Z(n1783) );
  XNOR U1996 ( .A(n2001), .B(n2002), .Z(n1976) );
  AND U1997 ( .A(n2003), .B(n2004), .Z(n2002) );
  XOR U1998 ( .A(n2001), .B(n2005), .Z(n2003) );
  XNOR U1999 ( .A(n1975), .B(n1973), .Z(n2000) );
  AND U2000 ( .A(n1831), .B(n2006), .Z(n1973) );
  XNOR U2001 ( .A(n2007), .B(n1970), .Z(n1975) );
  XOR U2002 ( .A(n2008), .B(n2009), .Z(n1970) );
  AND U2003 ( .A(n2010), .B(n2011), .Z(n2009) );
  XOR U2004 ( .A(n2008), .B(n2012), .Z(n2010) );
  XNOR U2005 ( .A(n2013), .B(n2014), .Z(n2007) );
  AND U2006 ( .A(n2015), .B(n2016), .Z(n2014) );
  XNOR U2007 ( .A(n2013), .B(n2017), .Z(n2015) );
  XOR U2008 ( .A(n2018), .B(n2019), .Z(n1977) );
  AND U2009 ( .A(n2020), .B(n2021), .Z(n2019) );
  XNOR U2010 ( .A(n2018), .B(n1993), .Z(n2021) );
  IV U2011 ( .A(n1834), .Z(n1993) );
  XNOR U2012 ( .A(n2022), .B(n1986), .Z(n1834) );
  XNOR U2013 ( .A(n2023), .B(n1992), .Z(n1986) );
  XOR U2014 ( .A(n2024), .B(n2025), .Z(n1992) );
  AND U2015 ( .A(n2026), .B(n2027), .Z(n2025) );
  XOR U2016 ( .A(n2024), .B(n2028), .Z(n2026) );
  XNOR U2017 ( .A(n1991), .B(n1983), .Z(n2023) );
  XOR U2018 ( .A(n2029), .B(n2030), .Z(n1983) );
  AND U2019 ( .A(n2031), .B(n2032), .Z(n2030) );
  XNOR U2020 ( .A(n2033), .B(n2029), .Z(n2031) );
  XNOR U2021 ( .A(n2034), .B(n1988), .Z(n1991) );
  XOR U2022 ( .A(n2035), .B(n2036), .Z(n1988) );
  AND U2023 ( .A(n2037), .B(n2038), .Z(n2036) );
  XOR U2024 ( .A(n2035), .B(n2039), .Z(n2037) );
  XNOR U2025 ( .A(n2040), .B(n2041), .Z(n2034) );
  AND U2026 ( .A(n2042), .B(n2043), .Z(n2041) );
  XNOR U2027 ( .A(n2040), .B(n2044), .Z(n2042) );
  XNOR U2028 ( .A(n1987), .B(n1994), .Z(n2022) );
  AND U2029 ( .A(n1930), .B(n2045), .Z(n1994) );
  XOR U2030 ( .A(n1999), .B(n1998), .Z(n1987) );
  XNOR U2031 ( .A(n2046), .B(n1995), .Z(n1998) );
  XOR U2032 ( .A(n2047), .B(n2048), .Z(n1995) );
  AND U2033 ( .A(n2049), .B(n2050), .Z(n2048) );
  XOR U2034 ( .A(n2047), .B(n2051), .Z(n2049) );
  XNOR U2035 ( .A(n2052), .B(n2053), .Z(n2046) );
  AND U2036 ( .A(n2054), .B(n2055), .Z(n2053) );
  XOR U2037 ( .A(n2052), .B(n2056), .Z(n2054) );
  XOR U2038 ( .A(n2057), .B(n2058), .Z(n1999) );
  AND U2039 ( .A(n2059), .B(n2060), .Z(n2058) );
  XOR U2040 ( .A(n2057), .B(n2061), .Z(n2059) );
  XNOR U2041 ( .A(n2062), .B(n2018), .Z(n2020) );
  IV U2042 ( .A(n1831), .Z(n2062) );
  XOR U2043 ( .A(n2063), .B(n2012), .Z(n1831) );
  XOR U2044 ( .A(n2005), .B(n2004), .Z(n2012) );
  XNOR U2045 ( .A(n2064), .B(n2001), .Z(n2004) );
  XOR U2046 ( .A(n2065), .B(n2066), .Z(n2001) );
  AND U2047 ( .A(n2067), .B(n2068), .Z(n2066) );
  XOR U2048 ( .A(n2065), .B(n2069), .Z(n2067) );
  XNOR U2049 ( .A(n2070), .B(n2071), .Z(n2064) );
  AND U2050 ( .A(n2072), .B(n2073), .Z(n2071) );
  XOR U2051 ( .A(n2070), .B(n2074), .Z(n2072) );
  XOR U2052 ( .A(n2075), .B(n2076), .Z(n2005) );
  AND U2053 ( .A(n2077), .B(n2078), .Z(n2076) );
  XOR U2054 ( .A(n2075), .B(n2079), .Z(n2077) );
  XNOR U2055 ( .A(n2011), .B(n2006), .Z(n2063) );
  AND U2056 ( .A(n1927), .B(n2080), .Z(n2006) );
  XOR U2057 ( .A(n2081), .B(n2017), .Z(n2011) );
  XNOR U2058 ( .A(n2082), .B(n2083), .Z(n2017) );
  AND U2059 ( .A(n2084), .B(n2085), .Z(n2083) );
  XOR U2060 ( .A(n2082), .B(n2086), .Z(n2084) );
  XNOR U2061 ( .A(n2016), .B(n2008), .Z(n2081) );
  XOR U2062 ( .A(n2087), .B(n2088), .Z(n2008) );
  AND U2063 ( .A(n2089), .B(n2090), .Z(n2088) );
  XOR U2064 ( .A(n2087), .B(n2091), .Z(n2089) );
  XNOR U2065 ( .A(n2092), .B(n2013), .Z(n2016) );
  XOR U2066 ( .A(n2093), .B(n2094), .Z(n2013) );
  AND U2067 ( .A(n2095), .B(n2096), .Z(n2094) );
  XOR U2068 ( .A(n2093), .B(n2097), .Z(n2095) );
  XNOR U2069 ( .A(n2098), .B(n2099), .Z(n2092) );
  AND U2070 ( .A(n2100), .B(n2101), .Z(n2099) );
  XNOR U2071 ( .A(n2098), .B(n2102), .Z(n2100) );
  XOR U2072 ( .A(n2103), .B(n2104), .Z(n2018) );
  AND U2073 ( .A(n2105), .B(n2106), .Z(n2104) );
  XNOR U2074 ( .A(n2103), .B(n1930), .Z(n2106) );
  XOR U2075 ( .A(n2107), .B(n2032), .Z(n1930) );
  XNOR U2076 ( .A(n2108), .B(n2039), .Z(n2032) );
  XOR U2077 ( .A(n2028), .B(n2027), .Z(n2039) );
  XNOR U2078 ( .A(n2109), .B(n2024), .Z(n2027) );
  XOR U2079 ( .A(n2110), .B(n2111), .Z(n2024) );
  AND U2080 ( .A(n2112), .B(n2113), .Z(n2111) );
  XNOR U2081 ( .A(n2114), .B(n2115), .Z(n2112) );
  IV U2082 ( .A(n2110), .Z(n2114) );
  XNOR U2083 ( .A(n2116), .B(n2117), .Z(n2109) );
  NOR U2084 ( .A(n2118), .B(n2119), .Z(n2117) );
  XNOR U2085 ( .A(n2116), .B(n2120), .Z(n2118) );
  XOR U2086 ( .A(n2121), .B(n2122), .Z(n2028) );
  NOR U2087 ( .A(n2123), .B(n2124), .Z(n2122) );
  XNOR U2088 ( .A(n2121), .B(n2125), .Z(n2123) );
  XNOR U2089 ( .A(n2038), .B(n2029), .Z(n2108) );
  XOR U2090 ( .A(n2126), .B(n2127), .Z(n2029) );
  AND U2091 ( .A(n2128), .B(n2129), .Z(n2127) );
  XOR U2092 ( .A(n2126), .B(n2130), .Z(n2128) );
  XOR U2093 ( .A(n2131), .B(n2044), .Z(n2038) );
  XOR U2094 ( .A(n2132), .B(n2133), .Z(n2044) );
  NOR U2095 ( .A(n2134), .B(n2135), .Z(n2133) );
  XOR U2096 ( .A(n2132), .B(n2136), .Z(n2134) );
  XNOR U2097 ( .A(n2043), .B(n2035), .Z(n2131) );
  XOR U2098 ( .A(n2137), .B(n2138), .Z(n2035) );
  AND U2099 ( .A(n2139), .B(n2140), .Z(n2138) );
  XOR U2100 ( .A(n2137), .B(n2141), .Z(n2139) );
  XNOR U2101 ( .A(n2142), .B(n2040), .Z(n2043) );
  XOR U2102 ( .A(n2143), .B(n2144), .Z(n2040) );
  AND U2103 ( .A(n2145), .B(n2146), .Z(n2144) );
  XNOR U2104 ( .A(n2147), .B(n2148), .Z(n2145) );
  IV U2105 ( .A(n2143), .Z(n2147) );
  XNOR U2106 ( .A(n2149), .B(n2150), .Z(n2142) );
  NOR U2107 ( .A(n2151), .B(n2152), .Z(n2150) );
  XNOR U2108 ( .A(n2149), .B(n2153), .Z(n2151) );
  XOR U2109 ( .A(n2033), .B(n2045), .Z(n2107) );
  NOR U2110 ( .A(n1952), .B(n2154), .Z(n2045) );
  XNOR U2111 ( .A(n2051), .B(n2050), .Z(n2033) );
  XNOR U2112 ( .A(n2155), .B(n2056), .Z(n2050) );
  XNOR U2113 ( .A(n2156), .B(n2157), .Z(n2056) );
  NOR U2114 ( .A(n2158), .B(n2159), .Z(n2157) );
  XOR U2115 ( .A(n2156), .B(n2160), .Z(n2158) );
  XNOR U2116 ( .A(n2055), .B(n2047), .Z(n2155) );
  XOR U2117 ( .A(n2161), .B(n2162), .Z(n2047) );
  AND U2118 ( .A(n2163), .B(n2164), .Z(n2162) );
  XOR U2119 ( .A(n2161), .B(n2165), .Z(n2163) );
  XNOR U2120 ( .A(n2166), .B(n2052), .Z(n2055) );
  XOR U2121 ( .A(n2167), .B(n2168), .Z(n2052) );
  AND U2122 ( .A(n2169), .B(n2170), .Z(n2168) );
  XNOR U2123 ( .A(n2171), .B(n2172), .Z(n2169) );
  IV U2124 ( .A(n2167), .Z(n2171) );
  XNOR U2125 ( .A(n2173), .B(n2174), .Z(n2166) );
  NOR U2126 ( .A(n2175), .B(n2176), .Z(n2174) );
  XNOR U2127 ( .A(n2173), .B(n2177), .Z(n2175) );
  XOR U2128 ( .A(n2061), .B(n2060), .Z(n2051) );
  XNOR U2129 ( .A(n2178), .B(n2057), .Z(n2060) );
  XOR U2130 ( .A(n2179), .B(n2180), .Z(n2057) );
  AND U2131 ( .A(n2181), .B(n2182), .Z(n2180) );
  XNOR U2132 ( .A(n2183), .B(n2184), .Z(n2181) );
  XNOR U2133 ( .A(n2185), .B(n2186), .Z(n2178) );
  NOR U2134 ( .A(n2187), .B(n2188), .Z(n2186) );
  XNOR U2135 ( .A(n2185), .B(n2189), .Z(n2187) );
  XOR U2136 ( .A(n2190), .B(n2191), .Z(n2061) );
  NOR U2137 ( .A(n2192), .B(n2193), .Z(n2191) );
  XNOR U2138 ( .A(n2190), .B(n2194), .Z(n2192) );
  XNOR U2139 ( .A(n2195), .B(n2103), .Z(n2105) );
  IV U2140 ( .A(n1927), .Z(n2195) );
  XOR U2141 ( .A(n2196), .B(n2091), .Z(n1927) );
  XOR U2142 ( .A(n2069), .B(n2068), .Z(n2091) );
  XNOR U2143 ( .A(n2197), .B(n2074), .Z(n2068) );
  XOR U2144 ( .A(n2198), .B(n2199), .Z(n2074) );
  NOR U2145 ( .A(n2200), .B(n2201), .Z(n2199) );
  XNOR U2146 ( .A(n2198), .B(n2202), .Z(n2200) );
  XNOR U2147 ( .A(n2073), .B(n2065), .Z(n2197) );
  XOR U2148 ( .A(n2203), .B(n2204), .Z(n2065) );
  AND U2149 ( .A(n2205), .B(n2206), .Z(n2204) );
  XNOR U2150 ( .A(n2203), .B(n2207), .Z(n2205) );
  XNOR U2151 ( .A(n2208), .B(n2070), .Z(n2073) );
  XOR U2152 ( .A(n2209), .B(n2210), .Z(n2070) );
  AND U2153 ( .A(n2211), .B(n2212), .Z(n2210) );
  XOR U2154 ( .A(n2209), .B(n2213), .Z(n2211) );
  XNOR U2155 ( .A(n2214), .B(n2215), .Z(n2208) );
  NOR U2156 ( .A(n2216), .B(n2217), .Z(n2215) );
  XOR U2157 ( .A(n2214), .B(n2218), .Z(n2216) );
  XOR U2158 ( .A(n2079), .B(n2078), .Z(n2069) );
  XNOR U2159 ( .A(n2219), .B(n2075), .Z(n2078) );
  XOR U2160 ( .A(n2220), .B(n2221), .Z(n2075) );
  AND U2161 ( .A(n2222), .B(n2223), .Z(n2221) );
  XOR U2162 ( .A(n2220), .B(n2224), .Z(n2222) );
  XNOR U2163 ( .A(n2225), .B(n2226), .Z(n2219) );
  NOR U2164 ( .A(n2227), .B(n2228), .Z(n2226) );
  XNOR U2165 ( .A(n2225), .B(n2229), .Z(n2227) );
  XOR U2166 ( .A(n2230), .B(n2231), .Z(n2079) );
  NOR U2167 ( .A(n2232), .B(n2233), .Z(n2231) );
  XNOR U2168 ( .A(n2230), .B(n2234), .Z(n2232) );
  XNOR U2169 ( .A(n2090), .B(n2080), .Z(n2196) );
  AND U2170 ( .A(n1949), .B(n2235), .Z(n2080) );
  XNOR U2171 ( .A(n2236), .B(n2097), .Z(n2090) );
  XOR U2172 ( .A(n2086), .B(n2085), .Z(n2097) );
  XNOR U2173 ( .A(n2237), .B(n2082), .Z(n2085) );
  XOR U2174 ( .A(n2238), .B(n2239), .Z(n2082) );
  AND U2175 ( .A(n2240), .B(n2241), .Z(n2239) );
  XOR U2176 ( .A(n2238), .B(n2242), .Z(n2240) );
  XNOR U2177 ( .A(n2243), .B(n2244), .Z(n2237) );
  NOR U2178 ( .A(n2245), .B(n2246), .Z(n2244) );
  XNOR U2179 ( .A(n2243), .B(n2247), .Z(n2245) );
  XOR U2180 ( .A(n2248), .B(n2249), .Z(n2086) );
  NOR U2181 ( .A(n2250), .B(n2251), .Z(n2249) );
  XNOR U2182 ( .A(n2248), .B(n2252), .Z(n2250) );
  XNOR U2183 ( .A(n2096), .B(n2087), .Z(n2236) );
  XOR U2184 ( .A(n2253), .B(n2254), .Z(n2087) );
  NOR U2185 ( .A(n2255), .B(n2256), .Z(n2254) );
  XNOR U2186 ( .A(n2253), .B(n2257), .Z(n2255) );
  XOR U2187 ( .A(n2258), .B(n2102), .Z(n2096) );
  XNOR U2188 ( .A(n2259), .B(n2260), .Z(n2102) );
  NOR U2189 ( .A(n2261), .B(n2262), .Z(n2260) );
  XNOR U2190 ( .A(n2259), .B(n2263), .Z(n2261) );
  XNOR U2191 ( .A(n2101), .B(n2093), .Z(n2258) );
  XOR U2192 ( .A(n2264), .B(n2265), .Z(n2093) );
  AND U2193 ( .A(n2266), .B(n2267), .Z(n2265) );
  XOR U2194 ( .A(n2264), .B(n2268), .Z(n2266) );
  XNOR U2195 ( .A(n2269), .B(n2098), .Z(n2101) );
  XOR U2196 ( .A(n2270), .B(n2271), .Z(n2098) );
  AND U2197 ( .A(n2272), .B(n2273), .Z(n2271) );
  XOR U2198 ( .A(n2270), .B(n2274), .Z(n2272) );
  XNOR U2199 ( .A(n2275), .B(n2276), .Z(n2269) );
  NOR U2200 ( .A(n2277), .B(n2278), .Z(n2276) );
  XOR U2201 ( .A(n2275), .B(n2279), .Z(n2277) );
  AND U2202 ( .A(n1949), .B(n1952), .Z(n2103) );
  XOR U2203 ( .A(n2280), .B(n2154), .Z(n1952) );
  XNOR U2204 ( .A(p_input[192]), .B(p_input[256]), .Z(n2154) );
  XNOR U2205 ( .A(n2130), .B(n2129), .Z(n2280) );
  XNOR U2206 ( .A(n2281), .B(n2141), .Z(n2129) );
  XOR U2207 ( .A(n2115), .B(n2113), .Z(n2141) );
  XNOR U2208 ( .A(n2282), .B(n2120), .Z(n2113) );
  XOR U2209 ( .A(p_input[216]), .B(p_input[280]), .Z(n2120) );
  XOR U2210 ( .A(n2110), .B(n2119), .Z(n2282) );
  XOR U2211 ( .A(n2283), .B(n2116), .Z(n2119) );
  XOR U2212 ( .A(p_input[214]), .B(p_input[278]), .Z(n2116) );
  XOR U2213 ( .A(p_input[215]), .B(n855), .Z(n2283) );
  XOR U2214 ( .A(p_input[210]), .B(p_input[274]), .Z(n2110) );
  XNOR U2215 ( .A(n2125), .B(n2124), .Z(n2115) );
  XOR U2216 ( .A(n2284), .B(n2121), .Z(n2124) );
  XOR U2217 ( .A(p_input[211]), .B(p_input[275]), .Z(n2121) );
  XOR U2218 ( .A(p_input[212]), .B(n857), .Z(n2284) );
  XOR U2219 ( .A(p_input[213]), .B(p_input[277]), .Z(n2125) );
  XOR U2220 ( .A(n2140), .B(n2285), .Z(n2281) );
  IV U2221 ( .A(n2126), .Z(n2285) );
  XOR U2222 ( .A(p_input[193]), .B(p_input[257]), .Z(n2126) );
  XNOR U2223 ( .A(n2286), .B(n2148), .Z(n2140) );
  XNOR U2224 ( .A(n2136), .B(n2135), .Z(n2148) );
  XNOR U2225 ( .A(n2287), .B(n2132), .Z(n2135) );
  XNOR U2226 ( .A(p_input[218]), .B(p_input[282]), .Z(n2132) );
  XOR U2227 ( .A(p_input[219]), .B(n861), .Z(n2287) );
  XOR U2228 ( .A(p_input[220]), .B(p_input[284]), .Z(n2136) );
  XOR U2229 ( .A(n2146), .B(n2288), .Z(n2286) );
  IV U2230 ( .A(n2137), .Z(n2288) );
  XOR U2231 ( .A(p_input[209]), .B(p_input[273]), .Z(n2137) );
  XNOR U2232 ( .A(n2289), .B(n2153), .Z(n2146) );
  XNOR U2233 ( .A(p_input[223]), .B(n1508), .Z(n2153) );
  IV U2234 ( .A(p_input[287]), .Z(n1508) );
  XOR U2235 ( .A(n2143), .B(n2152), .Z(n2289) );
  XOR U2236 ( .A(n2290), .B(n2149), .Z(n2152) );
  XOR U2237 ( .A(p_input[221]), .B(p_input[285]), .Z(n2149) );
  XNOR U2238 ( .A(p_input[222]), .B(p_input[286]), .Z(n2290) );
  XOR U2239 ( .A(p_input[217]), .B(p_input[281]), .Z(n2143) );
  XOR U2240 ( .A(n2165), .B(n2164), .Z(n2130) );
  XNOR U2241 ( .A(n2291), .B(n2172), .Z(n2164) );
  XNOR U2242 ( .A(n2160), .B(n2159), .Z(n2172) );
  XNOR U2243 ( .A(n2292), .B(n2156), .Z(n2159) );
  XNOR U2244 ( .A(p_input[203]), .B(p_input[267]), .Z(n2156) );
  XOR U2245 ( .A(p_input[204]), .B(n867), .Z(n2292) );
  XOR U2246 ( .A(p_input[205]), .B(p_input[269]), .Z(n2160) );
  XNOR U2247 ( .A(n2170), .B(n2161), .Z(n2291) );
  XOR U2248 ( .A(p_input[194]), .B(p_input[258]), .Z(n2161) );
  XNOR U2249 ( .A(n2293), .B(n2177), .Z(n2170) );
  XNOR U2250 ( .A(p_input[208]), .B(n869), .Z(n2177) );
  IV U2251 ( .A(p_input[272]), .Z(n869) );
  XOR U2252 ( .A(n2167), .B(n2176), .Z(n2293) );
  XOR U2253 ( .A(n2294), .B(n2173), .Z(n2176) );
  XOR U2254 ( .A(p_input[206]), .B(p_input[270]), .Z(n2173) );
  XOR U2255 ( .A(p_input[207]), .B(n871), .Z(n2294) );
  XOR U2256 ( .A(p_input[202]), .B(p_input[266]), .Z(n2167) );
  XOR U2257 ( .A(n2184), .B(n2182), .Z(n2165) );
  XNOR U2258 ( .A(n2295), .B(n2189), .Z(n2182) );
  XOR U2259 ( .A(p_input[201]), .B(p_input[265]), .Z(n2189) );
  XOR U2260 ( .A(n2179), .B(n2188), .Z(n2295) );
  XOR U2261 ( .A(n2296), .B(n2185), .Z(n2188) );
  XOR U2262 ( .A(p_input[199]), .B(p_input[263]), .Z(n2185) );
  XNOR U2263 ( .A(p_input[200]), .B(p_input[264]), .Z(n2296) );
  IV U2264 ( .A(n2183), .Z(n2179) );
  XNOR U2265 ( .A(p_input[195]), .B(p_input[259]), .Z(n2183) );
  XNOR U2266 ( .A(n2194), .B(n2193), .Z(n2184) );
  XOR U2267 ( .A(n2297), .B(n2190), .Z(n2193) );
  XOR U2268 ( .A(p_input[196]), .B(p_input[260]), .Z(n2190) );
  XNOR U2269 ( .A(p_input[197]), .B(p_input[261]), .Z(n2297) );
  XOR U2270 ( .A(p_input[198]), .B(p_input[262]), .Z(n2194) );
  XOR U2271 ( .A(n2298), .B(n2257), .Z(n1949) );
  XNOR U2272 ( .A(n2207), .B(n2206), .Z(n2257) );
  XNOR U2273 ( .A(n2299), .B(n2213), .Z(n2206) );
  XNOR U2274 ( .A(n2202), .B(n2201), .Z(n2213) );
  XOR U2275 ( .A(n2300), .B(n2198), .Z(n2201) );
  XNOR U2276 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n1086), .Z(n2198) );
  IV U2277 ( .A(p_input[267]), .Z(n1086) );
  XOR U2278 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n867), .Z(n2300) );
  IV U2279 ( .A(p_input[268]), .Z(n867) );
  XOR U2280 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[269]), .Z(n2202)
         );
  XNOR U2281 ( .A(n2212), .B(n2203), .Z(n2299) );
  XOR U2282 ( .A(\knn_comb_/min_val_out[0][2] ), .B(p_input[258]), .Z(n2203)
         );
  XOR U2283 ( .A(n2301), .B(n2218), .Z(n2212) );
  XNOR U2284 ( .A(\knn_comb_/min_val_out[0][16] ), .B(p_input[272]), .Z(n2218)
         );
  XOR U2285 ( .A(n2209), .B(n2217), .Z(n2301) );
  XOR U2286 ( .A(n2302), .B(n2214), .Z(n2217) );
  XOR U2287 ( .A(\knn_comb_/min_val_out[0][14] ), .B(p_input[270]), .Z(n2214)
         );
  XOR U2288 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n871), .Z(n2302) );
  IV U2289 ( .A(p_input[271]), .Z(n871) );
  XNOR U2290 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n1089), .Z(n2209) );
  IV U2291 ( .A(p_input[266]), .Z(n1089) );
  XNOR U2292 ( .A(n2224), .B(n2223), .Z(n2207) );
  XNOR U2293 ( .A(n2303), .B(n2229), .Z(n2223) );
  XOR U2294 ( .A(\knn_comb_/min_val_out[0][9] ), .B(p_input[265]), .Z(n2229)
         );
  XOR U2295 ( .A(n2220), .B(n2228), .Z(n2303) );
  XOR U2296 ( .A(n2304), .B(n2225), .Z(n2228) );
  XOR U2297 ( .A(\knn_comb_/min_val_out[0][7] ), .B(p_input[263]), .Z(n2225)
         );
  XNOR U2298 ( .A(\knn_comb_/min_val_out[0][8] ), .B(p_input[264]), .Z(n2304)
         );
  XOR U2299 ( .A(\knn_comb_/min_val_out[0][3] ), .B(p_input[259]), .Z(n2220)
         );
  XNOR U2300 ( .A(n2234), .B(n2233), .Z(n2224) );
  XOR U2301 ( .A(n2305), .B(n2230), .Z(n2233) );
  XOR U2302 ( .A(\knn_comb_/min_val_out[0][4] ), .B(p_input[260]), .Z(n2230)
         );
  XNOR U2303 ( .A(\knn_comb_/min_val_out[0][5] ), .B(p_input[261]), .Z(n2305)
         );
  XOR U2304 ( .A(\knn_comb_/min_val_out[0][6] ), .B(p_input[262]), .Z(n2234)
         );
  XOR U2305 ( .A(n2256), .B(n2235), .Z(n2298) );
  XOR U2306 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[256]), .Z(n2235)
         );
  XOR U2307 ( .A(n2306), .B(n2268), .Z(n2256) );
  XOR U2308 ( .A(n2242), .B(n2241), .Z(n2268) );
  XNOR U2309 ( .A(n2307), .B(n2247), .Z(n2241) );
  XOR U2310 ( .A(\knn_comb_/min_val_out[0][24] ), .B(p_input[280]), .Z(n2247)
         );
  XOR U2311 ( .A(n2238), .B(n2246), .Z(n2307) );
  XOR U2312 ( .A(n2308), .B(n2243), .Z(n2246) );
  XOR U2313 ( .A(\knn_comb_/min_val_out[0][22] ), .B(p_input[278]), .Z(n2243)
         );
  XOR U2314 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n855), .Z(n2308) );
  IV U2315 ( .A(p_input[279]), .Z(n855) );
  XNOR U2316 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n1074), .Z(n2238) );
  IV U2317 ( .A(p_input[274]), .Z(n1074) );
  XNOR U2318 ( .A(n2252), .B(n2251), .Z(n2242) );
  XOR U2319 ( .A(n2309), .B(n2248), .Z(n2251) );
  XOR U2320 ( .A(\knn_comb_/min_val_out[0][19] ), .B(p_input[275]), .Z(n2248)
         );
  XOR U2321 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n857), .Z(n2309) );
  IV U2322 ( .A(p_input[276]), .Z(n857) );
  XOR U2323 ( .A(\knn_comb_/min_val_out[0][21] ), .B(p_input[277]), .Z(n2252)
         );
  XNOR U2324 ( .A(n2267), .B(n2253), .Z(n2306) );
  XNOR U2325 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n1076), .Z(n2253) );
  IV U2326 ( .A(p_input[257]), .Z(n1076) );
  XNOR U2327 ( .A(n2310), .B(n2274), .Z(n2267) );
  XNOR U2328 ( .A(n2263), .B(n2262), .Z(n2274) );
  XOR U2329 ( .A(n2311), .B(n2259), .Z(n2262) );
  XNOR U2330 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n1079), .Z(n2259) );
  IV U2331 ( .A(p_input[282]), .Z(n1079) );
  XOR U2332 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n861), .Z(n2311) );
  IV U2333 ( .A(p_input[283]), .Z(n861) );
  XOR U2334 ( .A(\knn_comb_/min_val_out[0][28] ), .B(p_input[284]), .Z(n2263)
         );
  XNOR U2335 ( .A(n2273), .B(n2264), .Z(n2310) );
  XNOR U2336 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n1080), .Z(n2264) );
  IV U2337 ( .A(p_input[273]), .Z(n1080) );
  XOR U2338 ( .A(n2312), .B(n2279), .Z(n2273) );
  XNOR U2339 ( .A(\knn_comb_/min_val_out[0][31] ), .B(p_input[287]), .Z(n2279)
         );
  XOR U2340 ( .A(n2270), .B(n2278), .Z(n2312) );
  XOR U2341 ( .A(n2313), .B(n2275), .Z(n2278) );
  XOR U2342 ( .A(\knn_comb_/min_val_out[0][29] ), .B(p_input[285]), .Z(n2275)
         );
  XNOR U2343 ( .A(\knn_comb_/min_val_out[0][30] ), .B(p_input[286]), .Z(n2313)
         );
  XNOR U2344 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n1083), .Z(n2270) );
  IV U2345 ( .A(p_input[281]), .Z(n1083) );
endmodule

