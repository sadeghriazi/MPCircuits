
module knn_comb_BMR_W32_K2_N8 ( p_input, o );
  input [287:0] p_input;
  output [63:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/min_val_out[0][16] , \knn_comb_/min_val_out[0][17] ,
         \knn_comb_/min_val_out[0][18] , \knn_comb_/min_val_out[0][19] ,
         \knn_comb_/min_val_out[0][20] , \knn_comb_/min_val_out[0][21] ,
         \knn_comb_/min_val_out[0][22] , \knn_comb_/min_val_out[0][23] ,
         \knn_comb_/min_val_out[0][24] , \knn_comb_/min_val_out[0][25] ,
         \knn_comb_/min_val_out[0][26] , \knn_comb_/min_val_out[0][27] ,
         \knn_comb_/min_val_out[0][28] , \knn_comb_/min_val_out[0][29] ,
         \knn_comb_/min_val_out[0][30] , \knn_comb_/min_val_out[0][31] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][31] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741;
  assign \knn_comb_/min_val_out[0][0]  = p_input[224];
  assign \knn_comb_/min_val_out[0][1]  = p_input[225];
  assign \knn_comb_/min_val_out[0][2]  = p_input[226];
  assign \knn_comb_/min_val_out[0][3]  = p_input[227];
  assign \knn_comb_/min_val_out[0][4]  = p_input[228];
  assign \knn_comb_/min_val_out[0][5]  = p_input[229];
  assign \knn_comb_/min_val_out[0][6]  = p_input[230];
  assign \knn_comb_/min_val_out[0][7]  = p_input[231];
  assign \knn_comb_/min_val_out[0][8]  = p_input[232];
  assign \knn_comb_/min_val_out[0][9]  = p_input[233];
  assign \knn_comb_/min_val_out[0][10]  = p_input[234];
  assign \knn_comb_/min_val_out[0][11]  = p_input[235];
  assign \knn_comb_/min_val_out[0][12]  = p_input[236];
  assign \knn_comb_/min_val_out[0][13]  = p_input[237];
  assign \knn_comb_/min_val_out[0][14]  = p_input[238];
  assign \knn_comb_/min_val_out[0][15]  = p_input[239];
  assign \knn_comb_/min_val_out[0][16]  = p_input[240];
  assign \knn_comb_/min_val_out[0][17]  = p_input[241];
  assign \knn_comb_/min_val_out[0][18]  = p_input[242];
  assign \knn_comb_/min_val_out[0][19]  = p_input[243];
  assign \knn_comb_/min_val_out[0][20]  = p_input[244];
  assign \knn_comb_/min_val_out[0][21]  = p_input[245];
  assign \knn_comb_/min_val_out[0][22]  = p_input[246];
  assign \knn_comb_/min_val_out[0][23]  = p_input[247];
  assign \knn_comb_/min_val_out[0][24]  = p_input[248];
  assign \knn_comb_/min_val_out[0][25]  = p_input[249];
  assign \knn_comb_/min_val_out[0][26]  = p_input[250];
  assign \knn_comb_/min_val_out[0][27]  = p_input[251];
  assign \knn_comb_/min_val_out[0][28]  = p_input[252];
  assign \knn_comb_/min_val_out[0][29]  = p_input[253];
  assign \knn_comb_/min_val_out[0][30]  = p_input[254];
  assign \knn_comb_/min_val_out[0][31]  = p_input[255];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][0]  = p_input[192];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][1]  = p_input[193];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][2]  = p_input[194];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][3]  = p_input[195];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][4]  = p_input[196];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][5]  = p_input[197];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][6]  = p_input[198];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][7]  = p_input[199];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][8]  = p_input[200];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][9]  = p_input[201];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][10]  = p_input[202];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][11]  = p_input[203];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][12]  = p_input[204];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][13]  = p_input[205];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][14]  = p_input[206];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][15]  = p_input[207];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][16]  = p_input[208];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][17]  = p_input[209];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][18]  = p_input[210];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][19]  = p_input[211];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][20]  = p_input[212];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][21]  = p_input[213];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][22]  = p_input[214];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][23]  = p_input[215];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][24]  = p_input[216];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][25]  = p_input[217];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][26]  = p_input[218];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][27]  = p_input[219];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][28]  = p_input[220];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][29]  = p_input[221];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][30]  = p_input[222];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][31]  = p_input[223];

  XOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  XOR U2 ( .A(n3), .B(n4), .Z(o[8]) );
  XOR U3 ( .A(n5), .B(n6), .Z(o[7]) );
  XOR U4 ( .A(n7), .B(n8), .Z(o[6]) );
  XOR U5 ( .A(n9), .B(n10), .Z(o[63]) );
  XOR U6 ( .A(n11), .B(n12), .Z(o[62]) );
  XOR U7 ( .A(n13), .B(n14), .Z(o[61]) );
  XOR U8 ( .A(n15), .B(n16), .Z(o[60]) );
  XOR U9 ( .A(n17), .B(n18), .Z(o[5]) );
  XOR U10 ( .A(n19), .B(n20), .Z(o[59]) );
  XOR U11 ( .A(n21), .B(n22), .Z(o[58]) );
  XOR U12 ( .A(n23), .B(n24), .Z(o[57]) );
  XOR U13 ( .A(n25), .B(n26), .Z(o[56]) );
  XOR U14 ( .A(n27), .B(n28), .Z(o[55]) );
  XOR U15 ( .A(n29), .B(n30), .Z(o[54]) );
  XOR U16 ( .A(n31), .B(n32), .Z(o[53]) );
  XOR U17 ( .A(n33), .B(n34), .Z(o[52]) );
  XOR U18 ( .A(n35), .B(n36), .Z(o[51]) );
  XOR U19 ( .A(n37), .B(n38), .Z(o[50]) );
  XOR U20 ( .A(n39), .B(n40), .Z(o[4]) );
  XOR U21 ( .A(n41), .B(n42), .Z(o[49]) );
  XOR U22 ( .A(n43), .B(n44), .Z(o[48]) );
  XOR U23 ( .A(n45), .B(n46), .Z(o[47]) );
  XOR U24 ( .A(n47), .B(n48), .Z(o[46]) );
  XOR U25 ( .A(n49), .B(n50), .Z(o[45]) );
  XOR U26 ( .A(n51), .B(n52), .Z(o[44]) );
  XOR U27 ( .A(n53), .B(n54), .Z(o[43]) );
  XOR U28 ( .A(n55), .B(n56), .Z(o[42]) );
  XOR U29 ( .A(n1), .B(n57), .Z(o[41]) );
  AND U30 ( .A(n58), .B(n59), .Z(n1) );
  XOR U31 ( .A(n2), .B(n57), .Z(n59) );
  XOR U32 ( .A(n60), .B(n61), .Z(n57) );
  AND U33 ( .A(n62), .B(n63), .Z(n61) );
  XOR U34 ( .A(p_input[9]), .B(n60), .Z(n63) );
  XOR U35 ( .A(n64), .B(n65), .Z(n60) );
  AND U36 ( .A(n66), .B(n67), .Z(n65) );
  XOR U37 ( .A(n68), .B(n69), .Z(n2) );
  AND U38 ( .A(n70), .B(n67), .Z(n69) );
  XNOR U39 ( .A(n71), .B(n64), .Z(n67) );
  XOR U40 ( .A(n72), .B(n73), .Z(n64) );
  AND U41 ( .A(n74), .B(n75), .Z(n73) );
  XOR U42 ( .A(p_input[41]), .B(n72), .Z(n75) );
  XOR U43 ( .A(n76), .B(n77), .Z(n72) );
  AND U44 ( .A(n78), .B(n79), .Z(n77) );
  IV U45 ( .A(n68), .Z(n71) );
  XNOR U46 ( .A(n80), .B(n81), .Z(n68) );
  AND U47 ( .A(n82), .B(n79), .Z(n81) );
  XNOR U48 ( .A(n80), .B(n76), .Z(n79) );
  XOR U49 ( .A(n83), .B(n84), .Z(n76) );
  AND U50 ( .A(n85), .B(n86), .Z(n84) );
  XOR U51 ( .A(p_input[73]), .B(n83), .Z(n86) );
  XOR U52 ( .A(n87), .B(n88), .Z(n83) );
  AND U53 ( .A(n89), .B(n90), .Z(n88) );
  XOR U54 ( .A(n91), .B(n92), .Z(n80) );
  AND U55 ( .A(n93), .B(n90), .Z(n92) );
  XNOR U56 ( .A(n91), .B(n87), .Z(n90) );
  XOR U57 ( .A(n94), .B(n95), .Z(n87) );
  AND U58 ( .A(n96), .B(n97), .Z(n95) );
  XOR U59 ( .A(p_input[105]), .B(n94), .Z(n97) );
  XOR U60 ( .A(n98), .B(n99), .Z(n94) );
  AND U61 ( .A(n100), .B(n101), .Z(n99) );
  XOR U62 ( .A(n102), .B(n103), .Z(n91) );
  AND U63 ( .A(n104), .B(n101), .Z(n103) );
  XNOR U64 ( .A(n102), .B(n98), .Z(n101) );
  XOR U65 ( .A(n105), .B(n106), .Z(n98) );
  AND U66 ( .A(n107), .B(n108), .Z(n106) );
  XOR U67 ( .A(p_input[137]), .B(n105), .Z(n108) );
  XOR U68 ( .A(n109), .B(n110), .Z(n105) );
  AND U69 ( .A(n111), .B(n112), .Z(n110) );
  XOR U70 ( .A(n113), .B(n114), .Z(n102) );
  AND U71 ( .A(n115), .B(n112), .Z(n114) );
  XNOR U72 ( .A(n113), .B(n109), .Z(n112) );
  XOR U73 ( .A(n116), .B(n117), .Z(n109) );
  AND U74 ( .A(n118), .B(n119), .Z(n117) );
  XOR U75 ( .A(p_input[169]), .B(n116), .Z(n119) );
  XNOR U76 ( .A(n120), .B(n121), .Z(n116) );
  AND U77 ( .A(n122), .B(n123), .Z(n121) );
  XNOR U78 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n124), .Z(n113) );
  AND U79 ( .A(n125), .B(n123), .Z(n124) );
  XOR U80 ( .A(n126), .B(n120), .Z(n123) );
  XOR U81 ( .A(n3), .B(n127), .Z(o[40]) );
  AND U82 ( .A(n58), .B(n128), .Z(n3) );
  XOR U83 ( .A(n4), .B(n127), .Z(n128) );
  XOR U84 ( .A(n129), .B(n130), .Z(n127) );
  AND U85 ( .A(n62), .B(n131), .Z(n130) );
  XOR U86 ( .A(p_input[8]), .B(n129), .Z(n131) );
  XOR U87 ( .A(n132), .B(n133), .Z(n129) );
  AND U88 ( .A(n66), .B(n134), .Z(n133) );
  XOR U89 ( .A(n135), .B(n136), .Z(n4) );
  AND U90 ( .A(n70), .B(n134), .Z(n136) );
  XNOR U91 ( .A(n137), .B(n132), .Z(n134) );
  XOR U92 ( .A(n138), .B(n139), .Z(n132) );
  AND U93 ( .A(n74), .B(n140), .Z(n139) );
  XOR U94 ( .A(p_input[40]), .B(n138), .Z(n140) );
  XOR U95 ( .A(n141), .B(n142), .Z(n138) );
  AND U96 ( .A(n78), .B(n143), .Z(n142) );
  IV U97 ( .A(n135), .Z(n137) );
  XNOR U98 ( .A(n144), .B(n145), .Z(n135) );
  AND U99 ( .A(n82), .B(n143), .Z(n145) );
  XNOR U100 ( .A(n144), .B(n141), .Z(n143) );
  XOR U101 ( .A(n146), .B(n147), .Z(n141) );
  AND U102 ( .A(n85), .B(n148), .Z(n147) );
  XOR U103 ( .A(p_input[72]), .B(n146), .Z(n148) );
  XOR U104 ( .A(n149), .B(n150), .Z(n146) );
  AND U105 ( .A(n89), .B(n151), .Z(n150) );
  XOR U106 ( .A(n152), .B(n153), .Z(n144) );
  AND U107 ( .A(n93), .B(n151), .Z(n153) );
  XNOR U108 ( .A(n152), .B(n149), .Z(n151) );
  XOR U109 ( .A(n154), .B(n155), .Z(n149) );
  AND U110 ( .A(n96), .B(n156), .Z(n155) );
  XOR U111 ( .A(p_input[104]), .B(n154), .Z(n156) );
  XOR U112 ( .A(n157), .B(n158), .Z(n154) );
  AND U113 ( .A(n100), .B(n159), .Z(n158) );
  XOR U114 ( .A(n160), .B(n161), .Z(n152) );
  AND U115 ( .A(n104), .B(n159), .Z(n161) );
  XNOR U116 ( .A(n160), .B(n157), .Z(n159) );
  XOR U117 ( .A(n162), .B(n163), .Z(n157) );
  AND U118 ( .A(n107), .B(n164), .Z(n163) );
  XOR U119 ( .A(p_input[136]), .B(n162), .Z(n164) );
  XOR U120 ( .A(n165), .B(n166), .Z(n162) );
  AND U121 ( .A(n111), .B(n167), .Z(n166) );
  XOR U122 ( .A(n168), .B(n169), .Z(n160) );
  AND U123 ( .A(n115), .B(n167), .Z(n169) );
  XNOR U124 ( .A(n168), .B(n165), .Z(n167) );
  XOR U125 ( .A(n170), .B(n171), .Z(n165) );
  AND U126 ( .A(n118), .B(n172), .Z(n171) );
  XOR U127 ( .A(p_input[168]), .B(n170), .Z(n172) );
  XNOR U128 ( .A(n173), .B(n174), .Z(n170) );
  AND U129 ( .A(n122), .B(n175), .Z(n174) );
  XNOR U130 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n176), .Z(n168) );
  AND U131 ( .A(n125), .B(n175), .Z(n176) );
  XOR U132 ( .A(n177), .B(n173), .Z(n175) );
  IV U133 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .Z(n173) );
  IV U134 ( .A(\knn_comb_/min_val_out[0][8] ), .Z(n177) );
  XOR U135 ( .A(n178), .B(n179), .Z(o[3]) );
  XOR U136 ( .A(n5), .B(n180), .Z(o[39]) );
  AND U137 ( .A(n58), .B(n181), .Z(n5) );
  XOR U138 ( .A(n6), .B(n180), .Z(n181) );
  XOR U139 ( .A(n182), .B(n183), .Z(n180) );
  AND U140 ( .A(n62), .B(n184), .Z(n183) );
  XOR U141 ( .A(p_input[7]), .B(n182), .Z(n184) );
  XOR U142 ( .A(n185), .B(n186), .Z(n182) );
  AND U143 ( .A(n66), .B(n187), .Z(n186) );
  XOR U144 ( .A(n188), .B(n189), .Z(n6) );
  AND U145 ( .A(n70), .B(n187), .Z(n189) );
  XNOR U146 ( .A(n190), .B(n185), .Z(n187) );
  XOR U147 ( .A(n191), .B(n192), .Z(n185) );
  AND U148 ( .A(n74), .B(n193), .Z(n192) );
  XOR U149 ( .A(p_input[39]), .B(n191), .Z(n193) );
  XOR U150 ( .A(n194), .B(n195), .Z(n191) );
  AND U151 ( .A(n78), .B(n196), .Z(n195) );
  IV U152 ( .A(n188), .Z(n190) );
  XNOR U153 ( .A(n197), .B(n198), .Z(n188) );
  AND U154 ( .A(n82), .B(n196), .Z(n198) );
  XNOR U155 ( .A(n197), .B(n194), .Z(n196) );
  XOR U156 ( .A(n199), .B(n200), .Z(n194) );
  AND U157 ( .A(n85), .B(n201), .Z(n200) );
  XOR U158 ( .A(p_input[71]), .B(n199), .Z(n201) );
  XOR U159 ( .A(n202), .B(n203), .Z(n199) );
  AND U160 ( .A(n89), .B(n204), .Z(n203) );
  XOR U161 ( .A(n205), .B(n206), .Z(n197) );
  AND U162 ( .A(n93), .B(n204), .Z(n206) );
  XNOR U163 ( .A(n205), .B(n202), .Z(n204) );
  XOR U164 ( .A(n207), .B(n208), .Z(n202) );
  AND U165 ( .A(n96), .B(n209), .Z(n208) );
  XOR U166 ( .A(p_input[103]), .B(n207), .Z(n209) );
  XOR U167 ( .A(n210), .B(n211), .Z(n207) );
  AND U168 ( .A(n100), .B(n212), .Z(n211) );
  XOR U169 ( .A(n213), .B(n214), .Z(n205) );
  AND U170 ( .A(n104), .B(n212), .Z(n214) );
  XNOR U171 ( .A(n213), .B(n210), .Z(n212) );
  XOR U172 ( .A(n215), .B(n216), .Z(n210) );
  AND U173 ( .A(n107), .B(n217), .Z(n216) );
  XOR U174 ( .A(p_input[135]), .B(n215), .Z(n217) );
  XOR U175 ( .A(n218), .B(n219), .Z(n215) );
  AND U176 ( .A(n111), .B(n220), .Z(n219) );
  XOR U177 ( .A(n221), .B(n222), .Z(n213) );
  AND U178 ( .A(n115), .B(n220), .Z(n222) );
  XNOR U179 ( .A(n221), .B(n218), .Z(n220) );
  XOR U180 ( .A(n223), .B(n224), .Z(n218) );
  AND U181 ( .A(n118), .B(n225), .Z(n224) );
  XOR U182 ( .A(p_input[167]), .B(n223), .Z(n225) );
  XNOR U183 ( .A(n226), .B(n227), .Z(n223) );
  AND U184 ( .A(n122), .B(n228), .Z(n227) );
  XNOR U185 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n229), .Z(n221) );
  AND U186 ( .A(n125), .B(n228), .Z(n229) );
  XOR U187 ( .A(n230), .B(n226), .Z(n228) );
  XOR U188 ( .A(n7), .B(n231), .Z(o[38]) );
  AND U189 ( .A(n58), .B(n232), .Z(n7) );
  XOR U190 ( .A(n8), .B(n231), .Z(n232) );
  XOR U191 ( .A(n233), .B(n234), .Z(n231) );
  AND U192 ( .A(n62), .B(n235), .Z(n234) );
  XOR U193 ( .A(p_input[6]), .B(n233), .Z(n235) );
  XOR U194 ( .A(n236), .B(n237), .Z(n233) );
  AND U195 ( .A(n66), .B(n238), .Z(n237) );
  XOR U196 ( .A(n239), .B(n240), .Z(n8) );
  AND U197 ( .A(n70), .B(n238), .Z(n240) );
  XNOR U198 ( .A(n241), .B(n236), .Z(n238) );
  XOR U199 ( .A(n242), .B(n243), .Z(n236) );
  AND U200 ( .A(n74), .B(n244), .Z(n243) );
  XOR U201 ( .A(p_input[38]), .B(n242), .Z(n244) );
  XOR U202 ( .A(n245), .B(n246), .Z(n242) );
  AND U203 ( .A(n78), .B(n247), .Z(n246) );
  IV U204 ( .A(n239), .Z(n241) );
  XNOR U205 ( .A(n248), .B(n249), .Z(n239) );
  AND U206 ( .A(n82), .B(n247), .Z(n249) );
  XNOR U207 ( .A(n248), .B(n245), .Z(n247) );
  XOR U208 ( .A(n250), .B(n251), .Z(n245) );
  AND U209 ( .A(n85), .B(n252), .Z(n251) );
  XOR U210 ( .A(p_input[70]), .B(n250), .Z(n252) );
  XOR U211 ( .A(n253), .B(n254), .Z(n250) );
  AND U212 ( .A(n89), .B(n255), .Z(n254) );
  XOR U213 ( .A(n256), .B(n257), .Z(n248) );
  AND U214 ( .A(n93), .B(n255), .Z(n257) );
  XNOR U215 ( .A(n256), .B(n253), .Z(n255) );
  XOR U216 ( .A(n258), .B(n259), .Z(n253) );
  AND U217 ( .A(n96), .B(n260), .Z(n259) );
  XOR U218 ( .A(p_input[102]), .B(n258), .Z(n260) );
  XOR U219 ( .A(n261), .B(n262), .Z(n258) );
  AND U220 ( .A(n100), .B(n263), .Z(n262) );
  XOR U221 ( .A(n264), .B(n265), .Z(n256) );
  AND U222 ( .A(n104), .B(n263), .Z(n265) );
  XNOR U223 ( .A(n264), .B(n261), .Z(n263) );
  XOR U224 ( .A(n266), .B(n267), .Z(n261) );
  AND U225 ( .A(n107), .B(n268), .Z(n267) );
  XOR U226 ( .A(p_input[134]), .B(n266), .Z(n268) );
  XOR U227 ( .A(n269), .B(n270), .Z(n266) );
  AND U228 ( .A(n111), .B(n271), .Z(n270) );
  XOR U229 ( .A(n272), .B(n273), .Z(n264) );
  AND U230 ( .A(n115), .B(n271), .Z(n273) );
  XNOR U231 ( .A(n272), .B(n269), .Z(n271) );
  XOR U232 ( .A(n274), .B(n275), .Z(n269) );
  AND U233 ( .A(n118), .B(n276), .Z(n275) );
  XOR U234 ( .A(p_input[166]), .B(n274), .Z(n276) );
  XNOR U235 ( .A(n277), .B(n278), .Z(n274) );
  AND U236 ( .A(n122), .B(n279), .Z(n278) );
  XNOR U237 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n280), .Z(n272) );
  AND U238 ( .A(n125), .B(n279), .Z(n280) );
  XOR U239 ( .A(n281), .B(n277), .Z(n279) );
  XOR U240 ( .A(n17), .B(n282), .Z(o[37]) );
  AND U241 ( .A(n58), .B(n283), .Z(n17) );
  XOR U242 ( .A(n18), .B(n282), .Z(n283) );
  XOR U243 ( .A(n284), .B(n285), .Z(n282) );
  AND U244 ( .A(n62), .B(n286), .Z(n285) );
  XOR U245 ( .A(p_input[5]), .B(n284), .Z(n286) );
  XOR U246 ( .A(n287), .B(n288), .Z(n284) );
  AND U247 ( .A(n66), .B(n289), .Z(n288) );
  XOR U248 ( .A(n290), .B(n291), .Z(n18) );
  AND U249 ( .A(n70), .B(n289), .Z(n291) );
  XNOR U250 ( .A(n292), .B(n287), .Z(n289) );
  XOR U251 ( .A(n293), .B(n294), .Z(n287) );
  AND U252 ( .A(n74), .B(n295), .Z(n294) );
  XOR U253 ( .A(p_input[37]), .B(n293), .Z(n295) );
  XOR U254 ( .A(n296), .B(n297), .Z(n293) );
  AND U255 ( .A(n78), .B(n298), .Z(n297) );
  IV U256 ( .A(n290), .Z(n292) );
  XNOR U257 ( .A(n299), .B(n300), .Z(n290) );
  AND U258 ( .A(n82), .B(n298), .Z(n300) );
  XNOR U259 ( .A(n299), .B(n296), .Z(n298) );
  XOR U260 ( .A(n301), .B(n302), .Z(n296) );
  AND U261 ( .A(n85), .B(n303), .Z(n302) );
  XOR U262 ( .A(p_input[69]), .B(n301), .Z(n303) );
  XOR U263 ( .A(n304), .B(n305), .Z(n301) );
  AND U264 ( .A(n89), .B(n306), .Z(n305) );
  XOR U265 ( .A(n307), .B(n308), .Z(n299) );
  AND U266 ( .A(n93), .B(n306), .Z(n308) );
  XNOR U267 ( .A(n307), .B(n304), .Z(n306) );
  XOR U268 ( .A(n309), .B(n310), .Z(n304) );
  AND U269 ( .A(n96), .B(n311), .Z(n310) );
  XOR U270 ( .A(p_input[101]), .B(n309), .Z(n311) );
  XOR U271 ( .A(n312), .B(n313), .Z(n309) );
  AND U272 ( .A(n100), .B(n314), .Z(n313) );
  XOR U273 ( .A(n315), .B(n316), .Z(n307) );
  AND U274 ( .A(n104), .B(n314), .Z(n316) );
  XNOR U275 ( .A(n315), .B(n312), .Z(n314) );
  XOR U276 ( .A(n317), .B(n318), .Z(n312) );
  AND U277 ( .A(n107), .B(n319), .Z(n318) );
  XOR U278 ( .A(p_input[133]), .B(n317), .Z(n319) );
  XOR U279 ( .A(n320), .B(n321), .Z(n317) );
  AND U280 ( .A(n111), .B(n322), .Z(n321) );
  XOR U281 ( .A(n323), .B(n324), .Z(n315) );
  AND U282 ( .A(n115), .B(n322), .Z(n324) );
  XNOR U283 ( .A(n323), .B(n320), .Z(n322) );
  XOR U284 ( .A(n325), .B(n326), .Z(n320) );
  AND U285 ( .A(n118), .B(n327), .Z(n326) );
  XOR U286 ( .A(p_input[165]), .B(n325), .Z(n327) );
  XNOR U287 ( .A(n328), .B(n329), .Z(n325) );
  AND U288 ( .A(n122), .B(n330), .Z(n329) );
  XNOR U289 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n331), .Z(n323) );
  AND U290 ( .A(n125), .B(n330), .Z(n331) );
  XOR U291 ( .A(n332), .B(n328), .Z(n330) );
  IV U292 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .Z(n328) );
  IV U293 ( .A(\knn_comb_/min_val_out[0][5] ), .Z(n332) );
  XOR U294 ( .A(n39), .B(n333), .Z(o[36]) );
  AND U295 ( .A(n58), .B(n334), .Z(n39) );
  XOR U296 ( .A(n40), .B(n333), .Z(n334) );
  XOR U297 ( .A(n335), .B(n336), .Z(n333) );
  AND U298 ( .A(n62), .B(n337), .Z(n336) );
  XOR U299 ( .A(p_input[4]), .B(n335), .Z(n337) );
  XOR U300 ( .A(n338), .B(n339), .Z(n335) );
  AND U301 ( .A(n66), .B(n340), .Z(n339) );
  XOR U302 ( .A(n341), .B(n342), .Z(n40) );
  AND U303 ( .A(n70), .B(n340), .Z(n342) );
  XNOR U304 ( .A(n343), .B(n338), .Z(n340) );
  XOR U305 ( .A(n344), .B(n345), .Z(n338) );
  AND U306 ( .A(n74), .B(n346), .Z(n345) );
  XOR U307 ( .A(p_input[36]), .B(n344), .Z(n346) );
  XOR U308 ( .A(n347), .B(n348), .Z(n344) );
  AND U309 ( .A(n78), .B(n349), .Z(n348) );
  IV U310 ( .A(n341), .Z(n343) );
  XNOR U311 ( .A(n350), .B(n351), .Z(n341) );
  AND U312 ( .A(n82), .B(n349), .Z(n351) );
  XNOR U313 ( .A(n350), .B(n347), .Z(n349) );
  XOR U314 ( .A(n352), .B(n353), .Z(n347) );
  AND U315 ( .A(n85), .B(n354), .Z(n353) );
  XOR U316 ( .A(p_input[68]), .B(n352), .Z(n354) );
  XOR U317 ( .A(n355), .B(n356), .Z(n352) );
  AND U318 ( .A(n89), .B(n357), .Z(n356) );
  XOR U319 ( .A(n358), .B(n359), .Z(n350) );
  AND U320 ( .A(n93), .B(n357), .Z(n359) );
  XNOR U321 ( .A(n358), .B(n355), .Z(n357) );
  XOR U322 ( .A(n360), .B(n361), .Z(n355) );
  AND U323 ( .A(n96), .B(n362), .Z(n361) );
  XOR U324 ( .A(p_input[100]), .B(n360), .Z(n362) );
  XOR U325 ( .A(n363), .B(n364), .Z(n360) );
  AND U326 ( .A(n100), .B(n365), .Z(n364) );
  XOR U327 ( .A(n366), .B(n367), .Z(n358) );
  AND U328 ( .A(n104), .B(n365), .Z(n367) );
  XNOR U329 ( .A(n366), .B(n363), .Z(n365) );
  XOR U330 ( .A(n368), .B(n369), .Z(n363) );
  AND U331 ( .A(n107), .B(n370), .Z(n369) );
  XOR U332 ( .A(p_input[132]), .B(n368), .Z(n370) );
  XOR U333 ( .A(n371), .B(n372), .Z(n368) );
  AND U334 ( .A(n111), .B(n373), .Z(n372) );
  XOR U335 ( .A(n374), .B(n375), .Z(n366) );
  AND U336 ( .A(n115), .B(n373), .Z(n375) );
  XNOR U337 ( .A(n374), .B(n371), .Z(n373) );
  XOR U338 ( .A(n376), .B(n377), .Z(n371) );
  AND U339 ( .A(n118), .B(n378), .Z(n377) );
  XOR U340 ( .A(p_input[164]), .B(n376), .Z(n378) );
  XNOR U341 ( .A(n379), .B(n380), .Z(n376) );
  AND U342 ( .A(n122), .B(n381), .Z(n380) );
  XNOR U343 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n382), .Z(n374) );
  AND U344 ( .A(n125), .B(n381), .Z(n382) );
  XOR U345 ( .A(n383), .B(n379), .Z(n381) );
  XOR U346 ( .A(n178), .B(n384), .Z(o[35]) );
  AND U347 ( .A(n58), .B(n385), .Z(n178) );
  XOR U348 ( .A(n179), .B(n384), .Z(n385) );
  XOR U349 ( .A(n386), .B(n387), .Z(n384) );
  AND U350 ( .A(n62), .B(n388), .Z(n387) );
  XOR U351 ( .A(p_input[3]), .B(n386), .Z(n388) );
  XOR U352 ( .A(n389), .B(n390), .Z(n386) );
  AND U353 ( .A(n66), .B(n391), .Z(n390) );
  XOR U354 ( .A(n392), .B(n393), .Z(n179) );
  AND U355 ( .A(n70), .B(n391), .Z(n393) );
  XNOR U356 ( .A(n394), .B(n389), .Z(n391) );
  XOR U357 ( .A(n395), .B(n396), .Z(n389) );
  AND U358 ( .A(n74), .B(n397), .Z(n396) );
  XOR U359 ( .A(p_input[35]), .B(n395), .Z(n397) );
  XOR U360 ( .A(n398), .B(n399), .Z(n395) );
  AND U361 ( .A(n78), .B(n400), .Z(n399) );
  IV U362 ( .A(n392), .Z(n394) );
  XNOR U363 ( .A(n401), .B(n402), .Z(n392) );
  AND U364 ( .A(n82), .B(n400), .Z(n402) );
  XNOR U365 ( .A(n401), .B(n398), .Z(n400) );
  XOR U366 ( .A(n403), .B(n404), .Z(n398) );
  AND U367 ( .A(n85), .B(n405), .Z(n404) );
  XOR U368 ( .A(p_input[67]), .B(n403), .Z(n405) );
  XOR U369 ( .A(n406), .B(n407), .Z(n403) );
  AND U370 ( .A(n89), .B(n408), .Z(n407) );
  XOR U371 ( .A(n409), .B(n410), .Z(n401) );
  AND U372 ( .A(n93), .B(n408), .Z(n410) );
  XNOR U373 ( .A(n409), .B(n406), .Z(n408) );
  XOR U374 ( .A(n411), .B(n412), .Z(n406) );
  AND U375 ( .A(n96), .B(n413), .Z(n412) );
  XOR U376 ( .A(p_input[99]), .B(n411), .Z(n413) );
  XOR U377 ( .A(n414), .B(n415), .Z(n411) );
  AND U378 ( .A(n100), .B(n416), .Z(n415) );
  XOR U379 ( .A(n417), .B(n418), .Z(n409) );
  AND U380 ( .A(n104), .B(n416), .Z(n418) );
  XNOR U381 ( .A(n417), .B(n414), .Z(n416) );
  XOR U382 ( .A(n419), .B(n420), .Z(n414) );
  AND U383 ( .A(n107), .B(n421), .Z(n420) );
  XOR U384 ( .A(p_input[131]), .B(n419), .Z(n421) );
  XOR U385 ( .A(n422), .B(n423), .Z(n419) );
  AND U386 ( .A(n111), .B(n424), .Z(n423) );
  XOR U387 ( .A(n425), .B(n426), .Z(n417) );
  AND U388 ( .A(n115), .B(n424), .Z(n426) );
  XNOR U389 ( .A(n425), .B(n422), .Z(n424) );
  XOR U390 ( .A(n427), .B(n428), .Z(n422) );
  AND U391 ( .A(n118), .B(n429), .Z(n428) );
  XOR U392 ( .A(p_input[163]), .B(n427), .Z(n429) );
  XNOR U393 ( .A(n430), .B(n431), .Z(n427) );
  AND U394 ( .A(n122), .B(n432), .Z(n431) );
  XNOR U395 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n433), .Z(n425) );
  AND U396 ( .A(n125), .B(n432), .Z(n433) );
  XOR U397 ( .A(n434), .B(n430), .Z(n432) );
  XOR U398 ( .A(n435), .B(n436), .Z(o[34]) );
  XOR U399 ( .A(n437), .B(n438), .Z(o[33]) );
  XOR U400 ( .A(n439), .B(n440), .Z(o[32]) );
  XOR U401 ( .A(n9), .B(n441), .Z(o[31]) );
  AND U402 ( .A(n58), .B(n442), .Z(n9) );
  XOR U403 ( .A(n10), .B(n441), .Z(n442) );
  XOR U404 ( .A(n443), .B(n444), .Z(n441) );
  AND U405 ( .A(n70), .B(n445), .Z(n444) );
  XOR U406 ( .A(n446), .B(n447), .Z(n10) );
  AND U407 ( .A(n62), .B(n448), .Z(n447) );
  XOR U408 ( .A(p_input[31]), .B(n446), .Z(n448) );
  XNOR U409 ( .A(n449), .B(n450), .Z(n446) );
  AND U410 ( .A(n66), .B(n445), .Z(n450) );
  XNOR U411 ( .A(n449), .B(n443), .Z(n445) );
  XOR U412 ( .A(n451), .B(n452), .Z(n443) );
  AND U413 ( .A(n82), .B(n453), .Z(n452) );
  XNOR U414 ( .A(n454), .B(n455), .Z(n449) );
  AND U415 ( .A(n74), .B(n456), .Z(n455) );
  XOR U416 ( .A(p_input[63]), .B(n454), .Z(n456) );
  XNOR U417 ( .A(n457), .B(n458), .Z(n454) );
  AND U418 ( .A(n78), .B(n453), .Z(n458) );
  XNOR U419 ( .A(n457), .B(n451), .Z(n453) );
  XOR U420 ( .A(n459), .B(n460), .Z(n451) );
  AND U421 ( .A(n93), .B(n461), .Z(n460) );
  XNOR U422 ( .A(n462), .B(n463), .Z(n457) );
  AND U423 ( .A(n85), .B(n464), .Z(n463) );
  XOR U424 ( .A(p_input[95]), .B(n462), .Z(n464) );
  XNOR U425 ( .A(n465), .B(n466), .Z(n462) );
  AND U426 ( .A(n89), .B(n461), .Z(n466) );
  XNOR U427 ( .A(n465), .B(n459), .Z(n461) );
  XOR U428 ( .A(n467), .B(n468), .Z(n459) );
  AND U429 ( .A(n104), .B(n469), .Z(n468) );
  XNOR U430 ( .A(n470), .B(n471), .Z(n465) );
  AND U431 ( .A(n96), .B(n472), .Z(n471) );
  XOR U432 ( .A(p_input[127]), .B(n470), .Z(n472) );
  XNOR U433 ( .A(n473), .B(n474), .Z(n470) );
  AND U434 ( .A(n100), .B(n469), .Z(n474) );
  XNOR U435 ( .A(n473), .B(n467), .Z(n469) );
  XOR U436 ( .A(n475), .B(n476), .Z(n467) );
  AND U437 ( .A(n115), .B(n477), .Z(n476) );
  XNOR U438 ( .A(n478), .B(n479), .Z(n473) );
  AND U439 ( .A(n107), .B(n480), .Z(n479) );
  XOR U440 ( .A(p_input[159]), .B(n478), .Z(n480) );
  XNOR U441 ( .A(n481), .B(n482), .Z(n478) );
  AND U442 ( .A(n111), .B(n477), .Z(n482) );
  XNOR U443 ( .A(n481), .B(n475), .Z(n477) );
  XOR U444 ( .A(\knn_comb_/min_val_out[0][31] ), .B(n483), .Z(n475) );
  AND U445 ( .A(n125), .B(n484), .Z(n483) );
  XNOR U446 ( .A(n485), .B(n486), .Z(n481) );
  AND U447 ( .A(n118), .B(n487), .Z(n486) );
  XOR U448 ( .A(p_input[191]), .B(n485), .Z(n487) );
  XNOR U449 ( .A(n488), .B(n489), .Z(n485) );
  AND U450 ( .A(n122), .B(n484), .Z(n489) );
  XOR U451 ( .A(n490), .B(n488), .Z(n484) );
  IV U452 ( .A(\knn_comb_/min_val_out[0][31] ), .Z(n490) );
  IV U453 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .Z(n488) );
  XOR U454 ( .A(n11), .B(n491), .Z(o[30]) );
  AND U455 ( .A(n58), .B(n492), .Z(n11) );
  XOR U456 ( .A(n12), .B(n491), .Z(n492) );
  XOR U457 ( .A(n493), .B(n494), .Z(n491) );
  AND U458 ( .A(n70), .B(n495), .Z(n494) );
  XOR U459 ( .A(n496), .B(n497), .Z(n12) );
  AND U460 ( .A(n62), .B(n498), .Z(n497) );
  XOR U461 ( .A(p_input[30]), .B(n496), .Z(n498) );
  XNOR U462 ( .A(n499), .B(n500), .Z(n496) );
  AND U463 ( .A(n66), .B(n495), .Z(n500) );
  XNOR U464 ( .A(n499), .B(n493), .Z(n495) );
  XOR U465 ( .A(n501), .B(n502), .Z(n493) );
  AND U466 ( .A(n82), .B(n503), .Z(n502) );
  XNOR U467 ( .A(n504), .B(n505), .Z(n499) );
  AND U468 ( .A(n74), .B(n506), .Z(n505) );
  XOR U469 ( .A(p_input[62]), .B(n504), .Z(n506) );
  XNOR U470 ( .A(n507), .B(n508), .Z(n504) );
  AND U471 ( .A(n78), .B(n503), .Z(n508) );
  XNOR U472 ( .A(n507), .B(n501), .Z(n503) );
  XOR U473 ( .A(n509), .B(n510), .Z(n501) );
  AND U474 ( .A(n93), .B(n511), .Z(n510) );
  XNOR U475 ( .A(n512), .B(n513), .Z(n507) );
  AND U476 ( .A(n85), .B(n514), .Z(n513) );
  XOR U477 ( .A(p_input[94]), .B(n512), .Z(n514) );
  XNOR U478 ( .A(n515), .B(n516), .Z(n512) );
  AND U479 ( .A(n89), .B(n511), .Z(n516) );
  XNOR U480 ( .A(n515), .B(n509), .Z(n511) );
  XOR U481 ( .A(n517), .B(n518), .Z(n509) );
  AND U482 ( .A(n104), .B(n519), .Z(n518) );
  XNOR U483 ( .A(n520), .B(n521), .Z(n515) );
  AND U484 ( .A(n96), .B(n522), .Z(n521) );
  XOR U485 ( .A(p_input[126]), .B(n520), .Z(n522) );
  XNOR U486 ( .A(n523), .B(n524), .Z(n520) );
  AND U487 ( .A(n100), .B(n519), .Z(n524) );
  XNOR U488 ( .A(n523), .B(n517), .Z(n519) );
  XOR U489 ( .A(n525), .B(n526), .Z(n517) );
  AND U490 ( .A(n115), .B(n527), .Z(n526) );
  XNOR U491 ( .A(n528), .B(n529), .Z(n523) );
  AND U492 ( .A(n107), .B(n530), .Z(n529) );
  XOR U493 ( .A(p_input[158]), .B(n528), .Z(n530) );
  XNOR U494 ( .A(n531), .B(n532), .Z(n528) );
  AND U495 ( .A(n111), .B(n527), .Z(n532) );
  XNOR U496 ( .A(n531), .B(n525), .Z(n527) );
  XOR U497 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n533), .Z(n525) );
  AND U498 ( .A(n125), .B(n534), .Z(n533) );
  XNOR U499 ( .A(n535), .B(n536), .Z(n531) );
  AND U500 ( .A(n118), .B(n537), .Z(n536) );
  XOR U501 ( .A(p_input[190]), .B(n535), .Z(n537) );
  XNOR U502 ( .A(n538), .B(n539), .Z(n535) );
  AND U503 ( .A(n122), .B(n534), .Z(n539) );
  XOR U504 ( .A(n540), .B(n538), .Z(n534) );
  IV U505 ( .A(\knn_comb_/min_val_out[0][30] ), .Z(n540) );
  IV U506 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .Z(n538) );
  XOR U507 ( .A(n435), .B(n541), .Z(o[2]) );
  AND U508 ( .A(n58), .B(n542), .Z(n435) );
  XOR U509 ( .A(n436), .B(n541), .Z(n542) );
  XOR U510 ( .A(n543), .B(n544), .Z(n541) );
  AND U511 ( .A(n70), .B(n545), .Z(n544) );
  XOR U512 ( .A(n546), .B(n547), .Z(n436) );
  AND U513 ( .A(n62), .B(n548), .Z(n547) );
  XOR U514 ( .A(p_input[2]), .B(n546), .Z(n548) );
  XNOR U515 ( .A(n549), .B(n550), .Z(n546) );
  AND U516 ( .A(n66), .B(n545), .Z(n550) );
  XNOR U517 ( .A(n549), .B(n543), .Z(n545) );
  XOR U518 ( .A(n551), .B(n552), .Z(n543) );
  AND U519 ( .A(n82), .B(n553), .Z(n552) );
  XNOR U520 ( .A(n554), .B(n555), .Z(n549) );
  AND U521 ( .A(n74), .B(n556), .Z(n555) );
  XOR U522 ( .A(p_input[34]), .B(n554), .Z(n556) );
  XNOR U523 ( .A(n557), .B(n558), .Z(n554) );
  AND U524 ( .A(n78), .B(n553), .Z(n558) );
  XNOR U525 ( .A(n557), .B(n551), .Z(n553) );
  XOR U526 ( .A(n559), .B(n560), .Z(n551) );
  AND U527 ( .A(n93), .B(n561), .Z(n560) );
  XNOR U528 ( .A(n562), .B(n563), .Z(n557) );
  AND U529 ( .A(n85), .B(n564), .Z(n563) );
  XOR U530 ( .A(p_input[66]), .B(n562), .Z(n564) );
  XNOR U531 ( .A(n565), .B(n566), .Z(n562) );
  AND U532 ( .A(n89), .B(n561), .Z(n566) );
  XNOR U533 ( .A(n565), .B(n559), .Z(n561) );
  XOR U534 ( .A(n567), .B(n568), .Z(n559) );
  AND U535 ( .A(n104), .B(n569), .Z(n568) );
  XNOR U536 ( .A(n570), .B(n571), .Z(n565) );
  AND U537 ( .A(n96), .B(n572), .Z(n571) );
  XOR U538 ( .A(p_input[98]), .B(n570), .Z(n572) );
  XNOR U539 ( .A(n573), .B(n574), .Z(n570) );
  AND U540 ( .A(n100), .B(n569), .Z(n574) );
  XNOR U541 ( .A(n573), .B(n567), .Z(n569) );
  XOR U542 ( .A(n575), .B(n576), .Z(n567) );
  AND U543 ( .A(n115), .B(n577), .Z(n576) );
  XNOR U544 ( .A(n578), .B(n579), .Z(n573) );
  AND U545 ( .A(n107), .B(n580), .Z(n579) );
  XOR U546 ( .A(p_input[130]), .B(n578), .Z(n580) );
  XNOR U547 ( .A(n581), .B(n582), .Z(n578) );
  AND U548 ( .A(n111), .B(n577), .Z(n582) );
  XNOR U549 ( .A(n581), .B(n575), .Z(n577) );
  XOR U550 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n583), .Z(n575) );
  AND U551 ( .A(n125), .B(n584), .Z(n583) );
  XNOR U552 ( .A(n585), .B(n586), .Z(n581) );
  AND U553 ( .A(n118), .B(n587), .Z(n586) );
  XOR U554 ( .A(p_input[162]), .B(n585), .Z(n587) );
  XNOR U555 ( .A(n588), .B(n589), .Z(n585) );
  AND U556 ( .A(n122), .B(n584), .Z(n589) );
  XOR U557 ( .A(\knn_comb_/min_val_out[0][2] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n584) );
  XOR U558 ( .A(n13), .B(n590), .Z(o[29]) );
  AND U559 ( .A(n58), .B(n591), .Z(n13) );
  XOR U560 ( .A(n14), .B(n590), .Z(n591) );
  XOR U561 ( .A(n592), .B(n593), .Z(n590) );
  AND U562 ( .A(n70), .B(n594), .Z(n593) );
  XOR U563 ( .A(n595), .B(n596), .Z(n14) );
  AND U564 ( .A(n62), .B(n597), .Z(n596) );
  XOR U565 ( .A(p_input[29]), .B(n595), .Z(n597) );
  XNOR U566 ( .A(n598), .B(n599), .Z(n595) );
  AND U567 ( .A(n66), .B(n594), .Z(n599) );
  XNOR U568 ( .A(n598), .B(n592), .Z(n594) );
  XOR U569 ( .A(n600), .B(n601), .Z(n592) );
  AND U570 ( .A(n82), .B(n602), .Z(n601) );
  XNOR U571 ( .A(n603), .B(n604), .Z(n598) );
  AND U572 ( .A(n74), .B(n605), .Z(n604) );
  XOR U573 ( .A(p_input[61]), .B(n603), .Z(n605) );
  XNOR U574 ( .A(n606), .B(n607), .Z(n603) );
  AND U575 ( .A(n78), .B(n602), .Z(n607) );
  XNOR U576 ( .A(n606), .B(n600), .Z(n602) );
  XOR U577 ( .A(n608), .B(n609), .Z(n600) );
  AND U578 ( .A(n93), .B(n610), .Z(n609) );
  XNOR U579 ( .A(n611), .B(n612), .Z(n606) );
  AND U580 ( .A(n85), .B(n613), .Z(n612) );
  XOR U581 ( .A(p_input[93]), .B(n611), .Z(n613) );
  XNOR U582 ( .A(n614), .B(n615), .Z(n611) );
  AND U583 ( .A(n89), .B(n610), .Z(n615) );
  XNOR U584 ( .A(n614), .B(n608), .Z(n610) );
  XOR U585 ( .A(n616), .B(n617), .Z(n608) );
  AND U586 ( .A(n104), .B(n618), .Z(n617) );
  XNOR U587 ( .A(n619), .B(n620), .Z(n614) );
  AND U588 ( .A(n96), .B(n621), .Z(n620) );
  XOR U589 ( .A(p_input[125]), .B(n619), .Z(n621) );
  XNOR U590 ( .A(n622), .B(n623), .Z(n619) );
  AND U591 ( .A(n100), .B(n618), .Z(n623) );
  XNOR U592 ( .A(n622), .B(n616), .Z(n618) );
  XOR U593 ( .A(n624), .B(n625), .Z(n616) );
  AND U594 ( .A(n115), .B(n626), .Z(n625) );
  XNOR U595 ( .A(n627), .B(n628), .Z(n622) );
  AND U596 ( .A(n107), .B(n629), .Z(n628) );
  XOR U597 ( .A(p_input[157]), .B(n627), .Z(n629) );
  XNOR U598 ( .A(n630), .B(n631), .Z(n627) );
  AND U599 ( .A(n111), .B(n626), .Z(n631) );
  XNOR U600 ( .A(n630), .B(n624), .Z(n626) );
  XOR U601 ( .A(\knn_comb_/min_val_out[0][29] ), .B(n632), .Z(n624) );
  AND U602 ( .A(n125), .B(n633), .Z(n632) );
  XNOR U603 ( .A(n634), .B(n635), .Z(n630) );
  AND U604 ( .A(n118), .B(n636), .Z(n635) );
  XOR U605 ( .A(p_input[189]), .B(n634), .Z(n636) );
  XNOR U606 ( .A(n637), .B(n638), .Z(n634) );
  AND U607 ( .A(n122), .B(n633), .Z(n638) );
  XOR U608 ( .A(\knn_comb_/min_val_out[0][29] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .Z(n633) );
  XOR U609 ( .A(n15), .B(n639), .Z(o[28]) );
  AND U610 ( .A(n58), .B(n640), .Z(n15) );
  XOR U611 ( .A(n16), .B(n639), .Z(n640) );
  XOR U612 ( .A(n641), .B(n642), .Z(n639) );
  AND U613 ( .A(n70), .B(n643), .Z(n642) );
  XOR U614 ( .A(n644), .B(n645), .Z(n16) );
  AND U615 ( .A(n62), .B(n646), .Z(n645) );
  XOR U616 ( .A(p_input[28]), .B(n644), .Z(n646) );
  XNOR U617 ( .A(n647), .B(n648), .Z(n644) );
  AND U618 ( .A(n66), .B(n643), .Z(n648) );
  XNOR U619 ( .A(n647), .B(n641), .Z(n643) );
  XOR U620 ( .A(n649), .B(n650), .Z(n641) );
  AND U621 ( .A(n82), .B(n651), .Z(n650) );
  XNOR U622 ( .A(n652), .B(n653), .Z(n647) );
  AND U623 ( .A(n74), .B(n654), .Z(n653) );
  XOR U624 ( .A(p_input[60]), .B(n652), .Z(n654) );
  XNOR U625 ( .A(n655), .B(n656), .Z(n652) );
  AND U626 ( .A(n78), .B(n651), .Z(n656) );
  XNOR U627 ( .A(n655), .B(n649), .Z(n651) );
  XOR U628 ( .A(n657), .B(n658), .Z(n649) );
  AND U629 ( .A(n93), .B(n659), .Z(n658) );
  XNOR U630 ( .A(n660), .B(n661), .Z(n655) );
  AND U631 ( .A(n85), .B(n662), .Z(n661) );
  XOR U632 ( .A(p_input[92]), .B(n660), .Z(n662) );
  XNOR U633 ( .A(n663), .B(n664), .Z(n660) );
  AND U634 ( .A(n89), .B(n659), .Z(n664) );
  XNOR U635 ( .A(n663), .B(n657), .Z(n659) );
  XOR U636 ( .A(n665), .B(n666), .Z(n657) );
  AND U637 ( .A(n104), .B(n667), .Z(n666) );
  XNOR U638 ( .A(n668), .B(n669), .Z(n663) );
  AND U639 ( .A(n96), .B(n670), .Z(n669) );
  XOR U640 ( .A(p_input[124]), .B(n668), .Z(n670) );
  XNOR U641 ( .A(n671), .B(n672), .Z(n668) );
  AND U642 ( .A(n100), .B(n667), .Z(n672) );
  XNOR U643 ( .A(n671), .B(n665), .Z(n667) );
  XOR U644 ( .A(n673), .B(n674), .Z(n665) );
  AND U645 ( .A(n115), .B(n675), .Z(n674) );
  XNOR U646 ( .A(n676), .B(n677), .Z(n671) );
  AND U647 ( .A(n107), .B(n678), .Z(n677) );
  XOR U648 ( .A(p_input[156]), .B(n676), .Z(n678) );
  XNOR U649 ( .A(n679), .B(n680), .Z(n676) );
  AND U650 ( .A(n111), .B(n675), .Z(n680) );
  XNOR U651 ( .A(n679), .B(n673), .Z(n675) );
  XOR U652 ( .A(\knn_comb_/min_val_out[0][28] ), .B(n681), .Z(n673) );
  AND U653 ( .A(n125), .B(n682), .Z(n681) );
  XNOR U654 ( .A(n683), .B(n684), .Z(n679) );
  AND U655 ( .A(n118), .B(n685), .Z(n684) );
  XOR U656 ( .A(p_input[188]), .B(n683), .Z(n685) );
  XNOR U657 ( .A(n686), .B(n687), .Z(n683) );
  AND U658 ( .A(n122), .B(n682), .Z(n687) );
  XOR U659 ( .A(\knn_comb_/min_val_out[0][28] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .Z(n682) );
  XOR U660 ( .A(n19), .B(n688), .Z(o[27]) );
  AND U661 ( .A(n58), .B(n689), .Z(n19) );
  XOR U662 ( .A(n20), .B(n688), .Z(n689) );
  XOR U663 ( .A(n690), .B(n691), .Z(n688) );
  AND U664 ( .A(n70), .B(n692), .Z(n691) );
  XOR U665 ( .A(n693), .B(n694), .Z(n20) );
  AND U666 ( .A(n62), .B(n695), .Z(n694) );
  XOR U667 ( .A(p_input[27]), .B(n693), .Z(n695) );
  XNOR U668 ( .A(n696), .B(n697), .Z(n693) );
  AND U669 ( .A(n66), .B(n692), .Z(n697) );
  XNOR U670 ( .A(n696), .B(n690), .Z(n692) );
  XOR U671 ( .A(n698), .B(n699), .Z(n690) );
  AND U672 ( .A(n82), .B(n700), .Z(n699) );
  XNOR U673 ( .A(n701), .B(n702), .Z(n696) );
  AND U674 ( .A(n74), .B(n703), .Z(n702) );
  XOR U675 ( .A(p_input[59]), .B(n701), .Z(n703) );
  XNOR U676 ( .A(n704), .B(n705), .Z(n701) );
  AND U677 ( .A(n78), .B(n700), .Z(n705) );
  XNOR U678 ( .A(n704), .B(n698), .Z(n700) );
  XOR U679 ( .A(n706), .B(n707), .Z(n698) );
  AND U680 ( .A(n93), .B(n708), .Z(n707) );
  XNOR U681 ( .A(n709), .B(n710), .Z(n704) );
  AND U682 ( .A(n85), .B(n711), .Z(n710) );
  XOR U683 ( .A(p_input[91]), .B(n709), .Z(n711) );
  XNOR U684 ( .A(n712), .B(n713), .Z(n709) );
  AND U685 ( .A(n89), .B(n708), .Z(n713) );
  XNOR U686 ( .A(n712), .B(n706), .Z(n708) );
  XOR U687 ( .A(n714), .B(n715), .Z(n706) );
  AND U688 ( .A(n104), .B(n716), .Z(n715) );
  XNOR U689 ( .A(n717), .B(n718), .Z(n712) );
  AND U690 ( .A(n96), .B(n719), .Z(n718) );
  XOR U691 ( .A(p_input[123]), .B(n717), .Z(n719) );
  XNOR U692 ( .A(n720), .B(n721), .Z(n717) );
  AND U693 ( .A(n100), .B(n716), .Z(n721) );
  XNOR U694 ( .A(n720), .B(n714), .Z(n716) );
  XOR U695 ( .A(n722), .B(n723), .Z(n714) );
  AND U696 ( .A(n115), .B(n724), .Z(n723) );
  XNOR U697 ( .A(n725), .B(n726), .Z(n720) );
  AND U698 ( .A(n107), .B(n727), .Z(n726) );
  XOR U699 ( .A(p_input[155]), .B(n725), .Z(n727) );
  XNOR U700 ( .A(n728), .B(n729), .Z(n725) );
  AND U701 ( .A(n111), .B(n724), .Z(n729) );
  XNOR U702 ( .A(n728), .B(n722), .Z(n724) );
  XOR U703 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n730), .Z(n722) );
  AND U704 ( .A(n125), .B(n731), .Z(n730) );
  XNOR U705 ( .A(n732), .B(n733), .Z(n728) );
  AND U706 ( .A(n118), .B(n734), .Z(n733) );
  XOR U707 ( .A(p_input[187]), .B(n732), .Z(n734) );
  XNOR U708 ( .A(n735), .B(n736), .Z(n732) );
  AND U709 ( .A(n122), .B(n731), .Z(n736) );
  XOR U710 ( .A(n737), .B(n735), .Z(n731) );
  IV U711 ( .A(\knn_comb_/min_val_out[0][27] ), .Z(n737) );
  IV U712 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .Z(n735) );
  XOR U713 ( .A(n21), .B(n738), .Z(o[26]) );
  AND U714 ( .A(n58), .B(n739), .Z(n21) );
  XOR U715 ( .A(n22), .B(n738), .Z(n739) );
  XOR U716 ( .A(n740), .B(n741), .Z(n738) );
  AND U717 ( .A(n70), .B(n742), .Z(n741) );
  XOR U718 ( .A(n743), .B(n744), .Z(n22) );
  AND U719 ( .A(n62), .B(n745), .Z(n744) );
  XOR U720 ( .A(p_input[26]), .B(n743), .Z(n745) );
  XNOR U721 ( .A(n746), .B(n747), .Z(n743) );
  AND U722 ( .A(n66), .B(n742), .Z(n747) );
  XNOR U723 ( .A(n746), .B(n740), .Z(n742) );
  XOR U724 ( .A(n748), .B(n749), .Z(n740) );
  AND U725 ( .A(n82), .B(n750), .Z(n749) );
  XNOR U726 ( .A(n751), .B(n752), .Z(n746) );
  AND U727 ( .A(n74), .B(n753), .Z(n752) );
  XOR U728 ( .A(p_input[58]), .B(n751), .Z(n753) );
  XNOR U729 ( .A(n754), .B(n755), .Z(n751) );
  AND U730 ( .A(n78), .B(n750), .Z(n755) );
  XNOR U731 ( .A(n754), .B(n748), .Z(n750) );
  XOR U732 ( .A(n756), .B(n757), .Z(n748) );
  AND U733 ( .A(n93), .B(n758), .Z(n757) );
  XNOR U734 ( .A(n759), .B(n760), .Z(n754) );
  AND U735 ( .A(n85), .B(n761), .Z(n760) );
  XOR U736 ( .A(p_input[90]), .B(n759), .Z(n761) );
  XNOR U737 ( .A(n762), .B(n763), .Z(n759) );
  AND U738 ( .A(n89), .B(n758), .Z(n763) );
  XNOR U739 ( .A(n762), .B(n756), .Z(n758) );
  XOR U740 ( .A(n764), .B(n765), .Z(n756) );
  AND U741 ( .A(n104), .B(n766), .Z(n765) );
  XNOR U742 ( .A(n767), .B(n768), .Z(n762) );
  AND U743 ( .A(n96), .B(n769), .Z(n768) );
  XOR U744 ( .A(p_input[122]), .B(n767), .Z(n769) );
  XNOR U745 ( .A(n770), .B(n771), .Z(n767) );
  AND U746 ( .A(n100), .B(n766), .Z(n771) );
  XNOR U747 ( .A(n770), .B(n764), .Z(n766) );
  XOR U748 ( .A(n772), .B(n773), .Z(n764) );
  AND U749 ( .A(n115), .B(n774), .Z(n773) );
  XNOR U750 ( .A(n775), .B(n776), .Z(n770) );
  AND U751 ( .A(n107), .B(n777), .Z(n776) );
  XOR U752 ( .A(p_input[154]), .B(n775), .Z(n777) );
  XNOR U753 ( .A(n778), .B(n779), .Z(n775) );
  AND U754 ( .A(n111), .B(n774), .Z(n779) );
  XNOR U755 ( .A(n778), .B(n772), .Z(n774) );
  XOR U756 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n780), .Z(n772) );
  AND U757 ( .A(n125), .B(n781), .Z(n780) );
  XNOR U758 ( .A(n782), .B(n783), .Z(n778) );
  AND U759 ( .A(n118), .B(n784), .Z(n783) );
  XOR U760 ( .A(p_input[186]), .B(n782), .Z(n784) );
  XNOR U761 ( .A(n785), .B(n786), .Z(n782) );
  AND U762 ( .A(n122), .B(n781), .Z(n786) );
  XOR U763 ( .A(\knn_comb_/min_val_out[0][26] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .Z(n781) );
  XOR U764 ( .A(n23), .B(n787), .Z(o[25]) );
  AND U765 ( .A(n58), .B(n788), .Z(n23) );
  XOR U766 ( .A(n24), .B(n787), .Z(n788) );
  XOR U767 ( .A(n789), .B(n790), .Z(n787) );
  AND U768 ( .A(n70), .B(n791), .Z(n790) );
  XOR U769 ( .A(n792), .B(n793), .Z(n24) );
  AND U770 ( .A(n62), .B(n794), .Z(n793) );
  XOR U771 ( .A(p_input[25]), .B(n792), .Z(n794) );
  XNOR U772 ( .A(n795), .B(n796), .Z(n792) );
  AND U773 ( .A(n66), .B(n791), .Z(n796) );
  XNOR U774 ( .A(n795), .B(n789), .Z(n791) );
  XOR U775 ( .A(n797), .B(n798), .Z(n789) );
  AND U776 ( .A(n82), .B(n799), .Z(n798) );
  XNOR U777 ( .A(n800), .B(n801), .Z(n795) );
  AND U778 ( .A(n74), .B(n802), .Z(n801) );
  XOR U779 ( .A(p_input[57]), .B(n800), .Z(n802) );
  XNOR U780 ( .A(n803), .B(n804), .Z(n800) );
  AND U781 ( .A(n78), .B(n799), .Z(n804) );
  XNOR U782 ( .A(n803), .B(n797), .Z(n799) );
  XOR U783 ( .A(n805), .B(n806), .Z(n797) );
  AND U784 ( .A(n93), .B(n807), .Z(n806) );
  XNOR U785 ( .A(n808), .B(n809), .Z(n803) );
  AND U786 ( .A(n85), .B(n810), .Z(n809) );
  XOR U787 ( .A(p_input[89]), .B(n808), .Z(n810) );
  XNOR U788 ( .A(n811), .B(n812), .Z(n808) );
  AND U789 ( .A(n89), .B(n807), .Z(n812) );
  XNOR U790 ( .A(n811), .B(n805), .Z(n807) );
  XOR U791 ( .A(n813), .B(n814), .Z(n805) );
  AND U792 ( .A(n104), .B(n815), .Z(n814) );
  XNOR U793 ( .A(n816), .B(n817), .Z(n811) );
  AND U794 ( .A(n96), .B(n818), .Z(n817) );
  XOR U795 ( .A(p_input[121]), .B(n816), .Z(n818) );
  XNOR U796 ( .A(n819), .B(n820), .Z(n816) );
  AND U797 ( .A(n100), .B(n815), .Z(n820) );
  XNOR U798 ( .A(n819), .B(n813), .Z(n815) );
  XOR U799 ( .A(n821), .B(n822), .Z(n813) );
  AND U800 ( .A(n115), .B(n823), .Z(n822) );
  XNOR U801 ( .A(n824), .B(n825), .Z(n819) );
  AND U802 ( .A(n107), .B(n826), .Z(n825) );
  XOR U803 ( .A(p_input[153]), .B(n824), .Z(n826) );
  XNOR U804 ( .A(n827), .B(n828), .Z(n824) );
  AND U805 ( .A(n111), .B(n823), .Z(n828) );
  XNOR U806 ( .A(n827), .B(n821), .Z(n823) );
  XOR U807 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n829), .Z(n821) );
  AND U808 ( .A(n125), .B(n830), .Z(n829) );
  XNOR U809 ( .A(n831), .B(n832), .Z(n827) );
  AND U810 ( .A(n118), .B(n833), .Z(n832) );
  XOR U811 ( .A(p_input[185]), .B(n831), .Z(n833) );
  XNOR U812 ( .A(n834), .B(n835), .Z(n831) );
  AND U813 ( .A(n122), .B(n830), .Z(n835) );
  XOR U814 ( .A(\knn_comb_/min_val_out[0][25] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .Z(n830) );
  XOR U815 ( .A(n25), .B(n836), .Z(o[24]) );
  AND U816 ( .A(n58), .B(n837), .Z(n25) );
  XOR U817 ( .A(n26), .B(n836), .Z(n837) );
  XOR U818 ( .A(n838), .B(n839), .Z(n836) );
  AND U819 ( .A(n70), .B(n840), .Z(n839) );
  XOR U820 ( .A(n841), .B(n842), .Z(n26) );
  AND U821 ( .A(n62), .B(n843), .Z(n842) );
  XOR U822 ( .A(p_input[24]), .B(n841), .Z(n843) );
  XNOR U823 ( .A(n844), .B(n845), .Z(n841) );
  AND U824 ( .A(n66), .B(n840), .Z(n845) );
  XNOR U825 ( .A(n844), .B(n838), .Z(n840) );
  XOR U826 ( .A(n846), .B(n847), .Z(n838) );
  AND U827 ( .A(n82), .B(n848), .Z(n847) );
  XNOR U828 ( .A(n849), .B(n850), .Z(n844) );
  AND U829 ( .A(n74), .B(n851), .Z(n850) );
  XOR U830 ( .A(p_input[56]), .B(n849), .Z(n851) );
  XNOR U831 ( .A(n852), .B(n853), .Z(n849) );
  AND U832 ( .A(n78), .B(n848), .Z(n853) );
  XNOR U833 ( .A(n852), .B(n846), .Z(n848) );
  XOR U834 ( .A(n854), .B(n855), .Z(n846) );
  AND U835 ( .A(n93), .B(n856), .Z(n855) );
  XNOR U836 ( .A(n857), .B(n858), .Z(n852) );
  AND U837 ( .A(n85), .B(n859), .Z(n858) );
  XOR U838 ( .A(p_input[88]), .B(n857), .Z(n859) );
  XNOR U839 ( .A(n860), .B(n861), .Z(n857) );
  AND U840 ( .A(n89), .B(n856), .Z(n861) );
  XNOR U841 ( .A(n860), .B(n854), .Z(n856) );
  XOR U842 ( .A(n862), .B(n863), .Z(n854) );
  AND U843 ( .A(n104), .B(n864), .Z(n863) );
  XNOR U844 ( .A(n865), .B(n866), .Z(n860) );
  AND U845 ( .A(n96), .B(n867), .Z(n866) );
  XOR U846 ( .A(p_input[120]), .B(n865), .Z(n867) );
  XNOR U847 ( .A(n868), .B(n869), .Z(n865) );
  AND U848 ( .A(n100), .B(n864), .Z(n869) );
  XNOR U849 ( .A(n868), .B(n862), .Z(n864) );
  XOR U850 ( .A(n870), .B(n871), .Z(n862) );
  AND U851 ( .A(n115), .B(n872), .Z(n871) );
  XNOR U852 ( .A(n873), .B(n874), .Z(n868) );
  AND U853 ( .A(n107), .B(n875), .Z(n874) );
  XOR U854 ( .A(p_input[152]), .B(n873), .Z(n875) );
  XNOR U855 ( .A(n876), .B(n877), .Z(n873) );
  AND U856 ( .A(n111), .B(n872), .Z(n877) );
  XNOR U857 ( .A(n876), .B(n870), .Z(n872) );
  XOR U858 ( .A(\knn_comb_/min_val_out[0][24] ), .B(n878), .Z(n870) );
  AND U859 ( .A(n125), .B(n879), .Z(n878) );
  XNOR U860 ( .A(n880), .B(n881), .Z(n876) );
  AND U861 ( .A(n118), .B(n882), .Z(n881) );
  XOR U862 ( .A(p_input[184]), .B(n880), .Z(n882) );
  XNOR U863 ( .A(n883), .B(n884), .Z(n880) );
  AND U864 ( .A(n122), .B(n879), .Z(n884) );
  XOR U865 ( .A(\knn_comb_/min_val_out[0][24] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .Z(n879) );
  XOR U866 ( .A(n27), .B(n885), .Z(o[23]) );
  AND U867 ( .A(n58), .B(n886), .Z(n27) );
  XOR U868 ( .A(n28), .B(n885), .Z(n886) );
  XOR U869 ( .A(n887), .B(n888), .Z(n885) );
  AND U870 ( .A(n70), .B(n889), .Z(n888) );
  XOR U871 ( .A(n890), .B(n891), .Z(n28) );
  AND U872 ( .A(n62), .B(n892), .Z(n891) );
  XOR U873 ( .A(p_input[23]), .B(n890), .Z(n892) );
  XNOR U874 ( .A(n893), .B(n894), .Z(n890) );
  AND U875 ( .A(n66), .B(n889), .Z(n894) );
  XNOR U876 ( .A(n893), .B(n887), .Z(n889) );
  XOR U877 ( .A(n895), .B(n896), .Z(n887) );
  AND U878 ( .A(n82), .B(n897), .Z(n896) );
  XNOR U879 ( .A(n898), .B(n899), .Z(n893) );
  AND U880 ( .A(n74), .B(n900), .Z(n899) );
  XOR U881 ( .A(p_input[55]), .B(n898), .Z(n900) );
  XNOR U882 ( .A(n901), .B(n902), .Z(n898) );
  AND U883 ( .A(n78), .B(n897), .Z(n902) );
  XNOR U884 ( .A(n901), .B(n895), .Z(n897) );
  XOR U885 ( .A(n903), .B(n904), .Z(n895) );
  AND U886 ( .A(n93), .B(n905), .Z(n904) );
  XNOR U887 ( .A(n906), .B(n907), .Z(n901) );
  AND U888 ( .A(n85), .B(n908), .Z(n907) );
  XOR U889 ( .A(p_input[87]), .B(n906), .Z(n908) );
  XNOR U890 ( .A(n909), .B(n910), .Z(n906) );
  AND U891 ( .A(n89), .B(n905), .Z(n910) );
  XNOR U892 ( .A(n909), .B(n903), .Z(n905) );
  XOR U893 ( .A(n911), .B(n912), .Z(n903) );
  AND U894 ( .A(n104), .B(n913), .Z(n912) );
  XNOR U895 ( .A(n914), .B(n915), .Z(n909) );
  AND U896 ( .A(n96), .B(n916), .Z(n915) );
  XOR U897 ( .A(p_input[119]), .B(n914), .Z(n916) );
  XNOR U898 ( .A(n917), .B(n918), .Z(n914) );
  AND U899 ( .A(n100), .B(n913), .Z(n918) );
  XNOR U900 ( .A(n917), .B(n911), .Z(n913) );
  XOR U901 ( .A(n919), .B(n920), .Z(n911) );
  AND U902 ( .A(n115), .B(n921), .Z(n920) );
  XNOR U903 ( .A(n922), .B(n923), .Z(n917) );
  AND U904 ( .A(n107), .B(n924), .Z(n923) );
  XOR U905 ( .A(p_input[151]), .B(n922), .Z(n924) );
  XNOR U906 ( .A(n925), .B(n926), .Z(n922) );
  AND U907 ( .A(n111), .B(n921), .Z(n926) );
  XNOR U908 ( .A(n925), .B(n919), .Z(n921) );
  XOR U909 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n927), .Z(n919) );
  AND U910 ( .A(n125), .B(n928), .Z(n927) );
  XNOR U911 ( .A(n929), .B(n930), .Z(n925) );
  AND U912 ( .A(n118), .B(n931), .Z(n930) );
  XOR U913 ( .A(p_input[183]), .B(n929), .Z(n931) );
  XNOR U914 ( .A(n932), .B(n933), .Z(n929) );
  AND U915 ( .A(n122), .B(n928), .Z(n933) );
  XOR U916 ( .A(n934), .B(n932), .Z(n928) );
  IV U917 ( .A(\knn_comb_/min_val_out[0][23] ), .Z(n934) );
  IV U918 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .Z(n932) );
  XOR U919 ( .A(n29), .B(n935), .Z(o[22]) );
  AND U920 ( .A(n58), .B(n936), .Z(n29) );
  XOR U921 ( .A(n30), .B(n935), .Z(n936) );
  XOR U922 ( .A(n937), .B(n938), .Z(n935) );
  AND U923 ( .A(n70), .B(n939), .Z(n938) );
  XOR U924 ( .A(n940), .B(n941), .Z(n30) );
  AND U925 ( .A(n62), .B(n942), .Z(n941) );
  XOR U926 ( .A(p_input[22]), .B(n940), .Z(n942) );
  XNOR U927 ( .A(n943), .B(n944), .Z(n940) );
  AND U928 ( .A(n66), .B(n939), .Z(n944) );
  XNOR U929 ( .A(n943), .B(n937), .Z(n939) );
  XOR U930 ( .A(n945), .B(n946), .Z(n937) );
  AND U931 ( .A(n82), .B(n947), .Z(n946) );
  XNOR U932 ( .A(n948), .B(n949), .Z(n943) );
  AND U933 ( .A(n74), .B(n950), .Z(n949) );
  XOR U934 ( .A(p_input[54]), .B(n948), .Z(n950) );
  XNOR U935 ( .A(n951), .B(n952), .Z(n948) );
  AND U936 ( .A(n78), .B(n947), .Z(n952) );
  XNOR U937 ( .A(n951), .B(n945), .Z(n947) );
  XOR U938 ( .A(n953), .B(n954), .Z(n945) );
  AND U939 ( .A(n93), .B(n955), .Z(n954) );
  XNOR U940 ( .A(n956), .B(n957), .Z(n951) );
  AND U941 ( .A(n85), .B(n958), .Z(n957) );
  XOR U942 ( .A(p_input[86]), .B(n956), .Z(n958) );
  XNOR U943 ( .A(n959), .B(n960), .Z(n956) );
  AND U944 ( .A(n89), .B(n955), .Z(n960) );
  XNOR U945 ( .A(n959), .B(n953), .Z(n955) );
  XOR U946 ( .A(n961), .B(n962), .Z(n953) );
  AND U947 ( .A(n104), .B(n963), .Z(n962) );
  XNOR U948 ( .A(n964), .B(n965), .Z(n959) );
  AND U949 ( .A(n96), .B(n966), .Z(n965) );
  XOR U950 ( .A(p_input[118]), .B(n964), .Z(n966) );
  XNOR U951 ( .A(n967), .B(n968), .Z(n964) );
  AND U952 ( .A(n100), .B(n963), .Z(n968) );
  XNOR U953 ( .A(n967), .B(n961), .Z(n963) );
  XOR U954 ( .A(n969), .B(n970), .Z(n961) );
  AND U955 ( .A(n115), .B(n971), .Z(n970) );
  XNOR U956 ( .A(n972), .B(n973), .Z(n967) );
  AND U957 ( .A(n107), .B(n974), .Z(n973) );
  XOR U958 ( .A(p_input[150]), .B(n972), .Z(n974) );
  XNOR U959 ( .A(n975), .B(n976), .Z(n972) );
  AND U960 ( .A(n111), .B(n971), .Z(n976) );
  XNOR U961 ( .A(n975), .B(n969), .Z(n971) );
  XOR U962 ( .A(\knn_comb_/min_val_out[0][22] ), .B(n977), .Z(n969) );
  AND U963 ( .A(n125), .B(n978), .Z(n977) );
  XNOR U964 ( .A(n979), .B(n980), .Z(n975) );
  AND U965 ( .A(n118), .B(n981), .Z(n980) );
  XOR U966 ( .A(p_input[182]), .B(n979), .Z(n981) );
  XNOR U967 ( .A(n982), .B(n983), .Z(n979) );
  AND U968 ( .A(n122), .B(n978), .Z(n983) );
  XOR U969 ( .A(\knn_comb_/min_val_out[0][22] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .Z(n978) );
  XOR U970 ( .A(n31), .B(n984), .Z(o[21]) );
  AND U971 ( .A(n58), .B(n985), .Z(n31) );
  XOR U972 ( .A(n32), .B(n984), .Z(n985) );
  XOR U973 ( .A(n986), .B(n987), .Z(n984) );
  AND U974 ( .A(n70), .B(n988), .Z(n987) );
  XOR U975 ( .A(n989), .B(n990), .Z(n32) );
  AND U976 ( .A(n62), .B(n991), .Z(n990) );
  XOR U977 ( .A(p_input[21]), .B(n989), .Z(n991) );
  XNOR U978 ( .A(n992), .B(n993), .Z(n989) );
  AND U979 ( .A(n66), .B(n988), .Z(n993) );
  XNOR U980 ( .A(n992), .B(n986), .Z(n988) );
  XOR U981 ( .A(n994), .B(n995), .Z(n986) );
  AND U982 ( .A(n82), .B(n996), .Z(n995) );
  XNOR U983 ( .A(n997), .B(n998), .Z(n992) );
  AND U984 ( .A(n74), .B(n999), .Z(n998) );
  XOR U985 ( .A(p_input[53]), .B(n997), .Z(n999) );
  XNOR U986 ( .A(n1000), .B(n1001), .Z(n997) );
  AND U987 ( .A(n78), .B(n996), .Z(n1001) );
  XNOR U988 ( .A(n1000), .B(n994), .Z(n996) );
  XOR U989 ( .A(n1002), .B(n1003), .Z(n994) );
  AND U990 ( .A(n93), .B(n1004), .Z(n1003) );
  XNOR U991 ( .A(n1005), .B(n1006), .Z(n1000) );
  AND U992 ( .A(n85), .B(n1007), .Z(n1006) );
  XOR U993 ( .A(p_input[85]), .B(n1005), .Z(n1007) );
  XNOR U994 ( .A(n1008), .B(n1009), .Z(n1005) );
  AND U995 ( .A(n89), .B(n1004), .Z(n1009) );
  XNOR U996 ( .A(n1008), .B(n1002), .Z(n1004) );
  XOR U997 ( .A(n1010), .B(n1011), .Z(n1002) );
  AND U998 ( .A(n104), .B(n1012), .Z(n1011) );
  XNOR U999 ( .A(n1013), .B(n1014), .Z(n1008) );
  AND U1000 ( .A(n96), .B(n1015), .Z(n1014) );
  XOR U1001 ( .A(p_input[117]), .B(n1013), .Z(n1015) );
  XNOR U1002 ( .A(n1016), .B(n1017), .Z(n1013) );
  AND U1003 ( .A(n100), .B(n1012), .Z(n1017) );
  XNOR U1004 ( .A(n1016), .B(n1010), .Z(n1012) );
  XOR U1005 ( .A(n1018), .B(n1019), .Z(n1010) );
  AND U1006 ( .A(n115), .B(n1020), .Z(n1019) );
  XNOR U1007 ( .A(n1021), .B(n1022), .Z(n1016) );
  AND U1008 ( .A(n107), .B(n1023), .Z(n1022) );
  XOR U1009 ( .A(p_input[149]), .B(n1021), .Z(n1023) );
  XNOR U1010 ( .A(n1024), .B(n1025), .Z(n1021) );
  AND U1011 ( .A(n111), .B(n1020), .Z(n1025) );
  XNOR U1012 ( .A(n1024), .B(n1018), .Z(n1020) );
  XOR U1013 ( .A(\knn_comb_/min_val_out[0][21] ), .B(n1026), .Z(n1018) );
  AND U1014 ( .A(n125), .B(n1027), .Z(n1026) );
  XNOR U1015 ( .A(n1028), .B(n1029), .Z(n1024) );
  AND U1016 ( .A(n118), .B(n1030), .Z(n1029) );
  XOR U1017 ( .A(p_input[181]), .B(n1028), .Z(n1030) );
  XNOR U1018 ( .A(n1031), .B(n1032), .Z(n1028) );
  AND U1019 ( .A(n122), .B(n1027), .Z(n1032) );
  XOR U1020 ( .A(\knn_comb_/min_val_out[0][21] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .Z(n1027) );
  XOR U1021 ( .A(n33), .B(n1033), .Z(o[20]) );
  AND U1022 ( .A(n58), .B(n1034), .Z(n33) );
  XOR U1023 ( .A(n34), .B(n1033), .Z(n1034) );
  XOR U1024 ( .A(n1035), .B(n1036), .Z(n1033) );
  AND U1025 ( .A(n70), .B(n1037), .Z(n1036) );
  XOR U1026 ( .A(n1038), .B(n1039), .Z(n34) );
  AND U1027 ( .A(n62), .B(n1040), .Z(n1039) );
  XOR U1028 ( .A(p_input[20]), .B(n1038), .Z(n1040) );
  XNOR U1029 ( .A(n1041), .B(n1042), .Z(n1038) );
  AND U1030 ( .A(n66), .B(n1037), .Z(n1042) );
  XNOR U1031 ( .A(n1041), .B(n1035), .Z(n1037) );
  XOR U1032 ( .A(n1043), .B(n1044), .Z(n1035) );
  AND U1033 ( .A(n82), .B(n1045), .Z(n1044) );
  XNOR U1034 ( .A(n1046), .B(n1047), .Z(n1041) );
  AND U1035 ( .A(n74), .B(n1048), .Z(n1047) );
  XOR U1036 ( .A(p_input[52]), .B(n1046), .Z(n1048) );
  XNOR U1037 ( .A(n1049), .B(n1050), .Z(n1046) );
  AND U1038 ( .A(n78), .B(n1045), .Z(n1050) );
  XNOR U1039 ( .A(n1049), .B(n1043), .Z(n1045) );
  XOR U1040 ( .A(n1051), .B(n1052), .Z(n1043) );
  AND U1041 ( .A(n93), .B(n1053), .Z(n1052) );
  XNOR U1042 ( .A(n1054), .B(n1055), .Z(n1049) );
  AND U1043 ( .A(n85), .B(n1056), .Z(n1055) );
  XOR U1044 ( .A(p_input[84]), .B(n1054), .Z(n1056) );
  XNOR U1045 ( .A(n1057), .B(n1058), .Z(n1054) );
  AND U1046 ( .A(n89), .B(n1053), .Z(n1058) );
  XNOR U1047 ( .A(n1057), .B(n1051), .Z(n1053) );
  XOR U1048 ( .A(n1059), .B(n1060), .Z(n1051) );
  AND U1049 ( .A(n104), .B(n1061), .Z(n1060) );
  XNOR U1050 ( .A(n1062), .B(n1063), .Z(n1057) );
  AND U1051 ( .A(n96), .B(n1064), .Z(n1063) );
  XOR U1052 ( .A(p_input[116]), .B(n1062), .Z(n1064) );
  XNOR U1053 ( .A(n1065), .B(n1066), .Z(n1062) );
  AND U1054 ( .A(n100), .B(n1061), .Z(n1066) );
  XNOR U1055 ( .A(n1065), .B(n1059), .Z(n1061) );
  XOR U1056 ( .A(n1067), .B(n1068), .Z(n1059) );
  AND U1057 ( .A(n115), .B(n1069), .Z(n1068) );
  XNOR U1058 ( .A(n1070), .B(n1071), .Z(n1065) );
  AND U1059 ( .A(n107), .B(n1072), .Z(n1071) );
  XOR U1060 ( .A(p_input[148]), .B(n1070), .Z(n1072) );
  XNOR U1061 ( .A(n1073), .B(n1074), .Z(n1070) );
  AND U1062 ( .A(n111), .B(n1069), .Z(n1074) );
  XNOR U1063 ( .A(n1073), .B(n1067), .Z(n1069) );
  XOR U1064 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n1075), .Z(n1067) );
  AND U1065 ( .A(n125), .B(n1076), .Z(n1075) );
  XNOR U1066 ( .A(n1077), .B(n1078), .Z(n1073) );
  AND U1067 ( .A(n118), .B(n1079), .Z(n1078) );
  XOR U1068 ( .A(p_input[180]), .B(n1077), .Z(n1079) );
  XNOR U1069 ( .A(n1080), .B(n1081), .Z(n1077) );
  AND U1070 ( .A(n122), .B(n1076), .Z(n1081) );
  XOR U1071 ( .A(n1082), .B(n1080), .Z(n1076) );
  IV U1072 ( .A(\knn_comb_/min_val_out[0][20] ), .Z(n1082) );
  IV U1073 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .Z(n1080) );
  XOR U1074 ( .A(n437), .B(n1083), .Z(o[1]) );
  AND U1075 ( .A(n58), .B(n1084), .Z(n437) );
  XOR U1076 ( .A(n438), .B(n1083), .Z(n1084) );
  XOR U1077 ( .A(n1085), .B(n1086), .Z(n1083) );
  AND U1078 ( .A(n70), .B(n1087), .Z(n1086) );
  XOR U1079 ( .A(n1088), .B(n1089), .Z(n438) );
  AND U1080 ( .A(n62), .B(n1090), .Z(n1089) );
  XOR U1081 ( .A(p_input[1]), .B(n1088), .Z(n1090) );
  XNOR U1082 ( .A(n1091), .B(n1092), .Z(n1088) );
  AND U1083 ( .A(n66), .B(n1087), .Z(n1092) );
  XNOR U1084 ( .A(n1091), .B(n1085), .Z(n1087) );
  XOR U1085 ( .A(n1093), .B(n1094), .Z(n1085) );
  AND U1086 ( .A(n82), .B(n1095), .Z(n1094) );
  XNOR U1087 ( .A(n1096), .B(n1097), .Z(n1091) );
  AND U1088 ( .A(n74), .B(n1098), .Z(n1097) );
  XOR U1089 ( .A(p_input[33]), .B(n1096), .Z(n1098) );
  XNOR U1090 ( .A(n1099), .B(n1100), .Z(n1096) );
  AND U1091 ( .A(n78), .B(n1095), .Z(n1100) );
  XNOR U1092 ( .A(n1099), .B(n1093), .Z(n1095) );
  XOR U1093 ( .A(n1101), .B(n1102), .Z(n1093) );
  AND U1094 ( .A(n93), .B(n1103), .Z(n1102) );
  XNOR U1095 ( .A(n1104), .B(n1105), .Z(n1099) );
  AND U1096 ( .A(n85), .B(n1106), .Z(n1105) );
  XOR U1097 ( .A(p_input[65]), .B(n1104), .Z(n1106) );
  XNOR U1098 ( .A(n1107), .B(n1108), .Z(n1104) );
  AND U1099 ( .A(n89), .B(n1103), .Z(n1108) );
  XNOR U1100 ( .A(n1107), .B(n1101), .Z(n1103) );
  XOR U1101 ( .A(n1109), .B(n1110), .Z(n1101) );
  AND U1102 ( .A(n104), .B(n1111), .Z(n1110) );
  XNOR U1103 ( .A(n1112), .B(n1113), .Z(n1107) );
  AND U1104 ( .A(n96), .B(n1114), .Z(n1113) );
  XOR U1105 ( .A(p_input[97]), .B(n1112), .Z(n1114) );
  XNOR U1106 ( .A(n1115), .B(n1116), .Z(n1112) );
  AND U1107 ( .A(n100), .B(n1111), .Z(n1116) );
  XNOR U1108 ( .A(n1115), .B(n1109), .Z(n1111) );
  XOR U1109 ( .A(n1117), .B(n1118), .Z(n1109) );
  AND U1110 ( .A(n115), .B(n1119), .Z(n1118) );
  XNOR U1111 ( .A(n1120), .B(n1121), .Z(n1115) );
  AND U1112 ( .A(n107), .B(n1122), .Z(n1121) );
  XOR U1113 ( .A(p_input[129]), .B(n1120), .Z(n1122) );
  XNOR U1114 ( .A(n1123), .B(n1124), .Z(n1120) );
  AND U1115 ( .A(n111), .B(n1119), .Z(n1124) );
  XNOR U1116 ( .A(n1123), .B(n1117), .Z(n1119) );
  XOR U1117 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n1125), .Z(n1117) );
  AND U1118 ( .A(n125), .B(n1126), .Z(n1125) );
  XNOR U1119 ( .A(n1127), .B(n1128), .Z(n1123) );
  AND U1120 ( .A(n118), .B(n1129), .Z(n1128) );
  XOR U1121 ( .A(p_input[161]), .B(n1127), .Z(n1129) );
  XNOR U1122 ( .A(n1130), .B(n1131), .Z(n1127) );
  AND U1123 ( .A(n122), .B(n1126), .Z(n1131) );
  XOR U1124 ( .A(\knn_comb_/min_val_out[0][1] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n1126) );
  XOR U1125 ( .A(n35), .B(n1132), .Z(o[19]) );
  AND U1126 ( .A(n58), .B(n1133), .Z(n35) );
  XOR U1127 ( .A(n36), .B(n1132), .Z(n1133) );
  XOR U1128 ( .A(n1134), .B(n1135), .Z(n1132) );
  AND U1129 ( .A(n70), .B(n1136), .Z(n1135) );
  XOR U1130 ( .A(n1137), .B(n1138), .Z(n36) );
  AND U1131 ( .A(n62), .B(n1139), .Z(n1138) );
  XOR U1132 ( .A(p_input[19]), .B(n1137), .Z(n1139) );
  XNOR U1133 ( .A(n1140), .B(n1141), .Z(n1137) );
  AND U1134 ( .A(n66), .B(n1136), .Z(n1141) );
  XNOR U1135 ( .A(n1140), .B(n1134), .Z(n1136) );
  XOR U1136 ( .A(n1142), .B(n1143), .Z(n1134) );
  AND U1137 ( .A(n82), .B(n1144), .Z(n1143) );
  XNOR U1138 ( .A(n1145), .B(n1146), .Z(n1140) );
  AND U1139 ( .A(n74), .B(n1147), .Z(n1146) );
  XOR U1140 ( .A(p_input[51]), .B(n1145), .Z(n1147) );
  XNOR U1141 ( .A(n1148), .B(n1149), .Z(n1145) );
  AND U1142 ( .A(n78), .B(n1144), .Z(n1149) );
  XNOR U1143 ( .A(n1148), .B(n1142), .Z(n1144) );
  XOR U1144 ( .A(n1150), .B(n1151), .Z(n1142) );
  AND U1145 ( .A(n93), .B(n1152), .Z(n1151) );
  XNOR U1146 ( .A(n1153), .B(n1154), .Z(n1148) );
  AND U1147 ( .A(n85), .B(n1155), .Z(n1154) );
  XOR U1148 ( .A(p_input[83]), .B(n1153), .Z(n1155) );
  XNOR U1149 ( .A(n1156), .B(n1157), .Z(n1153) );
  AND U1150 ( .A(n89), .B(n1152), .Z(n1157) );
  XNOR U1151 ( .A(n1156), .B(n1150), .Z(n1152) );
  XOR U1152 ( .A(n1158), .B(n1159), .Z(n1150) );
  AND U1153 ( .A(n104), .B(n1160), .Z(n1159) );
  XNOR U1154 ( .A(n1161), .B(n1162), .Z(n1156) );
  AND U1155 ( .A(n96), .B(n1163), .Z(n1162) );
  XOR U1156 ( .A(p_input[115]), .B(n1161), .Z(n1163) );
  XNOR U1157 ( .A(n1164), .B(n1165), .Z(n1161) );
  AND U1158 ( .A(n100), .B(n1160), .Z(n1165) );
  XNOR U1159 ( .A(n1164), .B(n1158), .Z(n1160) );
  XOR U1160 ( .A(n1166), .B(n1167), .Z(n1158) );
  AND U1161 ( .A(n115), .B(n1168), .Z(n1167) );
  XNOR U1162 ( .A(n1169), .B(n1170), .Z(n1164) );
  AND U1163 ( .A(n107), .B(n1171), .Z(n1170) );
  XOR U1164 ( .A(p_input[147]), .B(n1169), .Z(n1171) );
  XNOR U1165 ( .A(n1172), .B(n1173), .Z(n1169) );
  AND U1166 ( .A(n111), .B(n1168), .Z(n1173) );
  XNOR U1167 ( .A(n1172), .B(n1166), .Z(n1168) );
  XOR U1168 ( .A(\knn_comb_/min_val_out[0][19] ), .B(n1174), .Z(n1166) );
  AND U1169 ( .A(n125), .B(n1175), .Z(n1174) );
  XNOR U1170 ( .A(n1176), .B(n1177), .Z(n1172) );
  AND U1171 ( .A(n118), .B(n1178), .Z(n1177) );
  XOR U1172 ( .A(p_input[179]), .B(n1176), .Z(n1178) );
  XNOR U1173 ( .A(n1179), .B(n1180), .Z(n1176) );
  AND U1174 ( .A(n122), .B(n1175), .Z(n1180) );
  XOR U1175 ( .A(\knn_comb_/min_val_out[0][19] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .Z(n1175) );
  XOR U1176 ( .A(n37), .B(n1181), .Z(o[18]) );
  AND U1177 ( .A(n58), .B(n1182), .Z(n37) );
  XOR U1178 ( .A(n38), .B(n1181), .Z(n1182) );
  XOR U1179 ( .A(n1183), .B(n1184), .Z(n1181) );
  AND U1180 ( .A(n70), .B(n1185), .Z(n1184) );
  XOR U1181 ( .A(n1186), .B(n1187), .Z(n38) );
  AND U1182 ( .A(n62), .B(n1188), .Z(n1187) );
  XOR U1183 ( .A(p_input[18]), .B(n1186), .Z(n1188) );
  XNOR U1184 ( .A(n1189), .B(n1190), .Z(n1186) );
  AND U1185 ( .A(n66), .B(n1185), .Z(n1190) );
  XNOR U1186 ( .A(n1189), .B(n1183), .Z(n1185) );
  XOR U1187 ( .A(n1191), .B(n1192), .Z(n1183) );
  AND U1188 ( .A(n82), .B(n1193), .Z(n1192) );
  XNOR U1189 ( .A(n1194), .B(n1195), .Z(n1189) );
  AND U1190 ( .A(n74), .B(n1196), .Z(n1195) );
  XOR U1191 ( .A(p_input[50]), .B(n1194), .Z(n1196) );
  XNOR U1192 ( .A(n1197), .B(n1198), .Z(n1194) );
  AND U1193 ( .A(n78), .B(n1193), .Z(n1198) );
  XNOR U1194 ( .A(n1197), .B(n1191), .Z(n1193) );
  XOR U1195 ( .A(n1199), .B(n1200), .Z(n1191) );
  AND U1196 ( .A(n93), .B(n1201), .Z(n1200) );
  XNOR U1197 ( .A(n1202), .B(n1203), .Z(n1197) );
  AND U1198 ( .A(n85), .B(n1204), .Z(n1203) );
  XOR U1199 ( .A(p_input[82]), .B(n1202), .Z(n1204) );
  XNOR U1200 ( .A(n1205), .B(n1206), .Z(n1202) );
  AND U1201 ( .A(n89), .B(n1201), .Z(n1206) );
  XNOR U1202 ( .A(n1205), .B(n1199), .Z(n1201) );
  XOR U1203 ( .A(n1207), .B(n1208), .Z(n1199) );
  AND U1204 ( .A(n104), .B(n1209), .Z(n1208) );
  XNOR U1205 ( .A(n1210), .B(n1211), .Z(n1205) );
  AND U1206 ( .A(n96), .B(n1212), .Z(n1211) );
  XOR U1207 ( .A(p_input[114]), .B(n1210), .Z(n1212) );
  XNOR U1208 ( .A(n1213), .B(n1214), .Z(n1210) );
  AND U1209 ( .A(n100), .B(n1209), .Z(n1214) );
  XNOR U1210 ( .A(n1213), .B(n1207), .Z(n1209) );
  XOR U1211 ( .A(n1215), .B(n1216), .Z(n1207) );
  AND U1212 ( .A(n115), .B(n1217), .Z(n1216) );
  XNOR U1213 ( .A(n1218), .B(n1219), .Z(n1213) );
  AND U1214 ( .A(n107), .B(n1220), .Z(n1219) );
  XOR U1215 ( .A(p_input[146]), .B(n1218), .Z(n1220) );
  XNOR U1216 ( .A(n1221), .B(n1222), .Z(n1218) );
  AND U1217 ( .A(n111), .B(n1217), .Z(n1222) );
  XNOR U1218 ( .A(n1221), .B(n1215), .Z(n1217) );
  XOR U1219 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n1223), .Z(n1215) );
  AND U1220 ( .A(n125), .B(n1224), .Z(n1223) );
  XNOR U1221 ( .A(n1225), .B(n1226), .Z(n1221) );
  AND U1222 ( .A(n118), .B(n1227), .Z(n1226) );
  XOR U1223 ( .A(p_input[178]), .B(n1225), .Z(n1227) );
  XNOR U1224 ( .A(n1228), .B(n1229), .Z(n1225) );
  AND U1225 ( .A(n122), .B(n1224), .Z(n1229) );
  XOR U1226 ( .A(\knn_comb_/min_val_out[0][18] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .Z(n1224) );
  XOR U1227 ( .A(n41), .B(n1230), .Z(o[17]) );
  AND U1228 ( .A(n58), .B(n1231), .Z(n41) );
  XOR U1229 ( .A(n42), .B(n1230), .Z(n1231) );
  XOR U1230 ( .A(n1232), .B(n1233), .Z(n1230) );
  AND U1231 ( .A(n70), .B(n1234), .Z(n1233) );
  XOR U1232 ( .A(n1235), .B(n1236), .Z(n42) );
  AND U1233 ( .A(n62), .B(n1237), .Z(n1236) );
  XOR U1234 ( .A(p_input[17]), .B(n1235), .Z(n1237) );
  XNOR U1235 ( .A(n1238), .B(n1239), .Z(n1235) );
  AND U1236 ( .A(n66), .B(n1234), .Z(n1239) );
  XNOR U1237 ( .A(n1238), .B(n1232), .Z(n1234) );
  XOR U1238 ( .A(n1240), .B(n1241), .Z(n1232) );
  AND U1239 ( .A(n82), .B(n1242), .Z(n1241) );
  XNOR U1240 ( .A(n1243), .B(n1244), .Z(n1238) );
  AND U1241 ( .A(n74), .B(n1245), .Z(n1244) );
  XOR U1242 ( .A(p_input[49]), .B(n1243), .Z(n1245) );
  XNOR U1243 ( .A(n1246), .B(n1247), .Z(n1243) );
  AND U1244 ( .A(n78), .B(n1242), .Z(n1247) );
  XNOR U1245 ( .A(n1246), .B(n1240), .Z(n1242) );
  XOR U1246 ( .A(n1248), .B(n1249), .Z(n1240) );
  AND U1247 ( .A(n93), .B(n1250), .Z(n1249) );
  XNOR U1248 ( .A(n1251), .B(n1252), .Z(n1246) );
  AND U1249 ( .A(n85), .B(n1253), .Z(n1252) );
  XOR U1250 ( .A(p_input[81]), .B(n1251), .Z(n1253) );
  XNOR U1251 ( .A(n1254), .B(n1255), .Z(n1251) );
  AND U1252 ( .A(n89), .B(n1250), .Z(n1255) );
  XNOR U1253 ( .A(n1254), .B(n1248), .Z(n1250) );
  XOR U1254 ( .A(n1256), .B(n1257), .Z(n1248) );
  AND U1255 ( .A(n104), .B(n1258), .Z(n1257) );
  XNOR U1256 ( .A(n1259), .B(n1260), .Z(n1254) );
  AND U1257 ( .A(n96), .B(n1261), .Z(n1260) );
  XOR U1258 ( .A(p_input[113]), .B(n1259), .Z(n1261) );
  XNOR U1259 ( .A(n1262), .B(n1263), .Z(n1259) );
  AND U1260 ( .A(n100), .B(n1258), .Z(n1263) );
  XNOR U1261 ( .A(n1262), .B(n1256), .Z(n1258) );
  XOR U1262 ( .A(n1264), .B(n1265), .Z(n1256) );
  AND U1263 ( .A(n115), .B(n1266), .Z(n1265) );
  XNOR U1264 ( .A(n1267), .B(n1268), .Z(n1262) );
  AND U1265 ( .A(n107), .B(n1269), .Z(n1268) );
  XOR U1266 ( .A(p_input[145]), .B(n1267), .Z(n1269) );
  XNOR U1267 ( .A(n1270), .B(n1271), .Z(n1267) );
  AND U1268 ( .A(n111), .B(n1266), .Z(n1271) );
  XNOR U1269 ( .A(n1270), .B(n1264), .Z(n1266) );
  XOR U1270 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n1272), .Z(n1264) );
  AND U1271 ( .A(n125), .B(n1273), .Z(n1272) );
  XNOR U1272 ( .A(n1274), .B(n1275), .Z(n1270) );
  AND U1273 ( .A(n118), .B(n1276), .Z(n1275) );
  XOR U1274 ( .A(p_input[177]), .B(n1274), .Z(n1276) );
  XNOR U1275 ( .A(n1277), .B(n1278), .Z(n1274) );
  AND U1276 ( .A(n122), .B(n1273), .Z(n1278) );
  XOR U1277 ( .A(\knn_comb_/min_val_out[0][17] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .Z(n1273) );
  XOR U1278 ( .A(n43), .B(n1279), .Z(o[16]) );
  AND U1279 ( .A(n58), .B(n1280), .Z(n43) );
  XOR U1280 ( .A(n44), .B(n1279), .Z(n1280) );
  XOR U1281 ( .A(n1281), .B(n1282), .Z(n1279) );
  AND U1282 ( .A(n70), .B(n1283), .Z(n1282) );
  XOR U1283 ( .A(n1284), .B(n1285), .Z(n44) );
  AND U1284 ( .A(n62), .B(n1286), .Z(n1285) );
  XOR U1285 ( .A(p_input[16]), .B(n1284), .Z(n1286) );
  XNOR U1286 ( .A(n1287), .B(n1288), .Z(n1284) );
  AND U1287 ( .A(n66), .B(n1283), .Z(n1288) );
  XNOR U1288 ( .A(n1287), .B(n1281), .Z(n1283) );
  XOR U1289 ( .A(n1289), .B(n1290), .Z(n1281) );
  AND U1290 ( .A(n82), .B(n1291), .Z(n1290) );
  XNOR U1291 ( .A(n1292), .B(n1293), .Z(n1287) );
  AND U1292 ( .A(n74), .B(n1294), .Z(n1293) );
  XOR U1293 ( .A(p_input[48]), .B(n1292), .Z(n1294) );
  XNOR U1294 ( .A(n1295), .B(n1296), .Z(n1292) );
  AND U1295 ( .A(n78), .B(n1291), .Z(n1296) );
  XNOR U1296 ( .A(n1295), .B(n1289), .Z(n1291) );
  XOR U1297 ( .A(n1297), .B(n1298), .Z(n1289) );
  AND U1298 ( .A(n93), .B(n1299), .Z(n1298) );
  XNOR U1299 ( .A(n1300), .B(n1301), .Z(n1295) );
  AND U1300 ( .A(n85), .B(n1302), .Z(n1301) );
  XOR U1301 ( .A(p_input[80]), .B(n1300), .Z(n1302) );
  XNOR U1302 ( .A(n1303), .B(n1304), .Z(n1300) );
  AND U1303 ( .A(n89), .B(n1299), .Z(n1304) );
  XNOR U1304 ( .A(n1303), .B(n1297), .Z(n1299) );
  XOR U1305 ( .A(n1305), .B(n1306), .Z(n1297) );
  AND U1306 ( .A(n104), .B(n1307), .Z(n1306) );
  XNOR U1307 ( .A(n1308), .B(n1309), .Z(n1303) );
  AND U1308 ( .A(n96), .B(n1310), .Z(n1309) );
  XOR U1309 ( .A(p_input[112]), .B(n1308), .Z(n1310) );
  XNOR U1310 ( .A(n1311), .B(n1312), .Z(n1308) );
  AND U1311 ( .A(n100), .B(n1307), .Z(n1312) );
  XNOR U1312 ( .A(n1311), .B(n1305), .Z(n1307) );
  XOR U1313 ( .A(n1313), .B(n1314), .Z(n1305) );
  AND U1314 ( .A(n115), .B(n1315), .Z(n1314) );
  XNOR U1315 ( .A(n1316), .B(n1317), .Z(n1311) );
  AND U1316 ( .A(n107), .B(n1318), .Z(n1317) );
  XOR U1317 ( .A(p_input[144]), .B(n1316), .Z(n1318) );
  XNOR U1318 ( .A(n1319), .B(n1320), .Z(n1316) );
  AND U1319 ( .A(n111), .B(n1315), .Z(n1320) );
  XNOR U1320 ( .A(n1319), .B(n1313), .Z(n1315) );
  XOR U1321 ( .A(\knn_comb_/min_val_out[0][16] ), .B(n1321), .Z(n1313) );
  AND U1322 ( .A(n125), .B(n1322), .Z(n1321) );
  XNOR U1323 ( .A(n1323), .B(n1324), .Z(n1319) );
  AND U1324 ( .A(n118), .B(n1325), .Z(n1324) );
  XOR U1325 ( .A(p_input[176]), .B(n1323), .Z(n1325) );
  XNOR U1326 ( .A(n1326), .B(n1327), .Z(n1323) );
  AND U1327 ( .A(n122), .B(n1322), .Z(n1327) );
  XOR U1328 ( .A(n1328), .B(n1326), .Z(n1322) );
  IV U1329 ( .A(\knn_comb_/min_val_out[0][16] ), .Z(n1328) );
  IV U1330 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .Z(n1326) );
  XOR U1331 ( .A(n45), .B(n1329), .Z(o[15]) );
  AND U1332 ( .A(n58), .B(n1330), .Z(n45) );
  XOR U1333 ( .A(n46), .B(n1329), .Z(n1330) );
  XOR U1334 ( .A(n1331), .B(n1332), .Z(n1329) );
  AND U1335 ( .A(n70), .B(n1333), .Z(n1332) );
  XOR U1336 ( .A(n1334), .B(n1335), .Z(n46) );
  AND U1337 ( .A(n62), .B(n1336), .Z(n1335) );
  XOR U1338 ( .A(p_input[15]), .B(n1334), .Z(n1336) );
  XNOR U1339 ( .A(n1337), .B(n1338), .Z(n1334) );
  AND U1340 ( .A(n66), .B(n1333), .Z(n1338) );
  XNOR U1341 ( .A(n1337), .B(n1331), .Z(n1333) );
  XOR U1342 ( .A(n1339), .B(n1340), .Z(n1331) );
  AND U1343 ( .A(n82), .B(n1341), .Z(n1340) );
  XNOR U1344 ( .A(n1342), .B(n1343), .Z(n1337) );
  AND U1345 ( .A(n74), .B(n1344), .Z(n1343) );
  XOR U1346 ( .A(p_input[47]), .B(n1342), .Z(n1344) );
  XNOR U1347 ( .A(n1345), .B(n1346), .Z(n1342) );
  AND U1348 ( .A(n78), .B(n1341), .Z(n1346) );
  XNOR U1349 ( .A(n1345), .B(n1339), .Z(n1341) );
  XOR U1350 ( .A(n1347), .B(n1348), .Z(n1339) );
  AND U1351 ( .A(n93), .B(n1349), .Z(n1348) );
  XNOR U1352 ( .A(n1350), .B(n1351), .Z(n1345) );
  AND U1353 ( .A(n85), .B(n1352), .Z(n1351) );
  XOR U1354 ( .A(p_input[79]), .B(n1350), .Z(n1352) );
  XNOR U1355 ( .A(n1353), .B(n1354), .Z(n1350) );
  AND U1356 ( .A(n89), .B(n1349), .Z(n1354) );
  XNOR U1357 ( .A(n1353), .B(n1347), .Z(n1349) );
  XOR U1358 ( .A(n1355), .B(n1356), .Z(n1347) );
  AND U1359 ( .A(n104), .B(n1357), .Z(n1356) );
  XNOR U1360 ( .A(n1358), .B(n1359), .Z(n1353) );
  AND U1361 ( .A(n96), .B(n1360), .Z(n1359) );
  XOR U1362 ( .A(p_input[111]), .B(n1358), .Z(n1360) );
  XNOR U1363 ( .A(n1361), .B(n1362), .Z(n1358) );
  AND U1364 ( .A(n100), .B(n1357), .Z(n1362) );
  XNOR U1365 ( .A(n1361), .B(n1355), .Z(n1357) );
  XOR U1366 ( .A(n1363), .B(n1364), .Z(n1355) );
  AND U1367 ( .A(n115), .B(n1365), .Z(n1364) );
  XNOR U1368 ( .A(n1366), .B(n1367), .Z(n1361) );
  AND U1369 ( .A(n107), .B(n1368), .Z(n1367) );
  XOR U1370 ( .A(p_input[143]), .B(n1366), .Z(n1368) );
  XNOR U1371 ( .A(n1369), .B(n1370), .Z(n1366) );
  AND U1372 ( .A(n111), .B(n1365), .Z(n1370) );
  XNOR U1373 ( .A(n1369), .B(n1363), .Z(n1365) );
  XOR U1374 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n1371), .Z(n1363) );
  AND U1375 ( .A(n125), .B(n1372), .Z(n1371) );
  XNOR U1376 ( .A(n1373), .B(n1374), .Z(n1369) );
  AND U1377 ( .A(n118), .B(n1375), .Z(n1374) );
  XOR U1378 ( .A(p_input[175]), .B(n1373), .Z(n1375) );
  XNOR U1379 ( .A(n1376), .B(n1377), .Z(n1373) );
  AND U1380 ( .A(n122), .B(n1372), .Z(n1377) );
  XOR U1381 ( .A(n1378), .B(n1376), .Z(n1372) );
  IV U1382 ( .A(\knn_comb_/min_val_out[0][15] ), .Z(n1378) );
  IV U1383 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .Z(n1376) );
  XOR U1384 ( .A(n47), .B(n1379), .Z(o[14]) );
  AND U1385 ( .A(n58), .B(n1380), .Z(n47) );
  XOR U1386 ( .A(n48), .B(n1379), .Z(n1380) );
  XOR U1387 ( .A(n1381), .B(n1382), .Z(n1379) );
  AND U1388 ( .A(n70), .B(n1383), .Z(n1382) );
  XOR U1389 ( .A(n1384), .B(n1385), .Z(n48) );
  AND U1390 ( .A(n62), .B(n1386), .Z(n1385) );
  XOR U1391 ( .A(p_input[14]), .B(n1384), .Z(n1386) );
  XNOR U1392 ( .A(n1387), .B(n1388), .Z(n1384) );
  AND U1393 ( .A(n66), .B(n1383), .Z(n1388) );
  XNOR U1394 ( .A(n1387), .B(n1381), .Z(n1383) );
  XOR U1395 ( .A(n1389), .B(n1390), .Z(n1381) );
  AND U1396 ( .A(n82), .B(n1391), .Z(n1390) );
  XNOR U1397 ( .A(n1392), .B(n1393), .Z(n1387) );
  AND U1398 ( .A(n74), .B(n1394), .Z(n1393) );
  XOR U1399 ( .A(p_input[46]), .B(n1392), .Z(n1394) );
  XNOR U1400 ( .A(n1395), .B(n1396), .Z(n1392) );
  AND U1401 ( .A(n78), .B(n1391), .Z(n1396) );
  XNOR U1402 ( .A(n1395), .B(n1389), .Z(n1391) );
  XOR U1403 ( .A(n1397), .B(n1398), .Z(n1389) );
  AND U1404 ( .A(n93), .B(n1399), .Z(n1398) );
  XNOR U1405 ( .A(n1400), .B(n1401), .Z(n1395) );
  AND U1406 ( .A(n85), .B(n1402), .Z(n1401) );
  XOR U1407 ( .A(p_input[78]), .B(n1400), .Z(n1402) );
  XNOR U1408 ( .A(n1403), .B(n1404), .Z(n1400) );
  AND U1409 ( .A(n89), .B(n1399), .Z(n1404) );
  XNOR U1410 ( .A(n1403), .B(n1397), .Z(n1399) );
  XOR U1411 ( .A(n1405), .B(n1406), .Z(n1397) );
  AND U1412 ( .A(n104), .B(n1407), .Z(n1406) );
  XNOR U1413 ( .A(n1408), .B(n1409), .Z(n1403) );
  AND U1414 ( .A(n96), .B(n1410), .Z(n1409) );
  XOR U1415 ( .A(p_input[110]), .B(n1408), .Z(n1410) );
  XNOR U1416 ( .A(n1411), .B(n1412), .Z(n1408) );
  AND U1417 ( .A(n100), .B(n1407), .Z(n1412) );
  XNOR U1418 ( .A(n1411), .B(n1405), .Z(n1407) );
  XOR U1419 ( .A(n1413), .B(n1414), .Z(n1405) );
  AND U1420 ( .A(n115), .B(n1415), .Z(n1414) );
  XNOR U1421 ( .A(n1416), .B(n1417), .Z(n1411) );
  AND U1422 ( .A(n107), .B(n1418), .Z(n1417) );
  XOR U1423 ( .A(p_input[142]), .B(n1416), .Z(n1418) );
  XNOR U1424 ( .A(n1419), .B(n1420), .Z(n1416) );
  AND U1425 ( .A(n111), .B(n1415), .Z(n1420) );
  XNOR U1426 ( .A(n1419), .B(n1413), .Z(n1415) );
  XOR U1427 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n1421), .Z(n1413) );
  AND U1428 ( .A(n125), .B(n1422), .Z(n1421) );
  XNOR U1429 ( .A(n1423), .B(n1424), .Z(n1419) );
  AND U1430 ( .A(n118), .B(n1425), .Z(n1424) );
  XOR U1431 ( .A(p_input[174]), .B(n1423), .Z(n1425) );
  XNOR U1432 ( .A(n1426), .B(n1427), .Z(n1423) );
  AND U1433 ( .A(n122), .B(n1422), .Z(n1427) );
  XOR U1434 ( .A(\knn_comb_/min_val_out[0][14] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n1422) );
  XOR U1435 ( .A(n49), .B(n1428), .Z(o[13]) );
  AND U1436 ( .A(n58), .B(n1429), .Z(n49) );
  XOR U1437 ( .A(n50), .B(n1428), .Z(n1429) );
  XOR U1438 ( .A(n1430), .B(n1431), .Z(n1428) );
  AND U1439 ( .A(n70), .B(n1432), .Z(n1431) );
  XOR U1440 ( .A(n1433), .B(n1434), .Z(n50) );
  AND U1441 ( .A(n62), .B(n1435), .Z(n1434) );
  XOR U1442 ( .A(p_input[13]), .B(n1433), .Z(n1435) );
  XNOR U1443 ( .A(n1436), .B(n1437), .Z(n1433) );
  AND U1444 ( .A(n66), .B(n1432), .Z(n1437) );
  XNOR U1445 ( .A(n1436), .B(n1430), .Z(n1432) );
  XOR U1446 ( .A(n1438), .B(n1439), .Z(n1430) );
  AND U1447 ( .A(n82), .B(n1440), .Z(n1439) );
  XNOR U1448 ( .A(n1441), .B(n1442), .Z(n1436) );
  AND U1449 ( .A(n74), .B(n1443), .Z(n1442) );
  XOR U1450 ( .A(p_input[45]), .B(n1441), .Z(n1443) );
  XNOR U1451 ( .A(n1444), .B(n1445), .Z(n1441) );
  AND U1452 ( .A(n78), .B(n1440), .Z(n1445) );
  XNOR U1453 ( .A(n1444), .B(n1438), .Z(n1440) );
  XOR U1454 ( .A(n1446), .B(n1447), .Z(n1438) );
  AND U1455 ( .A(n93), .B(n1448), .Z(n1447) );
  XNOR U1456 ( .A(n1449), .B(n1450), .Z(n1444) );
  AND U1457 ( .A(n85), .B(n1451), .Z(n1450) );
  XOR U1458 ( .A(p_input[77]), .B(n1449), .Z(n1451) );
  XNOR U1459 ( .A(n1452), .B(n1453), .Z(n1449) );
  AND U1460 ( .A(n89), .B(n1448), .Z(n1453) );
  XNOR U1461 ( .A(n1452), .B(n1446), .Z(n1448) );
  XOR U1462 ( .A(n1454), .B(n1455), .Z(n1446) );
  AND U1463 ( .A(n104), .B(n1456), .Z(n1455) );
  XNOR U1464 ( .A(n1457), .B(n1458), .Z(n1452) );
  AND U1465 ( .A(n96), .B(n1459), .Z(n1458) );
  XOR U1466 ( .A(p_input[109]), .B(n1457), .Z(n1459) );
  XNOR U1467 ( .A(n1460), .B(n1461), .Z(n1457) );
  AND U1468 ( .A(n100), .B(n1456), .Z(n1461) );
  XNOR U1469 ( .A(n1460), .B(n1454), .Z(n1456) );
  XOR U1470 ( .A(n1462), .B(n1463), .Z(n1454) );
  AND U1471 ( .A(n115), .B(n1464), .Z(n1463) );
  XNOR U1472 ( .A(n1465), .B(n1466), .Z(n1460) );
  AND U1473 ( .A(n107), .B(n1467), .Z(n1466) );
  XOR U1474 ( .A(p_input[141]), .B(n1465), .Z(n1467) );
  XNOR U1475 ( .A(n1468), .B(n1469), .Z(n1465) );
  AND U1476 ( .A(n111), .B(n1464), .Z(n1469) );
  XNOR U1477 ( .A(n1468), .B(n1462), .Z(n1464) );
  XOR U1478 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n1470), .Z(n1462) );
  AND U1479 ( .A(n125), .B(n1471), .Z(n1470) );
  XNOR U1480 ( .A(n1472), .B(n1473), .Z(n1468) );
  AND U1481 ( .A(n118), .B(n1474), .Z(n1473) );
  XOR U1482 ( .A(p_input[173]), .B(n1472), .Z(n1474) );
  XNOR U1483 ( .A(n1475), .B(n1476), .Z(n1472) );
  AND U1484 ( .A(n122), .B(n1471), .Z(n1476) );
  XOR U1485 ( .A(\knn_comb_/min_val_out[0][13] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n1471) );
  XOR U1486 ( .A(n51), .B(n1477), .Z(o[12]) );
  AND U1487 ( .A(n58), .B(n1478), .Z(n51) );
  XOR U1488 ( .A(n52), .B(n1477), .Z(n1478) );
  XOR U1489 ( .A(n1479), .B(n1480), .Z(n1477) );
  AND U1490 ( .A(n70), .B(n1481), .Z(n1480) );
  XOR U1491 ( .A(n1482), .B(n1483), .Z(n52) );
  AND U1492 ( .A(n62), .B(n1484), .Z(n1483) );
  XOR U1493 ( .A(p_input[12]), .B(n1482), .Z(n1484) );
  XNOR U1494 ( .A(n1485), .B(n1486), .Z(n1482) );
  AND U1495 ( .A(n66), .B(n1481), .Z(n1486) );
  XNOR U1496 ( .A(n1485), .B(n1479), .Z(n1481) );
  XOR U1497 ( .A(n1487), .B(n1488), .Z(n1479) );
  AND U1498 ( .A(n82), .B(n1489), .Z(n1488) );
  XNOR U1499 ( .A(n1490), .B(n1491), .Z(n1485) );
  AND U1500 ( .A(n74), .B(n1492), .Z(n1491) );
  XOR U1501 ( .A(p_input[44]), .B(n1490), .Z(n1492) );
  XNOR U1502 ( .A(n1493), .B(n1494), .Z(n1490) );
  AND U1503 ( .A(n78), .B(n1489), .Z(n1494) );
  XNOR U1504 ( .A(n1493), .B(n1487), .Z(n1489) );
  XOR U1505 ( .A(n1495), .B(n1496), .Z(n1487) );
  AND U1506 ( .A(n93), .B(n1497), .Z(n1496) );
  XNOR U1507 ( .A(n1498), .B(n1499), .Z(n1493) );
  AND U1508 ( .A(n85), .B(n1500), .Z(n1499) );
  XOR U1509 ( .A(p_input[76]), .B(n1498), .Z(n1500) );
  XNOR U1510 ( .A(n1501), .B(n1502), .Z(n1498) );
  AND U1511 ( .A(n89), .B(n1497), .Z(n1502) );
  XNOR U1512 ( .A(n1501), .B(n1495), .Z(n1497) );
  XOR U1513 ( .A(n1503), .B(n1504), .Z(n1495) );
  AND U1514 ( .A(n104), .B(n1505), .Z(n1504) );
  XNOR U1515 ( .A(n1506), .B(n1507), .Z(n1501) );
  AND U1516 ( .A(n96), .B(n1508), .Z(n1507) );
  XOR U1517 ( .A(p_input[108]), .B(n1506), .Z(n1508) );
  XNOR U1518 ( .A(n1509), .B(n1510), .Z(n1506) );
  AND U1519 ( .A(n100), .B(n1505), .Z(n1510) );
  XNOR U1520 ( .A(n1509), .B(n1503), .Z(n1505) );
  XOR U1521 ( .A(n1511), .B(n1512), .Z(n1503) );
  AND U1522 ( .A(n115), .B(n1513), .Z(n1512) );
  XNOR U1523 ( .A(n1514), .B(n1515), .Z(n1509) );
  AND U1524 ( .A(n107), .B(n1516), .Z(n1515) );
  XOR U1525 ( .A(p_input[140]), .B(n1514), .Z(n1516) );
  XNOR U1526 ( .A(n1517), .B(n1518), .Z(n1514) );
  AND U1527 ( .A(n111), .B(n1513), .Z(n1518) );
  XNOR U1528 ( .A(n1517), .B(n1511), .Z(n1513) );
  XOR U1529 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n1519), .Z(n1511) );
  AND U1530 ( .A(n125), .B(n1520), .Z(n1519) );
  XNOR U1531 ( .A(n1521), .B(n1522), .Z(n1517) );
  AND U1532 ( .A(n118), .B(n1523), .Z(n1522) );
  XOR U1533 ( .A(p_input[172]), .B(n1521), .Z(n1523) );
  XNOR U1534 ( .A(n1524), .B(n1525), .Z(n1521) );
  AND U1535 ( .A(n122), .B(n1520), .Z(n1525) );
  XOR U1536 ( .A(n1526), .B(n1524), .Z(n1520) );
  IV U1537 ( .A(\knn_comb_/min_val_out[0][12] ), .Z(n1526) );
  IV U1538 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n1524) );
  XOR U1539 ( .A(n53), .B(n1527), .Z(o[11]) );
  AND U1540 ( .A(n58), .B(n1528), .Z(n53) );
  XOR U1541 ( .A(n54), .B(n1527), .Z(n1528) );
  XOR U1542 ( .A(n1529), .B(n1530), .Z(n1527) );
  AND U1543 ( .A(n70), .B(n1531), .Z(n1530) );
  XOR U1544 ( .A(n1532), .B(n1533), .Z(n54) );
  AND U1545 ( .A(n62), .B(n1534), .Z(n1533) );
  XOR U1546 ( .A(p_input[11]), .B(n1532), .Z(n1534) );
  XNOR U1547 ( .A(n1535), .B(n1536), .Z(n1532) );
  AND U1548 ( .A(n66), .B(n1531), .Z(n1536) );
  XNOR U1549 ( .A(n1535), .B(n1529), .Z(n1531) );
  XOR U1550 ( .A(n1537), .B(n1538), .Z(n1529) );
  AND U1551 ( .A(n82), .B(n1539), .Z(n1538) );
  XNOR U1552 ( .A(n1540), .B(n1541), .Z(n1535) );
  AND U1553 ( .A(n74), .B(n1542), .Z(n1541) );
  XOR U1554 ( .A(p_input[43]), .B(n1540), .Z(n1542) );
  XNOR U1555 ( .A(n1543), .B(n1544), .Z(n1540) );
  AND U1556 ( .A(n78), .B(n1539), .Z(n1544) );
  XNOR U1557 ( .A(n1543), .B(n1537), .Z(n1539) );
  XOR U1558 ( .A(n1545), .B(n1546), .Z(n1537) );
  AND U1559 ( .A(n93), .B(n1547), .Z(n1546) );
  XNOR U1560 ( .A(n1548), .B(n1549), .Z(n1543) );
  AND U1561 ( .A(n85), .B(n1550), .Z(n1549) );
  XOR U1562 ( .A(p_input[75]), .B(n1548), .Z(n1550) );
  XNOR U1563 ( .A(n1551), .B(n1552), .Z(n1548) );
  AND U1564 ( .A(n89), .B(n1547), .Z(n1552) );
  XNOR U1565 ( .A(n1551), .B(n1545), .Z(n1547) );
  XOR U1566 ( .A(n1553), .B(n1554), .Z(n1545) );
  AND U1567 ( .A(n104), .B(n1555), .Z(n1554) );
  XNOR U1568 ( .A(n1556), .B(n1557), .Z(n1551) );
  AND U1569 ( .A(n96), .B(n1558), .Z(n1557) );
  XOR U1570 ( .A(p_input[107]), .B(n1556), .Z(n1558) );
  XNOR U1571 ( .A(n1559), .B(n1560), .Z(n1556) );
  AND U1572 ( .A(n100), .B(n1555), .Z(n1560) );
  XNOR U1573 ( .A(n1559), .B(n1553), .Z(n1555) );
  XOR U1574 ( .A(n1561), .B(n1562), .Z(n1553) );
  AND U1575 ( .A(n115), .B(n1563), .Z(n1562) );
  XNOR U1576 ( .A(n1564), .B(n1565), .Z(n1559) );
  AND U1577 ( .A(n107), .B(n1566), .Z(n1565) );
  XOR U1578 ( .A(p_input[139]), .B(n1564), .Z(n1566) );
  XNOR U1579 ( .A(n1567), .B(n1568), .Z(n1564) );
  AND U1580 ( .A(n111), .B(n1563), .Z(n1568) );
  XNOR U1581 ( .A(n1567), .B(n1561), .Z(n1563) );
  XOR U1582 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n1569), .Z(n1561) );
  AND U1583 ( .A(n125), .B(n1570), .Z(n1569) );
  XNOR U1584 ( .A(n1571), .B(n1572), .Z(n1567) );
  AND U1585 ( .A(n118), .B(n1573), .Z(n1572) );
  XOR U1586 ( .A(p_input[171]), .B(n1571), .Z(n1573) );
  XNOR U1587 ( .A(n1574), .B(n1575), .Z(n1571) );
  AND U1588 ( .A(n122), .B(n1570), .Z(n1575) );
  XOR U1589 ( .A(\knn_comb_/min_val_out[0][11] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n1570) );
  XOR U1590 ( .A(n55), .B(n1576), .Z(o[10]) );
  AND U1591 ( .A(n58), .B(n1577), .Z(n55) );
  XOR U1592 ( .A(n56), .B(n1576), .Z(n1577) );
  XOR U1593 ( .A(n1578), .B(n1579), .Z(n1576) );
  AND U1594 ( .A(n70), .B(n1580), .Z(n1579) );
  XOR U1595 ( .A(n1581), .B(n1582), .Z(n56) );
  AND U1596 ( .A(n62), .B(n1583), .Z(n1582) );
  XOR U1597 ( .A(p_input[10]), .B(n1581), .Z(n1583) );
  XNOR U1598 ( .A(n1584), .B(n1585), .Z(n1581) );
  AND U1599 ( .A(n66), .B(n1580), .Z(n1585) );
  XNOR U1600 ( .A(n1584), .B(n1578), .Z(n1580) );
  XOR U1601 ( .A(n1586), .B(n1587), .Z(n1578) );
  AND U1602 ( .A(n82), .B(n1588), .Z(n1587) );
  XNOR U1603 ( .A(n1589), .B(n1590), .Z(n1584) );
  AND U1604 ( .A(n74), .B(n1591), .Z(n1590) );
  XOR U1605 ( .A(p_input[42]), .B(n1589), .Z(n1591) );
  XNOR U1606 ( .A(n1592), .B(n1593), .Z(n1589) );
  AND U1607 ( .A(n78), .B(n1588), .Z(n1593) );
  XNOR U1608 ( .A(n1592), .B(n1586), .Z(n1588) );
  XOR U1609 ( .A(n1594), .B(n1595), .Z(n1586) );
  AND U1610 ( .A(n93), .B(n1596), .Z(n1595) );
  XNOR U1611 ( .A(n1597), .B(n1598), .Z(n1592) );
  AND U1612 ( .A(n85), .B(n1599), .Z(n1598) );
  XOR U1613 ( .A(p_input[74]), .B(n1597), .Z(n1599) );
  XNOR U1614 ( .A(n1600), .B(n1601), .Z(n1597) );
  AND U1615 ( .A(n89), .B(n1596), .Z(n1601) );
  XNOR U1616 ( .A(n1600), .B(n1594), .Z(n1596) );
  XOR U1617 ( .A(n1602), .B(n1603), .Z(n1594) );
  AND U1618 ( .A(n104), .B(n1604), .Z(n1603) );
  XNOR U1619 ( .A(n1605), .B(n1606), .Z(n1600) );
  AND U1620 ( .A(n96), .B(n1607), .Z(n1606) );
  XOR U1621 ( .A(p_input[106]), .B(n1605), .Z(n1607) );
  XNOR U1622 ( .A(n1608), .B(n1609), .Z(n1605) );
  AND U1623 ( .A(n100), .B(n1604), .Z(n1609) );
  XNOR U1624 ( .A(n1608), .B(n1602), .Z(n1604) );
  XOR U1625 ( .A(n1610), .B(n1611), .Z(n1602) );
  AND U1626 ( .A(n115), .B(n1612), .Z(n1611) );
  XNOR U1627 ( .A(n1613), .B(n1614), .Z(n1608) );
  AND U1628 ( .A(n107), .B(n1615), .Z(n1614) );
  XOR U1629 ( .A(p_input[138]), .B(n1613), .Z(n1615) );
  XNOR U1630 ( .A(n1616), .B(n1617), .Z(n1613) );
  AND U1631 ( .A(n111), .B(n1612), .Z(n1617) );
  XNOR U1632 ( .A(n1616), .B(n1610), .Z(n1612) );
  XOR U1633 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n1618), .Z(n1610) );
  AND U1634 ( .A(n125), .B(n1619), .Z(n1618) );
  XNOR U1635 ( .A(n1620), .B(n1621), .Z(n1616) );
  AND U1636 ( .A(n118), .B(n1622), .Z(n1621) );
  XOR U1637 ( .A(p_input[170]), .B(n1620), .Z(n1622) );
  XNOR U1638 ( .A(n1623), .B(n1624), .Z(n1620) );
  AND U1639 ( .A(n122), .B(n1619), .Z(n1624) );
  XOR U1640 ( .A(\knn_comb_/min_val_out[0][10] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n1619) );
  XOR U1641 ( .A(n439), .B(n1625), .Z(o[0]) );
  AND U1642 ( .A(n58), .B(n1626), .Z(n439) );
  XOR U1643 ( .A(n440), .B(n1625), .Z(n1626) );
  XOR U1644 ( .A(n1627), .B(n1628), .Z(n1625) );
  AND U1645 ( .A(n70), .B(n1629), .Z(n1628) );
  XOR U1646 ( .A(n1630), .B(n1631), .Z(n440) );
  AND U1647 ( .A(n62), .B(n1632), .Z(n1631) );
  XOR U1648 ( .A(p_input[0]), .B(n1630), .Z(n1632) );
  XNOR U1649 ( .A(n1633), .B(n1634), .Z(n1630) );
  AND U1650 ( .A(n66), .B(n1629), .Z(n1634) );
  XNOR U1651 ( .A(n1633), .B(n1627), .Z(n1629) );
  XOR U1652 ( .A(n1635), .B(n1636), .Z(n1627) );
  AND U1653 ( .A(n82), .B(n1637), .Z(n1636) );
  XNOR U1654 ( .A(n1638), .B(n1639), .Z(n1633) );
  AND U1655 ( .A(n74), .B(n1640), .Z(n1639) );
  XOR U1656 ( .A(p_input[32]), .B(n1638), .Z(n1640) );
  XNOR U1657 ( .A(n1641), .B(n1642), .Z(n1638) );
  AND U1658 ( .A(n78), .B(n1637), .Z(n1642) );
  XNOR U1659 ( .A(n1641), .B(n1635), .Z(n1637) );
  XOR U1660 ( .A(n1643), .B(n1644), .Z(n1635) );
  AND U1661 ( .A(n93), .B(n1645), .Z(n1644) );
  XNOR U1662 ( .A(n1646), .B(n1647), .Z(n1641) );
  AND U1663 ( .A(n85), .B(n1648), .Z(n1647) );
  XOR U1664 ( .A(p_input[64]), .B(n1646), .Z(n1648) );
  XNOR U1665 ( .A(n1649), .B(n1650), .Z(n1646) );
  AND U1666 ( .A(n89), .B(n1645), .Z(n1650) );
  XNOR U1667 ( .A(n1649), .B(n1643), .Z(n1645) );
  XOR U1668 ( .A(n1651), .B(n1652), .Z(n1643) );
  AND U1669 ( .A(n104), .B(n1653), .Z(n1652) );
  XNOR U1670 ( .A(n1654), .B(n1655), .Z(n1649) );
  AND U1671 ( .A(n96), .B(n1656), .Z(n1655) );
  XOR U1672 ( .A(p_input[96]), .B(n1654), .Z(n1656) );
  XNOR U1673 ( .A(n1657), .B(n1658), .Z(n1654) );
  AND U1674 ( .A(n100), .B(n1653), .Z(n1658) );
  XNOR U1675 ( .A(n1657), .B(n1651), .Z(n1653) );
  XOR U1676 ( .A(n1659), .B(n1660), .Z(n1651) );
  AND U1677 ( .A(n115), .B(n1661), .Z(n1660) );
  XNOR U1678 ( .A(n1662), .B(n1663), .Z(n1657) );
  AND U1679 ( .A(n107), .B(n1664), .Z(n1663) );
  XOR U1680 ( .A(p_input[128]), .B(n1662), .Z(n1664) );
  XNOR U1681 ( .A(n1665), .B(n1666), .Z(n1662) );
  AND U1682 ( .A(n111), .B(n1661), .Z(n1666) );
  XNOR U1683 ( .A(n1665), .B(n1659), .Z(n1661) );
  XOR U1684 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n1667), .Z(n1659) );
  AND U1685 ( .A(n125), .B(n1668), .Z(n1667) );
  XNOR U1686 ( .A(n1669), .B(n1670), .Z(n1665) );
  AND U1687 ( .A(n118), .B(n1671), .Z(n1670) );
  XOR U1688 ( .A(p_input[160]), .B(n1669), .Z(n1671) );
  XNOR U1689 ( .A(n1672), .B(n1673), .Z(n1669) );
  AND U1690 ( .A(n122), .B(n1668), .Z(n1673) );
  XOR U1691 ( .A(\knn_comb_/min_val_out[0][0] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n1668) );
  IV U1692 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n1672) );
  XNOR U1693 ( .A(n1674), .B(n1675), .Z(n58) );
  AND U1694 ( .A(n1676), .B(n1677), .Z(n1675) );
  XNOR U1695 ( .A(n1674), .B(n1678), .Z(n1677) );
  XOR U1696 ( .A(n1679), .B(n1680), .Z(n1678) );
  AND U1697 ( .A(n62), .B(n1681), .Z(n1680) );
  XNOR U1698 ( .A(n1679), .B(n1682), .Z(n1681) );
  XNOR U1699 ( .A(n1674), .B(n1683), .Z(n1676) );
  XOR U1700 ( .A(n1684), .B(n1685), .Z(n1683) );
  AND U1701 ( .A(n70), .B(n1686), .Z(n1685) );
  XOR U1702 ( .A(n1687), .B(n1688), .Z(n1674) );
  AND U1703 ( .A(n1689), .B(n1690), .Z(n1688) );
  XOR U1704 ( .A(n1691), .B(n1687), .Z(n1690) );
  XOR U1705 ( .A(n1692), .B(n1693), .Z(n1691) );
  AND U1706 ( .A(n62), .B(n1694), .Z(n1693) );
  XOR U1707 ( .A(n1695), .B(n1692), .Z(n1694) );
  XNOR U1708 ( .A(n1687), .B(n1696), .Z(n1689) );
  XOR U1709 ( .A(n1697), .B(n1698), .Z(n1696) );
  AND U1710 ( .A(n70), .B(n1699), .Z(n1698) );
  XOR U1711 ( .A(n1700), .B(n1701), .Z(n1687) );
  AND U1712 ( .A(n1702), .B(n1703), .Z(n1701) );
  XOR U1713 ( .A(n1704), .B(n1700), .Z(n1703) );
  XOR U1714 ( .A(n1705), .B(n1706), .Z(n1704) );
  AND U1715 ( .A(n62), .B(n1707), .Z(n1706) );
  XNOR U1716 ( .A(n1708), .B(n1705), .Z(n1707) );
  XNOR U1717 ( .A(n1700), .B(n1709), .Z(n1702) );
  XOR U1718 ( .A(n1710), .B(n1711), .Z(n1709) );
  AND U1719 ( .A(n70), .B(n1712), .Z(n1711) );
  XOR U1720 ( .A(n1713), .B(n1714), .Z(n1700) );
  AND U1721 ( .A(n1715), .B(n1716), .Z(n1714) );
  XOR U1722 ( .A(n1717), .B(n1713), .Z(n1716) );
  XOR U1723 ( .A(n1718), .B(n1719), .Z(n1717) );
  AND U1724 ( .A(n62), .B(n1720), .Z(n1719) );
  XOR U1725 ( .A(n1721), .B(n1718), .Z(n1720) );
  XNOR U1726 ( .A(n1713), .B(n1722), .Z(n1715) );
  XOR U1727 ( .A(n1723), .B(n1724), .Z(n1722) );
  AND U1728 ( .A(n70), .B(n1725), .Z(n1724) );
  XOR U1729 ( .A(n1726), .B(n1727), .Z(n1713) );
  AND U1730 ( .A(n1728), .B(n1729), .Z(n1727) );
  XOR U1731 ( .A(n1726), .B(n1730), .Z(n1729) );
  XOR U1732 ( .A(n1731), .B(n1732), .Z(n1730) );
  AND U1733 ( .A(n62), .B(n1733), .Z(n1732) );
  XNOR U1734 ( .A(n1734), .B(n1731), .Z(n1733) );
  XNOR U1735 ( .A(n1735), .B(n1726), .Z(n1728) );
  XNOR U1736 ( .A(n1736), .B(n1737), .Z(n1735) );
  AND U1737 ( .A(n70), .B(n1738), .Z(n1737) );
  AND U1738 ( .A(n1739), .B(n1740), .Z(n1726) );
  XNOR U1739 ( .A(n1741), .B(n1742), .Z(n1740) );
  AND U1740 ( .A(n62), .B(n1743), .Z(n1742) );
  XNOR U1741 ( .A(n1744), .B(n1741), .Z(n1743) );
  XNOR U1742 ( .A(n1745), .B(n1746), .Z(n62) );
  AND U1743 ( .A(n1747), .B(n1748), .Z(n1746) );
  XOR U1744 ( .A(n1682), .B(n1745), .Z(n1748) );
  AND U1745 ( .A(n1749), .B(n1750), .Z(n1682) );
  XOR U1746 ( .A(n1745), .B(n1679), .Z(n1747) );
  XNOR U1747 ( .A(n1751), .B(n1752), .Z(n1679) );
  AND U1748 ( .A(n66), .B(n1686), .Z(n1752) );
  XOR U1749 ( .A(n1684), .B(n1751), .Z(n1686) );
  XOR U1750 ( .A(n1753), .B(n1754), .Z(n1745) );
  AND U1751 ( .A(n1755), .B(n1756), .Z(n1754) );
  XNOR U1752 ( .A(n1753), .B(n1749), .Z(n1756) );
  IV U1753 ( .A(n1695), .Z(n1749) );
  XOR U1754 ( .A(n1757), .B(n1758), .Z(n1695) );
  XOR U1755 ( .A(n1759), .B(n1750), .Z(n1758) );
  AND U1756 ( .A(n1708), .B(n1760), .Z(n1750) );
  AND U1757 ( .A(n1761), .B(n1762), .Z(n1759) );
  XOR U1758 ( .A(n1763), .B(n1757), .Z(n1761) );
  XNOR U1759 ( .A(n1692), .B(n1753), .Z(n1755) );
  XNOR U1760 ( .A(n1764), .B(n1765), .Z(n1692) );
  AND U1761 ( .A(n66), .B(n1699), .Z(n1765) );
  XOR U1762 ( .A(n1764), .B(n1766), .Z(n1699) );
  XOR U1763 ( .A(n1767), .B(n1768), .Z(n1753) );
  AND U1764 ( .A(n1769), .B(n1770), .Z(n1768) );
  XNOR U1765 ( .A(n1767), .B(n1708), .Z(n1770) );
  XOR U1766 ( .A(n1771), .B(n1762), .Z(n1708) );
  XNOR U1767 ( .A(n1772), .B(n1757), .Z(n1762) );
  XOR U1768 ( .A(n1773), .B(n1774), .Z(n1757) );
  AND U1769 ( .A(n1775), .B(n1776), .Z(n1774) );
  XOR U1770 ( .A(n1777), .B(n1773), .Z(n1775) );
  XNOR U1771 ( .A(n1778), .B(n1779), .Z(n1772) );
  AND U1772 ( .A(n1780), .B(n1781), .Z(n1779) );
  XOR U1773 ( .A(n1778), .B(n1782), .Z(n1780) );
  XNOR U1774 ( .A(n1763), .B(n1760), .Z(n1771) );
  AND U1775 ( .A(n1783), .B(n1784), .Z(n1760) );
  XOR U1776 ( .A(n1785), .B(n1786), .Z(n1763) );
  AND U1777 ( .A(n1787), .B(n1788), .Z(n1786) );
  XOR U1778 ( .A(n1785), .B(n1789), .Z(n1787) );
  XNOR U1779 ( .A(n1705), .B(n1767), .Z(n1769) );
  XNOR U1780 ( .A(n1790), .B(n1791), .Z(n1705) );
  AND U1781 ( .A(n66), .B(n1712), .Z(n1791) );
  XOR U1782 ( .A(n1790), .B(n1792), .Z(n1712) );
  XOR U1783 ( .A(n1793), .B(n1794), .Z(n1767) );
  AND U1784 ( .A(n1795), .B(n1796), .Z(n1794) );
  XNOR U1785 ( .A(n1793), .B(n1783), .Z(n1796) );
  IV U1786 ( .A(n1721), .Z(n1783) );
  XNOR U1787 ( .A(n1797), .B(n1776), .Z(n1721) );
  XNOR U1788 ( .A(n1798), .B(n1782), .Z(n1776) );
  XOR U1789 ( .A(n1799), .B(n1800), .Z(n1782) );
  AND U1790 ( .A(n1801), .B(n1802), .Z(n1800) );
  XOR U1791 ( .A(n1799), .B(n1803), .Z(n1801) );
  XNOR U1792 ( .A(n1781), .B(n1773), .Z(n1798) );
  XOR U1793 ( .A(n1804), .B(n1805), .Z(n1773) );
  AND U1794 ( .A(n1806), .B(n1807), .Z(n1805) );
  XNOR U1795 ( .A(n1808), .B(n1804), .Z(n1806) );
  XNOR U1796 ( .A(n1809), .B(n1778), .Z(n1781) );
  XOR U1797 ( .A(n1810), .B(n1811), .Z(n1778) );
  AND U1798 ( .A(n1812), .B(n1813), .Z(n1811) );
  XOR U1799 ( .A(n1810), .B(n1814), .Z(n1812) );
  XNOR U1800 ( .A(n1815), .B(n1816), .Z(n1809) );
  AND U1801 ( .A(n1817), .B(n1818), .Z(n1816) );
  XNOR U1802 ( .A(n1815), .B(n1819), .Z(n1817) );
  XNOR U1803 ( .A(n1777), .B(n1784), .Z(n1797) );
  AND U1804 ( .A(n1734), .B(n1820), .Z(n1784) );
  XOR U1805 ( .A(n1789), .B(n1788), .Z(n1777) );
  XNOR U1806 ( .A(n1821), .B(n1785), .Z(n1788) );
  XOR U1807 ( .A(n1822), .B(n1823), .Z(n1785) );
  AND U1808 ( .A(n1824), .B(n1825), .Z(n1823) );
  XOR U1809 ( .A(n1822), .B(n1826), .Z(n1824) );
  XNOR U1810 ( .A(n1827), .B(n1828), .Z(n1821) );
  AND U1811 ( .A(n1829), .B(n1830), .Z(n1828) );
  XOR U1812 ( .A(n1827), .B(n1831), .Z(n1829) );
  XOR U1813 ( .A(n1832), .B(n1833), .Z(n1789) );
  AND U1814 ( .A(n1834), .B(n1835), .Z(n1833) );
  XOR U1815 ( .A(n1832), .B(n1836), .Z(n1834) );
  XNOR U1816 ( .A(n1718), .B(n1793), .Z(n1795) );
  XNOR U1817 ( .A(n1837), .B(n1838), .Z(n1718) );
  AND U1818 ( .A(n66), .B(n1725), .Z(n1838) );
  XOR U1819 ( .A(n1837), .B(n1839), .Z(n1725) );
  XOR U1820 ( .A(n1840), .B(n1841), .Z(n1793) );
  AND U1821 ( .A(n1842), .B(n1843), .Z(n1841) );
  XNOR U1822 ( .A(n1840), .B(n1734), .Z(n1843) );
  XOR U1823 ( .A(n1844), .B(n1807), .Z(n1734) );
  XNOR U1824 ( .A(n1845), .B(n1814), .Z(n1807) );
  XOR U1825 ( .A(n1803), .B(n1802), .Z(n1814) );
  XNOR U1826 ( .A(n1846), .B(n1799), .Z(n1802) );
  XOR U1827 ( .A(n1847), .B(n1848), .Z(n1799) );
  AND U1828 ( .A(n1849), .B(n1850), .Z(n1848) );
  XNOR U1829 ( .A(n1851), .B(n1852), .Z(n1849) );
  IV U1830 ( .A(n1847), .Z(n1851) );
  XNOR U1831 ( .A(n1853), .B(n1854), .Z(n1846) );
  NOR U1832 ( .A(n1855), .B(n1856), .Z(n1854) );
  XNOR U1833 ( .A(n1853), .B(n1857), .Z(n1855) );
  XOR U1834 ( .A(n1858), .B(n1859), .Z(n1803) );
  NOR U1835 ( .A(n1860), .B(n1861), .Z(n1859) );
  XNOR U1836 ( .A(n1858), .B(n1862), .Z(n1860) );
  XNOR U1837 ( .A(n1813), .B(n1804), .Z(n1845) );
  XOR U1838 ( .A(n1863), .B(n1864), .Z(n1804) );
  AND U1839 ( .A(n1865), .B(n1866), .Z(n1864) );
  XOR U1840 ( .A(n1863), .B(n1867), .Z(n1865) );
  XOR U1841 ( .A(n1868), .B(n1819), .Z(n1813) );
  XOR U1842 ( .A(n1869), .B(n1870), .Z(n1819) );
  NOR U1843 ( .A(n1871), .B(n1872), .Z(n1870) );
  XOR U1844 ( .A(n1869), .B(n1873), .Z(n1871) );
  XNOR U1845 ( .A(n1818), .B(n1810), .Z(n1868) );
  XOR U1846 ( .A(n1874), .B(n1875), .Z(n1810) );
  AND U1847 ( .A(n1876), .B(n1877), .Z(n1875) );
  XOR U1848 ( .A(n1874), .B(n1878), .Z(n1876) );
  XNOR U1849 ( .A(n1879), .B(n1815), .Z(n1818) );
  XOR U1850 ( .A(n1880), .B(n1881), .Z(n1815) );
  AND U1851 ( .A(n1882), .B(n1883), .Z(n1881) );
  XNOR U1852 ( .A(n1884), .B(n1885), .Z(n1882) );
  IV U1853 ( .A(n1880), .Z(n1884) );
  XNOR U1854 ( .A(n1886), .B(n1887), .Z(n1879) );
  NOR U1855 ( .A(n1888), .B(n1889), .Z(n1887) );
  XOR U1856 ( .A(n1886), .B(n1890), .Z(n1888) );
  XOR U1857 ( .A(n1808), .B(n1820), .Z(n1844) );
  NOR U1858 ( .A(n1744), .B(n1891), .Z(n1820) );
  XNOR U1859 ( .A(n1826), .B(n1825), .Z(n1808) );
  XNOR U1860 ( .A(n1892), .B(n1831), .Z(n1825) );
  XNOR U1861 ( .A(n1893), .B(n1894), .Z(n1831) );
  NOR U1862 ( .A(n1895), .B(n1896), .Z(n1894) );
  XOR U1863 ( .A(n1893), .B(n1897), .Z(n1895) );
  XNOR U1864 ( .A(n1830), .B(n1822), .Z(n1892) );
  XOR U1865 ( .A(n1898), .B(n1899), .Z(n1822) );
  AND U1866 ( .A(n1900), .B(n1901), .Z(n1899) );
  XNOR U1867 ( .A(n1898), .B(n1902), .Z(n1900) );
  XNOR U1868 ( .A(n1903), .B(n1827), .Z(n1830) );
  XOR U1869 ( .A(n1904), .B(n1905), .Z(n1827) );
  AND U1870 ( .A(n1906), .B(n1907), .Z(n1905) );
  XNOR U1871 ( .A(n1908), .B(n1909), .Z(n1906) );
  IV U1872 ( .A(n1904), .Z(n1908) );
  XNOR U1873 ( .A(n1910), .B(n1911), .Z(n1903) );
  NOR U1874 ( .A(n1912), .B(n1913), .Z(n1911) );
  XNOR U1875 ( .A(n1910), .B(n1914), .Z(n1912) );
  XOR U1876 ( .A(n1836), .B(n1835), .Z(n1826) );
  XNOR U1877 ( .A(n1915), .B(n1832), .Z(n1835) );
  XOR U1878 ( .A(n1916), .B(n1917), .Z(n1832) );
  AND U1879 ( .A(n1918), .B(n1919), .Z(n1917) );
  XOR U1880 ( .A(n1916), .B(n1920), .Z(n1918) );
  XNOR U1881 ( .A(n1921), .B(n1922), .Z(n1915) );
  NOR U1882 ( .A(n1923), .B(n1924), .Z(n1922) );
  XNOR U1883 ( .A(n1921), .B(n1925), .Z(n1923) );
  XOR U1884 ( .A(n1926), .B(n1927), .Z(n1836) );
  NOR U1885 ( .A(n1928), .B(n1929), .Z(n1927) );
  XNOR U1886 ( .A(n1926), .B(n1930), .Z(n1928) );
  XNOR U1887 ( .A(n1731), .B(n1840), .Z(n1842) );
  XNOR U1888 ( .A(n1931), .B(n1932), .Z(n1731) );
  AND U1889 ( .A(n66), .B(n1738), .Z(n1932) );
  XOR U1890 ( .A(n1931), .B(n1736), .Z(n1738) );
  AND U1891 ( .A(n1741), .B(n1744), .Z(n1840) );
  XOR U1892 ( .A(n1933), .B(n1891), .Z(n1744) );
  XNOR U1893 ( .A(p_input[0]), .B(p_input[256]), .Z(n1891) );
  XNOR U1894 ( .A(n1867), .B(n1866), .Z(n1933) );
  XNOR U1895 ( .A(n1934), .B(n1878), .Z(n1866) );
  XOR U1896 ( .A(n1852), .B(n1850), .Z(n1878) );
  XNOR U1897 ( .A(n1935), .B(n1857), .Z(n1850) );
  XOR U1898 ( .A(p_input[24]), .B(p_input[280]), .Z(n1857) );
  XOR U1899 ( .A(n1847), .B(n1856), .Z(n1935) );
  XOR U1900 ( .A(n1936), .B(n1853), .Z(n1856) );
  XOR U1901 ( .A(p_input[22]), .B(p_input[278]), .Z(n1853) );
  XOR U1902 ( .A(p_input[23]), .B(n1937), .Z(n1936) );
  XOR U1903 ( .A(p_input[18]), .B(p_input[274]), .Z(n1847) );
  XNOR U1904 ( .A(n1862), .B(n1861), .Z(n1852) );
  XOR U1905 ( .A(n1938), .B(n1858), .Z(n1861) );
  XOR U1906 ( .A(p_input[19]), .B(p_input[275]), .Z(n1858) );
  XOR U1907 ( .A(p_input[20]), .B(n1939), .Z(n1938) );
  XOR U1908 ( .A(p_input[21]), .B(p_input[277]), .Z(n1862) );
  XOR U1909 ( .A(n1877), .B(n1940), .Z(n1934) );
  IV U1910 ( .A(n1863), .Z(n1940) );
  XOR U1911 ( .A(p_input[1]), .B(p_input[257]), .Z(n1863) );
  XNOR U1912 ( .A(n1941), .B(n1885), .Z(n1877) );
  XNOR U1913 ( .A(n1873), .B(n1872), .Z(n1885) );
  XNOR U1914 ( .A(n1942), .B(n1869), .Z(n1872) );
  XNOR U1915 ( .A(p_input[26]), .B(p_input[282]), .Z(n1869) );
  XOR U1916 ( .A(p_input[27]), .B(n1943), .Z(n1942) );
  XOR U1917 ( .A(p_input[284]), .B(p_input[28]), .Z(n1873) );
  XOR U1918 ( .A(n1883), .B(n1944), .Z(n1941) );
  IV U1919 ( .A(n1874), .Z(n1944) );
  XOR U1920 ( .A(p_input[17]), .B(p_input[273]), .Z(n1874) );
  XOR U1921 ( .A(n1945), .B(n1890), .Z(n1883) );
  XNOR U1922 ( .A(p_input[287]), .B(p_input[31]), .Z(n1890) );
  XOR U1923 ( .A(n1880), .B(n1889), .Z(n1945) );
  XOR U1924 ( .A(n1946), .B(n1886), .Z(n1889) );
  XOR U1925 ( .A(p_input[285]), .B(p_input[29]), .Z(n1886) );
  XNOR U1926 ( .A(p_input[286]), .B(p_input[30]), .Z(n1946) );
  XOR U1927 ( .A(p_input[25]), .B(p_input[281]), .Z(n1880) );
  XNOR U1928 ( .A(n1902), .B(n1901), .Z(n1867) );
  XNOR U1929 ( .A(n1947), .B(n1909), .Z(n1901) );
  XNOR U1930 ( .A(n1897), .B(n1896), .Z(n1909) );
  XNOR U1931 ( .A(n1948), .B(n1893), .Z(n1896) );
  XNOR U1932 ( .A(p_input[11]), .B(p_input[267]), .Z(n1893) );
  XOR U1933 ( .A(p_input[12]), .B(n1949), .Z(n1948) );
  XOR U1934 ( .A(p_input[13]), .B(p_input[269]), .Z(n1897) );
  XNOR U1935 ( .A(n1907), .B(n1898), .Z(n1947) );
  XOR U1936 ( .A(p_input[258]), .B(p_input[2]), .Z(n1898) );
  XNOR U1937 ( .A(n1950), .B(n1914), .Z(n1907) );
  XNOR U1938 ( .A(p_input[16]), .B(n1951), .Z(n1914) );
  XOR U1939 ( .A(n1904), .B(n1913), .Z(n1950) );
  XOR U1940 ( .A(n1952), .B(n1910), .Z(n1913) );
  XOR U1941 ( .A(p_input[14]), .B(p_input[270]), .Z(n1910) );
  XOR U1942 ( .A(p_input[15]), .B(n1953), .Z(n1952) );
  XOR U1943 ( .A(p_input[10]), .B(p_input[266]), .Z(n1904) );
  XNOR U1944 ( .A(n1920), .B(n1919), .Z(n1902) );
  XNOR U1945 ( .A(n1954), .B(n1925), .Z(n1919) );
  XOR U1946 ( .A(p_input[265]), .B(p_input[9]), .Z(n1925) );
  XOR U1947 ( .A(n1916), .B(n1924), .Z(n1954) );
  XOR U1948 ( .A(n1955), .B(n1921), .Z(n1924) );
  XOR U1949 ( .A(p_input[263]), .B(p_input[7]), .Z(n1921) );
  XNOR U1950 ( .A(p_input[264]), .B(p_input[8]), .Z(n1955) );
  XOR U1951 ( .A(p_input[259]), .B(p_input[3]), .Z(n1916) );
  XNOR U1952 ( .A(n1930), .B(n1929), .Z(n1920) );
  XOR U1953 ( .A(n1956), .B(n1926), .Z(n1929) );
  XOR U1954 ( .A(p_input[260]), .B(p_input[4]), .Z(n1926) );
  XNOR U1955 ( .A(p_input[261]), .B(p_input[5]), .Z(n1956) );
  XOR U1956 ( .A(p_input[262]), .B(p_input[6]), .Z(n1930) );
  XNOR U1957 ( .A(n1957), .B(n1958), .Z(n1741) );
  AND U1958 ( .A(n66), .B(n1959), .Z(n1958) );
  XNOR U1959 ( .A(n1960), .B(n1961), .Z(n66) );
  AND U1960 ( .A(n1962), .B(n1963), .Z(n1961) );
  XOR U1961 ( .A(n1960), .B(n1751), .Z(n1963) );
  XNOR U1962 ( .A(n1960), .B(n1684), .Z(n1962) );
  XOR U1963 ( .A(n1964), .B(n1965), .Z(n1960) );
  AND U1964 ( .A(n1966), .B(n1967), .Z(n1965) );
  XNOR U1965 ( .A(n1764), .B(n1964), .Z(n1967) );
  XOR U1966 ( .A(n1964), .B(n1766), .Z(n1966) );
  XOR U1967 ( .A(n1968), .B(n1969), .Z(n1964) );
  AND U1968 ( .A(n1970), .B(n1971), .Z(n1969) );
  XNOR U1969 ( .A(n1790), .B(n1968), .Z(n1971) );
  XOR U1970 ( .A(n1968), .B(n1792), .Z(n1970) );
  IV U1971 ( .A(n1710), .Z(n1792) );
  XOR U1972 ( .A(n1972), .B(n1973), .Z(n1968) );
  AND U1973 ( .A(n1974), .B(n1975), .Z(n1973) );
  XOR U1974 ( .A(n1972), .B(n1839), .Z(n1974) );
  XOR U1975 ( .A(n1976), .B(n1977), .Z(n1739) );
  AND U1976 ( .A(n70), .B(n1959), .Z(n1977) );
  XNOR U1977 ( .A(n1957), .B(n1976), .Z(n1959) );
  XNOR U1978 ( .A(n1978), .B(n1979), .Z(n70) );
  AND U1979 ( .A(n1980), .B(n1981), .Z(n1979) );
  XNOR U1980 ( .A(n1982), .B(n1978), .Z(n1981) );
  IV U1981 ( .A(n1751), .Z(n1982) );
  XNOR U1982 ( .A(n1983), .B(n1984), .Z(n1751) );
  AND U1983 ( .A(n74), .B(n1985), .Z(n1984) );
  XNOR U1984 ( .A(n1983), .B(n1986), .Z(n1985) );
  XNOR U1985 ( .A(n1684), .B(n1978), .Z(n1980) );
  XNOR U1986 ( .A(n1987), .B(n1988), .Z(n1684) );
  AND U1987 ( .A(n82), .B(n1989), .Z(n1988) );
  XNOR U1988 ( .A(n1990), .B(n1991), .Z(n1989) );
  XOR U1989 ( .A(n1992), .B(n1993), .Z(n1978) );
  AND U1990 ( .A(n1994), .B(n1995), .Z(n1993) );
  XNOR U1991 ( .A(n1992), .B(n1764), .Z(n1995) );
  XNOR U1992 ( .A(n1996), .B(n1997), .Z(n1764) );
  AND U1993 ( .A(n74), .B(n1998), .Z(n1997) );
  XOR U1994 ( .A(n1999), .B(n1996), .Z(n1998) );
  XNOR U1995 ( .A(n1697), .B(n1992), .Z(n1994) );
  IV U1996 ( .A(n1766), .Z(n1697) );
  XOR U1997 ( .A(n2000), .B(n2001), .Z(n1766) );
  AND U1998 ( .A(n82), .B(n2002), .Z(n2001) );
  XOR U1999 ( .A(n2003), .B(n2004), .Z(n1992) );
  AND U2000 ( .A(n2005), .B(n2006), .Z(n2004) );
  XNOR U2001 ( .A(n2003), .B(n1790), .Z(n2006) );
  XNOR U2002 ( .A(n2007), .B(n2008), .Z(n1790) );
  AND U2003 ( .A(n74), .B(n2009), .Z(n2008) );
  XNOR U2004 ( .A(n2010), .B(n2007), .Z(n2009) );
  XNOR U2005 ( .A(n1710), .B(n2003), .Z(n2005) );
  XNOR U2006 ( .A(n2011), .B(n2012), .Z(n1710) );
  AND U2007 ( .A(n82), .B(n2013), .Z(n2012) );
  XOR U2008 ( .A(n1972), .B(n2014), .Z(n2003) );
  AND U2009 ( .A(n2015), .B(n1975), .Z(n2014) );
  XNOR U2010 ( .A(n1837), .B(n1972), .Z(n1975) );
  XNOR U2011 ( .A(n2016), .B(n2017), .Z(n1837) );
  AND U2012 ( .A(n74), .B(n2018), .Z(n2017) );
  XOR U2013 ( .A(n2019), .B(n2016), .Z(n2018) );
  XNOR U2014 ( .A(n1723), .B(n1972), .Z(n2015) );
  IV U2015 ( .A(n1839), .Z(n1723) );
  XOR U2016 ( .A(n2020), .B(n2021), .Z(n1839) );
  AND U2017 ( .A(n82), .B(n2022), .Z(n2021) );
  XOR U2018 ( .A(n2023), .B(n2024), .Z(n1972) );
  AND U2019 ( .A(n2025), .B(n2026), .Z(n2024) );
  XNOR U2020 ( .A(n2023), .B(n1931), .Z(n2026) );
  XNOR U2021 ( .A(n2027), .B(n2028), .Z(n1931) );
  AND U2022 ( .A(n74), .B(n2029), .Z(n2028) );
  XNOR U2023 ( .A(n2030), .B(n2027), .Z(n2029) );
  XNOR U2024 ( .A(n2031), .B(n2023), .Z(n2025) );
  IV U2025 ( .A(n1736), .Z(n2031) );
  XOR U2026 ( .A(n2032), .B(n2033), .Z(n1736) );
  AND U2027 ( .A(n82), .B(n2034), .Z(n2033) );
  AND U2028 ( .A(n1976), .B(n1957), .Z(n2023) );
  XNOR U2029 ( .A(n2035), .B(n2036), .Z(n1957) );
  AND U2030 ( .A(n74), .B(n2037), .Z(n2036) );
  XNOR U2031 ( .A(n2038), .B(n2035), .Z(n2037) );
  XNOR U2032 ( .A(n2039), .B(n2040), .Z(n74) );
  AND U2033 ( .A(n2041), .B(n2042), .Z(n2040) );
  XOR U2034 ( .A(n1986), .B(n2039), .Z(n2042) );
  AND U2035 ( .A(n2043), .B(n2044), .Z(n1986) );
  XOR U2036 ( .A(n2039), .B(n1983), .Z(n2041) );
  XOR U2037 ( .A(n1990), .B(n2045), .Z(n1983) );
  AND U2038 ( .A(n78), .B(n2046), .Z(n2045) );
  XOR U2039 ( .A(n1990), .B(n1987), .Z(n2046) );
  XOR U2040 ( .A(n2047), .B(n2048), .Z(n2039) );
  AND U2041 ( .A(n2049), .B(n2050), .Z(n2048) );
  XNOR U2042 ( .A(n2047), .B(n2043), .Z(n2050) );
  IV U2043 ( .A(n1999), .Z(n2043) );
  XOR U2044 ( .A(n2051), .B(n2052), .Z(n1999) );
  XOR U2045 ( .A(n2053), .B(n2044), .Z(n2052) );
  AND U2046 ( .A(n2010), .B(n2054), .Z(n2044) );
  AND U2047 ( .A(n2055), .B(n2056), .Z(n2053) );
  XOR U2048 ( .A(n2057), .B(n2051), .Z(n2055) );
  XNOR U2049 ( .A(n1996), .B(n2047), .Z(n2049) );
  XNOR U2050 ( .A(n2058), .B(n2059), .Z(n1996) );
  AND U2051 ( .A(n78), .B(n2002), .Z(n2059) );
  XOR U2052 ( .A(n2058), .B(n2000), .Z(n2002) );
  XOR U2053 ( .A(n2060), .B(n2061), .Z(n2047) );
  AND U2054 ( .A(n2062), .B(n2063), .Z(n2061) );
  XNOR U2055 ( .A(n2060), .B(n2010), .Z(n2063) );
  XOR U2056 ( .A(n2064), .B(n2056), .Z(n2010) );
  XNOR U2057 ( .A(n2065), .B(n2051), .Z(n2056) );
  XOR U2058 ( .A(n2066), .B(n2067), .Z(n2051) );
  AND U2059 ( .A(n2068), .B(n2069), .Z(n2067) );
  XOR U2060 ( .A(n2070), .B(n2066), .Z(n2068) );
  XNOR U2061 ( .A(n2071), .B(n2072), .Z(n2065) );
  AND U2062 ( .A(n2073), .B(n2074), .Z(n2072) );
  XOR U2063 ( .A(n2071), .B(n2075), .Z(n2073) );
  XNOR U2064 ( .A(n2057), .B(n2054), .Z(n2064) );
  AND U2065 ( .A(n2076), .B(n2077), .Z(n2054) );
  XOR U2066 ( .A(n2078), .B(n2079), .Z(n2057) );
  AND U2067 ( .A(n2080), .B(n2081), .Z(n2079) );
  XOR U2068 ( .A(n2078), .B(n2082), .Z(n2080) );
  XNOR U2069 ( .A(n2007), .B(n2060), .Z(n2062) );
  XNOR U2070 ( .A(n2083), .B(n2084), .Z(n2007) );
  AND U2071 ( .A(n78), .B(n2013), .Z(n2084) );
  XOR U2072 ( .A(n2083), .B(n2011), .Z(n2013) );
  XOR U2073 ( .A(n2085), .B(n2086), .Z(n2060) );
  AND U2074 ( .A(n2087), .B(n2088), .Z(n2086) );
  XNOR U2075 ( .A(n2085), .B(n2076), .Z(n2088) );
  IV U2076 ( .A(n2019), .Z(n2076) );
  XNOR U2077 ( .A(n2089), .B(n2069), .Z(n2019) );
  XNOR U2078 ( .A(n2090), .B(n2075), .Z(n2069) );
  XOR U2079 ( .A(n2091), .B(n2092), .Z(n2075) );
  AND U2080 ( .A(n2093), .B(n2094), .Z(n2092) );
  XOR U2081 ( .A(n2091), .B(n2095), .Z(n2093) );
  XNOR U2082 ( .A(n2074), .B(n2066), .Z(n2090) );
  XOR U2083 ( .A(n2096), .B(n2097), .Z(n2066) );
  AND U2084 ( .A(n2098), .B(n2099), .Z(n2097) );
  XNOR U2085 ( .A(n2100), .B(n2096), .Z(n2098) );
  XNOR U2086 ( .A(n2101), .B(n2071), .Z(n2074) );
  XOR U2087 ( .A(n2102), .B(n2103), .Z(n2071) );
  AND U2088 ( .A(n2104), .B(n2105), .Z(n2103) );
  XOR U2089 ( .A(n2102), .B(n2106), .Z(n2104) );
  XNOR U2090 ( .A(n2107), .B(n2108), .Z(n2101) );
  AND U2091 ( .A(n2109), .B(n2110), .Z(n2108) );
  XNOR U2092 ( .A(n2107), .B(n2111), .Z(n2109) );
  XNOR U2093 ( .A(n2070), .B(n2077), .Z(n2089) );
  AND U2094 ( .A(n2030), .B(n2112), .Z(n2077) );
  XOR U2095 ( .A(n2082), .B(n2081), .Z(n2070) );
  XNOR U2096 ( .A(n2113), .B(n2078), .Z(n2081) );
  XOR U2097 ( .A(n2114), .B(n2115), .Z(n2078) );
  AND U2098 ( .A(n2116), .B(n2117), .Z(n2115) );
  XOR U2099 ( .A(n2114), .B(n2118), .Z(n2116) );
  XNOR U2100 ( .A(n2119), .B(n2120), .Z(n2113) );
  AND U2101 ( .A(n2121), .B(n2122), .Z(n2120) );
  XOR U2102 ( .A(n2119), .B(n2123), .Z(n2121) );
  XOR U2103 ( .A(n2124), .B(n2125), .Z(n2082) );
  AND U2104 ( .A(n2126), .B(n2127), .Z(n2125) );
  XOR U2105 ( .A(n2124), .B(n2128), .Z(n2126) );
  XNOR U2106 ( .A(n2016), .B(n2085), .Z(n2087) );
  XNOR U2107 ( .A(n2129), .B(n2130), .Z(n2016) );
  AND U2108 ( .A(n78), .B(n2022), .Z(n2130) );
  XOR U2109 ( .A(n2129), .B(n2020), .Z(n2022) );
  XOR U2110 ( .A(n2131), .B(n2132), .Z(n2085) );
  AND U2111 ( .A(n2133), .B(n2134), .Z(n2132) );
  XNOR U2112 ( .A(n2131), .B(n2030), .Z(n2134) );
  XOR U2113 ( .A(n2135), .B(n2099), .Z(n2030) );
  XNOR U2114 ( .A(n2136), .B(n2106), .Z(n2099) );
  XOR U2115 ( .A(n2095), .B(n2094), .Z(n2106) );
  XNOR U2116 ( .A(n2137), .B(n2091), .Z(n2094) );
  XOR U2117 ( .A(n2138), .B(n2139), .Z(n2091) );
  AND U2118 ( .A(n2140), .B(n2141), .Z(n2139) );
  XOR U2119 ( .A(n2138), .B(n2142), .Z(n2140) );
  XNOR U2120 ( .A(n2143), .B(n2144), .Z(n2137) );
  NOR U2121 ( .A(n2145), .B(n2146), .Z(n2144) );
  XNOR U2122 ( .A(n2143), .B(n2147), .Z(n2145) );
  XOR U2123 ( .A(n2148), .B(n2149), .Z(n2095) );
  NOR U2124 ( .A(n2150), .B(n2151), .Z(n2149) );
  XNOR U2125 ( .A(n2148), .B(n2152), .Z(n2150) );
  XNOR U2126 ( .A(n2105), .B(n2096), .Z(n2136) );
  XOR U2127 ( .A(n2153), .B(n2154), .Z(n2096) );
  NOR U2128 ( .A(n2155), .B(n2156), .Z(n2154) );
  XNOR U2129 ( .A(n2153), .B(n2157), .Z(n2155) );
  XOR U2130 ( .A(n2158), .B(n2111), .Z(n2105) );
  XNOR U2131 ( .A(n2159), .B(n2160), .Z(n2111) );
  NOR U2132 ( .A(n2161), .B(n2162), .Z(n2160) );
  XNOR U2133 ( .A(n2159), .B(n2163), .Z(n2161) );
  XNOR U2134 ( .A(n2110), .B(n2102), .Z(n2158) );
  XOR U2135 ( .A(n2164), .B(n2165), .Z(n2102) );
  AND U2136 ( .A(n2166), .B(n2167), .Z(n2165) );
  XOR U2137 ( .A(n2164), .B(n2168), .Z(n2166) );
  XNOR U2138 ( .A(n2169), .B(n2107), .Z(n2110) );
  XOR U2139 ( .A(n2170), .B(n2171), .Z(n2107) );
  AND U2140 ( .A(n2172), .B(n2173), .Z(n2171) );
  XOR U2141 ( .A(n2170), .B(n2174), .Z(n2172) );
  XNOR U2142 ( .A(n2175), .B(n2176), .Z(n2169) );
  NOR U2143 ( .A(n2177), .B(n2178), .Z(n2176) );
  XOR U2144 ( .A(n2175), .B(n2179), .Z(n2177) );
  XOR U2145 ( .A(n2100), .B(n2112), .Z(n2135) );
  NOR U2146 ( .A(n2038), .B(n2180), .Z(n2112) );
  XNOR U2147 ( .A(n2118), .B(n2117), .Z(n2100) );
  XNOR U2148 ( .A(n2181), .B(n2123), .Z(n2117) );
  XOR U2149 ( .A(n2182), .B(n2183), .Z(n2123) );
  NOR U2150 ( .A(n2184), .B(n2185), .Z(n2183) );
  XNOR U2151 ( .A(n2182), .B(n2186), .Z(n2184) );
  XNOR U2152 ( .A(n2122), .B(n2114), .Z(n2181) );
  XOR U2153 ( .A(n2187), .B(n2188), .Z(n2114) );
  AND U2154 ( .A(n2189), .B(n2190), .Z(n2188) );
  XNOR U2155 ( .A(n2187), .B(n2191), .Z(n2189) );
  XNOR U2156 ( .A(n2192), .B(n2119), .Z(n2122) );
  XOR U2157 ( .A(n2193), .B(n2194), .Z(n2119) );
  AND U2158 ( .A(n2195), .B(n2196), .Z(n2194) );
  XOR U2159 ( .A(n2193), .B(n2197), .Z(n2195) );
  XNOR U2160 ( .A(n2198), .B(n2199), .Z(n2192) );
  NOR U2161 ( .A(n2200), .B(n2201), .Z(n2199) );
  XOR U2162 ( .A(n2198), .B(n2202), .Z(n2200) );
  XOR U2163 ( .A(n2128), .B(n2127), .Z(n2118) );
  XNOR U2164 ( .A(n2203), .B(n2124), .Z(n2127) );
  XOR U2165 ( .A(n2204), .B(n2205), .Z(n2124) );
  AND U2166 ( .A(n2206), .B(n2207), .Z(n2205) );
  XOR U2167 ( .A(n2204), .B(n2208), .Z(n2206) );
  XNOR U2168 ( .A(n2209), .B(n2210), .Z(n2203) );
  NOR U2169 ( .A(n2211), .B(n2212), .Z(n2210) );
  XNOR U2170 ( .A(n2209), .B(n2213), .Z(n2211) );
  XOR U2171 ( .A(n2214), .B(n2215), .Z(n2128) );
  NOR U2172 ( .A(n2216), .B(n2217), .Z(n2215) );
  XNOR U2173 ( .A(n2214), .B(n2218), .Z(n2216) );
  XNOR U2174 ( .A(n2027), .B(n2131), .Z(n2133) );
  XNOR U2175 ( .A(n2219), .B(n2220), .Z(n2027) );
  AND U2176 ( .A(n78), .B(n2034), .Z(n2220) );
  XOR U2177 ( .A(n2219), .B(n2032), .Z(n2034) );
  AND U2178 ( .A(n2035), .B(n2038), .Z(n2131) );
  XOR U2179 ( .A(n2221), .B(n2180), .Z(n2038) );
  XNOR U2180 ( .A(p_input[256]), .B(p_input[32]), .Z(n2180) );
  XOR U2181 ( .A(n2157), .B(n2156), .Z(n2221) );
  XOR U2182 ( .A(n2222), .B(n2168), .Z(n2156) );
  XOR U2183 ( .A(n2142), .B(n2141), .Z(n2168) );
  XNOR U2184 ( .A(n2223), .B(n2147), .Z(n2141) );
  XOR U2185 ( .A(p_input[280]), .B(p_input[56]), .Z(n2147) );
  XOR U2186 ( .A(n2138), .B(n2146), .Z(n2223) );
  XOR U2187 ( .A(n2224), .B(n2143), .Z(n2146) );
  XOR U2188 ( .A(p_input[278]), .B(p_input[54]), .Z(n2143) );
  XNOR U2189 ( .A(p_input[279]), .B(p_input[55]), .Z(n2224) );
  XNOR U2190 ( .A(n2225), .B(p_input[50]), .Z(n2138) );
  XNOR U2191 ( .A(n2152), .B(n2151), .Z(n2142) );
  XOR U2192 ( .A(n2226), .B(n2148), .Z(n2151) );
  XOR U2193 ( .A(p_input[275]), .B(p_input[51]), .Z(n2148) );
  XNOR U2194 ( .A(p_input[276]), .B(p_input[52]), .Z(n2226) );
  XOR U2195 ( .A(p_input[277]), .B(p_input[53]), .Z(n2152) );
  XNOR U2196 ( .A(n2167), .B(n2153), .Z(n2222) );
  XNOR U2197 ( .A(n2227), .B(p_input[33]), .Z(n2153) );
  XNOR U2198 ( .A(n2228), .B(n2174), .Z(n2167) );
  XNOR U2199 ( .A(n2163), .B(n2162), .Z(n2174) );
  XOR U2200 ( .A(n2229), .B(n2159), .Z(n2162) );
  XNOR U2201 ( .A(n2230), .B(p_input[58]), .Z(n2159) );
  XNOR U2202 ( .A(p_input[283]), .B(p_input[59]), .Z(n2229) );
  XOR U2203 ( .A(p_input[284]), .B(p_input[60]), .Z(n2163) );
  XNOR U2204 ( .A(n2173), .B(n2164), .Z(n2228) );
  XNOR U2205 ( .A(n2231), .B(p_input[49]), .Z(n2164) );
  XOR U2206 ( .A(n2232), .B(n2179), .Z(n2173) );
  XNOR U2207 ( .A(p_input[287]), .B(p_input[63]), .Z(n2179) );
  XOR U2208 ( .A(n2170), .B(n2178), .Z(n2232) );
  XOR U2209 ( .A(n2233), .B(n2175), .Z(n2178) );
  XOR U2210 ( .A(p_input[285]), .B(p_input[61]), .Z(n2175) );
  XNOR U2211 ( .A(p_input[286]), .B(p_input[62]), .Z(n2233) );
  XNOR U2212 ( .A(n2234), .B(p_input[57]), .Z(n2170) );
  XNOR U2213 ( .A(n2191), .B(n2190), .Z(n2157) );
  XNOR U2214 ( .A(n2235), .B(n2197), .Z(n2190) );
  XNOR U2215 ( .A(n2186), .B(n2185), .Z(n2197) );
  XOR U2216 ( .A(n2236), .B(n2182), .Z(n2185) );
  XNOR U2217 ( .A(n2237), .B(p_input[43]), .Z(n2182) );
  XNOR U2218 ( .A(p_input[268]), .B(p_input[44]), .Z(n2236) );
  XOR U2219 ( .A(p_input[269]), .B(p_input[45]), .Z(n2186) );
  XNOR U2220 ( .A(n2196), .B(n2187), .Z(n2235) );
  XOR U2221 ( .A(p_input[258]), .B(p_input[34]), .Z(n2187) );
  XOR U2222 ( .A(n2238), .B(n2202), .Z(n2196) );
  XNOR U2223 ( .A(p_input[272]), .B(p_input[48]), .Z(n2202) );
  XOR U2224 ( .A(n2193), .B(n2201), .Z(n2238) );
  XOR U2225 ( .A(n2239), .B(n2198), .Z(n2201) );
  XOR U2226 ( .A(p_input[270]), .B(p_input[46]), .Z(n2198) );
  XNOR U2227 ( .A(p_input[271]), .B(p_input[47]), .Z(n2239) );
  XNOR U2228 ( .A(n2240), .B(p_input[42]), .Z(n2193) );
  XNOR U2229 ( .A(n2208), .B(n2207), .Z(n2191) );
  XNOR U2230 ( .A(n2241), .B(n2213), .Z(n2207) );
  XOR U2231 ( .A(p_input[265]), .B(p_input[41]), .Z(n2213) );
  XOR U2232 ( .A(n2204), .B(n2212), .Z(n2241) );
  XOR U2233 ( .A(n2242), .B(n2209), .Z(n2212) );
  XOR U2234 ( .A(p_input[263]), .B(p_input[39]), .Z(n2209) );
  XNOR U2235 ( .A(p_input[264]), .B(p_input[40]), .Z(n2242) );
  XOR U2236 ( .A(p_input[259]), .B(p_input[35]), .Z(n2204) );
  XNOR U2237 ( .A(n2218), .B(n2217), .Z(n2208) );
  XOR U2238 ( .A(n2243), .B(n2214), .Z(n2217) );
  XOR U2239 ( .A(p_input[260]), .B(p_input[36]), .Z(n2214) );
  XNOR U2240 ( .A(p_input[261]), .B(p_input[37]), .Z(n2243) );
  XOR U2241 ( .A(p_input[262]), .B(p_input[38]), .Z(n2218) );
  XNOR U2242 ( .A(n2244), .B(n2245), .Z(n2035) );
  AND U2243 ( .A(n78), .B(n2246), .Z(n2245) );
  XNOR U2244 ( .A(n2247), .B(n2248), .Z(n78) );
  AND U2245 ( .A(n2249), .B(n2250), .Z(n2248) );
  XNOR U2246 ( .A(n2247), .B(n1990), .Z(n2250) );
  XOR U2247 ( .A(n2247), .B(n1987), .Z(n2249) );
  XOR U2248 ( .A(n2251), .B(n2252), .Z(n2247) );
  AND U2249 ( .A(n2253), .B(n2254), .Z(n2252) );
  XNOR U2250 ( .A(n2058), .B(n2251), .Z(n2254) );
  XOR U2251 ( .A(n2251), .B(n2000), .Z(n2253) );
  XOR U2252 ( .A(n2255), .B(n2256), .Z(n2251) );
  AND U2253 ( .A(n2257), .B(n2258), .Z(n2256) );
  XNOR U2254 ( .A(n2083), .B(n2255), .Z(n2258) );
  XOR U2255 ( .A(n2255), .B(n2011), .Z(n2257) );
  XOR U2256 ( .A(n2259), .B(n2260), .Z(n2255) );
  AND U2257 ( .A(n2261), .B(n2262), .Z(n2260) );
  XOR U2258 ( .A(n2259), .B(n2020), .Z(n2261) );
  XOR U2259 ( .A(n2263), .B(n2264), .Z(n1976) );
  AND U2260 ( .A(n82), .B(n2246), .Z(n2264) );
  XNOR U2261 ( .A(n2244), .B(n2263), .Z(n2246) );
  XNOR U2262 ( .A(n2265), .B(n2266), .Z(n82) );
  AND U2263 ( .A(n2267), .B(n2268), .Z(n2266) );
  XNOR U2264 ( .A(n1990), .B(n2265), .Z(n2268) );
  XOR U2265 ( .A(n2269), .B(n2270), .Z(n1990) );
  AND U2266 ( .A(n2271), .B(n85), .Z(n2270) );
  NOR U2267 ( .A(n2272), .B(n2269), .Z(n2271) );
  XOR U2268 ( .A(n2265), .B(n1987), .Z(n2267) );
  IV U2269 ( .A(n1991), .Z(n1987) );
  AND U2270 ( .A(n2273), .B(n2274), .Z(n1991) );
  XOR U2271 ( .A(n2275), .B(n2276), .Z(n2265) );
  AND U2272 ( .A(n2277), .B(n2278), .Z(n2276) );
  XNOR U2273 ( .A(n2275), .B(n2058), .Z(n2278) );
  XNOR U2274 ( .A(n2279), .B(n2280), .Z(n2058) );
  AND U2275 ( .A(n85), .B(n2281), .Z(n2280) );
  XOR U2276 ( .A(n2282), .B(n2279), .Z(n2281) );
  XNOR U2277 ( .A(n2283), .B(n2275), .Z(n2277) );
  IV U2278 ( .A(n2000), .Z(n2283) );
  XOR U2279 ( .A(n2284), .B(n2285), .Z(n2000) );
  AND U2280 ( .A(n93), .B(n2286), .Z(n2285) );
  XOR U2281 ( .A(n2287), .B(n2288), .Z(n2275) );
  AND U2282 ( .A(n2289), .B(n2290), .Z(n2288) );
  XNOR U2283 ( .A(n2287), .B(n2083), .Z(n2290) );
  XNOR U2284 ( .A(n2291), .B(n2292), .Z(n2083) );
  AND U2285 ( .A(n85), .B(n2293), .Z(n2292) );
  XNOR U2286 ( .A(n2294), .B(n2291), .Z(n2293) );
  XOR U2287 ( .A(n2011), .B(n2287), .Z(n2289) );
  XOR U2288 ( .A(n2295), .B(n2296), .Z(n2011) );
  AND U2289 ( .A(n93), .B(n2297), .Z(n2296) );
  XOR U2290 ( .A(n2259), .B(n2298), .Z(n2287) );
  AND U2291 ( .A(n2299), .B(n2262), .Z(n2298) );
  XNOR U2292 ( .A(n2129), .B(n2259), .Z(n2262) );
  XNOR U2293 ( .A(n2300), .B(n2301), .Z(n2129) );
  AND U2294 ( .A(n85), .B(n2302), .Z(n2301) );
  XOR U2295 ( .A(n2303), .B(n2300), .Z(n2302) );
  XNOR U2296 ( .A(n2304), .B(n2259), .Z(n2299) );
  IV U2297 ( .A(n2020), .Z(n2304) );
  XOR U2298 ( .A(n2305), .B(n2306), .Z(n2020) );
  AND U2299 ( .A(n93), .B(n2307), .Z(n2306) );
  XOR U2300 ( .A(n2308), .B(n2309), .Z(n2259) );
  AND U2301 ( .A(n2310), .B(n2311), .Z(n2309) );
  XNOR U2302 ( .A(n2308), .B(n2219), .Z(n2311) );
  XNOR U2303 ( .A(n2312), .B(n2313), .Z(n2219) );
  AND U2304 ( .A(n85), .B(n2314), .Z(n2313) );
  XNOR U2305 ( .A(n2315), .B(n2312), .Z(n2314) );
  XNOR U2306 ( .A(n2316), .B(n2308), .Z(n2310) );
  IV U2307 ( .A(n2032), .Z(n2316) );
  XOR U2308 ( .A(n2317), .B(n2318), .Z(n2032) );
  AND U2309 ( .A(n93), .B(n2319), .Z(n2318) );
  AND U2310 ( .A(n2263), .B(n2244), .Z(n2308) );
  XNOR U2311 ( .A(n2320), .B(n2321), .Z(n2244) );
  AND U2312 ( .A(n85), .B(n2322), .Z(n2321) );
  XNOR U2313 ( .A(n2323), .B(n2320), .Z(n2322) );
  XNOR U2314 ( .A(n2324), .B(n2325), .Z(n85) );
  NOR U2315 ( .A(n2326), .B(n2327), .Z(n2325) );
  XNOR U2316 ( .A(n2324), .B(n2269), .Z(n2327) );
  NOR U2317 ( .A(n2273), .B(n2274), .Z(n2269) );
  NOR U2318 ( .A(n2324), .B(n2272), .Z(n2326) );
  AND U2319 ( .A(n2328), .B(n2329), .Z(n2272) );
  XOR U2320 ( .A(n2330), .B(n2331), .Z(n2324) );
  AND U2321 ( .A(n2332), .B(n2333), .Z(n2331) );
  XNOR U2322 ( .A(n2330), .B(n2328), .Z(n2333) );
  IV U2323 ( .A(n2282), .Z(n2328) );
  XOR U2324 ( .A(n2334), .B(n2335), .Z(n2282) );
  XOR U2325 ( .A(n2336), .B(n2329), .Z(n2335) );
  AND U2326 ( .A(n2294), .B(n2337), .Z(n2329) );
  AND U2327 ( .A(n2338), .B(n2339), .Z(n2336) );
  XOR U2328 ( .A(n2340), .B(n2334), .Z(n2338) );
  XNOR U2329 ( .A(n2279), .B(n2330), .Z(n2332) );
  XNOR U2330 ( .A(n2341), .B(n2342), .Z(n2279) );
  AND U2331 ( .A(n89), .B(n2286), .Z(n2342) );
  XOR U2332 ( .A(n2341), .B(n2284), .Z(n2286) );
  XOR U2333 ( .A(n2343), .B(n2344), .Z(n2330) );
  AND U2334 ( .A(n2345), .B(n2346), .Z(n2344) );
  XNOR U2335 ( .A(n2343), .B(n2294), .Z(n2346) );
  XOR U2336 ( .A(n2347), .B(n2339), .Z(n2294) );
  XNOR U2337 ( .A(n2348), .B(n2334), .Z(n2339) );
  XOR U2338 ( .A(n2349), .B(n2350), .Z(n2334) );
  AND U2339 ( .A(n2351), .B(n2352), .Z(n2350) );
  XOR U2340 ( .A(n2353), .B(n2349), .Z(n2351) );
  XNOR U2341 ( .A(n2354), .B(n2355), .Z(n2348) );
  AND U2342 ( .A(n2356), .B(n2357), .Z(n2355) );
  XOR U2343 ( .A(n2354), .B(n2358), .Z(n2356) );
  XNOR U2344 ( .A(n2340), .B(n2337), .Z(n2347) );
  AND U2345 ( .A(n2359), .B(n2360), .Z(n2337) );
  XOR U2346 ( .A(n2361), .B(n2362), .Z(n2340) );
  AND U2347 ( .A(n2363), .B(n2364), .Z(n2362) );
  XOR U2348 ( .A(n2361), .B(n2365), .Z(n2363) );
  XNOR U2349 ( .A(n2291), .B(n2343), .Z(n2345) );
  XNOR U2350 ( .A(n2366), .B(n2367), .Z(n2291) );
  AND U2351 ( .A(n89), .B(n2297), .Z(n2367) );
  XOR U2352 ( .A(n2366), .B(n2295), .Z(n2297) );
  XOR U2353 ( .A(n2368), .B(n2369), .Z(n2343) );
  AND U2354 ( .A(n2370), .B(n2371), .Z(n2369) );
  XNOR U2355 ( .A(n2368), .B(n2359), .Z(n2371) );
  IV U2356 ( .A(n2303), .Z(n2359) );
  XNOR U2357 ( .A(n2372), .B(n2352), .Z(n2303) );
  XNOR U2358 ( .A(n2373), .B(n2358), .Z(n2352) );
  XOR U2359 ( .A(n2374), .B(n2375), .Z(n2358) );
  AND U2360 ( .A(n2376), .B(n2377), .Z(n2375) );
  XOR U2361 ( .A(n2374), .B(n2378), .Z(n2376) );
  XNOR U2362 ( .A(n2357), .B(n2349), .Z(n2373) );
  XOR U2363 ( .A(n2379), .B(n2380), .Z(n2349) );
  AND U2364 ( .A(n2381), .B(n2382), .Z(n2380) );
  XNOR U2365 ( .A(n2383), .B(n2379), .Z(n2381) );
  XNOR U2366 ( .A(n2384), .B(n2354), .Z(n2357) );
  XOR U2367 ( .A(n2385), .B(n2386), .Z(n2354) );
  AND U2368 ( .A(n2387), .B(n2388), .Z(n2386) );
  XOR U2369 ( .A(n2385), .B(n2389), .Z(n2387) );
  XNOR U2370 ( .A(n2390), .B(n2391), .Z(n2384) );
  AND U2371 ( .A(n2392), .B(n2393), .Z(n2391) );
  XNOR U2372 ( .A(n2390), .B(n2394), .Z(n2392) );
  XNOR U2373 ( .A(n2353), .B(n2360), .Z(n2372) );
  AND U2374 ( .A(n2315), .B(n2395), .Z(n2360) );
  XOR U2375 ( .A(n2365), .B(n2364), .Z(n2353) );
  XNOR U2376 ( .A(n2396), .B(n2361), .Z(n2364) );
  XOR U2377 ( .A(n2397), .B(n2398), .Z(n2361) );
  AND U2378 ( .A(n2399), .B(n2400), .Z(n2398) );
  XOR U2379 ( .A(n2397), .B(n2401), .Z(n2399) );
  XNOR U2380 ( .A(n2402), .B(n2403), .Z(n2396) );
  AND U2381 ( .A(n2404), .B(n2405), .Z(n2403) );
  XOR U2382 ( .A(n2402), .B(n2406), .Z(n2404) );
  XOR U2383 ( .A(n2407), .B(n2408), .Z(n2365) );
  AND U2384 ( .A(n2409), .B(n2410), .Z(n2408) );
  XOR U2385 ( .A(n2407), .B(n2411), .Z(n2409) );
  XNOR U2386 ( .A(n2300), .B(n2368), .Z(n2370) );
  XNOR U2387 ( .A(n2412), .B(n2413), .Z(n2300) );
  AND U2388 ( .A(n89), .B(n2307), .Z(n2413) );
  XOR U2389 ( .A(n2412), .B(n2305), .Z(n2307) );
  XOR U2390 ( .A(n2414), .B(n2415), .Z(n2368) );
  AND U2391 ( .A(n2416), .B(n2417), .Z(n2415) );
  XNOR U2392 ( .A(n2414), .B(n2315), .Z(n2417) );
  XOR U2393 ( .A(n2418), .B(n2382), .Z(n2315) );
  XNOR U2394 ( .A(n2419), .B(n2389), .Z(n2382) );
  XOR U2395 ( .A(n2378), .B(n2377), .Z(n2389) );
  XNOR U2396 ( .A(n2420), .B(n2374), .Z(n2377) );
  XOR U2397 ( .A(n2421), .B(n2422), .Z(n2374) );
  AND U2398 ( .A(n2423), .B(n2424), .Z(n2422) );
  XOR U2399 ( .A(n2421), .B(n2425), .Z(n2423) );
  XNOR U2400 ( .A(n2426), .B(n2427), .Z(n2420) );
  NOR U2401 ( .A(n2428), .B(n2429), .Z(n2427) );
  XNOR U2402 ( .A(n2426), .B(n2430), .Z(n2428) );
  XOR U2403 ( .A(n2431), .B(n2432), .Z(n2378) );
  NOR U2404 ( .A(n2433), .B(n2434), .Z(n2432) );
  XNOR U2405 ( .A(n2431), .B(n2435), .Z(n2433) );
  XNOR U2406 ( .A(n2388), .B(n2379), .Z(n2419) );
  XOR U2407 ( .A(n2436), .B(n2437), .Z(n2379) );
  NOR U2408 ( .A(n2438), .B(n2439), .Z(n2437) );
  XNOR U2409 ( .A(n2436), .B(n2440), .Z(n2438) );
  XOR U2410 ( .A(n2441), .B(n2394), .Z(n2388) );
  XNOR U2411 ( .A(n2442), .B(n2443), .Z(n2394) );
  NOR U2412 ( .A(n2444), .B(n2445), .Z(n2443) );
  XNOR U2413 ( .A(n2442), .B(n2446), .Z(n2444) );
  XNOR U2414 ( .A(n2393), .B(n2385), .Z(n2441) );
  XOR U2415 ( .A(n2447), .B(n2448), .Z(n2385) );
  AND U2416 ( .A(n2449), .B(n2450), .Z(n2448) );
  XOR U2417 ( .A(n2447), .B(n2451), .Z(n2449) );
  XNOR U2418 ( .A(n2452), .B(n2390), .Z(n2393) );
  XOR U2419 ( .A(n2453), .B(n2454), .Z(n2390) );
  AND U2420 ( .A(n2455), .B(n2456), .Z(n2454) );
  XOR U2421 ( .A(n2453), .B(n2457), .Z(n2455) );
  XNOR U2422 ( .A(n2458), .B(n2459), .Z(n2452) );
  NOR U2423 ( .A(n2460), .B(n2461), .Z(n2459) );
  XOR U2424 ( .A(n2458), .B(n2462), .Z(n2460) );
  XOR U2425 ( .A(n2383), .B(n2395), .Z(n2418) );
  NOR U2426 ( .A(n2323), .B(n2463), .Z(n2395) );
  XNOR U2427 ( .A(n2401), .B(n2400), .Z(n2383) );
  XNOR U2428 ( .A(n2464), .B(n2406), .Z(n2400) );
  XOR U2429 ( .A(n2465), .B(n2466), .Z(n2406) );
  NOR U2430 ( .A(n2467), .B(n2468), .Z(n2466) );
  XNOR U2431 ( .A(n2465), .B(n2469), .Z(n2467) );
  XNOR U2432 ( .A(n2405), .B(n2397), .Z(n2464) );
  XOR U2433 ( .A(n2470), .B(n2471), .Z(n2397) );
  AND U2434 ( .A(n2472), .B(n2473), .Z(n2471) );
  XNOR U2435 ( .A(n2470), .B(n2474), .Z(n2472) );
  XNOR U2436 ( .A(n2475), .B(n2402), .Z(n2405) );
  XOR U2437 ( .A(n2476), .B(n2477), .Z(n2402) );
  AND U2438 ( .A(n2478), .B(n2479), .Z(n2477) );
  XOR U2439 ( .A(n2476), .B(n2480), .Z(n2478) );
  XNOR U2440 ( .A(n2481), .B(n2482), .Z(n2475) );
  NOR U2441 ( .A(n2483), .B(n2484), .Z(n2482) );
  XOR U2442 ( .A(n2481), .B(n2485), .Z(n2483) );
  XOR U2443 ( .A(n2411), .B(n2410), .Z(n2401) );
  XNOR U2444 ( .A(n2486), .B(n2407), .Z(n2410) );
  XOR U2445 ( .A(n2487), .B(n2488), .Z(n2407) );
  AND U2446 ( .A(n2489), .B(n2490), .Z(n2488) );
  XOR U2447 ( .A(n2487), .B(n2491), .Z(n2489) );
  XNOR U2448 ( .A(n2492), .B(n2493), .Z(n2486) );
  NOR U2449 ( .A(n2494), .B(n2495), .Z(n2493) );
  XNOR U2450 ( .A(n2492), .B(n2496), .Z(n2494) );
  XOR U2451 ( .A(n2497), .B(n2498), .Z(n2411) );
  NOR U2452 ( .A(n2499), .B(n2500), .Z(n2498) );
  XNOR U2453 ( .A(n2497), .B(n2501), .Z(n2499) );
  XNOR U2454 ( .A(n2312), .B(n2414), .Z(n2416) );
  XNOR U2455 ( .A(n2502), .B(n2503), .Z(n2312) );
  AND U2456 ( .A(n89), .B(n2319), .Z(n2503) );
  XOR U2457 ( .A(n2502), .B(n2317), .Z(n2319) );
  AND U2458 ( .A(n2320), .B(n2323), .Z(n2414) );
  XOR U2459 ( .A(n2504), .B(n2463), .Z(n2323) );
  XNOR U2460 ( .A(p_input[256]), .B(p_input[64]), .Z(n2463) );
  XOR U2461 ( .A(n2440), .B(n2439), .Z(n2504) );
  XOR U2462 ( .A(n2505), .B(n2451), .Z(n2439) );
  XOR U2463 ( .A(n2425), .B(n2424), .Z(n2451) );
  XNOR U2464 ( .A(n2506), .B(n2430), .Z(n2424) );
  XOR U2465 ( .A(p_input[280]), .B(p_input[88]), .Z(n2430) );
  XOR U2466 ( .A(n2421), .B(n2429), .Z(n2506) );
  XOR U2467 ( .A(n2507), .B(n2426), .Z(n2429) );
  XOR U2468 ( .A(p_input[278]), .B(p_input[86]), .Z(n2426) );
  XNOR U2469 ( .A(p_input[279]), .B(p_input[87]), .Z(n2507) );
  XNOR U2470 ( .A(n2225), .B(p_input[82]), .Z(n2421) );
  XNOR U2471 ( .A(n2435), .B(n2434), .Z(n2425) );
  XOR U2472 ( .A(n2508), .B(n2431), .Z(n2434) );
  XOR U2473 ( .A(p_input[275]), .B(p_input[83]), .Z(n2431) );
  XNOR U2474 ( .A(p_input[276]), .B(p_input[84]), .Z(n2508) );
  XOR U2475 ( .A(p_input[277]), .B(p_input[85]), .Z(n2435) );
  XNOR U2476 ( .A(n2450), .B(n2436), .Z(n2505) );
  XNOR U2477 ( .A(n2227), .B(p_input[65]), .Z(n2436) );
  XNOR U2478 ( .A(n2509), .B(n2457), .Z(n2450) );
  XNOR U2479 ( .A(n2446), .B(n2445), .Z(n2457) );
  XOR U2480 ( .A(n2510), .B(n2442), .Z(n2445) );
  XNOR U2481 ( .A(n2230), .B(p_input[90]), .Z(n2442) );
  XNOR U2482 ( .A(p_input[283]), .B(p_input[91]), .Z(n2510) );
  XOR U2483 ( .A(p_input[284]), .B(p_input[92]), .Z(n2446) );
  XNOR U2484 ( .A(n2456), .B(n2447), .Z(n2509) );
  XNOR U2485 ( .A(n2231), .B(p_input[81]), .Z(n2447) );
  XOR U2486 ( .A(n2511), .B(n2462), .Z(n2456) );
  XNOR U2487 ( .A(p_input[287]), .B(p_input[95]), .Z(n2462) );
  XOR U2488 ( .A(n2453), .B(n2461), .Z(n2511) );
  XOR U2489 ( .A(n2512), .B(n2458), .Z(n2461) );
  XOR U2490 ( .A(p_input[285]), .B(p_input[93]), .Z(n2458) );
  XNOR U2491 ( .A(p_input[286]), .B(p_input[94]), .Z(n2512) );
  XNOR U2492 ( .A(n2234), .B(p_input[89]), .Z(n2453) );
  XNOR U2493 ( .A(n2474), .B(n2473), .Z(n2440) );
  XNOR U2494 ( .A(n2513), .B(n2480), .Z(n2473) );
  XNOR U2495 ( .A(n2469), .B(n2468), .Z(n2480) );
  XOR U2496 ( .A(n2514), .B(n2465), .Z(n2468) );
  XNOR U2497 ( .A(n2237), .B(p_input[75]), .Z(n2465) );
  XNOR U2498 ( .A(p_input[268]), .B(p_input[76]), .Z(n2514) );
  XOR U2499 ( .A(p_input[269]), .B(p_input[77]), .Z(n2469) );
  XNOR U2500 ( .A(n2479), .B(n2470), .Z(n2513) );
  XOR U2501 ( .A(p_input[258]), .B(p_input[66]), .Z(n2470) );
  XOR U2502 ( .A(n2515), .B(n2485), .Z(n2479) );
  XNOR U2503 ( .A(p_input[272]), .B(p_input[80]), .Z(n2485) );
  XOR U2504 ( .A(n2476), .B(n2484), .Z(n2515) );
  XOR U2505 ( .A(n2516), .B(n2481), .Z(n2484) );
  XOR U2506 ( .A(p_input[270]), .B(p_input[78]), .Z(n2481) );
  XNOR U2507 ( .A(p_input[271]), .B(p_input[79]), .Z(n2516) );
  XNOR U2508 ( .A(n2240), .B(p_input[74]), .Z(n2476) );
  XNOR U2509 ( .A(n2491), .B(n2490), .Z(n2474) );
  XNOR U2510 ( .A(n2517), .B(n2496), .Z(n2490) );
  XOR U2511 ( .A(p_input[265]), .B(p_input[73]), .Z(n2496) );
  XOR U2512 ( .A(n2487), .B(n2495), .Z(n2517) );
  XOR U2513 ( .A(n2518), .B(n2492), .Z(n2495) );
  XOR U2514 ( .A(p_input[263]), .B(p_input[71]), .Z(n2492) );
  XNOR U2515 ( .A(p_input[264]), .B(p_input[72]), .Z(n2518) );
  XOR U2516 ( .A(p_input[259]), .B(p_input[67]), .Z(n2487) );
  XNOR U2517 ( .A(n2501), .B(n2500), .Z(n2491) );
  XOR U2518 ( .A(n2519), .B(n2497), .Z(n2500) );
  XOR U2519 ( .A(p_input[260]), .B(p_input[68]), .Z(n2497) );
  XNOR U2520 ( .A(p_input[261]), .B(p_input[69]), .Z(n2519) );
  XOR U2521 ( .A(p_input[262]), .B(p_input[70]), .Z(n2501) );
  XNOR U2522 ( .A(n2520), .B(n2521), .Z(n2320) );
  AND U2523 ( .A(n89), .B(n2522), .Z(n2521) );
  XNOR U2524 ( .A(n2523), .B(n2524), .Z(n89) );
  NOR U2525 ( .A(n2525), .B(n2526), .Z(n2524) );
  XOR U2526 ( .A(n2274), .B(n2523), .Z(n2526) );
  NOR U2527 ( .A(n2523), .B(n2273), .Z(n2525) );
  XOR U2528 ( .A(n2527), .B(n2528), .Z(n2523) );
  AND U2529 ( .A(n2529), .B(n2530), .Z(n2528) );
  XNOR U2530 ( .A(n2341), .B(n2527), .Z(n2530) );
  XOR U2531 ( .A(n2527), .B(n2284), .Z(n2529) );
  XOR U2532 ( .A(n2531), .B(n2532), .Z(n2527) );
  AND U2533 ( .A(n2533), .B(n2534), .Z(n2532) );
  XNOR U2534 ( .A(n2366), .B(n2531), .Z(n2534) );
  XOR U2535 ( .A(n2531), .B(n2295), .Z(n2533) );
  XOR U2536 ( .A(n2535), .B(n2536), .Z(n2531) );
  AND U2537 ( .A(n2537), .B(n2538), .Z(n2536) );
  XOR U2538 ( .A(n2535), .B(n2305), .Z(n2537) );
  XOR U2539 ( .A(n2539), .B(n2540), .Z(n2263) );
  AND U2540 ( .A(n93), .B(n2522), .Z(n2540) );
  XNOR U2541 ( .A(n2520), .B(n2539), .Z(n2522) );
  XNOR U2542 ( .A(n2541), .B(n2542), .Z(n93) );
  NOR U2543 ( .A(n2543), .B(n2544), .Z(n2542) );
  XNOR U2544 ( .A(n2274), .B(n2545), .Z(n2544) );
  IV U2545 ( .A(n2541), .Z(n2545) );
  AND U2546 ( .A(n2546), .B(n2547), .Z(n2274) );
  NOR U2547 ( .A(n2541), .B(n2273), .Z(n2543) );
  AND U2548 ( .A(n2548), .B(n2549), .Z(n2273) );
  IV U2549 ( .A(n2550), .Z(n2548) );
  XOR U2550 ( .A(n2551), .B(n2552), .Z(n2541) );
  AND U2551 ( .A(n2553), .B(n2554), .Z(n2552) );
  XNOR U2552 ( .A(n2551), .B(n2341), .Z(n2554) );
  XNOR U2553 ( .A(n2555), .B(n2556), .Z(n2341) );
  AND U2554 ( .A(n96), .B(n2557), .Z(n2556) );
  XOR U2555 ( .A(n2558), .B(n2555), .Z(n2557) );
  XNOR U2556 ( .A(n2559), .B(n2551), .Z(n2553) );
  IV U2557 ( .A(n2284), .Z(n2559) );
  XOR U2558 ( .A(n2560), .B(n2561), .Z(n2284) );
  AND U2559 ( .A(n104), .B(n2562), .Z(n2561) );
  XOR U2560 ( .A(n2563), .B(n2564), .Z(n2551) );
  AND U2561 ( .A(n2565), .B(n2566), .Z(n2564) );
  XNOR U2562 ( .A(n2563), .B(n2366), .Z(n2566) );
  XNOR U2563 ( .A(n2567), .B(n2568), .Z(n2366) );
  AND U2564 ( .A(n96), .B(n2569), .Z(n2568) );
  XNOR U2565 ( .A(n2570), .B(n2567), .Z(n2569) );
  XOR U2566 ( .A(n2295), .B(n2563), .Z(n2565) );
  XOR U2567 ( .A(n2571), .B(n2572), .Z(n2295) );
  AND U2568 ( .A(n104), .B(n2573), .Z(n2572) );
  XOR U2569 ( .A(n2535), .B(n2574), .Z(n2563) );
  AND U2570 ( .A(n2575), .B(n2538), .Z(n2574) );
  XNOR U2571 ( .A(n2412), .B(n2535), .Z(n2538) );
  XNOR U2572 ( .A(n2576), .B(n2577), .Z(n2412) );
  AND U2573 ( .A(n96), .B(n2578), .Z(n2577) );
  XOR U2574 ( .A(n2579), .B(n2576), .Z(n2578) );
  XNOR U2575 ( .A(n2580), .B(n2535), .Z(n2575) );
  IV U2576 ( .A(n2305), .Z(n2580) );
  XOR U2577 ( .A(n2581), .B(n2582), .Z(n2305) );
  AND U2578 ( .A(n104), .B(n2583), .Z(n2582) );
  XOR U2579 ( .A(n2584), .B(n2585), .Z(n2535) );
  AND U2580 ( .A(n2586), .B(n2587), .Z(n2585) );
  XNOR U2581 ( .A(n2584), .B(n2502), .Z(n2587) );
  XNOR U2582 ( .A(n2588), .B(n2589), .Z(n2502) );
  AND U2583 ( .A(n96), .B(n2590), .Z(n2589) );
  XNOR U2584 ( .A(n2591), .B(n2588), .Z(n2590) );
  XNOR U2585 ( .A(n2592), .B(n2584), .Z(n2586) );
  IV U2586 ( .A(n2317), .Z(n2592) );
  XOR U2587 ( .A(n2593), .B(n2594), .Z(n2317) );
  AND U2588 ( .A(n104), .B(n2595), .Z(n2594) );
  AND U2589 ( .A(n2539), .B(n2520), .Z(n2584) );
  XNOR U2590 ( .A(n2596), .B(n2597), .Z(n2520) );
  AND U2591 ( .A(n96), .B(n2598), .Z(n2597) );
  XNOR U2592 ( .A(n2599), .B(n2596), .Z(n2598) );
  XNOR U2593 ( .A(n2600), .B(n2601), .Z(n96) );
  NOR U2594 ( .A(n2602), .B(n2603), .Z(n2601) );
  XNOR U2595 ( .A(n2600), .B(n2550), .Z(n2603) );
  NOR U2596 ( .A(n2546), .B(n2547), .Z(n2550) );
  NOR U2597 ( .A(n2600), .B(n2549), .Z(n2602) );
  AND U2598 ( .A(n2604), .B(n2605), .Z(n2549) );
  XOR U2599 ( .A(n2606), .B(n2607), .Z(n2600) );
  AND U2600 ( .A(n2608), .B(n2609), .Z(n2607) );
  XNOR U2601 ( .A(n2606), .B(n2604), .Z(n2609) );
  IV U2602 ( .A(n2558), .Z(n2604) );
  XOR U2603 ( .A(n2610), .B(n2611), .Z(n2558) );
  XOR U2604 ( .A(n2612), .B(n2605), .Z(n2611) );
  AND U2605 ( .A(n2570), .B(n2613), .Z(n2605) );
  AND U2606 ( .A(n2614), .B(n2615), .Z(n2612) );
  XOR U2607 ( .A(n2616), .B(n2610), .Z(n2614) );
  XNOR U2608 ( .A(n2555), .B(n2606), .Z(n2608) );
  XNOR U2609 ( .A(n2617), .B(n2618), .Z(n2555) );
  AND U2610 ( .A(n100), .B(n2562), .Z(n2618) );
  XOR U2611 ( .A(n2617), .B(n2560), .Z(n2562) );
  XOR U2612 ( .A(n2619), .B(n2620), .Z(n2606) );
  AND U2613 ( .A(n2621), .B(n2622), .Z(n2620) );
  XNOR U2614 ( .A(n2619), .B(n2570), .Z(n2622) );
  XOR U2615 ( .A(n2623), .B(n2615), .Z(n2570) );
  XNOR U2616 ( .A(n2624), .B(n2610), .Z(n2615) );
  XOR U2617 ( .A(n2625), .B(n2626), .Z(n2610) );
  AND U2618 ( .A(n2627), .B(n2628), .Z(n2626) );
  XOR U2619 ( .A(n2629), .B(n2625), .Z(n2627) );
  XNOR U2620 ( .A(n2630), .B(n2631), .Z(n2624) );
  AND U2621 ( .A(n2632), .B(n2633), .Z(n2631) );
  XOR U2622 ( .A(n2630), .B(n2634), .Z(n2632) );
  XNOR U2623 ( .A(n2616), .B(n2613), .Z(n2623) );
  AND U2624 ( .A(n2635), .B(n2636), .Z(n2613) );
  XOR U2625 ( .A(n2637), .B(n2638), .Z(n2616) );
  AND U2626 ( .A(n2639), .B(n2640), .Z(n2638) );
  XOR U2627 ( .A(n2637), .B(n2641), .Z(n2639) );
  XNOR U2628 ( .A(n2567), .B(n2619), .Z(n2621) );
  XNOR U2629 ( .A(n2642), .B(n2643), .Z(n2567) );
  AND U2630 ( .A(n100), .B(n2573), .Z(n2643) );
  XOR U2631 ( .A(n2642), .B(n2571), .Z(n2573) );
  XOR U2632 ( .A(n2644), .B(n2645), .Z(n2619) );
  AND U2633 ( .A(n2646), .B(n2647), .Z(n2645) );
  XNOR U2634 ( .A(n2644), .B(n2635), .Z(n2647) );
  IV U2635 ( .A(n2579), .Z(n2635) );
  XNOR U2636 ( .A(n2648), .B(n2628), .Z(n2579) );
  XNOR U2637 ( .A(n2649), .B(n2634), .Z(n2628) );
  XOR U2638 ( .A(n2650), .B(n2651), .Z(n2634) );
  AND U2639 ( .A(n2652), .B(n2653), .Z(n2651) );
  XOR U2640 ( .A(n2650), .B(n2654), .Z(n2652) );
  XNOR U2641 ( .A(n2633), .B(n2625), .Z(n2649) );
  XOR U2642 ( .A(n2655), .B(n2656), .Z(n2625) );
  AND U2643 ( .A(n2657), .B(n2658), .Z(n2656) );
  XNOR U2644 ( .A(n2659), .B(n2655), .Z(n2657) );
  XNOR U2645 ( .A(n2660), .B(n2630), .Z(n2633) );
  XOR U2646 ( .A(n2661), .B(n2662), .Z(n2630) );
  AND U2647 ( .A(n2663), .B(n2664), .Z(n2662) );
  XOR U2648 ( .A(n2661), .B(n2665), .Z(n2663) );
  XNOR U2649 ( .A(n2666), .B(n2667), .Z(n2660) );
  AND U2650 ( .A(n2668), .B(n2669), .Z(n2667) );
  XNOR U2651 ( .A(n2666), .B(n2670), .Z(n2668) );
  XNOR U2652 ( .A(n2629), .B(n2636), .Z(n2648) );
  AND U2653 ( .A(n2591), .B(n2671), .Z(n2636) );
  XOR U2654 ( .A(n2641), .B(n2640), .Z(n2629) );
  XNOR U2655 ( .A(n2672), .B(n2637), .Z(n2640) );
  XOR U2656 ( .A(n2673), .B(n2674), .Z(n2637) );
  AND U2657 ( .A(n2675), .B(n2676), .Z(n2674) );
  XOR U2658 ( .A(n2673), .B(n2677), .Z(n2675) );
  XNOR U2659 ( .A(n2678), .B(n2679), .Z(n2672) );
  AND U2660 ( .A(n2680), .B(n2681), .Z(n2679) );
  XOR U2661 ( .A(n2678), .B(n2682), .Z(n2680) );
  XOR U2662 ( .A(n2683), .B(n2684), .Z(n2641) );
  AND U2663 ( .A(n2685), .B(n2686), .Z(n2684) );
  XOR U2664 ( .A(n2683), .B(n2687), .Z(n2685) );
  XNOR U2665 ( .A(n2576), .B(n2644), .Z(n2646) );
  XNOR U2666 ( .A(n2688), .B(n2689), .Z(n2576) );
  AND U2667 ( .A(n100), .B(n2583), .Z(n2689) );
  XOR U2668 ( .A(n2688), .B(n2581), .Z(n2583) );
  XOR U2669 ( .A(n2690), .B(n2691), .Z(n2644) );
  AND U2670 ( .A(n2692), .B(n2693), .Z(n2691) );
  XNOR U2671 ( .A(n2690), .B(n2591), .Z(n2693) );
  XOR U2672 ( .A(n2694), .B(n2658), .Z(n2591) );
  XNOR U2673 ( .A(n2695), .B(n2665), .Z(n2658) );
  XOR U2674 ( .A(n2654), .B(n2653), .Z(n2665) );
  XNOR U2675 ( .A(n2696), .B(n2650), .Z(n2653) );
  XOR U2676 ( .A(n2697), .B(n2698), .Z(n2650) );
  AND U2677 ( .A(n2699), .B(n2700), .Z(n2698) );
  XNOR U2678 ( .A(n2701), .B(n2702), .Z(n2699) );
  IV U2679 ( .A(n2697), .Z(n2701) );
  XNOR U2680 ( .A(n2703), .B(n2704), .Z(n2696) );
  NOR U2681 ( .A(n2705), .B(n2706), .Z(n2704) );
  XNOR U2682 ( .A(n2703), .B(n2707), .Z(n2705) );
  XOR U2683 ( .A(n2708), .B(n2709), .Z(n2654) );
  NOR U2684 ( .A(n2710), .B(n2711), .Z(n2709) );
  XNOR U2685 ( .A(n2708), .B(n2712), .Z(n2710) );
  XNOR U2686 ( .A(n2664), .B(n2655), .Z(n2695) );
  XOR U2687 ( .A(n2713), .B(n2714), .Z(n2655) );
  AND U2688 ( .A(n2715), .B(n2716), .Z(n2714) );
  XOR U2689 ( .A(n2713), .B(n2717), .Z(n2715) );
  XOR U2690 ( .A(n2718), .B(n2670), .Z(n2664) );
  XOR U2691 ( .A(n2719), .B(n2720), .Z(n2670) );
  NOR U2692 ( .A(n2721), .B(n2722), .Z(n2720) );
  XOR U2693 ( .A(n2719), .B(n2723), .Z(n2721) );
  XNOR U2694 ( .A(n2669), .B(n2661), .Z(n2718) );
  XOR U2695 ( .A(n2724), .B(n2725), .Z(n2661) );
  AND U2696 ( .A(n2726), .B(n2727), .Z(n2725) );
  XOR U2697 ( .A(n2724), .B(n2728), .Z(n2726) );
  XNOR U2698 ( .A(n2729), .B(n2666), .Z(n2669) );
  XNOR U2699 ( .A(n2730), .B(n2731), .Z(n2666) );
  NOR U2700 ( .A(n2732), .B(n2733), .Z(n2731) );
  XOR U2701 ( .A(n2730), .B(n2734), .Z(n2732) );
  XNOR U2702 ( .A(n2735), .B(n2736), .Z(n2729) );
  NOR U2703 ( .A(n2737), .B(n2738), .Z(n2736) );
  XNOR U2704 ( .A(n2735), .B(n2739), .Z(n2737) );
  XOR U2705 ( .A(n2659), .B(n2671), .Z(n2694) );
  NOR U2706 ( .A(n2599), .B(n2740), .Z(n2671) );
  XNOR U2707 ( .A(n2677), .B(n2676), .Z(n2659) );
  XNOR U2708 ( .A(n2741), .B(n2682), .Z(n2676) );
  XNOR U2709 ( .A(n2742), .B(n2743), .Z(n2682) );
  NOR U2710 ( .A(n2744), .B(n2745), .Z(n2743) );
  XOR U2711 ( .A(n2742), .B(n2746), .Z(n2744) );
  XNOR U2712 ( .A(n2681), .B(n2673), .Z(n2741) );
  XOR U2713 ( .A(n2747), .B(n2748), .Z(n2673) );
  AND U2714 ( .A(n2749), .B(n2750), .Z(n2748) );
  XOR U2715 ( .A(n2747), .B(n2751), .Z(n2749) );
  XNOR U2716 ( .A(n2752), .B(n2678), .Z(n2681) );
  XOR U2717 ( .A(n2753), .B(n2754), .Z(n2678) );
  AND U2718 ( .A(n2755), .B(n2756), .Z(n2754) );
  XNOR U2719 ( .A(n2757), .B(n2758), .Z(n2755) );
  IV U2720 ( .A(n2753), .Z(n2757) );
  XNOR U2721 ( .A(n2759), .B(n2760), .Z(n2752) );
  NOR U2722 ( .A(n2761), .B(n2762), .Z(n2760) );
  XNOR U2723 ( .A(n2759), .B(n2763), .Z(n2761) );
  XOR U2724 ( .A(n2687), .B(n2686), .Z(n2677) );
  XNOR U2725 ( .A(n2764), .B(n2683), .Z(n2686) );
  XOR U2726 ( .A(n2765), .B(n2766), .Z(n2683) );
  NOR U2727 ( .A(n2767), .B(n2768), .Z(n2766) );
  XNOR U2728 ( .A(n2765), .B(n2769), .Z(n2767) );
  XNOR U2729 ( .A(n2770), .B(n2771), .Z(n2764) );
  NOR U2730 ( .A(n2772), .B(n2773), .Z(n2771) );
  XNOR U2731 ( .A(n2770), .B(n2774), .Z(n2772) );
  XOR U2732 ( .A(n2775), .B(n2776), .Z(n2687) );
  NOR U2733 ( .A(n2777), .B(n2778), .Z(n2776) );
  XNOR U2734 ( .A(n2775), .B(n2779), .Z(n2777) );
  XNOR U2735 ( .A(n2588), .B(n2690), .Z(n2692) );
  XNOR U2736 ( .A(n2780), .B(n2781), .Z(n2588) );
  AND U2737 ( .A(n100), .B(n2595), .Z(n2781) );
  XOR U2738 ( .A(n2780), .B(n2593), .Z(n2595) );
  AND U2739 ( .A(n2596), .B(n2599), .Z(n2690) );
  XOR U2740 ( .A(n2782), .B(n2740), .Z(n2599) );
  XNOR U2741 ( .A(p_input[256]), .B(p_input[96]), .Z(n2740) );
  XNOR U2742 ( .A(n2717), .B(n2716), .Z(n2782) );
  XNOR U2743 ( .A(n2783), .B(n2728), .Z(n2716) );
  XOR U2744 ( .A(n2702), .B(n2700), .Z(n2728) );
  XNOR U2745 ( .A(n2784), .B(n2707), .Z(n2700) );
  XOR U2746 ( .A(p_input[120]), .B(p_input[280]), .Z(n2707) );
  XOR U2747 ( .A(n2697), .B(n2706), .Z(n2784) );
  XOR U2748 ( .A(n2785), .B(n2703), .Z(n2706) );
  XOR U2749 ( .A(p_input[118]), .B(p_input[278]), .Z(n2703) );
  XOR U2750 ( .A(p_input[119]), .B(n1937), .Z(n2785) );
  XOR U2751 ( .A(p_input[114]), .B(p_input[274]), .Z(n2697) );
  XNOR U2752 ( .A(n2712), .B(n2711), .Z(n2702) );
  XOR U2753 ( .A(n2786), .B(n2708), .Z(n2711) );
  XOR U2754 ( .A(p_input[115]), .B(p_input[275]), .Z(n2708) );
  XOR U2755 ( .A(p_input[116]), .B(n1939), .Z(n2786) );
  XOR U2756 ( .A(p_input[117]), .B(p_input[277]), .Z(n2712) );
  XNOR U2757 ( .A(n2727), .B(n2713), .Z(n2783) );
  XNOR U2758 ( .A(n2227), .B(p_input[97]), .Z(n2713) );
  XNOR U2759 ( .A(n2787), .B(n2734), .Z(n2727) );
  XNOR U2760 ( .A(n2723), .B(n2722), .Z(n2734) );
  XNOR U2761 ( .A(n2788), .B(n2719), .Z(n2722) );
  XNOR U2762 ( .A(p_input[122]), .B(p_input[282]), .Z(n2719) );
  XOR U2763 ( .A(p_input[123]), .B(n1943), .Z(n2788) );
  XOR U2764 ( .A(p_input[124]), .B(p_input[284]), .Z(n2723) );
  XNOR U2765 ( .A(n2733), .B(n2789), .Z(n2787) );
  IV U2766 ( .A(n2724), .Z(n2789) );
  XOR U2767 ( .A(p_input[113]), .B(p_input[273]), .Z(n2724) );
  XOR U2768 ( .A(n2790), .B(n2739), .Z(n2733) );
  XOR U2769 ( .A(p_input[127]), .B(p_input[287]), .Z(n2739) );
  XNOR U2770 ( .A(n2730), .B(n2738), .Z(n2790) );
  XOR U2771 ( .A(n2791), .B(n2735), .Z(n2738) );
  XOR U2772 ( .A(p_input[125]), .B(p_input[285]), .Z(n2735) );
  XNOR U2773 ( .A(p_input[126]), .B(p_input[286]), .Z(n2791) );
  XNOR U2774 ( .A(p_input[121]), .B(p_input[281]), .Z(n2730) );
  XOR U2775 ( .A(n2751), .B(n2750), .Z(n2717) );
  XNOR U2776 ( .A(n2792), .B(n2758), .Z(n2750) );
  XNOR U2777 ( .A(n2746), .B(n2745), .Z(n2758) );
  XNOR U2778 ( .A(n2793), .B(n2742), .Z(n2745) );
  XNOR U2779 ( .A(p_input[107]), .B(p_input[267]), .Z(n2742) );
  XOR U2780 ( .A(p_input[108]), .B(n1949), .Z(n2793) );
  XOR U2781 ( .A(p_input[109]), .B(p_input[269]), .Z(n2746) );
  XNOR U2782 ( .A(n2756), .B(n2747), .Z(n2792) );
  XOR U2783 ( .A(p_input[258]), .B(p_input[98]), .Z(n2747) );
  XNOR U2784 ( .A(n2794), .B(n2763), .Z(n2756) );
  XNOR U2785 ( .A(p_input[112]), .B(n1951), .Z(n2763) );
  XOR U2786 ( .A(n2753), .B(n2762), .Z(n2794) );
  XOR U2787 ( .A(n2795), .B(n2759), .Z(n2762) );
  XOR U2788 ( .A(p_input[110]), .B(p_input[270]), .Z(n2759) );
  XOR U2789 ( .A(p_input[111]), .B(n1953), .Z(n2795) );
  XOR U2790 ( .A(p_input[106]), .B(p_input[266]), .Z(n2753) );
  XNOR U2791 ( .A(n2769), .B(n2768), .Z(n2751) );
  XOR U2792 ( .A(n2796), .B(n2774), .Z(n2768) );
  XOR U2793 ( .A(p_input[105]), .B(p_input[265]), .Z(n2774) );
  XOR U2794 ( .A(n2765), .B(n2773), .Z(n2796) );
  XOR U2795 ( .A(n2797), .B(n2770), .Z(n2773) );
  XOR U2796 ( .A(p_input[103]), .B(p_input[263]), .Z(n2770) );
  XNOR U2797 ( .A(p_input[104]), .B(p_input[264]), .Z(n2797) );
  XOR U2798 ( .A(p_input[259]), .B(p_input[99]), .Z(n2765) );
  XNOR U2799 ( .A(n2779), .B(n2778), .Z(n2769) );
  XOR U2800 ( .A(n2798), .B(n2775), .Z(n2778) );
  XOR U2801 ( .A(p_input[100]), .B(p_input[260]), .Z(n2775) );
  XNOR U2802 ( .A(p_input[101]), .B(p_input[261]), .Z(n2798) );
  XOR U2803 ( .A(p_input[102]), .B(p_input[262]), .Z(n2779) );
  XNOR U2804 ( .A(n2799), .B(n2800), .Z(n2596) );
  AND U2805 ( .A(n100), .B(n2801), .Z(n2800) );
  XNOR U2806 ( .A(n2802), .B(n2803), .Z(n100) );
  NOR U2807 ( .A(n2804), .B(n2805), .Z(n2803) );
  XOR U2808 ( .A(n2547), .B(n2802), .Z(n2805) );
  NOR U2809 ( .A(n2802), .B(n2546), .Z(n2804) );
  XOR U2810 ( .A(n2806), .B(n2807), .Z(n2802) );
  AND U2811 ( .A(n2808), .B(n2809), .Z(n2807) );
  XNOR U2812 ( .A(n2617), .B(n2806), .Z(n2809) );
  XOR U2813 ( .A(n2806), .B(n2560), .Z(n2808) );
  XOR U2814 ( .A(n2810), .B(n2811), .Z(n2806) );
  AND U2815 ( .A(n2812), .B(n2813), .Z(n2811) );
  XNOR U2816 ( .A(n2642), .B(n2810), .Z(n2813) );
  XOR U2817 ( .A(n2810), .B(n2571), .Z(n2812) );
  XOR U2818 ( .A(n2814), .B(n2815), .Z(n2810) );
  AND U2819 ( .A(n2816), .B(n2817), .Z(n2815) );
  XOR U2820 ( .A(n2814), .B(n2581), .Z(n2816) );
  XOR U2821 ( .A(n2818), .B(n2819), .Z(n2539) );
  AND U2822 ( .A(n104), .B(n2801), .Z(n2819) );
  XNOR U2823 ( .A(n2799), .B(n2818), .Z(n2801) );
  XNOR U2824 ( .A(n2820), .B(n2821), .Z(n104) );
  NOR U2825 ( .A(n2822), .B(n2823), .Z(n2821) );
  XNOR U2826 ( .A(n2547), .B(n2824), .Z(n2823) );
  IV U2827 ( .A(n2820), .Z(n2824) );
  AND U2828 ( .A(n2825), .B(n2826), .Z(n2547) );
  NOR U2829 ( .A(n2820), .B(n2546), .Z(n2822) );
  AND U2830 ( .A(n2827), .B(n2828), .Z(n2546) );
  IV U2831 ( .A(n2829), .Z(n2827) );
  XOR U2832 ( .A(n2830), .B(n2831), .Z(n2820) );
  AND U2833 ( .A(n2832), .B(n2833), .Z(n2831) );
  XNOR U2834 ( .A(n2830), .B(n2617), .Z(n2833) );
  XNOR U2835 ( .A(n2834), .B(n2835), .Z(n2617) );
  AND U2836 ( .A(n107), .B(n2836), .Z(n2835) );
  XOR U2837 ( .A(n2837), .B(n2834), .Z(n2836) );
  XNOR U2838 ( .A(n2838), .B(n2830), .Z(n2832) );
  IV U2839 ( .A(n2560), .Z(n2838) );
  XOR U2840 ( .A(n2839), .B(n2840), .Z(n2560) );
  AND U2841 ( .A(n115), .B(n2841), .Z(n2840) );
  XOR U2842 ( .A(n2842), .B(n2843), .Z(n2830) );
  AND U2843 ( .A(n2844), .B(n2845), .Z(n2843) );
  XNOR U2844 ( .A(n2842), .B(n2642), .Z(n2845) );
  XNOR U2845 ( .A(n2846), .B(n2847), .Z(n2642) );
  AND U2846 ( .A(n107), .B(n2848), .Z(n2847) );
  XNOR U2847 ( .A(n2849), .B(n2846), .Z(n2848) );
  XOR U2848 ( .A(n2571), .B(n2842), .Z(n2844) );
  XOR U2849 ( .A(n2850), .B(n2851), .Z(n2571) );
  AND U2850 ( .A(n115), .B(n2852), .Z(n2851) );
  XOR U2851 ( .A(n2814), .B(n2853), .Z(n2842) );
  AND U2852 ( .A(n2854), .B(n2817), .Z(n2853) );
  XNOR U2853 ( .A(n2688), .B(n2814), .Z(n2817) );
  XNOR U2854 ( .A(n2855), .B(n2856), .Z(n2688) );
  AND U2855 ( .A(n107), .B(n2857), .Z(n2856) );
  XOR U2856 ( .A(n2858), .B(n2855), .Z(n2857) );
  XNOR U2857 ( .A(n2859), .B(n2814), .Z(n2854) );
  IV U2858 ( .A(n2581), .Z(n2859) );
  XOR U2859 ( .A(n2860), .B(n2861), .Z(n2581) );
  AND U2860 ( .A(n115), .B(n2862), .Z(n2861) );
  XOR U2861 ( .A(n2863), .B(n2864), .Z(n2814) );
  AND U2862 ( .A(n2865), .B(n2866), .Z(n2864) );
  XNOR U2863 ( .A(n2863), .B(n2780), .Z(n2866) );
  XNOR U2864 ( .A(n2867), .B(n2868), .Z(n2780) );
  AND U2865 ( .A(n107), .B(n2869), .Z(n2868) );
  XNOR U2866 ( .A(n2870), .B(n2867), .Z(n2869) );
  XNOR U2867 ( .A(n2871), .B(n2863), .Z(n2865) );
  IV U2868 ( .A(n2593), .Z(n2871) );
  XOR U2869 ( .A(n2872), .B(n2873), .Z(n2593) );
  AND U2870 ( .A(n115), .B(n2874), .Z(n2873) );
  AND U2871 ( .A(n2818), .B(n2799), .Z(n2863) );
  XNOR U2872 ( .A(n2875), .B(n2876), .Z(n2799) );
  AND U2873 ( .A(n107), .B(n2877), .Z(n2876) );
  XNOR U2874 ( .A(n2878), .B(n2875), .Z(n2877) );
  XNOR U2875 ( .A(n2879), .B(n2880), .Z(n107) );
  NOR U2876 ( .A(n2881), .B(n2882), .Z(n2880) );
  XNOR U2877 ( .A(n2879), .B(n2829), .Z(n2882) );
  NOR U2878 ( .A(n2825), .B(n2826), .Z(n2829) );
  NOR U2879 ( .A(n2879), .B(n2828), .Z(n2881) );
  AND U2880 ( .A(n2883), .B(n2884), .Z(n2828) );
  XOR U2881 ( .A(n2885), .B(n2886), .Z(n2879) );
  AND U2882 ( .A(n2887), .B(n2888), .Z(n2886) );
  XNOR U2883 ( .A(n2885), .B(n2883), .Z(n2888) );
  IV U2884 ( .A(n2837), .Z(n2883) );
  XOR U2885 ( .A(n2889), .B(n2890), .Z(n2837) );
  XOR U2886 ( .A(n2891), .B(n2884), .Z(n2890) );
  AND U2887 ( .A(n2849), .B(n2892), .Z(n2884) );
  AND U2888 ( .A(n2893), .B(n2894), .Z(n2891) );
  XOR U2889 ( .A(n2895), .B(n2889), .Z(n2893) );
  XNOR U2890 ( .A(n2834), .B(n2885), .Z(n2887) );
  XNOR U2891 ( .A(n2896), .B(n2897), .Z(n2834) );
  AND U2892 ( .A(n111), .B(n2841), .Z(n2897) );
  XOR U2893 ( .A(n2896), .B(n2839), .Z(n2841) );
  XOR U2894 ( .A(n2898), .B(n2899), .Z(n2885) );
  AND U2895 ( .A(n2900), .B(n2901), .Z(n2899) );
  XNOR U2896 ( .A(n2898), .B(n2849), .Z(n2901) );
  XOR U2897 ( .A(n2902), .B(n2894), .Z(n2849) );
  XNOR U2898 ( .A(n2903), .B(n2889), .Z(n2894) );
  XOR U2899 ( .A(n2904), .B(n2905), .Z(n2889) );
  AND U2900 ( .A(n2906), .B(n2907), .Z(n2905) );
  XOR U2901 ( .A(n2908), .B(n2904), .Z(n2906) );
  XNOR U2902 ( .A(n2909), .B(n2910), .Z(n2903) );
  AND U2903 ( .A(n2911), .B(n2912), .Z(n2910) );
  XOR U2904 ( .A(n2909), .B(n2913), .Z(n2911) );
  XNOR U2905 ( .A(n2895), .B(n2892), .Z(n2902) );
  AND U2906 ( .A(n2914), .B(n2915), .Z(n2892) );
  XOR U2907 ( .A(n2916), .B(n2917), .Z(n2895) );
  AND U2908 ( .A(n2918), .B(n2919), .Z(n2917) );
  XOR U2909 ( .A(n2916), .B(n2920), .Z(n2918) );
  XNOR U2910 ( .A(n2846), .B(n2898), .Z(n2900) );
  XNOR U2911 ( .A(n2921), .B(n2922), .Z(n2846) );
  AND U2912 ( .A(n111), .B(n2852), .Z(n2922) );
  XOR U2913 ( .A(n2921), .B(n2850), .Z(n2852) );
  XOR U2914 ( .A(n2923), .B(n2924), .Z(n2898) );
  AND U2915 ( .A(n2925), .B(n2926), .Z(n2924) );
  XNOR U2916 ( .A(n2923), .B(n2914), .Z(n2926) );
  IV U2917 ( .A(n2858), .Z(n2914) );
  XNOR U2918 ( .A(n2927), .B(n2907), .Z(n2858) );
  XNOR U2919 ( .A(n2928), .B(n2913), .Z(n2907) );
  XOR U2920 ( .A(n2929), .B(n2930), .Z(n2913) );
  AND U2921 ( .A(n2931), .B(n2932), .Z(n2930) );
  XOR U2922 ( .A(n2929), .B(n2933), .Z(n2931) );
  XNOR U2923 ( .A(n2912), .B(n2904), .Z(n2928) );
  XOR U2924 ( .A(n2934), .B(n2935), .Z(n2904) );
  AND U2925 ( .A(n2936), .B(n2937), .Z(n2935) );
  XNOR U2926 ( .A(n2938), .B(n2934), .Z(n2936) );
  XNOR U2927 ( .A(n2939), .B(n2909), .Z(n2912) );
  XOR U2928 ( .A(n2940), .B(n2941), .Z(n2909) );
  AND U2929 ( .A(n2942), .B(n2943), .Z(n2941) );
  XOR U2930 ( .A(n2940), .B(n2944), .Z(n2942) );
  XNOR U2931 ( .A(n2945), .B(n2946), .Z(n2939) );
  AND U2932 ( .A(n2947), .B(n2948), .Z(n2946) );
  XNOR U2933 ( .A(n2945), .B(n2949), .Z(n2947) );
  XNOR U2934 ( .A(n2908), .B(n2915), .Z(n2927) );
  AND U2935 ( .A(n2870), .B(n2950), .Z(n2915) );
  XOR U2936 ( .A(n2920), .B(n2919), .Z(n2908) );
  XNOR U2937 ( .A(n2951), .B(n2916), .Z(n2919) );
  XOR U2938 ( .A(n2952), .B(n2953), .Z(n2916) );
  AND U2939 ( .A(n2954), .B(n2955), .Z(n2953) );
  XOR U2940 ( .A(n2952), .B(n2956), .Z(n2954) );
  XNOR U2941 ( .A(n2957), .B(n2958), .Z(n2951) );
  AND U2942 ( .A(n2959), .B(n2960), .Z(n2958) );
  XOR U2943 ( .A(n2957), .B(n2961), .Z(n2959) );
  XOR U2944 ( .A(n2962), .B(n2963), .Z(n2920) );
  AND U2945 ( .A(n2964), .B(n2965), .Z(n2963) );
  XOR U2946 ( .A(n2962), .B(n2966), .Z(n2964) );
  XNOR U2947 ( .A(n2855), .B(n2923), .Z(n2925) );
  XNOR U2948 ( .A(n2967), .B(n2968), .Z(n2855) );
  AND U2949 ( .A(n111), .B(n2862), .Z(n2968) );
  XOR U2950 ( .A(n2967), .B(n2860), .Z(n2862) );
  XOR U2951 ( .A(n2969), .B(n2970), .Z(n2923) );
  AND U2952 ( .A(n2971), .B(n2972), .Z(n2970) );
  XNOR U2953 ( .A(n2969), .B(n2870), .Z(n2972) );
  XOR U2954 ( .A(n2973), .B(n2937), .Z(n2870) );
  XNOR U2955 ( .A(n2974), .B(n2944), .Z(n2937) );
  XOR U2956 ( .A(n2933), .B(n2932), .Z(n2944) );
  XNOR U2957 ( .A(n2975), .B(n2929), .Z(n2932) );
  XOR U2958 ( .A(n2976), .B(n2977), .Z(n2929) );
  AND U2959 ( .A(n2978), .B(n2979), .Z(n2977) );
  XNOR U2960 ( .A(n2980), .B(n2981), .Z(n2978) );
  IV U2961 ( .A(n2976), .Z(n2980) );
  XNOR U2962 ( .A(n2982), .B(n2983), .Z(n2975) );
  NOR U2963 ( .A(n2984), .B(n2985), .Z(n2983) );
  XNOR U2964 ( .A(n2982), .B(n2986), .Z(n2984) );
  XOR U2965 ( .A(n2987), .B(n2988), .Z(n2933) );
  NOR U2966 ( .A(n2989), .B(n2990), .Z(n2988) );
  XNOR U2967 ( .A(n2987), .B(n2991), .Z(n2989) );
  XNOR U2968 ( .A(n2943), .B(n2934), .Z(n2974) );
  XOR U2969 ( .A(n2992), .B(n2993), .Z(n2934) );
  AND U2970 ( .A(n2994), .B(n2995), .Z(n2993) );
  XOR U2971 ( .A(n2992), .B(n2996), .Z(n2994) );
  XOR U2972 ( .A(n2997), .B(n2949), .Z(n2943) );
  XOR U2973 ( .A(n2998), .B(n2999), .Z(n2949) );
  NOR U2974 ( .A(n3000), .B(n3001), .Z(n2999) );
  XOR U2975 ( .A(n2998), .B(n3002), .Z(n3000) );
  XNOR U2976 ( .A(n2948), .B(n2940), .Z(n2997) );
  XOR U2977 ( .A(n3003), .B(n3004), .Z(n2940) );
  AND U2978 ( .A(n3005), .B(n3006), .Z(n3004) );
  XOR U2979 ( .A(n3003), .B(n3007), .Z(n3005) );
  XNOR U2980 ( .A(n3008), .B(n2945), .Z(n2948) );
  XOR U2981 ( .A(n3009), .B(n3010), .Z(n2945) );
  AND U2982 ( .A(n3011), .B(n3012), .Z(n3010) );
  XNOR U2983 ( .A(n3013), .B(n3014), .Z(n3011) );
  IV U2984 ( .A(n3009), .Z(n3013) );
  XNOR U2985 ( .A(n3015), .B(n3016), .Z(n3008) );
  NOR U2986 ( .A(n3017), .B(n3018), .Z(n3016) );
  XNOR U2987 ( .A(n3015), .B(n3019), .Z(n3017) );
  XOR U2988 ( .A(n2938), .B(n2950), .Z(n2973) );
  NOR U2989 ( .A(n2878), .B(n3020), .Z(n2950) );
  XNOR U2990 ( .A(n2956), .B(n2955), .Z(n2938) );
  XNOR U2991 ( .A(n3021), .B(n2961), .Z(n2955) );
  XNOR U2992 ( .A(n3022), .B(n3023), .Z(n2961) );
  NOR U2993 ( .A(n3024), .B(n3025), .Z(n3023) );
  XOR U2994 ( .A(n3022), .B(n3026), .Z(n3024) );
  XNOR U2995 ( .A(n2960), .B(n2952), .Z(n3021) );
  XOR U2996 ( .A(n3027), .B(n3028), .Z(n2952) );
  AND U2997 ( .A(n3029), .B(n3030), .Z(n3028) );
  XNOR U2998 ( .A(n3031), .B(n3032), .Z(n3029) );
  XNOR U2999 ( .A(n3033), .B(n2957), .Z(n2960) );
  XOR U3000 ( .A(n3034), .B(n3035), .Z(n2957) );
  AND U3001 ( .A(n3036), .B(n3037), .Z(n3035) );
  XNOR U3002 ( .A(n3038), .B(n3039), .Z(n3036) );
  IV U3003 ( .A(n3034), .Z(n3038) );
  XNOR U3004 ( .A(n3040), .B(n3041), .Z(n3033) );
  NOR U3005 ( .A(n3042), .B(n3043), .Z(n3041) );
  XNOR U3006 ( .A(n3040), .B(n3044), .Z(n3042) );
  XOR U3007 ( .A(n2966), .B(n2965), .Z(n2956) );
  XNOR U3008 ( .A(n3045), .B(n2962), .Z(n2965) );
  XOR U3009 ( .A(n3046), .B(n3047), .Z(n2962) );
  AND U3010 ( .A(n3048), .B(n3049), .Z(n3047) );
  XOR U3011 ( .A(n3046), .B(n3050), .Z(n3048) );
  XNOR U3012 ( .A(n3051), .B(n3052), .Z(n3045) );
  NOR U3013 ( .A(n3053), .B(n3054), .Z(n3052) );
  XNOR U3014 ( .A(n3051), .B(n3055), .Z(n3053) );
  XOR U3015 ( .A(n3056), .B(n3057), .Z(n2966) );
  NOR U3016 ( .A(n3058), .B(n3059), .Z(n3057) );
  XNOR U3017 ( .A(n3056), .B(n3060), .Z(n3058) );
  XNOR U3018 ( .A(n2867), .B(n2969), .Z(n2971) );
  XNOR U3019 ( .A(n3061), .B(n3062), .Z(n2867) );
  AND U3020 ( .A(n111), .B(n2874), .Z(n3062) );
  XOR U3021 ( .A(n3061), .B(n2872), .Z(n2874) );
  AND U3022 ( .A(n2875), .B(n2878), .Z(n2969) );
  XOR U3023 ( .A(n3063), .B(n3020), .Z(n2878) );
  XNOR U3024 ( .A(p_input[128]), .B(p_input[256]), .Z(n3020) );
  XNOR U3025 ( .A(n2996), .B(n2995), .Z(n3063) );
  XNOR U3026 ( .A(n3064), .B(n3007), .Z(n2995) );
  XOR U3027 ( .A(n2981), .B(n2979), .Z(n3007) );
  XNOR U3028 ( .A(n3065), .B(n2986), .Z(n2979) );
  XOR U3029 ( .A(p_input[152]), .B(p_input[280]), .Z(n2986) );
  XOR U3030 ( .A(n2976), .B(n2985), .Z(n3065) );
  XOR U3031 ( .A(n3066), .B(n2982), .Z(n2985) );
  XOR U3032 ( .A(p_input[150]), .B(p_input[278]), .Z(n2982) );
  XOR U3033 ( .A(p_input[151]), .B(n1937), .Z(n3066) );
  XOR U3034 ( .A(p_input[146]), .B(p_input[274]), .Z(n2976) );
  XNOR U3035 ( .A(n2991), .B(n2990), .Z(n2981) );
  XOR U3036 ( .A(n3067), .B(n2987), .Z(n2990) );
  XOR U3037 ( .A(p_input[147]), .B(p_input[275]), .Z(n2987) );
  XOR U3038 ( .A(p_input[148]), .B(n1939), .Z(n3067) );
  XOR U3039 ( .A(p_input[149]), .B(p_input[277]), .Z(n2991) );
  XOR U3040 ( .A(n3006), .B(n3068), .Z(n3064) );
  IV U3041 ( .A(n2992), .Z(n3068) );
  XOR U3042 ( .A(p_input[129]), .B(p_input[257]), .Z(n2992) );
  XNOR U3043 ( .A(n3069), .B(n3014), .Z(n3006) );
  XNOR U3044 ( .A(n3002), .B(n3001), .Z(n3014) );
  XNOR U3045 ( .A(n3070), .B(n2998), .Z(n3001) );
  XNOR U3046 ( .A(p_input[154]), .B(p_input[282]), .Z(n2998) );
  XOR U3047 ( .A(p_input[155]), .B(n1943), .Z(n3070) );
  XOR U3048 ( .A(p_input[156]), .B(p_input[284]), .Z(n3002) );
  XOR U3049 ( .A(n3012), .B(n3071), .Z(n3069) );
  IV U3050 ( .A(n3003), .Z(n3071) );
  XOR U3051 ( .A(p_input[145]), .B(p_input[273]), .Z(n3003) );
  XNOR U3052 ( .A(n3072), .B(n3019), .Z(n3012) );
  XOR U3053 ( .A(p_input[159]), .B(p_input[287]), .Z(n3019) );
  XOR U3054 ( .A(n3009), .B(n3018), .Z(n3072) );
  XOR U3055 ( .A(n3073), .B(n3015), .Z(n3018) );
  XOR U3056 ( .A(p_input[157]), .B(p_input[285]), .Z(n3015) );
  XOR U3057 ( .A(p_input[158]), .B(n3074), .Z(n3073) );
  XOR U3058 ( .A(p_input[153]), .B(p_input[281]), .Z(n3009) );
  XOR U3059 ( .A(n3032), .B(n3030), .Z(n2996) );
  XNOR U3060 ( .A(n3075), .B(n3039), .Z(n3030) );
  XNOR U3061 ( .A(n3026), .B(n3025), .Z(n3039) );
  XNOR U3062 ( .A(n3076), .B(n3022), .Z(n3025) );
  XNOR U3063 ( .A(p_input[139]), .B(p_input[267]), .Z(n3022) );
  XOR U3064 ( .A(p_input[140]), .B(n1949), .Z(n3076) );
  XOR U3065 ( .A(p_input[141]), .B(p_input[269]), .Z(n3026) );
  XOR U3066 ( .A(n3037), .B(n3031), .Z(n3075) );
  IV U3067 ( .A(n3027), .Z(n3031) );
  XOR U3068 ( .A(p_input[130]), .B(p_input[258]), .Z(n3027) );
  XNOR U3069 ( .A(n3077), .B(n3044), .Z(n3037) );
  XNOR U3070 ( .A(p_input[144]), .B(n1951), .Z(n3044) );
  XOR U3071 ( .A(n3034), .B(n3043), .Z(n3077) );
  XOR U3072 ( .A(n3078), .B(n3040), .Z(n3043) );
  XOR U3073 ( .A(p_input[142]), .B(p_input[270]), .Z(n3040) );
  XOR U3074 ( .A(p_input[143]), .B(n1953), .Z(n3078) );
  XOR U3075 ( .A(p_input[138]), .B(p_input[266]), .Z(n3034) );
  XOR U3076 ( .A(n3050), .B(n3049), .Z(n3032) );
  XNOR U3077 ( .A(n3079), .B(n3055), .Z(n3049) );
  XOR U3078 ( .A(p_input[137]), .B(p_input[265]), .Z(n3055) );
  XOR U3079 ( .A(n3046), .B(n3054), .Z(n3079) );
  XOR U3080 ( .A(n3080), .B(n3051), .Z(n3054) );
  XOR U3081 ( .A(p_input[135]), .B(p_input[263]), .Z(n3051) );
  XOR U3082 ( .A(p_input[136]), .B(n3081), .Z(n3080) );
  XOR U3083 ( .A(p_input[131]), .B(p_input[259]), .Z(n3046) );
  XNOR U3084 ( .A(n3060), .B(n3059), .Z(n3050) );
  XOR U3085 ( .A(n3082), .B(n3056), .Z(n3059) );
  XOR U3086 ( .A(p_input[132]), .B(p_input[260]), .Z(n3056) );
  XOR U3087 ( .A(p_input[133]), .B(n3083), .Z(n3082) );
  XOR U3088 ( .A(p_input[134]), .B(p_input[262]), .Z(n3060) );
  XNOR U3089 ( .A(n3084), .B(n3085), .Z(n2875) );
  AND U3090 ( .A(n111), .B(n3086), .Z(n3085) );
  XNOR U3091 ( .A(n3087), .B(n3088), .Z(n111) );
  NOR U3092 ( .A(n3089), .B(n3090), .Z(n3088) );
  XOR U3093 ( .A(n2826), .B(n3087), .Z(n3090) );
  NOR U3094 ( .A(n3087), .B(n2825), .Z(n3089) );
  XOR U3095 ( .A(n3091), .B(n3092), .Z(n3087) );
  AND U3096 ( .A(n3093), .B(n3094), .Z(n3092) );
  XNOR U3097 ( .A(n2896), .B(n3091), .Z(n3094) );
  XOR U3098 ( .A(n3091), .B(n2839), .Z(n3093) );
  XOR U3099 ( .A(n3095), .B(n3096), .Z(n3091) );
  AND U3100 ( .A(n3097), .B(n3098), .Z(n3096) );
  XNOR U3101 ( .A(n2921), .B(n3095), .Z(n3098) );
  XOR U3102 ( .A(n3095), .B(n2850), .Z(n3097) );
  XOR U3103 ( .A(n3099), .B(n3100), .Z(n3095) );
  AND U3104 ( .A(n3101), .B(n3102), .Z(n3100) );
  XOR U3105 ( .A(n3099), .B(n2860), .Z(n3101) );
  XOR U3106 ( .A(n3103), .B(n3104), .Z(n2818) );
  AND U3107 ( .A(n115), .B(n3086), .Z(n3104) );
  XNOR U3108 ( .A(n3084), .B(n3103), .Z(n3086) );
  XNOR U3109 ( .A(n3105), .B(n3106), .Z(n115) );
  NOR U3110 ( .A(n3107), .B(n3108), .Z(n3106) );
  XNOR U3111 ( .A(n2826), .B(n3109), .Z(n3108) );
  IV U3112 ( .A(n3105), .Z(n3109) );
  AND U3113 ( .A(n3110), .B(n3111), .Z(n2826) );
  NOR U3114 ( .A(n3105), .B(n2825), .Z(n3107) );
  AND U3115 ( .A(n3112), .B(n3113), .Z(n2825) );
  IV U3116 ( .A(n3114), .Z(n3112) );
  XOR U3117 ( .A(n3115), .B(n3116), .Z(n3105) );
  AND U3118 ( .A(n3117), .B(n3118), .Z(n3116) );
  XNOR U3119 ( .A(n3115), .B(n2896), .Z(n3118) );
  XNOR U3120 ( .A(n3119), .B(n3120), .Z(n2896) );
  AND U3121 ( .A(n118), .B(n3121), .Z(n3120) );
  XOR U3122 ( .A(n3122), .B(n3119), .Z(n3121) );
  XNOR U3123 ( .A(n3123), .B(n3115), .Z(n3117) );
  IV U3124 ( .A(n2839), .Z(n3123) );
  XOR U3125 ( .A(n3124), .B(n3125), .Z(n2839) );
  AND U3126 ( .A(n125), .B(n3126), .Z(n3125) );
  XOR U3127 ( .A(n3127), .B(n3128), .Z(n3115) );
  AND U3128 ( .A(n3129), .B(n3130), .Z(n3128) );
  XNOR U3129 ( .A(n3127), .B(n2921), .Z(n3130) );
  XNOR U3130 ( .A(n3131), .B(n3132), .Z(n2921) );
  AND U3131 ( .A(n118), .B(n3133), .Z(n3132) );
  XNOR U3132 ( .A(n3134), .B(n3131), .Z(n3133) );
  XOR U3133 ( .A(n2850), .B(n3127), .Z(n3129) );
  XOR U3134 ( .A(n3135), .B(n3136), .Z(n2850) );
  AND U3135 ( .A(n125), .B(n3137), .Z(n3136) );
  XOR U3136 ( .A(n3099), .B(n3138), .Z(n3127) );
  AND U3137 ( .A(n3139), .B(n3102), .Z(n3138) );
  XNOR U3138 ( .A(n2967), .B(n3099), .Z(n3102) );
  XNOR U3139 ( .A(n3140), .B(n3141), .Z(n2967) );
  AND U3140 ( .A(n118), .B(n3142), .Z(n3141) );
  XOR U3141 ( .A(n3143), .B(n3140), .Z(n3142) );
  XNOR U3142 ( .A(n3144), .B(n3099), .Z(n3139) );
  IV U3143 ( .A(n2860), .Z(n3144) );
  XOR U3144 ( .A(n3145), .B(n3146), .Z(n2860) );
  AND U3145 ( .A(n125), .B(n3147), .Z(n3146) );
  XOR U3146 ( .A(n3148), .B(n3149), .Z(n3099) );
  AND U3147 ( .A(n3150), .B(n3151), .Z(n3149) );
  XNOR U3148 ( .A(n3148), .B(n3061), .Z(n3151) );
  XNOR U3149 ( .A(n3152), .B(n3153), .Z(n3061) );
  AND U3150 ( .A(n118), .B(n3154), .Z(n3153) );
  XNOR U3151 ( .A(n3155), .B(n3152), .Z(n3154) );
  XNOR U3152 ( .A(n3156), .B(n3148), .Z(n3150) );
  IV U3153 ( .A(n2872), .Z(n3156) );
  XOR U3154 ( .A(n3157), .B(n3158), .Z(n2872) );
  AND U3155 ( .A(n125), .B(n3159), .Z(n3158) );
  AND U3156 ( .A(n3103), .B(n3084), .Z(n3148) );
  XNOR U3157 ( .A(n3160), .B(n3161), .Z(n3084) );
  AND U3158 ( .A(n118), .B(n3162), .Z(n3161) );
  XNOR U3159 ( .A(n3163), .B(n3160), .Z(n3162) );
  XNOR U3160 ( .A(n3164), .B(n3165), .Z(n118) );
  NOR U3161 ( .A(n3166), .B(n3167), .Z(n3165) );
  XNOR U3162 ( .A(n3164), .B(n3114), .Z(n3167) );
  NOR U3163 ( .A(n3110), .B(n3111), .Z(n3114) );
  NOR U3164 ( .A(n3164), .B(n3113), .Z(n3166) );
  AND U3165 ( .A(n3168), .B(n3169), .Z(n3113) );
  XOR U3166 ( .A(n3170), .B(n3171), .Z(n3164) );
  AND U3167 ( .A(n3172), .B(n3173), .Z(n3171) );
  XNOR U3168 ( .A(n3170), .B(n3168), .Z(n3173) );
  IV U3169 ( .A(n3122), .Z(n3168) );
  XOR U3170 ( .A(n3174), .B(n3175), .Z(n3122) );
  XOR U3171 ( .A(n3176), .B(n3169), .Z(n3175) );
  AND U3172 ( .A(n3134), .B(n3177), .Z(n3169) );
  AND U3173 ( .A(n3178), .B(n3179), .Z(n3176) );
  XOR U3174 ( .A(n3180), .B(n3174), .Z(n3178) );
  XNOR U3175 ( .A(n3119), .B(n3170), .Z(n3172) );
  XNOR U3176 ( .A(n3181), .B(n3182), .Z(n3119) );
  AND U3177 ( .A(n122), .B(n3126), .Z(n3182) );
  XOR U3178 ( .A(n3181), .B(n3124), .Z(n3126) );
  XOR U3179 ( .A(n3183), .B(n3184), .Z(n3170) );
  AND U3180 ( .A(n3185), .B(n3186), .Z(n3184) );
  XNOR U3181 ( .A(n3183), .B(n3134), .Z(n3186) );
  XOR U3182 ( .A(n3187), .B(n3179), .Z(n3134) );
  XNOR U3183 ( .A(n3188), .B(n3174), .Z(n3179) );
  XOR U3184 ( .A(n3189), .B(n3190), .Z(n3174) );
  AND U3185 ( .A(n3191), .B(n3192), .Z(n3190) );
  XOR U3186 ( .A(n3193), .B(n3189), .Z(n3191) );
  XNOR U3187 ( .A(n3194), .B(n3195), .Z(n3188) );
  AND U3188 ( .A(n3196), .B(n3197), .Z(n3195) );
  XOR U3189 ( .A(n3194), .B(n3198), .Z(n3196) );
  XNOR U3190 ( .A(n3180), .B(n3177), .Z(n3187) );
  AND U3191 ( .A(n3199), .B(n3200), .Z(n3177) );
  XOR U3192 ( .A(n3201), .B(n3202), .Z(n3180) );
  AND U3193 ( .A(n3203), .B(n3204), .Z(n3202) );
  XOR U3194 ( .A(n3201), .B(n3205), .Z(n3203) );
  XNOR U3195 ( .A(n3131), .B(n3183), .Z(n3185) );
  XNOR U3196 ( .A(n3206), .B(n3207), .Z(n3131) );
  AND U3197 ( .A(n122), .B(n3137), .Z(n3207) );
  XOR U3198 ( .A(n3206), .B(n3135), .Z(n3137) );
  XOR U3199 ( .A(n3208), .B(n3209), .Z(n3183) );
  AND U3200 ( .A(n3210), .B(n3211), .Z(n3209) );
  XNOR U3201 ( .A(n3208), .B(n3199), .Z(n3211) );
  IV U3202 ( .A(n3143), .Z(n3199) );
  XNOR U3203 ( .A(n3212), .B(n3192), .Z(n3143) );
  XNOR U3204 ( .A(n3213), .B(n3198), .Z(n3192) );
  XOR U3205 ( .A(n3214), .B(n3215), .Z(n3198) );
  AND U3206 ( .A(n3216), .B(n3217), .Z(n3215) );
  XOR U3207 ( .A(n3214), .B(n3218), .Z(n3216) );
  XNOR U3208 ( .A(n3197), .B(n3189), .Z(n3213) );
  XOR U3209 ( .A(n3219), .B(n3220), .Z(n3189) );
  AND U3210 ( .A(n3221), .B(n3222), .Z(n3220) );
  XNOR U3211 ( .A(n3223), .B(n3219), .Z(n3221) );
  XNOR U3212 ( .A(n3224), .B(n3194), .Z(n3197) );
  XOR U3213 ( .A(n3225), .B(n3226), .Z(n3194) );
  AND U3214 ( .A(n3227), .B(n3228), .Z(n3226) );
  XOR U3215 ( .A(n3225), .B(n3229), .Z(n3227) );
  XNOR U3216 ( .A(n3230), .B(n3231), .Z(n3224) );
  AND U3217 ( .A(n3232), .B(n3233), .Z(n3231) );
  XNOR U3218 ( .A(n3230), .B(n3234), .Z(n3232) );
  XNOR U3219 ( .A(n3193), .B(n3200), .Z(n3212) );
  AND U3220 ( .A(n3155), .B(n3235), .Z(n3200) );
  XOR U3221 ( .A(n3205), .B(n3204), .Z(n3193) );
  XNOR U3222 ( .A(n3236), .B(n3201), .Z(n3204) );
  XOR U3223 ( .A(n3237), .B(n3238), .Z(n3201) );
  AND U3224 ( .A(n3239), .B(n3240), .Z(n3238) );
  XOR U3225 ( .A(n3237), .B(n3241), .Z(n3239) );
  XNOR U3226 ( .A(n3242), .B(n3243), .Z(n3236) );
  AND U3227 ( .A(n3244), .B(n3245), .Z(n3243) );
  XOR U3228 ( .A(n3242), .B(n3246), .Z(n3244) );
  XOR U3229 ( .A(n3247), .B(n3248), .Z(n3205) );
  AND U3230 ( .A(n3249), .B(n3250), .Z(n3248) );
  XOR U3231 ( .A(n3247), .B(n3251), .Z(n3249) );
  XNOR U3232 ( .A(n3140), .B(n3208), .Z(n3210) );
  XNOR U3233 ( .A(n3252), .B(n3253), .Z(n3140) );
  AND U3234 ( .A(n122), .B(n3147), .Z(n3253) );
  XOR U3235 ( .A(n3252), .B(n3145), .Z(n3147) );
  XOR U3236 ( .A(n3254), .B(n3255), .Z(n3208) );
  AND U3237 ( .A(n3256), .B(n3257), .Z(n3255) );
  XNOR U3238 ( .A(n3254), .B(n3155), .Z(n3257) );
  XOR U3239 ( .A(n3258), .B(n3222), .Z(n3155) );
  XNOR U3240 ( .A(n3259), .B(n3229), .Z(n3222) );
  XOR U3241 ( .A(n3218), .B(n3217), .Z(n3229) );
  XNOR U3242 ( .A(n3260), .B(n3214), .Z(n3217) );
  XOR U3243 ( .A(n3261), .B(n3262), .Z(n3214) );
  AND U3244 ( .A(n3263), .B(n3264), .Z(n3262) );
  XNOR U3245 ( .A(n3265), .B(n3266), .Z(n3263) );
  IV U3246 ( .A(n3261), .Z(n3265) );
  XNOR U3247 ( .A(n3267), .B(n3268), .Z(n3260) );
  NOR U3248 ( .A(n3269), .B(n3270), .Z(n3268) );
  XNOR U3249 ( .A(n3267), .B(n3271), .Z(n3269) );
  XOR U3250 ( .A(n3272), .B(n3273), .Z(n3218) );
  NOR U3251 ( .A(n3274), .B(n3275), .Z(n3273) );
  XNOR U3252 ( .A(n3272), .B(n3276), .Z(n3274) );
  XNOR U3253 ( .A(n3228), .B(n3219), .Z(n3259) );
  XOR U3254 ( .A(n3277), .B(n3278), .Z(n3219) );
  AND U3255 ( .A(n3279), .B(n3280), .Z(n3278) );
  XOR U3256 ( .A(n3277), .B(n3281), .Z(n3279) );
  XOR U3257 ( .A(n3282), .B(n3234), .Z(n3228) );
  XOR U3258 ( .A(n3283), .B(n3284), .Z(n3234) );
  NOR U3259 ( .A(n3285), .B(n3286), .Z(n3284) );
  XOR U3260 ( .A(n3283), .B(n3287), .Z(n3285) );
  XNOR U3261 ( .A(n3233), .B(n3225), .Z(n3282) );
  XOR U3262 ( .A(n3288), .B(n3289), .Z(n3225) );
  AND U3263 ( .A(n3290), .B(n3291), .Z(n3289) );
  XOR U3264 ( .A(n3288), .B(n3292), .Z(n3290) );
  XNOR U3265 ( .A(n3293), .B(n3230), .Z(n3233) );
  XOR U3266 ( .A(n3294), .B(n3295), .Z(n3230) );
  AND U3267 ( .A(n3296), .B(n3297), .Z(n3295) );
  XNOR U3268 ( .A(n3298), .B(n3299), .Z(n3296) );
  IV U3269 ( .A(n3294), .Z(n3298) );
  XNOR U3270 ( .A(n3300), .B(n3301), .Z(n3293) );
  NOR U3271 ( .A(n3302), .B(n3303), .Z(n3301) );
  XNOR U3272 ( .A(n3300), .B(n3304), .Z(n3302) );
  XOR U3273 ( .A(n3223), .B(n3235), .Z(n3258) );
  NOR U3274 ( .A(n3163), .B(n3305), .Z(n3235) );
  XNOR U3275 ( .A(n3241), .B(n3240), .Z(n3223) );
  XNOR U3276 ( .A(n3306), .B(n3246), .Z(n3240) );
  XNOR U3277 ( .A(n3307), .B(n3308), .Z(n3246) );
  NOR U3278 ( .A(n3309), .B(n3310), .Z(n3308) );
  XOR U3279 ( .A(n3307), .B(n3311), .Z(n3309) );
  XNOR U3280 ( .A(n3245), .B(n3237), .Z(n3306) );
  XOR U3281 ( .A(n3312), .B(n3313), .Z(n3237) );
  AND U3282 ( .A(n3314), .B(n3315), .Z(n3313) );
  XOR U3283 ( .A(n3312), .B(n3316), .Z(n3314) );
  XNOR U3284 ( .A(n3317), .B(n3242), .Z(n3245) );
  XOR U3285 ( .A(n3318), .B(n3319), .Z(n3242) );
  AND U3286 ( .A(n3320), .B(n3321), .Z(n3319) );
  XNOR U3287 ( .A(n3322), .B(n3323), .Z(n3320) );
  IV U3288 ( .A(n3318), .Z(n3322) );
  XNOR U3289 ( .A(n3324), .B(n3325), .Z(n3317) );
  NOR U3290 ( .A(n3326), .B(n3327), .Z(n3325) );
  XNOR U3291 ( .A(n3324), .B(n3328), .Z(n3326) );
  XOR U3292 ( .A(n3251), .B(n3250), .Z(n3241) );
  XNOR U3293 ( .A(n3329), .B(n3247), .Z(n3250) );
  XOR U3294 ( .A(n3330), .B(n3331), .Z(n3247) );
  AND U3295 ( .A(n3332), .B(n3333), .Z(n3331) );
  XNOR U3296 ( .A(n3334), .B(n3335), .Z(n3332) );
  XNOR U3297 ( .A(n3336), .B(n3337), .Z(n3329) );
  NOR U3298 ( .A(n3338), .B(n3339), .Z(n3337) );
  XNOR U3299 ( .A(n3336), .B(n3340), .Z(n3338) );
  XOR U3300 ( .A(n3341), .B(n3342), .Z(n3251) );
  NOR U3301 ( .A(n3343), .B(n3344), .Z(n3342) );
  XNOR U3302 ( .A(n3341), .B(n3345), .Z(n3343) );
  XNOR U3303 ( .A(n3152), .B(n3254), .Z(n3256) );
  XNOR U3304 ( .A(n3346), .B(n3347), .Z(n3152) );
  AND U3305 ( .A(n122), .B(n3159), .Z(n3347) );
  XOR U3306 ( .A(n3346), .B(n3157), .Z(n3159) );
  AND U3307 ( .A(n3160), .B(n3163), .Z(n3254) );
  XOR U3308 ( .A(n3348), .B(n3305), .Z(n3163) );
  XNOR U3309 ( .A(p_input[160]), .B(p_input[256]), .Z(n3305) );
  XNOR U3310 ( .A(n3281), .B(n3280), .Z(n3348) );
  XNOR U3311 ( .A(n3349), .B(n3292), .Z(n3280) );
  XOR U3312 ( .A(n3266), .B(n3264), .Z(n3292) );
  XNOR U3313 ( .A(n3350), .B(n3271), .Z(n3264) );
  XOR U3314 ( .A(p_input[184]), .B(p_input[280]), .Z(n3271) );
  XOR U3315 ( .A(n3261), .B(n3270), .Z(n3350) );
  XOR U3316 ( .A(n3351), .B(n3267), .Z(n3270) );
  XOR U3317 ( .A(p_input[182]), .B(p_input[278]), .Z(n3267) );
  XOR U3318 ( .A(p_input[183]), .B(n1937), .Z(n3351) );
  XOR U3319 ( .A(p_input[178]), .B(p_input[274]), .Z(n3261) );
  XNOR U3320 ( .A(n3276), .B(n3275), .Z(n3266) );
  XOR U3321 ( .A(n3352), .B(n3272), .Z(n3275) );
  XOR U3322 ( .A(p_input[179]), .B(p_input[275]), .Z(n3272) );
  XOR U3323 ( .A(p_input[180]), .B(n1939), .Z(n3352) );
  XOR U3324 ( .A(p_input[181]), .B(p_input[277]), .Z(n3276) );
  XOR U3325 ( .A(n3291), .B(n3353), .Z(n3349) );
  IV U3326 ( .A(n3277), .Z(n3353) );
  XOR U3327 ( .A(p_input[161]), .B(p_input[257]), .Z(n3277) );
  XNOR U3328 ( .A(n3354), .B(n3299), .Z(n3291) );
  XNOR U3329 ( .A(n3287), .B(n3286), .Z(n3299) );
  XNOR U3330 ( .A(n3355), .B(n3283), .Z(n3286) );
  XNOR U3331 ( .A(p_input[186]), .B(p_input[282]), .Z(n3283) );
  XOR U3332 ( .A(p_input[187]), .B(n1943), .Z(n3355) );
  XOR U3333 ( .A(p_input[188]), .B(p_input[284]), .Z(n3287) );
  XOR U3334 ( .A(n3297), .B(n3356), .Z(n3354) );
  IV U3335 ( .A(n3288), .Z(n3356) );
  XOR U3336 ( .A(p_input[177]), .B(p_input[273]), .Z(n3288) );
  XNOR U3337 ( .A(n3357), .B(n3304), .Z(n3297) );
  XOR U3338 ( .A(p_input[191]), .B(p_input[287]), .Z(n3304) );
  XOR U3339 ( .A(n3294), .B(n3303), .Z(n3357) );
  XOR U3340 ( .A(n3358), .B(n3300), .Z(n3303) );
  XOR U3341 ( .A(p_input[189]), .B(p_input[285]), .Z(n3300) );
  XOR U3342 ( .A(p_input[190]), .B(n3074), .Z(n3358) );
  XOR U3343 ( .A(p_input[185]), .B(p_input[281]), .Z(n3294) );
  XOR U3344 ( .A(n3316), .B(n3315), .Z(n3281) );
  XNOR U3345 ( .A(n3359), .B(n3323), .Z(n3315) );
  XNOR U3346 ( .A(n3311), .B(n3310), .Z(n3323) );
  XNOR U3347 ( .A(n3360), .B(n3307), .Z(n3310) );
  XNOR U3348 ( .A(p_input[171]), .B(p_input[267]), .Z(n3307) );
  XOR U3349 ( .A(p_input[172]), .B(n1949), .Z(n3360) );
  XOR U3350 ( .A(p_input[173]), .B(p_input[269]), .Z(n3311) );
  XNOR U3351 ( .A(n3321), .B(n3312), .Z(n3359) );
  XOR U3352 ( .A(p_input[162]), .B(p_input[258]), .Z(n3312) );
  XNOR U3353 ( .A(n3361), .B(n3328), .Z(n3321) );
  XNOR U3354 ( .A(p_input[176]), .B(n1951), .Z(n3328) );
  IV U3355 ( .A(p_input[272]), .Z(n1951) );
  XOR U3356 ( .A(n3318), .B(n3327), .Z(n3361) );
  XOR U3357 ( .A(n3362), .B(n3324), .Z(n3327) );
  XOR U3358 ( .A(p_input[174]), .B(p_input[270]), .Z(n3324) );
  XOR U3359 ( .A(p_input[175]), .B(n1953), .Z(n3362) );
  XOR U3360 ( .A(p_input[170]), .B(p_input[266]), .Z(n3318) );
  XOR U3361 ( .A(n3335), .B(n3333), .Z(n3316) );
  XNOR U3362 ( .A(n3363), .B(n3340), .Z(n3333) );
  XOR U3363 ( .A(p_input[169]), .B(p_input[265]), .Z(n3340) );
  XOR U3364 ( .A(n3330), .B(n3339), .Z(n3363) );
  XOR U3365 ( .A(n3364), .B(n3336), .Z(n3339) );
  XOR U3366 ( .A(p_input[167]), .B(p_input[263]), .Z(n3336) );
  XOR U3367 ( .A(p_input[168]), .B(n3081), .Z(n3364) );
  IV U3368 ( .A(n3334), .Z(n3330) );
  XNOR U3369 ( .A(p_input[163]), .B(p_input[259]), .Z(n3334) );
  XNOR U3370 ( .A(n3345), .B(n3344), .Z(n3335) );
  XOR U3371 ( .A(n3365), .B(n3341), .Z(n3344) );
  XOR U3372 ( .A(p_input[164]), .B(p_input[260]), .Z(n3341) );
  XOR U3373 ( .A(p_input[165]), .B(n3083), .Z(n3365) );
  XOR U3374 ( .A(p_input[166]), .B(p_input[262]), .Z(n3345) );
  XNOR U3375 ( .A(n3366), .B(n3367), .Z(n3160) );
  AND U3376 ( .A(n122), .B(n3368), .Z(n3367) );
  XNOR U3377 ( .A(n3369), .B(n3370), .Z(n122) );
  NOR U3378 ( .A(n3371), .B(n3372), .Z(n3370) );
  XOR U3379 ( .A(n3111), .B(n3369), .Z(n3372) );
  NOR U3380 ( .A(n3369), .B(n3110), .Z(n3371) );
  XOR U3381 ( .A(n3373), .B(n3374), .Z(n3369) );
  AND U3382 ( .A(n3375), .B(n3376), .Z(n3374) );
  XNOR U3383 ( .A(n3181), .B(n3373), .Z(n3376) );
  XOR U3384 ( .A(n3373), .B(n3124), .Z(n3375) );
  XOR U3385 ( .A(n3377), .B(n3378), .Z(n3373) );
  AND U3386 ( .A(n3379), .B(n3380), .Z(n3378) );
  XNOR U3387 ( .A(n3206), .B(n3377), .Z(n3380) );
  XOR U3388 ( .A(n3377), .B(n3135), .Z(n3379) );
  XOR U3389 ( .A(n3381), .B(n3382), .Z(n3377) );
  AND U3390 ( .A(n3383), .B(n3384), .Z(n3382) );
  XOR U3391 ( .A(n3381), .B(n3145), .Z(n3383) );
  XOR U3392 ( .A(n3385), .B(n3386), .Z(n3103) );
  AND U3393 ( .A(n125), .B(n3368), .Z(n3386) );
  XOR U3394 ( .A(n3387), .B(n3385), .Z(n3368) );
  XNOR U3395 ( .A(n3388), .B(n3389), .Z(n125) );
  NOR U3396 ( .A(n3390), .B(n3391), .Z(n3389) );
  XNOR U3397 ( .A(n3111), .B(n3392), .Z(n3391) );
  IV U3398 ( .A(n3388), .Z(n3392) );
  AND U3399 ( .A(n3124), .B(n3393), .Z(n3111) );
  NOR U3400 ( .A(n3388), .B(n3110), .Z(n3390) );
  AND U3401 ( .A(n3181), .B(n3394), .Z(n3110) );
  XOR U3402 ( .A(n3395), .B(n3396), .Z(n3388) );
  AND U3403 ( .A(n3397), .B(n3398), .Z(n3396) );
  XNOR U3404 ( .A(n3395), .B(n3181), .Z(n3398) );
  XNOR U3405 ( .A(n3399), .B(n3400), .Z(n3181) );
  XOR U3406 ( .A(n3401), .B(n3394), .Z(n3400) );
  AND U3407 ( .A(n3206), .B(n3402), .Z(n3394) );
  AND U3408 ( .A(n3403), .B(n3404), .Z(n3401) );
  XOR U3409 ( .A(n3405), .B(n3399), .Z(n3403) );
  XNOR U3410 ( .A(n3406), .B(n3395), .Z(n3397) );
  IV U3411 ( .A(n3124), .Z(n3406) );
  XNOR U3412 ( .A(n3407), .B(n3408), .Z(n3124) );
  XOR U3413 ( .A(n3409), .B(n3393), .Z(n3408) );
  AND U3414 ( .A(n3135), .B(n3410), .Z(n3393) );
  AND U3415 ( .A(n3411), .B(n3412), .Z(n3409) );
  XNOR U3416 ( .A(n3407), .B(n3413), .Z(n3411) );
  XOR U3417 ( .A(n3414), .B(n3415), .Z(n3395) );
  AND U3418 ( .A(n3416), .B(n3417), .Z(n3415) );
  XNOR U3419 ( .A(n3414), .B(n3206), .Z(n3417) );
  XOR U3420 ( .A(n3418), .B(n3404), .Z(n3206) );
  XNOR U3421 ( .A(n3419), .B(n3399), .Z(n3404) );
  XOR U3422 ( .A(n3420), .B(n3421), .Z(n3399) );
  AND U3423 ( .A(n3422), .B(n3423), .Z(n3421) );
  XOR U3424 ( .A(n3424), .B(n3420), .Z(n3422) );
  XNOR U3425 ( .A(n3425), .B(n3426), .Z(n3419) );
  AND U3426 ( .A(n3427), .B(n3428), .Z(n3426) );
  XOR U3427 ( .A(n3425), .B(n3429), .Z(n3427) );
  XNOR U3428 ( .A(n3405), .B(n3402), .Z(n3418) );
  AND U3429 ( .A(n3252), .B(n3430), .Z(n3402) );
  XOR U3430 ( .A(n3431), .B(n3432), .Z(n3405) );
  AND U3431 ( .A(n3433), .B(n3434), .Z(n3432) );
  XOR U3432 ( .A(n3431), .B(n3435), .Z(n3433) );
  XOR U3433 ( .A(n3135), .B(n3414), .Z(n3416) );
  XNOR U3434 ( .A(n3436), .B(n3413), .Z(n3135) );
  XNOR U3435 ( .A(n3437), .B(n3438), .Z(n3413) );
  AND U3436 ( .A(n3439), .B(n3440), .Z(n3438) );
  XOR U3437 ( .A(n3437), .B(n3441), .Z(n3439) );
  XNOR U3438 ( .A(n3412), .B(n3410), .Z(n3436) );
  AND U3439 ( .A(n3145), .B(n3442), .Z(n3410) );
  XNOR U3440 ( .A(n3443), .B(n3407), .Z(n3412) );
  XOR U3441 ( .A(n3444), .B(n3445), .Z(n3407) );
  AND U3442 ( .A(n3446), .B(n3447), .Z(n3445) );
  XOR U3443 ( .A(n3444), .B(n3448), .Z(n3446) );
  XNOR U3444 ( .A(n3449), .B(n3450), .Z(n3443) );
  AND U3445 ( .A(n3451), .B(n3452), .Z(n3450) );
  XNOR U3446 ( .A(n3449), .B(n3453), .Z(n3451) );
  XOR U3447 ( .A(n3381), .B(n3454), .Z(n3414) );
  AND U3448 ( .A(n3455), .B(n3384), .Z(n3454) );
  XNOR U3449 ( .A(n3252), .B(n3381), .Z(n3384) );
  XOR U3450 ( .A(n3456), .B(n3423), .Z(n3252) );
  XNOR U3451 ( .A(n3457), .B(n3429), .Z(n3423) );
  XOR U3452 ( .A(n3458), .B(n3459), .Z(n3429) );
  AND U3453 ( .A(n3460), .B(n3461), .Z(n3459) );
  XOR U3454 ( .A(n3458), .B(n3462), .Z(n3460) );
  XNOR U3455 ( .A(n3428), .B(n3420), .Z(n3457) );
  XOR U3456 ( .A(n3463), .B(n3464), .Z(n3420) );
  AND U3457 ( .A(n3465), .B(n3466), .Z(n3464) );
  XNOR U3458 ( .A(n3467), .B(n3463), .Z(n3465) );
  XNOR U3459 ( .A(n3468), .B(n3425), .Z(n3428) );
  XOR U3460 ( .A(n3469), .B(n3470), .Z(n3425) );
  AND U3461 ( .A(n3471), .B(n3472), .Z(n3470) );
  XOR U3462 ( .A(n3469), .B(n3473), .Z(n3471) );
  XNOR U3463 ( .A(n3474), .B(n3475), .Z(n3468) );
  AND U3464 ( .A(n3476), .B(n3477), .Z(n3475) );
  XNOR U3465 ( .A(n3474), .B(n3478), .Z(n3476) );
  XNOR U3466 ( .A(n3424), .B(n3430), .Z(n3456) );
  AND U3467 ( .A(n3346), .B(n3479), .Z(n3430) );
  XOR U3468 ( .A(n3435), .B(n3434), .Z(n3424) );
  XNOR U3469 ( .A(n3480), .B(n3431), .Z(n3434) );
  XOR U3470 ( .A(n3481), .B(n3482), .Z(n3431) );
  AND U3471 ( .A(n3483), .B(n3484), .Z(n3482) );
  XOR U3472 ( .A(n3481), .B(n3485), .Z(n3483) );
  XNOR U3473 ( .A(n3486), .B(n3487), .Z(n3480) );
  AND U3474 ( .A(n3488), .B(n3489), .Z(n3487) );
  XOR U3475 ( .A(n3486), .B(n3490), .Z(n3488) );
  XOR U3476 ( .A(n3491), .B(n3492), .Z(n3435) );
  AND U3477 ( .A(n3493), .B(n3494), .Z(n3492) );
  XOR U3478 ( .A(n3491), .B(n3495), .Z(n3493) );
  XNOR U3479 ( .A(n3496), .B(n3381), .Z(n3455) );
  IV U3480 ( .A(n3145), .Z(n3496) );
  XOR U3481 ( .A(n3497), .B(n3448), .Z(n3145) );
  XOR U3482 ( .A(n3441), .B(n3440), .Z(n3448) );
  XNOR U3483 ( .A(n3498), .B(n3437), .Z(n3440) );
  XOR U3484 ( .A(n3499), .B(n3500), .Z(n3437) );
  AND U3485 ( .A(n3501), .B(n3502), .Z(n3500) );
  XOR U3486 ( .A(n3499), .B(n3503), .Z(n3501) );
  XNOR U3487 ( .A(n3504), .B(n3505), .Z(n3498) );
  AND U3488 ( .A(n3506), .B(n3507), .Z(n3505) );
  XOR U3489 ( .A(n3504), .B(n3508), .Z(n3506) );
  XOR U3490 ( .A(n3509), .B(n3510), .Z(n3441) );
  AND U3491 ( .A(n3511), .B(n3512), .Z(n3510) );
  XOR U3492 ( .A(n3509), .B(n3513), .Z(n3511) );
  XNOR U3493 ( .A(n3447), .B(n3442), .Z(n3497) );
  AND U3494 ( .A(n3157), .B(n3514), .Z(n3442) );
  XOR U3495 ( .A(n3515), .B(n3453), .Z(n3447) );
  XNOR U3496 ( .A(n3516), .B(n3517), .Z(n3453) );
  AND U3497 ( .A(n3518), .B(n3519), .Z(n3517) );
  XOR U3498 ( .A(n3516), .B(n3520), .Z(n3518) );
  XNOR U3499 ( .A(n3452), .B(n3444), .Z(n3515) );
  XOR U3500 ( .A(n3521), .B(n3522), .Z(n3444) );
  AND U3501 ( .A(n3523), .B(n3524), .Z(n3522) );
  XOR U3502 ( .A(n3521), .B(n3525), .Z(n3523) );
  XNOR U3503 ( .A(n3526), .B(n3449), .Z(n3452) );
  XOR U3504 ( .A(n3527), .B(n3528), .Z(n3449) );
  AND U3505 ( .A(n3529), .B(n3530), .Z(n3528) );
  XOR U3506 ( .A(n3527), .B(n3531), .Z(n3529) );
  XNOR U3507 ( .A(n3532), .B(n3533), .Z(n3526) );
  AND U3508 ( .A(n3534), .B(n3535), .Z(n3533) );
  XNOR U3509 ( .A(n3532), .B(n3536), .Z(n3534) );
  XOR U3510 ( .A(n3537), .B(n3538), .Z(n3381) );
  AND U3511 ( .A(n3539), .B(n3540), .Z(n3538) );
  XNOR U3512 ( .A(n3537), .B(n3346), .Z(n3540) );
  XOR U3513 ( .A(n3541), .B(n3466), .Z(n3346) );
  XNOR U3514 ( .A(n3542), .B(n3473), .Z(n3466) );
  XOR U3515 ( .A(n3462), .B(n3461), .Z(n3473) );
  XNOR U3516 ( .A(n3543), .B(n3458), .Z(n3461) );
  XOR U3517 ( .A(n3544), .B(n3545), .Z(n3458) );
  AND U3518 ( .A(n3546), .B(n3547), .Z(n3545) );
  XOR U3519 ( .A(n3544), .B(n3548), .Z(n3546) );
  XNOR U3520 ( .A(n3549), .B(n3550), .Z(n3543) );
  NOR U3521 ( .A(n3551), .B(n3552), .Z(n3550) );
  XNOR U3522 ( .A(n3549), .B(n3553), .Z(n3551) );
  XOR U3523 ( .A(n3554), .B(n3555), .Z(n3462) );
  NOR U3524 ( .A(n3556), .B(n3557), .Z(n3555) );
  XNOR U3525 ( .A(n3554), .B(n3558), .Z(n3556) );
  XNOR U3526 ( .A(n3472), .B(n3463), .Z(n3542) );
  XOR U3527 ( .A(n3559), .B(n3560), .Z(n3463) );
  NOR U3528 ( .A(n3561), .B(n3562), .Z(n3560) );
  XNOR U3529 ( .A(n3559), .B(n3563), .Z(n3561) );
  XOR U3530 ( .A(n3564), .B(n3478), .Z(n3472) );
  XNOR U3531 ( .A(n3565), .B(n3566), .Z(n3478) );
  NOR U3532 ( .A(n3567), .B(n3568), .Z(n3566) );
  XNOR U3533 ( .A(n3565), .B(n3569), .Z(n3567) );
  XNOR U3534 ( .A(n3477), .B(n3469), .Z(n3564) );
  XOR U3535 ( .A(n3570), .B(n3571), .Z(n3469) );
  AND U3536 ( .A(n3572), .B(n3573), .Z(n3571) );
  XOR U3537 ( .A(n3570), .B(n3574), .Z(n3572) );
  XNOR U3538 ( .A(n3575), .B(n3474), .Z(n3477) );
  XOR U3539 ( .A(n3576), .B(n3577), .Z(n3474) );
  AND U3540 ( .A(n3578), .B(n3579), .Z(n3577) );
  XOR U3541 ( .A(n3576), .B(n3580), .Z(n3578) );
  XNOR U3542 ( .A(n3581), .B(n3582), .Z(n3575) );
  NOR U3543 ( .A(n3583), .B(n3584), .Z(n3582) );
  XOR U3544 ( .A(n3581), .B(n3585), .Z(n3583) );
  XOR U3545 ( .A(n3467), .B(n3479), .Z(n3541) );
  AND U3546 ( .A(n3387), .B(n3586), .Z(n3479) );
  IV U3547 ( .A(n3366), .Z(n3387) );
  XNOR U3548 ( .A(n3485), .B(n3484), .Z(n3467) );
  XNOR U3549 ( .A(n3587), .B(n3490), .Z(n3484) );
  XOR U3550 ( .A(n3588), .B(n3589), .Z(n3490) );
  NOR U3551 ( .A(n3590), .B(n3591), .Z(n3589) );
  XNOR U3552 ( .A(n3588), .B(n3592), .Z(n3590) );
  XNOR U3553 ( .A(n3489), .B(n3481), .Z(n3587) );
  XOR U3554 ( .A(n3593), .B(n3594), .Z(n3481) );
  AND U3555 ( .A(n3595), .B(n3596), .Z(n3594) );
  XNOR U3556 ( .A(n3593), .B(n3597), .Z(n3595) );
  XNOR U3557 ( .A(n3598), .B(n3486), .Z(n3489) );
  XOR U3558 ( .A(n3599), .B(n3600), .Z(n3486) );
  AND U3559 ( .A(n3601), .B(n3602), .Z(n3600) );
  XOR U3560 ( .A(n3599), .B(n3603), .Z(n3601) );
  XNOR U3561 ( .A(n3604), .B(n3605), .Z(n3598) );
  NOR U3562 ( .A(n3606), .B(n3607), .Z(n3605) );
  XOR U3563 ( .A(n3604), .B(n3608), .Z(n3606) );
  XOR U3564 ( .A(n3495), .B(n3494), .Z(n3485) );
  XNOR U3565 ( .A(n3609), .B(n3491), .Z(n3494) );
  XOR U3566 ( .A(n3610), .B(n3611), .Z(n3491) );
  AND U3567 ( .A(n3612), .B(n3613), .Z(n3611) );
  XOR U3568 ( .A(n3610), .B(n3614), .Z(n3612) );
  XNOR U3569 ( .A(n3615), .B(n3616), .Z(n3609) );
  NOR U3570 ( .A(n3617), .B(n3618), .Z(n3616) );
  XNOR U3571 ( .A(n3615), .B(n3619), .Z(n3617) );
  XOR U3572 ( .A(n3620), .B(n3621), .Z(n3495) );
  NOR U3573 ( .A(n3622), .B(n3623), .Z(n3621) );
  XNOR U3574 ( .A(n3620), .B(n3624), .Z(n3622) );
  XNOR U3575 ( .A(n3625), .B(n3537), .Z(n3539) );
  IV U3576 ( .A(n3157), .Z(n3625) );
  XOR U3577 ( .A(n3626), .B(n3525), .Z(n3157) );
  XOR U3578 ( .A(n3503), .B(n3502), .Z(n3525) );
  XNOR U3579 ( .A(n3627), .B(n3508), .Z(n3502) );
  XOR U3580 ( .A(n3628), .B(n3629), .Z(n3508) );
  NOR U3581 ( .A(n3630), .B(n3631), .Z(n3629) );
  XNOR U3582 ( .A(n3628), .B(n3632), .Z(n3630) );
  XNOR U3583 ( .A(n3507), .B(n3499), .Z(n3627) );
  XOR U3584 ( .A(n3633), .B(n3634), .Z(n3499) );
  AND U3585 ( .A(n3635), .B(n3636), .Z(n3634) );
  XNOR U3586 ( .A(n3633), .B(n3637), .Z(n3635) );
  XNOR U3587 ( .A(n3638), .B(n3504), .Z(n3507) );
  XOR U3588 ( .A(n3639), .B(n3640), .Z(n3504) );
  AND U3589 ( .A(n3641), .B(n3642), .Z(n3640) );
  XOR U3590 ( .A(n3639), .B(n3643), .Z(n3641) );
  XNOR U3591 ( .A(n3644), .B(n3645), .Z(n3638) );
  NOR U3592 ( .A(n3646), .B(n3647), .Z(n3645) );
  XOR U3593 ( .A(n3644), .B(n3648), .Z(n3646) );
  XOR U3594 ( .A(n3513), .B(n3512), .Z(n3503) );
  XNOR U3595 ( .A(n3649), .B(n3509), .Z(n3512) );
  XOR U3596 ( .A(n3650), .B(n3651), .Z(n3509) );
  AND U3597 ( .A(n3652), .B(n3653), .Z(n3651) );
  XOR U3598 ( .A(n3650), .B(n3654), .Z(n3652) );
  XNOR U3599 ( .A(n3655), .B(n3656), .Z(n3649) );
  NOR U3600 ( .A(n3657), .B(n3658), .Z(n3656) );
  XNOR U3601 ( .A(n3655), .B(n3659), .Z(n3657) );
  XOR U3602 ( .A(n3660), .B(n3661), .Z(n3513) );
  NOR U3603 ( .A(n3662), .B(n3663), .Z(n3661) );
  XNOR U3604 ( .A(n3660), .B(n3664), .Z(n3662) );
  XNOR U3605 ( .A(n3524), .B(n3514), .Z(n3626) );
  AND U3606 ( .A(n3385), .B(n3665), .Z(n3514) );
  XNOR U3607 ( .A(n3666), .B(n3531), .Z(n3524) );
  XOR U3608 ( .A(n3520), .B(n3519), .Z(n3531) );
  XNOR U3609 ( .A(n3667), .B(n3516), .Z(n3519) );
  XOR U3610 ( .A(n3668), .B(n3669), .Z(n3516) );
  AND U3611 ( .A(n3670), .B(n3671), .Z(n3669) );
  XOR U3612 ( .A(n3668), .B(n3672), .Z(n3670) );
  XNOR U3613 ( .A(n3673), .B(n3674), .Z(n3667) );
  NOR U3614 ( .A(n3675), .B(n3676), .Z(n3674) );
  XNOR U3615 ( .A(n3673), .B(n3677), .Z(n3675) );
  XOR U3616 ( .A(n3678), .B(n3679), .Z(n3520) );
  NOR U3617 ( .A(n3680), .B(n3681), .Z(n3679) );
  XNOR U3618 ( .A(n3678), .B(n3682), .Z(n3680) );
  XNOR U3619 ( .A(n3530), .B(n3521), .Z(n3666) );
  XOR U3620 ( .A(n3683), .B(n3684), .Z(n3521) );
  NOR U3621 ( .A(n3685), .B(n3686), .Z(n3684) );
  XNOR U3622 ( .A(n3683), .B(n3687), .Z(n3685) );
  XOR U3623 ( .A(n3688), .B(n3536), .Z(n3530) );
  XNOR U3624 ( .A(n3689), .B(n3690), .Z(n3536) );
  NOR U3625 ( .A(n3691), .B(n3692), .Z(n3690) );
  XNOR U3626 ( .A(n3689), .B(n3693), .Z(n3691) );
  XNOR U3627 ( .A(n3535), .B(n3527), .Z(n3688) );
  XOR U3628 ( .A(n3694), .B(n3695), .Z(n3527) );
  AND U3629 ( .A(n3696), .B(n3697), .Z(n3695) );
  XOR U3630 ( .A(n3694), .B(n3698), .Z(n3696) );
  XNOR U3631 ( .A(n3699), .B(n3532), .Z(n3535) );
  XOR U3632 ( .A(n3700), .B(n3701), .Z(n3532) );
  AND U3633 ( .A(n3702), .B(n3703), .Z(n3701) );
  XOR U3634 ( .A(n3700), .B(n3704), .Z(n3702) );
  XNOR U3635 ( .A(n3705), .B(n3706), .Z(n3699) );
  NOR U3636 ( .A(n3707), .B(n3708), .Z(n3706) );
  XOR U3637 ( .A(n3705), .B(n3709), .Z(n3707) );
  AND U3638 ( .A(n3385), .B(n3366), .Z(n3537) );
  XNOR U3639 ( .A(n3710), .B(n3586), .Z(n3366) );
  XOR U3640 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(
        p_input[256]), .Z(n3586) );
  XOR U3641 ( .A(n3563), .B(n3562), .Z(n3710) );
  XOR U3642 ( .A(n3711), .B(n3574), .Z(n3562) );
  XOR U3643 ( .A(n3548), .B(n3547), .Z(n3574) );
  XNOR U3644 ( .A(n3712), .B(n3553), .Z(n3547) );
  XNOR U3645 ( .A(n883), .B(p_input[280]), .Z(n3553) );
  IV U3646 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .Z(n883) );
  XOR U3647 ( .A(n3544), .B(n3552), .Z(n3712) );
  XOR U3648 ( .A(n3713), .B(n3549), .Z(n3552) );
  XNOR U3649 ( .A(n982), .B(p_input[278]), .Z(n3549) );
  IV U3650 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .Z(n982) );
  XOR U3651 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .B(n1937), 
        .Z(n3713) );
  XNOR U3652 ( .A(n1228), .B(p_input[274]), .Z(n3544) );
  IV U3653 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .Z(n1228) );
  XNOR U3654 ( .A(n3558), .B(n3557), .Z(n3548) );
  XOR U3655 ( .A(n3714), .B(n3554), .Z(n3557) );
  XNOR U3656 ( .A(n1179), .B(p_input[275]), .Z(n3554) );
  IV U3657 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .Z(n1179) );
  XOR U3658 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .B(n1939), 
        .Z(n3714) );
  XNOR U3659 ( .A(n1031), .B(p_input[277]), .Z(n3558) );
  IV U3660 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .Z(n1031) );
  XNOR U3661 ( .A(n3573), .B(n3559), .Z(n3711) );
  XNOR U3662 ( .A(n1130), .B(p_input[257]), .Z(n3559) );
  IV U3663 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n1130) );
  XNOR U3664 ( .A(n3715), .B(n3580), .Z(n3573) );
  XNOR U3665 ( .A(n3569), .B(n3568), .Z(n3580) );
  XOR U3666 ( .A(n3716), .B(n3565), .Z(n3568) );
  XNOR U3667 ( .A(n785), .B(p_input[282]), .Z(n3565) );
  IV U3668 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .Z(n785) );
  XOR U3669 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .B(n1943), 
        .Z(n3716) );
  XNOR U3670 ( .A(n686), .B(p_input[284]), .Z(n3569) );
  IV U3671 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .Z(n686) );
  XNOR U3672 ( .A(n3579), .B(n3570), .Z(n3715) );
  XNOR U3673 ( .A(n1277), .B(p_input[273]), .Z(n3570) );
  IV U3674 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .Z(n1277) );
  XOR U3675 ( .A(n3717), .B(n3585), .Z(n3579) );
  XNOR U3676 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .B(
        p_input[287]), .Z(n3585) );
  XOR U3677 ( .A(n3576), .B(n3584), .Z(n3717) );
  XOR U3678 ( .A(n3718), .B(n3581), .Z(n3584) );
  XNOR U3679 ( .A(n637), .B(p_input[285]), .Z(n3581) );
  IV U3680 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .Z(n637) );
  XOR U3681 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .B(n3074), 
        .Z(n3718) );
  XNOR U3682 ( .A(n834), .B(p_input[281]), .Z(n3576) );
  IV U3683 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .Z(n834) );
  XNOR U3684 ( .A(n3597), .B(n3596), .Z(n3563) );
  XNOR U3685 ( .A(n3719), .B(n3603), .Z(n3596) );
  XNOR U3686 ( .A(n3592), .B(n3591), .Z(n3603) );
  XOR U3687 ( .A(n3720), .B(n3588), .Z(n3591) );
  XNOR U3688 ( .A(n1574), .B(p_input[267]), .Z(n3588) );
  IV U3689 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n1574) );
  XOR U3690 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(n1949), 
        .Z(n3720) );
  XNOR U3691 ( .A(n1475), .B(p_input[269]), .Z(n3592) );
  IV U3692 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n1475) );
  XNOR U3693 ( .A(n3602), .B(n3593), .Z(n3719) );
  XNOR U3694 ( .A(n588), .B(p_input[258]), .Z(n3593) );
  IV U3695 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n588) );
  XOR U3696 ( .A(n3721), .B(n3608), .Z(n3602) );
  XNOR U3697 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .B(
        p_input[272]), .Z(n3608) );
  XOR U3698 ( .A(n3599), .B(n3607), .Z(n3721) );
  XOR U3699 ( .A(n3722), .B(n3604), .Z(n3607) );
  XNOR U3700 ( .A(n1426), .B(p_input[270]), .Z(n3604) );
  IV U3701 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n1426) );
  XOR U3702 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(n1953), 
        .Z(n3722) );
  XNOR U3703 ( .A(n1623), .B(p_input[266]), .Z(n3599) );
  IV U3704 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n1623) );
  XNOR U3705 ( .A(n3614), .B(n3613), .Z(n3597) );
  XNOR U3706 ( .A(n3723), .B(n3619), .Z(n3613) );
  XNOR U3707 ( .A(n120), .B(p_input[265]), .Z(n3619) );
  IV U3708 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .Z(n120) );
  XOR U3709 ( .A(n3610), .B(n3618), .Z(n3723) );
  XOR U3710 ( .A(n3724), .B(n3615), .Z(n3618) );
  XNOR U3711 ( .A(n226), .B(p_input[263]), .Z(n3615) );
  IV U3712 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .Z(n226) );
  XOR U3713 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .B(n3081), 
        .Z(n3724) );
  XNOR U3714 ( .A(n430), .B(p_input[259]), .Z(n3610) );
  IV U3715 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .Z(n430) );
  XNOR U3716 ( .A(n3624), .B(n3623), .Z(n3614) );
  XOR U3717 ( .A(n3725), .B(n3620), .Z(n3623) );
  XNOR U3718 ( .A(n379), .B(p_input[260]), .Z(n3620) );
  IV U3719 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .Z(n379) );
  XOR U3720 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(n3083), 
        .Z(n3725) );
  XNOR U3721 ( .A(n277), .B(p_input[262]), .Z(n3624) );
  IV U3722 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .Z(n277) );
  XOR U3723 ( .A(n3726), .B(n3687), .Z(n3385) );
  XNOR U3724 ( .A(n3637), .B(n3636), .Z(n3687) );
  XNOR U3725 ( .A(n3727), .B(n3643), .Z(n3636) );
  XNOR U3726 ( .A(n3632), .B(n3631), .Z(n3643) );
  XOR U3727 ( .A(n3728), .B(n3628), .Z(n3631) );
  XNOR U3728 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n2237), .Z(n3628) );
  IV U3729 ( .A(p_input[267]), .Z(n2237) );
  XOR U3730 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n1949), .Z(n3728) );
  IV U3731 ( .A(p_input[268]), .Z(n1949) );
  XOR U3732 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[269]), .Z(n3632)
         );
  XNOR U3733 ( .A(n3642), .B(n3633), .Z(n3727) );
  XOR U3734 ( .A(\knn_comb_/min_val_out[0][2] ), .B(p_input[258]), .Z(n3633)
         );
  XOR U3735 ( .A(n3729), .B(n3648), .Z(n3642) );
  XNOR U3736 ( .A(\knn_comb_/min_val_out[0][16] ), .B(p_input[272]), .Z(n3648)
         );
  XOR U3737 ( .A(n3639), .B(n3647), .Z(n3729) );
  XOR U3738 ( .A(n3730), .B(n3644), .Z(n3647) );
  XOR U3739 ( .A(\knn_comb_/min_val_out[0][14] ), .B(p_input[270]), .Z(n3644)
         );
  XOR U3740 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n1953), .Z(n3730) );
  IV U3741 ( .A(p_input[271]), .Z(n1953) );
  XNOR U3742 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n2240), .Z(n3639) );
  IV U3743 ( .A(p_input[266]), .Z(n2240) );
  XNOR U3744 ( .A(n3654), .B(n3653), .Z(n3637) );
  XNOR U3745 ( .A(n3731), .B(n3659), .Z(n3653) );
  XNOR U3746 ( .A(n126), .B(p_input[265]), .Z(n3659) );
  IV U3747 ( .A(\knn_comb_/min_val_out[0][9] ), .Z(n126) );
  XOR U3748 ( .A(n3650), .B(n3658), .Z(n3731) );
  XOR U3749 ( .A(n3732), .B(n3655), .Z(n3658) );
  XNOR U3750 ( .A(n230), .B(p_input[263]), .Z(n3655) );
  IV U3751 ( .A(\knn_comb_/min_val_out[0][7] ), .Z(n230) );
  XOR U3752 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n3081), .Z(n3732) );
  IV U3753 ( .A(p_input[264]), .Z(n3081) );
  XNOR U3754 ( .A(n434), .B(p_input[259]), .Z(n3650) );
  IV U3755 ( .A(\knn_comb_/min_val_out[0][3] ), .Z(n434) );
  XNOR U3756 ( .A(n3664), .B(n3663), .Z(n3654) );
  XOR U3757 ( .A(n3733), .B(n3660), .Z(n3663) );
  XNOR U3758 ( .A(n383), .B(p_input[260]), .Z(n3660) );
  IV U3759 ( .A(\knn_comb_/min_val_out[0][4] ), .Z(n383) );
  XOR U3760 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n3083), .Z(n3733) );
  IV U3761 ( .A(p_input[261]), .Z(n3083) );
  XNOR U3762 ( .A(n281), .B(p_input[262]), .Z(n3664) );
  IV U3763 ( .A(\knn_comb_/min_val_out[0][6] ), .Z(n281) );
  XOR U3764 ( .A(n3686), .B(n3665), .Z(n3726) );
  XOR U3765 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[256]), .Z(n3665)
         );
  XOR U3766 ( .A(n3734), .B(n3698), .Z(n3686) );
  XOR U3767 ( .A(n3672), .B(n3671), .Z(n3698) );
  XNOR U3768 ( .A(n3735), .B(n3677), .Z(n3671) );
  XOR U3769 ( .A(\knn_comb_/min_val_out[0][24] ), .B(p_input[280]), .Z(n3677)
         );
  XOR U3770 ( .A(n3668), .B(n3676), .Z(n3735) );
  XOR U3771 ( .A(n3736), .B(n3673), .Z(n3676) );
  XOR U3772 ( .A(\knn_comb_/min_val_out[0][22] ), .B(p_input[278]), .Z(n3673)
         );
  XOR U3773 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n1937), .Z(n3736) );
  IV U3774 ( .A(p_input[279]), .Z(n1937) );
  XNOR U3775 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n2225), .Z(n3668) );
  IV U3776 ( .A(p_input[274]), .Z(n2225) );
  XNOR U3777 ( .A(n3682), .B(n3681), .Z(n3672) );
  XOR U3778 ( .A(n3737), .B(n3678), .Z(n3681) );
  XOR U3779 ( .A(\knn_comb_/min_val_out[0][19] ), .B(p_input[275]), .Z(n3678)
         );
  XOR U3780 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n1939), .Z(n3737) );
  IV U3781 ( .A(p_input[276]), .Z(n1939) );
  XOR U3782 ( .A(\knn_comb_/min_val_out[0][21] ), .B(p_input[277]), .Z(n3682)
         );
  XNOR U3783 ( .A(n3697), .B(n3683), .Z(n3734) );
  XNOR U3784 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n2227), .Z(n3683) );
  IV U3785 ( .A(p_input[257]), .Z(n2227) );
  XNOR U3786 ( .A(n3738), .B(n3704), .Z(n3697) );
  XNOR U3787 ( .A(n3693), .B(n3692), .Z(n3704) );
  XOR U3788 ( .A(n3739), .B(n3689), .Z(n3692) );
  XNOR U3789 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n2230), .Z(n3689) );
  IV U3790 ( .A(p_input[282]), .Z(n2230) );
  XOR U3791 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n1943), .Z(n3739) );
  IV U3792 ( .A(p_input[283]), .Z(n1943) );
  XOR U3793 ( .A(\knn_comb_/min_val_out[0][28] ), .B(p_input[284]), .Z(n3693)
         );
  XNOR U3794 ( .A(n3703), .B(n3694), .Z(n3738) );
  XNOR U3795 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n2231), .Z(n3694) );
  IV U3796 ( .A(p_input[273]), .Z(n2231) );
  XOR U3797 ( .A(n3740), .B(n3709), .Z(n3703) );
  XNOR U3798 ( .A(\knn_comb_/min_val_out[0][31] ), .B(p_input[287]), .Z(n3709)
         );
  XOR U3799 ( .A(n3700), .B(n3708), .Z(n3740) );
  XOR U3800 ( .A(n3741), .B(n3705), .Z(n3708) );
  XOR U3801 ( .A(\knn_comb_/min_val_out[0][29] ), .B(p_input[285]), .Z(n3705)
         );
  XOR U3802 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n3074), .Z(n3741) );
  IV U3803 ( .A(p_input[286]), .Z(n3074) );
  XNOR U3804 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n2234), .Z(n3700) );
  IV U3805 ( .A(p_input[281]), .Z(n2234) );
endmodule

