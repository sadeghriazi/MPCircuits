
module knn_comb_BMR_W32_K3_N64 ( p_input, o );
  input [2079:0] p_input;
  output [95:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/min_val_out[0][16] , \knn_comb_/min_val_out[0][17] ,
         \knn_comb_/min_val_out[0][18] , \knn_comb_/min_val_out[0][19] ,
         \knn_comb_/min_val_out[0][20] , \knn_comb_/min_val_out[0][21] ,
         \knn_comb_/min_val_out[0][22] , \knn_comb_/min_val_out[0][23] ,
         \knn_comb_/min_val_out[0][24] , \knn_comb_/min_val_out[0][25] ,
         \knn_comb_/min_val_out[0][26] , \knn_comb_/min_val_out[0][27] ,
         \knn_comb_/min_val_out[0][28] , \knn_comb_/min_val_out[0][29] ,
         \knn_comb_/min_val_out[0][30] , \knn_comb_/min_val_out[0][31] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][16] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][17] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][18] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][19] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][20] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][21] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][22] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][23] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][24] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][25] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][26] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][27] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][28] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][29] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][30] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][31] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][31] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401, n18402, n18403,
         n18404, n18405, n18406, n18407, n18408, n18409, n18410, n18411,
         n18412, n18413, n18414, n18415, n18416, n18417, n18418, n18419,
         n18420, n18421, n18422, n18423, n18424, n18425, n18426, n18427,
         n18428, n18429, n18430, n18431, n18432, n18433, n18434, n18435,
         n18436, n18437, n18438, n18439, n18440, n18441, n18442, n18443,
         n18444, n18445, n18446, n18447, n18448, n18449, n18450, n18451,
         n18452, n18453, n18454, n18455, n18456, n18457, n18458, n18459,
         n18460, n18461, n18462, n18463, n18464, n18465, n18466, n18467,
         n18468, n18469, n18470, n18471, n18472, n18473, n18474, n18475,
         n18476, n18477, n18478, n18479, n18480, n18481, n18482, n18483,
         n18484, n18485, n18486, n18487, n18488, n18489, n18490, n18491,
         n18492, n18493, n18494, n18495, n18496, n18497, n18498, n18499,
         n18500, n18501, n18502, n18503, n18504, n18505, n18506, n18507,
         n18508, n18509, n18510, n18511, n18512, n18513, n18514, n18515,
         n18516, n18517, n18518, n18519, n18520, n18521, n18522, n18523,
         n18524, n18525, n18526, n18527, n18528, n18529, n18530, n18531,
         n18532, n18533, n18534, n18535, n18536, n18537, n18538, n18539,
         n18540, n18541, n18542, n18543, n18544, n18545, n18546, n18547,
         n18548, n18549, n18550, n18551, n18552, n18553, n18554, n18555,
         n18556, n18557, n18558, n18559, n18560, n18561, n18562, n18563,
         n18564, n18565, n18566, n18567, n18568, n18569, n18570, n18571,
         n18572, n18573, n18574, n18575, n18576, n18577, n18578, n18579,
         n18580, n18581, n18582, n18583, n18584, n18585, n18586, n18587,
         n18588, n18589, n18590, n18591, n18592, n18593, n18594, n18595,
         n18596, n18597, n18598, n18599, n18600, n18601, n18602, n18603,
         n18604, n18605, n18606, n18607, n18608, n18609, n18610, n18611,
         n18612, n18613, n18614, n18615, n18616, n18617, n18618, n18619,
         n18620, n18621, n18622, n18623, n18624, n18625, n18626, n18627,
         n18628, n18629, n18630, n18631, n18632, n18633, n18634, n18635,
         n18636, n18637, n18638, n18639, n18640, n18641, n18642, n18643,
         n18644, n18645, n18646, n18647, n18648, n18649, n18650, n18651,
         n18652, n18653, n18654, n18655, n18656, n18657, n18658, n18659,
         n18660, n18661, n18662, n18663, n18664, n18665, n18666, n18667,
         n18668, n18669, n18670, n18671, n18672, n18673, n18674, n18675,
         n18676, n18677, n18678, n18679, n18680, n18681, n18682, n18683,
         n18684, n18685, n18686, n18687, n18688, n18689, n18690, n18691,
         n18692, n18693, n18694, n18695, n18696, n18697, n18698, n18699,
         n18700, n18701, n18702, n18703, n18704, n18705, n18706, n18707,
         n18708, n18709, n18710, n18711, n18712, n18713, n18714, n18715,
         n18716, n18717, n18718, n18719, n18720, n18721, n18722, n18723,
         n18724, n18725, n18726, n18727, n18728, n18729, n18730, n18731,
         n18732, n18733, n18734, n18735, n18736, n18737, n18738, n18739,
         n18740, n18741, n18742, n18743, n18744, n18745, n18746, n18747,
         n18748, n18749, n18750, n18751, n18752, n18753, n18754, n18755,
         n18756, n18757, n18758, n18759, n18760, n18761, n18762, n18763,
         n18764, n18765, n18766, n18767, n18768, n18769, n18770, n18771,
         n18772, n18773, n18774, n18775, n18776, n18777, n18778, n18779,
         n18780, n18781, n18782, n18783, n18784, n18785, n18786, n18787,
         n18788, n18789, n18790, n18791, n18792, n18793, n18794, n18795,
         n18796, n18797, n18798, n18799, n18800, n18801, n18802, n18803,
         n18804, n18805, n18806, n18807, n18808, n18809, n18810, n18811,
         n18812, n18813, n18814, n18815, n18816, n18817, n18818, n18819,
         n18820, n18821, n18822, n18823, n18824, n18825, n18826, n18827,
         n18828, n18829, n18830, n18831, n18832, n18833, n18834, n18835,
         n18836, n18837, n18838, n18839, n18840, n18841, n18842, n18843,
         n18844, n18845, n18846, n18847, n18848, n18849, n18850, n18851,
         n18852, n18853, n18854, n18855, n18856, n18857, n18858, n18859,
         n18860, n18861, n18862, n18863, n18864, n18865, n18866, n18867,
         n18868, n18869, n18870, n18871, n18872, n18873, n18874, n18875,
         n18876, n18877, n18878, n18879, n18880, n18881, n18882, n18883,
         n18884, n18885, n18886, n18887, n18888, n18889, n18890, n18891,
         n18892, n18893, n18894, n18895, n18896, n18897, n18898, n18899,
         n18900, n18901, n18902, n18903, n18904, n18905, n18906, n18907,
         n18908, n18909, n18910, n18911, n18912, n18913, n18914, n18915,
         n18916, n18917, n18918, n18919, n18920, n18921, n18922, n18923,
         n18924, n18925, n18926, n18927, n18928, n18929, n18930, n18931,
         n18932, n18933, n18934, n18935, n18936, n18937, n18938, n18939,
         n18940, n18941, n18942, n18943, n18944, n18945, n18946, n18947,
         n18948, n18949, n18950, n18951, n18952, n18953, n18954, n18955,
         n18956, n18957, n18958, n18959, n18960, n18961, n18962, n18963,
         n18964, n18965, n18966, n18967, n18968, n18969, n18970, n18971,
         n18972, n18973, n18974, n18975, n18976, n18977, n18978, n18979,
         n18980, n18981, n18982, n18983, n18984, n18985, n18986, n18987,
         n18988, n18989, n18990, n18991, n18992, n18993, n18994, n18995,
         n18996, n18997, n18998, n18999, n19000, n19001, n19002, n19003,
         n19004, n19005, n19006, n19007, n19008, n19009, n19010, n19011,
         n19012, n19013, n19014, n19015, n19016, n19017, n19018, n19019,
         n19020, n19021, n19022, n19023, n19024, n19025, n19026, n19027,
         n19028, n19029, n19030, n19031, n19032, n19033, n19034, n19035,
         n19036, n19037, n19038, n19039, n19040, n19041, n19042, n19043,
         n19044, n19045, n19046, n19047, n19048, n19049, n19050, n19051,
         n19052, n19053, n19054, n19055, n19056, n19057, n19058, n19059,
         n19060, n19061, n19062, n19063, n19064, n19065, n19066, n19067,
         n19068, n19069, n19070, n19071, n19072, n19073, n19074, n19075,
         n19076, n19077, n19078, n19079, n19080, n19081, n19082, n19083,
         n19084, n19085, n19086, n19087, n19088, n19089, n19090, n19091,
         n19092, n19093, n19094, n19095, n19096, n19097, n19098, n19099,
         n19100, n19101, n19102, n19103, n19104, n19105, n19106, n19107,
         n19108, n19109, n19110, n19111, n19112, n19113, n19114, n19115,
         n19116, n19117, n19118, n19119, n19120, n19121, n19122, n19123,
         n19124, n19125, n19126, n19127, n19128, n19129, n19130, n19131,
         n19132, n19133, n19134, n19135, n19136, n19137, n19138, n19139,
         n19140, n19141, n19142, n19143, n19144, n19145, n19146, n19147,
         n19148, n19149, n19150, n19151, n19152, n19153, n19154, n19155,
         n19156, n19157, n19158, n19159, n19160, n19161, n19162, n19163,
         n19164, n19165, n19166, n19167, n19168, n19169, n19170, n19171,
         n19172, n19173, n19174, n19175, n19176, n19177, n19178, n19179,
         n19180, n19181, n19182, n19183, n19184, n19185, n19186, n19187,
         n19188, n19189, n19190, n19191, n19192, n19193, n19194, n19195,
         n19196, n19197, n19198, n19199, n19200, n19201, n19202, n19203,
         n19204, n19205, n19206, n19207, n19208, n19209, n19210, n19211,
         n19212, n19213, n19214, n19215, n19216, n19217, n19218, n19219,
         n19220, n19221, n19222, n19223, n19224, n19225, n19226, n19227,
         n19228, n19229, n19230, n19231, n19232, n19233, n19234, n19235,
         n19236, n19237, n19238, n19239, n19240, n19241, n19242, n19243,
         n19244, n19245, n19246, n19247, n19248, n19249, n19250, n19251,
         n19252, n19253, n19254, n19255, n19256, n19257, n19258, n19259,
         n19260, n19261, n19262, n19263, n19264, n19265, n19266, n19267,
         n19268, n19269, n19270, n19271, n19272, n19273, n19274, n19275,
         n19276, n19277, n19278, n19279, n19280, n19281, n19282, n19283,
         n19284, n19285, n19286, n19287, n19288, n19289, n19290, n19291,
         n19292, n19293, n19294, n19295, n19296, n19297, n19298, n19299,
         n19300, n19301, n19302, n19303, n19304, n19305, n19306, n19307,
         n19308, n19309, n19310, n19311, n19312, n19313, n19314, n19315,
         n19316, n19317, n19318, n19319, n19320, n19321, n19322, n19323,
         n19324, n19325, n19326, n19327, n19328, n19329, n19330, n19331,
         n19332, n19333, n19334, n19335, n19336, n19337, n19338, n19339,
         n19340, n19341, n19342, n19343, n19344, n19345, n19346, n19347,
         n19348, n19349, n19350, n19351, n19352, n19353, n19354, n19355,
         n19356, n19357, n19358, n19359, n19360, n19361, n19362, n19363,
         n19364, n19365, n19366, n19367, n19368, n19369, n19370, n19371,
         n19372, n19373, n19374, n19375, n19376, n19377, n19378, n19379,
         n19380, n19381, n19382, n19383, n19384, n19385, n19386, n19387,
         n19388, n19389, n19390, n19391, n19392, n19393, n19394, n19395,
         n19396, n19397, n19398, n19399, n19400, n19401, n19402, n19403,
         n19404, n19405, n19406, n19407, n19408, n19409, n19410, n19411,
         n19412, n19413, n19414, n19415, n19416, n19417, n19418, n19419,
         n19420, n19421, n19422, n19423, n19424, n19425, n19426, n19427,
         n19428, n19429, n19430, n19431, n19432, n19433, n19434, n19435,
         n19436, n19437, n19438, n19439, n19440, n19441, n19442, n19443,
         n19444, n19445, n19446, n19447, n19448, n19449, n19450, n19451,
         n19452, n19453, n19454, n19455, n19456, n19457, n19458, n19459,
         n19460, n19461, n19462, n19463, n19464, n19465, n19466, n19467,
         n19468, n19469, n19470, n19471, n19472, n19473, n19474, n19475,
         n19476, n19477, n19478, n19479, n19480, n19481, n19482, n19483,
         n19484, n19485, n19486, n19487, n19488, n19489, n19490, n19491,
         n19492, n19493, n19494, n19495, n19496, n19497, n19498, n19499,
         n19500, n19501, n19502, n19503, n19504, n19505, n19506, n19507,
         n19508, n19509, n19510, n19511, n19512, n19513, n19514, n19515,
         n19516, n19517, n19518, n19519, n19520, n19521, n19522, n19523,
         n19524, n19525, n19526, n19527, n19528, n19529, n19530, n19531,
         n19532, n19533, n19534, n19535, n19536, n19537, n19538, n19539,
         n19540, n19541, n19542, n19543, n19544, n19545, n19546, n19547,
         n19548, n19549, n19550, n19551, n19552, n19553, n19554, n19555,
         n19556, n19557, n19558, n19559, n19560, n19561, n19562, n19563,
         n19564, n19565, n19566, n19567, n19568, n19569, n19570, n19571,
         n19572, n19573, n19574, n19575, n19576, n19577, n19578, n19579,
         n19580, n19581, n19582, n19583, n19584, n19585, n19586, n19587,
         n19588, n19589, n19590, n19591, n19592, n19593, n19594, n19595,
         n19596, n19597, n19598, n19599, n19600, n19601, n19602, n19603,
         n19604, n19605, n19606, n19607, n19608, n19609, n19610, n19611,
         n19612, n19613, n19614, n19615, n19616, n19617, n19618, n19619,
         n19620, n19621, n19622, n19623, n19624, n19625, n19626, n19627,
         n19628, n19629, n19630, n19631, n19632, n19633, n19634, n19635,
         n19636, n19637, n19638, n19639, n19640, n19641, n19642, n19643,
         n19644, n19645, n19646, n19647, n19648, n19649, n19650, n19651,
         n19652, n19653, n19654, n19655, n19656, n19657, n19658, n19659,
         n19660, n19661, n19662, n19663, n19664, n19665, n19666, n19667,
         n19668, n19669, n19670, n19671, n19672, n19673, n19674, n19675,
         n19676, n19677, n19678, n19679, n19680, n19681, n19682, n19683,
         n19684, n19685, n19686, n19687, n19688, n19689, n19690, n19691,
         n19692, n19693, n19694, n19695, n19696, n19697, n19698, n19699,
         n19700, n19701, n19702, n19703, n19704, n19705, n19706, n19707,
         n19708, n19709, n19710, n19711, n19712, n19713, n19714, n19715,
         n19716, n19717, n19718, n19719, n19720, n19721, n19722, n19723,
         n19724, n19725, n19726, n19727, n19728, n19729, n19730, n19731,
         n19732, n19733, n19734, n19735, n19736, n19737, n19738, n19739,
         n19740, n19741, n19742, n19743, n19744, n19745, n19746, n19747,
         n19748, n19749, n19750, n19751, n19752, n19753, n19754, n19755,
         n19756, n19757, n19758, n19759, n19760, n19761, n19762, n19763,
         n19764, n19765, n19766, n19767, n19768, n19769, n19770, n19771,
         n19772, n19773, n19774, n19775, n19776, n19777, n19778, n19779,
         n19780, n19781, n19782, n19783, n19784, n19785, n19786, n19787,
         n19788, n19789, n19790, n19791, n19792, n19793, n19794, n19795,
         n19796, n19797, n19798, n19799, n19800, n19801, n19802, n19803,
         n19804, n19805, n19806, n19807, n19808, n19809, n19810, n19811,
         n19812, n19813, n19814, n19815, n19816, n19817, n19818, n19819,
         n19820, n19821, n19822, n19823, n19824, n19825, n19826, n19827,
         n19828, n19829, n19830, n19831, n19832, n19833, n19834, n19835,
         n19836, n19837, n19838, n19839, n19840, n19841, n19842, n19843,
         n19844, n19845, n19846, n19847, n19848, n19849, n19850, n19851,
         n19852, n19853, n19854, n19855, n19856, n19857, n19858, n19859,
         n19860, n19861, n19862, n19863, n19864, n19865, n19866, n19867,
         n19868, n19869, n19870, n19871, n19872, n19873, n19874, n19875,
         n19876, n19877, n19878, n19879, n19880, n19881, n19882, n19883,
         n19884, n19885, n19886, n19887, n19888, n19889, n19890, n19891,
         n19892, n19893, n19894, n19895, n19896, n19897, n19898, n19899,
         n19900, n19901, n19902, n19903, n19904, n19905, n19906, n19907,
         n19908, n19909, n19910, n19911, n19912, n19913, n19914, n19915,
         n19916, n19917, n19918, n19919, n19920, n19921, n19922, n19923,
         n19924, n19925, n19926, n19927, n19928, n19929, n19930, n19931,
         n19932, n19933, n19934, n19935, n19936, n19937, n19938, n19939,
         n19940, n19941, n19942, n19943, n19944, n19945, n19946, n19947,
         n19948, n19949, n19950, n19951, n19952, n19953, n19954, n19955,
         n19956, n19957, n19958, n19959, n19960, n19961, n19962, n19963,
         n19964, n19965, n19966, n19967, n19968, n19969, n19970, n19971,
         n19972, n19973, n19974, n19975, n19976, n19977, n19978, n19979,
         n19980, n19981, n19982, n19983, n19984, n19985, n19986, n19987,
         n19988, n19989, n19990, n19991, n19992, n19993, n19994, n19995,
         n19996, n19997, n19998, n19999, n20000, n20001, n20002, n20003,
         n20004, n20005, n20006, n20007, n20008, n20009, n20010, n20011,
         n20012, n20013, n20014, n20015, n20016, n20017, n20018, n20019,
         n20020, n20021, n20022, n20023, n20024, n20025, n20026, n20027,
         n20028, n20029, n20030, n20031, n20032, n20033, n20034, n20035,
         n20036, n20037, n20038, n20039, n20040, n20041, n20042, n20043,
         n20044, n20045, n20046, n20047, n20048, n20049, n20050, n20051,
         n20052, n20053, n20054, n20055, n20056, n20057, n20058, n20059,
         n20060, n20061, n20062, n20063, n20064, n20065, n20066, n20067,
         n20068, n20069, n20070, n20071, n20072, n20073, n20074, n20075,
         n20076, n20077, n20078, n20079, n20080, n20081, n20082, n20083,
         n20084, n20085, n20086, n20087, n20088, n20089, n20090, n20091,
         n20092, n20093, n20094, n20095, n20096, n20097, n20098, n20099,
         n20100, n20101, n20102, n20103, n20104, n20105, n20106, n20107,
         n20108, n20109, n20110, n20111, n20112, n20113, n20114, n20115,
         n20116, n20117, n20118, n20119, n20120, n20121, n20122, n20123,
         n20124, n20125, n20126, n20127, n20128, n20129, n20130, n20131,
         n20132, n20133, n20134, n20135, n20136, n20137, n20138, n20139,
         n20140, n20141, n20142, n20143, n20144, n20145, n20146, n20147,
         n20148, n20149, n20150, n20151, n20152, n20153, n20154, n20155,
         n20156, n20157, n20158, n20159, n20160, n20161, n20162, n20163,
         n20164, n20165, n20166, n20167, n20168, n20169, n20170, n20171,
         n20172, n20173, n20174, n20175, n20176, n20177, n20178, n20179,
         n20180, n20181, n20182, n20183, n20184, n20185, n20186, n20187,
         n20188, n20189, n20190, n20191, n20192, n20193, n20194, n20195,
         n20196, n20197, n20198, n20199, n20200, n20201, n20202, n20203,
         n20204, n20205, n20206, n20207, n20208, n20209, n20210, n20211,
         n20212, n20213, n20214, n20215, n20216, n20217, n20218, n20219,
         n20220, n20221, n20222, n20223, n20224, n20225, n20226, n20227,
         n20228, n20229, n20230, n20231, n20232, n20233, n20234, n20235,
         n20236, n20237, n20238, n20239, n20240, n20241, n20242, n20243,
         n20244, n20245, n20246, n20247, n20248, n20249, n20250, n20251,
         n20252, n20253, n20254, n20255, n20256, n20257, n20258, n20259,
         n20260, n20261, n20262, n20263, n20264, n20265, n20266, n20267,
         n20268, n20269, n20270, n20271, n20272, n20273, n20274, n20275,
         n20276, n20277, n20278, n20279, n20280, n20281, n20282, n20283,
         n20284, n20285, n20286, n20287, n20288, n20289, n20290, n20291,
         n20292, n20293, n20294, n20295, n20296, n20297, n20298, n20299,
         n20300, n20301, n20302, n20303, n20304, n20305, n20306, n20307,
         n20308, n20309, n20310, n20311, n20312, n20313, n20314, n20315,
         n20316, n20317, n20318, n20319, n20320, n20321, n20322, n20323,
         n20324, n20325, n20326, n20327, n20328, n20329, n20330, n20331,
         n20332, n20333, n20334, n20335, n20336, n20337, n20338, n20339,
         n20340, n20341, n20342, n20343, n20344, n20345, n20346, n20347,
         n20348, n20349, n20350, n20351, n20352, n20353, n20354, n20355,
         n20356, n20357, n20358, n20359, n20360, n20361, n20362, n20363,
         n20364, n20365, n20366, n20367, n20368, n20369, n20370, n20371,
         n20372, n20373, n20374, n20375, n20376, n20377, n20378, n20379,
         n20380, n20381, n20382, n20383, n20384, n20385, n20386, n20387,
         n20388, n20389, n20390, n20391, n20392, n20393, n20394, n20395,
         n20396, n20397, n20398, n20399, n20400, n20401, n20402, n20403,
         n20404, n20405, n20406, n20407, n20408, n20409, n20410, n20411,
         n20412, n20413, n20414, n20415, n20416, n20417, n20418, n20419,
         n20420, n20421, n20422, n20423, n20424, n20425, n20426, n20427,
         n20428, n20429, n20430, n20431, n20432, n20433, n20434, n20435,
         n20436, n20437, n20438, n20439, n20440, n20441, n20442, n20443,
         n20444, n20445, n20446, n20447, n20448, n20449, n20450, n20451,
         n20452, n20453, n20454, n20455, n20456, n20457, n20458, n20459,
         n20460, n20461, n20462, n20463, n20464, n20465, n20466, n20467,
         n20468, n20469, n20470, n20471, n20472, n20473, n20474, n20475,
         n20476, n20477, n20478, n20479, n20480, n20481, n20482, n20483,
         n20484, n20485, n20486, n20487, n20488, n20489, n20490, n20491,
         n20492, n20493, n20494, n20495, n20496, n20497, n20498, n20499,
         n20500, n20501, n20502, n20503, n20504, n20505, n20506, n20507,
         n20508, n20509, n20510, n20511, n20512, n20513, n20514, n20515,
         n20516, n20517, n20518, n20519, n20520, n20521, n20522, n20523,
         n20524, n20525, n20526, n20527, n20528, n20529, n20530, n20531,
         n20532, n20533, n20534, n20535, n20536, n20537, n20538, n20539,
         n20540, n20541, n20542, n20543, n20544, n20545, n20546, n20547,
         n20548, n20549, n20550, n20551, n20552, n20553, n20554, n20555,
         n20556, n20557, n20558, n20559, n20560, n20561, n20562, n20563,
         n20564, n20565, n20566, n20567, n20568, n20569, n20570, n20571,
         n20572, n20573, n20574, n20575, n20576, n20577, n20578, n20579,
         n20580, n20581, n20582, n20583, n20584, n20585, n20586, n20587,
         n20588, n20589, n20590, n20591, n20592, n20593, n20594, n20595,
         n20596, n20597, n20598, n20599, n20600, n20601, n20602, n20603,
         n20604, n20605, n20606, n20607, n20608, n20609, n20610, n20611,
         n20612, n20613, n20614, n20615, n20616, n20617, n20618, n20619,
         n20620, n20621, n20622, n20623, n20624, n20625, n20626, n20627,
         n20628, n20629, n20630, n20631, n20632, n20633, n20634, n20635,
         n20636, n20637, n20638, n20639, n20640, n20641, n20642, n20643,
         n20644, n20645, n20646, n20647, n20648, n20649, n20650, n20651,
         n20652, n20653, n20654, n20655, n20656, n20657, n20658, n20659,
         n20660, n20661, n20662, n20663, n20664, n20665, n20666, n20667,
         n20668, n20669, n20670, n20671, n20672, n20673, n20674, n20675,
         n20676, n20677, n20678, n20679, n20680, n20681, n20682, n20683,
         n20684, n20685, n20686, n20687, n20688, n20689, n20690, n20691,
         n20692, n20693, n20694, n20695, n20696, n20697, n20698, n20699,
         n20700, n20701, n20702, n20703, n20704, n20705, n20706, n20707,
         n20708, n20709, n20710, n20711, n20712, n20713, n20714, n20715,
         n20716, n20717, n20718, n20719, n20720, n20721, n20722, n20723,
         n20724, n20725, n20726, n20727, n20728, n20729, n20730, n20731,
         n20732, n20733, n20734, n20735, n20736, n20737, n20738, n20739,
         n20740, n20741, n20742, n20743, n20744, n20745, n20746, n20747,
         n20748, n20749, n20750, n20751, n20752, n20753, n20754, n20755,
         n20756, n20757, n20758, n20759, n20760, n20761, n20762, n20763,
         n20764, n20765, n20766, n20767, n20768, n20769, n20770, n20771,
         n20772, n20773, n20774, n20775, n20776, n20777, n20778, n20779,
         n20780, n20781, n20782, n20783, n20784, n20785, n20786, n20787,
         n20788, n20789, n20790, n20791, n20792, n20793, n20794, n20795,
         n20796, n20797, n20798, n20799, n20800, n20801, n20802, n20803,
         n20804, n20805, n20806, n20807, n20808, n20809, n20810, n20811,
         n20812, n20813, n20814, n20815, n20816, n20817, n20818, n20819,
         n20820, n20821, n20822, n20823, n20824, n20825, n20826, n20827,
         n20828, n20829, n20830, n20831, n20832, n20833, n20834, n20835,
         n20836, n20837, n20838, n20839, n20840, n20841, n20842, n20843,
         n20844, n20845, n20846, n20847, n20848, n20849, n20850, n20851,
         n20852, n20853, n20854, n20855, n20856, n20857, n20858, n20859,
         n20860, n20861, n20862, n20863, n20864, n20865, n20866, n20867,
         n20868, n20869, n20870, n20871, n20872, n20873, n20874, n20875,
         n20876, n20877, n20878, n20879, n20880, n20881, n20882, n20883,
         n20884, n20885, n20886, n20887, n20888, n20889, n20890, n20891,
         n20892, n20893, n20894, n20895, n20896, n20897, n20898, n20899,
         n20900, n20901, n20902, n20903, n20904, n20905, n20906, n20907,
         n20908, n20909, n20910, n20911, n20912, n20913, n20914, n20915,
         n20916, n20917, n20918, n20919, n20920, n20921, n20922, n20923,
         n20924, n20925, n20926, n20927, n20928, n20929, n20930, n20931,
         n20932, n20933, n20934, n20935, n20936, n20937, n20938, n20939,
         n20940, n20941, n20942, n20943, n20944, n20945, n20946, n20947,
         n20948, n20949, n20950, n20951, n20952, n20953, n20954, n20955,
         n20956, n20957, n20958, n20959, n20960, n20961, n20962, n20963,
         n20964, n20965, n20966, n20967, n20968, n20969, n20970, n20971,
         n20972, n20973, n20974, n20975, n20976, n20977, n20978, n20979,
         n20980, n20981, n20982, n20983, n20984, n20985, n20986, n20987,
         n20988, n20989, n20990, n20991, n20992, n20993, n20994, n20995,
         n20996, n20997, n20998, n20999, n21000, n21001, n21002, n21003,
         n21004, n21005, n21006, n21007, n21008, n21009, n21010, n21011,
         n21012, n21013, n21014, n21015, n21016, n21017, n21018, n21019,
         n21020, n21021, n21022, n21023, n21024, n21025, n21026, n21027,
         n21028, n21029, n21030, n21031, n21032, n21033, n21034, n21035,
         n21036, n21037, n21038, n21039, n21040, n21041, n21042, n21043,
         n21044, n21045, n21046, n21047, n21048, n21049, n21050, n21051,
         n21052, n21053, n21054, n21055, n21056, n21057, n21058, n21059,
         n21060, n21061, n21062, n21063, n21064, n21065, n21066, n21067,
         n21068, n21069, n21070, n21071, n21072, n21073, n21074, n21075,
         n21076, n21077, n21078, n21079, n21080, n21081, n21082, n21083,
         n21084, n21085, n21086, n21087, n21088, n21089, n21090, n21091,
         n21092, n21093, n21094, n21095, n21096, n21097, n21098, n21099,
         n21100, n21101, n21102, n21103, n21104, n21105, n21106, n21107,
         n21108, n21109, n21110, n21111, n21112, n21113, n21114, n21115,
         n21116, n21117, n21118, n21119, n21120, n21121, n21122, n21123,
         n21124, n21125, n21126, n21127, n21128, n21129, n21130, n21131,
         n21132, n21133, n21134, n21135, n21136, n21137, n21138, n21139,
         n21140, n21141, n21142, n21143, n21144, n21145, n21146, n21147,
         n21148, n21149, n21150, n21151, n21152, n21153, n21154, n21155,
         n21156, n21157, n21158, n21159, n21160, n21161, n21162, n21163,
         n21164, n21165, n21166, n21167, n21168, n21169, n21170, n21171,
         n21172, n21173, n21174, n21175, n21176, n21177, n21178, n21179,
         n21180, n21181, n21182, n21183, n21184, n21185, n21186, n21187,
         n21188, n21189, n21190, n21191, n21192, n21193, n21194, n21195,
         n21196, n21197, n21198, n21199, n21200, n21201, n21202, n21203,
         n21204, n21205, n21206, n21207, n21208, n21209, n21210, n21211,
         n21212, n21213, n21214, n21215, n21216, n21217, n21218, n21219,
         n21220, n21221, n21222, n21223, n21224, n21225, n21226, n21227,
         n21228, n21229, n21230, n21231, n21232, n21233, n21234, n21235,
         n21236, n21237, n21238, n21239, n21240, n21241, n21242, n21243,
         n21244, n21245, n21246, n21247, n21248, n21249, n21250, n21251,
         n21252, n21253, n21254, n21255, n21256, n21257, n21258, n21259,
         n21260, n21261, n21262, n21263, n21264, n21265, n21266, n21267,
         n21268, n21269, n21270, n21271, n21272, n21273, n21274, n21275,
         n21276, n21277, n21278, n21279, n21280, n21281, n21282, n21283,
         n21284, n21285, n21286, n21287, n21288, n21289, n21290, n21291,
         n21292, n21293, n21294, n21295, n21296, n21297, n21298, n21299,
         n21300, n21301, n21302, n21303, n21304, n21305, n21306, n21307,
         n21308, n21309, n21310, n21311, n21312, n21313, n21314, n21315,
         n21316, n21317, n21318, n21319, n21320, n21321, n21322, n21323,
         n21324, n21325, n21326, n21327, n21328, n21329, n21330, n21331,
         n21332, n21333, n21334, n21335, n21336, n21337, n21338, n21339,
         n21340, n21341, n21342, n21343, n21344, n21345, n21346, n21347,
         n21348, n21349, n21350, n21351, n21352, n21353, n21354, n21355,
         n21356, n21357, n21358, n21359, n21360, n21361, n21362, n21363,
         n21364, n21365, n21366, n21367, n21368, n21369, n21370, n21371,
         n21372, n21373, n21374, n21375, n21376, n21377, n21378, n21379,
         n21380, n21381, n21382, n21383, n21384, n21385, n21386, n21387,
         n21388, n21389, n21390, n21391, n21392, n21393, n21394, n21395,
         n21396, n21397, n21398, n21399, n21400, n21401, n21402, n21403,
         n21404, n21405, n21406, n21407, n21408, n21409, n21410, n21411,
         n21412, n21413, n21414, n21415, n21416, n21417, n21418, n21419,
         n21420, n21421, n21422, n21423, n21424, n21425, n21426, n21427,
         n21428, n21429, n21430, n21431, n21432, n21433, n21434, n21435,
         n21436, n21437, n21438, n21439, n21440, n21441, n21442, n21443,
         n21444, n21445, n21446, n21447, n21448, n21449, n21450, n21451,
         n21452, n21453, n21454, n21455, n21456, n21457, n21458, n21459,
         n21460, n21461, n21462, n21463, n21464, n21465, n21466, n21467,
         n21468, n21469, n21470, n21471, n21472, n21473, n21474, n21475,
         n21476, n21477, n21478, n21479, n21480, n21481, n21482, n21483,
         n21484, n21485, n21486, n21487, n21488, n21489, n21490, n21491,
         n21492, n21493, n21494, n21495, n21496, n21497, n21498, n21499,
         n21500, n21501, n21502, n21503, n21504, n21505, n21506, n21507,
         n21508, n21509, n21510, n21511, n21512, n21513, n21514, n21515,
         n21516, n21517, n21518, n21519, n21520, n21521, n21522, n21523,
         n21524, n21525, n21526, n21527, n21528, n21529, n21530, n21531,
         n21532, n21533, n21534, n21535, n21536, n21537, n21538, n21539,
         n21540, n21541, n21542, n21543, n21544, n21545, n21546, n21547,
         n21548, n21549, n21550, n21551, n21552, n21553, n21554, n21555,
         n21556, n21557, n21558, n21559, n21560, n21561, n21562, n21563,
         n21564, n21565, n21566, n21567, n21568, n21569, n21570, n21571,
         n21572, n21573, n21574, n21575, n21576, n21577, n21578, n21579,
         n21580, n21581, n21582, n21583, n21584, n21585, n21586, n21587,
         n21588, n21589, n21590, n21591, n21592, n21593, n21594, n21595,
         n21596, n21597, n21598, n21599, n21600, n21601, n21602, n21603,
         n21604, n21605, n21606, n21607, n21608, n21609, n21610, n21611,
         n21612, n21613, n21614, n21615, n21616, n21617, n21618, n21619,
         n21620, n21621, n21622, n21623, n21624, n21625, n21626, n21627,
         n21628, n21629, n21630, n21631, n21632, n21633, n21634, n21635,
         n21636, n21637, n21638, n21639, n21640, n21641, n21642, n21643,
         n21644, n21645, n21646, n21647, n21648, n21649, n21650, n21651,
         n21652, n21653, n21654, n21655, n21656, n21657, n21658, n21659,
         n21660, n21661, n21662, n21663, n21664, n21665, n21666, n21667,
         n21668, n21669, n21670, n21671, n21672, n21673, n21674, n21675,
         n21676, n21677, n21678, n21679, n21680, n21681, n21682, n21683,
         n21684, n21685, n21686, n21687, n21688, n21689, n21690, n21691,
         n21692, n21693, n21694, n21695, n21696, n21697, n21698, n21699,
         n21700, n21701, n21702, n21703, n21704, n21705, n21706, n21707,
         n21708, n21709, n21710, n21711, n21712, n21713, n21714, n21715,
         n21716, n21717, n21718, n21719, n21720, n21721, n21722, n21723,
         n21724, n21725, n21726, n21727, n21728, n21729, n21730, n21731,
         n21732, n21733, n21734, n21735, n21736, n21737, n21738, n21739,
         n21740, n21741, n21742, n21743, n21744, n21745, n21746, n21747,
         n21748, n21749, n21750, n21751, n21752, n21753, n21754, n21755,
         n21756, n21757, n21758, n21759, n21760, n21761, n21762, n21763,
         n21764, n21765, n21766, n21767, n21768, n21769, n21770, n21771,
         n21772, n21773, n21774, n21775, n21776, n21777, n21778, n21779,
         n21780, n21781, n21782, n21783, n21784, n21785, n21786, n21787,
         n21788, n21789, n21790, n21791, n21792, n21793, n21794, n21795,
         n21796, n21797, n21798, n21799, n21800, n21801, n21802, n21803,
         n21804, n21805, n21806, n21807, n21808, n21809, n21810, n21811,
         n21812, n21813, n21814, n21815, n21816, n21817, n21818, n21819,
         n21820, n21821, n21822, n21823, n21824, n21825, n21826, n21827,
         n21828, n21829, n21830, n21831, n21832, n21833, n21834, n21835,
         n21836, n21837, n21838, n21839, n21840, n21841, n21842, n21843,
         n21844, n21845, n21846, n21847, n21848, n21849, n21850, n21851,
         n21852, n21853, n21854, n21855, n21856, n21857, n21858, n21859,
         n21860, n21861, n21862, n21863, n21864, n21865, n21866, n21867,
         n21868, n21869, n21870, n21871, n21872, n21873, n21874, n21875,
         n21876, n21877, n21878, n21879, n21880, n21881, n21882, n21883,
         n21884, n21885, n21886, n21887, n21888, n21889, n21890, n21891,
         n21892, n21893, n21894, n21895, n21896, n21897, n21898, n21899,
         n21900, n21901, n21902, n21903, n21904, n21905, n21906, n21907,
         n21908, n21909, n21910, n21911, n21912, n21913, n21914, n21915,
         n21916, n21917, n21918, n21919, n21920, n21921, n21922, n21923,
         n21924, n21925, n21926, n21927, n21928, n21929, n21930, n21931,
         n21932, n21933, n21934, n21935, n21936, n21937, n21938, n21939,
         n21940, n21941, n21942, n21943, n21944, n21945, n21946, n21947,
         n21948, n21949, n21950, n21951, n21952, n21953, n21954, n21955,
         n21956, n21957, n21958, n21959, n21960, n21961, n21962, n21963,
         n21964, n21965, n21966, n21967, n21968, n21969, n21970, n21971,
         n21972, n21973, n21974, n21975, n21976, n21977, n21978, n21979,
         n21980, n21981, n21982, n21983, n21984, n21985, n21986, n21987,
         n21988, n21989, n21990, n21991, n21992, n21993, n21994, n21995,
         n21996, n21997, n21998, n21999, n22000, n22001, n22002, n22003,
         n22004, n22005, n22006, n22007, n22008, n22009, n22010, n22011,
         n22012, n22013, n22014, n22015, n22016, n22017, n22018, n22019,
         n22020, n22021, n22022, n22023, n22024, n22025, n22026, n22027,
         n22028, n22029, n22030, n22031, n22032, n22033, n22034, n22035,
         n22036, n22037, n22038, n22039, n22040, n22041, n22042, n22043,
         n22044, n22045, n22046, n22047, n22048, n22049, n22050, n22051,
         n22052, n22053, n22054, n22055, n22056, n22057, n22058, n22059,
         n22060, n22061, n22062, n22063, n22064, n22065, n22066, n22067,
         n22068, n22069, n22070, n22071, n22072, n22073, n22074, n22075,
         n22076, n22077, n22078, n22079, n22080, n22081, n22082, n22083,
         n22084, n22085, n22086, n22087, n22088, n22089, n22090, n22091,
         n22092, n22093, n22094, n22095, n22096, n22097, n22098, n22099,
         n22100, n22101, n22102, n22103, n22104, n22105, n22106, n22107,
         n22108, n22109, n22110, n22111, n22112, n22113, n22114, n22115,
         n22116, n22117, n22118, n22119, n22120, n22121, n22122, n22123,
         n22124, n22125, n22126, n22127, n22128, n22129, n22130, n22131,
         n22132, n22133, n22134, n22135, n22136, n22137, n22138, n22139,
         n22140, n22141, n22142, n22143, n22144, n22145, n22146, n22147,
         n22148, n22149, n22150, n22151, n22152, n22153, n22154, n22155,
         n22156, n22157, n22158, n22159, n22160, n22161, n22162, n22163,
         n22164, n22165, n22166, n22167, n22168, n22169, n22170, n22171,
         n22172, n22173, n22174, n22175, n22176, n22177, n22178, n22179,
         n22180, n22181, n22182, n22183, n22184, n22185, n22186, n22187,
         n22188, n22189, n22190, n22191, n22192, n22193, n22194, n22195,
         n22196, n22197, n22198, n22199, n22200, n22201, n22202, n22203,
         n22204, n22205, n22206, n22207, n22208, n22209, n22210, n22211,
         n22212, n22213, n22214, n22215, n22216, n22217, n22218, n22219,
         n22220, n22221, n22222, n22223, n22224, n22225, n22226, n22227,
         n22228, n22229, n22230, n22231, n22232, n22233, n22234, n22235,
         n22236, n22237, n22238, n22239, n22240, n22241, n22242, n22243,
         n22244, n22245, n22246, n22247, n22248, n22249, n22250, n22251,
         n22252, n22253, n22254, n22255, n22256, n22257, n22258, n22259,
         n22260, n22261, n22262, n22263, n22264, n22265, n22266, n22267,
         n22268, n22269, n22270, n22271, n22272, n22273, n22274, n22275,
         n22276, n22277, n22278, n22279, n22280, n22281, n22282, n22283,
         n22284, n22285, n22286, n22287, n22288, n22289, n22290, n22291,
         n22292, n22293, n22294, n22295, n22296, n22297, n22298, n22299,
         n22300, n22301, n22302, n22303, n22304, n22305, n22306, n22307,
         n22308, n22309, n22310, n22311, n22312, n22313, n22314, n22315,
         n22316, n22317, n22318, n22319, n22320, n22321, n22322, n22323,
         n22324, n22325, n22326, n22327, n22328, n22329, n22330, n22331,
         n22332, n22333, n22334, n22335, n22336, n22337, n22338, n22339,
         n22340, n22341, n22342, n22343, n22344, n22345, n22346, n22347,
         n22348, n22349, n22350, n22351, n22352, n22353, n22354, n22355,
         n22356, n22357, n22358, n22359, n22360, n22361, n22362, n22363,
         n22364, n22365, n22366, n22367, n22368, n22369, n22370, n22371,
         n22372, n22373, n22374, n22375, n22376, n22377, n22378, n22379,
         n22380, n22381, n22382, n22383, n22384, n22385, n22386, n22387,
         n22388, n22389, n22390, n22391, n22392, n22393, n22394, n22395,
         n22396, n22397, n22398, n22399, n22400, n22401, n22402, n22403,
         n22404, n22405, n22406, n22407, n22408, n22409, n22410, n22411,
         n22412, n22413, n22414, n22415, n22416, n22417, n22418, n22419,
         n22420, n22421, n22422, n22423, n22424, n22425, n22426, n22427,
         n22428, n22429, n22430, n22431, n22432, n22433, n22434, n22435,
         n22436, n22437, n22438, n22439, n22440, n22441, n22442, n22443,
         n22444, n22445, n22446, n22447, n22448, n22449, n22450, n22451,
         n22452, n22453, n22454, n22455, n22456, n22457, n22458, n22459,
         n22460, n22461, n22462, n22463, n22464, n22465, n22466, n22467,
         n22468, n22469, n22470, n22471, n22472, n22473, n22474, n22475,
         n22476, n22477, n22478, n22479, n22480, n22481, n22482, n22483,
         n22484, n22485, n22486, n22487, n22488, n22489, n22490, n22491,
         n22492, n22493, n22494, n22495, n22496, n22497, n22498, n22499,
         n22500, n22501, n22502, n22503, n22504, n22505, n22506, n22507,
         n22508, n22509, n22510, n22511, n22512, n22513, n22514, n22515,
         n22516, n22517, n22518, n22519, n22520, n22521, n22522, n22523,
         n22524, n22525, n22526, n22527, n22528, n22529, n22530, n22531,
         n22532, n22533, n22534, n22535, n22536, n22537, n22538, n22539,
         n22540, n22541, n22542, n22543, n22544, n22545, n22546, n22547,
         n22548, n22549, n22550, n22551, n22552, n22553, n22554, n22555,
         n22556, n22557, n22558, n22559, n22560, n22561, n22562, n22563,
         n22564, n22565, n22566, n22567, n22568, n22569, n22570, n22571,
         n22572, n22573, n22574, n22575, n22576, n22577, n22578, n22579,
         n22580, n22581, n22582, n22583, n22584, n22585, n22586, n22587,
         n22588, n22589, n22590, n22591, n22592, n22593, n22594, n22595,
         n22596, n22597, n22598, n22599, n22600, n22601, n22602, n22603,
         n22604, n22605, n22606, n22607, n22608, n22609, n22610, n22611,
         n22612, n22613, n22614, n22615, n22616, n22617, n22618, n22619,
         n22620, n22621, n22622, n22623, n22624, n22625, n22626, n22627,
         n22628, n22629, n22630, n22631, n22632, n22633, n22634, n22635,
         n22636, n22637, n22638, n22639, n22640, n22641, n22642, n22643,
         n22644, n22645, n22646, n22647, n22648, n22649, n22650, n22651,
         n22652, n22653, n22654, n22655, n22656, n22657, n22658, n22659,
         n22660, n22661, n22662, n22663, n22664, n22665, n22666, n22667,
         n22668, n22669, n22670, n22671, n22672, n22673, n22674, n22675,
         n22676, n22677, n22678, n22679, n22680, n22681, n22682, n22683,
         n22684, n22685, n22686, n22687, n22688, n22689, n22690, n22691,
         n22692, n22693, n22694, n22695, n22696, n22697, n22698, n22699,
         n22700, n22701, n22702, n22703, n22704, n22705, n22706, n22707,
         n22708, n22709, n22710, n22711, n22712, n22713, n22714, n22715,
         n22716, n22717, n22718, n22719, n22720, n22721, n22722, n22723,
         n22724, n22725, n22726, n22727, n22728, n22729, n22730, n22731,
         n22732, n22733, n22734, n22735, n22736, n22737, n22738, n22739,
         n22740, n22741, n22742, n22743, n22744, n22745, n22746, n22747,
         n22748, n22749, n22750, n22751, n22752, n22753, n22754, n22755,
         n22756, n22757, n22758, n22759, n22760, n22761, n22762, n22763,
         n22764, n22765, n22766, n22767, n22768, n22769, n22770, n22771,
         n22772, n22773, n22774, n22775, n22776, n22777, n22778, n22779,
         n22780, n22781, n22782, n22783, n22784, n22785, n22786, n22787,
         n22788, n22789, n22790, n22791, n22792, n22793, n22794, n22795,
         n22796, n22797, n22798, n22799, n22800, n22801, n22802, n22803,
         n22804, n22805, n22806, n22807, n22808, n22809, n22810, n22811,
         n22812, n22813, n22814, n22815, n22816, n22817, n22818, n22819,
         n22820, n22821, n22822, n22823, n22824, n22825, n22826, n22827,
         n22828, n22829, n22830, n22831, n22832, n22833, n22834, n22835,
         n22836, n22837, n22838, n22839, n22840, n22841, n22842, n22843,
         n22844, n22845, n22846, n22847, n22848, n22849, n22850, n22851,
         n22852, n22853, n22854, n22855, n22856, n22857, n22858, n22859,
         n22860, n22861, n22862, n22863, n22864, n22865, n22866, n22867,
         n22868, n22869, n22870, n22871, n22872, n22873, n22874, n22875,
         n22876, n22877, n22878, n22879, n22880, n22881, n22882, n22883,
         n22884, n22885, n22886, n22887, n22888, n22889, n22890, n22891,
         n22892, n22893, n22894, n22895, n22896, n22897, n22898, n22899,
         n22900, n22901, n22902, n22903, n22904, n22905, n22906, n22907,
         n22908, n22909, n22910, n22911, n22912, n22913, n22914, n22915,
         n22916, n22917, n22918, n22919, n22920, n22921, n22922, n22923,
         n22924, n22925, n22926, n22927, n22928, n22929, n22930, n22931,
         n22932, n22933, n22934, n22935, n22936, n22937, n22938, n22939,
         n22940, n22941, n22942, n22943, n22944, n22945, n22946, n22947,
         n22948, n22949, n22950, n22951, n22952, n22953, n22954, n22955,
         n22956, n22957, n22958, n22959, n22960, n22961, n22962, n22963,
         n22964, n22965, n22966, n22967, n22968, n22969, n22970, n22971,
         n22972, n22973, n22974, n22975, n22976, n22977, n22978, n22979,
         n22980, n22981, n22982, n22983, n22984, n22985, n22986, n22987,
         n22988, n22989, n22990, n22991, n22992, n22993, n22994, n22995,
         n22996, n22997, n22998, n22999, n23000, n23001, n23002, n23003,
         n23004, n23005, n23006, n23007, n23008, n23009, n23010, n23011,
         n23012, n23013, n23014, n23015, n23016, n23017, n23018, n23019,
         n23020, n23021, n23022, n23023, n23024, n23025, n23026, n23027,
         n23028, n23029, n23030, n23031, n23032, n23033, n23034, n23035,
         n23036, n23037, n23038, n23039, n23040, n23041, n23042, n23043,
         n23044, n23045, n23046, n23047, n23048, n23049, n23050, n23051,
         n23052, n23053, n23054, n23055, n23056, n23057, n23058, n23059,
         n23060, n23061, n23062, n23063, n23064, n23065, n23066, n23067,
         n23068, n23069, n23070, n23071, n23072, n23073, n23074, n23075,
         n23076, n23077, n23078, n23079, n23080, n23081, n23082, n23083,
         n23084, n23085, n23086, n23087, n23088, n23089, n23090, n23091,
         n23092, n23093, n23094, n23095, n23096, n23097, n23098, n23099,
         n23100, n23101, n23102, n23103, n23104, n23105, n23106, n23107,
         n23108, n23109, n23110, n23111, n23112, n23113, n23114, n23115,
         n23116, n23117, n23118, n23119, n23120, n23121, n23122, n23123,
         n23124, n23125, n23126, n23127, n23128, n23129, n23130, n23131,
         n23132, n23133, n23134, n23135, n23136, n23137, n23138, n23139,
         n23140, n23141, n23142, n23143, n23144, n23145, n23146, n23147,
         n23148, n23149, n23150, n23151, n23152, n23153, n23154, n23155,
         n23156, n23157, n23158, n23159, n23160, n23161, n23162, n23163,
         n23164, n23165, n23166, n23167, n23168, n23169, n23170, n23171,
         n23172, n23173, n23174, n23175, n23176, n23177, n23178, n23179,
         n23180, n23181, n23182, n23183, n23184, n23185, n23186, n23187,
         n23188, n23189, n23190, n23191, n23192, n23193, n23194, n23195,
         n23196, n23197, n23198, n23199, n23200, n23201, n23202, n23203,
         n23204, n23205, n23206, n23207, n23208, n23209, n23210, n23211,
         n23212, n23213, n23214, n23215, n23216, n23217, n23218, n23219,
         n23220, n23221, n23222, n23223, n23224, n23225, n23226, n23227,
         n23228, n23229, n23230, n23231, n23232, n23233, n23234, n23235,
         n23236, n23237, n23238, n23239, n23240, n23241, n23242, n23243,
         n23244, n23245, n23246, n23247, n23248, n23249, n23250, n23251,
         n23252, n23253, n23254, n23255, n23256, n23257, n23258, n23259,
         n23260, n23261, n23262, n23263, n23264, n23265, n23266, n23267,
         n23268, n23269, n23270, n23271, n23272, n23273, n23274, n23275,
         n23276, n23277, n23278, n23279, n23280, n23281, n23282, n23283,
         n23284, n23285, n23286, n23287, n23288, n23289, n23290, n23291,
         n23292, n23293, n23294, n23295, n23296, n23297, n23298, n23299,
         n23300, n23301, n23302, n23303, n23304, n23305, n23306, n23307,
         n23308, n23309, n23310, n23311, n23312, n23313, n23314, n23315,
         n23316, n23317, n23318, n23319, n23320, n23321, n23322, n23323,
         n23324, n23325, n23326, n23327, n23328, n23329, n23330, n23331,
         n23332, n23333, n23334, n23335, n23336, n23337, n23338, n23339,
         n23340, n23341, n23342, n23343, n23344, n23345, n23346, n23347,
         n23348, n23349, n23350, n23351, n23352, n23353, n23354, n23355,
         n23356, n23357, n23358, n23359, n23360, n23361, n23362, n23363,
         n23364, n23365, n23366, n23367, n23368, n23369, n23370, n23371,
         n23372, n23373, n23374, n23375, n23376, n23377, n23378, n23379,
         n23380, n23381, n23382, n23383, n23384, n23385, n23386, n23387,
         n23388, n23389, n23390, n23391, n23392, n23393, n23394, n23395,
         n23396, n23397, n23398, n23399, n23400, n23401, n23402, n23403,
         n23404, n23405, n23406, n23407, n23408, n23409, n23410, n23411,
         n23412, n23413, n23414, n23415, n23416, n23417, n23418, n23419,
         n23420, n23421, n23422, n23423, n23424, n23425, n23426, n23427,
         n23428, n23429, n23430, n23431, n23432, n23433, n23434, n23435,
         n23436, n23437, n23438, n23439, n23440, n23441, n23442, n23443,
         n23444, n23445, n23446, n23447, n23448, n23449, n23450, n23451,
         n23452, n23453, n23454, n23455, n23456, n23457, n23458, n23459,
         n23460, n23461, n23462, n23463, n23464, n23465, n23466, n23467,
         n23468, n23469, n23470, n23471, n23472, n23473, n23474, n23475,
         n23476, n23477, n23478, n23479, n23480, n23481, n23482, n23483,
         n23484, n23485, n23486, n23487, n23488, n23489, n23490, n23491,
         n23492, n23493, n23494, n23495, n23496, n23497, n23498, n23499,
         n23500, n23501, n23502, n23503, n23504, n23505, n23506, n23507,
         n23508, n23509, n23510, n23511, n23512, n23513, n23514, n23515,
         n23516, n23517, n23518, n23519, n23520, n23521, n23522, n23523,
         n23524, n23525, n23526, n23527, n23528, n23529, n23530, n23531,
         n23532, n23533, n23534, n23535, n23536, n23537, n23538, n23539,
         n23540, n23541, n23542, n23543, n23544, n23545, n23546, n23547,
         n23548, n23549, n23550, n23551, n23552, n23553, n23554, n23555,
         n23556, n23557, n23558, n23559, n23560, n23561, n23562, n23563,
         n23564, n23565, n23566, n23567, n23568, n23569, n23570, n23571,
         n23572, n23573, n23574, n23575, n23576, n23577, n23578, n23579,
         n23580, n23581, n23582, n23583, n23584, n23585, n23586, n23587,
         n23588, n23589, n23590, n23591, n23592, n23593, n23594, n23595,
         n23596, n23597, n23598, n23599, n23600, n23601, n23602, n23603,
         n23604, n23605, n23606, n23607, n23608, n23609, n23610, n23611,
         n23612, n23613, n23614, n23615, n23616, n23617, n23618, n23619,
         n23620, n23621, n23622, n23623, n23624, n23625, n23626, n23627,
         n23628, n23629, n23630, n23631, n23632, n23633, n23634, n23635,
         n23636, n23637, n23638, n23639, n23640, n23641, n23642, n23643,
         n23644, n23645, n23646, n23647, n23648, n23649, n23650, n23651,
         n23652, n23653, n23654, n23655, n23656, n23657, n23658, n23659,
         n23660, n23661, n23662, n23663, n23664, n23665, n23666, n23667,
         n23668, n23669, n23670, n23671, n23672, n23673, n23674, n23675,
         n23676, n23677, n23678, n23679, n23680, n23681, n23682, n23683,
         n23684, n23685, n23686, n23687, n23688, n23689, n23690, n23691,
         n23692, n23693, n23694, n23695, n23696, n23697, n23698, n23699,
         n23700, n23701, n23702, n23703, n23704, n23705, n23706, n23707,
         n23708, n23709, n23710, n23711, n23712, n23713, n23714, n23715,
         n23716, n23717, n23718, n23719, n23720, n23721, n23722, n23723,
         n23724, n23725, n23726, n23727, n23728, n23729, n23730, n23731,
         n23732, n23733, n23734, n23735, n23736, n23737, n23738, n23739,
         n23740, n23741, n23742, n23743, n23744, n23745, n23746, n23747,
         n23748, n23749, n23750, n23751, n23752, n23753, n23754, n23755,
         n23756, n23757, n23758, n23759, n23760, n23761, n23762, n23763,
         n23764, n23765, n23766, n23767, n23768, n23769, n23770, n23771,
         n23772, n23773, n23774, n23775, n23776, n23777, n23778, n23779,
         n23780, n23781, n23782, n23783, n23784, n23785, n23786, n23787,
         n23788, n23789, n23790, n23791, n23792, n23793, n23794, n23795,
         n23796, n23797, n23798, n23799, n23800, n23801, n23802, n23803,
         n23804, n23805, n23806, n23807, n23808, n23809, n23810, n23811,
         n23812, n23813, n23814, n23815, n23816, n23817, n23818, n23819,
         n23820, n23821, n23822, n23823, n23824, n23825, n23826, n23827,
         n23828, n23829, n23830, n23831, n23832, n23833, n23834, n23835,
         n23836, n23837, n23838, n23839, n23840, n23841, n23842, n23843,
         n23844, n23845, n23846, n23847, n23848, n23849, n23850, n23851,
         n23852, n23853, n23854, n23855, n23856, n23857, n23858, n23859,
         n23860, n23861, n23862, n23863, n23864, n23865, n23866, n23867,
         n23868, n23869, n23870, n23871, n23872, n23873, n23874, n23875,
         n23876, n23877, n23878, n23879, n23880, n23881, n23882, n23883,
         n23884, n23885, n23886, n23887, n23888, n23889, n23890, n23891,
         n23892, n23893, n23894, n23895, n23896, n23897, n23898, n23899,
         n23900, n23901, n23902, n23903, n23904, n23905, n23906, n23907,
         n23908, n23909, n23910, n23911, n23912, n23913, n23914, n23915,
         n23916, n23917, n23918, n23919, n23920, n23921, n23922, n23923,
         n23924, n23925, n23926, n23927, n23928, n23929, n23930, n23931,
         n23932, n23933, n23934, n23935, n23936, n23937, n23938, n23939,
         n23940, n23941, n23942, n23943, n23944, n23945, n23946, n23947,
         n23948, n23949, n23950, n23951, n23952, n23953, n23954, n23955,
         n23956, n23957, n23958, n23959, n23960, n23961, n23962, n23963,
         n23964, n23965, n23966, n23967, n23968, n23969, n23970, n23971,
         n23972, n23973, n23974, n23975, n23976, n23977, n23978, n23979,
         n23980, n23981, n23982, n23983, n23984, n23985, n23986, n23987,
         n23988, n23989, n23990, n23991, n23992, n23993, n23994, n23995,
         n23996, n23997, n23998, n23999, n24000, n24001, n24002, n24003,
         n24004, n24005, n24006, n24007, n24008, n24009, n24010, n24011,
         n24012, n24013, n24014, n24015, n24016, n24017, n24018, n24019,
         n24020, n24021, n24022, n24023, n24024, n24025, n24026, n24027,
         n24028, n24029, n24030, n24031, n24032, n24033, n24034, n24035,
         n24036, n24037, n24038, n24039, n24040, n24041, n24042, n24043,
         n24044, n24045, n24046, n24047, n24048, n24049, n24050, n24051,
         n24052, n24053, n24054, n24055, n24056, n24057, n24058, n24059,
         n24060, n24061, n24062, n24063, n24064, n24065, n24066, n24067,
         n24068, n24069, n24070, n24071, n24072, n24073, n24074, n24075,
         n24076, n24077, n24078, n24079, n24080, n24081, n24082, n24083,
         n24084, n24085, n24086, n24087, n24088, n24089, n24090, n24091,
         n24092, n24093, n24094, n24095, n24096, n24097, n24098, n24099,
         n24100, n24101, n24102, n24103, n24104, n24105, n24106, n24107,
         n24108, n24109, n24110, n24111, n24112, n24113, n24114, n24115,
         n24116, n24117, n24118, n24119, n24120, n24121, n24122, n24123,
         n24124, n24125, n24126, n24127, n24128, n24129, n24130, n24131,
         n24132, n24133, n24134, n24135, n24136, n24137, n24138, n24139,
         n24140, n24141, n24142, n24143, n24144, n24145, n24146, n24147,
         n24148, n24149, n24150, n24151, n24152, n24153, n24154, n24155,
         n24156, n24157, n24158, n24159, n24160, n24161, n24162, n24163,
         n24164, n24165, n24166, n24167, n24168, n24169, n24170, n24171,
         n24172, n24173, n24174, n24175, n24176, n24177, n24178, n24179,
         n24180, n24181, n24182, n24183, n24184, n24185, n24186, n24187,
         n24188, n24189, n24190, n24191, n24192, n24193, n24194, n24195,
         n24196, n24197, n24198, n24199, n24200, n24201, n24202, n24203,
         n24204, n24205, n24206, n24207, n24208, n24209, n24210, n24211,
         n24212, n24213, n24214, n24215, n24216, n24217, n24218, n24219,
         n24220, n24221, n24222, n24223, n24224, n24225, n24226, n24227,
         n24228, n24229, n24230, n24231, n24232, n24233, n24234, n24235,
         n24236, n24237, n24238, n24239, n24240, n24241, n24242, n24243,
         n24244, n24245, n24246, n24247, n24248, n24249, n24250, n24251,
         n24252, n24253, n24254, n24255, n24256, n24257, n24258, n24259,
         n24260, n24261, n24262, n24263, n24264, n24265, n24266, n24267,
         n24268, n24269, n24270, n24271, n24272, n24273, n24274, n24275,
         n24276, n24277, n24278, n24279, n24280, n24281, n24282, n24283,
         n24284, n24285, n24286, n24287, n24288, n24289, n24290, n24291,
         n24292, n24293, n24294, n24295, n24296, n24297, n24298, n24299,
         n24300, n24301, n24302, n24303, n24304, n24305, n24306, n24307,
         n24308, n24309, n24310, n24311, n24312, n24313, n24314, n24315,
         n24316, n24317, n24318, n24319, n24320, n24321, n24322, n24323,
         n24324, n24325, n24326, n24327, n24328, n24329, n24330, n24331,
         n24332, n24333, n24334, n24335, n24336, n24337, n24338, n24339,
         n24340, n24341, n24342, n24343, n24344, n24345, n24346, n24347,
         n24348, n24349, n24350, n24351, n24352, n24353, n24354, n24355,
         n24356, n24357, n24358, n24359, n24360, n24361, n24362, n24363,
         n24364, n24365, n24366, n24367, n24368, n24369, n24370, n24371,
         n24372, n24373, n24374, n24375, n24376, n24377, n24378, n24379,
         n24380, n24381, n24382, n24383, n24384, n24385, n24386, n24387,
         n24388, n24389, n24390, n24391, n24392, n24393, n24394, n24395,
         n24396, n24397, n24398, n24399, n24400, n24401, n24402, n24403,
         n24404, n24405, n24406, n24407, n24408, n24409, n24410, n24411,
         n24412, n24413, n24414, n24415, n24416, n24417, n24418, n24419,
         n24420, n24421, n24422, n24423, n24424, n24425, n24426, n24427,
         n24428, n24429, n24430, n24431, n24432, n24433, n24434, n24435,
         n24436, n24437, n24438, n24439, n24440, n24441, n24442, n24443,
         n24444, n24445, n24446, n24447, n24448, n24449, n24450, n24451,
         n24452, n24453, n24454, n24455, n24456, n24457, n24458, n24459,
         n24460, n24461, n24462, n24463, n24464, n24465, n24466, n24467,
         n24468, n24469, n24470, n24471, n24472, n24473, n24474, n24475,
         n24476, n24477, n24478, n24479, n24480, n24481, n24482, n24483,
         n24484, n24485, n24486, n24487, n24488, n24489, n24490, n24491,
         n24492, n24493, n24494, n24495, n24496, n24497, n24498, n24499,
         n24500, n24501, n24502, n24503, n24504, n24505, n24506, n24507,
         n24508, n24509, n24510, n24511, n24512, n24513, n24514, n24515,
         n24516, n24517, n24518, n24519, n24520, n24521, n24522, n24523,
         n24524, n24525, n24526, n24527, n24528, n24529, n24530, n24531,
         n24532, n24533, n24534, n24535, n24536, n24537, n24538, n24539,
         n24540, n24541, n24542, n24543, n24544, n24545, n24546, n24547,
         n24548, n24549, n24550, n24551, n24552, n24553, n24554, n24555,
         n24556, n24557, n24558, n24559, n24560, n24561, n24562, n24563,
         n24564, n24565, n24566, n24567, n24568, n24569, n24570, n24571,
         n24572, n24573, n24574, n24575, n24576, n24577, n24578, n24579,
         n24580, n24581, n24582, n24583, n24584, n24585, n24586, n24587,
         n24588, n24589, n24590, n24591, n24592, n24593, n24594, n24595,
         n24596, n24597, n24598, n24599, n24600, n24601, n24602, n24603,
         n24604, n24605, n24606, n24607, n24608, n24609, n24610, n24611,
         n24612, n24613, n24614, n24615, n24616, n24617, n24618, n24619,
         n24620, n24621, n24622, n24623, n24624, n24625, n24626, n24627,
         n24628, n24629, n24630, n24631, n24632, n24633, n24634, n24635,
         n24636, n24637, n24638, n24639, n24640, n24641, n24642, n24643,
         n24644, n24645, n24646, n24647, n24648, n24649, n24650, n24651,
         n24652, n24653, n24654, n24655, n24656, n24657, n24658, n24659,
         n24660, n24661, n24662, n24663, n24664, n24665, n24666, n24667,
         n24668, n24669, n24670, n24671, n24672, n24673, n24674, n24675,
         n24676, n24677, n24678, n24679, n24680, n24681, n24682, n24683,
         n24684, n24685, n24686, n24687, n24688, n24689, n24690, n24691,
         n24692, n24693, n24694, n24695, n24696, n24697, n24698, n24699,
         n24700, n24701, n24702, n24703, n24704, n24705, n24706, n24707,
         n24708, n24709, n24710, n24711, n24712, n24713, n24714, n24715,
         n24716, n24717, n24718, n24719, n24720, n24721, n24722, n24723,
         n24724, n24725, n24726, n24727, n24728, n24729, n24730, n24731,
         n24732, n24733, n24734, n24735, n24736, n24737, n24738, n24739,
         n24740, n24741, n24742, n24743, n24744, n24745, n24746, n24747,
         n24748, n24749, n24750, n24751, n24752, n24753, n24754, n24755,
         n24756, n24757, n24758, n24759, n24760, n24761, n24762, n24763,
         n24764, n24765, n24766, n24767, n24768, n24769, n24770, n24771,
         n24772, n24773, n24774, n24775, n24776, n24777, n24778, n24779,
         n24780, n24781, n24782, n24783, n24784, n24785, n24786, n24787,
         n24788, n24789, n24790, n24791, n24792, n24793, n24794, n24795,
         n24796, n24797, n24798, n24799, n24800, n24801, n24802, n24803,
         n24804, n24805, n24806, n24807, n24808, n24809, n24810, n24811,
         n24812, n24813, n24814, n24815, n24816, n24817, n24818, n24819,
         n24820, n24821, n24822, n24823, n24824, n24825, n24826, n24827,
         n24828, n24829, n24830, n24831, n24832, n24833, n24834, n24835,
         n24836, n24837, n24838, n24839, n24840, n24841, n24842, n24843,
         n24844, n24845, n24846, n24847, n24848, n24849, n24850, n24851,
         n24852, n24853, n24854, n24855, n24856, n24857, n24858, n24859,
         n24860, n24861, n24862, n24863, n24864, n24865, n24866, n24867,
         n24868, n24869, n24870, n24871, n24872, n24873, n24874, n24875,
         n24876, n24877, n24878, n24879, n24880, n24881, n24882, n24883,
         n24884, n24885, n24886, n24887, n24888, n24889, n24890, n24891,
         n24892, n24893, n24894, n24895, n24896, n24897, n24898, n24899,
         n24900, n24901, n24902, n24903, n24904, n24905, n24906, n24907,
         n24908, n24909, n24910, n24911, n24912, n24913, n24914, n24915,
         n24916, n24917, n24918, n24919, n24920, n24921, n24922, n24923,
         n24924, n24925, n24926, n24927, n24928, n24929, n24930, n24931,
         n24932, n24933, n24934, n24935, n24936, n24937, n24938, n24939,
         n24940, n24941, n24942, n24943, n24944, n24945, n24946, n24947,
         n24948, n24949, n24950, n24951, n24952, n24953, n24954, n24955,
         n24956, n24957, n24958, n24959, n24960, n24961, n24962, n24963,
         n24964, n24965, n24966, n24967, n24968, n24969, n24970, n24971,
         n24972, n24973, n24974, n24975, n24976, n24977, n24978, n24979,
         n24980, n24981, n24982, n24983, n24984, n24985, n24986, n24987,
         n24988, n24989, n24990, n24991, n24992, n24993, n24994, n24995,
         n24996, n24997, n24998, n24999, n25000, n25001, n25002, n25003,
         n25004, n25005, n25006, n25007, n25008, n25009, n25010, n25011,
         n25012, n25013, n25014, n25015, n25016, n25017, n25018, n25019,
         n25020, n25021, n25022, n25023, n25024, n25025, n25026, n25027,
         n25028, n25029, n25030, n25031, n25032, n25033, n25034, n25035,
         n25036, n25037, n25038, n25039, n25040, n25041, n25042, n25043,
         n25044, n25045, n25046, n25047, n25048, n25049, n25050, n25051,
         n25052, n25053, n25054, n25055, n25056, n25057, n25058, n25059,
         n25060, n25061, n25062, n25063, n25064, n25065, n25066, n25067,
         n25068, n25069, n25070, n25071, n25072, n25073, n25074, n25075,
         n25076, n25077, n25078, n25079, n25080, n25081, n25082, n25083,
         n25084, n25085, n25086, n25087, n25088, n25089, n25090, n25091,
         n25092, n25093, n25094, n25095, n25096, n25097, n25098, n25099,
         n25100, n25101, n25102, n25103, n25104, n25105, n25106, n25107,
         n25108, n25109, n25110, n25111, n25112, n25113, n25114, n25115,
         n25116, n25117, n25118, n25119, n25120, n25121, n25122, n25123,
         n25124, n25125, n25126, n25127, n25128, n25129, n25130, n25131,
         n25132, n25133, n25134, n25135, n25136, n25137, n25138, n25139,
         n25140, n25141, n25142, n25143, n25144, n25145, n25146, n25147,
         n25148, n25149, n25150, n25151, n25152, n25153, n25154, n25155,
         n25156, n25157, n25158, n25159, n25160, n25161, n25162, n25163,
         n25164, n25165, n25166, n25167, n25168, n25169, n25170, n25171,
         n25172, n25173, n25174, n25175, n25176, n25177, n25178, n25179,
         n25180, n25181, n25182, n25183, n25184, n25185, n25186, n25187,
         n25188, n25189, n25190, n25191, n25192, n25193, n25194, n25195,
         n25196, n25197, n25198, n25199, n25200, n25201, n25202, n25203,
         n25204, n25205, n25206, n25207, n25208, n25209, n25210, n25211,
         n25212, n25213, n25214, n25215, n25216, n25217, n25218, n25219,
         n25220, n25221, n25222, n25223, n25224, n25225, n25226, n25227,
         n25228, n25229, n25230, n25231, n25232, n25233, n25234, n25235,
         n25236, n25237, n25238, n25239, n25240, n25241, n25242, n25243,
         n25244, n25245, n25246, n25247, n25248, n25249, n25250, n25251,
         n25252, n25253, n25254, n25255, n25256, n25257, n25258, n25259,
         n25260, n25261, n25262, n25263, n25264, n25265, n25266, n25267,
         n25268, n25269, n25270, n25271, n25272, n25273, n25274, n25275,
         n25276, n25277, n25278, n25279, n25280, n25281, n25282, n25283,
         n25284, n25285, n25286, n25287, n25288, n25289, n25290, n25291,
         n25292, n25293, n25294, n25295, n25296, n25297, n25298, n25299,
         n25300, n25301, n25302, n25303, n25304, n25305, n25306, n25307,
         n25308, n25309, n25310, n25311, n25312, n25313, n25314, n25315,
         n25316, n25317, n25318, n25319, n25320, n25321, n25322, n25323,
         n25324, n25325, n25326, n25327, n25328, n25329, n25330, n25331,
         n25332, n25333, n25334, n25335, n25336, n25337, n25338, n25339,
         n25340, n25341, n25342, n25343, n25344, n25345, n25346, n25347,
         n25348, n25349, n25350, n25351, n25352, n25353, n25354, n25355,
         n25356, n25357, n25358, n25359, n25360, n25361, n25362, n25363,
         n25364, n25365, n25366, n25367, n25368, n25369, n25370, n25371,
         n25372, n25373, n25374, n25375, n25376, n25377, n25378, n25379,
         n25380, n25381, n25382, n25383, n25384, n25385, n25386, n25387,
         n25388, n25389, n25390, n25391, n25392, n25393, n25394, n25395,
         n25396, n25397, n25398, n25399, n25400, n25401, n25402, n25403,
         n25404, n25405, n25406, n25407, n25408, n25409, n25410, n25411,
         n25412, n25413, n25414, n25415, n25416, n25417, n25418, n25419,
         n25420, n25421, n25422, n25423, n25424, n25425, n25426, n25427,
         n25428, n25429, n25430, n25431, n25432, n25433, n25434, n25435,
         n25436, n25437, n25438, n25439, n25440, n25441, n25442, n25443,
         n25444, n25445, n25446, n25447, n25448, n25449, n25450, n25451,
         n25452, n25453, n25454, n25455, n25456, n25457, n25458, n25459,
         n25460, n25461, n25462, n25463, n25464, n25465, n25466, n25467,
         n25468, n25469, n25470, n25471, n25472, n25473, n25474, n25475,
         n25476, n25477, n25478, n25479, n25480, n25481, n25482, n25483,
         n25484, n25485, n25486, n25487, n25488, n25489, n25490, n25491,
         n25492, n25493, n25494, n25495, n25496, n25497, n25498, n25499,
         n25500, n25501, n25502, n25503, n25504, n25505, n25506, n25507,
         n25508, n25509, n25510, n25511, n25512, n25513, n25514, n25515,
         n25516, n25517, n25518, n25519, n25520, n25521, n25522, n25523,
         n25524, n25525, n25526, n25527, n25528, n25529, n25530, n25531,
         n25532, n25533, n25534, n25535, n25536, n25537, n25538, n25539,
         n25540, n25541, n25542, n25543, n25544, n25545, n25546, n25547,
         n25548, n25549, n25550, n25551, n25552, n25553, n25554, n25555,
         n25556, n25557, n25558, n25559, n25560, n25561, n25562, n25563,
         n25564, n25565, n25566, n25567, n25568, n25569, n25570, n25571,
         n25572, n25573, n25574, n25575, n25576, n25577, n25578, n25579,
         n25580, n25581, n25582, n25583, n25584, n25585, n25586, n25587,
         n25588, n25589, n25590, n25591, n25592, n25593, n25594, n25595,
         n25596, n25597, n25598, n25599, n25600, n25601, n25602, n25603,
         n25604, n25605, n25606, n25607, n25608, n25609, n25610, n25611,
         n25612, n25613, n25614, n25615, n25616, n25617, n25618, n25619,
         n25620, n25621, n25622, n25623, n25624, n25625, n25626, n25627,
         n25628, n25629, n25630, n25631, n25632, n25633, n25634, n25635,
         n25636, n25637, n25638, n25639, n25640, n25641, n25642, n25643,
         n25644, n25645, n25646, n25647, n25648, n25649, n25650, n25651,
         n25652, n25653, n25654, n25655, n25656, n25657, n25658, n25659,
         n25660, n25661, n25662, n25663, n25664, n25665, n25666, n25667,
         n25668, n25669, n25670, n25671, n25672, n25673, n25674, n25675,
         n25676, n25677, n25678, n25679, n25680, n25681, n25682, n25683,
         n25684, n25685, n25686, n25687, n25688, n25689, n25690, n25691,
         n25692, n25693, n25694, n25695, n25696, n25697, n25698, n25699,
         n25700, n25701, n25702, n25703, n25704, n25705, n25706, n25707,
         n25708, n25709, n25710, n25711, n25712, n25713, n25714, n25715,
         n25716, n25717, n25718, n25719, n25720, n25721, n25722, n25723,
         n25724, n25725, n25726, n25727, n25728, n25729, n25730, n25731,
         n25732, n25733, n25734, n25735, n25736, n25737, n25738, n25739,
         n25740, n25741, n25742, n25743, n25744, n25745, n25746, n25747,
         n25748, n25749, n25750, n25751, n25752, n25753, n25754, n25755,
         n25756, n25757, n25758, n25759, n25760, n25761, n25762, n25763,
         n25764, n25765, n25766, n25767, n25768, n25769, n25770, n25771,
         n25772, n25773, n25774, n25775, n25776, n25777, n25778, n25779,
         n25780, n25781, n25782, n25783, n25784, n25785, n25786, n25787,
         n25788, n25789, n25790, n25791, n25792, n25793, n25794, n25795,
         n25796, n25797, n25798, n25799, n25800, n25801, n25802, n25803,
         n25804, n25805, n25806, n25807, n25808, n25809, n25810, n25811,
         n25812, n25813, n25814, n25815, n25816, n25817, n25818, n25819,
         n25820, n25821, n25822, n25823, n25824, n25825, n25826, n25827,
         n25828, n25829, n25830, n25831, n25832, n25833, n25834, n25835,
         n25836, n25837, n25838, n25839, n25840, n25841, n25842, n25843,
         n25844, n25845, n25846, n25847, n25848, n25849, n25850, n25851,
         n25852, n25853, n25854, n25855, n25856, n25857, n25858, n25859,
         n25860, n25861, n25862, n25863, n25864, n25865, n25866, n25867,
         n25868, n25869, n25870, n25871, n25872, n25873, n25874, n25875,
         n25876, n25877, n25878, n25879, n25880, n25881, n25882, n25883,
         n25884, n25885, n25886, n25887, n25888, n25889, n25890, n25891,
         n25892, n25893, n25894, n25895, n25896, n25897, n25898, n25899,
         n25900, n25901, n25902, n25903, n25904, n25905, n25906, n25907,
         n25908, n25909, n25910, n25911, n25912, n25913, n25914, n25915,
         n25916, n25917, n25918, n25919, n25920, n25921, n25922, n25923,
         n25924, n25925, n25926, n25927, n25928, n25929, n25930, n25931,
         n25932, n25933, n25934, n25935, n25936, n25937, n25938, n25939,
         n25940, n25941, n25942, n25943, n25944, n25945, n25946, n25947,
         n25948, n25949, n25950, n25951, n25952, n25953, n25954, n25955,
         n25956, n25957, n25958, n25959, n25960, n25961, n25962, n25963,
         n25964, n25965, n25966, n25967, n25968, n25969, n25970, n25971,
         n25972, n25973, n25974, n25975, n25976, n25977, n25978, n25979,
         n25980, n25981, n25982, n25983, n25984, n25985, n25986, n25987,
         n25988, n25989, n25990, n25991, n25992, n25993, n25994, n25995,
         n25996, n25997, n25998, n25999, n26000, n26001, n26002, n26003,
         n26004, n26005, n26006, n26007, n26008, n26009, n26010, n26011,
         n26012, n26013, n26014, n26015, n26016, n26017, n26018, n26019,
         n26020, n26021, n26022, n26023, n26024, n26025, n26026, n26027,
         n26028, n26029, n26030, n26031, n26032, n26033, n26034, n26035,
         n26036, n26037, n26038, n26039, n26040, n26041, n26042, n26043,
         n26044, n26045, n26046, n26047, n26048, n26049, n26050, n26051,
         n26052, n26053, n26054, n26055, n26056, n26057, n26058, n26059,
         n26060, n26061, n26062, n26063, n26064, n26065, n26066, n26067,
         n26068, n26069, n26070, n26071, n26072, n26073, n26074, n26075,
         n26076, n26077, n26078, n26079, n26080, n26081, n26082, n26083,
         n26084, n26085, n26086, n26087, n26088, n26089, n26090, n26091,
         n26092, n26093, n26094, n26095, n26096, n26097, n26098, n26099,
         n26100, n26101, n26102, n26103, n26104, n26105, n26106, n26107,
         n26108, n26109, n26110, n26111, n26112, n26113, n26114, n26115,
         n26116, n26117, n26118, n26119, n26120, n26121, n26122, n26123,
         n26124, n26125, n26126, n26127, n26128, n26129, n26130, n26131,
         n26132, n26133, n26134, n26135, n26136, n26137, n26138, n26139,
         n26140, n26141, n26142, n26143, n26144, n26145, n26146, n26147,
         n26148, n26149, n26150, n26151, n26152, n26153, n26154, n26155,
         n26156, n26157, n26158, n26159, n26160, n26161, n26162, n26163,
         n26164, n26165, n26166, n26167, n26168, n26169, n26170, n26171,
         n26172, n26173, n26174, n26175, n26176, n26177, n26178, n26179,
         n26180, n26181, n26182, n26183, n26184, n26185, n26186, n26187,
         n26188, n26189, n26190, n26191, n26192, n26193, n26194, n26195,
         n26196, n26197, n26198, n26199, n26200, n26201, n26202, n26203,
         n26204, n26205, n26206, n26207, n26208, n26209, n26210, n26211,
         n26212, n26213, n26214, n26215, n26216, n26217, n26218, n26219,
         n26220, n26221, n26222, n26223, n26224, n26225, n26226, n26227,
         n26228, n26229, n26230, n26231, n26232, n26233, n26234, n26235,
         n26236, n26237, n26238, n26239, n26240, n26241, n26242, n26243,
         n26244, n26245, n26246, n26247, n26248, n26249, n26250, n26251,
         n26252, n26253, n26254, n26255, n26256, n26257, n26258, n26259,
         n26260, n26261, n26262, n26263, n26264, n26265, n26266, n26267,
         n26268, n26269, n26270, n26271, n26272, n26273, n26274, n26275,
         n26276, n26277, n26278, n26279, n26280, n26281, n26282, n26283,
         n26284, n26285, n26286, n26287, n26288, n26289, n26290, n26291,
         n26292, n26293, n26294, n26295, n26296, n26297, n26298, n26299,
         n26300, n26301, n26302, n26303, n26304, n26305, n26306, n26307,
         n26308, n26309, n26310, n26311, n26312, n26313, n26314, n26315,
         n26316, n26317, n26318, n26319, n26320, n26321, n26322, n26323,
         n26324, n26325, n26326, n26327, n26328, n26329, n26330, n26331,
         n26332, n26333, n26334, n26335, n26336, n26337, n26338, n26339,
         n26340, n26341, n26342, n26343, n26344, n26345, n26346, n26347,
         n26348, n26349, n26350, n26351, n26352, n26353, n26354, n26355,
         n26356, n26357, n26358, n26359, n26360, n26361, n26362, n26363,
         n26364, n26365, n26366, n26367, n26368, n26369, n26370, n26371,
         n26372, n26373, n26374, n26375, n26376, n26377, n26378, n26379,
         n26380, n26381, n26382, n26383, n26384, n26385, n26386, n26387,
         n26388, n26389, n26390, n26391, n26392, n26393, n26394, n26395,
         n26396, n26397, n26398, n26399, n26400, n26401, n26402, n26403,
         n26404, n26405, n26406, n26407, n26408, n26409, n26410, n26411,
         n26412, n26413, n26414, n26415, n26416, n26417, n26418, n26419,
         n26420, n26421, n26422, n26423, n26424, n26425, n26426, n26427,
         n26428, n26429, n26430, n26431, n26432, n26433, n26434, n26435,
         n26436, n26437, n26438, n26439, n26440, n26441, n26442, n26443,
         n26444, n26445, n26446, n26447, n26448, n26449, n26450, n26451,
         n26452, n26453, n26454, n26455, n26456, n26457, n26458, n26459,
         n26460, n26461, n26462, n26463, n26464, n26465, n26466, n26467,
         n26468, n26469, n26470, n26471, n26472, n26473, n26474, n26475,
         n26476, n26477, n26478, n26479, n26480, n26481, n26482, n26483,
         n26484, n26485, n26486, n26487, n26488, n26489, n26490, n26491,
         n26492, n26493, n26494, n26495, n26496, n26497, n26498, n26499,
         n26500, n26501, n26502, n26503, n26504, n26505, n26506, n26507,
         n26508, n26509, n26510, n26511, n26512, n26513, n26514, n26515,
         n26516, n26517, n26518, n26519, n26520, n26521, n26522, n26523,
         n26524, n26525, n26526, n26527, n26528, n26529, n26530, n26531,
         n26532, n26533, n26534, n26535, n26536, n26537, n26538, n26539,
         n26540, n26541, n26542, n26543, n26544, n26545, n26546, n26547,
         n26548, n26549, n26550, n26551, n26552, n26553, n26554, n26555,
         n26556, n26557, n26558, n26559, n26560, n26561, n26562, n26563,
         n26564, n26565, n26566, n26567, n26568, n26569, n26570, n26571,
         n26572, n26573, n26574, n26575, n26576, n26577, n26578, n26579,
         n26580, n26581, n26582, n26583, n26584, n26585, n26586, n26587,
         n26588, n26589, n26590, n26591, n26592, n26593, n26594, n26595,
         n26596, n26597, n26598, n26599, n26600, n26601, n26602, n26603,
         n26604, n26605, n26606, n26607, n26608, n26609, n26610, n26611,
         n26612, n26613, n26614, n26615, n26616, n26617, n26618, n26619,
         n26620, n26621, n26622, n26623, n26624, n26625, n26626, n26627,
         n26628, n26629, n26630, n26631, n26632, n26633, n26634, n26635,
         n26636, n26637, n26638, n26639, n26640, n26641, n26642, n26643,
         n26644, n26645, n26646, n26647, n26648, n26649, n26650, n26651,
         n26652, n26653, n26654, n26655, n26656, n26657, n26658, n26659,
         n26660, n26661, n26662, n26663, n26664, n26665, n26666, n26667,
         n26668, n26669, n26670, n26671, n26672, n26673, n26674, n26675,
         n26676, n26677, n26678, n26679, n26680, n26681, n26682, n26683,
         n26684, n26685, n26686, n26687, n26688, n26689, n26690, n26691,
         n26692, n26693, n26694, n26695, n26696, n26697, n26698, n26699,
         n26700, n26701, n26702, n26703, n26704, n26705, n26706, n26707,
         n26708, n26709, n26710, n26711, n26712, n26713, n26714, n26715,
         n26716, n26717, n26718, n26719, n26720, n26721, n26722, n26723,
         n26724, n26725, n26726, n26727, n26728, n26729, n26730, n26731,
         n26732, n26733, n26734, n26735, n26736, n26737, n26738, n26739,
         n26740, n26741, n26742, n26743, n26744, n26745, n26746, n26747,
         n26748, n26749, n26750, n26751, n26752, n26753, n26754, n26755,
         n26756, n26757, n26758, n26759, n26760, n26761, n26762, n26763,
         n26764, n26765, n26766, n26767, n26768, n26769, n26770, n26771,
         n26772, n26773, n26774, n26775, n26776, n26777, n26778, n26779,
         n26780, n26781, n26782, n26783, n26784, n26785, n26786, n26787,
         n26788, n26789, n26790, n26791, n26792, n26793, n26794, n26795,
         n26796, n26797, n26798, n26799, n26800, n26801, n26802, n26803,
         n26804, n26805, n26806, n26807, n26808, n26809, n26810, n26811,
         n26812, n26813, n26814, n26815, n26816, n26817, n26818, n26819,
         n26820, n26821, n26822, n26823, n26824, n26825, n26826, n26827,
         n26828, n26829, n26830, n26831, n26832, n26833, n26834, n26835,
         n26836, n26837, n26838, n26839, n26840, n26841, n26842, n26843,
         n26844, n26845, n26846, n26847, n26848, n26849, n26850, n26851,
         n26852, n26853, n26854, n26855, n26856, n26857, n26858, n26859,
         n26860, n26861, n26862, n26863, n26864, n26865, n26866, n26867,
         n26868, n26869, n26870, n26871, n26872, n26873, n26874, n26875,
         n26876, n26877, n26878, n26879, n26880, n26881, n26882, n26883,
         n26884, n26885, n26886, n26887, n26888, n26889, n26890, n26891,
         n26892, n26893, n26894, n26895, n26896, n26897, n26898, n26899,
         n26900, n26901, n26902, n26903, n26904, n26905, n26906, n26907,
         n26908, n26909, n26910, n26911, n26912, n26913, n26914, n26915,
         n26916, n26917, n26918, n26919, n26920, n26921, n26922, n26923,
         n26924, n26925, n26926, n26927, n26928, n26929, n26930, n26931,
         n26932, n26933, n26934, n26935, n26936, n26937, n26938, n26939,
         n26940, n26941, n26942, n26943, n26944, n26945, n26946, n26947,
         n26948, n26949, n26950, n26951, n26952, n26953, n26954, n26955,
         n26956, n26957, n26958, n26959, n26960, n26961, n26962, n26963,
         n26964, n26965, n26966, n26967, n26968, n26969, n26970, n26971,
         n26972, n26973, n26974, n26975, n26976, n26977, n26978, n26979,
         n26980, n26981, n26982, n26983, n26984, n26985, n26986, n26987,
         n26988, n26989, n26990, n26991, n26992, n26993, n26994, n26995,
         n26996, n26997, n26998, n26999, n27000, n27001, n27002, n27003,
         n27004, n27005, n27006, n27007, n27008, n27009, n27010, n27011,
         n27012, n27013, n27014, n27015, n27016, n27017, n27018, n27019,
         n27020, n27021, n27022, n27023, n27024, n27025, n27026, n27027,
         n27028, n27029, n27030, n27031, n27032, n27033, n27034, n27035,
         n27036, n27037, n27038, n27039, n27040, n27041, n27042, n27043,
         n27044, n27045, n27046, n27047, n27048, n27049, n27050, n27051,
         n27052, n27053, n27054, n27055, n27056, n27057, n27058, n27059,
         n27060, n27061, n27062, n27063, n27064, n27065, n27066, n27067,
         n27068, n27069, n27070, n27071, n27072, n27073, n27074, n27075,
         n27076, n27077, n27078, n27079, n27080, n27081, n27082, n27083,
         n27084, n27085, n27086, n27087, n27088, n27089, n27090, n27091,
         n27092, n27093, n27094, n27095, n27096, n27097, n27098, n27099,
         n27100, n27101, n27102, n27103, n27104, n27105, n27106, n27107,
         n27108, n27109, n27110, n27111, n27112, n27113, n27114, n27115,
         n27116, n27117, n27118, n27119, n27120, n27121, n27122, n27123,
         n27124, n27125, n27126, n27127, n27128, n27129, n27130, n27131,
         n27132, n27133, n27134, n27135, n27136, n27137, n27138, n27139,
         n27140, n27141, n27142, n27143, n27144, n27145, n27146, n27147,
         n27148, n27149, n27150, n27151, n27152, n27153, n27154, n27155,
         n27156, n27157, n27158, n27159, n27160, n27161, n27162, n27163,
         n27164, n27165, n27166, n27167, n27168, n27169, n27170, n27171,
         n27172, n27173, n27174, n27175, n27176, n27177, n27178, n27179,
         n27180, n27181, n27182, n27183, n27184, n27185, n27186, n27187,
         n27188, n27189, n27190, n27191, n27192, n27193, n27194, n27195,
         n27196, n27197, n27198, n27199, n27200, n27201, n27202, n27203,
         n27204, n27205, n27206, n27207, n27208, n27209, n27210, n27211,
         n27212, n27213, n27214, n27215, n27216, n27217, n27218, n27219,
         n27220, n27221, n27222, n27223, n27224, n27225, n27226, n27227,
         n27228, n27229, n27230, n27231, n27232, n27233, n27234, n27235,
         n27236, n27237, n27238, n27239, n27240, n27241, n27242, n27243,
         n27244, n27245, n27246, n27247, n27248, n27249, n27250, n27251,
         n27252, n27253, n27254, n27255, n27256, n27257, n27258, n27259,
         n27260, n27261, n27262, n27263, n27264, n27265, n27266, n27267,
         n27268, n27269, n27270, n27271, n27272, n27273, n27274, n27275,
         n27276, n27277, n27278, n27279, n27280, n27281, n27282, n27283,
         n27284, n27285, n27286, n27287, n27288, n27289, n27290, n27291,
         n27292, n27293, n27294, n27295, n27296, n27297, n27298, n27299,
         n27300, n27301, n27302, n27303, n27304, n27305, n27306, n27307,
         n27308, n27309, n27310, n27311, n27312, n27313, n27314, n27315,
         n27316, n27317, n27318, n27319, n27320, n27321, n27322, n27323,
         n27324, n27325, n27326, n27327, n27328, n27329, n27330, n27331,
         n27332, n27333, n27334, n27335, n27336, n27337, n27338, n27339,
         n27340, n27341, n27342, n27343, n27344, n27345, n27346, n27347,
         n27348, n27349, n27350, n27351, n27352, n27353, n27354, n27355,
         n27356, n27357, n27358, n27359, n27360, n27361, n27362, n27363,
         n27364, n27365, n27366, n27367, n27368, n27369, n27370, n27371,
         n27372, n27373, n27374, n27375, n27376, n27377, n27378, n27379,
         n27380, n27381, n27382, n27383, n27384, n27385, n27386, n27387,
         n27388, n27389, n27390, n27391, n27392, n27393, n27394, n27395,
         n27396, n27397, n27398, n27399, n27400, n27401, n27402, n27403,
         n27404, n27405, n27406, n27407, n27408, n27409, n27410, n27411,
         n27412, n27413, n27414, n27415, n27416, n27417, n27418, n27419,
         n27420, n27421, n27422, n27423, n27424, n27425, n27426, n27427,
         n27428, n27429, n27430, n27431, n27432, n27433, n27434, n27435,
         n27436, n27437, n27438, n27439, n27440, n27441, n27442, n27443,
         n27444, n27445, n27446, n27447, n27448, n27449, n27450, n27451,
         n27452, n27453, n27454, n27455, n27456, n27457, n27458, n27459,
         n27460, n27461, n27462, n27463, n27464, n27465, n27466, n27467,
         n27468, n27469, n27470, n27471, n27472, n27473, n27474, n27475,
         n27476, n27477, n27478, n27479, n27480, n27481, n27482, n27483,
         n27484, n27485, n27486, n27487, n27488, n27489, n27490, n27491,
         n27492, n27493, n27494, n27495, n27496, n27497, n27498, n27499,
         n27500, n27501, n27502, n27503, n27504, n27505, n27506, n27507,
         n27508, n27509, n27510, n27511, n27512, n27513, n27514, n27515,
         n27516, n27517, n27518, n27519, n27520, n27521, n27522, n27523,
         n27524, n27525, n27526, n27527, n27528, n27529, n27530, n27531,
         n27532, n27533, n27534, n27535, n27536, n27537, n27538, n27539,
         n27540, n27541, n27542, n27543, n27544, n27545, n27546, n27547,
         n27548, n27549, n27550, n27551, n27552, n27553, n27554, n27555,
         n27556, n27557, n27558, n27559, n27560, n27561, n27562, n27563,
         n27564, n27565, n27566, n27567, n27568, n27569, n27570, n27571,
         n27572, n27573, n27574, n27575, n27576, n27577, n27578, n27579,
         n27580, n27581, n27582, n27583, n27584, n27585, n27586, n27587,
         n27588, n27589, n27590, n27591, n27592, n27593, n27594, n27595,
         n27596, n27597, n27598, n27599, n27600, n27601, n27602, n27603,
         n27604, n27605, n27606, n27607, n27608, n27609, n27610, n27611,
         n27612, n27613, n27614, n27615, n27616, n27617, n27618, n27619,
         n27620, n27621, n27622, n27623, n27624, n27625, n27626, n27627,
         n27628, n27629, n27630, n27631, n27632, n27633, n27634, n27635,
         n27636, n27637, n27638, n27639, n27640, n27641, n27642, n27643,
         n27644, n27645, n27646, n27647, n27648, n27649, n27650, n27651,
         n27652, n27653, n27654, n27655, n27656, n27657, n27658, n27659,
         n27660, n27661, n27662, n27663, n27664, n27665, n27666, n27667,
         n27668, n27669, n27670, n27671, n27672, n27673, n27674, n27675,
         n27676, n27677, n27678, n27679, n27680, n27681, n27682, n27683,
         n27684, n27685, n27686, n27687, n27688, n27689, n27690, n27691,
         n27692, n27693, n27694, n27695, n27696, n27697, n27698, n27699,
         n27700, n27701, n27702, n27703, n27704, n27705, n27706, n27707,
         n27708, n27709, n27710, n27711, n27712, n27713, n27714, n27715,
         n27716, n27717, n27718, n27719, n27720, n27721, n27722, n27723,
         n27724, n27725, n27726, n27727, n27728, n27729, n27730, n27731,
         n27732, n27733, n27734, n27735, n27736, n27737, n27738, n27739,
         n27740, n27741, n27742, n27743, n27744, n27745, n27746, n27747,
         n27748, n27749, n27750, n27751, n27752, n27753, n27754, n27755,
         n27756, n27757, n27758, n27759, n27760, n27761, n27762, n27763,
         n27764, n27765, n27766, n27767, n27768, n27769, n27770, n27771,
         n27772, n27773, n27774, n27775, n27776, n27777, n27778, n27779,
         n27780, n27781, n27782, n27783, n27784, n27785, n27786, n27787,
         n27788, n27789, n27790, n27791, n27792, n27793, n27794, n27795,
         n27796, n27797, n27798, n27799, n27800, n27801, n27802, n27803,
         n27804, n27805, n27806, n27807, n27808, n27809, n27810, n27811,
         n27812, n27813, n27814, n27815, n27816, n27817, n27818, n27819,
         n27820, n27821, n27822, n27823, n27824, n27825, n27826, n27827,
         n27828, n27829, n27830, n27831, n27832, n27833, n27834, n27835,
         n27836, n27837, n27838, n27839, n27840, n27841, n27842, n27843,
         n27844, n27845, n27846, n27847, n27848, n27849, n27850, n27851,
         n27852, n27853, n27854, n27855, n27856, n27857, n27858, n27859,
         n27860, n27861, n27862, n27863, n27864, n27865, n27866, n27867,
         n27868, n27869, n27870, n27871, n27872, n27873, n27874, n27875,
         n27876, n27877, n27878, n27879, n27880, n27881, n27882, n27883,
         n27884, n27885, n27886, n27887, n27888, n27889, n27890, n27891,
         n27892, n27893, n27894, n27895, n27896, n27897, n27898, n27899,
         n27900, n27901, n27902, n27903, n27904, n27905, n27906, n27907,
         n27908, n27909, n27910, n27911, n27912, n27913, n27914, n27915,
         n27916, n27917, n27918, n27919, n27920, n27921, n27922, n27923,
         n27924, n27925, n27926, n27927, n27928, n27929, n27930, n27931,
         n27932, n27933, n27934, n27935, n27936, n27937, n27938, n27939,
         n27940, n27941, n27942, n27943, n27944, n27945, n27946, n27947,
         n27948, n27949, n27950, n27951, n27952, n27953, n27954, n27955,
         n27956, n27957, n27958, n27959, n27960, n27961, n27962, n27963,
         n27964, n27965, n27966, n27967, n27968, n27969, n27970, n27971,
         n27972, n27973, n27974, n27975, n27976, n27977, n27978, n27979,
         n27980, n27981, n27982, n27983, n27984, n27985, n27986, n27987,
         n27988, n27989, n27990, n27991, n27992, n27993, n27994, n27995,
         n27996, n27997, n27998, n27999, n28000, n28001, n28002, n28003,
         n28004, n28005, n28006, n28007, n28008, n28009, n28010, n28011,
         n28012, n28013, n28014, n28015, n28016, n28017, n28018, n28019,
         n28020, n28021, n28022, n28023, n28024, n28025, n28026, n28027,
         n28028, n28029, n28030, n28031, n28032, n28033, n28034, n28035,
         n28036, n28037, n28038, n28039, n28040, n28041, n28042, n28043,
         n28044, n28045, n28046, n28047, n28048, n28049, n28050, n28051,
         n28052, n28053, n28054, n28055, n28056, n28057, n28058, n28059,
         n28060, n28061, n28062, n28063, n28064, n28065, n28066, n28067,
         n28068, n28069, n28070, n28071, n28072, n28073, n28074, n28075,
         n28076, n28077, n28078, n28079, n28080, n28081, n28082, n28083,
         n28084, n28085, n28086, n28087, n28088, n28089, n28090, n28091,
         n28092, n28093, n28094, n28095, n28096, n28097, n28098, n28099,
         n28100, n28101, n28102, n28103, n28104, n28105, n28106, n28107,
         n28108, n28109, n28110, n28111, n28112, n28113, n28114, n28115,
         n28116, n28117, n28118, n28119, n28120, n28121, n28122, n28123,
         n28124, n28125, n28126, n28127, n28128, n28129, n28130, n28131,
         n28132, n28133, n28134, n28135, n28136, n28137, n28138, n28139,
         n28140, n28141, n28142, n28143, n28144, n28145, n28146, n28147,
         n28148, n28149, n28150, n28151, n28152, n28153, n28154, n28155,
         n28156, n28157, n28158, n28159, n28160, n28161, n28162, n28163,
         n28164, n28165, n28166, n28167, n28168, n28169, n28170, n28171,
         n28172, n28173, n28174, n28175, n28176, n28177, n28178, n28179,
         n28180, n28181, n28182, n28183, n28184, n28185, n28186, n28187,
         n28188, n28189, n28190, n28191, n28192, n28193, n28194, n28195,
         n28196, n28197, n28198, n28199, n28200, n28201, n28202, n28203,
         n28204, n28205, n28206, n28207, n28208, n28209, n28210, n28211,
         n28212, n28213, n28214, n28215, n28216, n28217, n28218, n28219,
         n28220, n28221, n28222, n28223, n28224, n28225, n28226, n28227,
         n28228, n28229, n28230, n28231, n28232, n28233, n28234, n28235,
         n28236, n28237, n28238, n28239, n28240, n28241, n28242, n28243,
         n28244, n28245, n28246, n28247, n28248, n28249, n28250, n28251,
         n28252, n28253, n28254, n28255, n28256, n28257, n28258, n28259,
         n28260, n28261, n28262, n28263, n28264, n28265, n28266, n28267,
         n28268, n28269, n28270, n28271, n28272, n28273, n28274, n28275,
         n28276, n28277, n28278, n28279, n28280, n28281, n28282, n28283,
         n28284, n28285, n28286, n28287, n28288, n28289, n28290, n28291,
         n28292, n28293, n28294, n28295, n28296, n28297, n28298, n28299,
         n28300, n28301, n28302, n28303, n28304, n28305, n28306, n28307,
         n28308, n28309, n28310, n28311, n28312, n28313, n28314, n28315,
         n28316, n28317, n28318, n28319, n28320, n28321, n28322, n28323,
         n28324, n28325, n28326, n28327, n28328, n28329, n28330, n28331,
         n28332, n28333, n28334, n28335, n28336, n28337, n28338, n28339,
         n28340, n28341, n28342, n28343, n28344, n28345, n28346, n28347,
         n28348, n28349, n28350, n28351, n28352, n28353, n28354, n28355,
         n28356, n28357, n28358, n28359, n28360, n28361, n28362, n28363,
         n28364, n28365, n28366, n28367, n28368, n28369, n28370, n28371,
         n28372, n28373, n28374, n28375, n28376, n28377, n28378, n28379,
         n28380, n28381, n28382, n28383, n28384, n28385, n28386, n28387,
         n28388, n28389, n28390, n28391, n28392, n28393, n28394, n28395,
         n28396, n28397, n28398, n28399, n28400, n28401, n28402, n28403,
         n28404, n28405, n28406, n28407, n28408, n28409, n28410, n28411,
         n28412, n28413, n28414, n28415, n28416, n28417, n28418, n28419,
         n28420, n28421, n28422, n28423, n28424, n28425, n28426, n28427,
         n28428, n28429, n28430, n28431, n28432, n28433, n28434, n28435,
         n28436, n28437, n28438, n28439, n28440, n28441, n28442, n28443,
         n28444, n28445, n28446, n28447, n28448, n28449, n28450, n28451,
         n28452, n28453, n28454, n28455, n28456, n28457, n28458, n28459,
         n28460, n28461, n28462, n28463, n28464, n28465, n28466, n28467,
         n28468, n28469, n28470, n28471, n28472, n28473, n28474, n28475,
         n28476, n28477, n28478, n28479, n28480, n28481, n28482, n28483,
         n28484, n28485, n28486, n28487, n28488, n28489, n28490, n28491,
         n28492, n28493, n28494, n28495, n28496, n28497, n28498, n28499,
         n28500, n28501, n28502, n28503, n28504, n28505, n28506, n28507,
         n28508, n28509, n28510, n28511, n28512, n28513, n28514, n28515,
         n28516, n28517, n28518, n28519, n28520, n28521, n28522, n28523,
         n28524, n28525, n28526, n28527, n28528, n28529, n28530, n28531,
         n28532, n28533, n28534, n28535, n28536, n28537, n28538, n28539,
         n28540, n28541, n28542, n28543, n28544, n28545, n28546, n28547,
         n28548, n28549, n28550, n28551, n28552, n28553, n28554, n28555,
         n28556, n28557, n28558, n28559, n28560, n28561, n28562, n28563,
         n28564, n28565, n28566, n28567, n28568, n28569, n28570, n28571,
         n28572, n28573, n28574, n28575, n28576, n28577, n28578, n28579,
         n28580, n28581, n28582, n28583, n28584, n28585, n28586, n28587,
         n28588, n28589, n28590, n28591, n28592, n28593, n28594, n28595,
         n28596, n28597, n28598, n28599, n28600, n28601, n28602, n28603,
         n28604, n28605, n28606, n28607, n28608, n28609, n28610, n28611,
         n28612, n28613, n28614, n28615, n28616, n28617, n28618, n28619,
         n28620, n28621, n28622, n28623, n28624, n28625, n28626, n28627,
         n28628, n28629, n28630, n28631, n28632, n28633, n28634, n28635,
         n28636, n28637, n28638, n28639, n28640, n28641, n28642, n28643,
         n28644, n28645, n28646, n28647, n28648, n28649, n28650, n28651,
         n28652, n28653, n28654, n28655, n28656, n28657, n28658, n28659,
         n28660, n28661, n28662, n28663, n28664, n28665, n28666, n28667,
         n28668, n28669, n28670, n28671, n28672, n28673, n28674, n28675,
         n28676, n28677, n28678, n28679, n28680, n28681, n28682, n28683,
         n28684, n28685, n28686, n28687, n28688, n28689, n28690, n28691,
         n28692, n28693, n28694, n28695, n28696, n28697, n28698, n28699,
         n28700, n28701, n28702, n28703, n28704, n28705, n28706, n28707,
         n28708, n28709, n28710, n28711, n28712, n28713, n28714, n28715,
         n28716, n28717, n28718, n28719, n28720, n28721, n28722, n28723,
         n28724, n28725, n28726, n28727, n28728, n28729, n28730, n28731,
         n28732, n28733, n28734, n28735, n28736, n28737, n28738, n28739,
         n28740, n28741, n28742, n28743, n28744, n28745, n28746, n28747,
         n28748, n28749, n28750, n28751, n28752, n28753, n28754, n28755,
         n28756, n28757, n28758, n28759, n28760, n28761, n28762, n28763,
         n28764, n28765, n28766, n28767, n28768, n28769, n28770, n28771,
         n28772, n28773, n28774, n28775, n28776, n28777, n28778, n28779,
         n28780, n28781, n28782, n28783, n28784, n28785, n28786, n28787,
         n28788, n28789, n28790, n28791, n28792, n28793, n28794, n28795,
         n28796, n28797, n28798, n28799, n28800, n28801, n28802, n28803,
         n28804, n28805, n28806, n28807, n28808, n28809, n28810, n28811,
         n28812, n28813, n28814, n28815, n28816, n28817, n28818, n28819,
         n28820, n28821, n28822, n28823, n28824, n28825, n28826, n28827,
         n28828, n28829, n28830, n28831, n28832, n28833, n28834, n28835,
         n28836, n28837, n28838, n28839, n28840, n28841, n28842, n28843,
         n28844, n28845, n28846, n28847, n28848, n28849, n28850, n28851,
         n28852, n28853, n28854, n28855, n28856, n28857, n28858, n28859,
         n28860, n28861, n28862, n28863, n28864, n28865, n28866, n28867,
         n28868, n28869, n28870, n28871, n28872, n28873, n28874, n28875,
         n28876, n28877, n28878, n28879, n28880, n28881, n28882, n28883,
         n28884, n28885, n28886, n28887, n28888, n28889, n28890, n28891,
         n28892, n28893, n28894, n28895, n28896, n28897, n28898, n28899,
         n28900, n28901, n28902, n28903, n28904, n28905, n28906, n28907,
         n28908, n28909, n28910, n28911, n28912, n28913, n28914, n28915,
         n28916, n28917, n28918, n28919, n28920, n28921, n28922, n28923,
         n28924, n28925, n28926, n28927, n28928, n28929, n28930, n28931,
         n28932, n28933, n28934, n28935, n28936, n28937, n28938, n28939,
         n28940, n28941, n28942, n28943, n28944, n28945, n28946, n28947,
         n28948, n28949, n28950, n28951, n28952, n28953, n28954, n28955,
         n28956, n28957, n28958, n28959, n28960, n28961, n28962, n28963,
         n28964, n28965, n28966, n28967, n28968, n28969, n28970, n28971,
         n28972, n28973, n28974, n28975, n28976, n28977, n28978, n28979,
         n28980, n28981, n28982, n28983, n28984, n28985, n28986, n28987,
         n28988, n28989, n28990, n28991, n28992, n28993, n28994, n28995,
         n28996, n28997, n28998, n28999, n29000, n29001, n29002, n29003,
         n29004, n29005, n29006, n29007, n29008, n29009, n29010, n29011,
         n29012, n29013, n29014, n29015, n29016, n29017, n29018, n29019,
         n29020, n29021, n29022, n29023, n29024, n29025, n29026, n29027,
         n29028, n29029, n29030, n29031, n29032, n29033, n29034, n29035,
         n29036, n29037, n29038, n29039, n29040, n29041, n29042, n29043,
         n29044, n29045, n29046, n29047, n29048, n29049, n29050, n29051,
         n29052, n29053, n29054, n29055, n29056, n29057, n29058, n29059,
         n29060, n29061, n29062, n29063, n29064, n29065, n29066, n29067,
         n29068, n29069, n29070, n29071, n29072, n29073, n29074, n29075,
         n29076, n29077, n29078, n29079, n29080, n29081, n29082, n29083,
         n29084, n29085, n29086, n29087, n29088, n29089, n29090, n29091,
         n29092, n29093, n29094, n29095, n29096, n29097, n29098, n29099,
         n29100, n29101, n29102, n29103, n29104, n29105, n29106, n29107,
         n29108, n29109, n29110, n29111, n29112, n29113, n29114, n29115,
         n29116, n29117, n29118, n29119, n29120, n29121, n29122, n29123,
         n29124, n29125, n29126, n29127, n29128, n29129, n29130, n29131,
         n29132, n29133, n29134, n29135, n29136, n29137, n29138, n29139,
         n29140, n29141, n29142, n29143, n29144, n29145, n29146, n29147,
         n29148, n29149, n29150, n29151, n29152, n29153, n29154, n29155,
         n29156, n29157, n29158, n29159, n29160, n29161, n29162, n29163,
         n29164, n29165, n29166, n29167, n29168, n29169, n29170, n29171,
         n29172, n29173, n29174, n29175, n29176, n29177, n29178, n29179,
         n29180, n29181, n29182, n29183, n29184, n29185, n29186, n29187,
         n29188, n29189, n29190, n29191, n29192, n29193, n29194, n29195,
         n29196, n29197, n29198, n29199, n29200, n29201, n29202, n29203,
         n29204, n29205, n29206, n29207, n29208, n29209, n29210, n29211,
         n29212, n29213, n29214, n29215, n29216, n29217, n29218, n29219,
         n29220, n29221, n29222, n29223, n29224, n29225, n29226, n29227,
         n29228, n29229, n29230, n29231, n29232, n29233, n29234, n29235,
         n29236, n29237, n29238, n29239, n29240, n29241, n29242, n29243,
         n29244, n29245, n29246, n29247, n29248, n29249, n29250, n29251,
         n29252, n29253, n29254, n29255, n29256, n29257, n29258, n29259,
         n29260, n29261, n29262, n29263, n29264, n29265, n29266, n29267,
         n29268, n29269, n29270, n29271, n29272, n29273, n29274, n29275,
         n29276, n29277, n29278, n29279, n29280, n29281, n29282, n29283,
         n29284, n29285, n29286, n29287, n29288, n29289, n29290, n29291,
         n29292, n29293, n29294, n29295, n29296, n29297, n29298, n29299,
         n29300, n29301, n29302, n29303, n29304, n29305, n29306, n29307,
         n29308, n29309, n29310, n29311, n29312, n29313, n29314, n29315,
         n29316, n29317, n29318, n29319, n29320, n29321, n29322, n29323,
         n29324, n29325, n29326, n29327, n29328, n29329, n29330, n29331,
         n29332, n29333, n29334, n29335, n29336, n29337, n29338, n29339,
         n29340, n29341, n29342, n29343, n29344, n29345, n29346, n29347,
         n29348, n29349, n29350, n29351, n29352, n29353, n29354, n29355,
         n29356, n29357, n29358, n29359, n29360, n29361, n29362, n29363,
         n29364, n29365, n29366, n29367, n29368, n29369, n29370, n29371,
         n29372, n29373, n29374, n29375, n29376, n29377, n29378, n29379,
         n29380, n29381, n29382, n29383, n29384, n29385, n29386, n29387,
         n29388, n29389, n29390, n29391, n29392, n29393, n29394, n29395,
         n29396, n29397, n29398, n29399, n29400, n29401, n29402, n29403,
         n29404, n29405, n29406, n29407, n29408, n29409, n29410, n29411,
         n29412, n29413, n29414, n29415, n29416, n29417, n29418, n29419,
         n29420, n29421, n29422, n29423, n29424, n29425, n29426, n29427,
         n29428, n29429, n29430, n29431, n29432, n29433, n29434, n29435,
         n29436, n29437, n29438, n29439, n29440, n29441, n29442, n29443,
         n29444, n29445, n29446, n29447, n29448, n29449, n29450, n29451,
         n29452, n29453, n29454, n29455, n29456, n29457, n29458, n29459,
         n29460, n29461, n29462, n29463, n29464, n29465, n29466, n29467,
         n29468, n29469, n29470, n29471, n29472, n29473, n29474, n29475,
         n29476, n29477, n29478, n29479, n29480, n29481, n29482, n29483,
         n29484, n29485, n29486, n29487, n29488, n29489, n29490, n29491,
         n29492, n29493, n29494, n29495, n29496, n29497, n29498, n29499,
         n29500, n29501, n29502, n29503, n29504, n29505, n29506, n29507,
         n29508, n29509, n29510, n29511, n29512, n29513, n29514, n29515,
         n29516, n29517, n29518, n29519, n29520, n29521, n29522, n29523,
         n29524, n29525, n29526, n29527, n29528, n29529, n29530, n29531,
         n29532, n29533, n29534, n29535, n29536, n29537, n29538, n29539,
         n29540, n29541, n29542, n29543, n29544, n29545, n29546, n29547,
         n29548, n29549, n29550, n29551, n29552, n29553, n29554, n29555,
         n29556, n29557, n29558, n29559, n29560, n29561, n29562, n29563,
         n29564, n29565, n29566, n29567, n29568, n29569, n29570, n29571,
         n29572, n29573, n29574, n29575, n29576, n29577, n29578, n29579,
         n29580, n29581, n29582, n29583, n29584, n29585, n29586, n29587,
         n29588, n29589, n29590, n29591, n29592, n29593, n29594, n29595,
         n29596, n29597, n29598, n29599, n29600, n29601, n29602, n29603,
         n29604, n29605, n29606, n29607, n29608, n29609, n29610, n29611,
         n29612, n29613, n29614, n29615, n29616, n29617, n29618, n29619,
         n29620, n29621, n29622, n29623, n29624, n29625, n29626, n29627,
         n29628, n29629, n29630, n29631, n29632, n29633, n29634, n29635,
         n29636, n29637, n29638, n29639, n29640, n29641, n29642, n29643,
         n29644, n29645, n29646, n29647, n29648, n29649, n29650, n29651,
         n29652, n29653, n29654, n29655, n29656, n29657, n29658, n29659,
         n29660, n29661, n29662, n29663, n29664, n29665, n29666, n29667,
         n29668, n29669, n29670, n29671, n29672, n29673, n29674, n29675,
         n29676, n29677, n29678, n29679, n29680, n29681, n29682, n29683,
         n29684, n29685, n29686, n29687, n29688, n29689, n29690, n29691,
         n29692, n29693, n29694, n29695, n29696, n29697, n29698, n29699,
         n29700, n29701, n29702, n29703, n29704, n29705, n29706, n29707,
         n29708, n29709, n29710, n29711, n29712, n29713, n29714, n29715,
         n29716, n29717, n29718, n29719, n29720, n29721, n29722, n29723,
         n29724, n29725, n29726, n29727, n29728, n29729, n29730, n29731,
         n29732, n29733, n29734, n29735, n29736, n29737, n29738, n29739,
         n29740, n29741, n29742, n29743, n29744, n29745, n29746, n29747,
         n29748, n29749, n29750, n29751, n29752, n29753, n29754, n29755,
         n29756, n29757, n29758, n29759, n29760, n29761, n29762, n29763,
         n29764, n29765, n29766, n29767, n29768, n29769, n29770, n29771,
         n29772, n29773, n29774, n29775, n29776, n29777, n29778, n29779,
         n29780, n29781, n29782, n29783, n29784, n29785, n29786, n29787,
         n29788, n29789, n29790, n29791, n29792, n29793, n29794, n29795,
         n29796, n29797, n29798, n29799, n29800, n29801, n29802, n29803,
         n29804, n29805, n29806, n29807, n29808, n29809, n29810, n29811,
         n29812, n29813, n29814, n29815, n29816, n29817, n29818, n29819,
         n29820, n29821, n29822, n29823, n29824, n29825, n29826, n29827,
         n29828, n29829, n29830, n29831, n29832, n29833, n29834, n29835,
         n29836, n29837, n29838, n29839, n29840, n29841, n29842, n29843,
         n29844, n29845, n29846, n29847, n29848, n29849, n29850, n29851,
         n29852, n29853, n29854, n29855, n29856, n29857, n29858, n29859,
         n29860, n29861, n29862, n29863, n29864, n29865, n29866, n29867,
         n29868, n29869, n29870, n29871, n29872, n29873, n29874, n29875,
         n29876, n29877, n29878, n29879, n29880, n29881, n29882, n29883,
         n29884, n29885, n29886, n29887, n29888, n29889, n29890, n29891,
         n29892, n29893, n29894, n29895, n29896, n29897, n29898, n29899,
         n29900, n29901, n29902, n29903, n29904, n29905, n29906, n29907,
         n29908, n29909, n29910, n29911, n29912, n29913, n29914, n29915,
         n29916, n29917, n29918, n29919, n29920, n29921, n29922, n29923,
         n29924, n29925, n29926, n29927, n29928, n29929, n29930, n29931,
         n29932, n29933, n29934, n29935, n29936, n29937, n29938, n29939,
         n29940, n29941, n29942, n29943, n29944, n29945, n29946, n29947,
         n29948, n29949, n29950, n29951, n29952, n29953, n29954, n29955,
         n29956, n29957, n29958, n29959, n29960, n29961, n29962, n29963,
         n29964, n29965, n29966, n29967, n29968, n29969, n29970, n29971,
         n29972, n29973, n29974, n29975, n29976, n29977, n29978, n29979,
         n29980, n29981, n29982, n29983, n29984, n29985, n29986, n29987,
         n29988, n29989, n29990, n29991, n29992, n29993, n29994, n29995,
         n29996, n29997, n29998, n29999, n30000, n30001, n30002, n30003,
         n30004, n30005, n30006, n30007, n30008, n30009, n30010, n30011,
         n30012, n30013, n30014, n30015, n30016, n30017, n30018, n30019,
         n30020, n30021, n30022, n30023, n30024, n30025, n30026, n30027,
         n30028, n30029, n30030, n30031, n30032, n30033, n30034, n30035,
         n30036, n30037, n30038, n30039, n30040, n30041, n30042, n30043,
         n30044, n30045, n30046, n30047, n30048, n30049, n30050, n30051,
         n30052, n30053, n30054, n30055, n30056, n30057, n30058, n30059,
         n30060, n30061, n30062, n30063, n30064, n30065, n30066, n30067,
         n30068, n30069, n30070, n30071, n30072, n30073, n30074, n30075,
         n30076, n30077, n30078, n30079, n30080, n30081, n30082, n30083,
         n30084, n30085, n30086, n30087, n30088, n30089, n30090, n30091,
         n30092, n30093, n30094, n30095, n30096, n30097, n30098, n30099,
         n30100, n30101, n30102, n30103, n30104, n30105, n30106, n30107,
         n30108, n30109, n30110, n30111, n30112, n30113, n30114, n30115,
         n30116, n30117, n30118, n30119, n30120, n30121, n30122, n30123,
         n30124, n30125, n30126, n30127, n30128, n30129, n30130, n30131,
         n30132, n30133, n30134, n30135, n30136, n30137, n30138, n30139,
         n30140, n30141, n30142, n30143, n30144, n30145, n30146, n30147,
         n30148, n30149, n30150, n30151, n30152, n30153, n30154, n30155,
         n30156, n30157, n30158, n30159, n30160, n30161, n30162, n30163,
         n30164, n30165, n30166, n30167, n30168, n30169, n30170, n30171,
         n30172, n30173, n30174, n30175, n30176, n30177, n30178, n30179,
         n30180, n30181, n30182, n30183, n30184, n30185, n30186, n30187,
         n30188, n30189, n30190, n30191, n30192, n30193, n30194, n30195,
         n30196, n30197, n30198, n30199, n30200, n30201, n30202, n30203,
         n30204, n30205, n30206, n30207, n30208, n30209, n30210, n30211,
         n30212, n30213, n30214, n30215, n30216, n30217, n30218, n30219,
         n30220, n30221, n30222, n30223, n30224, n30225, n30226, n30227,
         n30228, n30229, n30230, n30231, n30232, n30233, n30234, n30235,
         n30236, n30237, n30238, n30239, n30240, n30241, n30242, n30243,
         n30244, n30245, n30246, n30247, n30248, n30249, n30250, n30251,
         n30252, n30253, n30254, n30255, n30256, n30257, n30258, n30259,
         n30260, n30261, n30262, n30263, n30264, n30265, n30266, n30267,
         n30268, n30269, n30270, n30271, n30272, n30273, n30274, n30275,
         n30276, n30277, n30278, n30279, n30280, n30281, n30282, n30283,
         n30284, n30285, n30286, n30287, n30288, n30289, n30290, n30291,
         n30292, n30293, n30294, n30295, n30296, n30297, n30298, n30299,
         n30300, n30301, n30302, n30303, n30304, n30305, n30306, n30307,
         n30308, n30309, n30310, n30311, n30312, n30313, n30314, n30315,
         n30316, n30317, n30318, n30319, n30320, n30321, n30322, n30323,
         n30324, n30325, n30326, n30327, n30328, n30329, n30330, n30331,
         n30332, n30333, n30334, n30335, n30336, n30337, n30338, n30339,
         n30340, n30341, n30342, n30343, n30344, n30345, n30346, n30347,
         n30348, n30349, n30350, n30351, n30352, n30353, n30354, n30355,
         n30356, n30357, n30358, n30359, n30360, n30361, n30362, n30363,
         n30364, n30365, n30366, n30367, n30368, n30369, n30370, n30371,
         n30372, n30373, n30374, n30375, n30376, n30377, n30378, n30379,
         n30380, n30381, n30382, n30383, n30384, n30385, n30386, n30387,
         n30388, n30389, n30390, n30391, n30392, n30393, n30394, n30395,
         n30396, n30397, n30398, n30399, n30400, n30401, n30402, n30403,
         n30404, n30405, n30406, n30407, n30408, n30409, n30410, n30411,
         n30412, n30413, n30414, n30415, n30416, n30417, n30418, n30419,
         n30420, n30421, n30422, n30423, n30424, n30425, n30426, n30427,
         n30428, n30429, n30430, n30431, n30432, n30433, n30434, n30435,
         n30436, n30437, n30438, n30439, n30440, n30441, n30442, n30443,
         n30444, n30445, n30446, n30447, n30448, n30449, n30450, n30451,
         n30452, n30453, n30454, n30455, n30456, n30457, n30458, n30459,
         n30460, n30461, n30462, n30463, n30464, n30465, n30466, n30467,
         n30468, n30469, n30470, n30471, n30472, n30473, n30474, n30475,
         n30476, n30477, n30478, n30479, n30480, n30481, n30482, n30483,
         n30484, n30485, n30486, n30487, n30488, n30489, n30490, n30491,
         n30492, n30493, n30494, n30495, n30496, n30497, n30498, n30499,
         n30500, n30501, n30502, n30503, n30504, n30505, n30506, n30507,
         n30508, n30509, n30510, n30511, n30512, n30513, n30514, n30515,
         n30516, n30517, n30518, n30519, n30520, n30521, n30522, n30523,
         n30524, n30525, n30526, n30527, n30528, n30529, n30530, n30531,
         n30532, n30533, n30534, n30535, n30536, n30537, n30538, n30539,
         n30540, n30541, n30542, n30543, n30544, n30545, n30546, n30547,
         n30548, n30549, n30550, n30551, n30552, n30553, n30554, n30555,
         n30556, n30557, n30558, n30559, n30560, n30561, n30562, n30563,
         n30564, n30565, n30566, n30567, n30568, n30569, n30570, n30571,
         n30572, n30573, n30574, n30575, n30576, n30577, n30578, n30579,
         n30580, n30581, n30582, n30583, n30584, n30585, n30586, n30587,
         n30588, n30589, n30590, n30591, n30592, n30593, n30594, n30595,
         n30596, n30597, n30598, n30599, n30600, n30601, n30602, n30603,
         n30604, n30605, n30606, n30607, n30608, n30609, n30610, n30611,
         n30612, n30613, n30614, n30615, n30616, n30617, n30618, n30619,
         n30620, n30621, n30622, n30623, n30624, n30625, n30626, n30627,
         n30628, n30629, n30630, n30631, n30632, n30633, n30634, n30635,
         n30636, n30637, n30638, n30639, n30640, n30641, n30642, n30643,
         n30644, n30645, n30646, n30647, n30648, n30649, n30650, n30651,
         n30652, n30653, n30654, n30655, n30656, n30657, n30658, n30659,
         n30660, n30661, n30662, n30663, n30664, n30665, n30666, n30667,
         n30668, n30669, n30670, n30671, n30672, n30673, n30674, n30675,
         n30676, n30677, n30678, n30679, n30680, n30681, n30682, n30683,
         n30684, n30685, n30686, n30687, n30688, n30689, n30690, n30691,
         n30692, n30693, n30694, n30695, n30696, n30697, n30698, n30699,
         n30700, n30701, n30702, n30703, n30704, n30705, n30706, n30707,
         n30708, n30709, n30710, n30711, n30712, n30713, n30714, n30715,
         n30716, n30717, n30718, n30719, n30720, n30721, n30722, n30723,
         n30724, n30725, n30726, n30727, n30728, n30729, n30730, n30731,
         n30732, n30733, n30734, n30735, n30736, n30737, n30738, n30739,
         n30740, n30741, n30742, n30743, n30744, n30745, n30746, n30747,
         n30748, n30749, n30750, n30751, n30752, n30753, n30754, n30755,
         n30756, n30757, n30758, n30759, n30760, n30761, n30762, n30763,
         n30764, n30765, n30766, n30767, n30768, n30769, n30770, n30771,
         n30772, n30773, n30774, n30775, n30776, n30777, n30778, n30779,
         n30780, n30781, n30782, n30783, n30784, n30785, n30786, n30787,
         n30788, n30789, n30790, n30791, n30792, n30793, n30794, n30795,
         n30796, n30797, n30798, n30799, n30800, n30801, n30802, n30803,
         n30804, n30805, n30806, n30807, n30808, n30809, n30810, n30811,
         n30812, n30813, n30814, n30815, n30816, n30817, n30818, n30819,
         n30820, n30821, n30822, n30823, n30824, n30825, n30826, n30827,
         n30828, n30829, n30830, n30831, n30832, n30833, n30834, n30835,
         n30836, n30837, n30838, n30839, n30840, n30841, n30842, n30843,
         n30844, n30845, n30846, n30847, n30848, n30849, n30850, n30851,
         n30852, n30853, n30854, n30855, n30856, n30857, n30858, n30859,
         n30860, n30861, n30862, n30863, n30864, n30865, n30866, n30867,
         n30868, n30869, n30870, n30871, n30872, n30873, n30874, n30875,
         n30876, n30877, n30878, n30879, n30880, n30881, n30882, n30883,
         n30884, n30885, n30886, n30887, n30888, n30889, n30890, n30891,
         n30892, n30893, n30894, n30895, n30896, n30897, n30898, n30899,
         n30900, n30901, n30902, n30903, n30904, n30905, n30906, n30907,
         n30908, n30909, n30910, n30911, n30912, n30913, n30914, n30915,
         n30916, n30917, n30918, n30919, n30920, n30921, n30922, n30923,
         n30924, n30925, n30926, n30927, n30928, n30929, n30930, n30931,
         n30932, n30933, n30934, n30935, n30936, n30937, n30938, n30939,
         n30940, n30941, n30942, n30943, n30944, n30945, n30946, n30947,
         n30948, n30949, n30950, n30951, n30952, n30953, n30954, n30955,
         n30956, n30957, n30958, n30959, n30960, n30961, n30962, n30963,
         n30964, n30965, n30966, n30967, n30968, n30969, n30970, n30971,
         n30972, n30973, n30974, n30975, n30976, n30977, n30978, n30979,
         n30980, n30981, n30982, n30983, n30984, n30985, n30986, n30987,
         n30988, n30989, n30990, n30991, n30992, n30993, n30994, n30995,
         n30996, n30997, n30998, n30999, n31000, n31001, n31002, n31003,
         n31004, n31005, n31006, n31007, n31008, n31009, n31010, n31011,
         n31012, n31013, n31014, n31015, n31016, n31017, n31018, n31019,
         n31020, n31021, n31022, n31023, n31024, n31025, n31026, n31027,
         n31028, n31029, n31030, n31031, n31032, n31033, n31034, n31035,
         n31036, n31037, n31038, n31039, n31040, n31041, n31042, n31043,
         n31044, n31045, n31046, n31047, n31048, n31049, n31050, n31051,
         n31052, n31053, n31054, n31055, n31056, n31057, n31058, n31059,
         n31060, n31061, n31062, n31063, n31064, n31065, n31066, n31067,
         n31068, n31069, n31070, n31071, n31072, n31073, n31074, n31075,
         n31076, n31077, n31078, n31079, n31080, n31081, n31082, n31083,
         n31084, n31085, n31086, n31087, n31088, n31089, n31090, n31091,
         n31092, n31093, n31094, n31095, n31096, n31097, n31098, n31099,
         n31100, n31101, n31102, n31103, n31104, n31105, n31106, n31107,
         n31108, n31109, n31110, n31111, n31112, n31113, n31114, n31115,
         n31116, n31117, n31118, n31119, n31120, n31121, n31122, n31123,
         n31124, n31125, n31126, n31127, n31128, n31129, n31130, n31131,
         n31132, n31133, n31134, n31135, n31136, n31137, n31138, n31139,
         n31140, n31141, n31142, n31143, n31144, n31145, n31146, n31147,
         n31148, n31149, n31150, n31151, n31152, n31153, n31154, n31155,
         n31156, n31157, n31158, n31159, n31160, n31161, n31162, n31163,
         n31164, n31165, n31166, n31167, n31168, n31169, n31170, n31171,
         n31172, n31173, n31174, n31175, n31176, n31177, n31178, n31179,
         n31180, n31181, n31182, n31183, n31184, n31185, n31186, n31187,
         n31188, n31189, n31190, n31191, n31192, n31193, n31194, n31195,
         n31196, n31197, n31198, n31199, n31200, n31201, n31202, n31203,
         n31204, n31205, n31206, n31207, n31208, n31209, n31210, n31211,
         n31212, n31213, n31214, n31215, n31216, n31217, n31218, n31219,
         n31220, n31221, n31222, n31223, n31224, n31225, n31226, n31227,
         n31228, n31229, n31230, n31231, n31232, n31233, n31234, n31235,
         n31236, n31237, n31238, n31239, n31240, n31241, n31242, n31243,
         n31244, n31245, n31246, n31247, n31248, n31249, n31250, n31251,
         n31252, n31253, n31254, n31255, n31256, n31257, n31258, n31259,
         n31260, n31261, n31262, n31263, n31264, n31265, n31266, n31267,
         n31268, n31269, n31270, n31271, n31272, n31273, n31274, n31275,
         n31276, n31277, n31278, n31279, n31280, n31281, n31282, n31283,
         n31284, n31285, n31286, n31287, n31288, n31289, n31290, n31291,
         n31292, n31293, n31294, n31295, n31296, n31297, n31298, n31299,
         n31300, n31301, n31302, n31303, n31304, n31305, n31306, n31307,
         n31308, n31309, n31310, n31311, n31312, n31313, n31314, n31315,
         n31316, n31317, n31318, n31319, n31320, n31321, n31322, n31323,
         n31324, n31325, n31326, n31327, n31328, n31329, n31330, n31331,
         n31332, n31333, n31334, n31335, n31336, n31337, n31338, n31339,
         n31340, n31341, n31342, n31343, n31344, n31345, n31346, n31347,
         n31348, n31349, n31350, n31351, n31352, n31353, n31354, n31355,
         n31356, n31357, n31358, n31359, n31360, n31361, n31362, n31363,
         n31364, n31365, n31366, n31367, n31368, n31369, n31370, n31371,
         n31372, n31373, n31374, n31375, n31376, n31377, n31378, n31379,
         n31380, n31381, n31382, n31383, n31384, n31385, n31386, n31387,
         n31388, n31389, n31390, n31391, n31392, n31393, n31394, n31395,
         n31396, n31397, n31398, n31399, n31400, n31401, n31402, n31403,
         n31404, n31405, n31406, n31407, n31408, n31409, n31410, n31411,
         n31412, n31413, n31414, n31415, n31416, n31417, n31418, n31419,
         n31420, n31421, n31422, n31423, n31424, n31425, n31426, n31427,
         n31428, n31429, n31430, n31431, n31432, n31433, n31434, n31435,
         n31436, n31437, n31438, n31439, n31440, n31441, n31442, n31443,
         n31444, n31445, n31446, n31447, n31448, n31449, n31450, n31451,
         n31452, n31453, n31454, n31455, n31456, n31457, n31458, n31459,
         n31460, n31461, n31462, n31463, n31464, n31465, n31466, n31467,
         n31468, n31469, n31470, n31471, n31472, n31473, n31474, n31475,
         n31476, n31477, n31478, n31479, n31480, n31481, n31482, n31483,
         n31484, n31485, n31486, n31487, n31488, n31489, n31490, n31491,
         n31492, n31493, n31494, n31495, n31496, n31497, n31498, n31499,
         n31500, n31501, n31502, n31503, n31504, n31505, n31506, n31507,
         n31508, n31509, n31510, n31511, n31512, n31513, n31514, n31515,
         n31516, n31517, n31518, n31519, n31520, n31521, n31522, n31523,
         n31524, n31525, n31526, n31527, n31528, n31529, n31530, n31531,
         n31532, n31533, n31534, n31535, n31536, n31537, n31538, n31539,
         n31540, n31541, n31542, n31543, n31544, n31545, n31546, n31547,
         n31548, n31549, n31550, n31551, n31552, n31553, n31554, n31555,
         n31556, n31557, n31558, n31559, n31560, n31561, n31562, n31563,
         n31564, n31565, n31566, n31567, n31568, n31569, n31570, n31571,
         n31572, n31573, n31574, n31575, n31576, n31577, n31578, n31579,
         n31580, n31581, n31582, n31583, n31584, n31585, n31586, n31587,
         n31588, n31589, n31590, n31591, n31592, n31593, n31594, n31595,
         n31596, n31597, n31598, n31599, n31600, n31601, n31602, n31603,
         n31604, n31605, n31606, n31607, n31608, n31609, n31610, n31611,
         n31612, n31613, n31614, n31615, n31616, n31617, n31618, n31619,
         n31620, n31621, n31622, n31623, n31624, n31625, n31626, n31627,
         n31628, n31629, n31630, n31631, n31632, n31633, n31634, n31635,
         n31636, n31637, n31638, n31639, n31640, n31641, n31642, n31643,
         n31644, n31645, n31646, n31647, n31648, n31649, n31650, n31651,
         n31652, n31653, n31654, n31655, n31656, n31657, n31658, n31659,
         n31660, n31661, n31662, n31663, n31664, n31665, n31666, n31667,
         n31668, n31669, n31670, n31671, n31672, n31673, n31674, n31675,
         n31676, n31677, n31678, n31679, n31680, n31681, n31682, n31683,
         n31684, n31685, n31686, n31687, n31688, n31689, n31690, n31691,
         n31692, n31693, n31694, n31695, n31696, n31697, n31698, n31699,
         n31700, n31701, n31702, n31703, n31704, n31705, n31706, n31707,
         n31708, n31709, n31710, n31711, n31712, n31713, n31714, n31715,
         n31716, n31717, n31718, n31719, n31720, n31721, n31722, n31723,
         n31724, n31725, n31726, n31727, n31728, n31729, n31730, n31731,
         n31732, n31733, n31734, n31735, n31736, n31737, n31738, n31739,
         n31740, n31741, n31742, n31743, n31744, n31745, n31746, n31747,
         n31748, n31749, n31750, n31751, n31752, n31753, n31754, n31755,
         n31756, n31757, n31758, n31759, n31760, n31761, n31762, n31763,
         n31764, n31765, n31766, n31767, n31768, n31769, n31770, n31771,
         n31772, n31773, n31774, n31775, n31776, n31777, n31778, n31779,
         n31780, n31781, n31782, n31783, n31784, n31785, n31786, n31787,
         n31788, n31789, n31790, n31791, n31792, n31793, n31794, n31795,
         n31796, n31797, n31798, n31799, n31800, n31801, n31802, n31803,
         n31804, n31805, n31806, n31807, n31808, n31809, n31810, n31811,
         n31812, n31813, n31814, n31815, n31816, n31817, n31818, n31819,
         n31820, n31821, n31822, n31823, n31824, n31825, n31826, n31827,
         n31828, n31829, n31830, n31831, n31832, n31833, n31834, n31835,
         n31836, n31837, n31838, n31839, n31840, n31841, n31842, n31843,
         n31844, n31845, n31846, n31847, n31848, n31849, n31850, n31851,
         n31852, n31853, n31854, n31855, n31856, n31857, n31858, n31859,
         n31860, n31861, n31862, n31863, n31864, n31865, n31866, n31867,
         n31868, n31869, n31870, n31871, n31872, n31873, n31874, n31875,
         n31876, n31877, n31878, n31879, n31880, n31881, n31882, n31883,
         n31884, n31885, n31886, n31887, n31888, n31889, n31890, n31891,
         n31892, n31893, n31894, n31895, n31896, n31897, n31898, n31899,
         n31900, n31901, n31902, n31903, n31904, n31905, n31906, n31907,
         n31908, n31909, n31910, n31911, n31912, n31913, n31914, n31915,
         n31916, n31917, n31918, n31919, n31920, n31921, n31922, n31923,
         n31924, n31925, n31926, n31927, n31928, n31929, n31930, n31931,
         n31932, n31933, n31934, n31935, n31936, n31937, n31938, n31939,
         n31940, n31941, n31942, n31943, n31944, n31945, n31946, n31947,
         n31948, n31949, n31950, n31951, n31952, n31953, n31954, n31955,
         n31956, n31957, n31958, n31959, n31960, n31961, n31962, n31963,
         n31964, n31965, n31966, n31967, n31968, n31969, n31970, n31971,
         n31972, n31973, n31974, n31975, n31976, n31977, n31978, n31979,
         n31980, n31981, n31982, n31983, n31984, n31985, n31986, n31987,
         n31988, n31989, n31990, n31991, n31992, n31993, n31994, n31995,
         n31996, n31997, n31998, n31999, n32000, n32001, n32002, n32003,
         n32004, n32005, n32006, n32007, n32008, n32009, n32010, n32011,
         n32012, n32013, n32014, n32015, n32016, n32017, n32018, n32019,
         n32020, n32021, n32022, n32023, n32024, n32025, n32026, n32027,
         n32028, n32029, n32030, n32031, n32032, n32033, n32034, n32035,
         n32036, n32037, n32038, n32039, n32040, n32041, n32042, n32043,
         n32044, n32045, n32046, n32047, n32048, n32049, n32050, n32051,
         n32052, n32053, n32054, n32055, n32056, n32057, n32058, n32059,
         n32060, n32061, n32062, n32063, n32064, n32065, n32066, n32067,
         n32068, n32069, n32070, n32071, n32072, n32073, n32074, n32075,
         n32076, n32077, n32078, n32079, n32080, n32081, n32082, n32083,
         n32084, n32085, n32086, n32087, n32088, n32089, n32090, n32091,
         n32092, n32093, n32094, n32095, n32096, n32097, n32098, n32099,
         n32100, n32101, n32102, n32103, n32104, n32105, n32106, n32107,
         n32108, n32109, n32110, n32111, n32112, n32113, n32114, n32115,
         n32116, n32117, n32118, n32119, n32120, n32121, n32122, n32123,
         n32124, n32125, n32126, n32127, n32128, n32129, n32130, n32131,
         n32132, n32133, n32134, n32135, n32136, n32137, n32138, n32139,
         n32140, n32141, n32142, n32143, n32144, n32145, n32146, n32147,
         n32148, n32149, n32150, n32151, n32152, n32153, n32154, n32155,
         n32156, n32157, n32158, n32159, n32160, n32161, n32162, n32163,
         n32164, n32165, n32166, n32167, n32168, n32169, n32170, n32171,
         n32172, n32173, n32174, n32175, n32176, n32177, n32178, n32179,
         n32180, n32181, n32182, n32183, n32184, n32185, n32186, n32187,
         n32188, n32189, n32190, n32191, n32192, n32193, n32194, n32195,
         n32196, n32197, n32198, n32199, n32200, n32201, n32202, n32203,
         n32204, n32205, n32206, n32207, n32208, n32209, n32210, n32211,
         n32212, n32213, n32214, n32215, n32216, n32217, n32218, n32219,
         n32220, n32221, n32222, n32223, n32224, n32225, n32226, n32227,
         n32228, n32229, n32230, n32231, n32232, n32233, n32234, n32235,
         n32236, n32237, n32238, n32239, n32240, n32241, n32242, n32243,
         n32244, n32245, n32246, n32247, n32248, n32249, n32250, n32251,
         n32252, n32253, n32254, n32255, n32256, n32257, n32258, n32259,
         n32260, n32261, n32262, n32263, n32264, n32265, n32266, n32267,
         n32268, n32269, n32270, n32271, n32272, n32273, n32274, n32275,
         n32276, n32277, n32278, n32279, n32280, n32281, n32282, n32283,
         n32284, n32285, n32286, n32287, n32288, n32289, n32290, n32291,
         n32292, n32293, n32294, n32295, n32296, n32297, n32298, n32299,
         n32300, n32301, n32302, n32303, n32304, n32305, n32306, n32307,
         n32308, n32309, n32310, n32311, n32312, n32313, n32314, n32315,
         n32316, n32317, n32318, n32319, n32320, n32321, n32322, n32323,
         n32324, n32325, n32326, n32327, n32328, n32329, n32330, n32331,
         n32332, n32333, n32334, n32335, n32336, n32337, n32338, n32339,
         n32340, n32341, n32342, n32343, n32344, n32345, n32346, n32347,
         n32348, n32349, n32350, n32351, n32352, n32353, n32354, n32355,
         n32356, n32357, n32358, n32359, n32360, n32361, n32362, n32363,
         n32364, n32365, n32366, n32367, n32368, n32369, n32370, n32371,
         n32372, n32373, n32374, n32375, n32376, n32377, n32378, n32379,
         n32380, n32381, n32382, n32383, n32384, n32385, n32386, n32387,
         n32388, n32389, n32390, n32391, n32392, n32393, n32394, n32395,
         n32396, n32397, n32398, n32399, n32400, n32401, n32402, n32403,
         n32404, n32405, n32406, n32407, n32408, n32409, n32410, n32411,
         n32412, n32413, n32414, n32415, n32416, n32417, n32418, n32419,
         n32420, n32421, n32422, n32423, n32424, n32425, n32426, n32427,
         n32428, n32429, n32430, n32431, n32432, n32433, n32434, n32435,
         n32436, n32437, n32438, n32439, n32440, n32441, n32442, n32443,
         n32444, n32445, n32446, n32447, n32448, n32449, n32450, n32451,
         n32452, n32453, n32454, n32455, n32456, n32457, n32458, n32459,
         n32460, n32461, n32462, n32463, n32464, n32465, n32466, n32467,
         n32468, n32469, n32470, n32471, n32472, n32473, n32474, n32475,
         n32476, n32477, n32478, n32479, n32480, n32481, n32482, n32483,
         n32484, n32485, n32486, n32487, n32488, n32489, n32490, n32491,
         n32492, n32493, n32494, n32495, n32496, n32497, n32498, n32499,
         n32500, n32501, n32502, n32503, n32504, n32505, n32506, n32507,
         n32508, n32509, n32510, n32511, n32512, n32513, n32514, n32515,
         n32516, n32517, n32518, n32519, n32520, n32521, n32522, n32523,
         n32524, n32525, n32526, n32527, n32528, n32529, n32530, n32531,
         n32532, n32533, n32534, n32535, n32536, n32537, n32538, n32539,
         n32540, n32541, n32542, n32543, n32544, n32545, n32546, n32547,
         n32548, n32549, n32550, n32551, n32552, n32553, n32554, n32555,
         n32556, n32557, n32558, n32559, n32560, n32561, n32562, n32563,
         n32564, n32565, n32566, n32567, n32568, n32569, n32570, n32571,
         n32572, n32573, n32574, n32575, n32576, n32577, n32578, n32579,
         n32580, n32581, n32582, n32583, n32584, n32585, n32586, n32587,
         n32588, n32589, n32590, n32591, n32592, n32593, n32594, n32595,
         n32596, n32597, n32598, n32599, n32600, n32601, n32602, n32603,
         n32604, n32605, n32606, n32607, n32608, n32609, n32610, n32611,
         n32612, n32613, n32614, n32615, n32616, n32617, n32618, n32619,
         n32620, n32621, n32622, n32623, n32624, n32625, n32626, n32627,
         n32628, n32629, n32630, n32631, n32632, n32633, n32634, n32635,
         n32636, n32637, n32638, n32639, n32640, n32641, n32642, n32643,
         n32644, n32645, n32646, n32647, n32648, n32649, n32650, n32651,
         n32652, n32653, n32654, n32655, n32656, n32657, n32658, n32659,
         n32660, n32661, n32662, n32663, n32664, n32665, n32666, n32667,
         n32668, n32669, n32670, n32671, n32672, n32673, n32674, n32675,
         n32676, n32677, n32678, n32679, n32680, n32681, n32682, n32683,
         n32684, n32685, n32686, n32687, n32688, n32689, n32690, n32691,
         n32692, n32693, n32694, n32695, n32696, n32697, n32698, n32699,
         n32700, n32701, n32702, n32703, n32704, n32705, n32706, n32707,
         n32708, n32709, n32710, n32711, n32712, n32713, n32714, n32715,
         n32716, n32717, n32718, n32719, n32720, n32721, n32722, n32723,
         n32724, n32725, n32726, n32727, n32728, n32729, n32730, n32731,
         n32732, n32733, n32734, n32735, n32736, n32737, n32738, n32739,
         n32740, n32741, n32742, n32743, n32744, n32745, n32746, n32747,
         n32748, n32749, n32750, n32751, n32752, n32753, n32754, n32755,
         n32756, n32757, n32758, n32759, n32760, n32761, n32762, n32763,
         n32764, n32765, n32766, n32767, n32768, n32769, n32770, n32771,
         n32772, n32773, n32774, n32775, n32776, n32777, n32778, n32779,
         n32780, n32781, n32782, n32783, n32784, n32785, n32786, n32787,
         n32788, n32789, n32790, n32791, n32792, n32793, n32794, n32795,
         n32796, n32797, n32798, n32799, n32800, n32801, n32802, n32803,
         n32804, n32805, n32806, n32807, n32808, n32809, n32810, n32811,
         n32812, n32813, n32814, n32815, n32816, n32817, n32818, n32819,
         n32820, n32821, n32822, n32823, n32824, n32825, n32826, n32827,
         n32828, n32829, n32830, n32831, n32832, n32833, n32834, n32835,
         n32836, n32837, n32838, n32839, n32840, n32841, n32842, n32843,
         n32844, n32845, n32846, n32847, n32848, n32849, n32850, n32851,
         n32852, n32853, n32854, n32855, n32856, n32857, n32858, n32859,
         n32860, n32861, n32862, n32863, n32864, n32865, n32866, n32867,
         n32868, n32869, n32870, n32871, n32872, n32873, n32874, n32875,
         n32876, n32877, n32878, n32879, n32880, n32881, n32882, n32883,
         n32884, n32885, n32886, n32887, n32888, n32889, n32890, n32891,
         n32892, n32893, n32894, n32895, n32896, n32897, n32898, n32899,
         n32900, n32901, n32902, n32903, n32904, n32905, n32906, n32907,
         n32908, n32909, n32910, n32911, n32912, n32913, n32914, n32915,
         n32916, n32917, n32918, n32919, n32920, n32921, n32922, n32923,
         n32924, n32925, n32926, n32927, n32928, n32929, n32930, n32931,
         n32932, n32933, n32934, n32935, n32936, n32937, n32938, n32939,
         n32940, n32941, n32942, n32943, n32944, n32945, n32946, n32947,
         n32948, n32949, n32950, n32951, n32952, n32953, n32954, n32955,
         n32956, n32957, n32958, n32959, n32960, n32961, n32962, n32963,
         n32964, n32965, n32966, n32967, n32968, n32969, n32970, n32971,
         n32972, n32973, n32974, n32975, n32976, n32977, n32978, n32979,
         n32980, n32981, n32982, n32983, n32984, n32985, n32986, n32987,
         n32988, n32989, n32990, n32991, n32992, n32993, n32994, n32995,
         n32996, n32997, n32998, n32999, n33000, n33001, n33002, n33003,
         n33004, n33005, n33006, n33007, n33008, n33009, n33010, n33011,
         n33012, n33013, n33014, n33015, n33016, n33017, n33018, n33019,
         n33020, n33021, n33022, n33023, n33024, n33025, n33026, n33027,
         n33028, n33029, n33030, n33031, n33032, n33033, n33034, n33035,
         n33036, n33037, n33038, n33039, n33040, n33041, n33042, n33043,
         n33044, n33045, n33046, n33047, n33048, n33049, n33050, n33051,
         n33052, n33053, n33054, n33055, n33056, n33057, n33058, n33059,
         n33060, n33061, n33062, n33063, n33064, n33065, n33066, n33067,
         n33068, n33069, n33070, n33071, n33072, n33073, n33074, n33075,
         n33076, n33077, n33078, n33079, n33080, n33081, n33082, n33083,
         n33084, n33085, n33086, n33087, n33088, n33089, n33090, n33091,
         n33092, n33093, n33094, n33095, n33096, n33097, n33098, n33099,
         n33100, n33101, n33102, n33103, n33104, n33105, n33106, n33107,
         n33108, n33109, n33110, n33111, n33112, n33113, n33114, n33115,
         n33116, n33117, n33118, n33119, n33120, n33121, n33122, n33123,
         n33124, n33125, n33126, n33127, n33128, n33129, n33130, n33131,
         n33132, n33133, n33134, n33135, n33136, n33137, n33138, n33139,
         n33140, n33141, n33142, n33143, n33144, n33145, n33146, n33147,
         n33148, n33149, n33150, n33151, n33152, n33153, n33154, n33155,
         n33156, n33157, n33158, n33159, n33160, n33161, n33162, n33163,
         n33164, n33165, n33166, n33167, n33168, n33169, n33170, n33171,
         n33172, n33173, n33174, n33175, n33176, n33177, n33178, n33179,
         n33180, n33181, n33182, n33183, n33184, n33185, n33186, n33187,
         n33188, n33189, n33190, n33191, n33192, n33193, n33194, n33195,
         n33196, n33197, n33198, n33199, n33200, n33201, n33202, n33203,
         n33204, n33205, n33206, n33207, n33208, n33209, n33210, n33211,
         n33212, n33213, n33214, n33215, n33216, n33217, n33218, n33219,
         n33220, n33221, n33222, n33223, n33224, n33225, n33226, n33227,
         n33228, n33229, n33230, n33231, n33232, n33233, n33234, n33235,
         n33236, n33237, n33238, n33239, n33240, n33241, n33242, n33243,
         n33244, n33245, n33246, n33247, n33248, n33249, n33250, n33251,
         n33252, n33253, n33254, n33255, n33256, n33257, n33258, n33259,
         n33260, n33261, n33262, n33263, n33264, n33265, n33266, n33267,
         n33268, n33269, n33270, n33271, n33272, n33273, n33274, n33275,
         n33276, n33277, n33278, n33279, n33280, n33281, n33282, n33283,
         n33284, n33285, n33286, n33287, n33288, n33289, n33290, n33291,
         n33292, n33293, n33294, n33295, n33296, n33297, n33298, n33299,
         n33300, n33301, n33302, n33303, n33304, n33305, n33306, n33307,
         n33308, n33309, n33310, n33311, n33312, n33313, n33314, n33315,
         n33316, n33317, n33318, n33319, n33320, n33321, n33322, n33323,
         n33324, n33325, n33326, n33327, n33328, n33329, n33330, n33331,
         n33332, n33333, n33334, n33335, n33336, n33337, n33338, n33339,
         n33340, n33341, n33342, n33343, n33344, n33345, n33346, n33347,
         n33348, n33349, n33350, n33351, n33352, n33353, n33354, n33355,
         n33356, n33357, n33358, n33359, n33360, n33361, n33362, n33363,
         n33364, n33365, n33366, n33367, n33368, n33369, n33370, n33371,
         n33372, n33373, n33374, n33375, n33376, n33377, n33378, n33379,
         n33380, n33381, n33382, n33383, n33384, n33385, n33386, n33387,
         n33388, n33389, n33390, n33391, n33392, n33393, n33394, n33395,
         n33396, n33397, n33398, n33399, n33400, n33401, n33402, n33403,
         n33404, n33405, n33406, n33407, n33408, n33409, n33410, n33411,
         n33412, n33413, n33414, n33415, n33416, n33417, n33418, n33419,
         n33420, n33421, n33422, n33423, n33424, n33425, n33426, n33427,
         n33428, n33429, n33430, n33431, n33432, n33433, n33434, n33435,
         n33436, n33437, n33438, n33439, n33440, n33441, n33442, n33443,
         n33444, n33445, n33446, n33447, n33448, n33449, n33450, n33451,
         n33452, n33453, n33454, n33455, n33456, n33457, n33458, n33459,
         n33460, n33461, n33462, n33463, n33464, n33465, n33466, n33467,
         n33468, n33469, n33470, n33471, n33472, n33473, n33474, n33475,
         n33476, n33477, n33478, n33479, n33480, n33481, n33482, n33483,
         n33484, n33485, n33486, n33487, n33488, n33489, n33490, n33491,
         n33492, n33493, n33494, n33495, n33496, n33497, n33498, n33499,
         n33500, n33501, n33502, n33503, n33504, n33505, n33506, n33507,
         n33508, n33509, n33510, n33511, n33512, n33513, n33514, n33515,
         n33516, n33517, n33518, n33519, n33520, n33521, n33522, n33523,
         n33524, n33525, n33526, n33527, n33528, n33529, n33530, n33531,
         n33532, n33533, n33534, n33535, n33536, n33537, n33538, n33539,
         n33540, n33541, n33542, n33543, n33544, n33545, n33546, n33547,
         n33548, n33549, n33550, n33551, n33552, n33553, n33554, n33555,
         n33556, n33557, n33558, n33559, n33560, n33561, n33562, n33563,
         n33564, n33565, n33566, n33567, n33568, n33569, n33570, n33571,
         n33572, n33573, n33574, n33575, n33576, n33577, n33578, n33579,
         n33580, n33581, n33582, n33583, n33584, n33585, n33586, n33587,
         n33588, n33589, n33590, n33591, n33592, n33593, n33594, n33595,
         n33596, n33597, n33598, n33599, n33600, n33601, n33602, n33603,
         n33604, n33605, n33606, n33607, n33608, n33609, n33610, n33611,
         n33612, n33613, n33614, n33615, n33616, n33617, n33618, n33619,
         n33620, n33621, n33622, n33623, n33624, n33625, n33626, n33627,
         n33628, n33629, n33630, n33631, n33632, n33633, n33634, n33635,
         n33636, n33637, n33638, n33639, n33640, n33641, n33642, n33643,
         n33644, n33645, n33646, n33647, n33648, n33649, n33650, n33651,
         n33652, n33653, n33654, n33655, n33656, n33657, n33658, n33659,
         n33660, n33661, n33662, n33663, n33664, n33665, n33666, n33667,
         n33668, n33669, n33670, n33671, n33672, n33673, n33674, n33675,
         n33676, n33677, n33678, n33679, n33680, n33681, n33682, n33683,
         n33684, n33685, n33686, n33687, n33688, n33689, n33690, n33691,
         n33692, n33693, n33694, n33695, n33696, n33697, n33698, n33699,
         n33700, n33701, n33702, n33703, n33704, n33705, n33706, n33707,
         n33708, n33709, n33710, n33711, n33712, n33713, n33714, n33715,
         n33716, n33717, n33718, n33719, n33720, n33721, n33722, n33723,
         n33724, n33725, n33726, n33727, n33728, n33729, n33730, n33731,
         n33732, n33733, n33734, n33735, n33736, n33737, n33738, n33739,
         n33740, n33741, n33742, n33743, n33744, n33745, n33746, n33747,
         n33748, n33749, n33750, n33751, n33752, n33753, n33754, n33755,
         n33756, n33757, n33758, n33759, n33760, n33761, n33762, n33763,
         n33764, n33765, n33766, n33767, n33768, n33769, n33770, n33771,
         n33772, n33773, n33774, n33775, n33776, n33777, n33778, n33779,
         n33780, n33781, n33782, n33783, n33784, n33785, n33786, n33787,
         n33788, n33789, n33790, n33791, n33792, n33793, n33794, n33795,
         n33796, n33797, n33798, n33799, n33800, n33801, n33802, n33803,
         n33804, n33805, n33806, n33807, n33808, n33809, n33810, n33811,
         n33812, n33813, n33814, n33815, n33816, n33817, n33818, n33819,
         n33820, n33821, n33822, n33823, n33824, n33825, n33826, n33827,
         n33828, n33829, n33830, n33831, n33832, n33833, n33834, n33835,
         n33836, n33837, n33838, n33839, n33840, n33841, n33842, n33843,
         n33844, n33845, n33846, n33847, n33848, n33849, n33850, n33851,
         n33852, n33853, n33854, n33855, n33856, n33857, n33858, n33859,
         n33860, n33861, n33862, n33863, n33864, n33865, n33866, n33867,
         n33868, n33869, n33870, n33871, n33872, n33873, n33874, n33875,
         n33876, n33877, n33878, n33879, n33880, n33881, n33882, n33883,
         n33884, n33885, n33886, n33887, n33888, n33889, n33890, n33891,
         n33892, n33893, n33894, n33895, n33896, n33897, n33898, n33899,
         n33900, n33901, n33902, n33903, n33904, n33905, n33906, n33907,
         n33908, n33909, n33910, n33911, n33912, n33913, n33914, n33915,
         n33916, n33917, n33918, n33919, n33920, n33921, n33922, n33923,
         n33924, n33925, n33926, n33927, n33928, n33929, n33930, n33931,
         n33932, n33933, n33934, n33935, n33936, n33937, n33938, n33939,
         n33940, n33941, n33942, n33943, n33944, n33945, n33946, n33947,
         n33948, n33949, n33950, n33951, n33952, n33953, n33954, n33955,
         n33956, n33957, n33958, n33959, n33960, n33961, n33962, n33963,
         n33964, n33965, n33966, n33967, n33968, n33969, n33970, n33971,
         n33972, n33973, n33974, n33975, n33976, n33977, n33978, n33979,
         n33980, n33981, n33982, n33983, n33984, n33985, n33986, n33987,
         n33988, n33989, n33990, n33991, n33992, n33993, n33994, n33995,
         n33996, n33997, n33998, n33999, n34000, n34001, n34002, n34003,
         n34004, n34005, n34006, n34007, n34008, n34009, n34010, n34011,
         n34012, n34013, n34014, n34015, n34016, n34017, n34018, n34019,
         n34020, n34021, n34022, n34023, n34024, n34025, n34026, n34027,
         n34028, n34029, n34030, n34031, n34032, n34033, n34034, n34035,
         n34036, n34037, n34038, n34039, n34040, n34041, n34042, n34043,
         n34044, n34045, n34046, n34047, n34048, n34049, n34050, n34051,
         n34052, n34053, n34054, n34055, n34056, n34057, n34058, n34059,
         n34060, n34061, n34062, n34063, n34064, n34065, n34066, n34067,
         n34068, n34069, n34070, n34071, n34072, n34073, n34074, n34075,
         n34076, n34077, n34078, n34079, n34080, n34081, n34082, n34083,
         n34084, n34085, n34086, n34087, n34088, n34089, n34090, n34091,
         n34092, n34093, n34094, n34095, n34096, n34097, n34098, n34099,
         n34100, n34101, n34102, n34103, n34104, n34105, n34106, n34107,
         n34108, n34109, n34110, n34111, n34112, n34113, n34114, n34115,
         n34116, n34117, n34118, n34119, n34120, n34121, n34122, n34123,
         n34124, n34125, n34126, n34127, n34128, n34129, n34130, n34131,
         n34132, n34133, n34134, n34135, n34136, n34137, n34138, n34139,
         n34140, n34141, n34142, n34143, n34144, n34145, n34146, n34147,
         n34148, n34149, n34150, n34151, n34152, n34153, n34154, n34155,
         n34156, n34157, n34158, n34159, n34160, n34161, n34162, n34163,
         n34164, n34165, n34166, n34167, n34168, n34169, n34170, n34171,
         n34172, n34173, n34174, n34175, n34176, n34177, n34178, n34179,
         n34180, n34181, n34182, n34183, n34184, n34185, n34186, n34187,
         n34188, n34189, n34190, n34191, n34192, n34193, n34194, n34195,
         n34196, n34197, n34198, n34199, n34200, n34201, n34202, n34203,
         n34204, n34205, n34206, n34207, n34208, n34209, n34210, n34211,
         n34212, n34213, n34214, n34215, n34216, n34217, n34218, n34219,
         n34220, n34221, n34222, n34223, n34224, n34225, n34226, n34227,
         n34228, n34229, n34230, n34231, n34232, n34233, n34234, n34235,
         n34236, n34237, n34238, n34239, n34240, n34241, n34242, n34243,
         n34244, n34245, n34246, n34247, n34248, n34249, n34250, n34251,
         n34252, n34253, n34254, n34255, n34256, n34257, n34258, n34259,
         n34260, n34261, n34262, n34263, n34264, n34265, n34266, n34267,
         n34268, n34269, n34270, n34271, n34272, n34273, n34274, n34275,
         n34276, n34277, n34278, n34279, n34280, n34281, n34282, n34283,
         n34284, n34285, n34286, n34287, n34288, n34289, n34290, n34291,
         n34292, n34293, n34294, n34295, n34296, n34297, n34298, n34299,
         n34300, n34301, n34302, n34303, n34304, n34305, n34306, n34307,
         n34308, n34309, n34310, n34311, n34312, n34313, n34314, n34315,
         n34316, n34317, n34318, n34319, n34320, n34321, n34322, n34323,
         n34324, n34325, n34326, n34327, n34328, n34329, n34330, n34331,
         n34332, n34333, n34334, n34335, n34336, n34337, n34338, n34339,
         n34340, n34341, n34342, n34343, n34344, n34345, n34346, n34347,
         n34348, n34349, n34350, n34351, n34352, n34353, n34354, n34355,
         n34356, n34357, n34358, n34359, n34360, n34361, n34362, n34363,
         n34364, n34365, n34366, n34367, n34368, n34369, n34370, n34371,
         n34372, n34373, n34374, n34375, n34376, n34377, n34378, n34379,
         n34380, n34381, n34382, n34383, n34384, n34385, n34386, n34387,
         n34388, n34389, n34390, n34391, n34392, n34393, n34394, n34395,
         n34396, n34397, n34398, n34399, n34400, n34401, n34402, n34403,
         n34404, n34405, n34406, n34407, n34408, n34409, n34410, n34411,
         n34412, n34413, n34414, n34415, n34416, n34417, n34418, n34419,
         n34420, n34421, n34422, n34423, n34424, n34425, n34426, n34427,
         n34428, n34429, n34430, n34431, n34432, n34433, n34434, n34435,
         n34436, n34437, n34438, n34439, n34440, n34441, n34442, n34443,
         n34444, n34445, n34446, n34447, n34448, n34449, n34450, n34451,
         n34452, n34453, n34454, n34455, n34456, n34457, n34458, n34459,
         n34460, n34461, n34462, n34463, n34464, n34465, n34466, n34467,
         n34468, n34469, n34470, n34471, n34472, n34473, n34474, n34475,
         n34476, n34477, n34478, n34479, n34480, n34481, n34482, n34483,
         n34484, n34485, n34486, n34487, n34488, n34489, n34490, n34491,
         n34492, n34493, n34494, n34495, n34496, n34497, n34498, n34499,
         n34500, n34501, n34502, n34503, n34504, n34505, n34506, n34507,
         n34508, n34509, n34510, n34511, n34512, n34513, n34514, n34515,
         n34516, n34517, n34518, n34519, n34520, n34521, n34522, n34523,
         n34524, n34525, n34526, n34527, n34528, n34529, n34530, n34531,
         n34532, n34533, n34534, n34535, n34536, n34537, n34538, n34539,
         n34540, n34541, n34542, n34543, n34544, n34545, n34546, n34547,
         n34548, n34549, n34550, n34551, n34552, n34553, n34554, n34555,
         n34556, n34557, n34558, n34559, n34560, n34561, n34562, n34563,
         n34564, n34565, n34566, n34567, n34568, n34569, n34570, n34571,
         n34572, n34573, n34574, n34575, n34576, n34577, n34578, n34579,
         n34580, n34581, n34582, n34583, n34584, n34585, n34586, n34587,
         n34588, n34589, n34590, n34591, n34592, n34593, n34594, n34595,
         n34596, n34597, n34598, n34599, n34600, n34601, n34602, n34603,
         n34604, n34605, n34606, n34607, n34608, n34609, n34610, n34611,
         n34612, n34613, n34614, n34615, n34616, n34617, n34618, n34619,
         n34620, n34621, n34622, n34623, n34624, n34625, n34626, n34627,
         n34628, n34629, n34630, n34631, n34632, n34633, n34634, n34635,
         n34636, n34637, n34638, n34639, n34640, n34641, n34642, n34643,
         n34644, n34645, n34646, n34647, n34648, n34649, n34650, n34651,
         n34652, n34653, n34654, n34655, n34656, n34657, n34658, n34659,
         n34660, n34661, n34662, n34663, n34664, n34665, n34666, n34667,
         n34668, n34669, n34670, n34671, n34672, n34673, n34674, n34675,
         n34676, n34677, n34678, n34679, n34680, n34681, n34682, n34683,
         n34684, n34685, n34686, n34687, n34688, n34689, n34690, n34691,
         n34692, n34693, n34694, n34695, n34696, n34697, n34698, n34699,
         n34700, n34701, n34702, n34703, n34704, n34705, n34706, n34707,
         n34708, n34709, n34710, n34711, n34712, n34713, n34714, n34715,
         n34716, n34717, n34718, n34719, n34720, n34721, n34722, n34723,
         n34724, n34725, n34726, n34727, n34728, n34729, n34730, n34731,
         n34732, n34733, n34734, n34735, n34736, n34737, n34738, n34739,
         n34740, n34741, n34742, n34743, n34744, n34745, n34746, n34747,
         n34748, n34749, n34750, n34751, n34752, n34753, n34754, n34755,
         n34756, n34757, n34758, n34759, n34760, n34761, n34762, n34763,
         n34764, n34765, n34766, n34767, n34768, n34769, n34770, n34771,
         n34772, n34773, n34774, n34775, n34776, n34777, n34778, n34779,
         n34780, n34781, n34782, n34783, n34784, n34785, n34786, n34787,
         n34788, n34789, n34790, n34791, n34792, n34793, n34794, n34795,
         n34796, n34797, n34798, n34799, n34800, n34801, n34802, n34803,
         n34804, n34805, n34806, n34807, n34808, n34809, n34810, n34811,
         n34812, n34813, n34814, n34815, n34816, n34817, n34818, n34819,
         n34820, n34821, n34822, n34823, n34824, n34825, n34826, n34827,
         n34828, n34829, n34830, n34831, n34832, n34833, n34834, n34835,
         n34836, n34837, n34838, n34839, n34840, n34841, n34842, n34843,
         n34844, n34845, n34846, n34847, n34848, n34849, n34850, n34851,
         n34852, n34853, n34854, n34855, n34856, n34857, n34858, n34859,
         n34860, n34861, n34862, n34863, n34864, n34865, n34866, n34867,
         n34868, n34869, n34870, n34871, n34872, n34873, n34874, n34875,
         n34876, n34877, n34878, n34879, n34880, n34881, n34882, n34883,
         n34884, n34885, n34886, n34887, n34888, n34889, n34890, n34891,
         n34892, n34893, n34894, n34895, n34896, n34897, n34898, n34899,
         n34900, n34901, n34902, n34903, n34904, n34905, n34906, n34907,
         n34908, n34909, n34910, n34911, n34912, n34913, n34914, n34915,
         n34916, n34917, n34918, n34919, n34920, n34921, n34922, n34923,
         n34924, n34925, n34926, n34927, n34928, n34929, n34930, n34931,
         n34932, n34933, n34934, n34935, n34936, n34937, n34938, n34939,
         n34940, n34941, n34942, n34943, n34944, n34945, n34946, n34947,
         n34948, n34949, n34950, n34951, n34952, n34953, n34954, n34955,
         n34956, n34957, n34958, n34959, n34960, n34961, n34962, n34963,
         n34964, n34965, n34966, n34967, n34968, n34969, n34970, n34971,
         n34972, n34973, n34974, n34975, n34976, n34977, n34978, n34979,
         n34980, n34981, n34982, n34983, n34984, n34985, n34986, n34987,
         n34988, n34989, n34990, n34991, n34992, n34993, n34994, n34995,
         n34996, n34997, n34998, n34999, n35000, n35001, n35002, n35003,
         n35004, n35005, n35006, n35007, n35008, n35009, n35010, n35011,
         n35012, n35013, n35014, n35015, n35016, n35017, n35018, n35019,
         n35020, n35021, n35022, n35023, n35024, n35025, n35026, n35027,
         n35028, n35029, n35030, n35031, n35032, n35033, n35034, n35035,
         n35036, n35037, n35038, n35039, n35040, n35041, n35042, n35043,
         n35044, n35045, n35046, n35047, n35048, n35049, n35050, n35051,
         n35052, n35053, n35054, n35055, n35056, n35057, n35058, n35059,
         n35060, n35061, n35062, n35063, n35064, n35065, n35066, n35067,
         n35068, n35069, n35070, n35071, n35072, n35073, n35074, n35075,
         n35076, n35077, n35078, n35079, n35080, n35081, n35082, n35083,
         n35084, n35085, n35086, n35087, n35088, n35089, n35090, n35091,
         n35092, n35093, n35094, n35095, n35096, n35097, n35098, n35099,
         n35100, n35101, n35102, n35103, n35104, n35105, n35106, n35107,
         n35108, n35109, n35110, n35111, n35112, n35113, n35114, n35115,
         n35116, n35117, n35118, n35119, n35120, n35121, n35122, n35123,
         n35124, n35125, n35126, n35127, n35128, n35129, n35130, n35131,
         n35132, n35133, n35134, n35135, n35136, n35137, n35138, n35139,
         n35140, n35141, n35142, n35143, n35144, n35145, n35146, n35147,
         n35148, n35149, n35150, n35151, n35152, n35153, n35154, n35155,
         n35156, n35157, n35158, n35159, n35160, n35161, n35162, n35163,
         n35164, n35165, n35166, n35167, n35168, n35169, n35170, n35171,
         n35172, n35173, n35174, n35175, n35176, n35177, n35178, n35179,
         n35180, n35181, n35182, n35183, n35184, n35185, n35186, n35187,
         n35188, n35189, n35190, n35191, n35192, n35193, n35194, n35195,
         n35196, n35197, n35198, n35199, n35200, n35201, n35202, n35203,
         n35204, n35205, n35206, n35207, n35208, n35209, n35210, n35211,
         n35212, n35213, n35214, n35215, n35216, n35217, n35218, n35219,
         n35220, n35221, n35222, n35223, n35224, n35225, n35226, n35227,
         n35228, n35229, n35230, n35231, n35232, n35233, n35234, n35235,
         n35236, n35237, n35238, n35239, n35240, n35241, n35242, n35243,
         n35244, n35245, n35246, n35247, n35248, n35249, n35250, n35251,
         n35252, n35253, n35254, n35255, n35256, n35257, n35258, n35259,
         n35260, n35261, n35262, n35263, n35264, n35265, n35266, n35267,
         n35268, n35269, n35270, n35271, n35272, n35273, n35274, n35275,
         n35276, n35277, n35278, n35279, n35280, n35281, n35282, n35283,
         n35284, n35285, n35286, n35287, n35288, n35289, n35290, n35291,
         n35292, n35293, n35294, n35295, n35296, n35297, n35298, n35299,
         n35300, n35301, n35302, n35303, n35304, n35305, n35306, n35307,
         n35308, n35309, n35310, n35311, n35312, n35313, n35314, n35315,
         n35316, n35317, n35318, n35319, n35320, n35321, n35322, n35323,
         n35324, n35325, n35326, n35327, n35328, n35329, n35330, n35331,
         n35332, n35333, n35334, n35335, n35336, n35337, n35338, n35339,
         n35340, n35341, n35342, n35343, n35344, n35345, n35346, n35347,
         n35348, n35349, n35350, n35351, n35352, n35353, n35354, n35355,
         n35356, n35357, n35358, n35359, n35360, n35361, n35362, n35363,
         n35364, n35365, n35366, n35367, n35368, n35369, n35370, n35371,
         n35372, n35373, n35374, n35375, n35376, n35377, n35378, n35379,
         n35380, n35381, n35382, n35383, n35384, n35385, n35386, n35387,
         n35388, n35389, n35390, n35391, n35392, n35393, n35394, n35395,
         n35396, n35397, n35398, n35399, n35400, n35401, n35402, n35403,
         n35404, n35405, n35406, n35407, n35408, n35409, n35410, n35411,
         n35412, n35413, n35414, n35415, n35416, n35417, n35418, n35419,
         n35420, n35421, n35422, n35423, n35424, n35425, n35426, n35427,
         n35428, n35429, n35430, n35431, n35432, n35433, n35434, n35435,
         n35436, n35437, n35438, n35439, n35440, n35441, n35442, n35443,
         n35444, n35445, n35446, n35447, n35448, n35449, n35450, n35451,
         n35452, n35453, n35454, n35455, n35456, n35457, n35458, n35459,
         n35460, n35461, n35462, n35463, n35464, n35465, n35466, n35467,
         n35468, n35469, n35470, n35471, n35472, n35473, n35474, n35475,
         n35476, n35477, n35478, n35479, n35480, n35481, n35482, n35483,
         n35484, n35485, n35486, n35487, n35488, n35489, n35490, n35491,
         n35492, n35493, n35494, n35495, n35496, n35497, n35498, n35499,
         n35500, n35501, n35502, n35503, n35504, n35505, n35506, n35507,
         n35508, n35509, n35510, n35511, n35512, n35513, n35514, n35515,
         n35516, n35517, n35518, n35519, n35520, n35521, n35522, n35523,
         n35524, n35525, n35526, n35527, n35528, n35529, n35530, n35531,
         n35532, n35533, n35534, n35535, n35536, n35537, n35538, n35539,
         n35540, n35541, n35542, n35543, n35544, n35545, n35546, n35547,
         n35548, n35549, n35550, n35551, n35552, n35553, n35554, n35555,
         n35556, n35557, n35558, n35559, n35560, n35561, n35562, n35563,
         n35564, n35565, n35566, n35567, n35568, n35569, n35570, n35571,
         n35572, n35573, n35574, n35575, n35576, n35577, n35578, n35579,
         n35580, n35581, n35582, n35583, n35584, n35585, n35586, n35587,
         n35588, n35589, n35590, n35591, n35592, n35593, n35594, n35595,
         n35596, n35597, n35598, n35599, n35600, n35601, n35602, n35603,
         n35604, n35605, n35606, n35607, n35608, n35609, n35610, n35611,
         n35612, n35613, n35614, n35615, n35616, n35617, n35618, n35619,
         n35620, n35621, n35622, n35623, n35624, n35625, n35626, n35627,
         n35628, n35629, n35630, n35631, n35632, n35633, n35634, n35635,
         n35636, n35637, n35638, n35639, n35640, n35641, n35642, n35643,
         n35644, n35645, n35646, n35647, n35648, n35649, n35650, n35651,
         n35652, n35653, n35654, n35655, n35656, n35657, n35658, n35659,
         n35660, n35661, n35662, n35663, n35664, n35665, n35666, n35667,
         n35668, n35669, n35670, n35671, n35672, n35673, n35674, n35675,
         n35676, n35677, n35678, n35679, n35680, n35681, n35682, n35683,
         n35684, n35685, n35686, n35687, n35688, n35689, n35690, n35691,
         n35692, n35693, n35694, n35695, n35696, n35697, n35698, n35699,
         n35700, n35701, n35702, n35703, n35704, n35705, n35706, n35707,
         n35708, n35709, n35710, n35711, n35712, n35713, n35714, n35715,
         n35716, n35717, n35718, n35719, n35720, n35721, n35722, n35723,
         n35724, n35725, n35726, n35727, n35728, n35729, n35730, n35731,
         n35732, n35733, n35734, n35735, n35736, n35737, n35738, n35739,
         n35740, n35741, n35742, n35743, n35744, n35745, n35746, n35747,
         n35748, n35749, n35750, n35751, n35752, n35753, n35754, n35755,
         n35756, n35757, n35758, n35759, n35760, n35761, n35762, n35763,
         n35764, n35765, n35766, n35767, n35768, n35769, n35770, n35771,
         n35772, n35773, n35774, n35775, n35776, n35777, n35778, n35779,
         n35780, n35781, n35782, n35783, n35784, n35785, n35786, n35787,
         n35788, n35789, n35790, n35791, n35792, n35793, n35794, n35795,
         n35796, n35797, n35798, n35799, n35800, n35801, n35802, n35803,
         n35804, n35805, n35806, n35807, n35808, n35809, n35810, n35811,
         n35812, n35813, n35814, n35815, n35816, n35817, n35818, n35819,
         n35820, n35821, n35822, n35823, n35824, n35825, n35826, n35827,
         n35828, n35829, n35830, n35831, n35832, n35833, n35834, n35835,
         n35836, n35837, n35838, n35839, n35840, n35841, n35842, n35843,
         n35844, n35845, n35846, n35847, n35848, n35849, n35850, n35851,
         n35852, n35853, n35854, n35855, n35856, n35857, n35858, n35859,
         n35860, n35861, n35862, n35863, n35864, n35865, n35866, n35867,
         n35868, n35869, n35870, n35871, n35872, n35873, n35874, n35875,
         n35876, n35877, n35878, n35879, n35880, n35881, n35882, n35883,
         n35884, n35885, n35886, n35887, n35888, n35889, n35890, n35891,
         n35892, n35893, n35894, n35895, n35896, n35897, n35898, n35899,
         n35900, n35901, n35902, n35903, n35904, n35905, n35906, n35907,
         n35908, n35909, n35910, n35911, n35912, n35913, n35914, n35915,
         n35916, n35917, n35918, n35919, n35920, n35921, n35922, n35923,
         n35924, n35925, n35926, n35927, n35928, n35929, n35930, n35931,
         n35932, n35933, n35934, n35935, n35936, n35937, n35938, n35939,
         n35940, n35941, n35942, n35943, n35944, n35945, n35946, n35947,
         n35948, n35949, n35950, n35951, n35952, n35953, n35954, n35955,
         n35956, n35957, n35958, n35959, n35960, n35961, n35962, n35963,
         n35964, n35965, n35966, n35967, n35968, n35969, n35970, n35971,
         n35972, n35973, n35974, n35975, n35976, n35977, n35978, n35979,
         n35980, n35981, n35982, n35983, n35984, n35985, n35986, n35987,
         n35988, n35989, n35990, n35991, n35992, n35993, n35994, n35995,
         n35996, n35997, n35998, n35999, n36000, n36001, n36002, n36003,
         n36004, n36005, n36006, n36007, n36008, n36009, n36010, n36011,
         n36012, n36013, n36014, n36015, n36016, n36017, n36018, n36019,
         n36020, n36021, n36022, n36023, n36024, n36025, n36026, n36027,
         n36028, n36029, n36030, n36031, n36032, n36033, n36034, n36035,
         n36036, n36037, n36038, n36039, n36040, n36041, n36042, n36043,
         n36044, n36045, n36046, n36047, n36048, n36049, n36050, n36051,
         n36052, n36053, n36054, n36055, n36056, n36057, n36058, n36059,
         n36060, n36061, n36062, n36063, n36064, n36065, n36066, n36067,
         n36068, n36069, n36070, n36071, n36072, n36073, n36074, n36075,
         n36076, n36077, n36078, n36079, n36080, n36081, n36082, n36083,
         n36084, n36085, n36086, n36087, n36088, n36089, n36090, n36091,
         n36092, n36093, n36094, n36095, n36096, n36097, n36098, n36099,
         n36100, n36101, n36102, n36103, n36104, n36105, n36106, n36107,
         n36108, n36109, n36110, n36111, n36112, n36113, n36114, n36115,
         n36116, n36117, n36118, n36119, n36120, n36121, n36122, n36123,
         n36124, n36125, n36126, n36127, n36128, n36129, n36130, n36131,
         n36132, n36133, n36134, n36135, n36136, n36137, n36138, n36139,
         n36140, n36141, n36142, n36143, n36144, n36145, n36146, n36147,
         n36148, n36149, n36150, n36151, n36152, n36153, n36154, n36155,
         n36156, n36157, n36158, n36159, n36160, n36161, n36162, n36163,
         n36164, n36165, n36166, n36167, n36168, n36169, n36170, n36171,
         n36172, n36173, n36174, n36175, n36176, n36177, n36178, n36179,
         n36180, n36181, n36182, n36183, n36184, n36185, n36186, n36187,
         n36188, n36189, n36190, n36191, n36192, n36193, n36194, n36195,
         n36196, n36197, n36198, n36199, n36200, n36201, n36202, n36203,
         n36204, n36205, n36206, n36207, n36208, n36209, n36210, n36211,
         n36212, n36213, n36214, n36215, n36216, n36217, n36218, n36219,
         n36220, n36221, n36222, n36223, n36224, n36225, n36226, n36227,
         n36228, n36229, n36230, n36231, n36232, n36233, n36234, n36235,
         n36236, n36237, n36238, n36239, n36240, n36241, n36242, n36243,
         n36244, n36245, n36246, n36247, n36248, n36249, n36250, n36251,
         n36252, n36253, n36254, n36255, n36256, n36257, n36258, n36259,
         n36260, n36261, n36262, n36263, n36264, n36265, n36266, n36267,
         n36268, n36269, n36270, n36271, n36272, n36273, n36274, n36275,
         n36276, n36277, n36278, n36279, n36280, n36281, n36282, n36283,
         n36284, n36285, n36286, n36287, n36288, n36289, n36290, n36291,
         n36292, n36293, n36294, n36295, n36296, n36297, n36298, n36299,
         n36300, n36301, n36302, n36303, n36304, n36305, n36306, n36307,
         n36308, n36309, n36310, n36311, n36312, n36313, n36314, n36315,
         n36316, n36317, n36318, n36319, n36320, n36321, n36322, n36323,
         n36324, n36325, n36326, n36327, n36328, n36329, n36330, n36331,
         n36332, n36333, n36334, n36335, n36336, n36337, n36338, n36339,
         n36340, n36341, n36342, n36343, n36344, n36345, n36346, n36347,
         n36348, n36349, n36350, n36351, n36352, n36353, n36354, n36355,
         n36356, n36357, n36358, n36359, n36360, n36361, n36362, n36363,
         n36364, n36365, n36366, n36367, n36368, n36369, n36370, n36371,
         n36372, n36373, n36374, n36375, n36376, n36377, n36378, n36379,
         n36380, n36381, n36382, n36383, n36384, n36385, n36386, n36387,
         n36388, n36389, n36390, n36391, n36392, n36393, n36394, n36395,
         n36396, n36397, n36398, n36399, n36400, n36401, n36402, n36403,
         n36404, n36405, n36406, n36407, n36408, n36409, n36410, n36411,
         n36412, n36413, n36414, n36415, n36416, n36417, n36418, n36419,
         n36420, n36421, n36422, n36423, n36424, n36425, n36426, n36427,
         n36428, n36429, n36430, n36431, n36432, n36433, n36434, n36435,
         n36436, n36437, n36438, n36439, n36440, n36441, n36442, n36443,
         n36444, n36445, n36446, n36447, n36448, n36449, n36450, n36451,
         n36452, n36453, n36454, n36455, n36456, n36457, n36458, n36459,
         n36460, n36461, n36462, n36463, n36464, n36465, n36466, n36467,
         n36468, n36469, n36470, n36471, n36472, n36473, n36474, n36475,
         n36476, n36477, n36478, n36479, n36480, n36481, n36482, n36483,
         n36484, n36485, n36486, n36487, n36488, n36489, n36490, n36491,
         n36492, n36493, n36494, n36495, n36496, n36497, n36498, n36499,
         n36500, n36501, n36502, n36503, n36504, n36505, n36506, n36507,
         n36508, n36509, n36510, n36511, n36512, n36513, n36514, n36515,
         n36516, n36517, n36518, n36519, n36520, n36521, n36522, n36523,
         n36524, n36525, n36526, n36527, n36528, n36529, n36530, n36531,
         n36532, n36533, n36534, n36535, n36536, n36537, n36538, n36539,
         n36540, n36541, n36542, n36543, n36544, n36545, n36546, n36547,
         n36548, n36549, n36550, n36551, n36552, n36553, n36554, n36555,
         n36556, n36557, n36558, n36559, n36560, n36561, n36562, n36563,
         n36564, n36565, n36566, n36567, n36568, n36569, n36570, n36571,
         n36572, n36573, n36574, n36575, n36576, n36577, n36578, n36579,
         n36580, n36581, n36582, n36583, n36584, n36585, n36586, n36587,
         n36588, n36589, n36590, n36591, n36592, n36593, n36594, n36595,
         n36596, n36597, n36598, n36599, n36600, n36601, n36602, n36603,
         n36604, n36605, n36606, n36607, n36608, n36609, n36610, n36611,
         n36612, n36613, n36614, n36615, n36616, n36617, n36618, n36619,
         n36620, n36621, n36622, n36623, n36624, n36625, n36626, n36627,
         n36628, n36629, n36630, n36631, n36632, n36633, n36634, n36635,
         n36636, n36637, n36638, n36639, n36640, n36641, n36642, n36643,
         n36644, n36645, n36646, n36647, n36648, n36649, n36650, n36651,
         n36652, n36653, n36654, n36655, n36656, n36657, n36658, n36659,
         n36660, n36661, n36662, n36663, n36664, n36665, n36666, n36667,
         n36668, n36669, n36670, n36671, n36672, n36673, n36674, n36675,
         n36676, n36677, n36678, n36679, n36680, n36681, n36682, n36683,
         n36684, n36685, n36686, n36687, n36688, n36689, n36690, n36691,
         n36692, n36693, n36694, n36695, n36696, n36697, n36698, n36699,
         n36700, n36701, n36702, n36703, n36704, n36705, n36706, n36707,
         n36708, n36709, n36710, n36711, n36712, n36713, n36714, n36715,
         n36716, n36717, n36718, n36719, n36720, n36721, n36722, n36723,
         n36724, n36725, n36726, n36727, n36728, n36729, n36730, n36731,
         n36732, n36733, n36734, n36735, n36736, n36737, n36738, n36739,
         n36740, n36741, n36742, n36743, n36744, n36745, n36746, n36747,
         n36748, n36749, n36750, n36751, n36752, n36753, n36754, n36755,
         n36756, n36757, n36758, n36759, n36760, n36761, n36762, n36763,
         n36764, n36765, n36766, n36767, n36768, n36769, n36770, n36771,
         n36772, n36773, n36774, n36775, n36776, n36777, n36778, n36779,
         n36780, n36781, n36782, n36783, n36784, n36785, n36786, n36787,
         n36788, n36789, n36790, n36791, n36792, n36793, n36794, n36795,
         n36796, n36797, n36798, n36799, n36800, n36801, n36802, n36803,
         n36804, n36805, n36806, n36807, n36808, n36809, n36810, n36811,
         n36812, n36813, n36814, n36815, n36816, n36817, n36818, n36819,
         n36820, n36821, n36822, n36823, n36824, n36825, n36826, n36827,
         n36828, n36829, n36830, n36831, n36832, n36833, n36834, n36835,
         n36836, n36837, n36838, n36839, n36840, n36841, n36842, n36843,
         n36844, n36845, n36846, n36847, n36848, n36849, n36850, n36851,
         n36852, n36853, n36854, n36855, n36856, n36857, n36858, n36859,
         n36860, n36861, n36862, n36863, n36864, n36865, n36866, n36867,
         n36868, n36869, n36870, n36871, n36872, n36873, n36874, n36875,
         n36876, n36877, n36878, n36879, n36880, n36881, n36882, n36883,
         n36884, n36885, n36886, n36887, n36888, n36889, n36890, n36891,
         n36892, n36893, n36894, n36895, n36896, n36897, n36898, n36899,
         n36900, n36901, n36902, n36903, n36904, n36905, n36906, n36907,
         n36908, n36909, n36910, n36911, n36912, n36913, n36914, n36915,
         n36916, n36917, n36918, n36919, n36920, n36921, n36922, n36923,
         n36924, n36925, n36926, n36927, n36928, n36929, n36930, n36931,
         n36932, n36933, n36934, n36935, n36936, n36937, n36938, n36939,
         n36940, n36941, n36942, n36943, n36944, n36945, n36946, n36947,
         n36948, n36949, n36950, n36951, n36952, n36953, n36954, n36955,
         n36956, n36957, n36958, n36959, n36960, n36961, n36962, n36963,
         n36964, n36965, n36966, n36967, n36968, n36969, n36970, n36971,
         n36972, n36973, n36974, n36975, n36976, n36977, n36978, n36979,
         n36980, n36981, n36982, n36983, n36984, n36985, n36986, n36987,
         n36988, n36989, n36990, n36991, n36992, n36993, n36994, n36995,
         n36996, n36997, n36998, n36999, n37000, n37001, n37002, n37003,
         n37004, n37005, n37006, n37007, n37008, n37009, n37010, n37011,
         n37012, n37013, n37014, n37015, n37016, n37017, n37018, n37019,
         n37020, n37021, n37022, n37023, n37024, n37025, n37026, n37027,
         n37028, n37029, n37030, n37031, n37032, n37033, n37034, n37035,
         n37036, n37037, n37038, n37039, n37040, n37041, n37042, n37043,
         n37044, n37045, n37046, n37047, n37048, n37049, n37050, n37051,
         n37052, n37053, n37054, n37055, n37056, n37057, n37058, n37059,
         n37060, n37061, n37062, n37063, n37064, n37065, n37066, n37067,
         n37068, n37069, n37070, n37071, n37072, n37073, n37074, n37075,
         n37076, n37077, n37078, n37079, n37080, n37081, n37082, n37083,
         n37084, n37085, n37086, n37087, n37088, n37089, n37090, n37091,
         n37092, n37093, n37094, n37095, n37096, n37097, n37098, n37099,
         n37100, n37101, n37102, n37103, n37104, n37105, n37106, n37107,
         n37108, n37109, n37110, n37111, n37112, n37113, n37114, n37115,
         n37116, n37117, n37118, n37119, n37120, n37121, n37122, n37123,
         n37124, n37125, n37126, n37127, n37128, n37129, n37130, n37131,
         n37132, n37133, n37134, n37135, n37136, n37137, n37138, n37139,
         n37140, n37141, n37142, n37143, n37144, n37145, n37146, n37147,
         n37148, n37149, n37150, n37151, n37152, n37153, n37154, n37155,
         n37156, n37157, n37158, n37159, n37160, n37161, n37162, n37163,
         n37164, n37165, n37166, n37167, n37168, n37169, n37170, n37171,
         n37172, n37173, n37174, n37175, n37176, n37177, n37178, n37179,
         n37180, n37181, n37182, n37183, n37184, n37185, n37186, n37187,
         n37188, n37189, n37190, n37191, n37192, n37193, n37194, n37195,
         n37196, n37197, n37198, n37199, n37200, n37201, n37202, n37203,
         n37204, n37205, n37206, n37207, n37208, n37209, n37210, n37211,
         n37212, n37213, n37214, n37215, n37216, n37217, n37218, n37219,
         n37220, n37221, n37222, n37223, n37224, n37225, n37226, n37227,
         n37228, n37229, n37230, n37231, n37232, n37233, n37234, n37235,
         n37236, n37237, n37238, n37239, n37240, n37241, n37242, n37243,
         n37244, n37245, n37246, n37247, n37248, n37249, n37250, n37251,
         n37252, n37253, n37254, n37255, n37256, n37257, n37258, n37259,
         n37260, n37261, n37262, n37263, n37264, n37265, n37266, n37267,
         n37268, n37269, n37270, n37271, n37272, n37273, n37274, n37275,
         n37276, n37277, n37278, n37279, n37280, n37281, n37282, n37283,
         n37284, n37285, n37286, n37287, n37288, n37289, n37290, n37291,
         n37292, n37293, n37294, n37295, n37296, n37297, n37298, n37299,
         n37300, n37301, n37302, n37303, n37304, n37305, n37306, n37307,
         n37308, n37309, n37310, n37311, n37312, n37313, n37314, n37315,
         n37316, n37317, n37318, n37319, n37320, n37321, n37322, n37323,
         n37324, n37325, n37326, n37327, n37328, n37329, n37330, n37331,
         n37332, n37333, n37334, n37335, n37336, n37337, n37338, n37339,
         n37340, n37341, n37342, n37343, n37344, n37345, n37346, n37347,
         n37348, n37349, n37350, n37351, n37352, n37353, n37354, n37355,
         n37356, n37357, n37358, n37359, n37360, n37361, n37362, n37363,
         n37364, n37365, n37366, n37367, n37368, n37369, n37370, n37371,
         n37372, n37373, n37374, n37375, n37376, n37377, n37378, n37379,
         n37380, n37381, n37382, n37383, n37384, n37385, n37386, n37387,
         n37388, n37389, n37390, n37391, n37392, n37393, n37394, n37395,
         n37396, n37397, n37398, n37399, n37400, n37401, n37402, n37403,
         n37404, n37405, n37406, n37407, n37408, n37409, n37410, n37411,
         n37412, n37413, n37414, n37415, n37416, n37417, n37418, n37419,
         n37420, n37421, n37422, n37423, n37424, n37425, n37426, n37427,
         n37428, n37429, n37430, n37431, n37432, n37433, n37434, n37435,
         n37436, n37437, n37438, n37439, n37440, n37441, n37442, n37443,
         n37444, n37445, n37446, n37447, n37448, n37449, n37450, n37451,
         n37452, n37453, n37454, n37455, n37456, n37457, n37458, n37459,
         n37460, n37461, n37462, n37463, n37464, n37465, n37466, n37467,
         n37468, n37469, n37470, n37471, n37472, n37473, n37474, n37475,
         n37476, n37477, n37478, n37479, n37480, n37481, n37482, n37483,
         n37484, n37485, n37486, n37487, n37488, n37489, n37490, n37491,
         n37492, n37493, n37494, n37495, n37496, n37497, n37498, n37499,
         n37500, n37501, n37502, n37503, n37504, n37505, n37506, n37507,
         n37508, n37509, n37510, n37511, n37512, n37513, n37514, n37515,
         n37516, n37517, n37518, n37519, n37520, n37521, n37522, n37523,
         n37524, n37525, n37526, n37527, n37528, n37529, n37530, n37531,
         n37532, n37533, n37534, n37535, n37536, n37537, n37538, n37539,
         n37540, n37541, n37542, n37543, n37544, n37545, n37546, n37547,
         n37548, n37549, n37550, n37551, n37552, n37553, n37554, n37555,
         n37556, n37557, n37558, n37559, n37560, n37561, n37562, n37563,
         n37564, n37565, n37566, n37567, n37568, n37569, n37570, n37571,
         n37572, n37573, n37574, n37575, n37576, n37577, n37578, n37579,
         n37580, n37581, n37582, n37583, n37584, n37585, n37586, n37587,
         n37588, n37589, n37590, n37591, n37592, n37593, n37594, n37595,
         n37596, n37597, n37598, n37599, n37600, n37601, n37602, n37603,
         n37604, n37605, n37606, n37607, n37608, n37609, n37610, n37611,
         n37612, n37613, n37614, n37615, n37616, n37617, n37618, n37619,
         n37620, n37621, n37622, n37623, n37624, n37625, n37626, n37627,
         n37628, n37629, n37630, n37631, n37632, n37633, n37634, n37635,
         n37636, n37637, n37638, n37639, n37640, n37641, n37642, n37643,
         n37644, n37645, n37646, n37647, n37648, n37649, n37650, n37651,
         n37652, n37653, n37654, n37655, n37656, n37657, n37658, n37659,
         n37660, n37661, n37662, n37663, n37664, n37665, n37666, n37667,
         n37668, n37669, n37670, n37671, n37672, n37673, n37674, n37675,
         n37676, n37677, n37678, n37679, n37680, n37681, n37682, n37683,
         n37684, n37685, n37686, n37687, n37688, n37689, n37690, n37691,
         n37692, n37693, n37694, n37695, n37696, n37697, n37698, n37699,
         n37700, n37701, n37702, n37703, n37704, n37705, n37706, n37707,
         n37708, n37709, n37710, n37711, n37712, n37713, n37714, n37715,
         n37716, n37717, n37718, n37719, n37720, n37721, n37722, n37723,
         n37724, n37725, n37726, n37727, n37728, n37729, n37730, n37731,
         n37732, n37733, n37734, n37735, n37736, n37737, n37738, n37739,
         n37740, n37741, n37742, n37743, n37744, n37745, n37746, n37747,
         n37748, n37749, n37750, n37751, n37752, n37753, n37754, n37755,
         n37756, n37757, n37758, n37759, n37760, n37761, n37762, n37763,
         n37764, n37765, n37766, n37767, n37768, n37769, n37770, n37771,
         n37772, n37773, n37774, n37775, n37776, n37777, n37778, n37779,
         n37780, n37781, n37782, n37783, n37784, n37785, n37786, n37787,
         n37788, n37789, n37790, n37791, n37792, n37793, n37794, n37795,
         n37796, n37797, n37798, n37799, n37800, n37801, n37802, n37803,
         n37804, n37805, n37806, n37807, n37808, n37809, n37810, n37811,
         n37812, n37813, n37814, n37815, n37816, n37817, n37818, n37819,
         n37820, n37821, n37822, n37823, n37824, n37825, n37826, n37827,
         n37828, n37829, n37830, n37831, n37832, n37833, n37834, n37835,
         n37836, n37837, n37838, n37839, n37840, n37841, n37842, n37843,
         n37844, n37845, n37846, n37847, n37848, n37849, n37850, n37851,
         n37852, n37853, n37854, n37855, n37856, n37857, n37858, n37859,
         n37860, n37861, n37862, n37863, n37864, n37865, n37866, n37867,
         n37868, n37869, n37870, n37871, n37872, n37873, n37874, n37875,
         n37876, n37877, n37878, n37879, n37880, n37881, n37882, n37883,
         n37884, n37885, n37886, n37887, n37888, n37889, n37890, n37891,
         n37892, n37893, n37894, n37895, n37896, n37897, n37898, n37899,
         n37900, n37901, n37902, n37903, n37904, n37905, n37906, n37907,
         n37908, n37909, n37910, n37911, n37912, n37913, n37914, n37915,
         n37916, n37917, n37918, n37919, n37920, n37921, n37922, n37923,
         n37924, n37925, n37926, n37927, n37928, n37929, n37930, n37931,
         n37932, n37933, n37934, n37935, n37936, n37937, n37938, n37939,
         n37940, n37941, n37942, n37943, n37944, n37945, n37946, n37947,
         n37948, n37949, n37950, n37951, n37952, n37953, n37954, n37955,
         n37956, n37957, n37958, n37959, n37960, n37961, n37962, n37963,
         n37964, n37965, n37966, n37967, n37968, n37969, n37970, n37971,
         n37972, n37973, n37974, n37975, n37976, n37977, n37978, n37979,
         n37980, n37981, n37982, n37983, n37984, n37985, n37986, n37987,
         n37988, n37989, n37990, n37991, n37992, n37993, n37994, n37995,
         n37996, n37997, n37998, n37999, n38000, n38001, n38002, n38003,
         n38004, n38005, n38006, n38007, n38008, n38009, n38010, n38011,
         n38012, n38013, n38014, n38015, n38016, n38017, n38018, n38019,
         n38020, n38021, n38022, n38023, n38024, n38025, n38026, n38027,
         n38028, n38029, n38030, n38031, n38032, n38033, n38034, n38035,
         n38036, n38037, n38038, n38039, n38040, n38041, n38042, n38043,
         n38044, n38045, n38046, n38047, n38048, n38049, n38050, n38051,
         n38052, n38053, n38054, n38055, n38056, n38057, n38058, n38059,
         n38060, n38061, n38062, n38063, n38064, n38065, n38066, n38067,
         n38068, n38069, n38070, n38071, n38072, n38073, n38074, n38075,
         n38076, n38077, n38078, n38079, n38080, n38081, n38082, n38083,
         n38084, n38085, n38086, n38087, n38088, n38089, n38090, n38091,
         n38092, n38093, n38094, n38095, n38096, n38097, n38098, n38099,
         n38100, n38101, n38102, n38103, n38104, n38105, n38106, n38107,
         n38108, n38109, n38110, n38111, n38112, n38113, n38114, n38115,
         n38116, n38117, n38118, n38119, n38120, n38121, n38122, n38123,
         n38124, n38125, n38126, n38127, n38128, n38129, n38130, n38131,
         n38132, n38133, n38134, n38135, n38136, n38137, n38138, n38139,
         n38140, n38141, n38142, n38143, n38144, n38145, n38146, n38147,
         n38148, n38149, n38150, n38151, n38152, n38153, n38154, n38155,
         n38156, n38157, n38158, n38159, n38160, n38161, n38162, n38163,
         n38164, n38165, n38166, n38167, n38168, n38169, n38170, n38171,
         n38172, n38173, n38174, n38175, n38176, n38177, n38178, n38179,
         n38180, n38181, n38182, n38183, n38184, n38185, n38186, n38187,
         n38188, n38189, n38190, n38191, n38192, n38193, n38194, n38195,
         n38196, n38197, n38198, n38199, n38200, n38201, n38202, n38203,
         n38204, n38205, n38206, n38207, n38208, n38209, n38210, n38211,
         n38212, n38213, n38214, n38215, n38216, n38217, n38218, n38219,
         n38220, n38221, n38222, n38223, n38224, n38225, n38226, n38227,
         n38228, n38229, n38230, n38231, n38232, n38233, n38234, n38235,
         n38236, n38237, n38238, n38239, n38240, n38241, n38242, n38243,
         n38244, n38245, n38246, n38247, n38248, n38249, n38250, n38251,
         n38252, n38253, n38254, n38255, n38256, n38257, n38258, n38259,
         n38260, n38261, n38262, n38263, n38264, n38265, n38266, n38267,
         n38268, n38269, n38270, n38271, n38272, n38273, n38274, n38275,
         n38276, n38277, n38278, n38279, n38280, n38281, n38282, n38283,
         n38284, n38285, n38286, n38287, n38288, n38289, n38290, n38291,
         n38292, n38293, n38294, n38295, n38296, n38297, n38298, n38299,
         n38300, n38301, n38302, n38303, n38304, n38305, n38306, n38307,
         n38308, n38309, n38310, n38311, n38312, n38313, n38314, n38315,
         n38316, n38317, n38318, n38319, n38320, n38321, n38322, n38323,
         n38324, n38325, n38326, n38327, n38328, n38329, n38330, n38331,
         n38332, n38333, n38334, n38335, n38336, n38337, n38338, n38339,
         n38340, n38341, n38342, n38343, n38344, n38345, n38346, n38347,
         n38348, n38349, n38350, n38351, n38352, n38353, n38354, n38355,
         n38356, n38357, n38358, n38359, n38360, n38361, n38362, n38363,
         n38364, n38365, n38366, n38367, n38368, n38369, n38370, n38371,
         n38372, n38373, n38374, n38375, n38376, n38377, n38378, n38379,
         n38380, n38381, n38382, n38383, n38384, n38385, n38386, n38387,
         n38388, n38389, n38390, n38391, n38392, n38393, n38394, n38395,
         n38396, n38397, n38398, n38399, n38400, n38401, n38402, n38403,
         n38404, n38405, n38406, n38407, n38408, n38409, n38410, n38411,
         n38412, n38413, n38414, n38415, n38416, n38417, n38418, n38419,
         n38420, n38421, n38422, n38423, n38424, n38425, n38426, n38427,
         n38428, n38429, n38430, n38431, n38432, n38433, n38434, n38435,
         n38436, n38437, n38438, n38439, n38440, n38441, n38442, n38443,
         n38444, n38445, n38446, n38447, n38448, n38449, n38450, n38451,
         n38452, n38453, n38454, n38455, n38456, n38457, n38458, n38459,
         n38460, n38461, n38462, n38463, n38464, n38465, n38466, n38467,
         n38468, n38469, n38470, n38471, n38472, n38473, n38474, n38475,
         n38476, n38477, n38478, n38479, n38480, n38481, n38482, n38483,
         n38484, n38485, n38486, n38487, n38488, n38489, n38490, n38491,
         n38492, n38493, n38494, n38495, n38496, n38497, n38498, n38499,
         n38500, n38501, n38502, n38503, n38504, n38505, n38506, n38507,
         n38508, n38509, n38510, n38511, n38512, n38513, n38514, n38515,
         n38516, n38517, n38518, n38519, n38520, n38521, n38522, n38523,
         n38524, n38525, n38526, n38527, n38528, n38529, n38530, n38531,
         n38532, n38533, n38534, n38535, n38536, n38537, n38538, n38539,
         n38540, n38541, n38542, n38543, n38544, n38545, n38546, n38547,
         n38548, n38549, n38550, n38551, n38552, n38553, n38554, n38555,
         n38556, n38557, n38558, n38559, n38560, n38561, n38562, n38563,
         n38564, n38565, n38566, n38567, n38568, n38569, n38570, n38571,
         n38572, n38573, n38574, n38575, n38576, n38577, n38578, n38579,
         n38580, n38581, n38582, n38583, n38584, n38585, n38586, n38587,
         n38588, n38589, n38590, n38591, n38592, n38593, n38594, n38595,
         n38596, n38597, n38598, n38599, n38600, n38601, n38602, n38603,
         n38604, n38605, n38606, n38607, n38608, n38609, n38610, n38611,
         n38612, n38613, n38614, n38615, n38616, n38617, n38618, n38619,
         n38620, n38621, n38622, n38623, n38624, n38625, n38626, n38627,
         n38628, n38629, n38630, n38631, n38632, n38633, n38634, n38635,
         n38636, n38637, n38638, n38639, n38640, n38641, n38642, n38643,
         n38644, n38645, n38646, n38647, n38648, n38649, n38650, n38651,
         n38652, n38653, n38654, n38655, n38656, n38657, n38658, n38659,
         n38660, n38661, n38662, n38663, n38664, n38665, n38666, n38667,
         n38668, n38669, n38670, n38671, n38672, n38673, n38674, n38675,
         n38676, n38677, n38678, n38679, n38680, n38681, n38682, n38683,
         n38684, n38685, n38686, n38687, n38688, n38689, n38690, n38691,
         n38692, n38693, n38694, n38695, n38696, n38697, n38698, n38699,
         n38700, n38701, n38702, n38703, n38704, n38705, n38706, n38707,
         n38708, n38709, n38710, n38711, n38712, n38713, n38714, n38715,
         n38716, n38717, n38718, n38719, n38720, n38721, n38722, n38723,
         n38724, n38725, n38726, n38727, n38728, n38729, n38730, n38731,
         n38732, n38733, n38734, n38735, n38736, n38737, n38738, n38739,
         n38740, n38741, n38742, n38743, n38744, n38745, n38746, n38747,
         n38748, n38749, n38750, n38751, n38752, n38753, n38754, n38755,
         n38756, n38757, n38758, n38759, n38760, n38761, n38762, n38763,
         n38764, n38765, n38766, n38767, n38768, n38769, n38770, n38771,
         n38772, n38773, n38774, n38775, n38776, n38777, n38778, n38779,
         n38780, n38781, n38782, n38783, n38784, n38785, n38786, n38787,
         n38788, n38789, n38790, n38791, n38792, n38793, n38794, n38795,
         n38796, n38797, n38798, n38799, n38800, n38801, n38802, n38803,
         n38804, n38805, n38806, n38807, n38808, n38809, n38810, n38811,
         n38812, n38813, n38814, n38815, n38816, n38817, n38818, n38819,
         n38820, n38821, n38822, n38823, n38824, n38825, n38826, n38827,
         n38828, n38829, n38830, n38831, n38832, n38833, n38834, n38835,
         n38836, n38837, n38838, n38839, n38840, n38841, n38842, n38843,
         n38844, n38845, n38846, n38847, n38848, n38849, n38850, n38851,
         n38852, n38853, n38854, n38855, n38856, n38857, n38858, n38859,
         n38860, n38861, n38862, n38863, n38864, n38865, n38866, n38867,
         n38868, n38869, n38870, n38871, n38872, n38873, n38874, n38875,
         n38876, n38877, n38878, n38879, n38880, n38881, n38882, n38883,
         n38884, n38885, n38886, n38887, n38888, n38889, n38890, n38891,
         n38892, n38893, n38894, n38895, n38896, n38897, n38898, n38899,
         n38900, n38901, n38902, n38903, n38904, n38905, n38906, n38907,
         n38908, n38909, n38910, n38911, n38912, n38913, n38914, n38915,
         n38916, n38917, n38918, n38919, n38920, n38921, n38922, n38923,
         n38924, n38925, n38926, n38927, n38928, n38929, n38930, n38931,
         n38932, n38933, n38934, n38935, n38936, n38937, n38938, n38939,
         n38940, n38941, n38942, n38943, n38944, n38945, n38946, n38947,
         n38948, n38949, n38950, n38951, n38952, n38953, n38954, n38955,
         n38956, n38957, n38958, n38959, n38960, n38961, n38962, n38963,
         n38964, n38965, n38966, n38967, n38968, n38969, n38970, n38971,
         n38972, n38973, n38974, n38975, n38976, n38977, n38978, n38979,
         n38980, n38981, n38982, n38983, n38984, n38985, n38986, n38987,
         n38988, n38989, n38990, n38991, n38992, n38993, n38994, n38995,
         n38996, n38997, n38998, n38999, n39000, n39001, n39002, n39003,
         n39004, n39005, n39006, n39007, n39008, n39009, n39010, n39011,
         n39012, n39013, n39014, n39015, n39016, n39017, n39018, n39019,
         n39020, n39021, n39022, n39023, n39024, n39025, n39026, n39027,
         n39028, n39029, n39030, n39031, n39032, n39033, n39034, n39035,
         n39036, n39037, n39038, n39039, n39040, n39041, n39042, n39043,
         n39044, n39045, n39046, n39047, n39048, n39049, n39050, n39051,
         n39052, n39053, n39054, n39055, n39056, n39057, n39058, n39059,
         n39060, n39061, n39062, n39063, n39064, n39065, n39066, n39067,
         n39068, n39069, n39070, n39071, n39072, n39073, n39074, n39075,
         n39076, n39077, n39078, n39079, n39080, n39081, n39082, n39083,
         n39084, n39085, n39086, n39087, n39088, n39089, n39090, n39091,
         n39092, n39093, n39094, n39095, n39096, n39097, n39098, n39099,
         n39100, n39101, n39102, n39103, n39104, n39105, n39106, n39107,
         n39108, n39109, n39110, n39111, n39112, n39113, n39114, n39115,
         n39116, n39117, n39118, n39119, n39120, n39121, n39122, n39123,
         n39124, n39125, n39126, n39127, n39128, n39129, n39130, n39131,
         n39132, n39133, n39134, n39135, n39136, n39137, n39138, n39139,
         n39140, n39141, n39142, n39143, n39144, n39145, n39146, n39147,
         n39148, n39149, n39150, n39151, n39152, n39153, n39154, n39155,
         n39156, n39157, n39158, n39159, n39160, n39161, n39162, n39163,
         n39164, n39165, n39166, n39167, n39168, n39169, n39170, n39171,
         n39172, n39173, n39174, n39175, n39176, n39177, n39178, n39179,
         n39180, n39181, n39182, n39183, n39184, n39185, n39186, n39187,
         n39188, n39189, n39190, n39191, n39192, n39193, n39194, n39195,
         n39196, n39197, n39198, n39199, n39200, n39201, n39202, n39203,
         n39204, n39205, n39206, n39207, n39208, n39209, n39210, n39211,
         n39212, n39213, n39214, n39215, n39216, n39217, n39218, n39219,
         n39220, n39221, n39222, n39223, n39224, n39225, n39226, n39227,
         n39228, n39229, n39230, n39231, n39232, n39233, n39234, n39235,
         n39236, n39237, n39238, n39239, n39240, n39241, n39242, n39243,
         n39244, n39245, n39246, n39247, n39248, n39249, n39250, n39251,
         n39252, n39253, n39254, n39255, n39256, n39257, n39258, n39259,
         n39260, n39261, n39262, n39263, n39264, n39265, n39266, n39267,
         n39268, n39269, n39270, n39271, n39272, n39273, n39274, n39275,
         n39276, n39277, n39278, n39279, n39280, n39281, n39282, n39283,
         n39284, n39285, n39286, n39287, n39288, n39289, n39290, n39291,
         n39292, n39293, n39294, n39295, n39296, n39297, n39298, n39299,
         n39300, n39301, n39302, n39303, n39304, n39305, n39306, n39307,
         n39308, n39309, n39310, n39311, n39312, n39313, n39314, n39315,
         n39316, n39317, n39318, n39319, n39320, n39321, n39322, n39323,
         n39324, n39325, n39326, n39327, n39328, n39329, n39330, n39331,
         n39332, n39333, n39334, n39335, n39336, n39337, n39338, n39339,
         n39340, n39341, n39342, n39343, n39344, n39345, n39346, n39347,
         n39348, n39349, n39350, n39351, n39352, n39353, n39354, n39355,
         n39356, n39357, n39358, n39359, n39360, n39361, n39362, n39363,
         n39364, n39365, n39366, n39367, n39368, n39369, n39370, n39371,
         n39372, n39373, n39374, n39375, n39376, n39377, n39378, n39379,
         n39380, n39381, n39382, n39383, n39384, n39385, n39386, n39387,
         n39388, n39389, n39390, n39391, n39392, n39393, n39394, n39395,
         n39396, n39397, n39398, n39399, n39400, n39401, n39402, n39403,
         n39404, n39405, n39406, n39407, n39408, n39409, n39410, n39411,
         n39412, n39413, n39414, n39415, n39416, n39417, n39418, n39419,
         n39420, n39421, n39422, n39423, n39424, n39425, n39426, n39427,
         n39428, n39429, n39430, n39431, n39432, n39433, n39434, n39435,
         n39436, n39437, n39438, n39439, n39440, n39441, n39442, n39443,
         n39444, n39445, n39446, n39447, n39448, n39449, n39450, n39451,
         n39452, n39453, n39454, n39455, n39456, n39457, n39458, n39459,
         n39460, n39461, n39462, n39463, n39464, n39465, n39466, n39467,
         n39468, n39469, n39470, n39471, n39472, n39473, n39474, n39475,
         n39476, n39477, n39478, n39479, n39480, n39481, n39482, n39483,
         n39484, n39485, n39486, n39487, n39488, n39489, n39490, n39491,
         n39492, n39493, n39494, n39495, n39496, n39497, n39498, n39499,
         n39500, n39501, n39502, n39503, n39504, n39505, n39506, n39507,
         n39508, n39509, n39510, n39511, n39512, n39513, n39514, n39515,
         n39516, n39517, n39518, n39519, n39520, n39521, n39522, n39523,
         n39524, n39525, n39526, n39527, n39528, n39529, n39530, n39531,
         n39532, n39533, n39534, n39535, n39536, n39537, n39538, n39539,
         n39540, n39541, n39542, n39543, n39544, n39545, n39546, n39547,
         n39548, n39549, n39550, n39551, n39552, n39553, n39554, n39555,
         n39556, n39557, n39558, n39559, n39560, n39561, n39562, n39563,
         n39564, n39565, n39566, n39567, n39568, n39569, n39570, n39571,
         n39572, n39573, n39574, n39575, n39576, n39577, n39578, n39579,
         n39580, n39581, n39582, n39583, n39584, n39585, n39586, n39587,
         n39588, n39589, n39590, n39591, n39592, n39593, n39594, n39595,
         n39596, n39597, n39598, n39599, n39600, n39601, n39602, n39603,
         n39604, n39605, n39606, n39607, n39608, n39609, n39610, n39611,
         n39612, n39613, n39614, n39615, n39616, n39617, n39618, n39619,
         n39620, n39621, n39622, n39623, n39624, n39625, n39626, n39627,
         n39628, n39629, n39630, n39631, n39632, n39633, n39634, n39635,
         n39636, n39637, n39638, n39639, n39640, n39641, n39642, n39643,
         n39644, n39645, n39646, n39647, n39648, n39649, n39650, n39651,
         n39652, n39653, n39654, n39655, n39656, n39657, n39658, n39659,
         n39660, n39661, n39662, n39663, n39664, n39665, n39666, n39667,
         n39668, n39669, n39670, n39671, n39672, n39673, n39674, n39675,
         n39676, n39677, n39678, n39679, n39680, n39681, n39682, n39683,
         n39684, n39685, n39686, n39687, n39688, n39689, n39690, n39691,
         n39692, n39693, n39694, n39695, n39696, n39697, n39698, n39699,
         n39700, n39701, n39702, n39703, n39704, n39705, n39706, n39707,
         n39708, n39709, n39710, n39711, n39712, n39713, n39714, n39715,
         n39716, n39717, n39718, n39719, n39720, n39721, n39722, n39723,
         n39724, n39725, n39726, n39727, n39728, n39729, n39730, n39731,
         n39732, n39733, n39734, n39735, n39736, n39737, n39738, n39739,
         n39740, n39741, n39742, n39743, n39744, n39745, n39746, n39747,
         n39748, n39749, n39750, n39751, n39752, n39753, n39754, n39755,
         n39756, n39757, n39758, n39759, n39760, n39761, n39762, n39763,
         n39764, n39765, n39766, n39767, n39768, n39769, n39770, n39771,
         n39772, n39773, n39774, n39775, n39776, n39777, n39778, n39779,
         n39780, n39781, n39782, n39783, n39784, n39785, n39786, n39787,
         n39788, n39789, n39790, n39791, n39792, n39793, n39794, n39795,
         n39796, n39797, n39798, n39799, n39800, n39801, n39802, n39803,
         n39804, n39805, n39806, n39807, n39808, n39809, n39810, n39811,
         n39812, n39813, n39814, n39815, n39816, n39817, n39818, n39819,
         n39820, n39821, n39822, n39823, n39824, n39825, n39826, n39827,
         n39828, n39829, n39830, n39831, n39832, n39833, n39834, n39835,
         n39836, n39837, n39838, n39839, n39840, n39841, n39842, n39843,
         n39844, n39845, n39846, n39847, n39848, n39849, n39850, n39851,
         n39852, n39853, n39854, n39855, n39856, n39857, n39858, n39859,
         n39860, n39861, n39862, n39863, n39864, n39865, n39866, n39867,
         n39868, n39869, n39870, n39871, n39872, n39873, n39874, n39875,
         n39876, n39877, n39878, n39879, n39880, n39881, n39882, n39883,
         n39884, n39885, n39886, n39887, n39888, n39889, n39890, n39891,
         n39892, n39893, n39894, n39895, n39896, n39897, n39898, n39899,
         n39900, n39901, n39902, n39903, n39904, n39905, n39906, n39907,
         n39908, n39909, n39910, n39911, n39912, n39913, n39914, n39915,
         n39916, n39917, n39918, n39919, n39920, n39921, n39922, n39923,
         n39924, n39925, n39926, n39927, n39928, n39929, n39930, n39931,
         n39932, n39933, n39934, n39935, n39936, n39937, n39938, n39939,
         n39940, n39941, n39942, n39943, n39944, n39945, n39946, n39947,
         n39948, n39949, n39950, n39951, n39952, n39953, n39954, n39955,
         n39956, n39957, n39958, n39959, n39960, n39961, n39962, n39963,
         n39964, n39965, n39966, n39967, n39968, n39969, n39970, n39971,
         n39972, n39973, n39974, n39975, n39976, n39977, n39978, n39979,
         n39980, n39981, n39982, n39983, n39984, n39985, n39986, n39987,
         n39988, n39989, n39990, n39991, n39992, n39993, n39994, n39995,
         n39996, n39997, n39998, n39999, n40000, n40001, n40002, n40003,
         n40004, n40005, n40006, n40007, n40008, n40009, n40010, n40011,
         n40012, n40013, n40014, n40015, n40016, n40017, n40018, n40019,
         n40020, n40021, n40022, n40023, n40024, n40025, n40026, n40027,
         n40028, n40029, n40030, n40031, n40032, n40033, n40034, n40035,
         n40036, n40037, n40038, n40039, n40040, n40041, n40042, n40043,
         n40044, n40045, n40046, n40047, n40048, n40049, n40050, n40051,
         n40052, n40053, n40054, n40055, n40056, n40057, n40058, n40059,
         n40060, n40061, n40062, n40063, n40064, n40065, n40066, n40067,
         n40068, n40069, n40070, n40071, n40072, n40073, n40074, n40075,
         n40076, n40077, n40078, n40079, n40080, n40081, n40082, n40083,
         n40084, n40085, n40086, n40087, n40088, n40089, n40090, n40091,
         n40092, n40093, n40094, n40095, n40096, n40097, n40098, n40099,
         n40100, n40101, n40102, n40103, n40104, n40105, n40106, n40107,
         n40108, n40109, n40110, n40111, n40112, n40113, n40114, n40115,
         n40116, n40117, n40118, n40119, n40120, n40121, n40122, n40123,
         n40124, n40125, n40126, n40127, n40128, n40129, n40130, n40131,
         n40132, n40133, n40134, n40135, n40136, n40137, n40138, n40139,
         n40140, n40141, n40142, n40143, n40144, n40145, n40146, n40147,
         n40148, n40149, n40150, n40151, n40152, n40153, n40154, n40155,
         n40156, n40157, n40158, n40159, n40160, n40161, n40162, n40163,
         n40164, n40165, n40166, n40167, n40168, n40169, n40170, n40171,
         n40172, n40173, n40174, n40175, n40176, n40177, n40178, n40179,
         n40180, n40181, n40182, n40183, n40184, n40185, n40186, n40187,
         n40188, n40189, n40190, n40191, n40192, n40193, n40194, n40195,
         n40196, n40197, n40198, n40199, n40200, n40201, n40202, n40203,
         n40204, n40205, n40206, n40207, n40208, n40209, n40210, n40211,
         n40212, n40213, n40214, n40215, n40216, n40217, n40218, n40219,
         n40220, n40221, n40222, n40223, n40224, n40225, n40226, n40227,
         n40228, n40229, n40230, n40231, n40232, n40233, n40234, n40235,
         n40236, n40237, n40238, n40239, n40240, n40241, n40242, n40243,
         n40244, n40245, n40246, n40247, n40248, n40249, n40250, n40251,
         n40252, n40253, n40254, n40255, n40256, n40257, n40258, n40259,
         n40260, n40261, n40262, n40263, n40264, n40265, n40266, n40267,
         n40268, n40269, n40270, n40271, n40272, n40273, n40274, n40275,
         n40276, n40277, n40278, n40279, n40280, n40281, n40282, n40283,
         n40284, n40285, n40286, n40287, n40288, n40289, n40290, n40291,
         n40292, n40293, n40294, n40295, n40296, n40297, n40298, n40299,
         n40300, n40301, n40302, n40303, n40304, n40305, n40306, n40307,
         n40308, n40309, n40310, n40311, n40312, n40313, n40314, n40315,
         n40316, n40317, n40318, n40319, n40320, n40321, n40322, n40323,
         n40324, n40325, n40326, n40327, n40328, n40329, n40330, n40331,
         n40332, n40333, n40334, n40335, n40336, n40337, n40338, n40339,
         n40340, n40341, n40342, n40343, n40344, n40345, n40346, n40347,
         n40348, n40349, n40350, n40351, n40352, n40353, n40354, n40355,
         n40356, n40357, n40358, n40359, n40360, n40361, n40362, n40363,
         n40364, n40365, n40366, n40367, n40368, n40369, n40370, n40371,
         n40372, n40373, n40374, n40375, n40376, n40377, n40378, n40379,
         n40380, n40381, n40382, n40383, n40384, n40385, n40386, n40387,
         n40388, n40389, n40390, n40391, n40392, n40393, n40394, n40395,
         n40396, n40397, n40398, n40399, n40400, n40401, n40402, n40403,
         n40404, n40405, n40406, n40407, n40408, n40409, n40410, n40411,
         n40412, n40413, n40414, n40415, n40416, n40417, n40418, n40419,
         n40420, n40421, n40422, n40423, n40424, n40425, n40426, n40427,
         n40428, n40429, n40430, n40431, n40432, n40433, n40434, n40435,
         n40436, n40437, n40438, n40439, n40440, n40441, n40442, n40443,
         n40444, n40445, n40446, n40447, n40448, n40449, n40450, n40451,
         n40452, n40453, n40454, n40455, n40456, n40457, n40458, n40459,
         n40460, n40461, n40462, n40463, n40464, n40465, n40466, n40467,
         n40468, n40469, n40470, n40471, n40472, n40473, n40474, n40475,
         n40476, n40477, n40478, n40479, n40480, n40481, n40482, n40483,
         n40484, n40485, n40486, n40487, n40488, n40489, n40490, n40491,
         n40492, n40493, n40494, n40495, n40496, n40497, n40498, n40499,
         n40500, n40501, n40502, n40503, n40504, n40505, n40506, n40507,
         n40508, n40509, n40510, n40511, n40512, n40513, n40514, n40515,
         n40516, n40517, n40518, n40519, n40520, n40521, n40522, n40523,
         n40524, n40525, n40526, n40527, n40528, n40529, n40530, n40531,
         n40532, n40533, n40534, n40535, n40536, n40537, n40538, n40539,
         n40540, n40541, n40542, n40543, n40544, n40545, n40546, n40547,
         n40548, n40549, n40550, n40551, n40552, n40553, n40554, n40555,
         n40556, n40557, n40558, n40559, n40560, n40561, n40562, n40563,
         n40564, n40565, n40566, n40567, n40568, n40569, n40570, n40571,
         n40572, n40573, n40574, n40575, n40576, n40577, n40578, n40579,
         n40580, n40581, n40582, n40583, n40584, n40585, n40586, n40587,
         n40588, n40589, n40590, n40591, n40592, n40593, n40594, n40595,
         n40596, n40597, n40598, n40599, n40600, n40601, n40602, n40603,
         n40604, n40605, n40606, n40607, n40608, n40609, n40610, n40611,
         n40612, n40613, n40614, n40615, n40616, n40617, n40618, n40619,
         n40620, n40621, n40622, n40623, n40624, n40625, n40626, n40627,
         n40628, n40629, n40630, n40631, n40632, n40633, n40634, n40635,
         n40636, n40637, n40638, n40639, n40640, n40641, n40642, n40643,
         n40644, n40645, n40646, n40647, n40648, n40649, n40650, n40651,
         n40652, n40653, n40654, n40655, n40656, n40657, n40658, n40659,
         n40660, n40661, n40662, n40663, n40664, n40665, n40666, n40667,
         n40668, n40669, n40670, n40671, n40672, n40673, n40674, n40675,
         n40676, n40677, n40678, n40679, n40680, n40681, n40682, n40683,
         n40684, n40685, n40686, n40687, n40688, n40689, n40690, n40691,
         n40692, n40693, n40694, n40695, n40696, n40697, n40698, n40699,
         n40700, n40701, n40702, n40703, n40704, n40705, n40706, n40707,
         n40708, n40709, n40710, n40711, n40712, n40713, n40714, n40715,
         n40716, n40717, n40718, n40719, n40720, n40721, n40722, n40723,
         n40724, n40725, n40726, n40727, n40728, n40729, n40730, n40731,
         n40732, n40733, n40734, n40735, n40736, n40737, n40738, n40739,
         n40740, n40741, n40742, n40743, n40744, n40745, n40746, n40747,
         n40748, n40749, n40750, n40751, n40752, n40753, n40754, n40755,
         n40756, n40757, n40758, n40759, n40760, n40761, n40762, n40763,
         n40764, n40765, n40766, n40767, n40768, n40769, n40770, n40771,
         n40772, n40773, n40774, n40775, n40776, n40777, n40778, n40779,
         n40780, n40781, n40782, n40783, n40784, n40785, n40786, n40787,
         n40788, n40789, n40790, n40791, n40792, n40793, n40794, n40795,
         n40796, n40797, n40798, n40799, n40800, n40801, n40802, n40803,
         n40804, n40805, n40806, n40807, n40808, n40809, n40810, n40811,
         n40812, n40813, n40814, n40815, n40816, n40817, n40818, n40819,
         n40820, n40821, n40822, n40823, n40824, n40825, n40826, n40827,
         n40828, n40829, n40830, n40831, n40832, n40833, n40834, n40835,
         n40836, n40837, n40838, n40839, n40840, n40841, n40842, n40843,
         n40844, n40845, n40846, n40847, n40848, n40849, n40850, n40851,
         n40852, n40853, n40854, n40855, n40856, n40857, n40858, n40859,
         n40860, n40861, n40862, n40863, n40864, n40865, n40866, n40867,
         n40868, n40869, n40870, n40871, n40872, n40873, n40874, n40875,
         n40876, n40877, n40878, n40879, n40880, n40881, n40882, n40883,
         n40884, n40885, n40886, n40887, n40888, n40889, n40890, n40891,
         n40892, n40893, n40894, n40895, n40896, n40897, n40898, n40899,
         n40900, n40901, n40902, n40903, n40904, n40905, n40906, n40907,
         n40908, n40909, n40910, n40911, n40912, n40913, n40914, n40915,
         n40916, n40917, n40918, n40919, n40920, n40921, n40922, n40923,
         n40924, n40925, n40926, n40927, n40928, n40929, n40930, n40931,
         n40932, n40933, n40934, n40935, n40936, n40937, n40938, n40939,
         n40940, n40941, n40942, n40943, n40944, n40945, n40946, n40947,
         n40948, n40949, n40950, n40951, n40952, n40953, n40954, n40955,
         n40956, n40957, n40958, n40959, n40960, n40961, n40962, n40963,
         n40964, n40965, n40966, n40967, n40968, n40969, n40970, n40971,
         n40972, n40973, n40974, n40975, n40976, n40977, n40978, n40979,
         n40980, n40981, n40982, n40983, n40984, n40985, n40986, n40987,
         n40988, n40989, n40990, n40991, n40992, n40993, n40994, n40995,
         n40996, n40997, n40998, n40999, n41000, n41001, n41002, n41003,
         n41004, n41005, n41006, n41007, n41008, n41009, n41010, n41011,
         n41012, n41013, n41014, n41015, n41016, n41017, n41018, n41019,
         n41020, n41021, n41022, n41023, n41024, n41025, n41026, n41027,
         n41028, n41029, n41030, n41031, n41032, n41033, n41034, n41035,
         n41036, n41037, n41038, n41039, n41040, n41041, n41042, n41043,
         n41044, n41045, n41046, n41047, n41048, n41049, n41050, n41051,
         n41052, n41053, n41054, n41055, n41056, n41057, n41058, n41059,
         n41060, n41061, n41062, n41063, n41064, n41065, n41066, n41067,
         n41068, n41069, n41070, n41071, n41072, n41073, n41074, n41075,
         n41076, n41077, n41078, n41079, n41080, n41081, n41082, n41083,
         n41084, n41085, n41086, n41087, n41088, n41089, n41090, n41091,
         n41092, n41093, n41094, n41095, n41096, n41097, n41098, n41099,
         n41100, n41101, n41102, n41103, n41104, n41105, n41106, n41107,
         n41108, n41109, n41110, n41111, n41112, n41113, n41114, n41115,
         n41116, n41117, n41118, n41119, n41120, n41121, n41122, n41123,
         n41124, n41125, n41126, n41127, n41128, n41129, n41130, n41131,
         n41132, n41133, n41134, n41135, n41136, n41137, n41138, n41139,
         n41140, n41141, n41142, n41143, n41144, n41145, n41146, n41147,
         n41148, n41149, n41150, n41151, n41152, n41153, n41154, n41155,
         n41156, n41157, n41158, n41159, n41160, n41161, n41162, n41163,
         n41164, n41165, n41166, n41167, n41168, n41169, n41170, n41171,
         n41172, n41173, n41174, n41175, n41176, n41177, n41178, n41179,
         n41180, n41181, n41182, n41183, n41184, n41185, n41186, n41187,
         n41188, n41189, n41190, n41191, n41192, n41193, n41194, n41195,
         n41196, n41197, n41198, n41199, n41200, n41201, n41202, n41203,
         n41204, n41205, n41206, n41207, n41208, n41209, n41210, n41211,
         n41212, n41213, n41214, n41215, n41216, n41217, n41218, n41219,
         n41220, n41221, n41222, n41223, n41224, n41225, n41226, n41227,
         n41228, n41229, n41230, n41231, n41232, n41233, n41234, n41235,
         n41236, n41237, n41238, n41239, n41240, n41241, n41242, n41243,
         n41244, n41245, n41246, n41247, n41248, n41249, n41250, n41251,
         n41252, n41253, n41254, n41255, n41256, n41257, n41258, n41259,
         n41260, n41261, n41262, n41263, n41264, n41265, n41266, n41267,
         n41268, n41269, n41270, n41271, n41272, n41273, n41274, n41275,
         n41276, n41277, n41278, n41279, n41280, n41281, n41282, n41283,
         n41284, n41285, n41286, n41287, n41288, n41289, n41290, n41291,
         n41292, n41293, n41294, n41295, n41296, n41297, n41298, n41299,
         n41300, n41301, n41302, n41303, n41304, n41305, n41306, n41307,
         n41308, n41309, n41310, n41311, n41312, n41313, n41314, n41315,
         n41316, n41317, n41318, n41319, n41320, n41321, n41322, n41323,
         n41324, n41325, n41326, n41327, n41328, n41329, n41330, n41331,
         n41332, n41333, n41334, n41335, n41336, n41337, n41338, n41339,
         n41340, n41341, n41342, n41343, n41344, n41345, n41346, n41347,
         n41348, n41349, n41350, n41351, n41352, n41353, n41354, n41355,
         n41356, n41357, n41358, n41359, n41360, n41361, n41362, n41363,
         n41364, n41365, n41366, n41367, n41368, n41369, n41370, n41371,
         n41372, n41373, n41374, n41375, n41376, n41377, n41378, n41379,
         n41380, n41381, n41382, n41383, n41384, n41385, n41386, n41387,
         n41388, n41389, n41390, n41391, n41392, n41393, n41394, n41395,
         n41396, n41397, n41398, n41399, n41400, n41401, n41402, n41403,
         n41404, n41405, n41406, n41407, n41408, n41409, n41410, n41411,
         n41412, n41413, n41414, n41415, n41416, n41417, n41418, n41419,
         n41420, n41421, n41422, n41423, n41424, n41425, n41426, n41427,
         n41428, n41429, n41430, n41431, n41432, n41433, n41434, n41435,
         n41436, n41437, n41438, n41439, n41440, n41441, n41442, n41443,
         n41444, n41445, n41446, n41447, n41448, n41449, n41450, n41451,
         n41452, n41453, n41454, n41455, n41456, n41457, n41458, n41459,
         n41460, n41461, n41462, n41463, n41464, n41465, n41466, n41467,
         n41468, n41469, n41470, n41471, n41472, n41473, n41474, n41475,
         n41476, n41477, n41478, n41479, n41480, n41481, n41482, n41483,
         n41484, n41485, n41486, n41487, n41488, n41489, n41490, n41491,
         n41492, n41493, n41494, n41495, n41496, n41497, n41498, n41499,
         n41500, n41501, n41502, n41503, n41504, n41505, n41506, n41507,
         n41508, n41509, n41510, n41511, n41512, n41513, n41514, n41515,
         n41516, n41517, n41518, n41519, n41520, n41521, n41522, n41523,
         n41524, n41525, n41526, n41527, n41528, n41529, n41530, n41531,
         n41532, n41533, n41534, n41535, n41536, n41537, n41538, n41539,
         n41540, n41541, n41542, n41543, n41544, n41545, n41546, n41547,
         n41548, n41549, n41550, n41551, n41552, n41553, n41554, n41555,
         n41556, n41557, n41558, n41559, n41560, n41561, n41562, n41563,
         n41564, n41565, n41566, n41567, n41568, n41569, n41570, n41571,
         n41572, n41573, n41574, n41575, n41576, n41577, n41578, n41579,
         n41580, n41581, n41582, n41583, n41584, n41585, n41586, n41587,
         n41588, n41589, n41590, n41591, n41592, n41593, n41594, n41595,
         n41596, n41597, n41598, n41599, n41600, n41601, n41602, n41603,
         n41604, n41605, n41606, n41607, n41608, n41609, n41610, n41611,
         n41612, n41613, n41614, n41615, n41616, n41617, n41618, n41619,
         n41620, n41621, n41622, n41623, n41624, n41625, n41626, n41627,
         n41628, n41629, n41630, n41631, n41632, n41633, n41634, n41635,
         n41636, n41637, n41638, n41639, n41640, n41641, n41642, n41643,
         n41644, n41645, n41646, n41647, n41648, n41649, n41650, n41651,
         n41652, n41653, n41654, n41655, n41656, n41657, n41658, n41659,
         n41660, n41661, n41662, n41663, n41664, n41665, n41666, n41667,
         n41668, n41669, n41670, n41671, n41672, n41673, n41674, n41675,
         n41676, n41677, n41678, n41679, n41680, n41681, n41682, n41683,
         n41684, n41685, n41686, n41687, n41688, n41689, n41690, n41691,
         n41692, n41693, n41694, n41695, n41696, n41697, n41698, n41699,
         n41700, n41701, n41702, n41703, n41704, n41705, n41706, n41707,
         n41708, n41709, n41710, n41711, n41712, n41713, n41714, n41715,
         n41716, n41717, n41718, n41719, n41720, n41721, n41722, n41723,
         n41724, n41725, n41726, n41727, n41728, n41729, n41730, n41731,
         n41732, n41733, n41734, n41735, n41736, n41737, n41738, n41739,
         n41740, n41741, n41742, n41743, n41744, n41745, n41746, n41747,
         n41748, n41749, n41750, n41751, n41752, n41753, n41754, n41755,
         n41756, n41757, n41758, n41759, n41760, n41761, n41762, n41763,
         n41764, n41765, n41766, n41767, n41768, n41769, n41770, n41771,
         n41772, n41773, n41774, n41775, n41776, n41777, n41778, n41779,
         n41780, n41781, n41782, n41783, n41784, n41785, n41786, n41787,
         n41788, n41789, n41790, n41791, n41792, n41793, n41794, n41795,
         n41796, n41797, n41798, n41799, n41800, n41801, n41802, n41803,
         n41804, n41805, n41806, n41807, n41808, n41809, n41810, n41811,
         n41812, n41813, n41814, n41815, n41816, n41817, n41818, n41819,
         n41820, n41821, n41822, n41823, n41824, n41825, n41826, n41827,
         n41828, n41829, n41830, n41831, n41832, n41833, n41834, n41835,
         n41836, n41837, n41838, n41839, n41840, n41841, n41842, n41843,
         n41844, n41845, n41846, n41847, n41848, n41849, n41850, n41851,
         n41852, n41853, n41854, n41855, n41856, n41857, n41858, n41859,
         n41860, n41861, n41862, n41863, n41864, n41865, n41866, n41867,
         n41868, n41869, n41870, n41871, n41872, n41873, n41874, n41875,
         n41876, n41877, n41878, n41879, n41880, n41881, n41882, n41883,
         n41884, n41885, n41886, n41887, n41888, n41889, n41890, n41891,
         n41892, n41893, n41894, n41895, n41896, n41897, n41898, n41899,
         n41900, n41901, n41902, n41903, n41904, n41905, n41906, n41907,
         n41908, n41909, n41910, n41911, n41912, n41913, n41914, n41915,
         n41916, n41917, n41918, n41919, n41920, n41921, n41922, n41923,
         n41924, n41925, n41926, n41927, n41928, n41929, n41930, n41931,
         n41932, n41933, n41934, n41935, n41936, n41937, n41938, n41939,
         n41940, n41941, n41942, n41943, n41944, n41945, n41946, n41947,
         n41948, n41949, n41950, n41951, n41952, n41953, n41954, n41955,
         n41956, n41957, n41958, n41959, n41960, n41961, n41962, n41963,
         n41964, n41965, n41966, n41967, n41968, n41969, n41970, n41971,
         n41972, n41973, n41974, n41975, n41976, n41977, n41978, n41979,
         n41980, n41981, n41982, n41983, n41984, n41985, n41986, n41987,
         n41988, n41989, n41990, n41991, n41992, n41993, n41994, n41995,
         n41996, n41997, n41998, n41999, n42000, n42001, n42002, n42003,
         n42004, n42005, n42006, n42007, n42008, n42009, n42010, n42011,
         n42012, n42013, n42014, n42015, n42016, n42017, n42018, n42019,
         n42020, n42021, n42022, n42023, n42024, n42025, n42026, n42027,
         n42028, n42029, n42030, n42031, n42032, n42033, n42034, n42035,
         n42036, n42037, n42038, n42039, n42040, n42041, n42042, n42043,
         n42044, n42045, n42046, n42047, n42048, n42049, n42050, n42051,
         n42052, n42053, n42054, n42055, n42056, n42057, n42058, n42059,
         n42060, n42061, n42062, n42063, n42064, n42065, n42066, n42067,
         n42068, n42069, n42070, n42071, n42072, n42073, n42074, n42075,
         n42076, n42077, n42078, n42079, n42080, n42081, n42082, n42083,
         n42084, n42085, n42086, n42087, n42088, n42089, n42090, n42091,
         n42092, n42093, n42094, n42095, n42096, n42097, n42098, n42099,
         n42100, n42101, n42102, n42103, n42104, n42105, n42106, n42107,
         n42108, n42109, n42110, n42111, n42112, n42113, n42114, n42115,
         n42116, n42117, n42118, n42119, n42120, n42121, n42122, n42123,
         n42124, n42125, n42126, n42127, n42128, n42129, n42130, n42131,
         n42132, n42133, n42134, n42135, n42136, n42137, n42138, n42139,
         n42140, n42141, n42142, n42143, n42144, n42145, n42146, n42147,
         n42148, n42149, n42150, n42151, n42152, n42153, n42154, n42155,
         n42156, n42157, n42158, n42159, n42160, n42161, n42162, n42163,
         n42164, n42165, n42166, n42167, n42168, n42169, n42170, n42171,
         n42172, n42173, n42174, n42175, n42176, n42177, n42178, n42179,
         n42180, n42181, n42182, n42183, n42184, n42185, n42186, n42187,
         n42188, n42189, n42190, n42191, n42192, n42193, n42194, n42195,
         n42196, n42197, n42198, n42199, n42200, n42201, n42202, n42203,
         n42204, n42205, n42206, n42207, n42208, n42209, n42210, n42211,
         n42212, n42213, n42214, n42215, n42216, n42217, n42218, n42219,
         n42220, n42221, n42222, n42223, n42224, n42225, n42226, n42227,
         n42228, n42229, n42230, n42231, n42232, n42233, n42234, n42235,
         n42236, n42237, n42238, n42239, n42240, n42241, n42242, n42243,
         n42244, n42245, n42246, n42247, n42248, n42249, n42250, n42251,
         n42252, n42253, n42254, n42255, n42256, n42257, n42258, n42259,
         n42260, n42261, n42262, n42263, n42264, n42265, n42266, n42267,
         n42268, n42269, n42270, n42271, n42272, n42273, n42274, n42275,
         n42276, n42277, n42278, n42279, n42280, n42281, n42282, n42283,
         n42284, n42285, n42286, n42287, n42288, n42289, n42290, n42291,
         n42292, n42293, n42294, n42295, n42296, n42297, n42298, n42299,
         n42300, n42301, n42302, n42303, n42304, n42305, n42306, n42307,
         n42308, n42309, n42310, n42311, n42312, n42313, n42314, n42315,
         n42316, n42317, n42318, n42319, n42320, n42321, n42322, n42323,
         n42324, n42325, n42326, n42327, n42328, n42329, n42330, n42331,
         n42332, n42333, n42334, n42335, n42336, n42337, n42338, n42339,
         n42340, n42341, n42342, n42343, n42344, n42345, n42346, n42347,
         n42348, n42349, n42350, n42351, n42352, n42353, n42354, n42355,
         n42356, n42357, n42358, n42359, n42360, n42361, n42362, n42363,
         n42364, n42365, n42366, n42367, n42368, n42369, n42370, n42371,
         n42372, n42373, n42374, n42375, n42376, n42377, n42378, n42379,
         n42380, n42381, n42382, n42383, n42384, n42385, n42386, n42387,
         n42388, n42389, n42390, n42391, n42392, n42393, n42394, n42395,
         n42396, n42397, n42398, n42399, n42400, n42401, n42402, n42403,
         n42404, n42405, n42406, n42407, n42408, n42409, n42410, n42411,
         n42412, n42413, n42414, n42415, n42416, n42417, n42418, n42419,
         n42420, n42421, n42422, n42423, n42424, n42425, n42426, n42427,
         n42428, n42429, n42430, n42431, n42432, n42433, n42434, n42435,
         n42436, n42437, n42438, n42439, n42440, n42441, n42442, n42443,
         n42444, n42445, n42446, n42447, n42448, n42449, n42450, n42451,
         n42452, n42453, n42454, n42455, n42456, n42457, n42458, n42459,
         n42460, n42461, n42462, n42463, n42464, n42465, n42466, n42467,
         n42468, n42469, n42470, n42471, n42472, n42473, n42474, n42475,
         n42476, n42477, n42478, n42479, n42480, n42481, n42482, n42483,
         n42484, n42485, n42486, n42487, n42488, n42489, n42490, n42491,
         n42492, n42493, n42494, n42495, n42496, n42497, n42498, n42499,
         n42500, n42501, n42502, n42503, n42504, n42505, n42506, n42507,
         n42508, n42509, n42510, n42511, n42512, n42513, n42514, n42515,
         n42516, n42517, n42518, n42519, n42520, n42521, n42522, n42523,
         n42524, n42525, n42526, n42527, n42528, n42529, n42530, n42531,
         n42532, n42533, n42534, n42535, n42536, n42537, n42538, n42539,
         n42540, n42541, n42542, n42543, n42544, n42545, n42546, n42547,
         n42548, n42549, n42550, n42551, n42552, n42553, n42554, n42555,
         n42556, n42557, n42558, n42559, n42560, n42561, n42562, n42563,
         n42564, n42565, n42566, n42567, n42568, n42569, n42570, n42571,
         n42572, n42573, n42574, n42575, n42576, n42577, n42578, n42579,
         n42580, n42581, n42582, n42583, n42584, n42585, n42586, n42587,
         n42588, n42589, n42590, n42591, n42592, n42593, n42594, n42595,
         n42596, n42597, n42598, n42599, n42600, n42601, n42602, n42603,
         n42604, n42605, n42606, n42607, n42608, n42609, n42610, n42611,
         n42612, n42613, n42614, n42615, n42616, n42617, n42618, n42619,
         n42620, n42621, n42622, n42623, n42624, n42625, n42626, n42627,
         n42628, n42629, n42630, n42631, n42632, n42633, n42634, n42635,
         n42636, n42637, n42638, n42639, n42640, n42641, n42642, n42643,
         n42644, n42645, n42646, n42647, n42648, n42649, n42650, n42651,
         n42652, n42653, n42654, n42655, n42656, n42657, n42658, n42659,
         n42660, n42661, n42662, n42663, n42664, n42665, n42666, n42667,
         n42668, n42669, n42670, n42671, n42672, n42673, n42674, n42675,
         n42676, n42677, n42678, n42679, n42680, n42681, n42682, n42683,
         n42684, n42685, n42686, n42687, n42688, n42689, n42690, n42691,
         n42692, n42693, n42694, n42695, n42696, n42697, n42698, n42699,
         n42700, n42701, n42702, n42703, n42704, n42705, n42706, n42707,
         n42708, n42709, n42710, n42711, n42712, n42713, n42714, n42715,
         n42716, n42717, n42718, n42719, n42720, n42721, n42722, n42723,
         n42724, n42725, n42726, n42727, n42728, n42729, n42730, n42731,
         n42732, n42733, n42734, n42735, n42736, n42737, n42738, n42739,
         n42740, n42741, n42742, n42743, n42744, n42745, n42746, n42747,
         n42748, n42749, n42750, n42751, n42752, n42753, n42754, n42755,
         n42756, n42757, n42758, n42759, n42760, n42761, n42762, n42763,
         n42764, n42765, n42766, n42767, n42768, n42769, n42770, n42771,
         n42772, n42773, n42774, n42775, n42776, n42777, n42778, n42779,
         n42780, n42781, n42782, n42783, n42784, n42785, n42786, n42787,
         n42788, n42789, n42790, n42791, n42792, n42793, n42794, n42795,
         n42796, n42797, n42798, n42799, n42800, n42801, n42802, n42803,
         n42804, n42805, n42806, n42807, n42808, n42809, n42810, n42811,
         n42812, n42813, n42814, n42815, n42816, n42817, n42818, n42819,
         n42820, n42821, n42822, n42823, n42824, n42825, n42826, n42827,
         n42828, n42829, n42830, n42831, n42832, n42833, n42834, n42835,
         n42836, n42837, n42838, n42839, n42840, n42841, n42842, n42843,
         n42844, n42845, n42846, n42847, n42848, n42849, n42850, n42851,
         n42852, n42853, n42854, n42855, n42856, n42857, n42858, n42859,
         n42860, n42861, n42862, n42863, n42864, n42865, n42866, n42867,
         n42868, n42869, n42870, n42871, n42872, n42873, n42874, n42875,
         n42876, n42877, n42878, n42879, n42880, n42881, n42882, n42883,
         n42884, n42885, n42886, n42887, n42888, n42889, n42890, n42891,
         n42892, n42893, n42894, n42895, n42896, n42897, n42898, n42899,
         n42900, n42901, n42902, n42903, n42904, n42905, n42906, n42907,
         n42908, n42909, n42910, n42911, n42912, n42913, n42914, n42915,
         n42916, n42917, n42918, n42919, n42920, n42921, n42922, n42923,
         n42924, n42925, n42926, n42927, n42928, n42929, n42930, n42931,
         n42932, n42933, n42934, n42935, n42936, n42937, n42938, n42939,
         n42940, n42941, n42942, n42943, n42944, n42945, n42946, n42947,
         n42948, n42949, n42950, n42951, n42952, n42953, n42954, n42955,
         n42956, n42957, n42958, n42959, n42960, n42961, n42962, n42963,
         n42964, n42965, n42966, n42967, n42968, n42969, n42970, n42971,
         n42972, n42973, n42974, n42975, n42976, n42977, n42978, n42979,
         n42980, n42981, n42982, n42983, n42984, n42985, n42986, n42987,
         n42988, n42989, n42990, n42991, n42992, n42993, n42994, n42995,
         n42996, n42997, n42998, n42999, n43000, n43001, n43002, n43003,
         n43004, n43005, n43006, n43007, n43008, n43009, n43010, n43011,
         n43012, n43013, n43014, n43015, n43016, n43017, n43018, n43019,
         n43020, n43021, n43022, n43023, n43024, n43025, n43026, n43027,
         n43028, n43029, n43030, n43031, n43032, n43033, n43034, n43035,
         n43036, n43037, n43038, n43039, n43040, n43041, n43042, n43043,
         n43044, n43045, n43046, n43047, n43048, n43049, n43050, n43051,
         n43052, n43053, n43054, n43055, n43056, n43057, n43058, n43059,
         n43060, n43061, n43062, n43063, n43064, n43065, n43066, n43067,
         n43068, n43069, n43070, n43071, n43072, n43073, n43074, n43075,
         n43076, n43077, n43078, n43079, n43080, n43081, n43082, n43083,
         n43084, n43085, n43086, n43087, n43088, n43089, n43090, n43091,
         n43092, n43093, n43094, n43095, n43096, n43097, n43098, n43099,
         n43100, n43101, n43102, n43103, n43104, n43105, n43106, n43107,
         n43108, n43109, n43110, n43111, n43112, n43113, n43114, n43115,
         n43116, n43117, n43118, n43119, n43120, n43121, n43122, n43123,
         n43124, n43125, n43126, n43127, n43128, n43129, n43130, n43131,
         n43132, n43133, n43134, n43135, n43136, n43137, n43138, n43139,
         n43140, n43141, n43142, n43143, n43144, n43145, n43146, n43147,
         n43148, n43149, n43150, n43151, n43152, n43153, n43154, n43155,
         n43156, n43157, n43158, n43159, n43160, n43161, n43162, n43163,
         n43164, n43165, n43166, n43167, n43168, n43169, n43170, n43171,
         n43172, n43173, n43174, n43175, n43176, n43177, n43178, n43179,
         n43180, n43181, n43182, n43183, n43184, n43185, n43186, n43187,
         n43188, n43189, n43190, n43191, n43192, n43193, n43194, n43195,
         n43196, n43197, n43198, n43199, n43200, n43201, n43202, n43203,
         n43204, n43205, n43206, n43207, n43208, n43209, n43210, n43211,
         n43212, n43213, n43214, n43215, n43216, n43217, n43218, n43219,
         n43220, n43221, n43222, n43223, n43224, n43225, n43226, n43227,
         n43228, n43229, n43230, n43231, n43232, n43233, n43234, n43235,
         n43236, n43237, n43238, n43239, n43240, n43241, n43242, n43243,
         n43244, n43245, n43246, n43247, n43248, n43249, n43250, n43251,
         n43252, n43253, n43254, n43255, n43256, n43257, n43258, n43259,
         n43260, n43261, n43262, n43263, n43264, n43265, n43266, n43267,
         n43268, n43269, n43270, n43271, n43272, n43273, n43274, n43275,
         n43276, n43277, n43278, n43279, n43280, n43281, n43282, n43283,
         n43284, n43285, n43286, n43287, n43288, n43289, n43290, n43291,
         n43292, n43293, n43294, n43295, n43296, n43297, n43298, n43299,
         n43300, n43301, n43302, n43303, n43304, n43305, n43306, n43307,
         n43308, n43309, n43310, n43311, n43312, n43313, n43314, n43315,
         n43316, n43317, n43318, n43319, n43320, n43321, n43322, n43323,
         n43324, n43325, n43326, n43327, n43328, n43329, n43330, n43331,
         n43332, n43333, n43334, n43335, n43336, n43337, n43338, n43339,
         n43340, n43341, n43342, n43343, n43344, n43345, n43346, n43347,
         n43348, n43349, n43350, n43351, n43352, n43353, n43354, n43355,
         n43356, n43357, n43358, n43359, n43360, n43361, n43362, n43363,
         n43364, n43365, n43366, n43367, n43368, n43369, n43370, n43371,
         n43372, n43373, n43374, n43375, n43376, n43377, n43378, n43379,
         n43380, n43381, n43382, n43383, n43384, n43385, n43386, n43387,
         n43388, n43389, n43390, n43391, n43392, n43393, n43394, n43395,
         n43396, n43397, n43398, n43399, n43400, n43401, n43402, n43403,
         n43404, n43405, n43406, n43407, n43408, n43409, n43410, n43411,
         n43412, n43413, n43414, n43415, n43416, n43417, n43418, n43419,
         n43420, n43421, n43422, n43423, n43424, n43425, n43426, n43427,
         n43428, n43429, n43430, n43431, n43432, n43433, n43434, n43435,
         n43436, n43437, n43438, n43439, n43440, n43441, n43442, n43443,
         n43444, n43445, n43446, n43447, n43448, n43449, n43450, n43451,
         n43452, n43453, n43454, n43455, n43456, n43457, n43458, n43459,
         n43460, n43461, n43462, n43463, n43464, n43465, n43466, n43467,
         n43468, n43469, n43470, n43471, n43472, n43473, n43474, n43475,
         n43476, n43477, n43478, n43479, n43480, n43481, n43482, n43483,
         n43484, n43485, n43486, n43487, n43488, n43489, n43490, n43491,
         n43492, n43493, n43494, n43495, n43496, n43497, n43498, n43499,
         n43500, n43501, n43502, n43503, n43504, n43505, n43506, n43507,
         n43508, n43509, n43510, n43511, n43512, n43513, n43514, n43515,
         n43516, n43517, n43518, n43519, n43520, n43521, n43522, n43523,
         n43524, n43525, n43526, n43527, n43528, n43529, n43530, n43531,
         n43532, n43533, n43534, n43535, n43536, n43537, n43538, n43539,
         n43540, n43541, n43542, n43543, n43544, n43545, n43546, n43547,
         n43548, n43549, n43550, n43551, n43552, n43553, n43554, n43555,
         n43556, n43557, n43558, n43559, n43560, n43561, n43562, n43563,
         n43564, n43565, n43566, n43567, n43568, n43569, n43570, n43571,
         n43572, n43573, n43574, n43575, n43576, n43577, n43578, n43579,
         n43580, n43581, n43582, n43583, n43584, n43585, n43586, n43587,
         n43588, n43589, n43590, n43591, n43592, n43593, n43594, n43595,
         n43596, n43597, n43598, n43599, n43600, n43601, n43602, n43603,
         n43604, n43605, n43606, n43607, n43608, n43609, n43610, n43611,
         n43612, n43613, n43614, n43615, n43616, n43617, n43618, n43619,
         n43620, n43621, n43622, n43623, n43624, n43625, n43626, n43627,
         n43628, n43629, n43630, n43631, n43632, n43633, n43634, n43635,
         n43636, n43637, n43638, n43639, n43640, n43641, n43642, n43643,
         n43644, n43645, n43646, n43647, n43648, n43649, n43650, n43651,
         n43652, n43653, n43654, n43655, n43656, n43657, n43658, n43659,
         n43660, n43661, n43662, n43663, n43664, n43665, n43666, n43667,
         n43668, n43669, n43670, n43671, n43672, n43673, n43674, n43675,
         n43676, n43677, n43678, n43679, n43680, n43681, n43682, n43683,
         n43684, n43685, n43686, n43687, n43688, n43689, n43690, n43691,
         n43692, n43693, n43694, n43695, n43696, n43697, n43698, n43699,
         n43700, n43701, n43702, n43703, n43704, n43705, n43706, n43707,
         n43708, n43709, n43710, n43711, n43712, n43713, n43714, n43715,
         n43716, n43717, n43718, n43719, n43720, n43721, n43722, n43723,
         n43724, n43725, n43726, n43727, n43728, n43729, n43730, n43731,
         n43732, n43733, n43734, n43735, n43736, n43737, n43738, n43739,
         n43740, n43741, n43742, n43743, n43744, n43745, n43746, n43747,
         n43748, n43749, n43750, n43751, n43752, n43753, n43754, n43755,
         n43756, n43757, n43758, n43759, n43760, n43761, n43762, n43763,
         n43764, n43765, n43766, n43767, n43768, n43769, n43770, n43771,
         n43772, n43773, n43774, n43775, n43776, n43777, n43778, n43779,
         n43780, n43781, n43782, n43783, n43784, n43785, n43786, n43787,
         n43788, n43789, n43790, n43791, n43792, n43793, n43794, n43795,
         n43796, n43797, n43798, n43799, n43800, n43801, n43802, n43803,
         n43804, n43805, n43806, n43807, n43808, n43809, n43810, n43811,
         n43812, n43813, n43814, n43815, n43816, n43817, n43818, n43819,
         n43820, n43821, n43822, n43823, n43824, n43825, n43826, n43827,
         n43828, n43829, n43830, n43831, n43832, n43833, n43834, n43835,
         n43836, n43837, n43838, n43839, n43840, n43841, n43842, n43843,
         n43844, n43845, n43846, n43847, n43848, n43849, n43850, n43851,
         n43852, n43853, n43854, n43855, n43856, n43857, n43858, n43859,
         n43860, n43861, n43862, n43863, n43864, n43865, n43866, n43867,
         n43868, n43869, n43870, n43871, n43872, n43873, n43874, n43875,
         n43876, n43877, n43878, n43879, n43880, n43881, n43882, n43883,
         n43884, n43885, n43886, n43887, n43888, n43889, n43890, n43891,
         n43892, n43893, n43894, n43895, n43896, n43897, n43898, n43899,
         n43900, n43901, n43902, n43903, n43904, n43905, n43906, n43907,
         n43908, n43909, n43910, n43911, n43912, n43913, n43914, n43915,
         n43916, n43917, n43918, n43919, n43920, n43921, n43922, n43923,
         n43924, n43925, n43926, n43927, n43928, n43929, n43930, n43931,
         n43932, n43933, n43934, n43935, n43936, n43937, n43938, n43939,
         n43940, n43941, n43942, n43943, n43944, n43945, n43946, n43947,
         n43948, n43949, n43950, n43951, n43952, n43953, n43954, n43955,
         n43956, n43957, n43958, n43959, n43960, n43961, n43962, n43963,
         n43964, n43965, n43966, n43967, n43968, n43969, n43970, n43971,
         n43972, n43973, n43974, n43975, n43976, n43977, n43978, n43979,
         n43980, n43981, n43982, n43983, n43984, n43985, n43986, n43987,
         n43988, n43989, n43990, n43991, n43992, n43993, n43994, n43995,
         n43996, n43997, n43998, n43999, n44000, n44001, n44002, n44003,
         n44004, n44005, n44006, n44007, n44008, n44009, n44010, n44011,
         n44012, n44013, n44014, n44015, n44016, n44017, n44018, n44019,
         n44020, n44021, n44022, n44023, n44024, n44025, n44026, n44027,
         n44028, n44029, n44030, n44031, n44032, n44033, n44034, n44035,
         n44036, n44037, n44038, n44039, n44040, n44041, n44042, n44043,
         n44044, n44045, n44046, n44047, n44048, n44049, n44050, n44051,
         n44052, n44053, n44054, n44055, n44056, n44057, n44058, n44059,
         n44060, n44061, n44062, n44063, n44064, n44065, n44066, n44067,
         n44068, n44069, n44070, n44071, n44072, n44073, n44074, n44075,
         n44076, n44077, n44078, n44079, n44080, n44081, n44082, n44083,
         n44084, n44085, n44086, n44087, n44088, n44089, n44090, n44091,
         n44092, n44093, n44094, n44095, n44096, n44097, n44098, n44099,
         n44100, n44101, n44102, n44103, n44104, n44105, n44106, n44107,
         n44108, n44109, n44110, n44111, n44112, n44113, n44114, n44115,
         n44116, n44117, n44118, n44119, n44120, n44121, n44122, n44123,
         n44124, n44125, n44126, n44127, n44128, n44129, n44130, n44131,
         n44132, n44133, n44134, n44135, n44136, n44137, n44138, n44139,
         n44140, n44141, n44142, n44143, n44144, n44145, n44146, n44147,
         n44148, n44149, n44150, n44151, n44152, n44153, n44154, n44155,
         n44156, n44157, n44158, n44159, n44160, n44161, n44162, n44163,
         n44164, n44165, n44166, n44167, n44168, n44169, n44170, n44171,
         n44172, n44173, n44174, n44175, n44176, n44177, n44178, n44179,
         n44180, n44181, n44182, n44183, n44184, n44185, n44186, n44187,
         n44188, n44189, n44190, n44191, n44192, n44193, n44194, n44195,
         n44196, n44197, n44198, n44199, n44200, n44201, n44202, n44203,
         n44204, n44205, n44206, n44207, n44208, n44209, n44210, n44211,
         n44212, n44213, n44214, n44215, n44216, n44217, n44218, n44219,
         n44220, n44221, n44222, n44223, n44224, n44225, n44226, n44227,
         n44228, n44229, n44230, n44231, n44232, n44233, n44234, n44235,
         n44236, n44237, n44238, n44239, n44240, n44241, n44242, n44243,
         n44244, n44245, n44246, n44247, n44248, n44249, n44250, n44251,
         n44252, n44253, n44254, n44255, n44256, n44257, n44258, n44259,
         n44260, n44261, n44262, n44263, n44264, n44265, n44266, n44267,
         n44268, n44269, n44270, n44271, n44272, n44273, n44274, n44275,
         n44276, n44277, n44278, n44279, n44280, n44281, n44282, n44283,
         n44284, n44285, n44286, n44287, n44288, n44289, n44290, n44291,
         n44292, n44293, n44294, n44295, n44296, n44297, n44298, n44299,
         n44300, n44301, n44302, n44303, n44304, n44305, n44306, n44307,
         n44308, n44309, n44310, n44311, n44312, n44313, n44314, n44315,
         n44316, n44317, n44318, n44319, n44320, n44321, n44322, n44323,
         n44324, n44325, n44326, n44327, n44328, n44329, n44330, n44331,
         n44332, n44333, n44334, n44335, n44336, n44337, n44338, n44339,
         n44340, n44341, n44342, n44343, n44344, n44345, n44346, n44347,
         n44348, n44349, n44350, n44351, n44352, n44353, n44354, n44355,
         n44356, n44357, n44358, n44359, n44360, n44361, n44362, n44363,
         n44364, n44365, n44366, n44367, n44368, n44369, n44370, n44371,
         n44372, n44373, n44374, n44375, n44376, n44377, n44378, n44379,
         n44380, n44381, n44382, n44383, n44384, n44385, n44386, n44387,
         n44388, n44389, n44390, n44391, n44392, n44393, n44394, n44395,
         n44396, n44397, n44398, n44399, n44400, n44401, n44402, n44403,
         n44404, n44405, n44406, n44407, n44408, n44409, n44410, n44411,
         n44412, n44413, n44414, n44415, n44416, n44417, n44418, n44419,
         n44420, n44421, n44422, n44423, n44424, n44425, n44426, n44427,
         n44428, n44429, n44430, n44431, n44432, n44433, n44434, n44435,
         n44436, n44437, n44438, n44439, n44440, n44441, n44442, n44443,
         n44444, n44445, n44446, n44447, n44448, n44449, n44450, n44451,
         n44452, n44453, n44454, n44455, n44456, n44457, n44458, n44459,
         n44460, n44461, n44462, n44463, n44464, n44465, n44466, n44467,
         n44468, n44469, n44470, n44471, n44472, n44473, n44474, n44475,
         n44476, n44477, n44478, n44479, n44480, n44481, n44482, n44483,
         n44484, n44485, n44486, n44487, n44488, n44489, n44490, n44491,
         n44492, n44493, n44494, n44495, n44496, n44497, n44498, n44499,
         n44500, n44501, n44502, n44503, n44504, n44505, n44506, n44507,
         n44508, n44509, n44510, n44511, n44512, n44513, n44514, n44515,
         n44516, n44517, n44518, n44519, n44520, n44521, n44522, n44523,
         n44524, n44525, n44526, n44527, n44528, n44529, n44530, n44531,
         n44532, n44533, n44534, n44535, n44536, n44537, n44538, n44539,
         n44540, n44541, n44542, n44543, n44544, n44545, n44546, n44547,
         n44548, n44549, n44550, n44551, n44552, n44553, n44554, n44555,
         n44556, n44557, n44558, n44559, n44560, n44561, n44562, n44563,
         n44564, n44565, n44566, n44567, n44568, n44569, n44570, n44571,
         n44572, n44573, n44574, n44575, n44576, n44577, n44578, n44579,
         n44580, n44581, n44582, n44583, n44584, n44585, n44586, n44587,
         n44588, n44589, n44590, n44591, n44592, n44593, n44594, n44595,
         n44596, n44597, n44598, n44599, n44600, n44601, n44602, n44603,
         n44604, n44605, n44606, n44607, n44608, n44609, n44610, n44611,
         n44612, n44613, n44614, n44615, n44616, n44617, n44618, n44619,
         n44620, n44621, n44622, n44623, n44624, n44625, n44626, n44627,
         n44628, n44629, n44630, n44631, n44632, n44633, n44634, n44635,
         n44636, n44637, n44638, n44639, n44640, n44641, n44642, n44643,
         n44644, n44645, n44646, n44647, n44648, n44649, n44650, n44651,
         n44652, n44653, n44654, n44655, n44656, n44657, n44658, n44659,
         n44660, n44661, n44662, n44663, n44664, n44665, n44666, n44667,
         n44668, n44669, n44670, n44671, n44672, n44673, n44674, n44675,
         n44676, n44677, n44678, n44679, n44680, n44681, n44682, n44683,
         n44684, n44685, n44686, n44687, n44688, n44689, n44690, n44691,
         n44692, n44693, n44694, n44695, n44696, n44697, n44698, n44699,
         n44700, n44701, n44702, n44703, n44704, n44705, n44706, n44707,
         n44708, n44709, n44710, n44711, n44712, n44713, n44714, n44715,
         n44716, n44717, n44718, n44719, n44720, n44721, n44722, n44723,
         n44724, n44725, n44726, n44727, n44728, n44729, n44730, n44731,
         n44732, n44733, n44734, n44735, n44736, n44737, n44738, n44739,
         n44740, n44741, n44742, n44743, n44744, n44745, n44746, n44747,
         n44748, n44749, n44750, n44751, n44752, n44753, n44754, n44755,
         n44756, n44757, n44758, n44759, n44760, n44761, n44762, n44763,
         n44764, n44765, n44766, n44767, n44768, n44769, n44770, n44771,
         n44772, n44773, n44774, n44775, n44776, n44777, n44778, n44779,
         n44780, n44781, n44782, n44783, n44784, n44785, n44786, n44787,
         n44788, n44789, n44790, n44791, n44792, n44793, n44794, n44795,
         n44796, n44797, n44798, n44799, n44800, n44801, n44802, n44803,
         n44804, n44805, n44806, n44807, n44808, n44809, n44810, n44811,
         n44812, n44813, n44814, n44815, n44816, n44817, n44818, n44819,
         n44820, n44821, n44822, n44823, n44824, n44825, n44826, n44827,
         n44828, n44829, n44830, n44831, n44832, n44833, n44834, n44835,
         n44836, n44837, n44838, n44839, n44840, n44841, n44842, n44843,
         n44844, n44845, n44846, n44847, n44848, n44849, n44850, n44851,
         n44852, n44853, n44854, n44855, n44856, n44857, n44858, n44859,
         n44860, n44861, n44862, n44863, n44864, n44865, n44866, n44867,
         n44868, n44869, n44870, n44871, n44872, n44873, n44874, n44875,
         n44876, n44877, n44878, n44879, n44880, n44881, n44882, n44883,
         n44884, n44885, n44886, n44887, n44888, n44889, n44890, n44891,
         n44892, n44893, n44894, n44895, n44896, n44897, n44898, n44899,
         n44900, n44901, n44902, n44903, n44904, n44905, n44906, n44907,
         n44908, n44909, n44910, n44911, n44912, n44913, n44914, n44915,
         n44916, n44917, n44918, n44919, n44920, n44921, n44922, n44923,
         n44924, n44925, n44926, n44927, n44928, n44929, n44930, n44931,
         n44932, n44933, n44934, n44935, n44936, n44937, n44938, n44939,
         n44940, n44941, n44942, n44943, n44944, n44945, n44946, n44947,
         n44948, n44949, n44950, n44951, n44952, n44953, n44954, n44955,
         n44956, n44957, n44958, n44959, n44960, n44961, n44962, n44963,
         n44964, n44965, n44966, n44967, n44968, n44969, n44970, n44971,
         n44972, n44973, n44974, n44975, n44976, n44977, n44978, n44979,
         n44980, n44981, n44982, n44983, n44984, n44985, n44986, n44987,
         n44988, n44989, n44990, n44991, n44992, n44993, n44994, n44995,
         n44996, n44997, n44998, n44999, n45000, n45001, n45002, n45003,
         n45004, n45005, n45006, n45007, n45008, n45009, n45010, n45011,
         n45012, n45013, n45014, n45015, n45016, n45017, n45018, n45019,
         n45020, n45021, n45022, n45023, n45024, n45025, n45026, n45027,
         n45028, n45029, n45030, n45031, n45032, n45033, n45034, n45035,
         n45036, n45037, n45038, n45039, n45040, n45041, n45042, n45043,
         n45044, n45045, n45046, n45047, n45048, n45049, n45050, n45051,
         n45052, n45053, n45054, n45055, n45056, n45057, n45058, n45059,
         n45060, n45061, n45062, n45063, n45064, n45065, n45066, n45067,
         n45068, n45069, n45070, n45071, n45072, n45073, n45074, n45075,
         n45076, n45077, n45078, n45079, n45080, n45081, n45082, n45083,
         n45084, n45085, n45086, n45087, n45088, n45089, n45090, n45091,
         n45092, n45093, n45094, n45095, n45096, n45097, n45098, n45099,
         n45100, n45101, n45102, n45103, n45104, n45105, n45106, n45107,
         n45108, n45109, n45110, n45111, n45112, n45113, n45114, n45115,
         n45116, n45117, n45118, n45119, n45120, n45121, n45122, n45123,
         n45124, n45125, n45126, n45127, n45128, n45129, n45130, n45131,
         n45132, n45133, n45134, n45135, n45136, n45137, n45138, n45139,
         n45140, n45141, n45142, n45143, n45144, n45145, n45146, n45147,
         n45148, n45149, n45150, n45151, n45152, n45153, n45154, n45155,
         n45156, n45157, n45158, n45159, n45160, n45161, n45162, n45163,
         n45164, n45165, n45166, n45167, n45168, n45169, n45170, n45171,
         n45172, n45173, n45174, n45175, n45176, n45177, n45178, n45179,
         n45180, n45181, n45182, n45183, n45184, n45185, n45186, n45187,
         n45188, n45189, n45190, n45191, n45192, n45193, n45194, n45195,
         n45196, n45197, n45198, n45199, n45200, n45201, n45202, n45203,
         n45204, n45205, n45206, n45207, n45208, n45209, n45210, n45211,
         n45212, n45213, n45214, n45215, n45216, n45217, n45218, n45219,
         n45220, n45221, n45222, n45223, n45224, n45225, n45226, n45227,
         n45228, n45229, n45230, n45231, n45232, n45233, n45234, n45235,
         n45236, n45237, n45238, n45239, n45240, n45241, n45242, n45243,
         n45244, n45245, n45246, n45247, n45248, n45249, n45250, n45251,
         n45252, n45253, n45254, n45255, n45256, n45257, n45258, n45259,
         n45260, n45261, n45262, n45263, n45264, n45265, n45266, n45267,
         n45268, n45269, n45270, n45271, n45272, n45273, n45274, n45275,
         n45276, n45277, n45278, n45279, n45280, n45281, n45282, n45283,
         n45284, n45285, n45286, n45287, n45288, n45289, n45290, n45291,
         n45292, n45293, n45294, n45295, n45296, n45297, n45298, n45299,
         n45300, n45301, n45302, n45303, n45304, n45305, n45306, n45307,
         n45308, n45309, n45310, n45311, n45312, n45313, n45314, n45315,
         n45316, n45317, n45318, n45319, n45320, n45321, n45322, n45323,
         n45324, n45325, n45326, n45327, n45328, n45329, n45330, n45331,
         n45332, n45333, n45334, n45335, n45336, n45337, n45338, n45339,
         n45340, n45341, n45342, n45343, n45344, n45345, n45346, n45347,
         n45348, n45349, n45350, n45351, n45352, n45353, n45354, n45355,
         n45356, n45357, n45358, n45359, n45360, n45361, n45362, n45363,
         n45364, n45365, n45366, n45367, n45368, n45369, n45370, n45371,
         n45372, n45373, n45374, n45375, n45376, n45377, n45378, n45379,
         n45380, n45381, n45382, n45383, n45384, n45385, n45386, n45387,
         n45388, n45389, n45390, n45391, n45392, n45393, n45394, n45395,
         n45396, n45397, n45398, n45399, n45400, n45401, n45402, n45403,
         n45404, n45405, n45406, n45407, n45408, n45409, n45410, n45411,
         n45412, n45413, n45414, n45415, n45416, n45417, n45418, n45419,
         n45420, n45421, n45422, n45423, n45424, n45425, n45426, n45427,
         n45428, n45429, n45430, n45431, n45432, n45433, n45434, n45435,
         n45436, n45437, n45438, n45439, n45440, n45441, n45442, n45443,
         n45444, n45445, n45446, n45447, n45448, n45449, n45450, n45451,
         n45452, n45453, n45454, n45455, n45456, n45457, n45458, n45459,
         n45460, n45461, n45462, n45463, n45464, n45465, n45466, n45467,
         n45468, n45469, n45470, n45471, n45472, n45473, n45474, n45475,
         n45476, n45477, n45478, n45479, n45480, n45481, n45482, n45483,
         n45484, n45485, n45486, n45487, n45488, n45489, n45490, n45491,
         n45492, n45493, n45494, n45495, n45496, n45497, n45498, n45499,
         n45500, n45501, n45502, n45503, n45504, n45505, n45506, n45507,
         n45508, n45509, n45510, n45511, n45512, n45513, n45514, n45515,
         n45516, n45517, n45518, n45519, n45520, n45521, n45522, n45523,
         n45524, n45525, n45526, n45527, n45528, n45529, n45530, n45531,
         n45532, n45533, n45534, n45535, n45536, n45537, n45538, n45539,
         n45540, n45541, n45542, n45543, n45544, n45545, n45546, n45547,
         n45548, n45549, n45550, n45551, n45552, n45553, n45554, n45555,
         n45556, n45557, n45558, n45559, n45560, n45561, n45562, n45563,
         n45564, n45565, n45566, n45567, n45568, n45569, n45570, n45571,
         n45572, n45573, n45574, n45575, n45576, n45577, n45578, n45579,
         n45580, n45581, n45582, n45583, n45584, n45585, n45586, n45587,
         n45588, n45589, n45590, n45591, n45592, n45593, n45594, n45595,
         n45596, n45597, n45598, n45599, n45600, n45601, n45602, n45603,
         n45604, n45605, n45606, n45607, n45608, n45609, n45610, n45611,
         n45612, n45613, n45614, n45615, n45616, n45617, n45618, n45619,
         n45620, n45621, n45622, n45623, n45624, n45625, n45626, n45627,
         n45628, n45629, n45630, n45631, n45632, n45633, n45634, n45635,
         n45636, n45637, n45638, n45639, n45640, n45641, n45642, n45643,
         n45644, n45645, n45646, n45647, n45648, n45649, n45650, n45651,
         n45652, n45653, n45654, n45655, n45656, n45657, n45658, n45659,
         n45660, n45661, n45662, n45663, n45664, n45665, n45666, n45667,
         n45668, n45669, n45670, n45671, n45672, n45673, n45674, n45675,
         n45676, n45677, n45678, n45679, n45680, n45681, n45682, n45683,
         n45684, n45685, n45686, n45687, n45688, n45689, n45690, n45691,
         n45692, n45693, n45694, n45695, n45696, n45697, n45698, n45699,
         n45700, n45701, n45702, n45703, n45704, n45705, n45706, n45707,
         n45708, n45709, n45710, n45711, n45712, n45713, n45714, n45715,
         n45716, n45717, n45718, n45719, n45720, n45721, n45722, n45723,
         n45724, n45725, n45726, n45727, n45728, n45729, n45730, n45731,
         n45732, n45733, n45734, n45735, n45736, n45737, n45738, n45739,
         n45740, n45741, n45742, n45743, n45744, n45745, n45746, n45747,
         n45748, n45749, n45750, n45751, n45752, n45753, n45754, n45755,
         n45756, n45757, n45758, n45759, n45760, n45761, n45762, n45763,
         n45764, n45765, n45766, n45767, n45768, n45769, n45770, n45771,
         n45772, n45773, n45774, n45775, n45776, n45777, n45778, n45779,
         n45780, n45781, n45782, n45783, n45784, n45785, n45786, n45787,
         n45788, n45789, n45790, n45791, n45792, n45793, n45794, n45795,
         n45796, n45797, n45798, n45799, n45800, n45801, n45802, n45803,
         n45804, n45805, n45806, n45807, n45808, n45809, n45810, n45811,
         n45812, n45813, n45814, n45815, n45816, n45817, n45818, n45819,
         n45820, n45821, n45822, n45823, n45824, n45825, n45826, n45827,
         n45828, n45829, n45830, n45831, n45832, n45833, n45834, n45835,
         n45836, n45837, n45838, n45839, n45840, n45841, n45842, n45843,
         n45844, n45845, n45846, n45847, n45848, n45849, n45850, n45851,
         n45852, n45853, n45854, n45855, n45856, n45857, n45858, n45859,
         n45860, n45861, n45862, n45863, n45864, n45865, n45866, n45867,
         n45868, n45869, n45870, n45871, n45872, n45873, n45874, n45875,
         n45876, n45877, n45878, n45879, n45880, n45881, n45882, n45883,
         n45884, n45885, n45886, n45887, n45888, n45889, n45890, n45891,
         n45892, n45893, n45894, n45895, n45896, n45897, n45898, n45899,
         n45900, n45901, n45902, n45903, n45904, n45905, n45906, n45907,
         n45908, n45909, n45910, n45911, n45912, n45913, n45914, n45915,
         n45916, n45917, n45918, n45919, n45920, n45921, n45922, n45923,
         n45924, n45925, n45926, n45927, n45928, n45929, n45930, n45931,
         n45932, n45933, n45934, n45935, n45936, n45937, n45938, n45939,
         n45940, n45941, n45942, n45943, n45944, n45945, n45946, n45947,
         n45948, n45949, n45950, n45951, n45952, n45953, n45954, n45955,
         n45956, n45957, n45958, n45959, n45960, n45961, n45962, n45963,
         n45964, n45965, n45966, n45967, n45968, n45969, n45970, n45971,
         n45972, n45973, n45974, n45975, n45976, n45977, n45978, n45979,
         n45980, n45981, n45982, n45983, n45984, n45985, n45986, n45987,
         n45988, n45989, n45990, n45991, n45992, n45993, n45994, n45995,
         n45996, n45997, n45998, n45999, n46000, n46001, n46002, n46003,
         n46004, n46005, n46006, n46007, n46008, n46009, n46010, n46011,
         n46012, n46013, n46014, n46015, n46016, n46017, n46018, n46019,
         n46020, n46021, n46022, n46023, n46024, n46025, n46026, n46027,
         n46028, n46029, n46030, n46031, n46032, n46033, n46034, n46035,
         n46036, n46037, n46038, n46039, n46040, n46041, n46042, n46043,
         n46044, n46045, n46046, n46047, n46048, n46049, n46050, n46051,
         n46052, n46053, n46054, n46055, n46056, n46057, n46058, n46059,
         n46060, n46061, n46062, n46063, n46064, n46065, n46066, n46067,
         n46068, n46069, n46070, n46071, n46072, n46073, n46074, n46075,
         n46076, n46077, n46078, n46079, n46080, n46081, n46082, n46083,
         n46084, n46085, n46086, n46087, n46088, n46089, n46090, n46091,
         n46092, n46093, n46094, n46095, n46096, n46097, n46098, n46099,
         n46100, n46101, n46102, n46103, n46104, n46105, n46106, n46107,
         n46108, n46109, n46110, n46111, n46112, n46113, n46114, n46115,
         n46116, n46117, n46118, n46119, n46120, n46121, n46122, n46123,
         n46124, n46125, n46126, n46127, n46128, n46129, n46130, n46131,
         n46132, n46133, n46134, n46135, n46136, n46137, n46138, n46139,
         n46140, n46141, n46142, n46143, n46144, n46145, n46146, n46147,
         n46148, n46149, n46150, n46151, n46152, n46153, n46154, n46155,
         n46156, n46157, n46158, n46159, n46160, n46161, n46162, n46163,
         n46164, n46165, n46166, n46167, n46168, n46169, n46170, n46171,
         n46172, n46173, n46174, n46175, n46176, n46177, n46178, n46179,
         n46180, n46181, n46182, n46183, n46184, n46185, n46186, n46187,
         n46188, n46189, n46190, n46191, n46192, n46193, n46194, n46195,
         n46196, n46197, n46198, n46199, n46200, n46201, n46202, n46203,
         n46204, n46205, n46206, n46207, n46208, n46209, n46210, n46211,
         n46212, n46213, n46214, n46215, n46216, n46217, n46218, n46219,
         n46220, n46221, n46222, n46223, n46224, n46225, n46226, n46227,
         n46228, n46229, n46230, n46231, n46232, n46233, n46234, n46235,
         n46236, n46237, n46238, n46239, n46240, n46241, n46242, n46243,
         n46244, n46245, n46246, n46247, n46248, n46249, n46250, n46251,
         n46252, n46253, n46254, n46255, n46256, n46257, n46258, n46259,
         n46260, n46261, n46262, n46263, n46264, n46265, n46266, n46267,
         n46268, n46269, n46270, n46271, n46272, n46273, n46274, n46275,
         n46276, n46277, n46278, n46279, n46280, n46281, n46282, n46283,
         n46284, n46285, n46286, n46287, n46288, n46289, n46290, n46291,
         n46292, n46293, n46294, n46295, n46296, n46297, n46298, n46299,
         n46300, n46301, n46302, n46303, n46304, n46305, n46306, n46307,
         n46308, n46309, n46310, n46311, n46312, n46313, n46314, n46315,
         n46316, n46317, n46318, n46319, n46320, n46321, n46322, n46323,
         n46324, n46325, n46326, n46327, n46328, n46329, n46330, n46331,
         n46332, n46333, n46334, n46335, n46336, n46337, n46338, n46339,
         n46340, n46341, n46342, n46343, n46344, n46345, n46346, n46347,
         n46348, n46349, n46350, n46351, n46352, n46353, n46354, n46355,
         n46356, n46357, n46358, n46359, n46360, n46361, n46362, n46363,
         n46364, n46365, n46366, n46367, n46368, n46369, n46370, n46371,
         n46372, n46373, n46374, n46375, n46376, n46377, n46378, n46379,
         n46380, n46381, n46382, n46383, n46384, n46385, n46386, n46387,
         n46388, n46389, n46390, n46391, n46392, n46393, n46394, n46395,
         n46396, n46397, n46398, n46399, n46400, n46401, n46402, n46403,
         n46404, n46405, n46406, n46407, n46408, n46409, n46410, n46411,
         n46412, n46413, n46414, n46415, n46416, n46417, n46418, n46419,
         n46420, n46421, n46422, n46423, n46424, n46425, n46426, n46427,
         n46428, n46429, n46430, n46431, n46432, n46433, n46434, n46435,
         n46436, n46437, n46438, n46439, n46440, n46441, n46442, n46443,
         n46444, n46445, n46446, n46447, n46448, n46449, n46450, n46451,
         n46452, n46453, n46454, n46455, n46456, n46457, n46458, n46459,
         n46460, n46461, n46462, n46463, n46464, n46465, n46466, n46467,
         n46468, n46469, n46470, n46471, n46472, n46473, n46474, n46475,
         n46476, n46477, n46478, n46479, n46480, n46481, n46482, n46483,
         n46484, n46485, n46486, n46487, n46488, n46489, n46490, n46491,
         n46492, n46493, n46494, n46495, n46496, n46497, n46498, n46499,
         n46500, n46501, n46502, n46503, n46504, n46505, n46506, n46507,
         n46508, n46509, n46510, n46511, n46512, n46513, n46514, n46515,
         n46516, n46517, n46518, n46519, n46520, n46521, n46522, n46523,
         n46524, n46525, n46526, n46527, n46528, n46529, n46530, n46531,
         n46532, n46533, n46534, n46535, n46536, n46537, n46538, n46539,
         n46540, n46541, n46542, n46543, n46544, n46545, n46546, n46547,
         n46548, n46549, n46550, n46551, n46552, n46553, n46554, n46555,
         n46556, n46557, n46558, n46559, n46560, n46561, n46562, n46563,
         n46564, n46565, n46566, n46567, n46568, n46569, n46570, n46571,
         n46572, n46573, n46574, n46575, n46576, n46577, n46578, n46579,
         n46580, n46581, n46582, n46583, n46584, n46585, n46586, n46587,
         n46588, n46589, n46590, n46591, n46592, n46593, n46594, n46595,
         n46596, n46597, n46598, n46599, n46600, n46601, n46602, n46603,
         n46604, n46605, n46606, n46607, n46608, n46609, n46610, n46611,
         n46612, n46613, n46614, n46615, n46616, n46617, n46618, n46619,
         n46620, n46621, n46622, n46623, n46624, n46625, n46626, n46627,
         n46628, n46629, n46630, n46631, n46632, n46633, n46634, n46635,
         n46636, n46637, n46638, n46639, n46640, n46641, n46642, n46643,
         n46644, n46645, n46646, n46647, n46648, n46649, n46650, n46651,
         n46652, n46653, n46654, n46655, n46656, n46657, n46658, n46659,
         n46660, n46661, n46662, n46663, n46664, n46665, n46666, n46667,
         n46668, n46669, n46670, n46671, n46672, n46673, n46674, n46675,
         n46676, n46677, n46678, n46679, n46680, n46681, n46682, n46683,
         n46684, n46685, n46686, n46687, n46688, n46689, n46690, n46691,
         n46692, n46693, n46694, n46695, n46696, n46697, n46698, n46699,
         n46700, n46701, n46702, n46703, n46704, n46705, n46706, n46707,
         n46708, n46709, n46710, n46711, n46712, n46713, n46714, n46715,
         n46716, n46717, n46718, n46719, n46720, n46721, n46722, n46723,
         n46724, n46725, n46726, n46727, n46728, n46729, n46730, n46731,
         n46732, n46733, n46734, n46735, n46736, n46737, n46738, n46739,
         n46740, n46741, n46742, n46743, n46744, n46745, n46746, n46747,
         n46748, n46749, n46750, n46751, n46752, n46753, n46754, n46755,
         n46756, n46757, n46758, n46759, n46760, n46761, n46762, n46763,
         n46764, n46765, n46766, n46767, n46768, n46769, n46770, n46771,
         n46772, n46773, n46774, n46775, n46776, n46777, n46778, n46779,
         n46780, n46781, n46782, n46783, n46784, n46785, n46786, n46787,
         n46788, n46789, n46790, n46791, n46792, n46793, n46794, n46795,
         n46796, n46797, n46798, n46799, n46800, n46801, n46802, n46803,
         n46804, n46805, n46806, n46807, n46808, n46809, n46810, n46811,
         n46812, n46813, n46814, n46815, n46816, n46817, n46818, n46819,
         n46820, n46821, n46822, n46823, n46824, n46825, n46826, n46827,
         n46828, n46829, n46830, n46831, n46832, n46833, n46834, n46835,
         n46836, n46837, n46838, n46839, n46840, n46841, n46842, n46843,
         n46844, n46845, n46846, n46847, n46848, n46849, n46850, n46851,
         n46852, n46853, n46854, n46855, n46856, n46857, n46858, n46859,
         n46860, n46861, n46862, n46863, n46864, n46865, n46866, n46867,
         n46868, n46869, n46870, n46871, n46872, n46873, n46874, n46875,
         n46876, n46877, n46878, n46879, n46880, n46881, n46882, n46883,
         n46884, n46885, n46886, n46887, n46888, n46889, n46890, n46891,
         n46892, n46893, n46894, n46895, n46896, n46897, n46898, n46899,
         n46900, n46901, n46902, n46903, n46904, n46905, n46906, n46907,
         n46908, n46909, n46910, n46911, n46912, n46913, n46914, n46915,
         n46916, n46917, n46918, n46919, n46920, n46921, n46922, n46923,
         n46924, n46925, n46926, n46927, n46928, n46929, n46930, n46931,
         n46932, n46933, n46934, n46935, n46936, n46937, n46938, n46939,
         n46940, n46941, n46942, n46943, n46944, n46945, n46946, n46947,
         n46948, n46949, n46950, n46951, n46952, n46953, n46954, n46955,
         n46956, n46957, n46958, n46959, n46960, n46961, n46962, n46963,
         n46964, n46965, n46966, n46967, n46968, n46969, n46970, n46971,
         n46972, n46973, n46974, n46975, n46976, n46977, n46978, n46979,
         n46980, n46981, n46982, n46983, n46984, n46985, n46986, n46987,
         n46988, n46989, n46990, n46991, n46992, n46993, n46994, n46995,
         n46996, n46997, n46998, n46999, n47000, n47001, n47002, n47003,
         n47004, n47005, n47006, n47007, n47008, n47009, n47010, n47011,
         n47012, n47013, n47014, n47015, n47016, n47017, n47018, n47019,
         n47020, n47021, n47022, n47023, n47024, n47025, n47026, n47027,
         n47028, n47029, n47030, n47031, n47032, n47033, n47034, n47035,
         n47036, n47037, n47038, n47039, n47040, n47041, n47042, n47043,
         n47044, n47045, n47046, n47047, n47048, n47049, n47050, n47051,
         n47052, n47053, n47054, n47055, n47056, n47057, n47058, n47059,
         n47060, n47061, n47062, n47063, n47064, n47065, n47066, n47067,
         n47068, n47069, n47070, n47071, n47072, n47073, n47074, n47075,
         n47076, n47077, n47078, n47079, n47080, n47081, n47082, n47083,
         n47084, n47085, n47086, n47087, n47088, n47089, n47090, n47091,
         n47092, n47093, n47094, n47095, n47096, n47097, n47098, n47099,
         n47100, n47101, n47102, n47103, n47104, n47105, n47106, n47107,
         n47108, n47109, n47110, n47111, n47112, n47113, n47114, n47115,
         n47116, n47117, n47118, n47119, n47120, n47121, n47122, n47123,
         n47124, n47125, n47126, n47127, n47128, n47129, n47130, n47131,
         n47132, n47133, n47134, n47135, n47136, n47137, n47138, n47139,
         n47140, n47141, n47142, n47143, n47144, n47145, n47146, n47147,
         n47148, n47149, n47150, n47151, n47152, n47153, n47154, n47155,
         n47156, n47157, n47158, n47159, n47160, n47161, n47162, n47163,
         n47164, n47165, n47166, n47167, n47168, n47169, n47170, n47171,
         n47172, n47173, n47174, n47175, n47176, n47177, n47178, n47179,
         n47180, n47181, n47182, n47183, n47184, n47185, n47186, n47187,
         n47188, n47189, n47190, n47191, n47192, n47193, n47194, n47195,
         n47196, n47197, n47198, n47199, n47200, n47201, n47202, n47203,
         n47204, n47205, n47206, n47207, n47208, n47209, n47210, n47211,
         n47212, n47213, n47214, n47215, n47216, n47217, n47218, n47219,
         n47220, n47221, n47222, n47223, n47224, n47225, n47226, n47227,
         n47228, n47229, n47230, n47231, n47232, n47233, n47234, n47235,
         n47236, n47237, n47238, n47239, n47240, n47241, n47242, n47243,
         n47244, n47245, n47246, n47247, n47248, n47249, n47250, n47251,
         n47252, n47253, n47254, n47255, n47256, n47257, n47258, n47259,
         n47260, n47261, n47262, n47263, n47264, n47265, n47266, n47267,
         n47268, n47269, n47270, n47271, n47272, n47273, n47274, n47275,
         n47276, n47277, n47278, n47279, n47280, n47281, n47282, n47283,
         n47284, n47285, n47286, n47287, n47288, n47289, n47290, n47291,
         n47292, n47293, n47294, n47295, n47296, n47297, n47298, n47299,
         n47300, n47301, n47302, n47303, n47304, n47305, n47306, n47307,
         n47308, n47309, n47310, n47311, n47312, n47313, n47314, n47315,
         n47316, n47317, n47318, n47319, n47320, n47321, n47322, n47323,
         n47324, n47325, n47326, n47327, n47328, n47329, n47330, n47331,
         n47332, n47333, n47334, n47335, n47336, n47337, n47338, n47339,
         n47340, n47341, n47342, n47343, n47344, n47345, n47346, n47347,
         n47348, n47349, n47350, n47351, n47352, n47353, n47354, n47355,
         n47356, n47357, n47358, n47359, n47360, n47361, n47362, n47363,
         n47364, n47365, n47366, n47367, n47368, n47369, n47370, n47371,
         n47372, n47373, n47374, n47375, n47376, n47377, n47378, n47379,
         n47380, n47381, n47382, n47383, n47384, n47385, n47386, n47387,
         n47388, n47389, n47390, n47391, n47392, n47393, n47394, n47395,
         n47396, n47397, n47398, n47399, n47400, n47401, n47402, n47403,
         n47404, n47405, n47406, n47407, n47408, n47409, n47410, n47411,
         n47412, n47413, n47414, n47415, n47416, n47417, n47418, n47419,
         n47420, n47421, n47422, n47423, n47424, n47425, n47426, n47427,
         n47428, n47429, n47430, n47431, n47432, n47433, n47434, n47435,
         n47436, n47437, n47438, n47439, n47440, n47441, n47442, n47443,
         n47444, n47445, n47446, n47447, n47448, n47449, n47450, n47451,
         n47452, n47453, n47454, n47455, n47456, n47457, n47458, n47459,
         n47460, n47461, n47462, n47463, n47464, n47465, n47466, n47467,
         n47468, n47469, n47470, n47471, n47472, n47473, n47474, n47475,
         n47476, n47477, n47478, n47479, n47480, n47481, n47482, n47483,
         n47484, n47485, n47486, n47487, n47488, n47489, n47490, n47491,
         n47492, n47493, n47494, n47495, n47496, n47497, n47498, n47499,
         n47500, n47501, n47502, n47503, n47504, n47505, n47506, n47507,
         n47508, n47509, n47510, n47511, n47512, n47513, n47514, n47515,
         n47516, n47517, n47518, n47519, n47520, n47521, n47522, n47523,
         n47524, n47525, n47526, n47527, n47528, n47529, n47530, n47531,
         n47532, n47533, n47534, n47535, n47536, n47537, n47538, n47539,
         n47540, n47541, n47542, n47543, n47544, n47545, n47546, n47547,
         n47548, n47549, n47550, n47551, n47552, n47553, n47554, n47555,
         n47556, n47557, n47558, n47559, n47560, n47561, n47562, n47563,
         n47564, n47565, n47566, n47567, n47568, n47569, n47570, n47571,
         n47572, n47573, n47574, n47575, n47576, n47577, n47578, n47579,
         n47580, n47581, n47582, n47583, n47584, n47585, n47586, n47587,
         n47588, n47589, n47590, n47591, n47592, n47593, n47594, n47595,
         n47596, n47597, n47598, n47599, n47600, n47601, n47602, n47603,
         n47604, n47605, n47606, n47607, n47608, n47609, n47610, n47611,
         n47612, n47613, n47614, n47615, n47616, n47617, n47618, n47619,
         n47620, n47621, n47622, n47623, n47624, n47625, n47626, n47627,
         n47628, n47629, n47630, n47631, n47632, n47633, n47634, n47635,
         n47636, n47637, n47638, n47639, n47640, n47641, n47642, n47643,
         n47644, n47645, n47646, n47647, n47648, n47649, n47650, n47651,
         n47652, n47653, n47654, n47655, n47656, n47657, n47658, n47659,
         n47660, n47661, n47662, n47663, n47664, n47665, n47666, n47667,
         n47668, n47669, n47670, n47671, n47672, n47673, n47674, n47675,
         n47676, n47677, n47678, n47679, n47680, n47681, n47682, n47683,
         n47684, n47685, n47686, n47687, n47688, n47689, n47690, n47691,
         n47692, n47693, n47694, n47695, n47696, n47697, n47698, n47699,
         n47700, n47701, n47702, n47703, n47704, n47705, n47706, n47707,
         n47708, n47709, n47710, n47711, n47712, n47713, n47714, n47715,
         n47716, n47717, n47718, n47719, n47720, n47721, n47722, n47723,
         n47724, n47725, n47726, n47727, n47728, n47729, n47730, n47731,
         n47732, n47733, n47734, n47735, n47736, n47737, n47738, n47739,
         n47740, n47741, n47742, n47743, n47744, n47745, n47746, n47747,
         n47748, n47749, n47750, n47751, n47752, n47753, n47754, n47755,
         n47756, n47757, n47758, n47759, n47760, n47761, n47762, n47763,
         n47764, n47765, n47766, n47767, n47768, n47769, n47770, n47771,
         n47772, n47773, n47774, n47775, n47776, n47777, n47778, n47779,
         n47780, n47781, n47782, n47783, n47784, n47785, n47786, n47787,
         n47788, n47789, n47790, n47791, n47792, n47793, n47794, n47795,
         n47796, n47797, n47798, n47799, n47800, n47801, n47802, n47803,
         n47804, n47805, n47806, n47807, n47808, n47809, n47810, n47811,
         n47812, n47813, n47814, n47815, n47816, n47817, n47818, n47819,
         n47820, n47821, n47822, n47823, n47824, n47825, n47826, n47827,
         n47828, n47829, n47830, n47831, n47832, n47833, n47834, n47835,
         n47836, n47837, n47838, n47839, n47840, n47841, n47842, n47843,
         n47844, n47845, n47846, n47847, n47848, n47849, n47850, n47851,
         n47852, n47853, n47854, n47855, n47856, n47857, n47858, n47859,
         n47860, n47861, n47862, n47863, n47864, n47865, n47866, n47867,
         n47868, n47869, n47870, n47871, n47872, n47873, n47874, n47875,
         n47876, n47877, n47878, n47879, n47880, n47881, n47882, n47883,
         n47884, n47885, n47886, n47887, n47888, n47889, n47890, n47891,
         n47892, n47893, n47894, n47895, n47896, n47897, n47898, n47899,
         n47900, n47901, n47902, n47903, n47904, n47905, n47906, n47907,
         n47908, n47909, n47910, n47911, n47912, n47913, n47914, n47915,
         n47916, n47917, n47918, n47919, n47920, n47921, n47922, n47923,
         n47924, n47925, n47926, n47927, n47928, n47929, n47930, n47931,
         n47932, n47933, n47934, n47935, n47936, n47937, n47938, n47939,
         n47940, n47941, n47942, n47943, n47944, n47945, n47946, n47947,
         n47948, n47949, n47950, n47951, n47952, n47953, n47954, n47955,
         n47956, n47957, n47958, n47959, n47960, n47961, n47962, n47963,
         n47964, n47965, n47966, n47967, n47968, n47969, n47970, n47971,
         n47972, n47973, n47974, n47975, n47976, n47977, n47978, n47979,
         n47980, n47981, n47982, n47983, n47984, n47985, n47986, n47987,
         n47988, n47989, n47990, n47991, n47992, n47993, n47994, n47995,
         n47996, n47997, n47998, n47999, n48000, n48001, n48002, n48003,
         n48004, n48005, n48006, n48007, n48008, n48009, n48010, n48011,
         n48012, n48013, n48014, n48015, n48016, n48017, n48018, n48019,
         n48020, n48021, n48022, n48023, n48024, n48025, n48026, n48027,
         n48028, n48029, n48030, n48031, n48032, n48033, n48034, n48035,
         n48036, n48037, n48038, n48039, n48040, n48041, n48042, n48043,
         n48044, n48045, n48046, n48047, n48048, n48049, n48050, n48051,
         n48052, n48053, n48054, n48055, n48056, n48057, n48058, n48059,
         n48060, n48061, n48062, n48063, n48064, n48065, n48066, n48067,
         n48068, n48069, n48070, n48071, n48072, n48073, n48074, n48075,
         n48076, n48077, n48078, n48079, n48080, n48081, n48082, n48083,
         n48084, n48085, n48086, n48087, n48088, n48089, n48090, n48091,
         n48092, n48093, n48094, n48095, n48096, n48097, n48098, n48099,
         n48100, n48101, n48102, n48103, n48104, n48105, n48106, n48107,
         n48108, n48109, n48110, n48111, n48112, n48113, n48114, n48115,
         n48116, n48117, n48118, n48119, n48120, n48121, n48122, n48123,
         n48124, n48125, n48126, n48127, n48128, n48129, n48130, n48131,
         n48132, n48133, n48134, n48135, n48136, n48137, n48138, n48139,
         n48140, n48141, n48142, n48143, n48144, n48145, n48146, n48147,
         n48148, n48149, n48150, n48151, n48152, n48153, n48154, n48155,
         n48156, n48157, n48158, n48159, n48160, n48161, n48162, n48163,
         n48164, n48165, n48166, n48167, n48168, n48169, n48170, n48171,
         n48172, n48173, n48174, n48175, n48176, n48177, n48178, n48179,
         n48180, n48181, n48182, n48183, n48184, n48185, n48186, n48187,
         n48188, n48189, n48190, n48191, n48192, n48193, n48194, n48195,
         n48196, n48197, n48198, n48199, n48200, n48201, n48202, n48203,
         n48204, n48205, n48206, n48207, n48208, n48209, n48210, n48211,
         n48212, n48213, n48214, n48215, n48216, n48217, n48218, n48219,
         n48220, n48221, n48222, n48223, n48224, n48225, n48226, n48227,
         n48228, n48229, n48230, n48231, n48232, n48233, n48234, n48235,
         n48236, n48237, n48238, n48239, n48240, n48241, n48242, n48243,
         n48244, n48245, n48246, n48247, n48248, n48249, n48250, n48251,
         n48252, n48253, n48254, n48255, n48256, n48257, n48258, n48259,
         n48260, n48261, n48262, n48263, n48264, n48265, n48266, n48267,
         n48268, n48269, n48270, n48271, n48272, n48273, n48274, n48275,
         n48276, n48277, n48278, n48279, n48280, n48281, n48282, n48283,
         n48284, n48285, n48286, n48287, n48288, n48289, n48290, n48291,
         n48292, n48293, n48294, n48295, n48296, n48297, n48298, n48299,
         n48300, n48301, n48302, n48303, n48304, n48305, n48306, n48307,
         n48308, n48309, n48310, n48311, n48312, n48313, n48314, n48315,
         n48316, n48317, n48318, n48319, n48320, n48321, n48322, n48323,
         n48324, n48325, n48326, n48327, n48328, n48329, n48330, n48331,
         n48332, n48333, n48334, n48335, n48336, n48337, n48338, n48339,
         n48340, n48341, n48342, n48343, n48344, n48345, n48346, n48347,
         n48348, n48349, n48350, n48351, n48352, n48353, n48354, n48355,
         n48356, n48357, n48358, n48359, n48360, n48361, n48362, n48363,
         n48364, n48365, n48366, n48367, n48368, n48369, n48370, n48371,
         n48372, n48373, n48374, n48375, n48376, n48377, n48378, n48379,
         n48380, n48381, n48382, n48383, n48384, n48385, n48386, n48387,
         n48388, n48389, n48390, n48391, n48392, n48393, n48394, n48395,
         n48396, n48397, n48398, n48399, n48400, n48401, n48402, n48403,
         n48404, n48405, n48406, n48407, n48408, n48409, n48410, n48411,
         n48412, n48413, n48414, n48415, n48416, n48417, n48418, n48419,
         n48420, n48421, n48422, n48423, n48424, n48425, n48426, n48427,
         n48428, n48429, n48430, n48431, n48432, n48433, n48434, n48435,
         n48436, n48437, n48438, n48439, n48440, n48441, n48442, n48443,
         n48444, n48445, n48446, n48447, n48448, n48449, n48450, n48451,
         n48452, n48453, n48454, n48455, n48456, n48457, n48458, n48459,
         n48460, n48461, n48462, n48463, n48464, n48465, n48466, n48467,
         n48468, n48469, n48470, n48471, n48472, n48473, n48474, n48475,
         n48476, n48477, n48478, n48479, n48480, n48481, n48482, n48483,
         n48484, n48485, n48486, n48487, n48488, n48489, n48490, n48491,
         n48492, n48493, n48494, n48495, n48496, n48497, n48498, n48499,
         n48500, n48501, n48502, n48503, n48504, n48505, n48506, n48507,
         n48508, n48509, n48510, n48511, n48512, n48513, n48514, n48515,
         n48516, n48517, n48518, n48519, n48520, n48521, n48522, n48523,
         n48524, n48525, n48526, n48527, n48528, n48529, n48530, n48531,
         n48532, n48533, n48534, n48535, n48536, n48537, n48538, n48539,
         n48540, n48541, n48542, n48543, n48544, n48545, n48546, n48547,
         n48548, n48549, n48550, n48551, n48552, n48553, n48554, n48555,
         n48556, n48557, n48558, n48559, n48560, n48561, n48562, n48563,
         n48564, n48565, n48566, n48567, n48568, n48569, n48570, n48571,
         n48572, n48573, n48574, n48575, n48576, n48577, n48578, n48579,
         n48580, n48581, n48582, n48583, n48584, n48585, n48586, n48587,
         n48588, n48589, n48590, n48591, n48592, n48593, n48594, n48595,
         n48596, n48597, n48598, n48599, n48600, n48601, n48602, n48603,
         n48604, n48605, n48606, n48607, n48608, n48609, n48610, n48611,
         n48612, n48613, n48614, n48615, n48616, n48617, n48618, n48619,
         n48620, n48621, n48622, n48623, n48624, n48625, n48626, n48627,
         n48628, n48629, n48630, n48631, n48632, n48633, n48634, n48635,
         n48636, n48637, n48638, n48639, n48640, n48641, n48642, n48643,
         n48644, n48645, n48646, n48647, n48648, n48649, n48650, n48651,
         n48652, n48653, n48654, n48655, n48656, n48657, n48658, n48659,
         n48660, n48661, n48662, n48663, n48664, n48665, n48666, n48667,
         n48668, n48669, n48670, n48671, n48672, n48673, n48674, n48675,
         n48676, n48677, n48678, n48679, n48680, n48681, n48682, n48683,
         n48684, n48685, n48686, n48687, n48688, n48689, n48690, n48691,
         n48692, n48693, n48694, n48695, n48696, n48697, n48698, n48699,
         n48700, n48701, n48702, n48703, n48704, n48705, n48706, n48707,
         n48708, n48709, n48710, n48711, n48712, n48713, n48714, n48715,
         n48716, n48717, n48718, n48719, n48720, n48721, n48722, n48723,
         n48724, n48725, n48726, n48727, n48728, n48729, n48730, n48731,
         n48732, n48733, n48734, n48735, n48736, n48737, n48738, n48739,
         n48740, n48741, n48742, n48743, n48744, n48745, n48746, n48747,
         n48748, n48749, n48750, n48751, n48752, n48753, n48754, n48755,
         n48756, n48757, n48758, n48759, n48760, n48761, n48762, n48763,
         n48764, n48765, n48766, n48767, n48768, n48769, n48770, n48771,
         n48772, n48773, n48774, n48775, n48776, n48777, n48778, n48779,
         n48780, n48781, n48782, n48783, n48784, n48785, n48786, n48787,
         n48788, n48789, n48790, n48791, n48792, n48793, n48794, n48795,
         n48796, n48797, n48798, n48799, n48800, n48801, n48802, n48803,
         n48804, n48805, n48806, n48807, n48808, n48809, n48810, n48811,
         n48812, n48813, n48814, n48815, n48816, n48817, n48818, n48819,
         n48820, n48821, n48822, n48823, n48824, n48825, n48826, n48827,
         n48828, n48829, n48830, n48831, n48832, n48833, n48834, n48835,
         n48836, n48837, n48838, n48839, n48840, n48841, n48842, n48843,
         n48844, n48845, n48846, n48847, n48848, n48849, n48850, n48851,
         n48852, n48853, n48854, n48855, n48856, n48857, n48858, n48859,
         n48860, n48861, n48862, n48863, n48864, n48865, n48866, n48867,
         n48868, n48869, n48870, n48871, n48872, n48873, n48874, n48875,
         n48876, n48877, n48878, n48879, n48880, n48881, n48882, n48883,
         n48884, n48885, n48886, n48887, n48888, n48889, n48890, n48891,
         n48892, n48893, n48894, n48895, n48896, n48897, n48898, n48899,
         n48900, n48901, n48902, n48903, n48904, n48905, n48906, n48907,
         n48908, n48909, n48910, n48911, n48912, n48913, n48914, n48915,
         n48916, n48917, n48918, n48919, n48920, n48921, n48922, n48923,
         n48924, n48925, n48926, n48927, n48928, n48929, n48930, n48931,
         n48932, n48933, n48934, n48935, n48936, n48937, n48938, n48939,
         n48940, n48941, n48942, n48943, n48944, n48945, n48946, n48947,
         n48948, n48949, n48950, n48951, n48952, n48953, n48954, n48955,
         n48956, n48957, n48958, n48959, n48960, n48961, n48962, n48963,
         n48964, n48965, n48966, n48967, n48968, n48969, n48970, n48971,
         n48972, n48973, n48974, n48975, n48976, n48977, n48978, n48979,
         n48980, n48981, n48982, n48983, n48984, n48985, n48986, n48987,
         n48988, n48989, n48990, n48991, n48992, n48993, n48994, n48995,
         n48996, n48997, n48998, n48999, n49000, n49001, n49002, n49003,
         n49004, n49005, n49006, n49007, n49008, n49009, n49010, n49011,
         n49012, n49013, n49014, n49015, n49016, n49017, n49018, n49019,
         n49020, n49021, n49022, n49023, n49024, n49025, n49026, n49027,
         n49028, n49029, n49030, n49031, n49032, n49033, n49034, n49035,
         n49036, n49037, n49038, n49039, n49040, n49041, n49042, n49043,
         n49044, n49045, n49046, n49047, n49048, n49049, n49050, n49051,
         n49052, n49053, n49054, n49055, n49056, n49057, n49058, n49059,
         n49060, n49061, n49062, n49063, n49064, n49065, n49066, n49067,
         n49068, n49069, n49070, n49071, n49072, n49073, n49074, n49075,
         n49076, n49077, n49078, n49079, n49080, n49081, n49082, n49083,
         n49084, n49085, n49086, n49087, n49088, n49089, n49090, n49091,
         n49092, n49093, n49094, n49095, n49096, n49097, n49098, n49099,
         n49100, n49101, n49102, n49103, n49104, n49105, n49106, n49107,
         n49108, n49109, n49110, n49111, n49112, n49113, n49114, n49115,
         n49116, n49117, n49118, n49119, n49120, n49121, n49122, n49123,
         n49124, n49125, n49126, n49127, n49128, n49129, n49130, n49131,
         n49132, n49133, n49134, n49135, n49136, n49137, n49138, n49139,
         n49140, n49141, n49142, n49143, n49144, n49145, n49146, n49147,
         n49148, n49149, n49150, n49151, n49152, n49153, n49154, n49155,
         n49156, n49157, n49158, n49159, n49160, n49161, n49162, n49163,
         n49164, n49165, n49166, n49167, n49168, n49169, n49170, n49171,
         n49172, n49173, n49174, n49175, n49176, n49177, n49178, n49179,
         n49180, n49181, n49182, n49183, n49184, n49185, n49186, n49187,
         n49188, n49189, n49190, n49191, n49192, n49193, n49194, n49195,
         n49196, n49197, n49198, n49199, n49200, n49201, n49202, n49203,
         n49204, n49205, n49206, n49207, n49208, n49209, n49210, n49211,
         n49212, n49213, n49214, n49215, n49216, n49217, n49218, n49219,
         n49220, n49221, n49222, n49223, n49224, n49225, n49226, n49227,
         n49228, n49229, n49230, n49231, n49232, n49233, n49234, n49235,
         n49236, n49237, n49238, n49239, n49240, n49241, n49242, n49243,
         n49244, n49245, n49246, n49247, n49248, n49249, n49250, n49251,
         n49252, n49253, n49254, n49255, n49256, n49257, n49258, n49259,
         n49260, n49261, n49262, n49263, n49264, n49265, n49266, n49267,
         n49268, n49269, n49270, n49271, n49272, n49273, n49274, n49275,
         n49276, n49277, n49278, n49279, n49280, n49281, n49282, n49283,
         n49284, n49285, n49286, n49287, n49288, n49289, n49290, n49291,
         n49292, n49293, n49294, n49295, n49296, n49297, n49298, n49299,
         n49300, n49301, n49302, n49303, n49304, n49305, n49306, n49307,
         n49308, n49309, n49310, n49311, n49312, n49313, n49314, n49315,
         n49316, n49317, n49318, n49319, n49320, n49321, n49322, n49323,
         n49324, n49325, n49326, n49327, n49328, n49329, n49330, n49331,
         n49332, n49333, n49334, n49335, n49336, n49337, n49338, n49339,
         n49340, n49341, n49342, n49343, n49344, n49345, n49346, n49347,
         n49348, n49349, n49350, n49351, n49352, n49353, n49354, n49355,
         n49356, n49357, n49358, n49359, n49360, n49361, n49362, n49363,
         n49364, n49365, n49366, n49367, n49368, n49369, n49370, n49371,
         n49372, n49373, n49374, n49375, n49376, n49377, n49378, n49379,
         n49380, n49381, n49382, n49383, n49384, n49385, n49386, n49387,
         n49388, n49389, n49390, n49391, n49392, n49393, n49394, n49395,
         n49396, n49397, n49398, n49399, n49400, n49401, n49402, n49403,
         n49404, n49405, n49406, n49407, n49408, n49409, n49410, n49411,
         n49412, n49413, n49414, n49415, n49416, n49417, n49418, n49419,
         n49420, n49421, n49422, n49423, n49424, n49425, n49426, n49427,
         n49428, n49429, n49430, n49431, n49432, n49433, n49434, n49435,
         n49436, n49437, n49438, n49439, n49440, n49441, n49442, n49443,
         n49444, n49445, n49446, n49447, n49448, n49449, n49450, n49451,
         n49452, n49453, n49454, n49455, n49456, n49457, n49458, n49459,
         n49460, n49461, n49462, n49463, n49464, n49465, n49466, n49467,
         n49468, n49469, n49470, n49471, n49472, n49473, n49474, n49475,
         n49476, n49477, n49478, n49479, n49480, n49481, n49482, n49483,
         n49484, n49485, n49486, n49487, n49488, n49489, n49490, n49491,
         n49492, n49493, n49494, n49495, n49496, n49497, n49498, n49499,
         n49500, n49501, n49502, n49503, n49504, n49505, n49506, n49507,
         n49508, n49509, n49510, n49511, n49512, n49513, n49514, n49515,
         n49516, n49517, n49518, n49519, n49520, n49521, n49522, n49523,
         n49524, n49525, n49526, n49527, n49528, n49529, n49530, n49531,
         n49532, n49533, n49534, n49535, n49536, n49537, n49538, n49539,
         n49540, n49541, n49542, n49543, n49544, n49545, n49546, n49547,
         n49548, n49549, n49550, n49551, n49552, n49553, n49554, n49555,
         n49556, n49557, n49558, n49559, n49560, n49561, n49562, n49563,
         n49564, n49565, n49566, n49567, n49568, n49569, n49570, n49571,
         n49572, n49573, n49574, n49575, n49576, n49577, n49578, n49579,
         n49580, n49581, n49582, n49583, n49584, n49585, n49586, n49587,
         n49588, n49589, n49590, n49591, n49592, n49593, n49594, n49595,
         n49596, n49597, n49598, n49599, n49600, n49601, n49602, n49603,
         n49604, n49605, n49606, n49607, n49608, n49609, n49610, n49611,
         n49612, n49613, n49614, n49615, n49616, n49617, n49618, n49619,
         n49620, n49621, n49622, n49623, n49624, n49625, n49626, n49627,
         n49628, n49629, n49630, n49631, n49632, n49633, n49634, n49635,
         n49636, n49637, n49638, n49639, n49640, n49641, n49642, n49643,
         n49644, n49645, n49646, n49647, n49648, n49649, n49650, n49651,
         n49652, n49653, n49654, n49655, n49656, n49657, n49658, n49659,
         n49660, n49661, n49662, n49663, n49664, n49665, n49666, n49667,
         n49668, n49669, n49670, n49671, n49672, n49673, n49674, n49675,
         n49676, n49677, n49678, n49679, n49680, n49681, n49682, n49683,
         n49684, n49685, n49686, n49687, n49688, n49689, n49690, n49691,
         n49692, n49693, n49694, n49695, n49696, n49697, n49698, n49699,
         n49700, n49701, n49702, n49703, n49704, n49705, n49706, n49707,
         n49708, n49709, n49710, n49711, n49712, n49713, n49714, n49715,
         n49716, n49717, n49718, n49719, n49720, n49721, n49722, n49723,
         n49724, n49725, n49726, n49727, n49728, n49729, n49730, n49731,
         n49732, n49733, n49734, n49735, n49736, n49737, n49738, n49739,
         n49740, n49741, n49742, n49743, n49744, n49745, n49746, n49747,
         n49748, n49749, n49750, n49751, n49752, n49753, n49754, n49755,
         n49756, n49757, n49758, n49759, n49760, n49761, n49762, n49763,
         n49764, n49765, n49766, n49767, n49768, n49769, n49770, n49771,
         n49772, n49773, n49774, n49775, n49776, n49777, n49778, n49779,
         n49780, n49781, n49782, n49783, n49784, n49785, n49786, n49787,
         n49788, n49789, n49790, n49791, n49792, n49793, n49794, n49795,
         n49796, n49797, n49798, n49799, n49800, n49801, n49802, n49803,
         n49804, n49805, n49806, n49807, n49808, n49809, n49810, n49811,
         n49812, n49813, n49814, n49815, n49816, n49817, n49818, n49819,
         n49820, n49821, n49822, n49823, n49824, n49825, n49826, n49827,
         n49828, n49829, n49830, n49831, n49832, n49833, n49834, n49835,
         n49836, n49837, n49838, n49839, n49840, n49841, n49842, n49843,
         n49844, n49845, n49846, n49847, n49848, n49849, n49850, n49851,
         n49852, n49853, n49854, n49855, n49856, n49857, n49858, n49859,
         n49860, n49861, n49862, n49863, n49864, n49865, n49866, n49867,
         n49868, n49869, n49870, n49871, n49872, n49873, n49874, n49875,
         n49876, n49877, n49878, n49879, n49880, n49881, n49882, n49883,
         n49884, n49885, n49886, n49887, n49888, n49889, n49890, n49891,
         n49892, n49893, n49894, n49895, n49896, n49897, n49898, n49899,
         n49900, n49901, n49902, n49903, n49904, n49905, n49906, n49907,
         n49908, n49909, n49910, n49911, n49912, n49913, n49914, n49915,
         n49916, n49917, n49918, n49919, n49920, n49921, n49922, n49923,
         n49924, n49925, n49926, n49927, n49928, n49929, n49930, n49931,
         n49932, n49933, n49934, n49935, n49936, n49937, n49938, n49939,
         n49940, n49941, n49942, n49943, n49944, n49945, n49946, n49947,
         n49948, n49949, n49950, n49951, n49952, n49953, n49954, n49955,
         n49956, n49957, n49958, n49959, n49960, n49961, n49962, n49963,
         n49964, n49965, n49966, n49967, n49968, n49969, n49970, n49971,
         n49972, n49973, n49974, n49975, n49976, n49977, n49978, n49979,
         n49980, n49981, n49982, n49983, n49984, n49985, n49986, n49987,
         n49988, n49989, n49990, n49991, n49992, n49993, n49994, n49995,
         n49996, n49997, n49998, n49999, n50000, n50001, n50002, n50003,
         n50004, n50005, n50006, n50007, n50008, n50009, n50010, n50011,
         n50012, n50013, n50014, n50015, n50016, n50017, n50018, n50019,
         n50020, n50021, n50022, n50023, n50024, n50025, n50026, n50027,
         n50028, n50029, n50030, n50031, n50032, n50033, n50034, n50035,
         n50036, n50037, n50038, n50039, n50040, n50041, n50042, n50043,
         n50044, n50045, n50046, n50047, n50048, n50049, n50050, n50051,
         n50052, n50053, n50054, n50055, n50056, n50057, n50058, n50059,
         n50060, n50061, n50062, n50063, n50064, n50065, n50066, n50067,
         n50068, n50069, n50070, n50071, n50072, n50073, n50074, n50075,
         n50076, n50077, n50078, n50079, n50080, n50081, n50082, n50083,
         n50084, n50085, n50086, n50087, n50088, n50089, n50090, n50091,
         n50092, n50093, n50094, n50095, n50096, n50097, n50098, n50099,
         n50100, n50101, n50102, n50103, n50104, n50105, n50106, n50107,
         n50108, n50109, n50110, n50111, n50112, n50113, n50114, n50115,
         n50116, n50117, n50118, n50119, n50120, n50121, n50122, n50123,
         n50124, n50125, n50126, n50127, n50128, n50129, n50130, n50131,
         n50132, n50133, n50134, n50135, n50136, n50137, n50138, n50139,
         n50140, n50141, n50142, n50143, n50144, n50145, n50146, n50147,
         n50148, n50149, n50150, n50151, n50152, n50153, n50154, n50155,
         n50156, n50157, n50158, n50159, n50160, n50161, n50162, n50163,
         n50164, n50165, n50166, n50167, n50168, n50169, n50170, n50171,
         n50172, n50173, n50174, n50175, n50176, n50177, n50178, n50179,
         n50180, n50181, n50182, n50183, n50184, n50185, n50186, n50187,
         n50188, n50189, n50190, n50191, n50192, n50193, n50194, n50195,
         n50196, n50197, n50198, n50199, n50200, n50201, n50202, n50203,
         n50204, n50205, n50206, n50207, n50208, n50209, n50210, n50211,
         n50212, n50213, n50214, n50215, n50216, n50217, n50218, n50219,
         n50220, n50221, n50222, n50223, n50224, n50225, n50226, n50227,
         n50228, n50229, n50230, n50231, n50232, n50233, n50234, n50235,
         n50236, n50237, n50238, n50239, n50240, n50241, n50242, n50243,
         n50244, n50245, n50246, n50247, n50248, n50249, n50250, n50251,
         n50252, n50253, n50254, n50255, n50256, n50257, n50258, n50259,
         n50260, n50261, n50262, n50263, n50264, n50265, n50266, n50267,
         n50268, n50269, n50270, n50271, n50272, n50273, n50274, n50275,
         n50276, n50277, n50278, n50279, n50280, n50281, n50282, n50283,
         n50284, n50285, n50286, n50287, n50288, n50289, n50290, n50291,
         n50292, n50293, n50294, n50295, n50296, n50297, n50298, n50299,
         n50300, n50301, n50302, n50303, n50304, n50305, n50306, n50307,
         n50308, n50309, n50310, n50311, n50312, n50313, n50314, n50315,
         n50316, n50317, n50318, n50319, n50320, n50321, n50322, n50323,
         n50324, n50325, n50326, n50327, n50328, n50329, n50330, n50331,
         n50332, n50333, n50334, n50335, n50336, n50337, n50338, n50339,
         n50340, n50341, n50342, n50343, n50344, n50345, n50346, n50347,
         n50348, n50349, n50350, n50351, n50352, n50353, n50354, n50355,
         n50356, n50357, n50358, n50359, n50360, n50361, n50362, n50363,
         n50364, n50365, n50366, n50367, n50368, n50369, n50370, n50371,
         n50372, n50373, n50374, n50375, n50376, n50377, n50378, n50379,
         n50380, n50381, n50382, n50383, n50384, n50385, n50386, n50387,
         n50388, n50389, n50390, n50391, n50392, n50393, n50394, n50395,
         n50396, n50397, n50398, n50399, n50400, n50401, n50402, n50403,
         n50404, n50405, n50406, n50407, n50408, n50409, n50410, n50411,
         n50412, n50413, n50414, n50415, n50416, n50417, n50418, n50419,
         n50420, n50421, n50422, n50423, n50424, n50425, n50426, n50427,
         n50428, n50429, n50430, n50431, n50432, n50433, n50434, n50435,
         n50436, n50437, n50438, n50439, n50440, n50441, n50442, n50443,
         n50444, n50445, n50446, n50447, n50448, n50449, n50450, n50451,
         n50452, n50453, n50454, n50455, n50456, n50457, n50458, n50459,
         n50460, n50461, n50462, n50463, n50464, n50465, n50466, n50467,
         n50468, n50469, n50470, n50471, n50472, n50473, n50474, n50475,
         n50476, n50477, n50478, n50479, n50480, n50481, n50482, n50483,
         n50484, n50485, n50486, n50487, n50488, n50489, n50490, n50491,
         n50492, n50493, n50494, n50495, n50496, n50497, n50498, n50499,
         n50500, n50501, n50502, n50503, n50504, n50505, n50506, n50507,
         n50508, n50509, n50510, n50511, n50512, n50513, n50514, n50515,
         n50516, n50517, n50518, n50519, n50520, n50521, n50522, n50523,
         n50524, n50525, n50526, n50527, n50528, n50529, n50530, n50531,
         n50532, n50533, n50534, n50535, n50536, n50537, n50538, n50539,
         n50540, n50541, n50542, n50543, n50544, n50545, n50546, n50547,
         n50548, n50549, n50550, n50551, n50552, n50553, n50554, n50555,
         n50556, n50557, n50558, n50559, n50560, n50561, n50562, n50563,
         n50564, n50565, n50566, n50567, n50568, n50569, n50570, n50571,
         n50572, n50573, n50574, n50575, n50576, n50577, n50578, n50579,
         n50580, n50581, n50582, n50583, n50584, n50585, n50586, n50587,
         n50588, n50589, n50590, n50591, n50592, n50593, n50594, n50595,
         n50596, n50597, n50598, n50599, n50600, n50601, n50602, n50603,
         n50604, n50605, n50606, n50607, n50608, n50609, n50610, n50611,
         n50612, n50613, n50614, n50615, n50616, n50617, n50618, n50619,
         n50620, n50621, n50622, n50623, n50624, n50625, n50626, n50627,
         n50628, n50629, n50630, n50631, n50632, n50633, n50634, n50635,
         n50636, n50637, n50638, n50639, n50640, n50641, n50642, n50643,
         n50644, n50645, n50646, n50647, n50648, n50649, n50650, n50651,
         n50652, n50653, n50654, n50655, n50656, n50657, n50658, n50659,
         n50660, n50661, n50662, n50663, n50664, n50665, n50666, n50667,
         n50668, n50669, n50670, n50671, n50672, n50673, n50674, n50675,
         n50676, n50677, n50678, n50679, n50680, n50681, n50682, n50683,
         n50684, n50685, n50686, n50687, n50688, n50689, n50690, n50691,
         n50692, n50693, n50694, n50695, n50696, n50697, n50698, n50699,
         n50700, n50701, n50702, n50703, n50704, n50705, n50706, n50707,
         n50708, n50709, n50710, n50711, n50712, n50713, n50714, n50715,
         n50716, n50717, n50718, n50719, n50720, n50721, n50722, n50723,
         n50724, n50725, n50726, n50727, n50728, n50729, n50730, n50731,
         n50732, n50733;
  assign \knn_comb_/min_val_out[0][0]  = p_input[2016];
  assign \knn_comb_/min_val_out[0][1]  = p_input[2017];
  assign \knn_comb_/min_val_out[0][2]  = p_input[2018];
  assign \knn_comb_/min_val_out[0][3]  = p_input[2019];
  assign \knn_comb_/min_val_out[0][4]  = p_input[2020];
  assign \knn_comb_/min_val_out[0][5]  = p_input[2021];
  assign \knn_comb_/min_val_out[0][6]  = p_input[2022];
  assign \knn_comb_/min_val_out[0][7]  = p_input[2023];
  assign \knn_comb_/min_val_out[0][8]  = p_input[2024];
  assign \knn_comb_/min_val_out[0][9]  = p_input[2025];
  assign \knn_comb_/min_val_out[0][10]  = p_input[2026];
  assign \knn_comb_/min_val_out[0][11]  = p_input[2027];
  assign \knn_comb_/min_val_out[0][12]  = p_input[2028];
  assign \knn_comb_/min_val_out[0][13]  = p_input[2029];
  assign \knn_comb_/min_val_out[0][14]  = p_input[2030];
  assign \knn_comb_/min_val_out[0][15]  = p_input[2031];
  assign \knn_comb_/min_val_out[0][16]  = p_input[2032];
  assign \knn_comb_/min_val_out[0][17]  = p_input[2033];
  assign \knn_comb_/min_val_out[0][18]  = p_input[2034];
  assign \knn_comb_/min_val_out[0][19]  = p_input[2035];
  assign \knn_comb_/min_val_out[0][20]  = p_input[2036];
  assign \knn_comb_/min_val_out[0][21]  = p_input[2037];
  assign \knn_comb_/min_val_out[0][22]  = p_input[2038];
  assign \knn_comb_/min_val_out[0][23]  = p_input[2039];
  assign \knn_comb_/min_val_out[0][24]  = p_input[2040];
  assign \knn_comb_/min_val_out[0][25]  = p_input[2041];
  assign \knn_comb_/min_val_out[0][26]  = p_input[2042];
  assign \knn_comb_/min_val_out[0][27]  = p_input[2043];
  assign \knn_comb_/min_val_out[0][28]  = p_input[2044];
  assign \knn_comb_/min_val_out[0][29]  = p_input[2045];
  assign \knn_comb_/min_val_out[0][30]  = p_input[2046];
  assign \knn_comb_/min_val_out[0][31]  = p_input[2047];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][0]  = p_input[1952];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][1]  = p_input[1953];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][2]  = p_input[1954];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][3]  = p_input[1955];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][4]  = p_input[1956];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][5]  = p_input[1957];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][6]  = p_input[1958];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][7]  = p_input[1959];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][8]  = p_input[1960];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][9]  = p_input[1961];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][10]  = p_input[1962];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][11]  = p_input[1963];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][12]  = p_input[1964];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][13]  = p_input[1965];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][14]  = p_input[1966];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][15]  = p_input[1967];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][16]  = p_input[1968];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][17]  = p_input[1969];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][18]  = p_input[1970];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][19]  = p_input[1971];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][20]  = p_input[1972];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][21]  = p_input[1973];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][22]  = p_input[1974];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][23]  = p_input[1975];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][24]  = p_input[1976];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][25]  = p_input[1977];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][26]  = p_input[1978];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][27]  = p_input[1979];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][28]  = p_input[1980];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][29]  = p_input[1981];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][30]  = p_input[1982];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][31]  = p_input[1983];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][0]  = p_input[1984];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][1]  = p_input[1985];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][2]  = p_input[1986];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][3]  = p_input[1987];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][4]  = p_input[1988];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][5]  = p_input[1989];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][6]  = p_input[1990];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][7]  = p_input[1991];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][8]  = p_input[1992];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][9]  = p_input[1993];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][10]  = p_input[1994];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][11]  = p_input[1995];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][12]  = p_input[1996];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][13]  = p_input[1997];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][14]  = p_input[1998];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][15]  = p_input[1999];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][16]  = p_input[2000];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][17]  = p_input[2001];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][18]  = p_input[2002];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][19]  = p_input[2003];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][20]  = p_input[2004];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][21]  = p_input[2005];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][22]  = p_input[2006];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][23]  = p_input[2007];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][24]  = p_input[2008];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][25]  = p_input[2009];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][26]  = p_input[2010];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][27]  = p_input[2011];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][28]  = p_input[2012];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][29]  = p_input[2013];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][30]  = p_input[2014];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][31]  = p_input[2015];

  XOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  XOR U2 ( .A(n3), .B(n4), .Z(o[95]) );
  XOR U3 ( .A(n5), .B(n6), .Z(o[94]) );
  XOR U4 ( .A(n7), .B(n8), .Z(o[93]) );
  XOR U5 ( .A(n9), .B(n10), .Z(o[92]) );
  XOR U6 ( .A(n11), .B(n12), .Z(o[91]) );
  XOR U7 ( .A(n13), .B(n14), .Z(o[90]) );
  XOR U8 ( .A(n15), .B(n16), .Z(o[8]) );
  XOR U9 ( .A(n17), .B(n18), .Z(o[89]) );
  XOR U10 ( .A(n19), .B(n20), .Z(o[88]) );
  XOR U11 ( .A(n21), .B(n22), .Z(o[87]) );
  XOR U12 ( .A(n23), .B(n24), .Z(o[86]) );
  XOR U13 ( .A(n25), .B(n26), .Z(o[85]) );
  XOR U14 ( .A(n27), .B(n28), .Z(o[84]) );
  XOR U15 ( .A(n29), .B(n30), .Z(o[83]) );
  XOR U16 ( .A(n31), .B(n32), .Z(o[82]) );
  XOR U17 ( .A(n33), .B(n34), .Z(o[81]) );
  XOR U18 ( .A(n35), .B(n36), .Z(o[80]) );
  XOR U19 ( .A(n37), .B(n38), .Z(o[7]) );
  XOR U20 ( .A(n39), .B(n40), .Z(o[79]) );
  XOR U21 ( .A(n41), .B(n42), .Z(o[78]) );
  XOR U22 ( .A(n43), .B(n44), .Z(o[77]) );
  XOR U23 ( .A(n45), .B(n46), .Z(o[76]) );
  XOR U24 ( .A(n47), .B(n48), .Z(o[75]) );
  XOR U25 ( .A(n49), .B(n50), .Z(o[74]) );
  XOR U26 ( .A(n51), .B(n52), .Z(o[73]) );
  XOR U27 ( .A(n53), .B(n54), .Z(o[72]) );
  XOR U28 ( .A(n55), .B(n56), .Z(o[71]) );
  XOR U29 ( .A(n57), .B(n58), .Z(o[70]) );
  XOR U30 ( .A(n59), .B(n60), .Z(o[6]) );
  XOR U31 ( .A(n61), .B(n62), .Z(o[69]) );
  XOR U32 ( .A(n63), .B(n64), .Z(o[68]) );
  XOR U33 ( .A(n65), .B(n66), .Z(o[67]) );
  XOR U34 ( .A(n67), .B(n68), .Z(o[66]) );
  XOR U35 ( .A(n69), .B(n70), .Z(o[65]) );
  XOR U36 ( .A(n71), .B(n72), .Z(o[64]) );
  XOR U37 ( .A(n73), .B(n74), .Z(o[63]) );
  XOR U38 ( .A(n75), .B(n76), .Z(o[62]) );
  XOR U39 ( .A(n77), .B(n78), .Z(o[61]) );
  XOR U40 ( .A(n79), .B(n80), .Z(o[60]) );
  XOR U41 ( .A(n81), .B(n82), .Z(o[5]) );
  XOR U42 ( .A(n83), .B(n84), .Z(o[59]) );
  XOR U43 ( .A(n85), .B(n86), .Z(o[58]) );
  XOR U44 ( .A(n87), .B(n88), .Z(o[57]) );
  XOR U45 ( .A(n89), .B(n90), .Z(o[56]) );
  XOR U46 ( .A(n91), .B(n92), .Z(o[55]) );
  XOR U47 ( .A(n93), .B(n94), .Z(o[54]) );
  XOR U48 ( .A(n95), .B(n96), .Z(o[53]) );
  XOR U49 ( .A(n97), .B(n98), .Z(o[52]) );
  XOR U50 ( .A(n99), .B(n100), .Z(o[51]) );
  XOR U51 ( .A(n101), .B(n102), .Z(o[50]) );
  XOR U52 ( .A(n103), .B(n104), .Z(o[4]) );
  XOR U53 ( .A(n105), .B(n106), .Z(o[49]) );
  XOR U54 ( .A(n107), .B(n108), .Z(o[48]) );
  XOR U55 ( .A(n109), .B(n110), .Z(o[47]) );
  XOR U56 ( .A(n111), .B(n112), .Z(o[46]) );
  XOR U57 ( .A(n113), .B(n114), .Z(o[45]) );
  XOR U58 ( .A(n115), .B(n116), .Z(o[44]) );
  XOR U59 ( .A(n117), .B(n118), .Z(o[43]) );
  XOR U60 ( .A(n119), .B(n120), .Z(o[42]) );
  XOR U61 ( .A(n1), .B(n121), .Z(o[41]) );
  AND U62 ( .A(n122), .B(n123), .Z(n1) );
  XOR U63 ( .A(n2), .B(n121), .Z(n123) );
  XOR U64 ( .A(n124), .B(n51), .Z(n121) );
  AND U65 ( .A(n125), .B(n126), .Z(n51) );
  XNOR U66 ( .A(n127), .B(n52), .Z(n126) );
  XOR U67 ( .A(n128), .B(n129), .Z(n52) );
  AND U68 ( .A(n130), .B(n131), .Z(n129) );
  XOR U69 ( .A(p_input[9]), .B(n128), .Z(n131) );
  XOR U70 ( .A(n132), .B(n133), .Z(n128) );
  AND U71 ( .A(n134), .B(n135), .Z(n133) );
  IV U72 ( .A(n124), .Z(n127) );
  XOR U73 ( .A(n136), .B(n137), .Z(n124) );
  AND U74 ( .A(n138), .B(n139), .Z(n137) );
  XOR U75 ( .A(n140), .B(n141), .Z(n2) );
  AND U76 ( .A(n142), .B(n139), .Z(n141) );
  XNOR U77 ( .A(n143), .B(n136), .Z(n139) );
  XOR U78 ( .A(n144), .B(n145), .Z(n136) );
  AND U79 ( .A(n146), .B(n135), .Z(n145) );
  XNOR U80 ( .A(n147), .B(n132), .Z(n135) );
  XOR U81 ( .A(n148), .B(n149), .Z(n132) );
  AND U82 ( .A(n150), .B(n151), .Z(n149) );
  XOR U83 ( .A(p_input[41]), .B(n148), .Z(n151) );
  XOR U84 ( .A(n152), .B(n153), .Z(n148) );
  AND U85 ( .A(n154), .B(n155), .Z(n153) );
  IV U86 ( .A(n144), .Z(n147) );
  XOR U87 ( .A(n156), .B(n157), .Z(n144) );
  AND U88 ( .A(n158), .B(n159), .Z(n157) );
  IV U89 ( .A(n140), .Z(n143) );
  XNOR U90 ( .A(n160), .B(n161), .Z(n140) );
  AND U91 ( .A(n162), .B(n159), .Z(n161) );
  XNOR U92 ( .A(n160), .B(n156), .Z(n159) );
  XOR U93 ( .A(n163), .B(n164), .Z(n156) );
  AND U94 ( .A(n165), .B(n155), .Z(n164) );
  XNOR U95 ( .A(n166), .B(n152), .Z(n155) );
  XOR U96 ( .A(n167), .B(n168), .Z(n152) );
  AND U97 ( .A(n169), .B(n170), .Z(n168) );
  XOR U98 ( .A(p_input[73]), .B(n167), .Z(n170) );
  XOR U99 ( .A(n171), .B(n172), .Z(n167) );
  AND U100 ( .A(n173), .B(n174), .Z(n172) );
  IV U101 ( .A(n163), .Z(n166) );
  XOR U102 ( .A(n175), .B(n176), .Z(n163) );
  AND U103 ( .A(n177), .B(n178), .Z(n176) );
  XOR U104 ( .A(n179), .B(n180), .Z(n160) );
  AND U105 ( .A(n181), .B(n178), .Z(n180) );
  XNOR U106 ( .A(n179), .B(n175), .Z(n178) );
  XOR U107 ( .A(n182), .B(n183), .Z(n175) );
  AND U108 ( .A(n184), .B(n174), .Z(n183) );
  XNOR U109 ( .A(n185), .B(n171), .Z(n174) );
  XOR U110 ( .A(n186), .B(n187), .Z(n171) );
  AND U111 ( .A(n188), .B(n189), .Z(n187) );
  XOR U112 ( .A(p_input[105]), .B(n186), .Z(n189) );
  XOR U113 ( .A(n190), .B(n191), .Z(n186) );
  AND U114 ( .A(n192), .B(n193), .Z(n191) );
  IV U115 ( .A(n182), .Z(n185) );
  XOR U116 ( .A(n194), .B(n195), .Z(n182) );
  AND U117 ( .A(n196), .B(n197), .Z(n195) );
  XOR U118 ( .A(n198), .B(n199), .Z(n179) );
  AND U119 ( .A(n200), .B(n197), .Z(n199) );
  XNOR U120 ( .A(n198), .B(n194), .Z(n197) );
  XOR U121 ( .A(n201), .B(n202), .Z(n194) );
  AND U122 ( .A(n203), .B(n193), .Z(n202) );
  XNOR U123 ( .A(n204), .B(n190), .Z(n193) );
  XOR U124 ( .A(n205), .B(n206), .Z(n190) );
  AND U125 ( .A(n207), .B(n208), .Z(n206) );
  XOR U126 ( .A(p_input[137]), .B(n205), .Z(n208) );
  XOR U127 ( .A(n209), .B(n210), .Z(n205) );
  AND U128 ( .A(n211), .B(n212), .Z(n210) );
  IV U129 ( .A(n201), .Z(n204) );
  XOR U130 ( .A(n213), .B(n214), .Z(n201) );
  AND U131 ( .A(n215), .B(n216), .Z(n214) );
  XOR U132 ( .A(n217), .B(n218), .Z(n198) );
  AND U133 ( .A(n219), .B(n216), .Z(n218) );
  XNOR U134 ( .A(n217), .B(n213), .Z(n216) );
  XOR U135 ( .A(n220), .B(n221), .Z(n213) );
  AND U136 ( .A(n222), .B(n212), .Z(n221) );
  XNOR U137 ( .A(n223), .B(n209), .Z(n212) );
  XOR U138 ( .A(n224), .B(n225), .Z(n209) );
  AND U139 ( .A(n226), .B(n227), .Z(n225) );
  XOR U140 ( .A(p_input[169]), .B(n224), .Z(n227) );
  XOR U141 ( .A(n228), .B(n229), .Z(n224) );
  AND U142 ( .A(n230), .B(n231), .Z(n229) );
  IV U143 ( .A(n220), .Z(n223) );
  XOR U144 ( .A(n232), .B(n233), .Z(n220) );
  AND U145 ( .A(n234), .B(n235), .Z(n233) );
  XOR U146 ( .A(n236), .B(n237), .Z(n217) );
  AND U147 ( .A(n238), .B(n235), .Z(n237) );
  XNOR U148 ( .A(n236), .B(n232), .Z(n235) );
  XOR U149 ( .A(n239), .B(n240), .Z(n232) );
  AND U150 ( .A(n241), .B(n231), .Z(n240) );
  XNOR U151 ( .A(n242), .B(n228), .Z(n231) );
  XOR U152 ( .A(n243), .B(n244), .Z(n228) );
  AND U153 ( .A(n245), .B(n246), .Z(n244) );
  XOR U154 ( .A(p_input[201]), .B(n243), .Z(n246) );
  XOR U155 ( .A(n247), .B(n248), .Z(n243) );
  AND U156 ( .A(n249), .B(n250), .Z(n248) );
  IV U157 ( .A(n239), .Z(n242) );
  XOR U158 ( .A(n251), .B(n252), .Z(n239) );
  AND U159 ( .A(n253), .B(n254), .Z(n252) );
  XOR U160 ( .A(n255), .B(n256), .Z(n236) );
  AND U161 ( .A(n257), .B(n254), .Z(n256) );
  XNOR U162 ( .A(n255), .B(n251), .Z(n254) );
  XOR U163 ( .A(n258), .B(n259), .Z(n251) );
  AND U164 ( .A(n260), .B(n250), .Z(n259) );
  XNOR U165 ( .A(n261), .B(n247), .Z(n250) );
  XOR U166 ( .A(n262), .B(n263), .Z(n247) );
  AND U167 ( .A(n264), .B(n265), .Z(n263) );
  XOR U168 ( .A(p_input[233]), .B(n262), .Z(n265) );
  XOR U169 ( .A(n266), .B(n267), .Z(n262) );
  AND U170 ( .A(n268), .B(n269), .Z(n267) );
  IV U171 ( .A(n258), .Z(n261) );
  XOR U172 ( .A(n270), .B(n271), .Z(n258) );
  AND U173 ( .A(n272), .B(n273), .Z(n271) );
  XOR U174 ( .A(n274), .B(n275), .Z(n255) );
  AND U175 ( .A(n276), .B(n273), .Z(n275) );
  XNOR U176 ( .A(n274), .B(n270), .Z(n273) );
  XOR U177 ( .A(n277), .B(n278), .Z(n270) );
  AND U178 ( .A(n279), .B(n269), .Z(n278) );
  XNOR U179 ( .A(n280), .B(n266), .Z(n269) );
  XOR U180 ( .A(n281), .B(n282), .Z(n266) );
  AND U181 ( .A(n283), .B(n284), .Z(n282) );
  XOR U182 ( .A(p_input[265]), .B(n281), .Z(n284) );
  XOR U183 ( .A(n285), .B(n286), .Z(n281) );
  AND U184 ( .A(n287), .B(n288), .Z(n286) );
  IV U185 ( .A(n277), .Z(n280) );
  XOR U186 ( .A(n289), .B(n290), .Z(n277) );
  AND U187 ( .A(n291), .B(n292), .Z(n290) );
  XOR U188 ( .A(n293), .B(n294), .Z(n274) );
  AND U189 ( .A(n295), .B(n292), .Z(n294) );
  XNOR U190 ( .A(n293), .B(n289), .Z(n292) );
  XOR U191 ( .A(n296), .B(n297), .Z(n289) );
  AND U192 ( .A(n298), .B(n288), .Z(n297) );
  XNOR U193 ( .A(n299), .B(n285), .Z(n288) );
  XOR U194 ( .A(n300), .B(n301), .Z(n285) );
  AND U195 ( .A(n302), .B(n303), .Z(n301) );
  XOR U196 ( .A(p_input[297]), .B(n300), .Z(n303) );
  XOR U197 ( .A(n304), .B(n305), .Z(n300) );
  AND U198 ( .A(n306), .B(n307), .Z(n305) );
  IV U199 ( .A(n296), .Z(n299) );
  XOR U200 ( .A(n308), .B(n309), .Z(n296) );
  AND U201 ( .A(n310), .B(n311), .Z(n309) );
  XOR U202 ( .A(n312), .B(n313), .Z(n293) );
  AND U203 ( .A(n314), .B(n311), .Z(n313) );
  XNOR U204 ( .A(n312), .B(n308), .Z(n311) );
  XOR U205 ( .A(n315), .B(n316), .Z(n308) );
  AND U206 ( .A(n317), .B(n307), .Z(n316) );
  XNOR U207 ( .A(n318), .B(n304), .Z(n307) );
  XOR U208 ( .A(n319), .B(n320), .Z(n304) );
  AND U209 ( .A(n321), .B(n322), .Z(n320) );
  XOR U210 ( .A(p_input[329]), .B(n319), .Z(n322) );
  XOR U211 ( .A(n323), .B(n324), .Z(n319) );
  AND U212 ( .A(n325), .B(n326), .Z(n324) );
  IV U213 ( .A(n315), .Z(n318) );
  XOR U214 ( .A(n327), .B(n328), .Z(n315) );
  AND U215 ( .A(n329), .B(n330), .Z(n328) );
  XOR U216 ( .A(n331), .B(n332), .Z(n312) );
  AND U217 ( .A(n333), .B(n330), .Z(n332) );
  XNOR U218 ( .A(n331), .B(n327), .Z(n330) );
  XOR U219 ( .A(n334), .B(n335), .Z(n327) );
  AND U220 ( .A(n336), .B(n326), .Z(n335) );
  XNOR U221 ( .A(n337), .B(n323), .Z(n326) );
  XOR U222 ( .A(n338), .B(n339), .Z(n323) );
  AND U223 ( .A(n340), .B(n341), .Z(n339) );
  XOR U224 ( .A(p_input[361]), .B(n338), .Z(n341) );
  XOR U225 ( .A(n342), .B(n343), .Z(n338) );
  AND U226 ( .A(n344), .B(n345), .Z(n343) );
  IV U227 ( .A(n334), .Z(n337) );
  XOR U228 ( .A(n346), .B(n347), .Z(n334) );
  AND U229 ( .A(n348), .B(n349), .Z(n347) );
  XOR U230 ( .A(n350), .B(n351), .Z(n331) );
  AND U231 ( .A(n352), .B(n349), .Z(n351) );
  XNOR U232 ( .A(n350), .B(n346), .Z(n349) );
  XOR U233 ( .A(n353), .B(n354), .Z(n346) );
  AND U234 ( .A(n355), .B(n345), .Z(n354) );
  XNOR U235 ( .A(n356), .B(n342), .Z(n345) );
  XOR U236 ( .A(n357), .B(n358), .Z(n342) );
  AND U237 ( .A(n359), .B(n360), .Z(n358) );
  XOR U238 ( .A(p_input[393]), .B(n357), .Z(n360) );
  XOR U239 ( .A(n361), .B(n362), .Z(n357) );
  AND U240 ( .A(n363), .B(n364), .Z(n362) );
  IV U241 ( .A(n353), .Z(n356) );
  XOR U242 ( .A(n365), .B(n366), .Z(n353) );
  AND U243 ( .A(n367), .B(n368), .Z(n366) );
  XOR U244 ( .A(n369), .B(n370), .Z(n350) );
  AND U245 ( .A(n371), .B(n368), .Z(n370) );
  XNOR U246 ( .A(n369), .B(n365), .Z(n368) );
  XOR U247 ( .A(n372), .B(n373), .Z(n365) );
  AND U248 ( .A(n374), .B(n364), .Z(n373) );
  XNOR U249 ( .A(n375), .B(n361), .Z(n364) );
  XOR U250 ( .A(n376), .B(n377), .Z(n361) );
  AND U251 ( .A(n378), .B(n379), .Z(n377) );
  XOR U252 ( .A(p_input[425]), .B(n376), .Z(n379) );
  XOR U253 ( .A(n380), .B(n381), .Z(n376) );
  AND U254 ( .A(n382), .B(n383), .Z(n381) );
  IV U255 ( .A(n372), .Z(n375) );
  XOR U256 ( .A(n384), .B(n385), .Z(n372) );
  AND U257 ( .A(n386), .B(n387), .Z(n385) );
  XOR U258 ( .A(n388), .B(n389), .Z(n369) );
  AND U259 ( .A(n390), .B(n387), .Z(n389) );
  XNOR U260 ( .A(n388), .B(n384), .Z(n387) );
  XOR U261 ( .A(n391), .B(n392), .Z(n384) );
  AND U262 ( .A(n393), .B(n383), .Z(n392) );
  XNOR U263 ( .A(n394), .B(n380), .Z(n383) );
  XOR U264 ( .A(n395), .B(n396), .Z(n380) );
  AND U265 ( .A(n397), .B(n398), .Z(n396) );
  XOR U266 ( .A(p_input[457]), .B(n395), .Z(n398) );
  XOR U267 ( .A(n399), .B(n400), .Z(n395) );
  AND U268 ( .A(n401), .B(n402), .Z(n400) );
  IV U269 ( .A(n391), .Z(n394) );
  XOR U270 ( .A(n403), .B(n404), .Z(n391) );
  AND U271 ( .A(n405), .B(n406), .Z(n404) );
  XOR U272 ( .A(n407), .B(n408), .Z(n388) );
  AND U273 ( .A(n409), .B(n406), .Z(n408) );
  XNOR U274 ( .A(n407), .B(n403), .Z(n406) );
  XOR U275 ( .A(n410), .B(n411), .Z(n403) );
  AND U276 ( .A(n412), .B(n402), .Z(n411) );
  XNOR U277 ( .A(n413), .B(n399), .Z(n402) );
  XOR U278 ( .A(n414), .B(n415), .Z(n399) );
  AND U279 ( .A(n416), .B(n417), .Z(n415) );
  XOR U280 ( .A(p_input[489]), .B(n414), .Z(n417) );
  XOR U281 ( .A(n418), .B(n419), .Z(n414) );
  AND U282 ( .A(n420), .B(n421), .Z(n419) );
  IV U283 ( .A(n410), .Z(n413) );
  XOR U284 ( .A(n422), .B(n423), .Z(n410) );
  AND U285 ( .A(n424), .B(n425), .Z(n423) );
  XOR U286 ( .A(n426), .B(n427), .Z(n407) );
  AND U287 ( .A(n428), .B(n425), .Z(n427) );
  XNOR U288 ( .A(n426), .B(n422), .Z(n425) );
  XOR U289 ( .A(n429), .B(n430), .Z(n422) );
  AND U290 ( .A(n431), .B(n421), .Z(n430) );
  XNOR U291 ( .A(n432), .B(n418), .Z(n421) );
  XOR U292 ( .A(n433), .B(n434), .Z(n418) );
  AND U293 ( .A(n435), .B(n436), .Z(n434) );
  XOR U294 ( .A(p_input[521]), .B(n433), .Z(n436) );
  XOR U295 ( .A(n437), .B(n438), .Z(n433) );
  AND U296 ( .A(n439), .B(n440), .Z(n438) );
  IV U297 ( .A(n429), .Z(n432) );
  XOR U298 ( .A(n441), .B(n442), .Z(n429) );
  AND U299 ( .A(n443), .B(n444), .Z(n442) );
  XOR U300 ( .A(n445), .B(n446), .Z(n426) );
  AND U301 ( .A(n447), .B(n444), .Z(n446) );
  XNOR U302 ( .A(n445), .B(n441), .Z(n444) );
  XOR U303 ( .A(n448), .B(n449), .Z(n441) );
  AND U304 ( .A(n450), .B(n440), .Z(n449) );
  XNOR U305 ( .A(n451), .B(n437), .Z(n440) );
  XOR U306 ( .A(n452), .B(n453), .Z(n437) );
  AND U307 ( .A(n454), .B(n455), .Z(n453) );
  XOR U308 ( .A(p_input[553]), .B(n452), .Z(n455) );
  XOR U309 ( .A(n456), .B(n457), .Z(n452) );
  AND U310 ( .A(n458), .B(n459), .Z(n457) );
  IV U311 ( .A(n448), .Z(n451) );
  XOR U312 ( .A(n460), .B(n461), .Z(n448) );
  AND U313 ( .A(n462), .B(n463), .Z(n461) );
  XOR U314 ( .A(n464), .B(n465), .Z(n445) );
  AND U315 ( .A(n466), .B(n463), .Z(n465) );
  XNOR U316 ( .A(n464), .B(n460), .Z(n463) );
  XOR U317 ( .A(n467), .B(n468), .Z(n460) );
  AND U318 ( .A(n469), .B(n459), .Z(n468) );
  XNOR U319 ( .A(n470), .B(n456), .Z(n459) );
  XOR U320 ( .A(n471), .B(n472), .Z(n456) );
  AND U321 ( .A(n473), .B(n474), .Z(n472) );
  XOR U322 ( .A(p_input[585]), .B(n471), .Z(n474) );
  XOR U323 ( .A(n475), .B(n476), .Z(n471) );
  AND U324 ( .A(n477), .B(n478), .Z(n476) );
  IV U325 ( .A(n467), .Z(n470) );
  XOR U326 ( .A(n479), .B(n480), .Z(n467) );
  AND U327 ( .A(n481), .B(n482), .Z(n480) );
  XOR U328 ( .A(n483), .B(n484), .Z(n464) );
  AND U329 ( .A(n485), .B(n482), .Z(n484) );
  XNOR U330 ( .A(n483), .B(n479), .Z(n482) );
  XOR U331 ( .A(n486), .B(n487), .Z(n479) );
  AND U332 ( .A(n488), .B(n478), .Z(n487) );
  XNOR U333 ( .A(n489), .B(n475), .Z(n478) );
  XOR U334 ( .A(n490), .B(n491), .Z(n475) );
  AND U335 ( .A(n492), .B(n493), .Z(n491) );
  XOR U336 ( .A(p_input[617]), .B(n490), .Z(n493) );
  XOR U337 ( .A(n494), .B(n495), .Z(n490) );
  AND U338 ( .A(n496), .B(n497), .Z(n495) );
  IV U339 ( .A(n486), .Z(n489) );
  XOR U340 ( .A(n498), .B(n499), .Z(n486) );
  AND U341 ( .A(n500), .B(n501), .Z(n499) );
  XOR U342 ( .A(n502), .B(n503), .Z(n483) );
  AND U343 ( .A(n504), .B(n501), .Z(n503) );
  XNOR U344 ( .A(n502), .B(n498), .Z(n501) );
  XOR U345 ( .A(n505), .B(n506), .Z(n498) );
  AND U346 ( .A(n507), .B(n497), .Z(n506) );
  XNOR U347 ( .A(n508), .B(n494), .Z(n497) );
  XOR U348 ( .A(n509), .B(n510), .Z(n494) );
  AND U349 ( .A(n511), .B(n512), .Z(n510) );
  XOR U350 ( .A(p_input[649]), .B(n509), .Z(n512) );
  XOR U351 ( .A(n513), .B(n514), .Z(n509) );
  AND U352 ( .A(n515), .B(n516), .Z(n514) );
  IV U353 ( .A(n505), .Z(n508) );
  XOR U354 ( .A(n517), .B(n518), .Z(n505) );
  AND U355 ( .A(n519), .B(n520), .Z(n518) );
  XOR U356 ( .A(n521), .B(n522), .Z(n502) );
  AND U357 ( .A(n523), .B(n520), .Z(n522) );
  XNOR U358 ( .A(n521), .B(n517), .Z(n520) );
  XOR U359 ( .A(n524), .B(n525), .Z(n517) );
  AND U360 ( .A(n526), .B(n516), .Z(n525) );
  XNOR U361 ( .A(n527), .B(n513), .Z(n516) );
  XOR U362 ( .A(n528), .B(n529), .Z(n513) );
  AND U363 ( .A(n530), .B(n531), .Z(n529) );
  XOR U364 ( .A(p_input[681]), .B(n528), .Z(n531) );
  XOR U365 ( .A(n532), .B(n533), .Z(n528) );
  AND U366 ( .A(n534), .B(n535), .Z(n533) );
  IV U367 ( .A(n524), .Z(n527) );
  XOR U368 ( .A(n536), .B(n537), .Z(n524) );
  AND U369 ( .A(n538), .B(n539), .Z(n537) );
  XOR U370 ( .A(n540), .B(n541), .Z(n521) );
  AND U371 ( .A(n542), .B(n539), .Z(n541) );
  XNOR U372 ( .A(n540), .B(n536), .Z(n539) );
  XOR U373 ( .A(n543), .B(n544), .Z(n536) );
  AND U374 ( .A(n545), .B(n535), .Z(n544) );
  XNOR U375 ( .A(n546), .B(n532), .Z(n535) );
  XOR U376 ( .A(n547), .B(n548), .Z(n532) );
  AND U377 ( .A(n549), .B(n550), .Z(n548) );
  XOR U378 ( .A(p_input[713]), .B(n547), .Z(n550) );
  XOR U379 ( .A(n551), .B(n552), .Z(n547) );
  AND U380 ( .A(n553), .B(n554), .Z(n552) );
  IV U381 ( .A(n543), .Z(n546) );
  XOR U382 ( .A(n555), .B(n556), .Z(n543) );
  AND U383 ( .A(n557), .B(n558), .Z(n556) );
  XOR U384 ( .A(n559), .B(n560), .Z(n540) );
  AND U385 ( .A(n561), .B(n558), .Z(n560) );
  XNOR U386 ( .A(n559), .B(n555), .Z(n558) );
  XOR U387 ( .A(n562), .B(n563), .Z(n555) );
  AND U388 ( .A(n564), .B(n554), .Z(n563) );
  XNOR U389 ( .A(n565), .B(n551), .Z(n554) );
  XOR U390 ( .A(n566), .B(n567), .Z(n551) );
  AND U391 ( .A(n568), .B(n569), .Z(n567) );
  XOR U392 ( .A(p_input[745]), .B(n566), .Z(n569) );
  XOR U393 ( .A(n570), .B(n571), .Z(n566) );
  AND U394 ( .A(n572), .B(n573), .Z(n571) );
  IV U395 ( .A(n562), .Z(n565) );
  XOR U396 ( .A(n574), .B(n575), .Z(n562) );
  AND U397 ( .A(n576), .B(n577), .Z(n575) );
  XOR U398 ( .A(n578), .B(n579), .Z(n559) );
  AND U399 ( .A(n580), .B(n577), .Z(n579) );
  XNOR U400 ( .A(n578), .B(n574), .Z(n577) );
  XOR U401 ( .A(n581), .B(n582), .Z(n574) );
  AND U402 ( .A(n583), .B(n573), .Z(n582) );
  XNOR U403 ( .A(n584), .B(n570), .Z(n573) );
  XOR U404 ( .A(n585), .B(n586), .Z(n570) );
  AND U405 ( .A(n587), .B(n588), .Z(n586) );
  XOR U406 ( .A(p_input[777]), .B(n585), .Z(n588) );
  XOR U407 ( .A(n589), .B(n590), .Z(n585) );
  AND U408 ( .A(n591), .B(n592), .Z(n590) );
  IV U409 ( .A(n581), .Z(n584) );
  XOR U410 ( .A(n593), .B(n594), .Z(n581) );
  AND U411 ( .A(n595), .B(n596), .Z(n594) );
  XOR U412 ( .A(n597), .B(n598), .Z(n578) );
  AND U413 ( .A(n599), .B(n596), .Z(n598) );
  XNOR U414 ( .A(n597), .B(n593), .Z(n596) );
  XOR U415 ( .A(n600), .B(n601), .Z(n593) );
  AND U416 ( .A(n602), .B(n592), .Z(n601) );
  XNOR U417 ( .A(n603), .B(n589), .Z(n592) );
  XOR U418 ( .A(n604), .B(n605), .Z(n589) );
  AND U419 ( .A(n606), .B(n607), .Z(n605) );
  XOR U420 ( .A(p_input[809]), .B(n604), .Z(n607) );
  XOR U421 ( .A(n608), .B(n609), .Z(n604) );
  AND U422 ( .A(n610), .B(n611), .Z(n609) );
  IV U423 ( .A(n600), .Z(n603) );
  XOR U424 ( .A(n612), .B(n613), .Z(n600) );
  AND U425 ( .A(n614), .B(n615), .Z(n613) );
  XOR U426 ( .A(n616), .B(n617), .Z(n597) );
  AND U427 ( .A(n618), .B(n615), .Z(n617) );
  XNOR U428 ( .A(n616), .B(n612), .Z(n615) );
  XOR U429 ( .A(n619), .B(n620), .Z(n612) );
  AND U430 ( .A(n621), .B(n611), .Z(n620) );
  XNOR U431 ( .A(n622), .B(n608), .Z(n611) );
  XOR U432 ( .A(n623), .B(n624), .Z(n608) );
  AND U433 ( .A(n625), .B(n626), .Z(n624) );
  XOR U434 ( .A(p_input[841]), .B(n623), .Z(n626) );
  XOR U435 ( .A(n627), .B(n628), .Z(n623) );
  AND U436 ( .A(n629), .B(n630), .Z(n628) );
  IV U437 ( .A(n619), .Z(n622) );
  XOR U438 ( .A(n631), .B(n632), .Z(n619) );
  AND U439 ( .A(n633), .B(n634), .Z(n632) );
  XOR U440 ( .A(n635), .B(n636), .Z(n616) );
  AND U441 ( .A(n637), .B(n634), .Z(n636) );
  XNOR U442 ( .A(n635), .B(n631), .Z(n634) );
  XOR U443 ( .A(n638), .B(n639), .Z(n631) );
  AND U444 ( .A(n640), .B(n630), .Z(n639) );
  XNOR U445 ( .A(n641), .B(n627), .Z(n630) );
  XOR U446 ( .A(n642), .B(n643), .Z(n627) );
  AND U447 ( .A(n644), .B(n645), .Z(n643) );
  XOR U448 ( .A(p_input[873]), .B(n642), .Z(n645) );
  XOR U449 ( .A(n646), .B(n647), .Z(n642) );
  AND U450 ( .A(n648), .B(n649), .Z(n647) );
  IV U451 ( .A(n638), .Z(n641) );
  XOR U452 ( .A(n650), .B(n651), .Z(n638) );
  AND U453 ( .A(n652), .B(n653), .Z(n651) );
  XOR U454 ( .A(n654), .B(n655), .Z(n635) );
  AND U455 ( .A(n656), .B(n653), .Z(n655) );
  XNOR U456 ( .A(n654), .B(n650), .Z(n653) );
  XOR U457 ( .A(n657), .B(n658), .Z(n650) );
  AND U458 ( .A(n659), .B(n649), .Z(n658) );
  XNOR U459 ( .A(n660), .B(n646), .Z(n649) );
  XOR U460 ( .A(n661), .B(n662), .Z(n646) );
  AND U461 ( .A(n663), .B(n664), .Z(n662) );
  XOR U462 ( .A(p_input[905]), .B(n661), .Z(n664) );
  XOR U463 ( .A(n665), .B(n666), .Z(n661) );
  AND U464 ( .A(n667), .B(n668), .Z(n666) );
  IV U465 ( .A(n657), .Z(n660) );
  XOR U466 ( .A(n669), .B(n670), .Z(n657) );
  AND U467 ( .A(n671), .B(n672), .Z(n670) );
  XOR U468 ( .A(n673), .B(n674), .Z(n654) );
  AND U469 ( .A(n675), .B(n672), .Z(n674) );
  XNOR U470 ( .A(n673), .B(n669), .Z(n672) );
  XOR U471 ( .A(n676), .B(n677), .Z(n669) );
  AND U472 ( .A(n678), .B(n668), .Z(n677) );
  XNOR U473 ( .A(n679), .B(n665), .Z(n668) );
  XOR U474 ( .A(n680), .B(n681), .Z(n665) );
  AND U475 ( .A(n682), .B(n683), .Z(n681) );
  XOR U476 ( .A(p_input[937]), .B(n680), .Z(n683) );
  XOR U477 ( .A(n684), .B(n685), .Z(n680) );
  AND U478 ( .A(n686), .B(n687), .Z(n685) );
  IV U479 ( .A(n676), .Z(n679) );
  XOR U480 ( .A(n688), .B(n689), .Z(n676) );
  AND U481 ( .A(n690), .B(n691), .Z(n689) );
  XOR U482 ( .A(n692), .B(n693), .Z(n673) );
  AND U483 ( .A(n694), .B(n691), .Z(n693) );
  XNOR U484 ( .A(n692), .B(n688), .Z(n691) );
  XOR U485 ( .A(n695), .B(n696), .Z(n688) );
  AND U486 ( .A(n697), .B(n687), .Z(n696) );
  XNOR U487 ( .A(n698), .B(n684), .Z(n687) );
  XOR U488 ( .A(n699), .B(n700), .Z(n684) );
  AND U489 ( .A(n701), .B(n702), .Z(n700) );
  XOR U490 ( .A(p_input[969]), .B(n699), .Z(n702) );
  XOR U491 ( .A(n703), .B(n704), .Z(n699) );
  AND U492 ( .A(n705), .B(n706), .Z(n704) );
  IV U493 ( .A(n695), .Z(n698) );
  XOR U494 ( .A(n707), .B(n708), .Z(n695) );
  AND U495 ( .A(n709), .B(n710), .Z(n708) );
  XOR U496 ( .A(n711), .B(n712), .Z(n692) );
  AND U497 ( .A(n713), .B(n710), .Z(n712) );
  XNOR U498 ( .A(n711), .B(n707), .Z(n710) );
  XOR U499 ( .A(n714), .B(n715), .Z(n707) );
  AND U500 ( .A(n716), .B(n706), .Z(n715) );
  XNOR U501 ( .A(n717), .B(n703), .Z(n706) );
  XOR U502 ( .A(n718), .B(n719), .Z(n703) );
  AND U503 ( .A(n720), .B(n721), .Z(n719) );
  XOR U504 ( .A(p_input[1001]), .B(n718), .Z(n721) );
  XOR U505 ( .A(n722), .B(n723), .Z(n718) );
  AND U506 ( .A(n724), .B(n725), .Z(n723) );
  IV U507 ( .A(n714), .Z(n717) );
  XOR U508 ( .A(n726), .B(n727), .Z(n714) );
  AND U509 ( .A(n728), .B(n729), .Z(n727) );
  XOR U510 ( .A(n730), .B(n731), .Z(n711) );
  AND U511 ( .A(n732), .B(n729), .Z(n731) );
  XNOR U512 ( .A(n730), .B(n726), .Z(n729) );
  XOR U513 ( .A(n733), .B(n734), .Z(n726) );
  AND U514 ( .A(n735), .B(n725), .Z(n734) );
  XNOR U515 ( .A(n736), .B(n722), .Z(n725) );
  XOR U516 ( .A(n737), .B(n738), .Z(n722) );
  AND U517 ( .A(n739), .B(n740), .Z(n738) );
  XOR U518 ( .A(p_input[1033]), .B(n737), .Z(n740) );
  XOR U519 ( .A(n741), .B(n742), .Z(n737) );
  AND U520 ( .A(n743), .B(n744), .Z(n742) );
  IV U521 ( .A(n733), .Z(n736) );
  XOR U522 ( .A(n745), .B(n746), .Z(n733) );
  AND U523 ( .A(n747), .B(n748), .Z(n746) );
  XOR U524 ( .A(n749), .B(n750), .Z(n730) );
  AND U525 ( .A(n751), .B(n748), .Z(n750) );
  XNOR U526 ( .A(n749), .B(n745), .Z(n748) );
  XOR U527 ( .A(n752), .B(n753), .Z(n745) );
  AND U528 ( .A(n754), .B(n744), .Z(n753) );
  XNOR U529 ( .A(n755), .B(n741), .Z(n744) );
  XOR U530 ( .A(n756), .B(n757), .Z(n741) );
  AND U531 ( .A(n758), .B(n759), .Z(n757) );
  XOR U532 ( .A(p_input[1065]), .B(n756), .Z(n759) );
  XOR U533 ( .A(n760), .B(n761), .Z(n756) );
  AND U534 ( .A(n762), .B(n763), .Z(n761) );
  IV U535 ( .A(n752), .Z(n755) );
  XOR U536 ( .A(n764), .B(n765), .Z(n752) );
  AND U537 ( .A(n766), .B(n767), .Z(n765) );
  XOR U538 ( .A(n768), .B(n769), .Z(n749) );
  AND U539 ( .A(n770), .B(n767), .Z(n769) );
  XNOR U540 ( .A(n768), .B(n764), .Z(n767) );
  XOR U541 ( .A(n771), .B(n772), .Z(n764) );
  AND U542 ( .A(n773), .B(n763), .Z(n772) );
  XNOR U543 ( .A(n774), .B(n760), .Z(n763) );
  XOR U544 ( .A(n775), .B(n776), .Z(n760) );
  AND U545 ( .A(n777), .B(n778), .Z(n776) );
  XOR U546 ( .A(p_input[1097]), .B(n775), .Z(n778) );
  XOR U547 ( .A(n779), .B(n780), .Z(n775) );
  AND U548 ( .A(n781), .B(n782), .Z(n780) );
  IV U549 ( .A(n771), .Z(n774) );
  XOR U550 ( .A(n783), .B(n784), .Z(n771) );
  AND U551 ( .A(n785), .B(n786), .Z(n784) );
  XOR U552 ( .A(n787), .B(n788), .Z(n768) );
  AND U553 ( .A(n789), .B(n786), .Z(n788) );
  XNOR U554 ( .A(n787), .B(n783), .Z(n786) );
  XOR U555 ( .A(n790), .B(n791), .Z(n783) );
  AND U556 ( .A(n792), .B(n782), .Z(n791) );
  XNOR U557 ( .A(n793), .B(n779), .Z(n782) );
  XOR U558 ( .A(n794), .B(n795), .Z(n779) );
  AND U559 ( .A(n796), .B(n797), .Z(n795) );
  XOR U560 ( .A(p_input[1129]), .B(n794), .Z(n797) );
  XOR U561 ( .A(n798), .B(n799), .Z(n794) );
  AND U562 ( .A(n800), .B(n801), .Z(n799) );
  IV U563 ( .A(n790), .Z(n793) );
  XOR U564 ( .A(n802), .B(n803), .Z(n790) );
  AND U565 ( .A(n804), .B(n805), .Z(n803) );
  XOR U566 ( .A(n806), .B(n807), .Z(n787) );
  AND U567 ( .A(n808), .B(n805), .Z(n807) );
  XNOR U568 ( .A(n806), .B(n802), .Z(n805) );
  XOR U569 ( .A(n809), .B(n810), .Z(n802) );
  AND U570 ( .A(n811), .B(n801), .Z(n810) );
  XNOR U571 ( .A(n812), .B(n798), .Z(n801) );
  XOR U572 ( .A(n813), .B(n814), .Z(n798) );
  AND U573 ( .A(n815), .B(n816), .Z(n814) );
  XOR U574 ( .A(p_input[1161]), .B(n813), .Z(n816) );
  XOR U575 ( .A(n817), .B(n818), .Z(n813) );
  AND U576 ( .A(n819), .B(n820), .Z(n818) );
  IV U577 ( .A(n809), .Z(n812) );
  XOR U578 ( .A(n821), .B(n822), .Z(n809) );
  AND U579 ( .A(n823), .B(n824), .Z(n822) );
  XOR U580 ( .A(n825), .B(n826), .Z(n806) );
  AND U581 ( .A(n827), .B(n824), .Z(n826) );
  XNOR U582 ( .A(n825), .B(n821), .Z(n824) );
  XOR U583 ( .A(n828), .B(n829), .Z(n821) );
  AND U584 ( .A(n830), .B(n820), .Z(n829) );
  XNOR U585 ( .A(n831), .B(n817), .Z(n820) );
  XOR U586 ( .A(n832), .B(n833), .Z(n817) );
  AND U587 ( .A(n834), .B(n835), .Z(n833) );
  XOR U588 ( .A(p_input[1193]), .B(n832), .Z(n835) );
  XOR U589 ( .A(n836), .B(n837), .Z(n832) );
  AND U590 ( .A(n838), .B(n839), .Z(n837) );
  IV U591 ( .A(n828), .Z(n831) );
  XOR U592 ( .A(n840), .B(n841), .Z(n828) );
  AND U593 ( .A(n842), .B(n843), .Z(n841) );
  XOR U594 ( .A(n844), .B(n845), .Z(n825) );
  AND U595 ( .A(n846), .B(n843), .Z(n845) );
  XNOR U596 ( .A(n844), .B(n840), .Z(n843) );
  XOR U597 ( .A(n847), .B(n848), .Z(n840) );
  AND U598 ( .A(n849), .B(n839), .Z(n848) );
  XNOR U599 ( .A(n850), .B(n836), .Z(n839) );
  XOR U600 ( .A(n851), .B(n852), .Z(n836) );
  AND U601 ( .A(n853), .B(n854), .Z(n852) );
  XOR U602 ( .A(p_input[1225]), .B(n851), .Z(n854) );
  XOR U603 ( .A(n855), .B(n856), .Z(n851) );
  AND U604 ( .A(n857), .B(n858), .Z(n856) );
  IV U605 ( .A(n847), .Z(n850) );
  XOR U606 ( .A(n859), .B(n860), .Z(n847) );
  AND U607 ( .A(n861), .B(n862), .Z(n860) );
  XOR U608 ( .A(n863), .B(n864), .Z(n844) );
  AND U609 ( .A(n865), .B(n862), .Z(n864) );
  XNOR U610 ( .A(n863), .B(n859), .Z(n862) );
  XOR U611 ( .A(n866), .B(n867), .Z(n859) );
  AND U612 ( .A(n868), .B(n858), .Z(n867) );
  XNOR U613 ( .A(n869), .B(n855), .Z(n858) );
  XOR U614 ( .A(n870), .B(n871), .Z(n855) );
  AND U615 ( .A(n872), .B(n873), .Z(n871) );
  XOR U616 ( .A(p_input[1257]), .B(n870), .Z(n873) );
  XOR U617 ( .A(n874), .B(n875), .Z(n870) );
  AND U618 ( .A(n876), .B(n877), .Z(n875) );
  IV U619 ( .A(n866), .Z(n869) );
  XOR U620 ( .A(n878), .B(n879), .Z(n866) );
  AND U621 ( .A(n880), .B(n881), .Z(n879) );
  XOR U622 ( .A(n882), .B(n883), .Z(n863) );
  AND U623 ( .A(n884), .B(n881), .Z(n883) );
  XNOR U624 ( .A(n882), .B(n878), .Z(n881) );
  XOR U625 ( .A(n885), .B(n886), .Z(n878) );
  AND U626 ( .A(n887), .B(n877), .Z(n886) );
  XNOR U627 ( .A(n888), .B(n874), .Z(n877) );
  XOR U628 ( .A(n889), .B(n890), .Z(n874) );
  AND U629 ( .A(n891), .B(n892), .Z(n890) );
  XOR U630 ( .A(p_input[1289]), .B(n889), .Z(n892) );
  XOR U631 ( .A(n893), .B(n894), .Z(n889) );
  AND U632 ( .A(n895), .B(n896), .Z(n894) );
  IV U633 ( .A(n885), .Z(n888) );
  XOR U634 ( .A(n897), .B(n898), .Z(n885) );
  AND U635 ( .A(n899), .B(n900), .Z(n898) );
  XOR U636 ( .A(n901), .B(n902), .Z(n882) );
  AND U637 ( .A(n903), .B(n900), .Z(n902) );
  XNOR U638 ( .A(n901), .B(n897), .Z(n900) );
  XOR U639 ( .A(n904), .B(n905), .Z(n897) );
  AND U640 ( .A(n906), .B(n896), .Z(n905) );
  XNOR U641 ( .A(n907), .B(n893), .Z(n896) );
  XOR U642 ( .A(n908), .B(n909), .Z(n893) );
  AND U643 ( .A(n910), .B(n911), .Z(n909) );
  XOR U644 ( .A(p_input[1321]), .B(n908), .Z(n911) );
  XOR U645 ( .A(n912), .B(n913), .Z(n908) );
  AND U646 ( .A(n914), .B(n915), .Z(n913) );
  IV U647 ( .A(n904), .Z(n907) );
  XOR U648 ( .A(n916), .B(n917), .Z(n904) );
  AND U649 ( .A(n918), .B(n919), .Z(n917) );
  XOR U650 ( .A(n920), .B(n921), .Z(n901) );
  AND U651 ( .A(n922), .B(n919), .Z(n921) );
  XNOR U652 ( .A(n920), .B(n916), .Z(n919) );
  XOR U653 ( .A(n923), .B(n924), .Z(n916) );
  AND U654 ( .A(n925), .B(n915), .Z(n924) );
  XNOR U655 ( .A(n926), .B(n912), .Z(n915) );
  XOR U656 ( .A(n927), .B(n928), .Z(n912) );
  AND U657 ( .A(n929), .B(n930), .Z(n928) );
  XOR U658 ( .A(p_input[1353]), .B(n927), .Z(n930) );
  XOR U659 ( .A(n931), .B(n932), .Z(n927) );
  AND U660 ( .A(n933), .B(n934), .Z(n932) );
  IV U661 ( .A(n923), .Z(n926) );
  XOR U662 ( .A(n935), .B(n936), .Z(n923) );
  AND U663 ( .A(n937), .B(n938), .Z(n936) );
  XOR U664 ( .A(n939), .B(n940), .Z(n920) );
  AND U665 ( .A(n941), .B(n938), .Z(n940) );
  XNOR U666 ( .A(n939), .B(n935), .Z(n938) );
  XOR U667 ( .A(n942), .B(n943), .Z(n935) );
  AND U668 ( .A(n944), .B(n934), .Z(n943) );
  XNOR U669 ( .A(n945), .B(n931), .Z(n934) );
  XOR U670 ( .A(n946), .B(n947), .Z(n931) );
  AND U671 ( .A(n948), .B(n949), .Z(n947) );
  XOR U672 ( .A(p_input[1385]), .B(n946), .Z(n949) );
  XOR U673 ( .A(n950), .B(n951), .Z(n946) );
  AND U674 ( .A(n952), .B(n953), .Z(n951) );
  IV U675 ( .A(n942), .Z(n945) );
  XOR U676 ( .A(n954), .B(n955), .Z(n942) );
  AND U677 ( .A(n956), .B(n957), .Z(n955) );
  XOR U678 ( .A(n958), .B(n959), .Z(n939) );
  AND U679 ( .A(n960), .B(n957), .Z(n959) );
  XNOR U680 ( .A(n958), .B(n954), .Z(n957) );
  XOR U681 ( .A(n961), .B(n962), .Z(n954) );
  AND U682 ( .A(n963), .B(n953), .Z(n962) );
  XNOR U683 ( .A(n964), .B(n950), .Z(n953) );
  XOR U684 ( .A(n965), .B(n966), .Z(n950) );
  AND U685 ( .A(n967), .B(n968), .Z(n966) );
  XOR U686 ( .A(p_input[1417]), .B(n965), .Z(n968) );
  XOR U687 ( .A(n969), .B(n970), .Z(n965) );
  AND U688 ( .A(n971), .B(n972), .Z(n970) );
  IV U689 ( .A(n961), .Z(n964) );
  XOR U690 ( .A(n973), .B(n974), .Z(n961) );
  AND U691 ( .A(n975), .B(n976), .Z(n974) );
  XOR U692 ( .A(n977), .B(n978), .Z(n958) );
  AND U693 ( .A(n979), .B(n976), .Z(n978) );
  XNOR U694 ( .A(n977), .B(n973), .Z(n976) );
  XOR U695 ( .A(n980), .B(n981), .Z(n973) );
  AND U696 ( .A(n982), .B(n972), .Z(n981) );
  XNOR U697 ( .A(n983), .B(n969), .Z(n972) );
  XOR U698 ( .A(n984), .B(n985), .Z(n969) );
  AND U699 ( .A(n986), .B(n987), .Z(n985) );
  XOR U700 ( .A(p_input[1449]), .B(n984), .Z(n987) );
  XOR U701 ( .A(n988), .B(n989), .Z(n984) );
  AND U702 ( .A(n990), .B(n991), .Z(n989) );
  IV U703 ( .A(n980), .Z(n983) );
  XOR U704 ( .A(n992), .B(n993), .Z(n980) );
  AND U705 ( .A(n994), .B(n995), .Z(n993) );
  XOR U706 ( .A(n996), .B(n997), .Z(n977) );
  AND U707 ( .A(n998), .B(n995), .Z(n997) );
  XNOR U708 ( .A(n996), .B(n992), .Z(n995) );
  XOR U709 ( .A(n999), .B(n1000), .Z(n992) );
  AND U710 ( .A(n1001), .B(n991), .Z(n1000) );
  XNOR U711 ( .A(n1002), .B(n988), .Z(n991) );
  XOR U712 ( .A(n1003), .B(n1004), .Z(n988) );
  AND U713 ( .A(n1005), .B(n1006), .Z(n1004) );
  XOR U714 ( .A(p_input[1481]), .B(n1003), .Z(n1006) );
  XOR U715 ( .A(n1007), .B(n1008), .Z(n1003) );
  AND U716 ( .A(n1009), .B(n1010), .Z(n1008) );
  IV U717 ( .A(n999), .Z(n1002) );
  XOR U718 ( .A(n1011), .B(n1012), .Z(n999) );
  AND U719 ( .A(n1013), .B(n1014), .Z(n1012) );
  XOR U720 ( .A(n1015), .B(n1016), .Z(n996) );
  AND U721 ( .A(n1017), .B(n1014), .Z(n1016) );
  XNOR U722 ( .A(n1015), .B(n1011), .Z(n1014) );
  XOR U723 ( .A(n1018), .B(n1019), .Z(n1011) );
  AND U724 ( .A(n1020), .B(n1010), .Z(n1019) );
  XNOR U725 ( .A(n1021), .B(n1007), .Z(n1010) );
  XOR U726 ( .A(n1022), .B(n1023), .Z(n1007) );
  AND U727 ( .A(n1024), .B(n1025), .Z(n1023) );
  XOR U728 ( .A(p_input[1513]), .B(n1022), .Z(n1025) );
  XOR U729 ( .A(n1026), .B(n1027), .Z(n1022) );
  AND U730 ( .A(n1028), .B(n1029), .Z(n1027) );
  IV U731 ( .A(n1018), .Z(n1021) );
  XOR U732 ( .A(n1030), .B(n1031), .Z(n1018) );
  AND U733 ( .A(n1032), .B(n1033), .Z(n1031) );
  XOR U734 ( .A(n1034), .B(n1035), .Z(n1015) );
  AND U735 ( .A(n1036), .B(n1033), .Z(n1035) );
  XNOR U736 ( .A(n1034), .B(n1030), .Z(n1033) );
  XOR U737 ( .A(n1037), .B(n1038), .Z(n1030) );
  AND U738 ( .A(n1039), .B(n1029), .Z(n1038) );
  XNOR U739 ( .A(n1040), .B(n1026), .Z(n1029) );
  XOR U740 ( .A(n1041), .B(n1042), .Z(n1026) );
  AND U741 ( .A(n1043), .B(n1044), .Z(n1042) );
  XOR U742 ( .A(p_input[1545]), .B(n1041), .Z(n1044) );
  XOR U743 ( .A(n1045), .B(n1046), .Z(n1041) );
  AND U744 ( .A(n1047), .B(n1048), .Z(n1046) );
  IV U745 ( .A(n1037), .Z(n1040) );
  XOR U746 ( .A(n1049), .B(n1050), .Z(n1037) );
  AND U747 ( .A(n1051), .B(n1052), .Z(n1050) );
  XOR U748 ( .A(n1053), .B(n1054), .Z(n1034) );
  AND U749 ( .A(n1055), .B(n1052), .Z(n1054) );
  XNOR U750 ( .A(n1053), .B(n1049), .Z(n1052) );
  XOR U751 ( .A(n1056), .B(n1057), .Z(n1049) );
  AND U752 ( .A(n1058), .B(n1048), .Z(n1057) );
  XNOR U753 ( .A(n1059), .B(n1045), .Z(n1048) );
  XOR U754 ( .A(n1060), .B(n1061), .Z(n1045) );
  AND U755 ( .A(n1062), .B(n1063), .Z(n1061) );
  XOR U756 ( .A(p_input[1577]), .B(n1060), .Z(n1063) );
  XOR U757 ( .A(n1064), .B(n1065), .Z(n1060) );
  AND U758 ( .A(n1066), .B(n1067), .Z(n1065) );
  IV U759 ( .A(n1056), .Z(n1059) );
  XOR U760 ( .A(n1068), .B(n1069), .Z(n1056) );
  AND U761 ( .A(n1070), .B(n1071), .Z(n1069) );
  XOR U762 ( .A(n1072), .B(n1073), .Z(n1053) );
  AND U763 ( .A(n1074), .B(n1071), .Z(n1073) );
  XNOR U764 ( .A(n1072), .B(n1068), .Z(n1071) );
  XOR U765 ( .A(n1075), .B(n1076), .Z(n1068) );
  AND U766 ( .A(n1077), .B(n1067), .Z(n1076) );
  XNOR U767 ( .A(n1078), .B(n1064), .Z(n1067) );
  XOR U768 ( .A(n1079), .B(n1080), .Z(n1064) );
  AND U769 ( .A(n1081), .B(n1082), .Z(n1080) );
  XOR U770 ( .A(p_input[1609]), .B(n1079), .Z(n1082) );
  XOR U771 ( .A(n1083), .B(n1084), .Z(n1079) );
  AND U772 ( .A(n1085), .B(n1086), .Z(n1084) );
  IV U773 ( .A(n1075), .Z(n1078) );
  XOR U774 ( .A(n1087), .B(n1088), .Z(n1075) );
  AND U775 ( .A(n1089), .B(n1090), .Z(n1088) );
  XOR U776 ( .A(n1091), .B(n1092), .Z(n1072) );
  AND U777 ( .A(n1093), .B(n1090), .Z(n1092) );
  XNOR U778 ( .A(n1091), .B(n1087), .Z(n1090) );
  XOR U779 ( .A(n1094), .B(n1095), .Z(n1087) );
  AND U780 ( .A(n1096), .B(n1086), .Z(n1095) );
  XNOR U781 ( .A(n1097), .B(n1083), .Z(n1086) );
  XOR U782 ( .A(n1098), .B(n1099), .Z(n1083) );
  AND U783 ( .A(n1100), .B(n1101), .Z(n1099) );
  XOR U784 ( .A(p_input[1641]), .B(n1098), .Z(n1101) );
  XOR U785 ( .A(n1102), .B(n1103), .Z(n1098) );
  AND U786 ( .A(n1104), .B(n1105), .Z(n1103) );
  IV U787 ( .A(n1094), .Z(n1097) );
  XOR U788 ( .A(n1106), .B(n1107), .Z(n1094) );
  AND U789 ( .A(n1108), .B(n1109), .Z(n1107) );
  XOR U790 ( .A(n1110), .B(n1111), .Z(n1091) );
  AND U791 ( .A(n1112), .B(n1109), .Z(n1111) );
  XNOR U792 ( .A(n1110), .B(n1106), .Z(n1109) );
  XOR U793 ( .A(n1113), .B(n1114), .Z(n1106) );
  AND U794 ( .A(n1115), .B(n1105), .Z(n1114) );
  XNOR U795 ( .A(n1116), .B(n1102), .Z(n1105) );
  XOR U796 ( .A(n1117), .B(n1118), .Z(n1102) );
  AND U797 ( .A(n1119), .B(n1120), .Z(n1118) );
  XOR U798 ( .A(p_input[1673]), .B(n1117), .Z(n1120) );
  XOR U799 ( .A(n1121), .B(n1122), .Z(n1117) );
  AND U800 ( .A(n1123), .B(n1124), .Z(n1122) );
  IV U801 ( .A(n1113), .Z(n1116) );
  XOR U802 ( .A(n1125), .B(n1126), .Z(n1113) );
  AND U803 ( .A(n1127), .B(n1128), .Z(n1126) );
  XOR U804 ( .A(n1129), .B(n1130), .Z(n1110) );
  AND U805 ( .A(n1131), .B(n1128), .Z(n1130) );
  XNOR U806 ( .A(n1129), .B(n1125), .Z(n1128) );
  XOR U807 ( .A(n1132), .B(n1133), .Z(n1125) );
  AND U808 ( .A(n1134), .B(n1124), .Z(n1133) );
  XNOR U809 ( .A(n1135), .B(n1121), .Z(n1124) );
  XOR U810 ( .A(n1136), .B(n1137), .Z(n1121) );
  AND U811 ( .A(n1138), .B(n1139), .Z(n1137) );
  XOR U812 ( .A(p_input[1705]), .B(n1136), .Z(n1139) );
  XOR U813 ( .A(n1140), .B(n1141), .Z(n1136) );
  AND U814 ( .A(n1142), .B(n1143), .Z(n1141) );
  IV U815 ( .A(n1132), .Z(n1135) );
  XOR U816 ( .A(n1144), .B(n1145), .Z(n1132) );
  AND U817 ( .A(n1146), .B(n1147), .Z(n1145) );
  XOR U818 ( .A(n1148), .B(n1149), .Z(n1129) );
  AND U819 ( .A(n1150), .B(n1147), .Z(n1149) );
  XNOR U820 ( .A(n1148), .B(n1144), .Z(n1147) );
  XOR U821 ( .A(n1151), .B(n1152), .Z(n1144) );
  AND U822 ( .A(n1153), .B(n1143), .Z(n1152) );
  XNOR U823 ( .A(n1154), .B(n1140), .Z(n1143) );
  XOR U824 ( .A(n1155), .B(n1156), .Z(n1140) );
  AND U825 ( .A(n1157), .B(n1158), .Z(n1156) );
  XOR U826 ( .A(p_input[1737]), .B(n1155), .Z(n1158) );
  XOR U827 ( .A(n1159), .B(n1160), .Z(n1155) );
  AND U828 ( .A(n1161), .B(n1162), .Z(n1160) );
  IV U829 ( .A(n1151), .Z(n1154) );
  XOR U830 ( .A(n1163), .B(n1164), .Z(n1151) );
  AND U831 ( .A(n1165), .B(n1166), .Z(n1164) );
  XOR U832 ( .A(n1167), .B(n1168), .Z(n1148) );
  AND U833 ( .A(n1169), .B(n1166), .Z(n1168) );
  XNOR U834 ( .A(n1167), .B(n1163), .Z(n1166) );
  XOR U835 ( .A(n1170), .B(n1171), .Z(n1163) );
  AND U836 ( .A(n1172), .B(n1162), .Z(n1171) );
  XNOR U837 ( .A(n1173), .B(n1159), .Z(n1162) );
  XOR U838 ( .A(n1174), .B(n1175), .Z(n1159) );
  AND U839 ( .A(n1176), .B(n1177), .Z(n1175) );
  XOR U840 ( .A(p_input[1769]), .B(n1174), .Z(n1177) );
  XOR U841 ( .A(n1178), .B(n1179), .Z(n1174) );
  AND U842 ( .A(n1180), .B(n1181), .Z(n1179) );
  IV U843 ( .A(n1170), .Z(n1173) );
  XOR U844 ( .A(n1182), .B(n1183), .Z(n1170) );
  AND U845 ( .A(n1184), .B(n1185), .Z(n1183) );
  XOR U846 ( .A(n1186), .B(n1187), .Z(n1167) );
  AND U847 ( .A(n1188), .B(n1185), .Z(n1187) );
  XNOR U848 ( .A(n1186), .B(n1182), .Z(n1185) );
  XOR U849 ( .A(n1189), .B(n1190), .Z(n1182) );
  AND U850 ( .A(n1191), .B(n1181), .Z(n1190) );
  XNOR U851 ( .A(n1192), .B(n1178), .Z(n1181) );
  XOR U852 ( .A(n1193), .B(n1194), .Z(n1178) );
  AND U853 ( .A(n1195), .B(n1196), .Z(n1194) );
  XOR U854 ( .A(p_input[1801]), .B(n1193), .Z(n1196) );
  XOR U855 ( .A(n1197), .B(n1198), .Z(n1193) );
  AND U856 ( .A(n1199), .B(n1200), .Z(n1198) );
  IV U857 ( .A(n1189), .Z(n1192) );
  XOR U858 ( .A(n1201), .B(n1202), .Z(n1189) );
  AND U859 ( .A(n1203), .B(n1204), .Z(n1202) );
  XOR U860 ( .A(n1205), .B(n1206), .Z(n1186) );
  AND U861 ( .A(n1207), .B(n1204), .Z(n1206) );
  XNOR U862 ( .A(n1205), .B(n1201), .Z(n1204) );
  XOR U863 ( .A(n1208), .B(n1209), .Z(n1201) );
  AND U864 ( .A(n1210), .B(n1200), .Z(n1209) );
  XNOR U865 ( .A(n1211), .B(n1197), .Z(n1200) );
  XOR U866 ( .A(n1212), .B(n1213), .Z(n1197) );
  AND U867 ( .A(n1214), .B(n1215), .Z(n1213) );
  XOR U868 ( .A(p_input[1833]), .B(n1212), .Z(n1215) );
  XOR U869 ( .A(n1216), .B(n1217), .Z(n1212) );
  AND U870 ( .A(n1218), .B(n1219), .Z(n1217) );
  IV U871 ( .A(n1208), .Z(n1211) );
  XOR U872 ( .A(n1220), .B(n1221), .Z(n1208) );
  AND U873 ( .A(n1222), .B(n1223), .Z(n1221) );
  XOR U874 ( .A(n1224), .B(n1225), .Z(n1205) );
  AND U875 ( .A(n1226), .B(n1223), .Z(n1225) );
  XNOR U876 ( .A(n1224), .B(n1220), .Z(n1223) );
  XOR U877 ( .A(n1227), .B(n1228), .Z(n1220) );
  AND U878 ( .A(n1229), .B(n1219), .Z(n1228) );
  XNOR U879 ( .A(n1230), .B(n1216), .Z(n1219) );
  XOR U880 ( .A(n1231), .B(n1232), .Z(n1216) );
  AND U881 ( .A(n1233), .B(n1234), .Z(n1232) );
  XOR U882 ( .A(p_input[1865]), .B(n1231), .Z(n1234) );
  XOR U883 ( .A(n1235), .B(n1236), .Z(n1231) );
  AND U884 ( .A(n1237), .B(n1238), .Z(n1236) );
  IV U885 ( .A(n1227), .Z(n1230) );
  XOR U886 ( .A(n1239), .B(n1240), .Z(n1227) );
  AND U887 ( .A(n1241), .B(n1242), .Z(n1240) );
  XOR U888 ( .A(n1243), .B(n1244), .Z(n1224) );
  AND U889 ( .A(n1245), .B(n1242), .Z(n1244) );
  XNOR U890 ( .A(n1243), .B(n1239), .Z(n1242) );
  XOR U891 ( .A(n1246), .B(n1247), .Z(n1239) );
  AND U892 ( .A(n1248), .B(n1238), .Z(n1247) );
  XNOR U893 ( .A(n1249), .B(n1235), .Z(n1238) );
  XOR U894 ( .A(n1250), .B(n1251), .Z(n1235) );
  AND U895 ( .A(n1252), .B(n1253), .Z(n1251) );
  XOR U896 ( .A(p_input[1897]), .B(n1250), .Z(n1253) );
  XOR U897 ( .A(n1254), .B(n1255), .Z(n1250) );
  AND U898 ( .A(n1256), .B(n1257), .Z(n1255) );
  IV U899 ( .A(n1246), .Z(n1249) );
  XOR U900 ( .A(n1258), .B(n1259), .Z(n1246) );
  AND U901 ( .A(n1260), .B(n1261), .Z(n1259) );
  XOR U902 ( .A(n1262), .B(n1263), .Z(n1243) );
  AND U903 ( .A(n1264), .B(n1261), .Z(n1263) );
  XNOR U904 ( .A(n1262), .B(n1258), .Z(n1261) );
  XOR U905 ( .A(n1265), .B(n1266), .Z(n1258) );
  AND U906 ( .A(n1267), .B(n1257), .Z(n1266) );
  XNOR U907 ( .A(n1268), .B(n1254), .Z(n1257) );
  XOR U908 ( .A(n1269), .B(n1270), .Z(n1254) );
  AND U909 ( .A(n1271), .B(n1272), .Z(n1270) );
  XOR U910 ( .A(p_input[1929]), .B(n1269), .Z(n1272) );
  XOR U911 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(n1273), .Z(
        n1269) );
  AND U912 ( .A(n1274), .B(n1275), .Z(n1273) );
  IV U913 ( .A(n1265), .Z(n1268) );
  XOR U914 ( .A(n1276), .B(n1277), .Z(n1265) );
  AND U915 ( .A(n1278), .B(n1279), .Z(n1277) );
  XOR U916 ( .A(n1280), .B(n1281), .Z(n1262) );
  AND U917 ( .A(n1282), .B(n1279), .Z(n1281) );
  XNOR U918 ( .A(n1280), .B(n1276), .Z(n1279) );
  XNOR U919 ( .A(n1283), .B(n1284), .Z(n1276) );
  AND U920 ( .A(n1285), .B(n1275), .Z(n1284) );
  XNOR U921 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(n1283), 
        .Z(n1275) );
  XNOR U922 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .B(n1286), 
        .Z(n1283) );
  AND U923 ( .A(n1287), .B(n1288), .Z(n1286) );
  XNOR U924 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n1289), .Z(n1280) );
  AND U925 ( .A(n1290), .B(n1288), .Z(n1289) );
  XOR U926 ( .A(n1291), .B(n1292), .Z(n1288) );
  XOR U927 ( .A(n15), .B(n1293), .Z(o[40]) );
  AND U928 ( .A(n122), .B(n1294), .Z(n15) );
  XOR U929 ( .A(n16), .B(n1293), .Z(n1294) );
  XOR U930 ( .A(n1295), .B(n53), .Z(n1293) );
  AND U931 ( .A(n125), .B(n1296), .Z(n53) );
  XNOR U932 ( .A(n1297), .B(n54), .Z(n1296) );
  XOR U933 ( .A(n1298), .B(n1299), .Z(n54) );
  AND U934 ( .A(n130), .B(n1300), .Z(n1299) );
  XOR U935 ( .A(p_input[8]), .B(n1298), .Z(n1300) );
  XOR U936 ( .A(n1301), .B(n1302), .Z(n1298) );
  AND U937 ( .A(n134), .B(n1303), .Z(n1302) );
  IV U938 ( .A(n1295), .Z(n1297) );
  XOR U939 ( .A(n1304), .B(n1305), .Z(n1295) );
  AND U940 ( .A(n138), .B(n1306), .Z(n1305) );
  XOR U941 ( .A(n1307), .B(n1308), .Z(n16) );
  AND U942 ( .A(n142), .B(n1306), .Z(n1308) );
  XNOR U943 ( .A(n1309), .B(n1304), .Z(n1306) );
  XOR U944 ( .A(n1310), .B(n1311), .Z(n1304) );
  AND U945 ( .A(n146), .B(n1303), .Z(n1311) );
  XNOR U946 ( .A(n1312), .B(n1301), .Z(n1303) );
  XOR U947 ( .A(n1313), .B(n1314), .Z(n1301) );
  AND U948 ( .A(n150), .B(n1315), .Z(n1314) );
  XOR U949 ( .A(p_input[40]), .B(n1313), .Z(n1315) );
  XOR U950 ( .A(n1316), .B(n1317), .Z(n1313) );
  AND U951 ( .A(n154), .B(n1318), .Z(n1317) );
  IV U952 ( .A(n1310), .Z(n1312) );
  XOR U953 ( .A(n1319), .B(n1320), .Z(n1310) );
  AND U954 ( .A(n158), .B(n1321), .Z(n1320) );
  IV U955 ( .A(n1307), .Z(n1309) );
  XNOR U956 ( .A(n1322), .B(n1323), .Z(n1307) );
  AND U957 ( .A(n162), .B(n1321), .Z(n1323) );
  XNOR U958 ( .A(n1322), .B(n1319), .Z(n1321) );
  XOR U959 ( .A(n1324), .B(n1325), .Z(n1319) );
  AND U960 ( .A(n165), .B(n1318), .Z(n1325) );
  XNOR U961 ( .A(n1326), .B(n1316), .Z(n1318) );
  XOR U962 ( .A(n1327), .B(n1328), .Z(n1316) );
  AND U963 ( .A(n169), .B(n1329), .Z(n1328) );
  XOR U964 ( .A(p_input[72]), .B(n1327), .Z(n1329) );
  XOR U965 ( .A(n1330), .B(n1331), .Z(n1327) );
  AND U966 ( .A(n173), .B(n1332), .Z(n1331) );
  IV U967 ( .A(n1324), .Z(n1326) );
  XOR U968 ( .A(n1333), .B(n1334), .Z(n1324) );
  AND U969 ( .A(n177), .B(n1335), .Z(n1334) );
  XOR U970 ( .A(n1336), .B(n1337), .Z(n1322) );
  AND U971 ( .A(n181), .B(n1335), .Z(n1337) );
  XNOR U972 ( .A(n1336), .B(n1333), .Z(n1335) );
  XOR U973 ( .A(n1338), .B(n1339), .Z(n1333) );
  AND U974 ( .A(n184), .B(n1332), .Z(n1339) );
  XNOR U975 ( .A(n1340), .B(n1330), .Z(n1332) );
  XOR U976 ( .A(n1341), .B(n1342), .Z(n1330) );
  AND U977 ( .A(n188), .B(n1343), .Z(n1342) );
  XOR U978 ( .A(p_input[104]), .B(n1341), .Z(n1343) );
  XOR U979 ( .A(n1344), .B(n1345), .Z(n1341) );
  AND U980 ( .A(n192), .B(n1346), .Z(n1345) );
  IV U981 ( .A(n1338), .Z(n1340) );
  XOR U982 ( .A(n1347), .B(n1348), .Z(n1338) );
  AND U983 ( .A(n196), .B(n1349), .Z(n1348) );
  XOR U984 ( .A(n1350), .B(n1351), .Z(n1336) );
  AND U985 ( .A(n200), .B(n1349), .Z(n1351) );
  XNOR U986 ( .A(n1350), .B(n1347), .Z(n1349) );
  XOR U987 ( .A(n1352), .B(n1353), .Z(n1347) );
  AND U988 ( .A(n203), .B(n1346), .Z(n1353) );
  XNOR U989 ( .A(n1354), .B(n1344), .Z(n1346) );
  XOR U990 ( .A(n1355), .B(n1356), .Z(n1344) );
  AND U991 ( .A(n207), .B(n1357), .Z(n1356) );
  XOR U992 ( .A(p_input[136]), .B(n1355), .Z(n1357) );
  XOR U993 ( .A(n1358), .B(n1359), .Z(n1355) );
  AND U994 ( .A(n211), .B(n1360), .Z(n1359) );
  IV U995 ( .A(n1352), .Z(n1354) );
  XOR U996 ( .A(n1361), .B(n1362), .Z(n1352) );
  AND U997 ( .A(n215), .B(n1363), .Z(n1362) );
  XOR U998 ( .A(n1364), .B(n1365), .Z(n1350) );
  AND U999 ( .A(n219), .B(n1363), .Z(n1365) );
  XNOR U1000 ( .A(n1364), .B(n1361), .Z(n1363) );
  XOR U1001 ( .A(n1366), .B(n1367), .Z(n1361) );
  AND U1002 ( .A(n222), .B(n1360), .Z(n1367) );
  XNOR U1003 ( .A(n1368), .B(n1358), .Z(n1360) );
  XOR U1004 ( .A(n1369), .B(n1370), .Z(n1358) );
  AND U1005 ( .A(n226), .B(n1371), .Z(n1370) );
  XOR U1006 ( .A(p_input[168]), .B(n1369), .Z(n1371) );
  XOR U1007 ( .A(n1372), .B(n1373), .Z(n1369) );
  AND U1008 ( .A(n230), .B(n1374), .Z(n1373) );
  IV U1009 ( .A(n1366), .Z(n1368) );
  XOR U1010 ( .A(n1375), .B(n1376), .Z(n1366) );
  AND U1011 ( .A(n234), .B(n1377), .Z(n1376) );
  XOR U1012 ( .A(n1378), .B(n1379), .Z(n1364) );
  AND U1013 ( .A(n238), .B(n1377), .Z(n1379) );
  XNOR U1014 ( .A(n1378), .B(n1375), .Z(n1377) );
  XOR U1015 ( .A(n1380), .B(n1381), .Z(n1375) );
  AND U1016 ( .A(n241), .B(n1374), .Z(n1381) );
  XNOR U1017 ( .A(n1382), .B(n1372), .Z(n1374) );
  XOR U1018 ( .A(n1383), .B(n1384), .Z(n1372) );
  AND U1019 ( .A(n245), .B(n1385), .Z(n1384) );
  XOR U1020 ( .A(p_input[200]), .B(n1383), .Z(n1385) );
  XOR U1021 ( .A(n1386), .B(n1387), .Z(n1383) );
  AND U1022 ( .A(n249), .B(n1388), .Z(n1387) );
  IV U1023 ( .A(n1380), .Z(n1382) );
  XOR U1024 ( .A(n1389), .B(n1390), .Z(n1380) );
  AND U1025 ( .A(n253), .B(n1391), .Z(n1390) );
  XOR U1026 ( .A(n1392), .B(n1393), .Z(n1378) );
  AND U1027 ( .A(n257), .B(n1391), .Z(n1393) );
  XNOR U1028 ( .A(n1392), .B(n1389), .Z(n1391) );
  XOR U1029 ( .A(n1394), .B(n1395), .Z(n1389) );
  AND U1030 ( .A(n260), .B(n1388), .Z(n1395) );
  XNOR U1031 ( .A(n1396), .B(n1386), .Z(n1388) );
  XOR U1032 ( .A(n1397), .B(n1398), .Z(n1386) );
  AND U1033 ( .A(n264), .B(n1399), .Z(n1398) );
  XOR U1034 ( .A(p_input[232]), .B(n1397), .Z(n1399) );
  XOR U1035 ( .A(n1400), .B(n1401), .Z(n1397) );
  AND U1036 ( .A(n268), .B(n1402), .Z(n1401) );
  IV U1037 ( .A(n1394), .Z(n1396) );
  XOR U1038 ( .A(n1403), .B(n1404), .Z(n1394) );
  AND U1039 ( .A(n272), .B(n1405), .Z(n1404) );
  XOR U1040 ( .A(n1406), .B(n1407), .Z(n1392) );
  AND U1041 ( .A(n276), .B(n1405), .Z(n1407) );
  XNOR U1042 ( .A(n1406), .B(n1403), .Z(n1405) );
  XOR U1043 ( .A(n1408), .B(n1409), .Z(n1403) );
  AND U1044 ( .A(n279), .B(n1402), .Z(n1409) );
  XNOR U1045 ( .A(n1410), .B(n1400), .Z(n1402) );
  XOR U1046 ( .A(n1411), .B(n1412), .Z(n1400) );
  AND U1047 ( .A(n283), .B(n1413), .Z(n1412) );
  XOR U1048 ( .A(p_input[264]), .B(n1411), .Z(n1413) );
  XOR U1049 ( .A(n1414), .B(n1415), .Z(n1411) );
  AND U1050 ( .A(n287), .B(n1416), .Z(n1415) );
  IV U1051 ( .A(n1408), .Z(n1410) );
  XOR U1052 ( .A(n1417), .B(n1418), .Z(n1408) );
  AND U1053 ( .A(n291), .B(n1419), .Z(n1418) );
  XOR U1054 ( .A(n1420), .B(n1421), .Z(n1406) );
  AND U1055 ( .A(n295), .B(n1419), .Z(n1421) );
  XNOR U1056 ( .A(n1420), .B(n1417), .Z(n1419) );
  XOR U1057 ( .A(n1422), .B(n1423), .Z(n1417) );
  AND U1058 ( .A(n298), .B(n1416), .Z(n1423) );
  XNOR U1059 ( .A(n1424), .B(n1414), .Z(n1416) );
  XOR U1060 ( .A(n1425), .B(n1426), .Z(n1414) );
  AND U1061 ( .A(n302), .B(n1427), .Z(n1426) );
  XOR U1062 ( .A(p_input[296]), .B(n1425), .Z(n1427) );
  XOR U1063 ( .A(n1428), .B(n1429), .Z(n1425) );
  AND U1064 ( .A(n306), .B(n1430), .Z(n1429) );
  IV U1065 ( .A(n1422), .Z(n1424) );
  XOR U1066 ( .A(n1431), .B(n1432), .Z(n1422) );
  AND U1067 ( .A(n310), .B(n1433), .Z(n1432) );
  XOR U1068 ( .A(n1434), .B(n1435), .Z(n1420) );
  AND U1069 ( .A(n314), .B(n1433), .Z(n1435) );
  XNOR U1070 ( .A(n1434), .B(n1431), .Z(n1433) );
  XOR U1071 ( .A(n1436), .B(n1437), .Z(n1431) );
  AND U1072 ( .A(n317), .B(n1430), .Z(n1437) );
  XNOR U1073 ( .A(n1438), .B(n1428), .Z(n1430) );
  XOR U1074 ( .A(n1439), .B(n1440), .Z(n1428) );
  AND U1075 ( .A(n321), .B(n1441), .Z(n1440) );
  XOR U1076 ( .A(p_input[328]), .B(n1439), .Z(n1441) );
  XOR U1077 ( .A(n1442), .B(n1443), .Z(n1439) );
  AND U1078 ( .A(n325), .B(n1444), .Z(n1443) );
  IV U1079 ( .A(n1436), .Z(n1438) );
  XOR U1080 ( .A(n1445), .B(n1446), .Z(n1436) );
  AND U1081 ( .A(n329), .B(n1447), .Z(n1446) );
  XOR U1082 ( .A(n1448), .B(n1449), .Z(n1434) );
  AND U1083 ( .A(n333), .B(n1447), .Z(n1449) );
  XNOR U1084 ( .A(n1448), .B(n1445), .Z(n1447) );
  XOR U1085 ( .A(n1450), .B(n1451), .Z(n1445) );
  AND U1086 ( .A(n336), .B(n1444), .Z(n1451) );
  XNOR U1087 ( .A(n1452), .B(n1442), .Z(n1444) );
  XOR U1088 ( .A(n1453), .B(n1454), .Z(n1442) );
  AND U1089 ( .A(n340), .B(n1455), .Z(n1454) );
  XOR U1090 ( .A(p_input[360]), .B(n1453), .Z(n1455) );
  XOR U1091 ( .A(n1456), .B(n1457), .Z(n1453) );
  AND U1092 ( .A(n344), .B(n1458), .Z(n1457) );
  IV U1093 ( .A(n1450), .Z(n1452) );
  XOR U1094 ( .A(n1459), .B(n1460), .Z(n1450) );
  AND U1095 ( .A(n348), .B(n1461), .Z(n1460) );
  XOR U1096 ( .A(n1462), .B(n1463), .Z(n1448) );
  AND U1097 ( .A(n352), .B(n1461), .Z(n1463) );
  XNOR U1098 ( .A(n1462), .B(n1459), .Z(n1461) );
  XOR U1099 ( .A(n1464), .B(n1465), .Z(n1459) );
  AND U1100 ( .A(n355), .B(n1458), .Z(n1465) );
  XNOR U1101 ( .A(n1466), .B(n1456), .Z(n1458) );
  XOR U1102 ( .A(n1467), .B(n1468), .Z(n1456) );
  AND U1103 ( .A(n359), .B(n1469), .Z(n1468) );
  XOR U1104 ( .A(p_input[392]), .B(n1467), .Z(n1469) );
  XOR U1105 ( .A(n1470), .B(n1471), .Z(n1467) );
  AND U1106 ( .A(n363), .B(n1472), .Z(n1471) );
  IV U1107 ( .A(n1464), .Z(n1466) );
  XOR U1108 ( .A(n1473), .B(n1474), .Z(n1464) );
  AND U1109 ( .A(n367), .B(n1475), .Z(n1474) );
  XOR U1110 ( .A(n1476), .B(n1477), .Z(n1462) );
  AND U1111 ( .A(n371), .B(n1475), .Z(n1477) );
  XNOR U1112 ( .A(n1476), .B(n1473), .Z(n1475) );
  XOR U1113 ( .A(n1478), .B(n1479), .Z(n1473) );
  AND U1114 ( .A(n374), .B(n1472), .Z(n1479) );
  XNOR U1115 ( .A(n1480), .B(n1470), .Z(n1472) );
  XOR U1116 ( .A(n1481), .B(n1482), .Z(n1470) );
  AND U1117 ( .A(n378), .B(n1483), .Z(n1482) );
  XOR U1118 ( .A(p_input[424]), .B(n1481), .Z(n1483) );
  XOR U1119 ( .A(n1484), .B(n1485), .Z(n1481) );
  AND U1120 ( .A(n382), .B(n1486), .Z(n1485) );
  IV U1121 ( .A(n1478), .Z(n1480) );
  XOR U1122 ( .A(n1487), .B(n1488), .Z(n1478) );
  AND U1123 ( .A(n386), .B(n1489), .Z(n1488) );
  XOR U1124 ( .A(n1490), .B(n1491), .Z(n1476) );
  AND U1125 ( .A(n390), .B(n1489), .Z(n1491) );
  XNOR U1126 ( .A(n1490), .B(n1487), .Z(n1489) );
  XOR U1127 ( .A(n1492), .B(n1493), .Z(n1487) );
  AND U1128 ( .A(n393), .B(n1486), .Z(n1493) );
  XNOR U1129 ( .A(n1494), .B(n1484), .Z(n1486) );
  XOR U1130 ( .A(n1495), .B(n1496), .Z(n1484) );
  AND U1131 ( .A(n397), .B(n1497), .Z(n1496) );
  XOR U1132 ( .A(p_input[456]), .B(n1495), .Z(n1497) );
  XOR U1133 ( .A(n1498), .B(n1499), .Z(n1495) );
  AND U1134 ( .A(n401), .B(n1500), .Z(n1499) );
  IV U1135 ( .A(n1492), .Z(n1494) );
  XOR U1136 ( .A(n1501), .B(n1502), .Z(n1492) );
  AND U1137 ( .A(n405), .B(n1503), .Z(n1502) );
  XOR U1138 ( .A(n1504), .B(n1505), .Z(n1490) );
  AND U1139 ( .A(n409), .B(n1503), .Z(n1505) );
  XNOR U1140 ( .A(n1504), .B(n1501), .Z(n1503) );
  XOR U1141 ( .A(n1506), .B(n1507), .Z(n1501) );
  AND U1142 ( .A(n412), .B(n1500), .Z(n1507) );
  XNOR U1143 ( .A(n1508), .B(n1498), .Z(n1500) );
  XOR U1144 ( .A(n1509), .B(n1510), .Z(n1498) );
  AND U1145 ( .A(n416), .B(n1511), .Z(n1510) );
  XOR U1146 ( .A(p_input[488]), .B(n1509), .Z(n1511) );
  XOR U1147 ( .A(n1512), .B(n1513), .Z(n1509) );
  AND U1148 ( .A(n420), .B(n1514), .Z(n1513) );
  IV U1149 ( .A(n1506), .Z(n1508) );
  XOR U1150 ( .A(n1515), .B(n1516), .Z(n1506) );
  AND U1151 ( .A(n424), .B(n1517), .Z(n1516) );
  XOR U1152 ( .A(n1518), .B(n1519), .Z(n1504) );
  AND U1153 ( .A(n428), .B(n1517), .Z(n1519) );
  XNOR U1154 ( .A(n1518), .B(n1515), .Z(n1517) );
  XOR U1155 ( .A(n1520), .B(n1521), .Z(n1515) );
  AND U1156 ( .A(n431), .B(n1514), .Z(n1521) );
  XNOR U1157 ( .A(n1522), .B(n1512), .Z(n1514) );
  XOR U1158 ( .A(n1523), .B(n1524), .Z(n1512) );
  AND U1159 ( .A(n435), .B(n1525), .Z(n1524) );
  XOR U1160 ( .A(p_input[520]), .B(n1523), .Z(n1525) );
  XOR U1161 ( .A(n1526), .B(n1527), .Z(n1523) );
  AND U1162 ( .A(n439), .B(n1528), .Z(n1527) );
  IV U1163 ( .A(n1520), .Z(n1522) );
  XOR U1164 ( .A(n1529), .B(n1530), .Z(n1520) );
  AND U1165 ( .A(n443), .B(n1531), .Z(n1530) );
  XOR U1166 ( .A(n1532), .B(n1533), .Z(n1518) );
  AND U1167 ( .A(n447), .B(n1531), .Z(n1533) );
  XNOR U1168 ( .A(n1532), .B(n1529), .Z(n1531) );
  XOR U1169 ( .A(n1534), .B(n1535), .Z(n1529) );
  AND U1170 ( .A(n450), .B(n1528), .Z(n1535) );
  XNOR U1171 ( .A(n1536), .B(n1526), .Z(n1528) );
  XOR U1172 ( .A(n1537), .B(n1538), .Z(n1526) );
  AND U1173 ( .A(n454), .B(n1539), .Z(n1538) );
  XOR U1174 ( .A(p_input[552]), .B(n1537), .Z(n1539) );
  XOR U1175 ( .A(n1540), .B(n1541), .Z(n1537) );
  AND U1176 ( .A(n458), .B(n1542), .Z(n1541) );
  IV U1177 ( .A(n1534), .Z(n1536) );
  XOR U1178 ( .A(n1543), .B(n1544), .Z(n1534) );
  AND U1179 ( .A(n462), .B(n1545), .Z(n1544) );
  XOR U1180 ( .A(n1546), .B(n1547), .Z(n1532) );
  AND U1181 ( .A(n466), .B(n1545), .Z(n1547) );
  XNOR U1182 ( .A(n1546), .B(n1543), .Z(n1545) );
  XOR U1183 ( .A(n1548), .B(n1549), .Z(n1543) );
  AND U1184 ( .A(n469), .B(n1542), .Z(n1549) );
  XNOR U1185 ( .A(n1550), .B(n1540), .Z(n1542) );
  XOR U1186 ( .A(n1551), .B(n1552), .Z(n1540) );
  AND U1187 ( .A(n473), .B(n1553), .Z(n1552) );
  XOR U1188 ( .A(p_input[584]), .B(n1551), .Z(n1553) );
  XOR U1189 ( .A(n1554), .B(n1555), .Z(n1551) );
  AND U1190 ( .A(n477), .B(n1556), .Z(n1555) );
  IV U1191 ( .A(n1548), .Z(n1550) );
  XOR U1192 ( .A(n1557), .B(n1558), .Z(n1548) );
  AND U1193 ( .A(n481), .B(n1559), .Z(n1558) );
  XOR U1194 ( .A(n1560), .B(n1561), .Z(n1546) );
  AND U1195 ( .A(n485), .B(n1559), .Z(n1561) );
  XNOR U1196 ( .A(n1560), .B(n1557), .Z(n1559) );
  XOR U1197 ( .A(n1562), .B(n1563), .Z(n1557) );
  AND U1198 ( .A(n488), .B(n1556), .Z(n1563) );
  XNOR U1199 ( .A(n1564), .B(n1554), .Z(n1556) );
  XOR U1200 ( .A(n1565), .B(n1566), .Z(n1554) );
  AND U1201 ( .A(n492), .B(n1567), .Z(n1566) );
  XOR U1202 ( .A(p_input[616]), .B(n1565), .Z(n1567) );
  XOR U1203 ( .A(n1568), .B(n1569), .Z(n1565) );
  AND U1204 ( .A(n496), .B(n1570), .Z(n1569) );
  IV U1205 ( .A(n1562), .Z(n1564) );
  XOR U1206 ( .A(n1571), .B(n1572), .Z(n1562) );
  AND U1207 ( .A(n500), .B(n1573), .Z(n1572) );
  XOR U1208 ( .A(n1574), .B(n1575), .Z(n1560) );
  AND U1209 ( .A(n504), .B(n1573), .Z(n1575) );
  XNOR U1210 ( .A(n1574), .B(n1571), .Z(n1573) );
  XOR U1211 ( .A(n1576), .B(n1577), .Z(n1571) );
  AND U1212 ( .A(n507), .B(n1570), .Z(n1577) );
  XNOR U1213 ( .A(n1578), .B(n1568), .Z(n1570) );
  XOR U1214 ( .A(n1579), .B(n1580), .Z(n1568) );
  AND U1215 ( .A(n511), .B(n1581), .Z(n1580) );
  XOR U1216 ( .A(p_input[648]), .B(n1579), .Z(n1581) );
  XOR U1217 ( .A(n1582), .B(n1583), .Z(n1579) );
  AND U1218 ( .A(n515), .B(n1584), .Z(n1583) );
  IV U1219 ( .A(n1576), .Z(n1578) );
  XOR U1220 ( .A(n1585), .B(n1586), .Z(n1576) );
  AND U1221 ( .A(n519), .B(n1587), .Z(n1586) );
  XOR U1222 ( .A(n1588), .B(n1589), .Z(n1574) );
  AND U1223 ( .A(n523), .B(n1587), .Z(n1589) );
  XNOR U1224 ( .A(n1588), .B(n1585), .Z(n1587) );
  XOR U1225 ( .A(n1590), .B(n1591), .Z(n1585) );
  AND U1226 ( .A(n526), .B(n1584), .Z(n1591) );
  XNOR U1227 ( .A(n1592), .B(n1582), .Z(n1584) );
  XOR U1228 ( .A(n1593), .B(n1594), .Z(n1582) );
  AND U1229 ( .A(n530), .B(n1595), .Z(n1594) );
  XOR U1230 ( .A(p_input[680]), .B(n1593), .Z(n1595) );
  XOR U1231 ( .A(n1596), .B(n1597), .Z(n1593) );
  AND U1232 ( .A(n534), .B(n1598), .Z(n1597) );
  IV U1233 ( .A(n1590), .Z(n1592) );
  XOR U1234 ( .A(n1599), .B(n1600), .Z(n1590) );
  AND U1235 ( .A(n538), .B(n1601), .Z(n1600) );
  XOR U1236 ( .A(n1602), .B(n1603), .Z(n1588) );
  AND U1237 ( .A(n542), .B(n1601), .Z(n1603) );
  XNOR U1238 ( .A(n1602), .B(n1599), .Z(n1601) );
  XOR U1239 ( .A(n1604), .B(n1605), .Z(n1599) );
  AND U1240 ( .A(n545), .B(n1598), .Z(n1605) );
  XNOR U1241 ( .A(n1606), .B(n1596), .Z(n1598) );
  XOR U1242 ( .A(n1607), .B(n1608), .Z(n1596) );
  AND U1243 ( .A(n549), .B(n1609), .Z(n1608) );
  XOR U1244 ( .A(p_input[712]), .B(n1607), .Z(n1609) );
  XOR U1245 ( .A(n1610), .B(n1611), .Z(n1607) );
  AND U1246 ( .A(n553), .B(n1612), .Z(n1611) );
  IV U1247 ( .A(n1604), .Z(n1606) );
  XOR U1248 ( .A(n1613), .B(n1614), .Z(n1604) );
  AND U1249 ( .A(n557), .B(n1615), .Z(n1614) );
  XOR U1250 ( .A(n1616), .B(n1617), .Z(n1602) );
  AND U1251 ( .A(n561), .B(n1615), .Z(n1617) );
  XNOR U1252 ( .A(n1616), .B(n1613), .Z(n1615) );
  XOR U1253 ( .A(n1618), .B(n1619), .Z(n1613) );
  AND U1254 ( .A(n564), .B(n1612), .Z(n1619) );
  XNOR U1255 ( .A(n1620), .B(n1610), .Z(n1612) );
  XOR U1256 ( .A(n1621), .B(n1622), .Z(n1610) );
  AND U1257 ( .A(n568), .B(n1623), .Z(n1622) );
  XOR U1258 ( .A(p_input[744]), .B(n1621), .Z(n1623) );
  XOR U1259 ( .A(n1624), .B(n1625), .Z(n1621) );
  AND U1260 ( .A(n572), .B(n1626), .Z(n1625) );
  IV U1261 ( .A(n1618), .Z(n1620) );
  XOR U1262 ( .A(n1627), .B(n1628), .Z(n1618) );
  AND U1263 ( .A(n576), .B(n1629), .Z(n1628) );
  XOR U1264 ( .A(n1630), .B(n1631), .Z(n1616) );
  AND U1265 ( .A(n580), .B(n1629), .Z(n1631) );
  XNOR U1266 ( .A(n1630), .B(n1627), .Z(n1629) );
  XOR U1267 ( .A(n1632), .B(n1633), .Z(n1627) );
  AND U1268 ( .A(n583), .B(n1626), .Z(n1633) );
  XNOR U1269 ( .A(n1634), .B(n1624), .Z(n1626) );
  XOR U1270 ( .A(n1635), .B(n1636), .Z(n1624) );
  AND U1271 ( .A(n587), .B(n1637), .Z(n1636) );
  XOR U1272 ( .A(p_input[776]), .B(n1635), .Z(n1637) );
  XOR U1273 ( .A(n1638), .B(n1639), .Z(n1635) );
  AND U1274 ( .A(n591), .B(n1640), .Z(n1639) );
  IV U1275 ( .A(n1632), .Z(n1634) );
  XOR U1276 ( .A(n1641), .B(n1642), .Z(n1632) );
  AND U1277 ( .A(n595), .B(n1643), .Z(n1642) );
  XOR U1278 ( .A(n1644), .B(n1645), .Z(n1630) );
  AND U1279 ( .A(n599), .B(n1643), .Z(n1645) );
  XNOR U1280 ( .A(n1644), .B(n1641), .Z(n1643) );
  XOR U1281 ( .A(n1646), .B(n1647), .Z(n1641) );
  AND U1282 ( .A(n602), .B(n1640), .Z(n1647) );
  XNOR U1283 ( .A(n1648), .B(n1638), .Z(n1640) );
  XOR U1284 ( .A(n1649), .B(n1650), .Z(n1638) );
  AND U1285 ( .A(n606), .B(n1651), .Z(n1650) );
  XOR U1286 ( .A(p_input[808]), .B(n1649), .Z(n1651) );
  XOR U1287 ( .A(n1652), .B(n1653), .Z(n1649) );
  AND U1288 ( .A(n610), .B(n1654), .Z(n1653) );
  IV U1289 ( .A(n1646), .Z(n1648) );
  XOR U1290 ( .A(n1655), .B(n1656), .Z(n1646) );
  AND U1291 ( .A(n614), .B(n1657), .Z(n1656) );
  XOR U1292 ( .A(n1658), .B(n1659), .Z(n1644) );
  AND U1293 ( .A(n618), .B(n1657), .Z(n1659) );
  XNOR U1294 ( .A(n1658), .B(n1655), .Z(n1657) );
  XOR U1295 ( .A(n1660), .B(n1661), .Z(n1655) );
  AND U1296 ( .A(n621), .B(n1654), .Z(n1661) );
  XNOR U1297 ( .A(n1662), .B(n1652), .Z(n1654) );
  XOR U1298 ( .A(n1663), .B(n1664), .Z(n1652) );
  AND U1299 ( .A(n625), .B(n1665), .Z(n1664) );
  XOR U1300 ( .A(p_input[840]), .B(n1663), .Z(n1665) );
  XOR U1301 ( .A(n1666), .B(n1667), .Z(n1663) );
  AND U1302 ( .A(n629), .B(n1668), .Z(n1667) );
  IV U1303 ( .A(n1660), .Z(n1662) );
  XOR U1304 ( .A(n1669), .B(n1670), .Z(n1660) );
  AND U1305 ( .A(n633), .B(n1671), .Z(n1670) );
  XOR U1306 ( .A(n1672), .B(n1673), .Z(n1658) );
  AND U1307 ( .A(n637), .B(n1671), .Z(n1673) );
  XNOR U1308 ( .A(n1672), .B(n1669), .Z(n1671) );
  XOR U1309 ( .A(n1674), .B(n1675), .Z(n1669) );
  AND U1310 ( .A(n640), .B(n1668), .Z(n1675) );
  XNOR U1311 ( .A(n1676), .B(n1666), .Z(n1668) );
  XOR U1312 ( .A(n1677), .B(n1678), .Z(n1666) );
  AND U1313 ( .A(n644), .B(n1679), .Z(n1678) );
  XOR U1314 ( .A(p_input[872]), .B(n1677), .Z(n1679) );
  XOR U1315 ( .A(n1680), .B(n1681), .Z(n1677) );
  AND U1316 ( .A(n648), .B(n1682), .Z(n1681) );
  IV U1317 ( .A(n1674), .Z(n1676) );
  XOR U1318 ( .A(n1683), .B(n1684), .Z(n1674) );
  AND U1319 ( .A(n652), .B(n1685), .Z(n1684) );
  XOR U1320 ( .A(n1686), .B(n1687), .Z(n1672) );
  AND U1321 ( .A(n656), .B(n1685), .Z(n1687) );
  XNOR U1322 ( .A(n1686), .B(n1683), .Z(n1685) );
  XOR U1323 ( .A(n1688), .B(n1689), .Z(n1683) );
  AND U1324 ( .A(n659), .B(n1682), .Z(n1689) );
  XNOR U1325 ( .A(n1690), .B(n1680), .Z(n1682) );
  XOR U1326 ( .A(n1691), .B(n1692), .Z(n1680) );
  AND U1327 ( .A(n663), .B(n1693), .Z(n1692) );
  XOR U1328 ( .A(p_input[904]), .B(n1691), .Z(n1693) );
  XOR U1329 ( .A(n1694), .B(n1695), .Z(n1691) );
  AND U1330 ( .A(n667), .B(n1696), .Z(n1695) );
  IV U1331 ( .A(n1688), .Z(n1690) );
  XOR U1332 ( .A(n1697), .B(n1698), .Z(n1688) );
  AND U1333 ( .A(n671), .B(n1699), .Z(n1698) );
  XOR U1334 ( .A(n1700), .B(n1701), .Z(n1686) );
  AND U1335 ( .A(n675), .B(n1699), .Z(n1701) );
  XNOR U1336 ( .A(n1700), .B(n1697), .Z(n1699) );
  XOR U1337 ( .A(n1702), .B(n1703), .Z(n1697) );
  AND U1338 ( .A(n678), .B(n1696), .Z(n1703) );
  XNOR U1339 ( .A(n1704), .B(n1694), .Z(n1696) );
  XOR U1340 ( .A(n1705), .B(n1706), .Z(n1694) );
  AND U1341 ( .A(n682), .B(n1707), .Z(n1706) );
  XOR U1342 ( .A(p_input[936]), .B(n1705), .Z(n1707) );
  XOR U1343 ( .A(n1708), .B(n1709), .Z(n1705) );
  AND U1344 ( .A(n686), .B(n1710), .Z(n1709) );
  IV U1345 ( .A(n1702), .Z(n1704) );
  XOR U1346 ( .A(n1711), .B(n1712), .Z(n1702) );
  AND U1347 ( .A(n690), .B(n1713), .Z(n1712) );
  XOR U1348 ( .A(n1714), .B(n1715), .Z(n1700) );
  AND U1349 ( .A(n694), .B(n1713), .Z(n1715) );
  XNOR U1350 ( .A(n1714), .B(n1711), .Z(n1713) );
  XOR U1351 ( .A(n1716), .B(n1717), .Z(n1711) );
  AND U1352 ( .A(n697), .B(n1710), .Z(n1717) );
  XNOR U1353 ( .A(n1718), .B(n1708), .Z(n1710) );
  XOR U1354 ( .A(n1719), .B(n1720), .Z(n1708) );
  AND U1355 ( .A(n701), .B(n1721), .Z(n1720) );
  XOR U1356 ( .A(p_input[968]), .B(n1719), .Z(n1721) );
  XOR U1357 ( .A(n1722), .B(n1723), .Z(n1719) );
  AND U1358 ( .A(n705), .B(n1724), .Z(n1723) );
  IV U1359 ( .A(n1716), .Z(n1718) );
  XOR U1360 ( .A(n1725), .B(n1726), .Z(n1716) );
  AND U1361 ( .A(n709), .B(n1727), .Z(n1726) );
  XOR U1362 ( .A(n1728), .B(n1729), .Z(n1714) );
  AND U1363 ( .A(n713), .B(n1727), .Z(n1729) );
  XNOR U1364 ( .A(n1728), .B(n1725), .Z(n1727) );
  XOR U1365 ( .A(n1730), .B(n1731), .Z(n1725) );
  AND U1366 ( .A(n716), .B(n1724), .Z(n1731) );
  XNOR U1367 ( .A(n1732), .B(n1722), .Z(n1724) );
  XOR U1368 ( .A(n1733), .B(n1734), .Z(n1722) );
  AND U1369 ( .A(n720), .B(n1735), .Z(n1734) );
  XOR U1370 ( .A(p_input[1000]), .B(n1733), .Z(n1735) );
  XOR U1371 ( .A(n1736), .B(n1737), .Z(n1733) );
  AND U1372 ( .A(n724), .B(n1738), .Z(n1737) );
  IV U1373 ( .A(n1730), .Z(n1732) );
  XOR U1374 ( .A(n1739), .B(n1740), .Z(n1730) );
  AND U1375 ( .A(n728), .B(n1741), .Z(n1740) );
  XOR U1376 ( .A(n1742), .B(n1743), .Z(n1728) );
  AND U1377 ( .A(n732), .B(n1741), .Z(n1743) );
  XNOR U1378 ( .A(n1742), .B(n1739), .Z(n1741) );
  XOR U1379 ( .A(n1744), .B(n1745), .Z(n1739) );
  AND U1380 ( .A(n735), .B(n1738), .Z(n1745) );
  XNOR U1381 ( .A(n1746), .B(n1736), .Z(n1738) );
  XOR U1382 ( .A(n1747), .B(n1748), .Z(n1736) );
  AND U1383 ( .A(n739), .B(n1749), .Z(n1748) );
  XOR U1384 ( .A(p_input[1032]), .B(n1747), .Z(n1749) );
  XOR U1385 ( .A(n1750), .B(n1751), .Z(n1747) );
  AND U1386 ( .A(n743), .B(n1752), .Z(n1751) );
  IV U1387 ( .A(n1744), .Z(n1746) );
  XOR U1388 ( .A(n1753), .B(n1754), .Z(n1744) );
  AND U1389 ( .A(n747), .B(n1755), .Z(n1754) );
  XOR U1390 ( .A(n1756), .B(n1757), .Z(n1742) );
  AND U1391 ( .A(n751), .B(n1755), .Z(n1757) );
  XNOR U1392 ( .A(n1756), .B(n1753), .Z(n1755) );
  XOR U1393 ( .A(n1758), .B(n1759), .Z(n1753) );
  AND U1394 ( .A(n754), .B(n1752), .Z(n1759) );
  XNOR U1395 ( .A(n1760), .B(n1750), .Z(n1752) );
  XOR U1396 ( .A(n1761), .B(n1762), .Z(n1750) );
  AND U1397 ( .A(n758), .B(n1763), .Z(n1762) );
  XOR U1398 ( .A(p_input[1064]), .B(n1761), .Z(n1763) );
  XOR U1399 ( .A(n1764), .B(n1765), .Z(n1761) );
  AND U1400 ( .A(n762), .B(n1766), .Z(n1765) );
  IV U1401 ( .A(n1758), .Z(n1760) );
  XOR U1402 ( .A(n1767), .B(n1768), .Z(n1758) );
  AND U1403 ( .A(n766), .B(n1769), .Z(n1768) );
  XOR U1404 ( .A(n1770), .B(n1771), .Z(n1756) );
  AND U1405 ( .A(n770), .B(n1769), .Z(n1771) );
  XNOR U1406 ( .A(n1770), .B(n1767), .Z(n1769) );
  XOR U1407 ( .A(n1772), .B(n1773), .Z(n1767) );
  AND U1408 ( .A(n773), .B(n1766), .Z(n1773) );
  XNOR U1409 ( .A(n1774), .B(n1764), .Z(n1766) );
  XOR U1410 ( .A(n1775), .B(n1776), .Z(n1764) );
  AND U1411 ( .A(n777), .B(n1777), .Z(n1776) );
  XOR U1412 ( .A(p_input[1096]), .B(n1775), .Z(n1777) );
  XOR U1413 ( .A(n1778), .B(n1779), .Z(n1775) );
  AND U1414 ( .A(n781), .B(n1780), .Z(n1779) );
  IV U1415 ( .A(n1772), .Z(n1774) );
  XOR U1416 ( .A(n1781), .B(n1782), .Z(n1772) );
  AND U1417 ( .A(n785), .B(n1783), .Z(n1782) );
  XOR U1418 ( .A(n1784), .B(n1785), .Z(n1770) );
  AND U1419 ( .A(n789), .B(n1783), .Z(n1785) );
  XNOR U1420 ( .A(n1784), .B(n1781), .Z(n1783) );
  XOR U1421 ( .A(n1786), .B(n1787), .Z(n1781) );
  AND U1422 ( .A(n792), .B(n1780), .Z(n1787) );
  XNOR U1423 ( .A(n1788), .B(n1778), .Z(n1780) );
  XOR U1424 ( .A(n1789), .B(n1790), .Z(n1778) );
  AND U1425 ( .A(n796), .B(n1791), .Z(n1790) );
  XOR U1426 ( .A(p_input[1128]), .B(n1789), .Z(n1791) );
  XOR U1427 ( .A(n1792), .B(n1793), .Z(n1789) );
  AND U1428 ( .A(n800), .B(n1794), .Z(n1793) );
  IV U1429 ( .A(n1786), .Z(n1788) );
  XOR U1430 ( .A(n1795), .B(n1796), .Z(n1786) );
  AND U1431 ( .A(n804), .B(n1797), .Z(n1796) );
  XOR U1432 ( .A(n1798), .B(n1799), .Z(n1784) );
  AND U1433 ( .A(n808), .B(n1797), .Z(n1799) );
  XNOR U1434 ( .A(n1798), .B(n1795), .Z(n1797) );
  XOR U1435 ( .A(n1800), .B(n1801), .Z(n1795) );
  AND U1436 ( .A(n811), .B(n1794), .Z(n1801) );
  XNOR U1437 ( .A(n1802), .B(n1792), .Z(n1794) );
  XOR U1438 ( .A(n1803), .B(n1804), .Z(n1792) );
  AND U1439 ( .A(n815), .B(n1805), .Z(n1804) );
  XOR U1440 ( .A(p_input[1160]), .B(n1803), .Z(n1805) );
  XOR U1441 ( .A(n1806), .B(n1807), .Z(n1803) );
  AND U1442 ( .A(n819), .B(n1808), .Z(n1807) );
  IV U1443 ( .A(n1800), .Z(n1802) );
  XOR U1444 ( .A(n1809), .B(n1810), .Z(n1800) );
  AND U1445 ( .A(n823), .B(n1811), .Z(n1810) );
  XOR U1446 ( .A(n1812), .B(n1813), .Z(n1798) );
  AND U1447 ( .A(n827), .B(n1811), .Z(n1813) );
  XNOR U1448 ( .A(n1812), .B(n1809), .Z(n1811) );
  XOR U1449 ( .A(n1814), .B(n1815), .Z(n1809) );
  AND U1450 ( .A(n830), .B(n1808), .Z(n1815) );
  XNOR U1451 ( .A(n1816), .B(n1806), .Z(n1808) );
  XOR U1452 ( .A(n1817), .B(n1818), .Z(n1806) );
  AND U1453 ( .A(n834), .B(n1819), .Z(n1818) );
  XOR U1454 ( .A(p_input[1192]), .B(n1817), .Z(n1819) );
  XOR U1455 ( .A(n1820), .B(n1821), .Z(n1817) );
  AND U1456 ( .A(n838), .B(n1822), .Z(n1821) );
  IV U1457 ( .A(n1814), .Z(n1816) );
  XOR U1458 ( .A(n1823), .B(n1824), .Z(n1814) );
  AND U1459 ( .A(n842), .B(n1825), .Z(n1824) );
  XOR U1460 ( .A(n1826), .B(n1827), .Z(n1812) );
  AND U1461 ( .A(n846), .B(n1825), .Z(n1827) );
  XNOR U1462 ( .A(n1826), .B(n1823), .Z(n1825) );
  XOR U1463 ( .A(n1828), .B(n1829), .Z(n1823) );
  AND U1464 ( .A(n849), .B(n1822), .Z(n1829) );
  XNOR U1465 ( .A(n1830), .B(n1820), .Z(n1822) );
  XOR U1466 ( .A(n1831), .B(n1832), .Z(n1820) );
  AND U1467 ( .A(n853), .B(n1833), .Z(n1832) );
  XOR U1468 ( .A(p_input[1224]), .B(n1831), .Z(n1833) );
  XOR U1469 ( .A(n1834), .B(n1835), .Z(n1831) );
  AND U1470 ( .A(n857), .B(n1836), .Z(n1835) );
  IV U1471 ( .A(n1828), .Z(n1830) );
  XOR U1472 ( .A(n1837), .B(n1838), .Z(n1828) );
  AND U1473 ( .A(n861), .B(n1839), .Z(n1838) );
  XOR U1474 ( .A(n1840), .B(n1841), .Z(n1826) );
  AND U1475 ( .A(n865), .B(n1839), .Z(n1841) );
  XNOR U1476 ( .A(n1840), .B(n1837), .Z(n1839) );
  XOR U1477 ( .A(n1842), .B(n1843), .Z(n1837) );
  AND U1478 ( .A(n868), .B(n1836), .Z(n1843) );
  XNOR U1479 ( .A(n1844), .B(n1834), .Z(n1836) );
  XOR U1480 ( .A(n1845), .B(n1846), .Z(n1834) );
  AND U1481 ( .A(n872), .B(n1847), .Z(n1846) );
  XOR U1482 ( .A(p_input[1256]), .B(n1845), .Z(n1847) );
  XOR U1483 ( .A(n1848), .B(n1849), .Z(n1845) );
  AND U1484 ( .A(n876), .B(n1850), .Z(n1849) );
  IV U1485 ( .A(n1842), .Z(n1844) );
  XOR U1486 ( .A(n1851), .B(n1852), .Z(n1842) );
  AND U1487 ( .A(n880), .B(n1853), .Z(n1852) );
  XOR U1488 ( .A(n1854), .B(n1855), .Z(n1840) );
  AND U1489 ( .A(n884), .B(n1853), .Z(n1855) );
  XNOR U1490 ( .A(n1854), .B(n1851), .Z(n1853) );
  XOR U1491 ( .A(n1856), .B(n1857), .Z(n1851) );
  AND U1492 ( .A(n887), .B(n1850), .Z(n1857) );
  XNOR U1493 ( .A(n1858), .B(n1848), .Z(n1850) );
  XOR U1494 ( .A(n1859), .B(n1860), .Z(n1848) );
  AND U1495 ( .A(n891), .B(n1861), .Z(n1860) );
  XOR U1496 ( .A(p_input[1288]), .B(n1859), .Z(n1861) );
  XOR U1497 ( .A(n1862), .B(n1863), .Z(n1859) );
  AND U1498 ( .A(n895), .B(n1864), .Z(n1863) );
  IV U1499 ( .A(n1856), .Z(n1858) );
  XOR U1500 ( .A(n1865), .B(n1866), .Z(n1856) );
  AND U1501 ( .A(n899), .B(n1867), .Z(n1866) );
  XOR U1502 ( .A(n1868), .B(n1869), .Z(n1854) );
  AND U1503 ( .A(n903), .B(n1867), .Z(n1869) );
  XNOR U1504 ( .A(n1868), .B(n1865), .Z(n1867) );
  XOR U1505 ( .A(n1870), .B(n1871), .Z(n1865) );
  AND U1506 ( .A(n906), .B(n1864), .Z(n1871) );
  XNOR U1507 ( .A(n1872), .B(n1862), .Z(n1864) );
  XOR U1508 ( .A(n1873), .B(n1874), .Z(n1862) );
  AND U1509 ( .A(n910), .B(n1875), .Z(n1874) );
  XOR U1510 ( .A(p_input[1320]), .B(n1873), .Z(n1875) );
  XOR U1511 ( .A(n1876), .B(n1877), .Z(n1873) );
  AND U1512 ( .A(n914), .B(n1878), .Z(n1877) );
  IV U1513 ( .A(n1870), .Z(n1872) );
  XOR U1514 ( .A(n1879), .B(n1880), .Z(n1870) );
  AND U1515 ( .A(n918), .B(n1881), .Z(n1880) );
  XOR U1516 ( .A(n1882), .B(n1883), .Z(n1868) );
  AND U1517 ( .A(n922), .B(n1881), .Z(n1883) );
  XNOR U1518 ( .A(n1882), .B(n1879), .Z(n1881) );
  XOR U1519 ( .A(n1884), .B(n1885), .Z(n1879) );
  AND U1520 ( .A(n925), .B(n1878), .Z(n1885) );
  XNOR U1521 ( .A(n1886), .B(n1876), .Z(n1878) );
  XOR U1522 ( .A(n1887), .B(n1888), .Z(n1876) );
  AND U1523 ( .A(n929), .B(n1889), .Z(n1888) );
  XOR U1524 ( .A(p_input[1352]), .B(n1887), .Z(n1889) );
  XOR U1525 ( .A(n1890), .B(n1891), .Z(n1887) );
  AND U1526 ( .A(n933), .B(n1892), .Z(n1891) );
  IV U1527 ( .A(n1884), .Z(n1886) );
  XOR U1528 ( .A(n1893), .B(n1894), .Z(n1884) );
  AND U1529 ( .A(n937), .B(n1895), .Z(n1894) );
  XOR U1530 ( .A(n1896), .B(n1897), .Z(n1882) );
  AND U1531 ( .A(n941), .B(n1895), .Z(n1897) );
  XNOR U1532 ( .A(n1896), .B(n1893), .Z(n1895) );
  XOR U1533 ( .A(n1898), .B(n1899), .Z(n1893) );
  AND U1534 ( .A(n944), .B(n1892), .Z(n1899) );
  XNOR U1535 ( .A(n1900), .B(n1890), .Z(n1892) );
  XOR U1536 ( .A(n1901), .B(n1902), .Z(n1890) );
  AND U1537 ( .A(n948), .B(n1903), .Z(n1902) );
  XOR U1538 ( .A(p_input[1384]), .B(n1901), .Z(n1903) );
  XOR U1539 ( .A(n1904), .B(n1905), .Z(n1901) );
  AND U1540 ( .A(n952), .B(n1906), .Z(n1905) );
  IV U1541 ( .A(n1898), .Z(n1900) );
  XOR U1542 ( .A(n1907), .B(n1908), .Z(n1898) );
  AND U1543 ( .A(n956), .B(n1909), .Z(n1908) );
  XOR U1544 ( .A(n1910), .B(n1911), .Z(n1896) );
  AND U1545 ( .A(n960), .B(n1909), .Z(n1911) );
  XNOR U1546 ( .A(n1910), .B(n1907), .Z(n1909) );
  XOR U1547 ( .A(n1912), .B(n1913), .Z(n1907) );
  AND U1548 ( .A(n963), .B(n1906), .Z(n1913) );
  XNOR U1549 ( .A(n1914), .B(n1904), .Z(n1906) );
  XOR U1550 ( .A(n1915), .B(n1916), .Z(n1904) );
  AND U1551 ( .A(n967), .B(n1917), .Z(n1916) );
  XOR U1552 ( .A(p_input[1416]), .B(n1915), .Z(n1917) );
  XOR U1553 ( .A(n1918), .B(n1919), .Z(n1915) );
  AND U1554 ( .A(n971), .B(n1920), .Z(n1919) );
  IV U1555 ( .A(n1912), .Z(n1914) );
  XOR U1556 ( .A(n1921), .B(n1922), .Z(n1912) );
  AND U1557 ( .A(n975), .B(n1923), .Z(n1922) );
  XOR U1558 ( .A(n1924), .B(n1925), .Z(n1910) );
  AND U1559 ( .A(n979), .B(n1923), .Z(n1925) );
  XNOR U1560 ( .A(n1924), .B(n1921), .Z(n1923) );
  XOR U1561 ( .A(n1926), .B(n1927), .Z(n1921) );
  AND U1562 ( .A(n982), .B(n1920), .Z(n1927) );
  XNOR U1563 ( .A(n1928), .B(n1918), .Z(n1920) );
  XOR U1564 ( .A(n1929), .B(n1930), .Z(n1918) );
  AND U1565 ( .A(n986), .B(n1931), .Z(n1930) );
  XOR U1566 ( .A(p_input[1448]), .B(n1929), .Z(n1931) );
  XOR U1567 ( .A(n1932), .B(n1933), .Z(n1929) );
  AND U1568 ( .A(n990), .B(n1934), .Z(n1933) );
  IV U1569 ( .A(n1926), .Z(n1928) );
  XOR U1570 ( .A(n1935), .B(n1936), .Z(n1926) );
  AND U1571 ( .A(n994), .B(n1937), .Z(n1936) );
  XOR U1572 ( .A(n1938), .B(n1939), .Z(n1924) );
  AND U1573 ( .A(n998), .B(n1937), .Z(n1939) );
  XNOR U1574 ( .A(n1938), .B(n1935), .Z(n1937) );
  XOR U1575 ( .A(n1940), .B(n1941), .Z(n1935) );
  AND U1576 ( .A(n1001), .B(n1934), .Z(n1941) );
  XNOR U1577 ( .A(n1942), .B(n1932), .Z(n1934) );
  XOR U1578 ( .A(n1943), .B(n1944), .Z(n1932) );
  AND U1579 ( .A(n1005), .B(n1945), .Z(n1944) );
  XOR U1580 ( .A(p_input[1480]), .B(n1943), .Z(n1945) );
  XOR U1581 ( .A(n1946), .B(n1947), .Z(n1943) );
  AND U1582 ( .A(n1009), .B(n1948), .Z(n1947) );
  IV U1583 ( .A(n1940), .Z(n1942) );
  XOR U1584 ( .A(n1949), .B(n1950), .Z(n1940) );
  AND U1585 ( .A(n1013), .B(n1951), .Z(n1950) );
  XOR U1586 ( .A(n1952), .B(n1953), .Z(n1938) );
  AND U1587 ( .A(n1017), .B(n1951), .Z(n1953) );
  XNOR U1588 ( .A(n1952), .B(n1949), .Z(n1951) );
  XOR U1589 ( .A(n1954), .B(n1955), .Z(n1949) );
  AND U1590 ( .A(n1020), .B(n1948), .Z(n1955) );
  XNOR U1591 ( .A(n1956), .B(n1946), .Z(n1948) );
  XOR U1592 ( .A(n1957), .B(n1958), .Z(n1946) );
  AND U1593 ( .A(n1024), .B(n1959), .Z(n1958) );
  XOR U1594 ( .A(p_input[1512]), .B(n1957), .Z(n1959) );
  XOR U1595 ( .A(n1960), .B(n1961), .Z(n1957) );
  AND U1596 ( .A(n1028), .B(n1962), .Z(n1961) );
  IV U1597 ( .A(n1954), .Z(n1956) );
  XOR U1598 ( .A(n1963), .B(n1964), .Z(n1954) );
  AND U1599 ( .A(n1032), .B(n1965), .Z(n1964) );
  XOR U1600 ( .A(n1966), .B(n1967), .Z(n1952) );
  AND U1601 ( .A(n1036), .B(n1965), .Z(n1967) );
  XNOR U1602 ( .A(n1966), .B(n1963), .Z(n1965) );
  XOR U1603 ( .A(n1968), .B(n1969), .Z(n1963) );
  AND U1604 ( .A(n1039), .B(n1962), .Z(n1969) );
  XNOR U1605 ( .A(n1970), .B(n1960), .Z(n1962) );
  XOR U1606 ( .A(n1971), .B(n1972), .Z(n1960) );
  AND U1607 ( .A(n1043), .B(n1973), .Z(n1972) );
  XOR U1608 ( .A(p_input[1544]), .B(n1971), .Z(n1973) );
  XOR U1609 ( .A(n1974), .B(n1975), .Z(n1971) );
  AND U1610 ( .A(n1047), .B(n1976), .Z(n1975) );
  IV U1611 ( .A(n1968), .Z(n1970) );
  XOR U1612 ( .A(n1977), .B(n1978), .Z(n1968) );
  AND U1613 ( .A(n1051), .B(n1979), .Z(n1978) );
  XOR U1614 ( .A(n1980), .B(n1981), .Z(n1966) );
  AND U1615 ( .A(n1055), .B(n1979), .Z(n1981) );
  XNOR U1616 ( .A(n1980), .B(n1977), .Z(n1979) );
  XOR U1617 ( .A(n1982), .B(n1983), .Z(n1977) );
  AND U1618 ( .A(n1058), .B(n1976), .Z(n1983) );
  XNOR U1619 ( .A(n1984), .B(n1974), .Z(n1976) );
  XOR U1620 ( .A(n1985), .B(n1986), .Z(n1974) );
  AND U1621 ( .A(n1062), .B(n1987), .Z(n1986) );
  XOR U1622 ( .A(p_input[1576]), .B(n1985), .Z(n1987) );
  XOR U1623 ( .A(n1988), .B(n1989), .Z(n1985) );
  AND U1624 ( .A(n1066), .B(n1990), .Z(n1989) );
  IV U1625 ( .A(n1982), .Z(n1984) );
  XOR U1626 ( .A(n1991), .B(n1992), .Z(n1982) );
  AND U1627 ( .A(n1070), .B(n1993), .Z(n1992) );
  XOR U1628 ( .A(n1994), .B(n1995), .Z(n1980) );
  AND U1629 ( .A(n1074), .B(n1993), .Z(n1995) );
  XNOR U1630 ( .A(n1994), .B(n1991), .Z(n1993) );
  XOR U1631 ( .A(n1996), .B(n1997), .Z(n1991) );
  AND U1632 ( .A(n1077), .B(n1990), .Z(n1997) );
  XNOR U1633 ( .A(n1998), .B(n1988), .Z(n1990) );
  XOR U1634 ( .A(n1999), .B(n2000), .Z(n1988) );
  AND U1635 ( .A(n1081), .B(n2001), .Z(n2000) );
  XOR U1636 ( .A(p_input[1608]), .B(n1999), .Z(n2001) );
  XOR U1637 ( .A(n2002), .B(n2003), .Z(n1999) );
  AND U1638 ( .A(n1085), .B(n2004), .Z(n2003) );
  IV U1639 ( .A(n1996), .Z(n1998) );
  XOR U1640 ( .A(n2005), .B(n2006), .Z(n1996) );
  AND U1641 ( .A(n1089), .B(n2007), .Z(n2006) );
  XOR U1642 ( .A(n2008), .B(n2009), .Z(n1994) );
  AND U1643 ( .A(n1093), .B(n2007), .Z(n2009) );
  XNOR U1644 ( .A(n2008), .B(n2005), .Z(n2007) );
  XOR U1645 ( .A(n2010), .B(n2011), .Z(n2005) );
  AND U1646 ( .A(n1096), .B(n2004), .Z(n2011) );
  XNOR U1647 ( .A(n2012), .B(n2002), .Z(n2004) );
  XOR U1648 ( .A(n2013), .B(n2014), .Z(n2002) );
  AND U1649 ( .A(n1100), .B(n2015), .Z(n2014) );
  XOR U1650 ( .A(p_input[1640]), .B(n2013), .Z(n2015) );
  XOR U1651 ( .A(n2016), .B(n2017), .Z(n2013) );
  AND U1652 ( .A(n1104), .B(n2018), .Z(n2017) );
  IV U1653 ( .A(n2010), .Z(n2012) );
  XOR U1654 ( .A(n2019), .B(n2020), .Z(n2010) );
  AND U1655 ( .A(n1108), .B(n2021), .Z(n2020) );
  XOR U1656 ( .A(n2022), .B(n2023), .Z(n2008) );
  AND U1657 ( .A(n1112), .B(n2021), .Z(n2023) );
  XNOR U1658 ( .A(n2022), .B(n2019), .Z(n2021) );
  XOR U1659 ( .A(n2024), .B(n2025), .Z(n2019) );
  AND U1660 ( .A(n1115), .B(n2018), .Z(n2025) );
  XNOR U1661 ( .A(n2026), .B(n2016), .Z(n2018) );
  XOR U1662 ( .A(n2027), .B(n2028), .Z(n2016) );
  AND U1663 ( .A(n1119), .B(n2029), .Z(n2028) );
  XOR U1664 ( .A(p_input[1672]), .B(n2027), .Z(n2029) );
  XOR U1665 ( .A(n2030), .B(n2031), .Z(n2027) );
  AND U1666 ( .A(n1123), .B(n2032), .Z(n2031) );
  IV U1667 ( .A(n2024), .Z(n2026) );
  XOR U1668 ( .A(n2033), .B(n2034), .Z(n2024) );
  AND U1669 ( .A(n1127), .B(n2035), .Z(n2034) );
  XOR U1670 ( .A(n2036), .B(n2037), .Z(n2022) );
  AND U1671 ( .A(n1131), .B(n2035), .Z(n2037) );
  XNOR U1672 ( .A(n2036), .B(n2033), .Z(n2035) );
  XOR U1673 ( .A(n2038), .B(n2039), .Z(n2033) );
  AND U1674 ( .A(n1134), .B(n2032), .Z(n2039) );
  XNOR U1675 ( .A(n2040), .B(n2030), .Z(n2032) );
  XOR U1676 ( .A(n2041), .B(n2042), .Z(n2030) );
  AND U1677 ( .A(n1138), .B(n2043), .Z(n2042) );
  XOR U1678 ( .A(p_input[1704]), .B(n2041), .Z(n2043) );
  XOR U1679 ( .A(n2044), .B(n2045), .Z(n2041) );
  AND U1680 ( .A(n1142), .B(n2046), .Z(n2045) );
  IV U1681 ( .A(n2038), .Z(n2040) );
  XOR U1682 ( .A(n2047), .B(n2048), .Z(n2038) );
  AND U1683 ( .A(n1146), .B(n2049), .Z(n2048) );
  XOR U1684 ( .A(n2050), .B(n2051), .Z(n2036) );
  AND U1685 ( .A(n1150), .B(n2049), .Z(n2051) );
  XNOR U1686 ( .A(n2050), .B(n2047), .Z(n2049) );
  XOR U1687 ( .A(n2052), .B(n2053), .Z(n2047) );
  AND U1688 ( .A(n1153), .B(n2046), .Z(n2053) );
  XNOR U1689 ( .A(n2054), .B(n2044), .Z(n2046) );
  XOR U1690 ( .A(n2055), .B(n2056), .Z(n2044) );
  AND U1691 ( .A(n1157), .B(n2057), .Z(n2056) );
  XOR U1692 ( .A(p_input[1736]), .B(n2055), .Z(n2057) );
  XOR U1693 ( .A(n2058), .B(n2059), .Z(n2055) );
  AND U1694 ( .A(n1161), .B(n2060), .Z(n2059) );
  IV U1695 ( .A(n2052), .Z(n2054) );
  XOR U1696 ( .A(n2061), .B(n2062), .Z(n2052) );
  AND U1697 ( .A(n1165), .B(n2063), .Z(n2062) );
  XOR U1698 ( .A(n2064), .B(n2065), .Z(n2050) );
  AND U1699 ( .A(n1169), .B(n2063), .Z(n2065) );
  XNOR U1700 ( .A(n2064), .B(n2061), .Z(n2063) );
  XOR U1701 ( .A(n2066), .B(n2067), .Z(n2061) );
  AND U1702 ( .A(n1172), .B(n2060), .Z(n2067) );
  XNOR U1703 ( .A(n2068), .B(n2058), .Z(n2060) );
  XOR U1704 ( .A(n2069), .B(n2070), .Z(n2058) );
  AND U1705 ( .A(n1176), .B(n2071), .Z(n2070) );
  XOR U1706 ( .A(p_input[1768]), .B(n2069), .Z(n2071) );
  XOR U1707 ( .A(n2072), .B(n2073), .Z(n2069) );
  AND U1708 ( .A(n1180), .B(n2074), .Z(n2073) );
  IV U1709 ( .A(n2066), .Z(n2068) );
  XOR U1710 ( .A(n2075), .B(n2076), .Z(n2066) );
  AND U1711 ( .A(n1184), .B(n2077), .Z(n2076) );
  XOR U1712 ( .A(n2078), .B(n2079), .Z(n2064) );
  AND U1713 ( .A(n1188), .B(n2077), .Z(n2079) );
  XNOR U1714 ( .A(n2078), .B(n2075), .Z(n2077) );
  XOR U1715 ( .A(n2080), .B(n2081), .Z(n2075) );
  AND U1716 ( .A(n1191), .B(n2074), .Z(n2081) );
  XNOR U1717 ( .A(n2082), .B(n2072), .Z(n2074) );
  XOR U1718 ( .A(n2083), .B(n2084), .Z(n2072) );
  AND U1719 ( .A(n1195), .B(n2085), .Z(n2084) );
  XOR U1720 ( .A(p_input[1800]), .B(n2083), .Z(n2085) );
  XOR U1721 ( .A(n2086), .B(n2087), .Z(n2083) );
  AND U1722 ( .A(n1199), .B(n2088), .Z(n2087) );
  IV U1723 ( .A(n2080), .Z(n2082) );
  XOR U1724 ( .A(n2089), .B(n2090), .Z(n2080) );
  AND U1725 ( .A(n1203), .B(n2091), .Z(n2090) );
  XOR U1726 ( .A(n2092), .B(n2093), .Z(n2078) );
  AND U1727 ( .A(n1207), .B(n2091), .Z(n2093) );
  XNOR U1728 ( .A(n2092), .B(n2089), .Z(n2091) );
  XOR U1729 ( .A(n2094), .B(n2095), .Z(n2089) );
  AND U1730 ( .A(n1210), .B(n2088), .Z(n2095) );
  XNOR U1731 ( .A(n2096), .B(n2086), .Z(n2088) );
  XOR U1732 ( .A(n2097), .B(n2098), .Z(n2086) );
  AND U1733 ( .A(n1214), .B(n2099), .Z(n2098) );
  XOR U1734 ( .A(p_input[1832]), .B(n2097), .Z(n2099) );
  XOR U1735 ( .A(n2100), .B(n2101), .Z(n2097) );
  AND U1736 ( .A(n1218), .B(n2102), .Z(n2101) );
  IV U1737 ( .A(n2094), .Z(n2096) );
  XOR U1738 ( .A(n2103), .B(n2104), .Z(n2094) );
  AND U1739 ( .A(n1222), .B(n2105), .Z(n2104) );
  XOR U1740 ( .A(n2106), .B(n2107), .Z(n2092) );
  AND U1741 ( .A(n1226), .B(n2105), .Z(n2107) );
  XNOR U1742 ( .A(n2106), .B(n2103), .Z(n2105) );
  XOR U1743 ( .A(n2108), .B(n2109), .Z(n2103) );
  AND U1744 ( .A(n1229), .B(n2102), .Z(n2109) );
  XNOR U1745 ( .A(n2110), .B(n2100), .Z(n2102) );
  XOR U1746 ( .A(n2111), .B(n2112), .Z(n2100) );
  AND U1747 ( .A(n1233), .B(n2113), .Z(n2112) );
  XOR U1748 ( .A(p_input[1864]), .B(n2111), .Z(n2113) );
  XOR U1749 ( .A(n2114), .B(n2115), .Z(n2111) );
  AND U1750 ( .A(n1237), .B(n2116), .Z(n2115) );
  IV U1751 ( .A(n2108), .Z(n2110) );
  XOR U1752 ( .A(n2117), .B(n2118), .Z(n2108) );
  AND U1753 ( .A(n1241), .B(n2119), .Z(n2118) );
  XOR U1754 ( .A(n2120), .B(n2121), .Z(n2106) );
  AND U1755 ( .A(n1245), .B(n2119), .Z(n2121) );
  XNOR U1756 ( .A(n2120), .B(n2117), .Z(n2119) );
  XOR U1757 ( .A(n2122), .B(n2123), .Z(n2117) );
  AND U1758 ( .A(n1248), .B(n2116), .Z(n2123) );
  XNOR U1759 ( .A(n2124), .B(n2114), .Z(n2116) );
  XOR U1760 ( .A(n2125), .B(n2126), .Z(n2114) );
  AND U1761 ( .A(n1252), .B(n2127), .Z(n2126) );
  XOR U1762 ( .A(p_input[1896]), .B(n2125), .Z(n2127) );
  XOR U1763 ( .A(n2128), .B(n2129), .Z(n2125) );
  AND U1764 ( .A(n1256), .B(n2130), .Z(n2129) );
  IV U1765 ( .A(n2122), .Z(n2124) );
  XOR U1766 ( .A(n2131), .B(n2132), .Z(n2122) );
  AND U1767 ( .A(n1260), .B(n2133), .Z(n2132) );
  XOR U1768 ( .A(n2134), .B(n2135), .Z(n2120) );
  AND U1769 ( .A(n1264), .B(n2133), .Z(n2135) );
  XNOR U1770 ( .A(n2134), .B(n2131), .Z(n2133) );
  XOR U1771 ( .A(n2136), .B(n2137), .Z(n2131) );
  AND U1772 ( .A(n1267), .B(n2130), .Z(n2137) );
  XNOR U1773 ( .A(n2138), .B(n2128), .Z(n2130) );
  XOR U1774 ( .A(n2139), .B(n2140), .Z(n2128) );
  AND U1775 ( .A(n1271), .B(n2141), .Z(n2140) );
  XOR U1776 ( .A(p_input[1928]), .B(n2139), .Z(n2141) );
  XOR U1777 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n2142), 
        .Z(n2139) );
  AND U1778 ( .A(n1274), .B(n2143), .Z(n2142) );
  IV U1779 ( .A(n2136), .Z(n2138) );
  XOR U1780 ( .A(n2144), .B(n2145), .Z(n2136) );
  AND U1781 ( .A(n1278), .B(n2146), .Z(n2145) );
  XOR U1782 ( .A(n2147), .B(n2148), .Z(n2134) );
  AND U1783 ( .A(n1282), .B(n2146), .Z(n2148) );
  XNOR U1784 ( .A(n2147), .B(n2144), .Z(n2146) );
  XNOR U1785 ( .A(n2149), .B(n2150), .Z(n2144) );
  AND U1786 ( .A(n1285), .B(n2143), .Z(n2150) );
  XNOR U1787 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n2149), 
        .Z(n2143) );
  XNOR U1788 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .B(n2151), 
        .Z(n2149) );
  AND U1789 ( .A(n1287), .B(n2152), .Z(n2151) );
  XNOR U1790 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n2153), .Z(n2147) );
  AND U1791 ( .A(n1290), .B(n2152), .Z(n2153) );
  XOR U1792 ( .A(n2154), .B(n2155), .Z(n2152) );
  IV U1793 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .Z(n2155) );
  IV U1794 ( .A(\knn_comb_/min_val_out[0][8] ), .Z(n2154) );
  XOR U1795 ( .A(n2156), .B(n2157), .Z(o[3]) );
  XOR U1796 ( .A(n37), .B(n2158), .Z(o[39]) );
  AND U1797 ( .A(n122), .B(n2159), .Z(n37) );
  XOR U1798 ( .A(n38), .B(n2158), .Z(n2159) );
  XOR U1799 ( .A(n2160), .B(n55), .Z(n2158) );
  AND U1800 ( .A(n125), .B(n2161), .Z(n55) );
  XNOR U1801 ( .A(n2162), .B(n56), .Z(n2161) );
  XOR U1802 ( .A(n2163), .B(n2164), .Z(n56) );
  AND U1803 ( .A(n130), .B(n2165), .Z(n2164) );
  XOR U1804 ( .A(p_input[7]), .B(n2163), .Z(n2165) );
  XOR U1805 ( .A(n2166), .B(n2167), .Z(n2163) );
  AND U1806 ( .A(n134), .B(n2168), .Z(n2167) );
  IV U1807 ( .A(n2160), .Z(n2162) );
  XOR U1808 ( .A(n2169), .B(n2170), .Z(n2160) );
  AND U1809 ( .A(n138), .B(n2171), .Z(n2170) );
  XOR U1810 ( .A(n2172), .B(n2173), .Z(n38) );
  AND U1811 ( .A(n142), .B(n2171), .Z(n2173) );
  XNOR U1812 ( .A(n2174), .B(n2169), .Z(n2171) );
  XOR U1813 ( .A(n2175), .B(n2176), .Z(n2169) );
  AND U1814 ( .A(n146), .B(n2168), .Z(n2176) );
  XNOR U1815 ( .A(n2177), .B(n2166), .Z(n2168) );
  XOR U1816 ( .A(n2178), .B(n2179), .Z(n2166) );
  AND U1817 ( .A(n150), .B(n2180), .Z(n2179) );
  XOR U1818 ( .A(p_input[39]), .B(n2178), .Z(n2180) );
  XOR U1819 ( .A(n2181), .B(n2182), .Z(n2178) );
  AND U1820 ( .A(n154), .B(n2183), .Z(n2182) );
  IV U1821 ( .A(n2175), .Z(n2177) );
  XOR U1822 ( .A(n2184), .B(n2185), .Z(n2175) );
  AND U1823 ( .A(n158), .B(n2186), .Z(n2185) );
  IV U1824 ( .A(n2172), .Z(n2174) );
  XNOR U1825 ( .A(n2187), .B(n2188), .Z(n2172) );
  AND U1826 ( .A(n162), .B(n2186), .Z(n2188) );
  XNOR U1827 ( .A(n2187), .B(n2184), .Z(n2186) );
  XOR U1828 ( .A(n2189), .B(n2190), .Z(n2184) );
  AND U1829 ( .A(n165), .B(n2183), .Z(n2190) );
  XNOR U1830 ( .A(n2191), .B(n2181), .Z(n2183) );
  XOR U1831 ( .A(n2192), .B(n2193), .Z(n2181) );
  AND U1832 ( .A(n169), .B(n2194), .Z(n2193) );
  XOR U1833 ( .A(p_input[71]), .B(n2192), .Z(n2194) );
  XOR U1834 ( .A(n2195), .B(n2196), .Z(n2192) );
  AND U1835 ( .A(n173), .B(n2197), .Z(n2196) );
  IV U1836 ( .A(n2189), .Z(n2191) );
  XOR U1837 ( .A(n2198), .B(n2199), .Z(n2189) );
  AND U1838 ( .A(n177), .B(n2200), .Z(n2199) );
  XOR U1839 ( .A(n2201), .B(n2202), .Z(n2187) );
  AND U1840 ( .A(n181), .B(n2200), .Z(n2202) );
  XNOR U1841 ( .A(n2201), .B(n2198), .Z(n2200) );
  XOR U1842 ( .A(n2203), .B(n2204), .Z(n2198) );
  AND U1843 ( .A(n184), .B(n2197), .Z(n2204) );
  XNOR U1844 ( .A(n2205), .B(n2195), .Z(n2197) );
  XOR U1845 ( .A(n2206), .B(n2207), .Z(n2195) );
  AND U1846 ( .A(n188), .B(n2208), .Z(n2207) );
  XOR U1847 ( .A(p_input[103]), .B(n2206), .Z(n2208) );
  XOR U1848 ( .A(n2209), .B(n2210), .Z(n2206) );
  AND U1849 ( .A(n192), .B(n2211), .Z(n2210) );
  IV U1850 ( .A(n2203), .Z(n2205) );
  XOR U1851 ( .A(n2212), .B(n2213), .Z(n2203) );
  AND U1852 ( .A(n196), .B(n2214), .Z(n2213) );
  XOR U1853 ( .A(n2215), .B(n2216), .Z(n2201) );
  AND U1854 ( .A(n200), .B(n2214), .Z(n2216) );
  XNOR U1855 ( .A(n2215), .B(n2212), .Z(n2214) );
  XOR U1856 ( .A(n2217), .B(n2218), .Z(n2212) );
  AND U1857 ( .A(n203), .B(n2211), .Z(n2218) );
  XNOR U1858 ( .A(n2219), .B(n2209), .Z(n2211) );
  XOR U1859 ( .A(n2220), .B(n2221), .Z(n2209) );
  AND U1860 ( .A(n207), .B(n2222), .Z(n2221) );
  XOR U1861 ( .A(p_input[135]), .B(n2220), .Z(n2222) );
  XOR U1862 ( .A(n2223), .B(n2224), .Z(n2220) );
  AND U1863 ( .A(n211), .B(n2225), .Z(n2224) );
  IV U1864 ( .A(n2217), .Z(n2219) );
  XOR U1865 ( .A(n2226), .B(n2227), .Z(n2217) );
  AND U1866 ( .A(n215), .B(n2228), .Z(n2227) );
  XOR U1867 ( .A(n2229), .B(n2230), .Z(n2215) );
  AND U1868 ( .A(n219), .B(n2228), .Z(n2230) );
  XNOR U1869 ( .A(n2229), .B(n2226), .Z(n2228) );
  XOR U1870 ( .A(n2231), .B(n2232), .Z(n2226) );
  AND U1871 ( .A(n222), .B(n2225), .Z(n2232) );
  XNOR U1872 ( .A(n2233), .B(n2223), .Z(n2225) );
  XOR U1873 ( .A(n2234), .B(n2235), .Z(n2223) );
  AND U1874 ( .A(n226), .B(n2236), .Z(n2235) );
  XOR U1875 ( .A(p_input[167]), .B(n2234), .Z(n2236) );
  XOR U1876 ( .A(n2237), .B(n2238), .Z(n2234) );
  AND U1877 ( .A(n230), .B(n2239), .Z(n2238) );
  IV U1878 ( .A(n2231), .Z(n2233) );
  XOR U1879 ( .A(n2240), .B(n2241), .Z(n2231) );
  AND U1880 ( .A(n234), .B(n2242), .Z(n2241) );
  XOR U1881 ( .A(n2243), .B(n2244), .Z(n2229) );
  AND U1882 ( .A(n238), .B(n2242), .Z(n2244) );
  XNOR U1883 ( .A(n2243), .B(n2240), .Z(n2242) );
  XOR U1884 ( .A(n2245), .B(n2246), .Z(n2240) );
  AND U1885 ( .A(n241), .B(n2239), .Z(n2246) );
  XNOR U1886 ( .A(n2247), .B(n2237), .Z(n2239) );
  XOR U1887 ( .A(n2248), .B(n2249), .Z(n2237) );
  AND U1888 ( .A(n245), .B(n2250), .Z(n2249) );
  XOR U1889 ( .A(p_input[199]), .B(n2248), .Z(n2250) );
  XOR U1890 ( .A(n2251), .B(n2252), .Z(n2248) );
  AND U1891 ( .A(n249), .B(n2253), .Z(n2252) );
  IV U1892 ( .A(n2245), .Z(n2247) );
  XOR U1893 ( .A(n2254), .B(n2255), .Z(n2245) );
  AND U1894 ( .A(n253), .B(n2256), .Z(n2255) );
  XOR U1895 ( .A(n2257), .B(n2258), .Z(n2243) );
  AND U1896 ( .A(n257), .B(n2256), .Z(n2258) );
  XNOR U1897 ( .A(n2257), .B(n2254), .Z(n2256) );
  XOR U1898 ( .A(n2259), .B(n2260), .Z(n2254) );
  AND U1899 ( .A(n260), .B(n2253), .Z(n2260) );
  XNOR U1900 ( .A(n2261), .B(n2251), .Z(n2253) );
  XOR U1901 ( .A(n2262), .B(n2263), .Z(n2251) );
  AND U1902 ( .A(n264), .B(n2264), .Z(n2263) );
  XOR U1903 ( .A(p_input[231]), .B(n2262), .Z(n2264) );
  XOR U1904 ( .A(n2265), .B(n2266), .Z(n2262) );
  AND U1905 ( .A(n268), .B(n2267), .Z(n2266) );
  IV U1906 ( .A(n2259), .Z(n2261) );
  XOR U1907 ( .A(n2268), .B(n2269), .Z(n2259) );
  AND U1908 ( .A(n272), .B(n2270), .Z(n2269) );
  XOR U1909 ( .A(n2271), .B(n2272), .Z(n2257) );
  AND U1910 ( .A(n276), .B(n2270), .Z(n2272) );
  XNOR U1911 ( .A(n2271), .B(n2268), .Z(n2270) );
  XOR U1912 ( .A(n2273), .B(n2274), .Z(n2268) );
  AND U1913 ( .A(n279), .B(n2267), .Z(n2274) );
  XNOR U1914 ( .A(n2275), .B(n2265), .Z(n2267) );
  XOR U1915 ( .A(n2276), .B(n2277), .Z(n2265) );
  AND U1916 ( .A(n283), .B(n2278), .Z(n2277) );
  XOR U1917 ( .A(p_input[263]), .B(n2276), .Z(n2278) );
  XOR U1918 ( .A(n2279), .B(n2280), .Z(n2276) );
  AND U1919 ( .A(n287), .B(n2281), .Z(n2280) );
  IV U1920 ( .A(n2273), .Z(n2275) );
  XOR U1921 ( .A(n2282), .B(n2283), .Z(n2273) );
  AND U1922 ( .A(n291), .B(n2284), .Z(n2283) );
  XOR U1923 ( .A(n2285), .B(n2286), .Z(n2271) );
  AND U1924 ( .A(n295), .B(n2284), .Z(n2286) );
  XNOR U1925 ( .A(n2285), .B(n2282), .Z(n2284) );
  XOR U1926 ( .A(n2287), .B(n2288), .Z(n2282) );
  AND U1927 ( .A(n298), .B(n2281), .Z(n2288) );
  XNOR U1928 ( .A(n2289), .B(n2279), .Z(n2281) );
  XOR U1929 ( .A(n2290), .B(n2291), .Z(n2279) );
  AND U1930 ( .A(n302), .B(n2292), .Z(n2291) );
  XOR U1931 ( .A(p_input[295]), .B(n2290), .Z(n2292) );
  XOR U1932 ( .A(n2293), .B(n2294), .Z(n2290) );
  AND U1933 ( .A(n306), .B(n2295), .Z(n2294) );
  IV U1934 ( .A(n2287), .Z(n2289) );
  XOR U1935 ( .A(n2296), .B(n2297), .Z(n2287) );
  AND U1936 ( .A(n310), .B(n2298), .Z(n2297) );
  XOR U1937 ( .A(n2299), .B(n2300), .Z(n2285) );
  AND U1938 ( .A(n314), .B(n2298), .Z(n2300) );
  XNOR U1939 ( .A(n2299), .B(n2296), .Z(n2298) );
  XOR U1940 ( .A(n2301), .B(n2302), .Z(n2296) );
  AND U1941 ( .A(n317), .B(n2295), .Z(n2302) );
  XNOR U1942 ( .A(n2303), .B(n2293), .Z(n2295) );
  XOR U1943 ( .A(n2304), .B(n2305), .Z(n2293) );
  AND U1944 ( .A(n321), .B(n2306), .Z(n2305) );
  XOR U1945 ( .A(p_input[327]), .B(n2304), .Z(n2306) );
  XOR U1946 ( .A(n2307), .B(n2308), .Z(n2304) );
  AND U1947 ( .A(n325), .B(n2309), .Z(n2308) );
  IV U1948 ( .A(n2301), .Z(n2303) );
  XOR U1949 ( .A(n2310), .B(n2311), .Z(n2301) );
  AND U1950 ( .A(n329), .B(n2312), .Z(n2311) );
  XOR U1951 ( .A(n2313), .B(n2314), .Z(n2299) );
  AND U1952 ( .A(n333), .B(n2312), .Z(n2314) );
  XNOR U1953 ( .A(n2313), .B(n2310), .Z(n2312) );
  XOR U1954 ( .A(n2315), .B(n2316), .Z(n2310) );
  AND U1955 ( .A(n336), .B(n2309), .Z(n2316) );
  XNOR U1956 ( .A(n2317), .B(n2307), .Z(n2309) );
  XOR U1957 ( .A(n2318), .B(n2319), .Z(n2307) );
  AND U1958 ( .A(n340), .B(n2320), .Z(n2319) );
  XOR U1959 ( .A(p_input[359]), .B(n2318), .Z(n2320) );
  XOR U1960 ( .A(n2321), .B(n2322), .Z(n2318) );
  AND U1961 ( .A(n344), .B(n2323), .Z(n2322) );
  IV U1962 ( .A(n2315), .Z(n2317) );
  XOR U1963 ( .A(n2324), .B(n2325), .Z(n2315) );
  AND U1964 ( .A(n348), .B(n2326), .Z(n2325) );
  XOR U1965 ( .A(n2327), .B(n2328), .Z(n2313) );
  AND U1966 ( .A(n352), .B(n2326), .Z(n2328) );
  XNOR U1967 ( .A(n2327), .B(n2324), .Z(n2326) );
  XOR U1968 ( .A(n2329), .B(n2330), .Z(n2324) );
  AND U1969 ( .A(n355), .B(n2323), .Z(n2330) );
  XNOR U1970 ( .A(n2331), .B(n2321), .Z(n2323) );
  XOR U1971 ( .A(n2332), .B(n2333), .Z(n2321) );
  AND U1972 ( .A(n359), .B(n2334), .Z(n2333) );
  XOR U1973 ( .A(p_input[391]), .B(n2332), .Z(n2334) );
  XOR U1974 ( .A(n2335), .B(n2336), .Z(n2332) );
  AND U1975 ( .A(n363), .B(n2337), .Z(n2336) );
  IV U1976 ( .A(n2329), .Z(n2331) );
  XOR U1977 ( .A(n2338), .B(n2339), .Z(n2329) );
  AND U1978 ( .A(n367), .B(n2340), .Z(n2339) );
  XOR U1979 ( .A(n2341), .B(n2342), .Z(n2327) );
  AND U1980 ( .A(n371), .B(n2340), .Z(n2342) );
  XNOR U1981 ( .A(n2341), .B(n2338), .Z(n2340) );
  XOR U1982 ( .A(n2343), .B(n2344), .Z(n2338) );
  AND U1983 ( .A(n374), .B(n2337), .Z(n2344) );
  XNOR U1984 ( .A(n2345), .B(n2335), .Z(n2337) );
  XOR U1985 ( .A(n2346), .B(n2347), .Z(n2335) );
  AND U1986 ( .A(n378), .B(n2348), .Z(n2347) );
  XOR U1987 ( .A(p_input[423]), .B(n2346), .Z(n2348) );
  XOR U1988 ( .A(n2349), .B(n2350), .Z(n2346) );
  AND U1989 ( .A(n382), .B(n2351), .Z(n2350) );
  IV U1990 ( .A(n2343), .Z(n2345) );
  XOR U1991 ( .A(n2352), .B(n2353), .Z(n2343) );
  AND U1992 ( .A(n386), .B(n2354), .Z(n2353) );
  XOR U1993 ( .A(n2355), .B(n2356), .Z(n2341) );
  AND U1994 ( .A(n390), .B(n2354), .Z(n2356) );
  XNOR U1995 ( .A(n2355), .B(n2352), .Z(n2354) );
  XOR U1996 ( .A(n2357), .B(n2358), .Z(n2352) );
  AND U1997 ( .A(n393), .B(n2351), .Z(n2358) );
  XNOR U1998 ( .A(n2359), .B(n2349), .Z(n2351) );
  XOR U1999 ( .A(n2360), .B(n2361), .Z(n2349) );
  AND U2000 ( .A(n397), .B(n2362), .Z(n2361) );
  XOR U2001 ( .A(p_input[455]), .B(n2360), .Z(n2362) );
  XOR U2002 ( .A(n2363), .B(n2364), .Z(n2360) );
  AND U2003 ( .A(n401), .B(n2365), .Z(n2364) );
  IV U2004 ( .A(n2357), .Z(n2359) );
  XOR U2005 ( .A(n2366), .B(n2367), .Z(n2357) );
  AND U2006 ( .A(n405), .B(n2368), .Z(n2367) );
  XOR U2007 ( .A(n2369), .B(n2370), .Z(n2355) );
  AND U2008 ( .A(n409), .B(n2368), .Z(n2370) );
  XNOR U2009 ( .A(n2369), .B(n2366), .Z(n2368) );
  XOR U2010 ( .A(n2371), .B(n2372), .Z(n2366) );
  AND U2011 ( .A(n412), .B(n2365), .Z(n2372) );
  XNOR U2012 ( .A(n2373), .B(n2363), .Z(n2365) );
  XOR U2013 ( .A(n2374), .B(n2375), .Z(n2363) );
  AND U2014 ( .A(n416), .B(n2376), .Z(n2375) );
  XOR U2015 ( .A(p_input[487]), .B(n2374), .Z(n2376) );
  XOR U2016 ( .A(n2377), .B(n2378), .Z(n2374) );
  AND U2017 ( .A(n420), .B(n2379), .Z(n2378) );
  IV U2018 ( .A(n2371), .Z(n2373) );
  XOR U2019 ( .A(n2380), .B(n2381), .Z(n2371) );
  AND U2020 ( .A(n424), .B(n2382), .Z(n2381) );
  XOR U2021 ( .A(n2383), .B(n2384), .Z(n2369) );
  AND U2022 ( .A(n428), .B(n2382), .Z(n2384) );
  XNOR U2023 ( .A(n2383), .B(n2380), .Z(n2382) );
  XOR U2024 ( .A(n2385), .B(n2386), .Z(n2380) );
  AND U2025 ( .A(n431), .B(n2379), .Z(n2386) );
  XNOR U2026 ( .A(n2387), .B(n2377), .Z(n2379) );
  XOR U2027 ( .A(n2388), .B(n2389), .Z(n2377) );
  AND U2028 ( .A(n435), .B(n2390), .Z(n2389) );
  XOR U2029 ( .A(p_input[519]), .B(n2388), .Z(n2390) );
  XOR U2030 ( .A(n2391), .B(n2392), .Z(n2388) );
  AND U2031 ( .A(n439), .B(n2393), .Z(n2392) );
  IV U2032 ( .A(n2385), .Z(n2387) );
  XOR U2033 ( .A(n2394), .B(n2395), .Z(n2385) );
  AND U2034 ( .A(n443), .B(n2396), .Z(n2395) );
  XOR U2035 ( .A(n2397), .B(n2398), .Z(n2383) );
  AND U2036 ( .A(n447), .B(n2396), .Z(n2398) );
  XNOR U2037 ( .A(n2397), .B(n2394), .Z(n2396) );
  XOR U2038 ( .A(n2399), .B(n2400), .Z(n2394) );
  AND U2039 ( .A(n450), .B(n2393), .Z(n2400) );
  XNOR U2040 ( .A(n2401), .B(n2391), .Z(n2393) );
  XOR U2041 ( .A(n2402), .B(n2403), .Z(n2391) );
  AND U2042 ( .A(n454), .B(n2404), .Z(n2403) );
  XOR U2043 ( .A(p_input[551]), .B(n2402), .Z(n2404) );
  XOR U2044 ( .A(n2405), .B(n2406), .Z(n2402) );
  AND U2045 ( .A(n458), .B(n2407), .Z(n2406) );
  IV U2046 ( .A(n2399), .Z(n2401) );
  XOR U2047 ( .A(n2408), .B(n2409), .Z(n2399) );
  AND U2048 ( .A(n462), .B(n2410), .Z(n2409) );
  XOR U2049 ( .A(n2411), .B(n2412), .Z(n2397) );
  AND U2050 ( .A(n466), .B(n2410), .Z(n2412) );
  XNOR U2051 ( .A(n2411), .B(n2408), .Z(n2410) );
  XOR U2052 ( .A(n2413), .B(n2414), .Z(n2408) );
  AND U2053 ( .A(n469), .B(n2407), .Z(n2414) );
  XNOR U2054 ( .A(n2415), .B(n2405), .Z(n2407) );
  XOR U2055 ( .A(n2416), .B(n2417), .Z(n2405) );
  AND U2056 ( .A(n473), .B(n2418), .Z(n2417) );
  XOR U2057 ( .A(p_input[583]), .B(n2416), .Z(n2418) );
  XOR U2058 ( .A(n2419), .B(n2420), .Z(n2416) );
  AND U2059 ( .A(n477), .B(n2421), .Z(n2420) );
  IV U2060 ( .A(n2413), .Z(n2415) );
  XOR U2061 ( .A(n2422), .B(n2423), .Z(n2413) );
  AND U2062 ( .A(n481), .B(n2424), .Z(n2423) );
  XOR U2063 ( .A(n2425), .B(n2426), .Z(n2411) );
  AND U2064 ( .A(n485), .B(n2424), .Z(n2426) );
  XNOR U2065 ( .A(n2425), .B(n2422), .Z(n2424) );
  XOR U2066 ( .A(n2427), .B(n2428), .Z(n2422) );
  AND U2067 ( .A(n488), .B(n2421), .Z(n2428) );
  XNOR U2068 ( .A(n2429), .B(n2419), .Z(n2421) );
  XOR U2069 ( .A(n2430), .B(n2431), .Z(n2419) );
  AND U2070 ( .A(n492), .B(n2432), .Z(n2431) );
  XOR U2071 ( .A(p_input[615]), .B(n2430), .Z(n2432) );
  XOR U2072 ( .A(n2433), .B(n2434), .Z(n2430) );
  AND U2073 ( .A(n496), .B(n2435), .Z(n2434) );
  IV U2074 ( .A(n2427), .Z(n2429) );
  XOR U2075 ( .A(n2436), .B(n2437), .Z(n2427) );
  AND U2076 ( .A(n500), .B(n2438), .Z(n2437) );
  XOR U2077 ( .A(n2439), .B(n2440), .Z(n2425) );
  AND U2078 ( .A(n504), .B(n2438), .Z(n2440) );
  XNOR U2079 ( .A(n2439), .B(n2436), .Z(n2438) );
  XOR U2080 ( .A(n2441), .B(n2442), .Z(n2436) );
  AND U2081 ( .A(n507), .B(n2435), .Z(n2442) );
  XNOR U2082 ( .A(n2443), .B(n2433), .Z(n2435) );
  XOR U2083 ( .A(n2444), .B(n2445), .Z(n2433) );
  AND U2084 ( .A(n511), .B(n2446), .Z(n2445) );
  XOR U2085 ( .A(p_input[647]), .B(n2444), .Z(n2446) );
  XOR U2086 ( .A(n2447), .B(n2448), .Z(n2444) );
  AND U2087 ( .A(n515), .B(n2449), .Z(n2448) );
  IV U2088 ( .A(n2441), .Z(n2443) );
  XOR U2089 ( .A(n2450), .B(n2451), .Z(n2441) );
  AND U2090 ( .A(n519), .B(n2452), .Z(n2451) );
  XOR U2091 ( .A(n2453), .B(n2454), .Z(n2439) );
  AND U2092 ( .A(n523), .B(n2452), .Z(n2454) );
  XNOR U2093 ( .A(n2453), .B(n2450), .Z(n2452) );
  XOR U2094 ( .A(n2455), .B(n2456), .Z(n2450) );
  AND U2095 ( .A(n526), .B(n2449), .Z(n2456) );
  XNOR U2096 ( .A(n2457), .B(n2447), .Z(n2449) );
  XOR U2097 ( .A(n2458), .B(n2459), .Z(n2447) );
  AND U2098 ( .A(n530), .B(n2460), .Z(n2459) );
  XOR U2099 ( .A(p_input[679]), .B(n2458), .Z(n2460) );
  XOR U2100 ( .A(n2461), .B(n2462), .Z(n2458) );
  AND U2101 ( .A(n534), .B(n2463), .Z(n2462) );
  IV U2102 ( .A(n2455), .Z(n2457) );
  XOR U2103 ( .A(n2464), .B(n2465), .Z(n2455) );
  AND U2104 ( .A(n538), .B(n2466), .Z(n2465) );
  XOR U2105 ( .A(n2467), .B(n2468), .Z(n2453) );
  AND U2106 ( .A(n542), .B(n2466), .Z(n2468) );
  XNOR U2107 ( .A(n2467), .B(n2464), .Z(n2466) );
  XOR U2108 ( .A(n2469), .B(n2470), .Z(n2464) );
  AND U2109 ( .A(n545), .B(n2463), .Z(n2470) );
  XNOR U2110 ( .A(n2471), .B(n2461), .Z(n2463) );
  XOR U2111 ( .A(n2472), .B(n2473), .Z(n2461) );
  AND U2112 ( .A(n549), .B(n2474), .Z(n2473) );
  XOR U2113 ( .A(p_input[711]), .B(n2472), .Z(n2474) );
  XOR U2114 ( .A(n2475), .B(n2476), .Z(n2472) );
  AND U2115 ( .A(n553), .B(n2477), .Z(n2476) );
  IV U2116 ( .A(n2469), .Z(n2471) );
  XOR U2117 ( .A(n2478), .B(n2479), .Z(n2469) );
  AND U2118 ( .A(n557), .B(n2480), .Z(n2479) );
  XOR U2119 ( .A(n2481), .B(n2482), .Z(n2467) );
  AND U2120 ( .A(n561), .B(n2480), .Z(n2482) );
  XNOR U2121 ( .A(n2481), .B(n2478), .Z(n2480) );
  XOR U2122 ( .A(n2483), .B(n2484), .Z(n2478) );
  AND U2123 ( .A(n564), .B(n2477), .Z(n2484) );
  XNOR U2124 ( .A(n2485), .B(n2475), .Z(n2477) );
  XOR U2125 ( .A(n2486), .B(n2487), .Z(n2475) );
  AND U2126 ( .A(n568), .B(n2488), .Z(n2487) );
  XOR U2127 ( .A(p_input[743]), .B(n2486), .Z(n2488) );
  XOR U2128 ( .A(n2489), .B(n2490), .Z(n2486) );
  AND U2129 ( .A(n572), .B(n2491), .Z(n2490) );
  IV U2130 ( .A(n2483), .Z(n2485) );
  XOR U2131 ( .A(n2492), .B(n2493), .Z(n2483) );
  AND U2132 ( .A(n576), .B(n2494), .Z(n2493) );
  XOR U2133 ( .A(n2495), .B(n2496), .Z(n2481) );
  AND U2134 ( .A(n580), .B(n2494), .Z(n2496) );
  XNOR U2135 ( .A(n2495), .B(n2492), .Z(n2494) );
  XOR U2136 ( .A(n2497), .B(n2498), .Z(n2492) );
  AND U2137 ( .A(n583), .B(n2491), .Z(n2498) );
  XNOR U2138 ( .A(n2499), .B(n2489), .Z(n2491) );
  XOR U2139 ( .A(n2500), .B(n2501), .Z(n2489) );
  AND U2140 ( .A(n587), .B(n2502), .Z(n2501) );
  XOR U2141 ( .A(p_input[775]), .B(n2500), .Z(n2502) );
  XOR U2142 ( .A(n2503), .B(n2504), .Z(n2500) );
  AND U2143 ( .A(n591), .B(n2505), .Z(n2504) );
  IV U2144 ( .A(n2497), .Z(n2499) );
  XOR U2145 ( .A(n2506), .B(n2507), .Z(n2497) );
  AND U2146 ( .A(n595), .B(n2508), .Z(n2507) );
  XOR U2147 ( .A(n2509), .B(n2510), .Z(n2495) );
  AND U2148 ( .A(n599), .B(n2508), .Z(n2510) );
  XNOR U2149 ( .A(n2509), .B(n2506), .Z(n2508) );
  XOR U2150 ( .A(n2511), .B(n2512), .Z(n2506) );
  AND U2151 ( .A(n602), .B(n2505), .Z(n2512) );
  XNOR U2152 ( .A(n2513), .B(n2503), .Z(n2505) );
  XOR U2153 ( .A(n2514), .B(n2515), .Z(n2503) );
  AND U2154 ( .A(n606), .B(n2516), .Z(n2515) );
  XOR U2155 ( .A(p_input[807]), .B(n2514), .Z(n2516) );
  XOR U2156 ( .A(n2517), .B(n2518), .Z(n2514) );
  AND U2157 ( .A(n610), .B(n2519), .Z(n2518) );
  IV U2158 ( .A(n2511), .Z(n2513) );
  XOR U2159 ( .A(n2520), .B(n2521), .Z(n2511) );
  AND U2160 ( .A(n614), .B(n2522), .Z(n2521) );
  XOR U2161 ( .A(n2523), .B(n2524), .Z(n2509) );
  AND U2162 ( .A(n618), .B(n2522), .Z(n2524) );
  XNOR U2163 ( .A(n2523), .B(n2520), .Z(n2522) );
  XOR U2164 ( .A(n2525), .B(n2526), .Z(n2520) );
  AND U2165 ( .A(n621), .B(n2519), .Z(n2526) );
  XNOR U2166 ( .A(n2527), .B(n2517), .Z(n2519) );
  XOR U2167 ( .A(n2528), .B(n2529), .Z(n2517) );
  AND U2168 ( .A(n625), .B(n2530), .Z(n2529) );
  XOR U2169 ( .A(p_input[839]), .B(n2528), .Z(n2530) );
  XOR U2170 ( .A(n2531), .B(n2532), .Z(n2528) );
  AND U2171 ( .A(n629), .B(n2533), .Z(n2532) );
  IV U2172 ( .A(n2525), .Z(n2527) );
  XOR U2173 ( .A(n2534), .B(n2535), .Z(n2525) );
  AND U2174 ( .A(n633), .B(n2536), .Z(n2535) );
  XOR U2175 ( .A(n2537), .B(n2538), .Z(n2523) );
  AND U2176 ( .A(n637), .B(n2536), .Z(n2538) );
  XNOR U2177 ( .A(n2537), .B(n2534), .Z(n2536) );
  XOR U2178 ( .A(n2539), .B(n2540), .Z(n2534) );
  AND U2179 ( .A(n640), .B(n2533), .Z(n2540) );
  XNOR U2180 ( .A(n2541), .B(n2531), .Z(n2533) );
  XOR U2181 ( .A(n2542), .B(n2543), .Z(n2531) );
  AND U2182 ( .A(n644), .B(n2544), .Z(n2543) );
  XOR U2183 ( .A(p_input[871]), .B(n2542), .Z(n2544) );
  XOR U2184 ( .A(n2545), .B(n2546), .Z(n2542) );
  AND U2185 ( .A(n648), .B(n2547), .Z(n2546) );
  IV U2186 ( .A(n2539), .Z(n2541) );
  XOR U2187 ( .A(n2548), .B(n2549), .Z(n2539) );
  AND U2188 ( .A(n652), .B(n2550), .Z(n2549) );
  XOR U2189 ( .A(n2551), .B(n2552), .Z(n2537) );
  AND U2190 ( .A(n656), .B(n2550), .Z(n2552) );
  XNOR U2191 ( .A(n2551), .B(n2548), .Z(n2550) );
  XOR U2192 ( .A(n2553), .B(n2554), .Z(n2548) );
  AND U2193 ( .A(n659), .B(n2547), .Z(n2554) );
  XNOR U2194 ( .A(n2555), .B(n2545), .Z(n2547) );
  XOR U2195 ( .A(n2556), .B(n2557), .Z(n2545) );
  AND U2196 ( .A(n663), .B(n2558), .Z(n2557) );
  XOR U2197 ( .A(p_input[903]), .B(n2556), .Z(n2558) );
  XOR U2198 ( .A(n2559), .B(n2560), .Z(n2556) );
  AND U2199 ( .A(n667), .B(n2561), .Z(n2560) );
  IV U2200 ( .A(n2553), .Z(n2555) );
  XOR U2201 ( .A(n2562), .B(n2563), .Z(n2553) );
  AND U2202 ( .A(n671), .B(n2564), .Z(n2563) );
  XOR U2203 ( .A(n2565), .B(n2566), .Z(n2551) );
  AND U2204 ( .A(n675), .B(n2564), .Z(n2566) );
  XNOR U2205 ( .A(n2565), .B(n2562), .Z(n2564) );
  XOR U2206 ( .A(n2567), .B(n2568), .Z(n2562) );
  AND U2207 ( .A(n678), .B(n2561), .Z(n2568) );
  XNOR U2208 ( .A(n2569), .B(n2559), .Z(n2561) );
  XOR U2209 ( .A(n2570), .B(n2571), .Z(n2559) );
  AND U2210 ( .A(n682), .B(n2572), .Z(n2571) );
  XOR U2211 ( .A(p_input[935]), .B(n2570), .Z(n2572) );
  XOR U2212 ( .A(n2573), .B(n2574), .Z(n2570) );
  AND U2213 ( .A(n686), .B(n2575), .Z(n2574) );
  IV U2214 ( .A(n2567), .Z(n2569) );
  XOR U2215 ( .A(n2576), .B(n2577), .Z(n2567) );
  AND U2216 ( .A(n690), .B(n2578), .Z(n2577) );
  XOR U2217 ( .A(n2579), .B(n2580), .Z(n2565) );
  AND U2218 ( .A(n694), .B(n2578), .Z(n2580) );
  XNOR U2219 ( .A(n2579), .B(n2576), .Z(n2578) );
  XOR U2220 ( .A(n2581), .B(n2582), .Z(n2576) );
  AND U2221 ( .A(n697), .B(n2575), .Z(n2582) );
  XNOR U2222 ( .A(n2583), .B(n2573), .Z(n2575) );
  XOR U2223 ( .A(n2584), .B(n2585), .Z(n2573) );
  AND U2224 ( .A(n701), .B(n2586), .Z(n2585) );
  XOR U2225 ( .A(p_input[967]), .B(n2584), .Z(n2586) );
  XOR U2226 ( .A(n2587), .B(n2588), .Z(n2584) );
  AND U2227 ( .A(n705), .B(n2589), .Z(n2588) );
  IV U2228 ( .A(n2581), .Z(n2583) );
  XOR U2229 ( .A(n2590), .B(n2591), .Z(n2581) );
  AND U2230 ( .A(n709), .B(n2592), .Z(n2591) );
  XOR U2231 ( .A(n2593), .B(n2594), .Z(n2579) );
  AND U2232 ( .A(n713), .B(n2592), .Z(n2594) );
  XNOR U2233 ( .A(n2593), .B(n2590), .Z(n2592) );
  XOR U2234 ( .A(n2595), .B(n2596), .Z(n2590) );
  AND U2235 ( .A(n716), .B(n2589), .Z(n2596) );
  XNOR U2236 ( .A(n2597), .B(n2587), .Z(n2589) );
  XOR U2237 ( .A(n2598), .B(n2599), .Z(n2587) );
  AND U2238 ( .A(n720), .B(n2600), .Z(n2599) );
  XOR U2239 ( .A(p_input[999]), .B(n2598), .Z(n2600) );
  XOR U2240 ( .A(n2601), .B(n2602), .Z(n2598) );
  AND U2241 ( .A(n724), .B(n2603), .Z(n2602) );
  IV U2242 ( .A(n2595), .Z(n2597) );
  XOR U2243 ( .A(n2604), .B(n2605), .Z(n2595) );
  AND U2244 ( .A(n728), .B(n2606), .Z(n2605) );
  XOR U2245 ( .A(n2607), .B(n2608), .Z(n2593) );
  AND U2246 ( .A(n732), .B(n2606), .Z(n2608) );
  XNOR U2247 ( .A(n2607), .B(n2604), .Z(n2606) );
  XOR U2248 ( .A(n2609), .B(n2610), .Z(n2604) );
  AND U2249 ( .A(n735), .B(n2603), .Z(n2610) );
  XNOR U2250 ( .A(n2611), .B(n2601), .Z(n2603) );
  XOR U2251 ( .A(n2612), .B(n2613), .Z(n2601) );
  AND U2252 ( .A(n739), .B(n2614), .Z(n2613) );
  XOR U2253 ( .A(p_input[1031]), .B(n2612), .Z(n2614) );
  XOR U2254 ( .A(n2615), .B(n2616), .Z(n2612) );
  AND U2255 ( .A(n743), .B(n2617), .Z(n2616) );
  IV U2256 ( .A(n2609), .Z(n2611) );
  XOR U2257 ( .A(n2618), .B(n2619), .Z(n2609) );
  AND U2258 ( .A(n747), .B(n2620), .Z(n2619) );
  XOR U2259 ( .A(n2621), .B(n2622), .Z(n2607) );
  AND U2260 ( .A(n751), .B(n2620), .Z(n2622) );
  XNOR U2261 ( .A(n2621), .B(n2618), .Z(n2620) );
  XOR U2262 ( .A(n2623), .B(n2624), .Z(n2618) );
  AND U2263 ( .A(n754), .B(n2617), .Z(n2624) );
  XNOR U2264 ( .A(n2625), .B(n2615), .Z(n2617) );
  XOR U2265 ( .A(n2626), .B(n2627), .Z(n2615) );
  AND U2266 ( .A(n758), .B(n2628), .Z(n2627) );
  XOR U2267 ( .A(p_input[1063]), .B(n2626), .Z(n2628) );
  XOR U2268 ( .A(n2629), .B(n2630), .Z(n2626) );
  AND U2269 ( .A(n762), .B(n2631), .Z(n2630) );
  IV U2270 ( .A(n2623), .Z(n2625) );
  XOR U2271 ( .A(n2632), .B(n2633), .Z(n2623) );
  AND U2272 ( .A(n766), .B(n2634), .Z(n2633) );
  XOR U2273 ( .A(n2635), .B(n2636), .Z(n2621) );
  AND U2274 ( .A(n770), .B(n2634), .Z(n2636) );
  XNOR U2275 ( .A(n2635), .B(n2632), .Z(n2634) );
  XOR U2276 ( .A(n2637), .B(n2638), .Z(n2632) );
  AND U2277 ( .A(n773), .B(n2631), .Z(n2638) );
  XNOR U2278 ( .A(n2639), .B(n2629), .Z(n2631) );
  XOR U2279 ( .A(n2640), .B(n2641), .Z(n2629) );
  AND U2280 ( .A(n777), .B(n2642), .Z(n2641) );
  XOR U2281 ( .A(p_input[1095]), .B(n2640), .Z(n2642) );
  XOR U2282 ( .A(n2643), .B(n2644), .Z(n2640) );
  AND U2283 ( .A(n781), .B(n2645), .Z(n2644) );
  IV U2284 ( .A(n2637), .Z(n2639) );
  XOR U2285 ( .A(n2646), .B(n2647), .Z(n2637) );
  AND U2286 ( .A(n785), .B(n2648), .Z(n2647) );
  XOR U2287 ( .A(n2649), .B(n2650), .Z(n2635) );
  AND U2288 ( .A(n789), .B(n2648), .Z(n2650) );
  XNOR U2289 ( .A(n2649), .B(n2646), .Z(n2648) );
  XOR U2290 ( .A(n2651), .B(n2652), .Z(n2646) );
  AND U2291 ( .A(n792), .B(n2645), .Z(n2652) );
  XNOR U2292 ( .A(n2653), .B(n2643), .Z(n2645) );
  XOR U2293 ( .A(n2654), .B(n2655), .Z(n2643) );
  AND U2294 ( .A(n796), .B(n2656), .Z(n2655) );
  XOR U2295 ( .A(p_input[1127]), .B(n2654), .Z(n2656) );
  XOR U2296 ( .A(n2657), .B(n2658), .Z(n2654) );
  AND U2297 ( .A(n800), .B(n2659), .Z(n2658) );
  IV U2298 ( .A(n2651), .Z(n2653) );
  XOR U2299 ( .A(n2660), .B(n2661), .Z(n2651) );
  AND U2300 ( .A(n804), .B(n2662), .Z(n2661) );
  XOR U2301 ( .A(n2663), .B(n2664), .Z(n2649) );
  AND U2302 ( .A(n808), .B(n2662), .Z(n2664) );
  XNOR U2303 ( .A(n2663), .B(n2660), .Z(n2662) );
  XOR U2304 ( .A(n2665), .B(n2666), .Z(n2660) );
  AND U2305 ( .A(n811), .B(n2659), .Z(n2666) );
  XNOR U2306 ( .A(n2667), .B(n2657), .Z(n2659) );
  XOR U2307 ( .A(n2668), .B(n2669), .Z(n2657) );
  AND U2308 ( .A(n815), .B(n2670), .Z(n2669) );
  XOR U2309 ( .A(p_input[1159]), .B(n2668), .Z(n2670) );
  XOR U2310 ( .A(n2671), .B(n2672), .Z(n2668) );
  AND U2311 ( .A(n819), .B(n2673), .Z(n2672) );
  IV U2312 ( .A(n2665), .Z(n2667) );
  XOR U2313 ( .A(n2674), .B(n2675), .Z(n2665) );
  AND U2314 ( .A(n823), .B(n2676), .Z(n2675) );
  XOR U2315 ( .A(n2677), .B(n2678), .Z(n2663) );
  AND U2316 ( .A(n827), .B(n2676), .Z(n2678) );
  XNOR U2317 ( .A(n2677), .B(n2674), .Z(n2676) );
  XOR U2318 ( .A(n2679), .B(n2680), .Z(n2674) );
  AND U2319 ( .A(n830), .B(n2673), .Z(n2680) );
  XNOR U2320 ( .A(n2681), .B(n2671), .Z(n2673) );
  XOR U2321 ( .A(n2682), .B(n2683), .Z(n2671) );
  AND U2322 ( .A(n834), .B(n2684), .Z(n2683) );
  XOR U2323 ( .A(p_input[1191]), .B(n2682), .Z(n2684) );
  XOR U2324 ( .A(n2685), .B(n2686), .Z(n2682) );
  AND U2325 ( .A(n838), .B(n2687), .Z(n2686) );
  IV U2326 ( .A(n2679), .Z(n2681) );
  XOR U2327 ( .A(n2688), .B(n2689), .Z(n2679) );
  AND U2328 ( .A(n842), .B(n2690), .Z(n2689) );
  XOR U2329 ( .A(n2691), .B(n2692), .Z(n2677) );
  AND U2330 ( .A(n846), .B(n2690), .Z(n2692) );
  XNOR U2331 ( .A(n2691), .B(n2688), .Z(n2690) );
  XOR U2332 ( .A(n2693), .B(n2694), .Z(n2688) );
  AND U2333 ( .A(n849), .B(n2687), .Z(n2694) );
  XNOR U2334 ( .A(n2695), .B(n2685), .Z(n2687) );
  XOR U2335 ( .A(n2696), .B(n2697), .Z(n2685) );
  AND U2336 ( .A(n853), .B(n2698), .Z(n2697) );
  XOR U2337 ( .A(p_input[1223]), .B(n2696), .Z(n2698) );
  XOR U2338 ( .A(n2699), .B(n2700), .Z(n2696) );
  AND U2339 ( .A(n857), .B(n2701), .Z(n2700) );
  IV U2340 ( .A(n2693), .Z(n2695) );
  XOR U2341 ( .A(n2702), .B(n2703), .Z(n2693) );
  AND U2342 ( .A(n861), .B(n2704), .Z(n2703) );
  XOR U2343 ( .A(n2705), .B(n2706), .Z(n2691) );
  AND U2344 ( .A(n865), .B(n2704), .Z(n2706) );
  XNOR U2345 ( .A(n2705), .B(n2702), .Z(n2704) );
  XOR U2346 ( .A(n2707), .B(n2708), .Z(n2702) );
  AND U2347 ( .A(n868), .B(n2701), .Z(n2708) );
  XNOR U2348 ( .A(n2709), .B(n2699), .Z(n2701) );
  XOR U2349 ( .A(n2710), .B(n2711), .Z(n2699) );
  AND U2350 ( .A(n872), .B(n2712), .Z(n2711) );
  XOR U2351 ( .A(p_input[1255]), .B(n2710), .Z(n2712) );
  XOR U2352 ( .A(n2713), .B(n2714), .Z(n2710) );
  AND U2353 ( .A(n876), .B(n2715), .Z(n2714) );
  IV U2354 ( .A(n2707), .Z(n2709) );
  XOR U2355 ( .A(n2716), .B(n2717), .Z(n2707) );
  AND U2356 ( .A(n880), .B(n2718), .Z(n2717) );
  XOR U2357 ( .A(n2719), .B(n2720), .Z(n2705) );
  AND U2358 ( .A(n884), .B(n2718), .Z(n2720) );
  XNOR U2359 ( .A(n2719), .B(n2716), .Z(n2718) );
  XOR U2360 ( .A(n2721), .B(n2722), .Z(n2716) );
  AND U2361 ( .A(n887), .B(n2715), .Z(n2722) );
  XNOR U2362 ( .A(n2723), .B(n2713), .Z(n2715) );
  XOR U2363 ( .A(n2724), .B(n2725), .Z(n2713) );
  AND U2364 ( .A(n891), .B(n2726), .Z(n2725) );
  XOR U2365 ( .A(p_input[1287]), .B(n2724), .Z(n2726) );
  XOR U2366 ( .A(n2727), .B(n2728), .Z(n2724) );
  AND U2367 ( .A(n895), .B(n2729), .Z(n2728) );
  IV U2368 ( .A(n2721), .Z(n2723) );
  XOR U2369 ( .A(n2730), .B(n2731), .Z(n2721) );
  AND U2370 ( .A(n899), .B(n2732), .Z(n2731) );
  XOR U2371 ( .A(n2733), .B(n2734), .Z(n2719) );
  AND U2372 ( .A(n903), .B(n2732), .Z(n2734) );
  XNOR U2373 ( .A(n2733), .B(n2730), .Z(n2732) );
  XOR U2374 ( .A(n2735), .B(n2736), .Z(n2730) );
  AND U2375 ( .A(n906), .B(n2729), .Z(n2736) );
  XNOR U2376 ( .A(n2737), .B(n2727), .Z(n2729) );
  XOR U2377 ( .A(n2738), .B(n2739), .Z(n2727) );
  AND U2378 ( .A(n910), .B(n2740), .Z(n2739) );
  XOR U2379 ( .A(p_input[1319]), .B(n2738), .Z(n2740) );
  XOR U2380 ( .A(n2741), .B(n2742), .Z(n2738) );
  AND U2381 ( .A(n914), .B(n2743), .Z(n2742) );
  IV U2382 ( .A(n2735), .Z(n2737) );
  XOR U2383 ( .A(n2744), .B(n2745), .Z(n2735) );
  AND U2384 ( .A(n918), .B(n2746), .Z(n2745) );
  XOR U2385 ( .A(n2747), .B(n2748), .Z(n2733) );
  AND U2386 ( .A(n922), .B(n2746), .Z(n2748) );
  XNOR U2387 ( .A(n2747), .B(n2744), .Z(n2746) );
  XOR U2388 ( .A(n2749), .B(n2750), .Z(n2744) );
  AND U2389 ( .A(n925), .B(n2743), .Z(n2750) );
  XNOR U2390 ( .A(n2751), .B(n2741), .Z(n2743) );
  XOR U2391 ( .A(n2752), .B(n2753), .Z(n2741) );
  AND U2392 ( .A(n929), .B(n2754), .Z(n2753) );
  XOR U2393 ( .A(p_input[1351]), .B(n2752), .Z(n2754) );
  XOR U2394 ( .A(n2755), .B(n2756), .Z(n2752) );
  AND U2395 ( .A(n933), .B(n2757), .Z(n2756) );
  IV U2396 ( .A(n2749), .Z(n2751) );
  XOR U2397 ( .A(n2758), .B(n2759), .Z(n2749) );
  AND U2398 ( .A(n937), .B(n2760), .Z(n2759) );
  XOR U2399 ( .A(n2761), .B(n2762), .Z(n2747) );
  AND U2400 ( .A(n941), .B(n2760), .Z(n2762) );
  XNOR U2401 ( .A(n2761), .B(n2758), .Z(n2760) );
  XOR U2402 ( .A(n2763), .B(n2764), .Z(n2758) );
  AND U2403 ( .A(n944), .B(n2757), .Z(n2764) );
  XNOR U2404 ( .A(n2765), .B(n2755), .Z(n2757) );
  XOR U2405 ( .A(n2766), .B(n2767), .Z(n2755) );
  AND U2406 ( .A(n948), .B(n2768), .Z(n2767) );
  XOR U2407 ( .A(p_input[1383]), .B(n2766), .Z(n2768) );
  XOR U2408 ( .A(n2769), .B(n2770), .Z(n2766) );
  AND U2409 ( .A(n952), .B(n2771), .Z(n2770) );
  IV U2410 ( .A(n2763), .Z(n2765) );
  XOR U2411 ( .A(n2772), .B(n2773), .Z(n2763) );
  AND U2412 ( .A(n956), .B(n2774), .Z(n2773) );
  XOR U2413 ( .A(n2775), .B(n2776), .Z(n2761) );
  AND U2414 ( .A(n960), .B(n2774), .Z(n2776) );
  XNOR U2415 ( .A(n2775), .B(n2772), .Z(n2774) );
  XOR U2416 ( .A(n2777), .B(n2778), .Z(n2772) );
  AND U2417 ( .A(n963), .B(n2771), .Z(n2778) );
  XNOR U2418 ( .A(n2779), .B(n2769), .Z(n2771) );
  XOR U2419 ( .A(n2780), .B(n2781), .Z(n2769) );
  AND U2420 ( .A(n967), .B(n2782), .Z(n2781) );
  XOR U2421 ( .A(p_input[1415]), .B(n2780), .Z(n2782) );
  XOR U2422 ( .A(n2783), .B(n2784), .Z(n2780) );
  AND U2423 ( .A(n971), .B(n2785), .Z(n2784) );
  IV U2424 ( .A(n2777), .Z(n2779) );
  XOR U2425 ( .A(n2786), .B(n2787), .Z(n2777) );
  AND U2426 ( .A(n975), .B(n2788), .Z(n2787) );
  XOR U2427 ( .A(n2789), .B(n2790), .Z(n2775) );
  AND U2428 ( .A(n979), .B(n2788), .Z(n2790) );
  XNOR U2429 ( .A(n2789), .B(n2786), .Z(n2788) );
  XOR U2430 ( .A(n2791), .B(n2792), .Z(n2786) );
  AND U2431 ( .A(n982), .B(n2785), .Z(n2792) );
  XNOR U2432 ( .A(n2793), .B(n2783), .Z(n2785) );
  XOR U2433 ( .A(n2794), .B(n2795), .Z(n2783) );
  AND U2434 ( .A(n986), .B(n2796), .Z(n2795) );
  XOR U2435 ( .A(p_input[1447]), .B(n2794), .Z(n2796) );
  XOR U2436 ( .A(n2797), .B(n2798), .Z(n2794) );
  AND U2437 ( .A(n990), .B(n2799), .Z(n2798) );
  IV U2438 ( .A(n2791), .Z(n2793) );
  XOR U2439 ( .A(n2800), .B(n2801), .Z(n2791) );
  AND U2440 ( .A(n994), .B(n2802), .Z(n2801) );
  XOR U2441 ( .A(n2803), .B(n2804), .Z(n2789) );
  AND U2442 ( .A(n998), .B(n2802), .Z(n2804) );
  XNOR U2443 ( .A(n2803), .B(n2800), .Z(n2802) );
  XOR U2444 ( .A(n2805), .B(n2806), .Z(n2800) );
  AND U2445 ( .A(n1001), .B(n2799), .Z(n2806) );
  XNOR U2446 ( .A(n2807), .B(n2797), .Z(n2799) );
  XOR U2447 ( .A(n2808), .B(n2809), .Z(n2797) );
  AND U2448 ( .A(n1005), .B(n2810), .Z(n2809) );
  XOR U2449 ( .A(p_input[1479]), .B(n2808), .Z(n2810) );
  XOR U2450 ( .A(n2811), .B(n2812), .Z(n2808) );
  AND U2451 ( .A(n1009), .B(n2813), .Z(n2812) );
  IV U2452 ( .A(n2805), .Z(n2807) );
  XOR U2453 ( .A(n2814), .B(n2815), .Z(n2805) );
  AND U2454 ( .A(n1013), .B(n2816), .Z(n2815) );
  XOR U2455 ( .A(n2817), .B(n2818), .Z(n2803) );
  AND U2456 ( .A(n1017), .B(n2816), .Z(n2818) );
  XNOR U2457 ( .A(n2817), .B(n2814), .Z(n2816) );
  XOR U2458 ( .A(n2819), .B(n2820), .Z(n2814) );
  AND U2459 ( .A(n1020), .B(n2813), .Z(n2820) );
  XNOR U2460 ( .A(n2821), .B(n2811), .Z(n2813) );
  XOR U2461 ( .A(n2822), .B(n2823), .Z(n2811) );
  AND U2462 ( .A(n1024), .B(n2824), .Z(n2823) );
  XOR U2463 ( .A(p_input[1511]), .B(n2822), .Z(n2824) );
  XOR U2464 ( .A(n2825), .B(n2826), .Z(n2822) );
  AND U2465 ( .A(n1028), .B(n2827), .Z(n2826) );
  IV U2466 ( .A(n2819), .Z(n2821) );
  XOR U2467 ( .A(n2828), .B(n2829), .Z(n2819) );
  AND U2468 ( .A(n1032), .B(n2830), .Z(n2829) );
  XOR U2469 ( .A(n2831), .B(n2832), .Z(n2817) );
  AND U2470 ( .A(n1036), .B(n2830), .Z(n2832) );
  XNOR U2471 ( .A(n2831), .B(n2828), .Z(n2830) );
  XOR U2472 ( .A(n2833), .B(n2834), .Z(n2828) );
  AND U2473 ( .A(n1039), .B(n2827), .Z(n2834) );
  XNOR U2474 ( .A(n2835), .B(n2825), .Z(n2827) );
  XOR U2475 ( .A(n2836), .B(n2837), .Z(n2825) );
  AND U2476 ( .A(n1043), .B(n2838), .Z(n2837) );
  XOR U2477 ( .A(p_input[1543]), .B(n2836), .Z(n2838) );
  XOR U2478 ( .A(n2839), .B(n2840), .Z(n2836) );
  AND U2479 ( .A(n1047), .B(n2841), .Z(n2840) );
  IV U2480 ( .A(n2833), .Z(n2835) );
  XOR U2481 ( .A(n2842), .B(n2843), .Z(n2833) );
  AND U2482 ( .A(n1051), .B(n2844), .Z(n2843) );
  XOR U2483 ( .A(n2845), .B(n2846), .Z(n2831) );
  AND U2484 ( .A(n1055), .B(n2844), .Z(n2846) );
  XNOR U2485 ( .A(n2845), .B(n2842), .Z(n2844) );
  XOR U2486 ( .A(n2847), .B(n2848), .Z(n2842) );
  AND U2487 ( .A(n1058), .B(n2841), .Z(n2848) );
  XNOR U2488 ( .A(n2849), .B(n2839), .Z(n2841) );
  XOR U2489 ( .A(n2850), .B(n2851), .Z(n2839) );
  AND U2490 ( .A(n1062), .B(n2852), .Z(n2851) );
  XOR U2491 ( .A(p_input[1575]), .B(n2850), .Z(n2852) );
  XOR U2492 ( .A(n2853), .B(n2854), .Z(n2850) );
  AND U2493 ( .A(n1066), .B(n2855), .Z(n2854) );
  IV U2494 ( .A(n2847), .Z(n2849) );
  XOR U2495 ( .A(n2856), .B(n2857), .Z(n2847) );
  AND U2496 ( .A(n1070), .B(n2858), .Z(n2857) );
  XOR U2497 ( .A(n2859), .B(n2860), .Z(n2845) );
  AND U2498 ( .A(n1074), .B(n2858), .Z(n2860) );
  XNOR U2499 ( .A(n2859), .B(n2856), .Z(n2858) );
  XOR U2500 ( .A(n2861), .B(n2862), .Z(n2856) );
  AND U2501 ( .A(n1077), .B(n2855), .Z(n2862) );
  XNOR U2502 ( .A(n2863), .B(n2853), .Z(n2855) );
  XOR U2503 ( .A(n2864), .B(n2865), .Z(n2853) );
  AND U2504 ( .A(n1081), .B(n2866), .Z(n2865) );
  XOR U2505 ( .A(p_input[1607]), .B(n2864), .Z(n2866) );
  XOR U2506 ( .A(n2867), .B(n2868), .Z(n2864) );
  AND U2507 ( .A(n1085), .B(n2869), .Z(n2868) );
  IV U2508 ( .A(n2861), .Z(n2863) );
  XOR U2509 ( .A(n2870), .B(n2871), .Z(n2861) );
  AND U2510 ( .A(n1089), .B(n2872), .Z(n2871) );
  XOR U2511 ( .A(n2873), .B(n2874), .Z(n2859) );
  AND U2512 ( .A(n1093), .B(n2872), .Z(n2874) );
  XNOR U2513 ( .A(n2873), .B(n2870), .Z(n2872) );
  XOR U2514 ( .A(n2875), .B(n2876), .Z(n2870) );
  AND U2515 ( .A(n1096), .B(n2869), .Z(n2876) );
  XNOR U2516 ( .A(n2877), .B(n2867), .Z(n2869) );
  XOR U2517 ( .A(n2878), .B(n2879), .Z(n2867) );
  AND U2518 ( .A(n1100), .B(n2880), .Z(n2879) );
  XOR U2519 ( .A(p_input[1639]), .B(n2878), .Z(n2880) );
  XOR U2520 ( .A(n2881), .B(n2882), .Z(n2878) );
  AND U2521 ( .A(n1104), .B(n2883), .Z(n2882) );
  IV U2522 ( .A(n2875), .Z(n2877) );
  XOR U2523 ( .A(n2884), .B(n2885), .Z(n2875) );
  AND U2524 ( .A(n1108), .B(n2886), .Z(n2885) );
  XOR U2525 ( .A(n2887), .B(n2888), .Z(n2873) );
  AND U2526 ( .A(n1112), .B(n2886), .Z(n2888) );
  XNOR U2527 ( .A(n2887), .B(n2884), .Z(n2886) );
  XOR U2528 ( .A(n2889), .B(n2890), .Z(n2884) );
  AND U2529 ( .A(n1115), .B(n2883), .Z(n2890) );
  XNOR U2530 ( .A(n2891), .B(n2881), .Z(n2883) );
  XOR U2531 ( .A(n2892), .B(n2893), .Z(n2881) );
  AND U2532 ( .A(n1119), .B(n2894), .Z(n2893) );
  XOR U2533 ( .A(p_input[1671]), .B(n2892), .Z(n2894) );
  XOR U2534 ( .A(n2895), .B(n2896), .Z(n2892) );
  AND U2535 ( .A(n1123), .B(n2897), .Z(n2896) );
  IV U2536 ( .A(n2889), .Z(n2891) );
  XOR U2537 ( .A(n2898), .B(n2899), .Z(n2889) );
  AND U2538 ( .A(n1127), .B(n2900), .Z(n2899) );
  XOR U2539 ( .A(n2901), .B(n2902), .Z(n2887) );
  AND U2540 ( .A(n1131), .B(n2900), .Z(n2902) );
  XNOR U2541 ( .A(n2901), .B(n2898), .Z(n2900) );
  XOR U2542 ( .A(n2903), .B(n2904), .Z(n2898) );
  AND U2543 ( .A(n1134), .B(n2897), .Z(n2904) );
  XNOR U2544 ( .A(n2905), .B(n2895), .Z(n2897) );
  XOR U2545 ( .A(n2906), .B(n2907), .Z(n2895) );
  AND U2546 ( .A(n1138), .B(n2908), .Z(n2907) );
  XOR U2547 ( .A(p_input[1703]), .B(n2906), .Z(n2908) );
  XOR U2548 ( .A(n2909), .B(n2910), .Z(n2906) );
  AND U2549 ( .A(n1142), .B(n2911), .Z(n2910) );
  IV U2550 ( .A(n2903), .Z(n2905) );
  XOR U2551 ( .A(n2912), .B(n2913), .Z(n2903) );
  AND U2552 ( .A(n1146), .B(n2914), .Z(n2913) );
  XOR U2553 ( .A(n2915), .B(n2916), .Z(n2901) );
  AND U2554 ( .A(n1150), .B(n2914), .Z(n2916) );
  XNOR U2555 ( .A(n2915), .B(n2912), .Z(n2914) );
  XOR U2556 ( .A(n2917), .B(n2918), .Z(n2912) );
  AND U2557 ( .A(n1153), .B(n2911), .Z(n2918) );
  XNOR U2558 ( .A(n2919), .B(n2909), .Z(n2911) );
  XOR U2559 ( .A(n2920), .B(n2921), .Z(n2909) );
  AND U2560 ( .A(n1157), .B(n2922), .Z(n2921) );
  XOR U2561 ( .A(p_input[1735]), .B(n2920), .Z(n2922) );
  XOR U2562 ( .A(n2923), .B(n2924), .Z(n2920) );
  AND U2563 ( .A(n1161), .B(n2925), .Z(n2924) );
  IV U2564 ( .A(n2917), .Z(n2919) );
  XOR U2565 ( .A(n2926), .B(n2927), .Z(n2917) );
  AND U2566 ( .A(n1165), .B(n2928), .Z(n2927) );
  XOR U2567 ( .A(n2929), .B(n2930), .Z(n2915) );
  AND U2568 ( .A(n1169), .B(n2928), .Z(n2930) );
  XNOR U2569 ( .A(n2929), .B(n2926), .Z(n2928) );
  XOR U2570 ( .A(n2931), .B(n2932), .Z(n2926) );
  AND U2571 ( .A(n1172), .B(n2925), .Z(n2932) );
  XNOR U2572 ( .A(n2933), .B(n2923), .Z(n2925) );
  XOR U2573 ( .A(n2934), .B(n2935), .Z(n2923) );
  AND U2574 ( .A(n1176), .B(n2936), .Z(n2935) );
  XOR U2575 ( .A(p_input[1767]), .B(n2934), .Z(n2936) );
  XOR U2576 ( .A(n2937), .B(n2938), .Z(n2934) );
  AND U2577 ( .A(n1180), .B(n2939), .Z(n2938) );
  IV U2578 ( .A(n2931), .Z(n2933) );
  XOR U2579 ( .A(n2940), .B(n2941), .Z(n2931) );
  AND U2580 ( .A(n1184), .B(n2942), .Z(n2941) );
  XOR U2581 ( .A(n2943), .B(n2944), .Z(n2929) );
  AND U2582 ( .A(n1188), .B(n2942), .Z(n2944) );
  XNOR U2583 ( .A(n2943), .B(n2940), .Z(n2942) );
  XOR U2584 ( .A(n2945), .B(n2946), .Z(n2940) );
  AND U2585 ( .A(n1191), .B(n2939), .Z(n2946) );
  XNOR U2586 ( .A(n2947), .B(n2937), .Z(n2939) );
  XOR U2587 ( .A(n2948), .B(n2949), .Z(n2937) );
  AND U2588 ( .A(n1195), .B(n2950), .Z(n2949) );
  XOR U2589 ( .A(p_input[1799]), .B(n2948), .Z(n2950) );
  XOR U2590 ( .A(n2951), .B(n2952), .Z(n2948) );
  AND U2591 ( .A(n1199), .B(n2953), .Z(n2952) );
  IV U2592 ( .A(n2945), .Z(n2947) );
  XOR U2593 ( .A(n2954), .B(n2955), .Z(n2945) );
  AND U2594 ( .A(n1203), .B(n2956), .Z(n2955) );
  XOR U2595 ( .A(n2957), .B(n2958), .Z(n2943) );
  AND U2596 ( .A(n1207), .B(n2956), .Z(n2958) );
  XNOR U2597 ( .A(n2957), .B(n2954), .Z(n2956) );
  XOR U2598 ( .A(n2959), .B(n2960), .Z(n2954) );
  AND U2599 ( .A(n1210), .B(n2953), .Z(n2960) );
  XNOR U2600 ( .A(n2961), .B(n2951), .Z(n2953) );
  XOR U2601 ( .A(n2962), .B(n2963), .Z(n2951) );
  AND U2602 ( .A(n1214), .B(n2964), .Z(n2963) );
  XOR U2603 ( .A(p_input[1831]), .B(n2962), .Z(n2964) );
  XOR U2604 ( .A(n2965), .B(n2966), .Z(n2962) );
  AND U2605 ( .A(n1218), .B(n2967), .Z(n2966) );
  IV U2606 ( .A(n2959), .Z(n2961) );
  XOR U2607 ( .A(n2968), .B(n2969), .Z(n2959) );
  AND U2608 ( .A(n1222), .B(n2970), .Z(n2969) );
  XOR U2609 ( .A(n2971), .B(n2972), .Z(n2957) );
  AND U2610 ( .A(n1226), .B(n2970), .Z(n2972) );
  XNOR U2611 ( .A(n2971), .B(n2968), .Z(n2970) );
  XOR U2612 ( .A(n2973), .B(n2974), .Z(n2968) );
  AND U2613 ( .A(n1229), .B(n2967), .Z(n2974) );
  XNOR U2614 ( .A(n2975), .B(n2965), .Z(n2967) );
  XOR U2615 ( .A(n2976), .B(n2977), .Z(n2965) );
  AND U2616 ( .A(n1233), .B(n2978), .Z(n2977) );
  XOR U2617 ( .A(p_input[1863]), .B(n2976), .Z(n2978) );
  XOR U2618 ( .A(n2979), .B(n2980), .Z(n2976) );
  AND U2619 ( .A(n1237), .B(n2981), .Z(n2980) );
  IV U2620 ( .A(n2973), .Z(n2975) );
  XOR U2621 ( .A(n2982), .B(n2983), .Z(n2973) );
  AND U2622 ( .A(n1241), .B(n2984), .Z(n2983) );
  XOR U2623 ( .A(n2985), .B(n2986), .Z(n2971) );
  AND U2624 ( .A(n1245), .B(n2984), .Z(n2986) );
  XNOR U2625 ( .A(n2985), .B(n2982), .Z(n2984) );
  XOR U2626 ( .A(n2987), .B(n2988), .Z(n2982) );
  AND U2627 ( .A(n1248), .B(n2981), .Z(n2988) );
  XNOR U2628 ( .A(n2989), .B(n2979), .Z(n2981) );
  XOR U2629 ( .A(n2990), .B(n2991), .Z(n2979) );
  AND U2630 ( .A(n1252), .B(n2992), .Z(n2991) );
  XOR U2631 ( .A(p_input[1895]), .B(n2990), .Z(n2992) );
  XOR U2632 ( .A(n2993), .B(n2994), .Z(n2990) );
  AND U2633 ( .A(n1256), .B(n2995), .Z(n2994) );
  IV U2634 ( .A(n2987), .Z(n2989) );
  XOR U2635 ( .A(n2996), .B(n2997), .Z(n2987) );
  AND U2636 ( .A(n1260), .B(n2998), .Z(n2997) );
  XOR U2637 ( .A(n2999), .B(n3000), .Z(n2985) );
  AND U2638 ( .A(n1264), .B(n2998), .Z(n3000) );
  XNOR U2639 ( .A(n2999), .B(n2996), .Z(n2998) );
  XOR U2640 ( .A(n3001), .B(n3002), .Z(n2996) );
  AND U2641 ( .A(n1267), .B(n2995), .Z(n3002) );
  XNOR U2642 ( .A(n3003), .B(n2993), .Z(n2995) );
  XOR U2643 ( .A(n3004), .B(n3005), .Z(n2993) );
  AND U2644 ( .A(n1271), .B(n3006), .Z(n3005) );
  XOR U2645 ( .A(p_input[1927]), .B(n3004), .Z(n3006) );
  XOR U2646 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(n3007), 
        .Z(n3004) );
  AND U2647 ( .A(n1274), .B(n3008), .Z(n3007) );
  IV U2648 ( .A(n3001), .Z(n3003) );
  XOR U2649 ( .A(n3009), .B(n3010), .Z(n3001) );
  AND U2650 ( .A(n1278), .B(n3011), .Z(n3010) );
  XOR U2651 ( .A(n3012), .B(n3013), .Z(n2999) );
  AND U2652 ( .A(n1282), .B(n3011), .Z(n3013) );
  XNOR U2653 ( .A(n3012), .B(n3009), .Z(n3011) );
  XNOR U2654 ( .A(n3014), .B(n3015), .Z(n3009) );
  AND U2655 ( .A(n1285), .B(n3008), .Z(n3015) );
  XNOR U2656 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(n3014), 
        .Z(n3008) );
  XNOR U2657 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(n3016), 
        .Z(n3014) );
  AND U2658 ( .A(n1287), .B(n3017), .Z(n3016) );
  XNOR U2659 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n3018), .Z(n3012) );
  AND U2660 ( .A(n1290), .B(n3017), .Z(n3018) );
  XOR U2661 ( .A(n3019), .B(n3020), .Z(n3017) );
  XOR U2662 ( .A(n59), .B(n3021), .Z(o[38]) );
  AND U2663 ( .A(n122), .B(n3022), .Z(n59) );
  XOR U2664 ( .A(n60), .B(n3021), .Z(n3022) );
  XOR U2665 ( .A(n3023), .B(n57), .Z(n3021) );
  AND U2666 ( .A(n125), .B(n3024), .Z(n57) );
  XOR U2667 ( .A(n58), .B(n3023), .Z(n3024) );
  XOR U2668 ( .A(n3025), .B(n3026), .Z(n58) );
  AND U2669 ( .A(n130), .B(n3027), .Z(n3026) );
  XOR U2670 ( .A(p_input[6]), .B(n3025), .Z(n3027) );
  XNOR U2671 ( .A(n3028), .B(n3029), .Z(n3025) );
  AND U2672 ( .A(n134), .B(n3030), .Z(n3029) );
  XOR U2673 ( .A(n3031), .B(n3032), .Z(n3023) );
  AND U2674 ( .A(n138), .B(n3033), .Z(n3032) );
  XOR U2675 ( .A(n3034), .B(n3035), .Z(n60) );
  AND U2676 ( .A(n142), .B(n3033), .Z(n3035) );
  XNOR U2677 ( .A(n3036), .B(n3034), .Z(n3033) );
  IV U2678 ( .A(n3031), .Z(n3036) );
  XOR U2679 ( .A(n3037), .B(n3038), .Z(n3031) );
  AND U2680 ( .A(n146), .B(n3030), .Z(n3038) );
  XNOR U2681 ( .A(n3028), .B(n3037), .Z(n3030) );
  XNOR U2682 ( .A(n3039), .B(n3040), .Z(n3028) );
  AND U2683 ( .A(n150), .B(n3041), .Z(n3040) );
  XOR U2684 ( .A(p_input[38]), .B(n3039), .Z(n3041) );
  XNOR U2685 ( .A(n3042), .B(n3043), .Z(n3039) );
  AND U2686 ( .A(n154), .B(n3044), .Z(n3043) );
  XOR U2687 ( .A(n3045), .B(n3046), .Z(n3037) );
  AND U2688 ( .A(n158), .B(n3047), .Z(n3046) );
  XOR U2689 ( .A(n3048), .B(n3049), .Z(n3034) );
  AND U2690 ( .A(n162), .B(n3047), .Z(n3049) );
  XNOR U2691 ( .A(n3050), .B(n3048), .Z(n3047) );
  IV U2692 ( .A(n3045), .Z(n3050) );
  XOR U2693 ( .A(n3051), .B(n3052), .Z(n3045) );
  AND U2694 ( .A(n165), .B(n3044), .Z(n3052) );
  XNOR U2695 ( .A(n3042), .B(n3051), .Z(n3044) );
  XNOR U2696 ( .A(n3053), .B(n3054), .Z(n3042) );
  AND U2697 ( .A(n169), .B(n3055), .Z(n3054) );
  XOR U2698 ( .A(p_input[70]), .B(n3053), .Z(n3055) );
  XNOR U2699 ( .A(n3056), .B(n3057), .Z(n3053) );
  AND U2700 ( .A(n173), .B(n3058), .Z(n3057) );
  XOR U2701 ( .A(n3059), .B(n3060), .Z(n3051) );
  AND U2702 ( .A(n177), .B(n3061), .Z(n3060) );
  XOR U2703 ( .A(n3062), .B(n3063), .Z(n3048) );
  AND U2704 ( .A(n181), .B(n3061), .Z(n3063) );
  XNOR U2705 ( .A(n3064), .B(n3062), .Z(n3061) );
  IV U2706 ( .A(n3059), .Z(n3064) );
  XOR U2707 ( .A(n3065), .B(n3066), .Z(n3059) );
  AND U2708 ( .A(n184), .B(n3058), .Z(n3066) );
  XNOR U2709 ( .A(n3056), .B(n3065), .Z(n3058) );
  XNOR U2710 ( .A(n3067), .B(n3068), .Z(n3056) );
  AND U2711 ( .A(n188), .B(n3069), .Z(n3068) );
  XOR U2712 ( .A(p_input[102]), .B(n3067), .Z(n3069) );
  XNOR U2713 ( .A(n3070), .B(n3071), .Z(n3067) );
  AND U2714 ( .A(n192), .B(n3072), .Z(n3071) );
  XOR U2715 ( .A(n3073), .B(n3074), .Z(n3065) );
  AND U2716 ( .A(n196), .B(n3075), .Z(n3074) );
  XOR U2717 ( .A(n3076), .B(n3077), .Z(n3062) );
  AND U2718 ( .A(n200), .B(n3075), .Z(n3077) );
  XNOR U2719 ( .A(n3078), .B(n3076), .Z(n3075) );
  IV U2720 ( .A(n3073), .Z(n3078) );
  XOR U2721 ( .A(n3079), .B(n3080), .Z(n3073) );
  AND U2722 ( .A(n203), .B(n3072), .Z(n3080) );
  XNOR U2723 ( .A(n3070), .B(n3079), .Z(n3072) );
  XNOR U2724 ( .A(n3081), .B(n3082), .Z(n3070) );
  AND U2725 ( .A(n207), .B(n3083), .Z(n3082) );
  XOR U2726 ( .A(p_input[134]), .B(n3081), .Z(n3083) );
  XNOR U2727 ( .A(n3084), .B(n3085), .Z(n3081) );
  AND U2728 ( .A(n211), .B(n3086), .Z(n3085) );
  XOR U2729 ( .A(n3087), .B(n3088), .Z(n3079) );
  AND U2730 ( .A(n215), .B(n3089), .Z(n3088) );
  XOR U2731 ( .A(n3090), .B(n3091), .Z(n3076) );
  AND U2732 ( .A(n219), .B(n3089), .Z(n3091) );
  XNOR U2733 ( .A(n3092), .B(n3090), .Z(n3089) );
  IV U2734 ( .A(n3087), .Z(n3092) );
  XOR U2735 ( .A(n3093), .B(n3094), .Z(n3087) );
  AND U2736 ( .A(n222), .B(n3086), .Z(n3094) );
  XNOR U2737 ( .A(n3084), .B(n3093), .Z(n3086) );
  XNOR U2738 ( .A(n3095), .B(n3096), .Z(n3084) );
  AND U2739 ( .A(n226), .B(n3097), .Z(n3096) );
  XOR U2740 ( .A(p_input[166]), .B(n3095), .Z(n3097) );
  XNOR U2741 ( .A(n3098), .B(n3099), .Z(n3095) );
  AND U2742 ( .A(n230), .B(n3100), .Z(n3099) );
  XOR U2743 ( .A(n3101), .B(n3102), .Z(n3093) );
  AND U2744 ( .A(n234), .B(n3103), .Z(n3102) );
  XOR U2745 ( .A(n3104), .B(n3105), .Z(n3090) );
  AND U2746 ( .A(n238), .B(n3103), .Z(n3105) );
  XNOR U2747 ( .A(n3106), .B(n3104), .Z(n3103) );
  IV U2748 ( .A(n3101), .Z(n3106) );
  XOR U2749 ( .A(n3107), .B(n3108), .Z(n3101) );
  AND U2750 ( .A(n241), .B(n3100), .Z(n3108) );
  XNOR U2751 ( .A(n3098), .B(n3107), .Z(n3100) );
  XNOR U2752 ( .A(n3109), .B(n3110), .Z(n3098) );
  AND U2753 ( .A(n245), .B(n3111), .Z(n3110) );
  XOR U2754 ( .A(p_input[198]), .B(n3109), .Z(n3111) );
  XNOR U2755 ( .A(n3112), .B(n3113), .Z(n3109) );
  AND U2756 ( .A(n249), .B(n3114), .Z(n3113) );
  XOR U2757 ( .A(n3115), .B(n3116), .Z(n3107) );
  AND U2758 ( .A(n253), .B(n3117), .Z(n3116) );
  XOR U2759 ( .A(n3118), .B(n3119), .Z(n3104) );
  AND U2760 ( .A(n257), .B(n3117), .Z(n3119) );
  XNOR U2761 ( .A(n3120), .B(n3118), .Z(n3117) );
  IV U2762 ( .A(n3115), .Z(n3120) );
  XOR U2763 ( .A(n3121), .B(n3122), .Z(n3115) );
  AND U2764 ( .A(n260), .B(n3114), .Z(n3122) );
  XNOR U2765 ( .A(n3112), .B(n3121), .Z(n3114) );
  XNOR U2766 ( .A(n3123), .B(n3124), .Z(n3112) );
  AND U2767 ( .A(n264), .B(n3125), .Z(n3124) );
  XOR U2768 ( .A(p_input[230]), .B(n3123), .Z(n3125) );
  XNOR U2769 ( .A(n3126), .B(n3127), .Z(n3123) );
  AND U2770 ( .A(n268), .B(n3128), .Z(n3127) );
  XOR U2771 ( .A(n3129), .B(n3130), .Z(n3121) );
  AND U2772 ( .A(n272), .B(n3131), .Z(n3130) );
  XOR U2773 ( .A(n3132), .B(n3133), .Z(n3118) );
  AND U2774 ( .A(n276), .B(n3131), .Z(n3133) );
  XNOR U2775 ( .A(n3134), .B(n3132), .Z(n3131) );
  IV U2776 ( .A(n3129), .Z(n3134) );
  XOR U2777 ( .A(n3135), .B(n3136), .Z(n3129) );
  AND U2778 ( .A(n279), .B(n3128), .Z(n3136) );
  XNOR U2779 ( .A(n3126), .B(n3135), .Z(n3128) );
  XNOR U2780 ( .A(n3137), .B(n3138), .Z(n3126) );
  AND U2781 ( .A(n283), .B(n3139), .Z(n3138) );
  XOR U2782 ( .A(p_input[262]), .B(n3137), .Z(n3139) );
  XNOR U2783 ( .A(n3140), .B(n3141), .Z(n3137) );
  AND U2784 ( .A(n287), .B(n3142), .Z(n3141) );
  XOR U2785 ( .A(n3143), .B(n3144), .Z(n3135) );
  AND U2786 ( .A(n291), .B(n3145), .Z(n3144) );
  XOR U2787 ( .A(n3146), .B(n3147), .Z(n3132) );
  AND U2788 ( .A(n295), .B(n3145), .Z(n3147) );
  XNOR U2789 ( .A(n3148), .B(n3146), .Z(n3145) );
  IV U2790 ( .A(n3143), .Z(n3148) );
  XOR U2791 ( .A(n3149), .B(n3150), .Z(n3143) );
  AND U2792 ( .A(n298), .B(n3142), .Z(n3150) );
  XNOR U2793 ( .A(n3140), .B(n3149), .Z(n3142) );
  XNOR U2794 ( .A(n3151), .B(n3152), .Z(n3140) );
  AND U2795 ( .A(n302), .B(n3153), .Z(n3152) );
  XOR U2796 ( .A(p_input[294]), .B(n3151), .Z(n3153) );
  XNOR U2797 ( .A(n3154), .B(n3155), .Z(n3151) );
  AND U2798 ( .A(n306), .B(n3156), .Z(n3155) );
  XOR U2799 ( .A(n3157), .B(n3158), .Z(n3149) );
  AND U2800 ( .A(n310), .B(n3159), .Z(n3158) );
  XOR U2801 ( .A(n3160), .B(n3161), .Z(n3146) );
  AND U2802 ( .A(n314), .B(n3159), .Z(n3161) );
  XNOR U2803 ( .A(n3162), .B(n3160), .Z(n3159) );
  IV U2804 ( .A(n3157), .Z(n3162) );
  XOR U2805 ( .A(n3163), .B(n3164), .Z(n3157) );
  AND U2806 ( .A(n317), .B(n3156), .Z(n3164) );
  XNOR U2807 ( .A(n3154), .B(n3163), .Z(n3156) );
  XNOR U2808 ( .A(n3165), .B(n3166), .Z(n3154) );
  AND U2809 ( .A(n321), .B(n3167), .Z(n3166) );
  XOR U2810 ( .A(p_input[326]), .B(n3165), .Z(n3167) );
  XNOR U2811 ( .A(n3168), .B(n3169), .Z(n3165) );
  AND U2812 ( .A(n325), .B(n3170), .Z(n3169) );
  XOR U2813 ( .A(n3171), .B(n3172), .Z(n3163) );
  AND U2814 ( .A(n329), .B(n3173), .Z(n3172) );
  XOR U2815 ( .A(n3174), .B(n3175), .Z(n3160) );
  AND U2816 ( .A(n333), .B(n3173), .Z(n3175) );
  XNOR U2817 ( .A(n3176), .B(n3174), .Z(n3173) );
  IV U2818 ( .A(n3171), .Z(n3176) );
  XOR U2819 ( .A(n3177), .B(n3178), .Z(n3171) );
  AND U2820 ( .A(n336), .B(n3170), .Z(n3178) );
  XNOR U2821 ( .A(n3168), .B(n3177), .Z(n3170) );
  XNOR U2822 ( .A(n3179), .B(n3180), .Z(n3168) );
  AND U2823 ( .A(n340), .B(n3181), .Z(n3180) );
  XOR U2824 ( .A(p_input[358]), .B(n3179), .Z(n3181) );
  XNOR U2825 ( .A(n3182), .B(n3183), .Z(n3179) );
  AND U2826 ( .A(n344), .B(n3184), .Z(n3183) );
  XOR U2827 ( .A(n3185), .B(n3186), .Z(n3177) );
  AND U2828 ( .A(n348), .B(n3187), .Z(n3186) );
  XOR U2829 ( .A(n3188), .B(n3189), .Z(n3174) );
  AND U2830 ( .A(n352), .B(n3187), .Z(n3189) );
  XNOR U2831 ( .A(n3190), .B(n3188), .Z(n3187) );
  IV U2832 ( .A(n3185), .Z(n3190) );
  XOR U2833 ( .A(n3191), .B(n3192), .Z(n3185) );
  AND U2834 ( .A(n355), .B(n3184), .Z(n3192) );
  XNOR U2835 ( .A(n3182), .B(n3191), .Z(n3184) );
  XNOR U2836 ( .A(n3193), .B(n3194), .Z(n3182) );
  AND U2837 ( .A(n359), .B(n3195), .Z(n3194) );
  XOR U2838 ( .A(p_input[390]), .B(n3193), .Z(n3195) );
  XNOR U2839 ( .A(n3196), .B(n3197), .Z(n3193) );
  AND U2840 ( .A(n363), .B(n3198), .Z(n3197) );
  XOR U2841 ( .A(n3199), .B(n3200), .Z(n3191) );
  AND U2842 ( .A(n367), .B(n3201), .Z(n3200) );
  XOR U2843 ( .A(n3202), .B(n3203), .Z(n3188) );
  AND U2844 ( .A(n371), .B(n3201), .Z(n3203) );
  XNOR U2845 ( .A(n3204), .B(n3202), .Z(n3201) );
  IV U2846 ( .A(n3199), .Z(n3204) );
  XOR U2847 ( .A(n3205), .B(n3206), .Z(n3199) );
  AND U2848 ( .A(n374), .B(n3198), .Z(n3206) );
  XNOR U2849 ( .A(n3196), .B(n3205), .Z(n3198) );
  XNOR U2850 ( .A(n3207), .B(n3208), .Z(n3196) );
  AND U2851 ( .A(n378), .B(n3209), .Z(n3208) );
  XOR U2852 ( .A(p_input[422]), .B(n3207), .Z(n3209) );
  XNOR U2853 ( .A(n3210), .B(n3211), .Z(n3207) );
  AND U2854 ( .A(n382), .B(n3212), .Z(n3211) );
  XOR U2855 ( .A(n3213), .B(n3214), .Z(n3205) );
  AND U2856 ( .A(n386), .B(n3215), .Z(n3214) );
  XOR U2857 ( .A(n3216), .B(n3217), .Z(n3202) );
  AND U2858 ( .A(n390), .B(n3215), .Z(n3217) );
  XNOR U2859 ( .A(n3218), .B(n3216), .Z(n3215) );
  IV U2860 ( .A(n3213), .Z(n3218) );
  XOR U2861 ( .A(n3219), .B(n3220), .Z(n3213) );
  AND U2862 ( .A(n393), .B(n3212), .Z(n3220) );
  XNOR U2863 ( .A(n3210), .B(n3219), .Z(n3212) );
  XNOR U2864 ( .A(n3221), .B(n3222), .Z(n3210) );
  AND U2865 ( .A(n397), .B(n3223), .Z(n3222) );
  XOR U2866 ( .A(p_input[454]), .B(n3221), .Z(n3223) );
  XNOR U2867 ( .A(n3224), .B(n3225), .Z(n3221) );
  AND U2868 ( .A(n401), .B(n3226), .Z(n3225) );
  XOR U2869 ( .A(n3227), .B(n3228), .Z(n3219) );
  AND U2870 ( .A(n405), .B(n3229), .Z(n3228) );
  XOR U2871 ( .A(n3230), .B(n3231), .Z(n3216) );
  AND U2872 ( .A(n409), .B(n3229), .Z(n3231) );
  XNOR U2873 ( .A(n3232), .B(n3230), .Z(n3229) );
  IV U2874 ( .A(n3227), .Z(n3232) );
  XOR U2875 ( .A(n3233), .B(n3234), .Z(n3227) );
  AND U2876 ( .A(n412), .B(n3226), .Z(n3234) );
  XNOR U2877 ( .A(n3224), .B(n3233), .Z(n3226) );
  XNOR U2878 ( .A(n3235), .B(n3236), .Z(n3224) );
  AND U2879 ( .A(n416), .B(n3237), .Z(n3236) );
  XOR U2880 ( .A(p_input[486]), .B(n3235), .Z(n3237) );
  XNOR U2881 ( .A(n3238), .B(n3239), .Z(n3235) );
  AND U2882 ( .A(n420), .B(n3240), .Z(n3239) );
  XOR U2883 ( .A(n3241), .B(n3242), .Z(n3233) );
  AND U2884 ( .A(n424), .B(n3243), .Z(n3242) );
  XOR U2885 ( .A(n3244), .B(n3245), .Z(n3230) );
  AND U2886 ( .A(n428), .B(n3243), .Z(n3245) );
  XNOR U2887 ( .A(n3246), .B(n3244), .Z(n3243) );
  IV U2888 ( .A(n3241), .Z(n3246) );
  XOR U2889 ( .A(n3247), .B(n3248), .Z(n3241) );
  AND U2890 ( .A(n431), .B(n3240), .Z(n3248) );
  XNOR U2891 ( .A(n3238), .B(n3247), .Z(n3240) );
  XNOR U2892 ( .A(n3249), .B(n3250), .Z(n3238) );
  AND U2893 ( .A(n435), .B(n3251), .Z(n3250) );
  XOR U2894 ( .A(p_input[518]), .B(n3249), .Z(n3251) );
  XNOR U2895 ( .A(n3252), .B(n3253), .Z(n3249) );
  AND U2896 ( .A(n439), .B(n3254), .Z(n3253) );
  XOR U2897 ( .A(n3255), .B(n3256), .Z(n3247) );
  AND U2898 ( .A(n443), .B(n3257), .Z(n3256) );
  XOR U2899 ( .A(n3258), .B(n3259), .Z(n3244) );
  AND U2900 ( .A(n447), .B(n3257), .Z(n3259) );
  XNOR U2901 ( .A(n3260), .B(n3258), .Z(n3257) );
  IV U2902 ( .A(n3255), .Z(n3260) );
  XOR U2903 ( .A(n3261), .B(n3262), .Z(n3255) );
  AND U2904 ( .A(n450), .B(n3254), .Z(n3262) );
  XNOR U2905 ( .A(n3252), .B(n3261), .Z(n3254) );
  XNOR U2906 ( .A(n3263), .B(n3264), .Z(n3252) );
  AND U2907 ( .A(n454), .B(n3265), .Z(n3264) );
  XOR U2908 ( .A(p_input[550]), .B(n3263), .Z(n3265) );
  XNOR U2909 ( .A(n3266), .B(n3267), .Z(n3263) );
  AND U2910 ( .A(n458), .B(n3268), .Z(n3267) );
  XOR U2911 ( .A(n3269), .B(n3270), .Z(n3261) );
  AND U2912 ( .A(n462), .B(n3271), .Z(n3270) );
  XOR U2913 ( .A(n3272), .B(n3273), .Z(n3258) );
  AND U2914 ( .A(n466), .B(n3271), .Z(n3273) );
  XNOR U2915 ( .A(n3274), .B(n3272), .Z(n3271) );
  IV U2916 ( .A(n3269), .Z(n3274) );
  XOR U2917 ( .A(n3275), .B(n3276), .Z(n3269) );
  AND U2918 ( .A(n469), .B(n3268), .Z(n3276) );
  XNOR U2919 ( .A(n3266), .B(n3275), .Z(n3268) );
  XNOR U2920 ( .A(n3277), .B(n3278), .Z(n3266) );
  AND U2921 ( .A(n473), .B(n3279), .Z(n3278) );
  XOR U2922 ( .A(p_input[582]), .B(n3277), .Z(n3279) );
  XNOR U2923 ( .A(n3280), .B(n3281), .Z(n3277) );
  AND U2924 ( .A(n477), .B(n3282), .Z(n3281) );
  XOR U2925 ( .A(n3283), .B(n3284), .Z(n3275) );
  AND U2926 ( .A(n481), .B(n3285), .Z(n3284) );
  XOR U2927 ( .A(n3286), .B(n3287), .Z(n3272) );
  AND U2928 ( .A(n485), .B(n3285), .Z(n3287) );
  XNOR U2929 ( .A(n3288), .B(n3286), .Z(n3285) );
  IV U2930 ( .A(n3283), .Z(n3288) );
  XOR U2931 ( .A(n3289), .B(n3290), .Z(n3283) );
  AND U2932 ( .A(n488), .B(n3282), .Z(n3290) );
  XNOR U2933 ( .A(n3280), .B(n3289), .Z(n3282) );
  XNOR U2934 ( .A(n3291), .B(n3292), .Z(n3280) );
  AND U2935 ( .A(n492), .B(n3293), .Z(n3292) );
  XOR U2936 ( .A(p_input[614]), .B(n3291), .Z(n3293) );
  XNOR U2937 ( .A(n3294), .B(n3295), .Z(n3291) );
  AND U2938 ( .A(n496), .B(n3296), .Z(n3295) );
  XOR U2939 ( .A(n3297), .B(n3298), .Z(n3289) );
  AND U2940 ( .A(n500), .B(n3299), .Z(n3298) );
  XOR U2941 ( .A(n3300), .B(n3301), .Z(n3286) );
  AND U2942 ( .A(n504), .B(n3299), .Z(n3301) );
  XNOR U2943 ( .A(n3302), .B(n3300), .Z(n3299) );
  IV U2944 ( .A(n3297), .Z(n3302) );
  XOR U2945 ( .A(n3303), .B(n3304), .Z(n3297) );
  AND U2946 ( .A(n507), .B(n3296), .Z(n3304) );
  XNOR U2947 ( .A(n3294), .B(n3303), .Z(n3296) );
  XNOR U2948 ( .A(n3305), .B(n3306), .Z(n3294) );
  AND U2949 ( .A(n511), .B(n3307), .Z(n3306) );
  XOR U2950 ( .A(p_input[646]), .B(n3305), .Z(n3307) );
  XNOR U2951 ( .A(n3308), .B(n3309), .Z(n3305) );
  AND U2952 ( .A(n515), .B(n3310), .Z(n3309) );
  XOR U2953 ( .A(n3311), .B(n3312), .Z(n3303) );
  AND U2954 ( .A(n519), .B(n3313), .Z(n3312) );
  XOR U2955 ( .A(n3314), .B(n3315), .Z(n3300) );
  AND U2956 ( .A(n523), .B(n3313), .Z(n3315) );
  XNOR U2957 ( .A(n3316), .B(n3314), .Z(n3313) );
  IV U2958 ( .A(n3311), .Z(n3316) );
  XOR U2959 ( .A(n3317), .B(n3318), .Z(n3311) );
  AND U2960 ( .A(n526), .B(n3310), .Z(n3318) );
  XNOR U2961 ( .A(n3308), .B(n3317), .Z(n3310) );
  XNOR U2962 ( .A(n3319), .B(n3320), .Z(n3308) );
  AND U2963 ( .A(n530), .B(n3321), .Z(n3320) );
  XOR U2964 ( .A(p_input[678]), .B(n3319), .Z(n3321) );
  XNOR U2965 ( .A(n3322), .B(n3323), .Z(n3319) );
  AND U2966 ( .A(n534), .B(n3324), .Z(n3323) );
  XOR U2967 ( .A(n3325), .B(n3326), .Z(n3317) );
  AND U2968 ( .A(n538), .B(n3327), .Z(n3326) );
  XOR U2969 ( .A(n3328), .B(n3329), .Z(n3314) );
  AND U2970 ( .A(n542), .B(n3327), .Z(n3329) );
  XNOR U2971 ( .A(n3330), .B(n3328), .Z(n3327) );
  IV U2972 ( .A(n3325), .Z(n3330) );
  XOR U2973 ( .A(n3331), .B(n3332), .Z(n3325) );
  AND U2974 ( .A(n545), .B(n3324), .Z(n3332) );
  XNOR U2975 ( .A(n3322), .B(n3331), .Z(n3324) );
  XNOR U2976 ( .A(n3333), .B(n3334), .Z(n3322) );
  AND U2977 ( .A(n549), .B(n3335), .Z(n3334) );
  XOR U2978 ( .A(p_input[710]), .B(n3333), .Z(n3335) );
  XNOR U2979 ( .A(n3336), .B(n3337), .Z(n3333) );
  AND U2980 ( .A(n553), .B(n3338), .Z(n3337) );
  XOR U2981 ( .A(n3339), .B(n3340), .Z(n3331) );
  AND U2982 ( .A(n557), .B(n3341), .Z(n3340) );
  XOR U2983 ( .A(n3342), .B(n3343), .Z(n3328) );
  AND U2984 ( .A(n561), .B(n3341), .Z(n3343) );
  XNOR U2985 ( .A(n3344), .B(n3342), .Z(n3341) );
  IV U2986 ( .A(n3339), .Z(n3344) );
  XOR U2987 ( .A(n3345), .B(n3346), .Z(n3339) );
  AND U2988 ( .A(n564), .B(n3338), .Z(n3346) );
  XNOR U2989 ( .A(n3336), .B(n3345), .Z(n3338) );
  XNOR U2990 ( .A(n3347), .B(n3348), .Z(n3336) );
  AND U2991 ( .A(n568), .B(n3349), .Z(n3348) );
  XOR U2992 ( .A(p_input[742]), .B(n3347), .Z(n3349) );
  XNOR U2993 ( .A(n3350), .B(n3351), .Z(n3347) );
  AND U2994 ( .A(n572), .B(n3352), .Z(n3351) );
  XOR U2995 ( .A(n3353), .B(n3354), .Z(n3345) );
  AND U2996 ( .A(n576), .B(n3355), .Z(n3354) );
  XOR U2997 ( .A(n3356), .B(n3357), .Z(n3342) );
  AND U2998 ( .A(n580), .B(n3355), .Z(n3357) );
  XNOR U2999 ( .A(n3358), .B(n3356), .Z(n3355) );
  IV U3000 ( .A(n3353), .Z(n3358) );
  XOR U3001 ( .A(n3359), .B(n3360), .Z(n3353) );
  AND U3002 ( .A(n583), .B(n3352), .Z(n3360) );
  XNOR U3003 ( .A(n3350), .B(n3359), .Z(n3352) );
  XNOR U3004 ( .A(n3361), .B(n3362), .Z(n3350) );
  AND U3005 ( .A(n587), .B(n3363), .Z(n3362) );
  XOR U3006 ( .A(p_input[774]), .B(n3361), .Z(n3363) );
  XNOR U3007 ( .A(n3364), .B(n3365), .Z(n3361) );
  AND U3008 ( .A(n591), .B(n3366), .Z(n3365) );
  XOR U3009 ( .A(n3367), .B(n3368), .Z(n3359) );
  AND U3010 ( .A(n595), .B(n3369), .Z(n3368) );
  XOR U3011 ( .A(n3370), .B(n3371), .Z(n3356) );
  AND U3012 ( .A(n599), .B(n3369), .Z(n3371) );
  XNOR U3013 ( .A(n3372), .B(n3370), .Z(n3369) );
  IV U3014 ( .A(n3367), .Z(n3372) );
  XOR U3015 ( .A(n3373), .B(n3374), .Z(n3367) );
  AND U3016 ( .A(n602), .B(n3366), .Z(n3374) );
  XNOR U3017 ( .A(n3364), .B(n3373), .Z(n3366) );
  XNOR U3018 ( .A(n3375), .B(n3376), .Z(n3364) );
  AND U3019 ( .A(n606), .B(n3377), .Z(n3376) );
  XOR U3020 ( .A(p_input[806]), .B(n3375), .Z(n3377) );
  XNOR U3021 ( .A(n3378), .B(n3379), .Z(n3375) );
  AND U3022 ( .A(n610), .B(n3380), .Z(n3379) );
  XOR U3023 ( .A(n3381), .B(n3382), .Z(n3373) );
  AND U3024 ( .A(n614), .B(n3383), .Z(n3382) );
  XOR U3025 ( .A(n3384), .B(n3385), .Z(n3370) );
  AND U3026 ( .A(n618), .B(n3383), .Z(n3385) );
  XNOR U3027 ( .A(n3386), .B(n3384), .Z(n3383) );
  IV U3028 ( .A(n3381), .Z(n3386) );
  XOR U3029 ( .A(n3387), .B(n3388), .Z(n3381) );
  AND U3030 ( .A(n621), .B(n3380), .Z(n3388) );
  XNOR U3031 ( .A(n3378), .B(n3387), .Z(n3380) );
  XNOR U3032 ( .A(n3389), .B(n3390), .Z(n3378) );
  AND U3033 ( .A(n625), .B(n3391), .Z(n3390) );
  XOR U3034 ( .A(p_input[838]), .B(n3389), .Z(n3391) );
  XNOR U3035 ( .A(n3392), .B(n3393), .Z(n3389) );
  AND U3036 ( .A(n629), .B(n3394), .Z(n3393) );
  XOR U3037 ( .A(n3395), .B(n3396), .Z(n3387) );
  AND U3038 ( .A(n633), .B(n3397), .Z(n3396) );
  XOR U3039 ( .A(n3398), .B(n3399), .Z(n3384) );
  AND U3040 ( .A(n637), .B(n3397), .Z(n3399) );
  XNOR U3041 ( .A(n3400), .B(n3398), .Z(n3397) );
  IV U3042 ( .A(n3395), .Z(n3400) );
  XOR U3043 ( .A(n3401), .B(n3402), .Z(n3395) );
  AND U3044 ( .A(n640), .B(n3394), .Z(n3402) );
  XNOR U3045 ( .A(n3392), .B(n3401), .Z(n3394) );
  XNOR U3046 ( .A(n3403), .B(n3404), .Z(n3392) );
  AND U3047 ( .A(n644), .B(n3405), .Z(n3404) );
  XOR U3048 ( .A(p_input[870]), .B(n3403), .Z(n3405) );
  XNOR U3049 ( .A(n3406), .B(n3407), .Z(n3403) );
  AND U3050 ( .A(n648), .B(n3408), .Z(n3407) );
  XOR U3051 ( .A(n3409), .B(n3410), .Z(n3401) );
  AND U3052 ( .A(n652), .B(n3411), .Z(n3410) );
  XOR U3053 ( .A(n3412), .B(n3413), .Z(n3398) );
  AND U3054 ( .A(n656), .B(n3411), .Z(n3413) );
  XNOR U3055 ( .A(n3414), .B(n3412), .Z(n3411) );
  IV U3056 ( .A(n3409), .Z(n3414) );
  XOR U3057 ( .A(n3415), .B(n3416), .Z(n3409) );
  AND U3058 ( .A(n659), .B(n3408), .Z(n3416) );
  XNOR U3059 ( .A(n3406), .B(n3415), .Z(n3408) );
  XNOR U3060 ( .A(n3417), .B(n3418), .Z(n3406) );
  AND U3061 ( .A(n663), .B(n3419), .Z(n3418) );
  XOR U3062 ( .A(p_input[902]), .B(n3417), .Z(n3419) );
  XNOR U3063 ( .A(n3420), .B(n3421), .Z(n3417) );
  AND U3064 ( .A(n667), .B(n3422), .Z(n3421) );
  XOR U3065 ( .A(n3423), .B(n3424), .Z(n3415) );
  AND U3066 ( .A(n671), .B(n3425), .Z(n3424) );
  XOR U3067 ( .A(n3426), .B(n3427), .Z(n3412) );
  AND U3068 ( .A(n675), .B(n3425), .Z(n3427) );
  XNOR U3069 ( .A(n3428), .B(n3426), .Z(n3425) );
  IV U3070 ( .A(n3423), .Z(n3428) );
  XOR U3071 ( .A(n3429), .B(n3430), .Z(n3423) );
  AND U3072 ( .A(n678), .B(n3422), .Z(n3430) );
  XNOR U3073 ( .A(n3420), .B(n3429), .Z(n3422) );
  XNOR U3074 ( .A(n3431), .B(n3432), .Z(n3420) );
  AND U3075 ( .A(n682), .B(n3433), .Z(n3432) );
  XOR U3076 ( .A(p_input[934]), .B(n3431), .Z(n3433) );
  XNOR U3077 ( .A(n3434), .B(n3435), .Z(n3431) );
  AND U3078 ( .A(n686), .B(n3436), .Z(n3435) );
  XOR U3079 ( .A(n3437), .B(n3438), .Z(n3429) );
  AND U3080 ( .A(n690), .B(n3439), .Z(n3438) );
  XOR U3081 ( .A(n3440), .B(n3441), .Z(n3426) );
  AND U3082 ( .A(n694), .B(n3439), .Z(n3441) );
  XNOR U3083 ( .A(n3442), .B(n3440), .Z(n3439) );
  IV U3084 ( .A(n3437), .Z(n3442) );
  XOR U3085 ( .A(n3443), .B(n3444), .Z(n3437) );
  AND U3086 ( .A(n697), .B(n3436), .Z(n3444) );
  XNOR U3087 ( .A(n3434), .B(n3443), .Z(n3436) );
  XNOR U3088 ( .A(n3445), .B(n3446), .Z(n3434) );
  AND U3089 ( .A(n701), .B(n3447), .Z(n3446) );
  XOR U3090 ( .A(p_input[966]), .B(n3445), .Z(n3447) );
  XNOR U3091 ( .A(n3448), .B(n3449), .Z(n3445) );
  AND U3092 ( .A(n705), .B(n3450), .Z(n3449) );
  XOR U3093 ( .A(n3451), .B(n3452), .Z(n3443) );
  AND U3094 ( .A(n709), .B(n3453), .Z(n3452) );
  XOR U3095 ( .A(n3454), .B(n3455), .Z(n3440) );
  AND U3096 ( .A(n713), .B(n3453), .Z(n3455) );
  XNOR U3097 ( .A(n3456), .B(n3454), .Z(n3453) );
  IV U3098 ( .A(n3451), .Z(n3456) );
  XOR U3099 ( .A(n3457), .B(n3458), .Z(n3451) );
  AND U3100 ( .A(n716), .B(n3450), .Z(n3458) );
  XNOR U3101 ( .A(n3448), .B(n3457), .Z(n3450) );
  XNOR U3102 ( .A(n3459), .B(n3460), .Z(n3448) );
  AND U3103 ( .A(n720), .B(n3461), .Z(n3460) );
  XOR U3104 ( .A(p_input[998]), .B(n3459), .Z(n3461) );
  XNOR U3105 ( .A(n3462), .B(n3463), .Z(n3459) );
  AND U3106 ( .A(n724), .B(n3464), .Z(n3463) );
  XOR U3107 ( .A(n3465), .B(n3466), .Z(n3457) );
  AND U3108 ( .A(n728), .B(n3467), .Z(n3466) );
  XOR U3109 ( .A(n3468), .B(n3469), .Z(n3454) );
  AND U3110 ( .A(n732), .B(n3467), .Z(n3469) );
  XNOR U3111 ( .A(n3470), .B(n3468), .Z(n3467) );
  IV U3112 ( .A(n3465), .Z(n3470) );
  XOR U3113 ( .A(n3471), .B(n3472), .Z(n3465) );
  AND U3114 ( .A(n735), .B(n3464), .Z(n3472) );
  XNOR U3115 ( .A(n3462), .B(n3471), .Z(n3464) );
  XNOR U3116 ( .A(n3473), .B(n3474), .Z(n3462) );
  AND U3117 ( .A(n739), .B(n3475), .Z(n3474) );
  XOR U3118 ( .A(p_input[1030]), .B(n3473), .Z(n3475) );
  XNOR U3119 ( .A(n3476), .B(n3477), .Z(n3473) );
  AND U3120 ( .A(n743), .B(n3478), .Z(n3477) );
  XOR U3121 ( .A(n3479), .B(n3480), .Z(n3471) );
  AND U3122 ( .A(n747), .B(n3481), .Z(n3480) );
  XOR U3123 ( .A(n3482), .B(n3483), .Z(n3468) );
  AND U3124 ( .A(n751), .B(n3481), .Z(n3483) );
  XNOR U3125 ( .A(n3484), .B(n3482), .Z(n3481) );
  IV U3126 ( .A(n3479), .Z(n3484) );
  XOR U3127 ( .A(n3485), .B(n3486), .Z(n3479) );
  AND U3128 ( .A(n754), .B(n3478), .Z(n3486) );
  XNOR U3129 ( .A(n3476), .B(n3485), .Z(n3478) );
  XNOR U3130 ( .A(n3487), .B(n3488), .Z(n3476) );
  AND U3131 ( .A(n758), .B(n3489), .Z(n3488) );
  XOR U3132 ( .A(p_input[1062]), .B(n3487), .Z(n3489) );
  XNOR U3133 ( .A(n3490), .B(n3491), .Z(n3487) );
  AND U3134 ( .A(n762), .B(n3492), .Z(n3491) );
  XOR U3135 ( .A(n3493), .B(n3494), .Z(n3485) );
  AND U3136 ( .A(n766), .B(n3495), .Z(n3494) );
  XOR U3137 ( .A(n3496), .B(n3497), .Z(n3482) );
  AND U3138 ( .A(n770), .B(n3495), .Z(n3497) );
  XNOR U3139 ( .A(n3498), .B(n3496), .Z(n3495) );
  IV U3140 ( .A(n3493), .Z(n3498) );
  XOR U3141 ( .A(n3499), .B(n3500), .Z(n3493) );
  AND U3142 ( .A(n773), .B(n3492), .Z(n3500) );
  XNOR U3143 ( .A(n3490), .B(n3499), .Z(n3492) );
  XNOR U3144 ( .A(n3501), .B(n3502), .Z(n3490) );
  AND U3145 ( .A(n777), .B(n3503), .Z(n3502) );
  XOR U3146 ( .A(p_input[1094]), .B(n3501), .Z(n3503) );
  XNOR U3147 ( .A(n3504), .B(n3505), .Z(n3501) );
  AND U3148 ( .A(n781), .B(n3506), .Z(n3505) );
  XOR U3149 ( .A(n3507), .B(n3508), .Z(n3499) );
  AND U3150 ( .A(n785), .B(n3509), .Z(n3508) );
  XOR U3151 ( .A(n3510), .B(n3511), .Z(n3496) );
  AND U3152 ( .A(n789), .B(n3509), .Z(n3511) );
  XNOR U3153 ( .A(n3512), .B(n3510), .Z(n3509) );
  IV U3154 ( .A(n3507), .Z(n3512) );
  XOR U3155 ( .A(n3513), .B(n3514), .Z(n3507) );
  AND U3156 ( .A(n792), .B(n3506), .Z(n3514) );
  XNOR U3157 ( .A(n3504), .B(n3513), .Z(n3506) );
  XNOR U3158 ( .A(n3515), .B(n3516), .Z(n3504) );
  AND U3159 ( .A(n796), .B(n3517), .Z(n3516) );
  XOR U3160 ( .A(p_input[1126]), .B(n3515), .Z(n3517) );
  XNOR U3161 ( .A(n3518), .B(n3519), .Z(n3515) );
  AND U3162 ( .A(n800), .B(n3520), .Z(n3519) );
  XOR U3163 ( .A(n3521), .B(n3522), .Z(n3513) );
  AND U3164 ( .A(n804), .B(n3523), .Z(n3522) );
  XOR U3165 ( .A(n3524), .B(n3525), .Z(n3510) );
  AND U3166 ( .A(n808), .B(n3523), .Z(n3525) );
  XNOR U3167 ( .A(n3526), .B(n3524), .Z(n3523) );
  IV U3168 ( .A(n3521), .Z(n3526) );
  XOR U3169 ( .A(n3527), .B(n3528), .Z(n3521) );
  AND U3170 ( .A(n811), .B(n3520), .Z(n3528) );
  XNOR U3171 ( .A(n3518), .B(n3527), .Z(n3520) );
  XNOR U3172 ( .A(n3529), .B(n3530), .Z(n3518) );
  AND U3173 ( .A(n815), .B(n3531), .Z(n3530) );
  XOR U3174 ( .A(p_input[1158]), .B(n3529), .Z(n3531) );
  XNOR U3175 ( .A(n3532), .B(n3533), .Z(n3529) );
  AND U3176 ( .A(n819), .B(n3534), .Z(n3533) );
  XOR U3177 ( .A(n3535), .B(n3536), .Z(n3527) );
  AND U3178 ( .A(n823), .B(n3537), .Z(n3536) );
  XOR U3179 ( .A(n3538), .B(n3539), .Z(n3524) );
  AND U3180 ( .A(n827), .B(n3537), .Z(n3539) );
  XNOR U3181 ( .A(n3540), .B(n3538), .Z(n3537) );
  IV U3182 ( .A(n3535), .Z(n3540) );
  XOR U3183 ( .A(n3541), .B(n3542), .Z(n3535) );
  AND U3184 ( .A(n830), .B(n3534), .Z(n3542) );
  XNOR U3185 ( .A(n3532), .B(n3541), .Z(n3534) );
  XNOR U3186 ( .A(n3543), .B(n3544), .Z(n3532) );
  AND U3187 ( .A(n834), .B(n3545), .Z(n3544) );
  XOR U3188 ( .A(p_input[1190]), .B(n3543), .Z(n3545) );
  XNOR U3189 ( .A(n3546), .B(n3547), .Z(n3543) );
  AND U3190 ( .A(n838), .B(n3548), .Z(n3547) );
  XOR U3191 ( .A(n3549), .B(n3550), .Z(n3541) );
  AND U3192 ( .A(n842), .B(n3551), .Z(n3550) );
  XOR U3193 ( .A(n3552), .B(n3553), .Z(n3538) );
  AND U3194 ( .A(n846), .B(n3551), .Z(n3553) );
  XNOR U3195 ( .A(n3554), .B(n3552), .Z(n3551) );
  IV U3196 ( .A(n3549), .Z(n3554) );
  XOR U3197 ( .A(n3555), .B(n3556), .Z(n3549) );
  AND U3198 ( .A(n849), .B(n3548), .Z(n3556) );
  XNOR U3199 ( .A(n3546), .B(n3555), .Z(n3548) );
  XNOR U3200 ( .A(n3557), .B(n3558), .Z(n3546) );
  AND U3201 ( .A(n853), .B(n3559), .Z(n3558) );
  XOR U3202 ( .A(p_input[1222]), .B(n3557), .Z(n3559) );
  XNOR U3203 ( .A(n3560), .B(n3561), .Z(n3557) );
  AND U3204 ( .A(n857), .B(n3562), .Z(n3561) );
  XOR U3205 ( .A(n3563), .B(n3564), .Z(n3555) );
  AND U3206 ( .A(n861), .B(n3565), .Z(n3564) );
  XOR U3207 ( .A(n3566), .B(n3567), .Z(n3552) );
  AND U3208 ( .A(n865), .B(n3565), .Z(n3567) );
  XNOR U3209 ( .A(n3568), .B(n3566), .Z(n3565) );
  IV U3210 ( .A(n3563), .Z(n3568) );
  XOR U3211 ( .A(n3569), .B(n3570), .Z(n3563) );
  AND U3212 ( .A(n868), .B(n3562), .Z(n3570) );
  XNOR U3213 ( .A(n3560), .B(n3569), .Z(n3562) );
  XNOR U3214 ( .A(n3571), .B(n3572), .Z(n3560) );
  AND U3215 ( .A(n872), .B(n3573), .Z(n3572) );
  XOR U3216 ( .A(p_input[1254]), .B(n3571), .Z(n3573) );
  XNOR U3217 ( .A(n3574), .B(n3575), .Z(n3571) );
  AND U3218 ( .A(n876), .B(n3576), .Z(n3575) );
  XOR U3219 ( .A(n3577), .B(n3578), .Z(n3569) );
  AND U3220 ( .A(n880), .B(n3579), .Z(n3578) );
  XOR U3221 ( .A(n3580), .B(n3581), .Z(n3566) );
  AND U3222 ( .A(n884), .B(n3579), .Z(n3581) );
  XNOR U3223 ( .A(n3582), .B(n3580), .Z(n3579) );
  IV U3224 ( .A(n3577), .Z(n3582) );
  XOR U3225 ( .A(n3583), .B(n3584), .Z(n3577) );
  AND U3226 ( .A(n887), .B(n3576), .Z(n3584) );
  XNOR U3227 ( .A(n3574), .B(n3583), .Z(n3576) );
  XNOR U3228 ( .A(n3585), .B(n3586), .Z(n3574) );
  AND U3229 ( .A(n891), .B(n3587), .Z(n3586) );
  XOR U3230 ( .A(p_input[1286]), .B(n3585), .Z(n3587) );
  XNOR U3231 ( .A(n3588), .B(n3589), .Z(n3585) );
  AND U3232 ( .A(n895), .B(n3590), .Z(n3589) );
  XOR U3233 ( .A(n3591), .B(n3592), .Z(n3583) );
  AND U3234 ( .A(n899), .B(n3593), .Z(n3592) );
  XOR U3235 ( .A(n3594), .B(n3595), .Z(n3580) );
  AND U3236 ( .A(n903), .B(n3593), .Z(n3595) );
  XNOR U3237 ( .A(n3596), .B(n3594), .Z(n3593) );
  IV U3238 ( .A(n3591), .Z(n3596) );
  XOR U3239 ( .A(n3597), .B(n3598), .Z(n3591) );
  AND U3240 ( .A(n906), .B(n3590), .Z(n3598) );
  XNOR U3241 ( .A(n3588), .B(n3597), .Z(n3590) );
  XNOR U3242 ( .A(n3599), .B(n3600), .Z(n3588) );
  AND U3243 ( .A(n910), .B(n3601), .Z(n3600) );
  XOR U3244 ( .A(p_input[1318]), .B(n3599), .Z(n3601) );
  XNOR U3245 ( .A(n3602), .B(n3603), .Z(n3599) );
  AND U3246 ( .A(n914), .B(n3604), .Z(n3603) );
  XOR U3247 ( .A(n3605), .B(n3606), .Z(n3597) );
  AND U3248 ( .A(n918), .B(n3607), .Z(n3606) );
  XOR U3249 ( .A(n3608), .B(n3609), .Z(n3594) );
  AND U3250 ( .A(n922), .B(n3607), .Z(n3609) );
  XNOR U3251 ( .A(n3610), .B(n3608), .Z(n3607) );
  IV U3252 ( .A(n3605), .Z(n3610) );
  XOR U3253 ( .A(n3611), .B(n3612), .Z(n3605) );
  AND U3254 ( .A(n925), .B(n3604), .Z(n3612) );
  XNOR U3255 ( .A(n3602), .B(n3611), .Z(n3604) );
  XNOR U3256 ( .A(n3613), .B(n3614), .Z(n3602) );
  AND U3257 ( .A(n929), .B(n3615), .Z(n3614) );
  XOR U3258 ( .A(p_input[1350]), .B(n3613), .Z(n3615) );
  XNOR U3259 ( .A(n3616), .B(n3617), .Z(n3613) );
  AND U3260 ( .A(n933), .B(n3618), .Z(n3617) );
  XOR U3261 ( .A(n3619), .B(n3620), .Z(n3611) );
  AND U3262 ( .A(n937), .B(n3621), .Z(n3620) );
  XOR U3263 ( .A(n3622), .B(n3623), .Z(n3608) );
  AND U3264 ( .A(n941), .B(n3621), .Z(n3623) );
  XNOR U3265 ( .A(n3624), .B(n3622), .Z(n3621) );
  IV U3266 ( .A(n3619), .Z(n3624) );
  XOR U3267 ( .A(n3625), .B(n3626), .Z(n3619) );
  AND U3268 ( .A(n944), .B(n3618), .Z(n3626) );
  XNOR U3269 ( .A(n3616), .B(n3625), .Z(n3618) );
  XNOR U3270 ( .A(n3627), .B(n3628), .Z(n3616) );
  AND U3271 ( .A(n948), .B(n3629), .Z(n3628) );
  XOR U3272 ( .A(p_input[1382]), .B(n3627), .Z(n3629) );
  XNOR U3273 ( .A(n3630), .B(n3631), .Z(n3627) );
  AND U3274 ( .A(n952), .B(n3632), .Z(n3631) );
  XOR U3275 ( .A(n3633), .B(n3634), .Z(n3625) );
  AND U3276 ( .A(n956), .B(n3635), .Z(n3634) );
  XOR U3277 ( .A(n3636), .B(n3637), .Z(n3622) );
  AND U3278 ( .A(n960), .B(n3635), .Z(n3637) );
  XNOR U3279 ( .A(n3638), .B(n3636), .Z(n3635) );
  IV U3280 ( .A(n3633), .Z(n3638) );
  XOR U3281 ( .A(n3639), .B(n3640), .Z(n3633) );
  AND U3282 ( .A(n963), .B(n3632), .Z(n3640) );
  XNOR U3283 ( .A(n3630), .B(n3639), .Z(n3632) );
  XNOR U3284 ( .A(n3641), .B(n3642), .Z(n3630) );
  AND U3285 ( .A(n967), .B(n3643), .Z(n3642) );
  XOR U3286 ( .A(p_input[1414]), .B(n3641), .Z(n3643) );
  XNOR U3287 ( .A(n3644), .B(n3645), .Z(n3641) );
  AND U3288 ( .A(n971), .B(n3646), .Z(n3645) );
  XOR U3289 ( .A(n3647), .B(n3648), .Z(n3639) );
  AND U3290 ( .A(n975), .B(n3649), .Z(n3648) );
  XOR U3291 ( .A(n3650), .B(n3651), .Z(n3636) );
  AND U3292 ( .A(n979), .B(n3649), .Z(n3651) );
  XNOR U3293 ( .A(n3652), .B(n3650), .Z(n3649) );
  IV U3294 ( .A(n3647), .Z(n3652) );
  XOR U3295 ( .A(n3653), .B(n3654), .Z(n3647) );
  AND U3296 ( .A(n982), .B(n3646), .Z(n3654) );
  XNOR U3297 ( .A(n3644), .B(n3653), .Z(n3646) );
  XNOR U3298 ( .A(n3655), .B(n3656), .Z(n3644) );
  AND U3299 ( .A(n986), .B(n3657), .Z(n3656) );
  XOR U3300 ( .A(p_input[1446]), .B(n3655), .Z(n3657) );
  XNOR U3301 ( .A(n3658), .B(n3659), .Z(n3655) );
  AND U3302 ( .A(n990), .B(n3660), .Z(n3659) );
  XOR U3303 ( .A(n3661), .B(n3662), .Z(n3653) );
  AND U3304 ( .A(n994), .B(n3663), .Z(n3662) );
  XOR U3305 ( .A(n3664), .B(n3665), .Z(n3650) );
  AND U3306 ( .A(n998), .B(n3663), .Z(n3665) );
  XNOR U3307 ( .A(n3666), .B(n3664), .Z(n3663) );
  IV U3308 ( .A(n3661), .Z(n3666) );
  XOR U3309 ( .A(n3667), .B(n3668), .Z(n3661) );
  AND U3310 ( .A(n1001), .B(n3660), .Z(n3668) );
  XNOR U3311 ( .A(n3658), .B(n3667), .Z(n3660) );
  XNOR U3312 ( .A(n3669), .B(n3670), .Z(n3658) );
  AND U3313 ( .A(n1005), .B(n3671), .Z(n3670) );
  XOR U3314 ( .A(p_input[1478]), .B(n3669), .Z(n3671) );
  XNOR U3315 ( .A(n3672), .B(n3673), .Z(n3669) );
  AND U3316 ( .A(n1009), .B(n3674), .Z(n3673) );
  XOR U3317 ( .A(n3675), .B(n3676), .Z(n3667) );
  AND U3318 ( .A(n1013), .B(n3677), .Z(n3676) );
  XOR U3319 ( .A(n3678), .B(n3679), .Z(n3664) );
  AND U3320 ( .A(n1017), .B(n3677), .Z(n3679) );
  XNOR U3321 ( .A(n3680), .B(n3678), .Z(n3677) );
  IV U3322 ( .A(n3675), .Z(n3680) );
  XOR U3323 ( .A(n3681), .B(n3682), .Z(n3675) );
  AND U3324 ( .A(n1020), .B(n3674), .Z(n3682) );
  XNOR U3325 ( .A(n3672), .B(n3681), .Z(n3674) );
  XNOR U3326 ( .A(n3683), .B(n3684), .Z(n3672) );
  AND U3327 ( .A(n1024), .B(n3685), .Z(n3684) );
  XOR U3328 ( .A(p_input[1510]), .B(n3683), .Z(n3685) );
  XNOR U3329 ( .A(n3686), .B(n3687), .Z(n3683) );
  AND U3330 ( .A(n1028), .B(n3688), .Z(n3687) );
  XOR U3331 ( .A(n3689), .B(n3690), .Z(n3681) );
  AND U3332 ( .A(n1032), .B(n3691), .Z(n3690) );
  XOR U3333 ( .A(n3692), .B(n3693), .Z(n3678) );
  AND U3334 ( .A(n1036), .B(n3691), .Z(n3693) );
  XNOR U3335 ( .A(n3694), .B(n3692), .Z(n3691) );
  IV U3336 ( .A(n3689), .Z(n3694) );
  XOR U3337 ( .A(n3695), .B(n3696), .Z(n3689) );
  AND U3338 ( .A(n1039), .B(n3688), .Z(n3696) );
  XNOR U3339 ( .A(n3686), .B(n3695), .Z(n3688) );
  XNOR U3340 ( .A(n3697), .B(n3698), .Z(n3686) );
  AND U3341 ( .A(n1043), .B(n3699), .Z(n3698) );
  XOR U3342 ( .A(p_input[1542]), .B(n3697), .Z(n3699) );
  XNOR U3343 ( .A(n3700), .B(n3701), .Z(n3697) );
  AND U3344 ( .A(n1047), .B(n3702), .Z(n3701) );
  XOR U3345 ( .A(n3703), .B(n3704), .Z(n3695) );
  AND U3346 ( .A(n1051), .B(n3705), .Z(n3704) );
  XOR U3347 ( .A(n3706), .B(n3707), .Z(n3692) );
  AND U3348 ( .A(n1055), .B(n3705), .Z(n3707) );
  XNOR U3349 ( .A(n3708), .B(n3706), .Z(n3705) );
  IV U3350 ( .A(n3703), .Z(n3708) );
  XOR U3351 ( .A(n3709), .B(n3710), .Z(n3703) );
  AND U3352 ( .A(n1058), .B(n3702), .Z(n3710) );
  XNOR U3353 ( .A(n3700), .B(n3709), .Z(n3702) );
  XNOR U3354 ( .A(n3711), .B(n3712), .Z(n3700) );
  AND U3355 ( .A(n1062), .B(n3713), .Z(n3712) );
  XOR U3356 ( .A(p_input[1574]), .B(n3711), .Z(n3713) );
  XNOR U3357 ( .A(n3714), .B(n3715), .Z(n3711) );
  AND U3358 ( .A(n1066), .B(n3716), .Z(n3715) );
  XOR U3359 ( .A(n3717), .B(n3718), .Z(n3709) );
  AND U3360 ( .A(n1070), .B(n3719), .Z(n3718) );
  XOR U3361 ( .A(n3720), .B(n3721), .Z(n3706) );
  AND U3362 ( .A(n1074), .B(n3719), .Z(n3721) );
  XNOR U3363 ( .A(n3722), .B(n3720), .Z(n3719) );
  IV U3364 ( .A(n3717), .Z(n3722) );
  XOR U3365 ( .A(n3723), .B(n3724), .Z(n3717) );
  AND U3366 ( .A(n1077), .B(n3716), .Z(n3724) );
  XNOR U3367 ( .A(n3714), .B(n3723), .Z(n3716) );
  XNOR U3368 ( .A(n3725), .B(n3726), .Z(n3714) );
  AND U3369 ( .A(n1081), .B(n3727), .Z(n3726) );
  XOR U3370 ( .A(p_input[1606]), .B(n3725), .Z(n3727) );
  XNOR U3371 ( .A(n3728), .B(n3729), .Z(n3725) );
  AND U3372 ( .A(n1085), .B(n3730), .Z(n3729) );
  XOR U3373 ( .A(n3731), .B(n3732), .Z(n3723) );
  AND U3374 ( .A(n1089), .B(n3733), .Z(n3732) );
  XOR U3375 ( .A(n3734), .B(n3735), .Z(n3720) );
  AND U3376 ( .A(n1093), .B(n3733), .Z(n3735) );
  XNOR U3377 ( .A(n3736), .B(n3734), .Z(n3733) );
  IV U3378 ( .A(n3731), .Z(n3736) );
  XOR U3379 ( .A(n3737), .B(n3738), .Z(n3731) );
  AND U3380 ( .A(n1096), .B(n3730), .Z(n3738) );
  XNOR U3381 ( .A(n3728), .B(n3737), .Z(n3730) );
  XNOR U3382 ( .A(n3739), .B(n3740), .Z(n3728) );
  AND U3383 ( .A(n1100), .B(n3741), .Z(n3740) );
  XOR U3384 ( .A(p_input[1638]), .B(n3739), .Z(n3741) );
  XNOR U3385 ( .A(n3742), .B(n3743), .Z(n3739) );
  AND U3386 ( .A(n1104), .B(n3744), .Z(n3743) );
  XOR U3387 ( .A(n3745), .B(n3746), .Z(n3737) );
  AND U3388 ( .A(n1108), .B(n3747), .Z(n3746) );
  XOR U3389 ( .A(n3748), .B(n3749), .Z(n3734) );
  AND U3390 ( .A(n1112), .B(n3747), .Z(n3749) );
  XNOR U3391 ( .A(n3750), .B(n3748), .Z(n3747) );
  IV U3392 ( .A(n3745), .Z(n3750) );
  XOR U3393 ( .A(n3751), .B(n3752), .Z(n3745) );
  AND U3394 ( .A(n1115), .B(n3744), .Z(n3752) );
  XNOR U3395 ( .A(n3742), .B(n3751), .Z(n3744) );
  XNOR U3396 ( .A(n3753), .B(n3754), .Z(n3742) );
  AND U3397 ( .A(n1119), .B(n3755), .Z(n3754) );
  XOR U3398 ( .A(p_input[1670]), .B(n3753), .Z(n3755) );
  XNOR U3399 ( .A(n3756), .B(n3757), .Z(n3753) );
  AND U3400 ( .A(n1123), .B(n3758), .Z(n3757) );
  XOR U3401 ( .A(n3759), .B(n3760), .Z(n3751) );
  AND U3402 ( .A(n1127), .B(n3761), .Z(n3760) );
  XOR U3403 ( .A(n3762), .B(n3763), .Z(n3748) );
  AND U3404 ( .A(n1131), .B(n3761), .Z(n3763) );
  XNOR U3405 ( .A(n3764), .B(n3762), .Z(n3761) );
  IV U3406 ( .A(n3759), .Z(n3764) );
  XOR U3407 ( .A(n3765), .B(n3766), .Z(n3759) );
  AND U3408 ( .A(n1134), .B(n3758), .Z(n3766) );
  XNOR U3409 ( .A(n3756), .B(n3765), .Z(n3758) );
  XNOR U3410 ( .A(n3767), .B(n3768), .Z(n3756) );
  AND U3411 ( .A(n1138), .B(n3769), .Z(n3768) );
  XOR U3412 ( .A(p_input[1702]), .B(n3767), .Z(n3769) );
  XNOR U3413 ( .A(n3770), .B(n3771), .Z(n3767) );
  AND U3414 ( .A(n1142), .B(n3772), .Z(n3771) );
  XOR U3415 ( .A(n3773), .B(n3774), .Z(n3765) );
  AND U3416 ( .A(n1146), .B(n3775), .Z(n3774) );
  XOR U3417 ( .A(n3776), .B(n3777), .Z(n3762) );
  AND U3418 ( .A(n1150), .B(n3775), .Z(n3777) );
  XNOR U3419 ( .A(n3778), .B(n3776), .Z(n3775) );
  IV U3420 ( .A(n3773), .Z(n3778) );
  XOR U3421 ( .A(n3779), .B(n3780), .Z(n3773) );
  AND U3422 ( .A(n1153), .B(n3772), .Z(n3780) );
  XNOR U3423 ( .A(n3770), .B(n3779), .Z(n3772) );
  XNOR U3424 ( .A(n3781), .B(n3782), .Z(n3770) );
  AND U3425 ( .A(n1157), .B(n3783), .Z(n3782) );
  XOR U3426 ( .A(p_input[1734]), .B(n3781), .Z(n3783) );
  XNOR U3427 ( .A(n3784), .B(n3785), .Z(n3781) );
  AND U3428 ( .A(n1161), .B(n3786), .Z(n3785) );
  XOR U3429 ( .A(n3787), .B(n3788), .Z(n3779) );
  AND U3430 ( .A(n1165), .B(n3789), .Z(n3788) );
  XOR U3431 ( .A(n3790), .B(n3791), .Z(n3776) );
  AND U3432 ( .A(n1169), .B(n3789), .Z(n3791) );
  XNOR U3433 ( .A(n3792), .B(n3790), .Z(n3789) );
  IV U3434 ( .A(n3787), .Z(n3792) );
  XOR U3435 ( .A(n3793), .B(n3794), .Z(n3787) );
  AND U3436 ( .A(n1172), .B(n3786), .Z(n3794) );
  XNOR U3437 ( .A(n3784), .B(n3793), .Z(n3786) );
  XNOR U3438 ( .A(n3795), .B(n3796), .Z(n3784) );
  AND U3439 ( .A(n1176), .B(n3797), .Z(n3796) );
  XOR U3440 ( .A(p_input[1766]), .B(n3795), .Z(n3797) );
  XNOR U3441 ( .A(n3798), .B(n3799), .Z(n3795) );
  AND U3442 ( .A(n1180), .B(n3800), .Z(n3799) );
  XOR U3443 ( .A(n3801), .B(n3802), .Z(n3793) );
  AND U3444 ( .A(n1184), .B(n3803), .Z(n3802) );
  XOR U3445 ( .A(n3804), .B(n3805), .Z(n3790) );
  AND U3446 ( .A(n1188), .B(n3803), .Z(n3805) );
  XNOR U3447 ( .A(n3806), .B(n3804), .Z(n3803) );
  IV U3448 ( .A(n3801), .Z(n3806) );
  XOR U3449 ( .A(n3807), .B(n3808), .Z(n3801) );
  AND U3450 ( .A(n1191), .B(n3800), .Z(n3808) );
  XNOR U3451 ( .A(n3798), .B(n3807), .Z(n3800) );
  XNOR U3452 ( .A(n3809), .B(n3810), .Z(n3798) );
  AND U3453 ( .A(n1195), .B(n3811), .Z(n3810) );
  XOR U3454 ( .A(p_input[1798]), .B(n3809), .Z(n3811) );
  XNOR U3455 ( .A(n3812), .B(n3813), .Z(n3809) );
  AND U3456 ( .A(n1199), .B(n3814), .Z(n3813) );
  XOR U3457 ( .A(n3815), .B(n3816), .Z(n3807) );
  AND U3458 ( .A(n1203), .B(n3817), .Z(n3816) );
  XOR U3459 ( .A(n3818), .B(n3819), .Z(n3804) );
  AND U3460 ( .A(n1207), .B(n3817), .Z(n3819) );
  XNOR U3461 ( .A(n3820), .B(n3818), .Z(n3817) );
  IV U3462 ( .A(n3815), .Z(n3820) );
  XOR U3463 ( .A(n3821), .B(n3822), .Z(n3815) );
  AND U3464 ( .A(n1210), .B(n3814), .Z(n3822) );
  XNOR U3465 ( .A(n3812), .B(n3821), .Z(n3814) );
  XNOR U3466 ( .A(n3823), .B(n3824), .Z(n3812) );
  AND U3467 ( .A(n1214), .B(n3825), .Z(n3824) );
  XOR U3468 ( .A(p_input[1830]), .B(n3823), .Z(n3825) );
  XNOR U3469 ( .A(n3826), .B(n3827), .Z(n3823) );
  AND U3470 ( .A(n1218), .B(n3828), .Z(n3827) );
  XOR U3471 ( .A(n3829), .B(n3830), .Z(n3821) );
  AND U3472 ( .A(n1222), .B(n3831), .Z(n3830) );
  XOR U3473 ( .A(n3832), .B(n3833), .Z(n3818) );
  AND U3474 ( .A(n1226), .B(n3831), .Z(n3833) );
  XNOR U3475 ( .A(n3834), .B(n3832), .Z(n3831) );
  IV U3476 ( .A(n3829), .Z(n3834) );
  XOR U3477 ( .A(n3835), .B(n3836), .Z(n3829) );
  AND U3478 ( .A(n1229), .B(n3828), .Z(n3836) );
  XNOR U3479 ( .A(n3826), .B(n3835), .Z(n3828) );
  XNOR U3480 ( .A(n3837), .B(n3838), .Z(n3826) );
  AND U3481 ( .A(n1233), .B(n3839), .Z(n3838) );
  XOR U3482 ( .A(p_input[1862]), .B(n3837), .Z(n3839) );
  XNOR U3483 ( .A(n3840), .B(n3841), .Z(n3837) );
  AND U3484 ( .A(n1237), .B(n3842), .Z(n3841) );
  XOR U3485 ( .A(n3843), .B(n3844), .Z(n3835) );
  AND U3486 ( .A(n1241), .B(n3845), .Z(n3844) );
  XOR U3487 ( .A(n3846), .B(n3847), .Z(n3832) );
  AND U3488 ( .A(n1245), .B(n3845), .Z(n3847) );
  XNOR U3489 ( .A(n3848), .B(n3846), .Z(n3845) );
  IV U3490 ( .A(n3843), .Z(n3848) );
  XOR U3491 ( .A(n3849), .B(n3850), .Z(n3843) );
  AND U3492 ( .A(n1248), .B(n3842), .Z(n3850) );
  XNOR U3493 ( .A(n3840), .B(n3849), .Z(n3842) );
  XNOR U3494 ( .A(n3851), .B(n3852), .Z(n3840) );
  AND U3495 ( .A(n1252), .B(n3853), .Z(n3852) );
  XOR U3496 ( .A(p_input[1894]), .B(n3851), .Z(n3853) );
  XNOR U3497 ( .A(n3854), .B(n3855), .Z(n3851) );
  AND U3498 ( .A(n1256), .B(n3856), .Z(n3855) );
  XOR U3499 ( .A(n3857), .B(n3858), .Z(n3849) );
  AND U3500 ( .A(n1260), .B(n3859), .Z(n3858) );
  XOR U3501 ( .A(n3860), .B(n3861), .Z(n3846) );
  AND U3502 ( .A(n1264), .B(n3859), .Z(n3861) );
  XNOR U3503 ( .A(n3862), .B(n3860), .Z(n3859) );
  IV U3504 ( .A(n3857), .Z(n3862) );
  XOR U3505 ( .A(n3863), .B(n3864), .Z(n3857) );
  AND U3506 ( .A(n1267), .B(n3856), .Z(n3864) );
  XNOR U3507 ( .A(n3854), .B(n3863), .Z(n3856) );
  XNOR U3508 ( .A(n3865), .B(n3866), .Z(n3854) );
  AND U3509 ( .A(n1271), .B(n3867), .Z(n3866) );
  XOR U3510 ( .A(p_input[1926]), .B(n3865), .Z(n3867) );
  XOR U3511 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(n3868), 
        .Z(n3865) );
  AND U3512 ( .A(n1274), .B(n3869), .Z(n3868) );
  XOR U3513 ( .A(n3870), .B(n3871), .Z(n3863) );
  AND U3514 ( .A(n1278), .B(n3872), .Z(n3871) );
  XOR U3515 ( .A(n3873), .B(n3874), .Z(n3860) );
  AND U3516 ( .A(n1282), .B(n3872), .Z(n3874) );
  XNOR U3517 ( .A(n3875), .B(n3873), .Z(n3872) );
  IV U3518 ( .A(n3870), .Z(n3875) );
  XOR U3519 ( .A(n3876), .B(n3877), .Z(n3870) );
  AND U3520 ( .A(n1285), .B(n3869), .Z(n3877) );
  XOR U3521 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(n3876), 
        .Z(n3869) );
  XOR U3522 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .B(n3878), 
        .Z(n3876) );
  AND U3523 ( .A(n1287), .B(n3879), .Z(n3878) );
  XOR U3524 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n3880), .Z(n3873) );
  AND U3525 ( .A(n1290), .B(n3879), .Z(n3880) );
  XOR U3526 ( .A(\knn_comb_/min_val_out[0][6] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .Z(n3879) );
  XOR U3527 ( .A(n81), .B(n3881), .Z(o[37]) );
  AND U3528 ( .A(n122), .B(n3882), .Z(n81) );
  XOR U3529 ( .A(n82), .B(n3881), .Z(n3882) );
  XOR U3530 ( .A(n3883), .B(n61), .Z(n3881) );
  AND U3531 ( .A(n125), .B(n3884), .Z(n61) );
  XOR U3532 ( .A(n62), .B(n3883), .Z(n3884) );
  XOR U3533 ( .A(n3885), .B(n3886), .Z(n62) );
  AND U3534 ( .A(n130), .B(n3887), .Z(n3886) );
  XOR U3535 ( .A(p_input[5]), .B(n3885), .Z(n3887) );
  XNOR U3536 ( .A(n3888), .B(n3889), .Z(n3885) );
  AND U3537 ( .A(n134), .B(n3890), .Z(n3889) );
  XOR U3538 ( .A(n3891), .B(n3892), .Z(n3883) );
  AND U3539 ( .A(n138), .B(n3893), .Z(n3892) );
  XOR U3540 ( .A(n3894), .B(n3895), .Z(n82) );
  AND U3541 ( .A(n142), .B(n3893), .Z(n3895) );
  XNOR U3542 ( .A(n3896), .B(n3894), .Z(n3893) );
  IV U3543 ( .A(n3891), .Z(n3896) );
  XOR U3544 ( .A(n3897), .B(n3898), .Z(n3891) );
  AND U3545 ( .A(n146), .B(n3890), .Z(n3898) );
  XNOR U3546 ( .A(n3888), .B(n3897), .Z(n3890) );
  XNOR U3547 ( .A(n3899), .B(n3900), .Z(n3888) );
  AND U3548 ( .A(n150), .B(n3901), .Z(n3900) );
  XOR U3549 ( .A(p_input[37]), .B(n3899), .Z(n3901) );
  XNOR U3550 ( .A(n3902), .B(n3903), .Z(n3899) );
  AND U3551 ( .A(n154), .B(n3904), .Z(n3903) );
  XOR U3552 ( .A(n3905), .B(n3906), .Z(n3897) );
  AND U3553 ( .A(n158), .B(n3907), .Z(n3906) );
  XOR U3554 ( .A(n3908), .B(n3909), .Z(n3894) );
  AND U3555 ( .A(n162), .B(n3907), .Z(n3909) );
  XNOR U3556 ( .A(n3910), .B(n3908), .Z(n3907) );
  IV U3557 ( .A(n3905), .Z(n3910) );
  XOR U3558 ( .A(n3911), .B(n3912), .Z(n3905) );
  AND U3559 ( .A(n165), .B(n3904), .Z(n3912) );
  XNOR U3560 ( .A(n3902), .B(n3911), .Z(n3904) );
  XNOR U3561 ( .A(n3913), .B(n3914), .Z(n3902) );
  AND U3562 ( .A(n169), .B(n3915), .Z(n3914) );
  XOR U3563 ( .A(p_input[69]), .B(n3913), .Z(n3915) );
  XNOR U3564 ( .A(n3916), .B(n3917), .Z(n3913) );
  AND U3565 ( .A(n173), .B(n3918), .Z(n3917) );
  XOR U3566 ( .A(n3919), .B(n3920), .Z(n3911) );
  AND U3567 ( .A(n177), .B(n3921), .Z(n3920) );
  XOR U3568 ( .A(n3922), .B(n3923), .Z(n3908) );
  AND U3569 ( .A(n181), .B(n3921), .Z(n3923) );
  XNOR U3570 ( .A(n3924), .B(n3922), .Z(n3921) );
  IV U3571 ( .A(n3919), .Z(n3924) );
  XOR U3572 ( .A(n3925), .B(n3926), .Z(n3919) );
  AND U3573 ( .A(n184), .B(n3918), .Z(n3926) );
  XNOR U3574 ( .A(n3916), .B(n3925), .Z(n3918) );
  XNOR U3575 ( .A(n3927), .B(n3928), .Z(n3916) );
  AND U3576 ( .A(n188), .B(n3929), .Z(n3928) );
  XOR U3577 ( .A(p_input[101]), .B(n3927), .Z(n3929) );
  XNOR U3578 ( .A(n3930), .B(n3931), .Z(n3927) );
  AND U3579 ( .A(n192), .B(n3932), .Z(n3931) );
  XOR U3580 ( .A(n3933), .B(n3934), .Z(n3925) );
  AND U3581 ( .A(n196), .B(n3935), .Z(n3934) );
  XOR U3582 ( .A(n3936), .B(n3937), .Z(n3922) );
  AND U3583 ( .A(n200), .B(n3935), .Z(n3937) );
  XNOR U3584 ( .A(n3938), .B(n3936), .Z(n3935) );
  IV U3585 ( .A(n3933), .Z(n3938) );
  XOR U3586 ( .A(n3939), .B(n3940), .Z(n3933) );
  AND U3587 ( .A(n203), .B(n3932), .Z(n3940) );
  XNOR U3588 ( .A(n3930), .B(n3939), .Z(n3932) );
  XNOR U3589 ( .A(n3941), .B(n3942), .Z(n3930) );
  AND U3590 ( .A(n207), .B(n3943), .Z(n3942) );
  XOR U3591 ( .A(p_input[133]), .B(n3941), .Z(n3943) );
  XNOR U3592 ( .A(n3944), .B(n3945), .Z(n3941) );
  AND U3593 ( .A(n211), .B(n3946), .Z(n3945) );
  XOR U3594 ( .A(n3947), .B(n3948), .Z(n3939) );
  AND U3595 ( .A(n215), .B(n3949), .Z(n3948) );
  XOR U3596 ( .A(n3950), .B(n3951), .Z(n3936) );
  AND U3597 ( .A(n219), .B(n3949), .Z(n3951) );
  XNOR U3598 ( .A(n3952), .B(n3950), .Z(n3949) );
  IV U3599 ( .A(n3947), .Z(n3952) );
  XOR U3600 ( .A(n3953), .B(n3954), .Z(n3947) );
  AND U3601 ( .A(n222), .B(n3946), .Z(n3954) );
  XNOR U3602 ( .A(n3944), .B(n3953), .Z(n3946) );
  XNOR U3603 ( .A(n3955), .B(n3956), .Z(n3944) );
  AND U3604 ( .A(n226), .B(n3957), .Z(n3956) );
  XOR U3605 ( .A(p_input[165]), .B(n3955), .Z(n3957) );
  XNOR U3606 ( .A(n3958), .B(n3959), .Z(n3955) );
  AND U3607 ( .A(n230), .B(n3960), .Z(n3959) );
  XOR U3608 ( .A(n3961), .B(n3962), .Z(n3953) );
  AND U3609 ( .A(n234), .B(n3963), .Z(n3962) );
  XOR U3610 ( .A(n3964), .B(n3965), .Z(n3950) );
  AND U3611 ( .A(n238), .B(n3963), .Z(n3965) );
  XNOR U3612 ( .A(n3966), .B(n3964), .Z(n3963) );
  IV U3613 ( .A(n3961), .Z(n3966) );
  XOR U3614 ( .A(n3967), .B(n3968), .Z(n3961) );
  AND U3615 ( .A(n241), .B(n3960), .Z(n3968) );
  XNOR U3616 ( .A(n3958), .B(n3967), .Z(n3960) );
  XNOR U3617 ( .A(n3969), .B(n3970), .Z(n3958) );
  AND U3618 ( .A(n245), .B(n3971), .Z(n3970) );
  XOR U3619 ( .A(p_input[197]), .B(n3969), .Z(n3971) );
  XNOR U3620 ( .A(n3972), .B(n3973), .Z(n3969) );
  AND U3621 ( .A(n249), .B(n3974), .Z(n3973) );
  XOR U3622 ( .A(n3975), .B(n3976), .Z(n3967) );
  AND U3623 ( .A(n253), .B(n3977), .Z(n3976) );
  XOR U3624 ( .A(n3978), .B(n3979), .Z(n3964) );
  AND U3625 ( .A(n257), .B(n3977), .Z(n3979) );
  XNOR U3626 ( .A(n3980), .B(n3978), .Z(n3977) );
  IV U3627 ( .A(n3975), .Z(n3980) );
  XOR U3628 ( .A(n3981), .B(n3982), .Z(n3975) );
  AND U3629 ( .A(n260), .B(n3974), .Z(n3982) );
  XNOR U3630 ( .A(n3972), .B(n3981), .Z(n3974) );
  XNOR U3631 ( .A(n3983), .B(n3984), .Z(n3972) );
  AND U3632 ( .A(n264), .B(n3985), .Z(n3984) );
  XOR U3633 ( .A(p_input[229]), .B(n3983), .Z(n3985) );
  XNOR U3634 ( .A(n3986), .B(n3987), .Z(n3983) );
  AND U3635 ( .A(n268), .B(n3988), .Z(n3987) );
  XOR U3636 ( .A(n3989), .B(n3990), .Z(n3981) );
  AND U3637 ( .A(n272), .B(n3991), .Z(n3990) );
  XOR U3638 ( .A(n3992), .B(n3993), .Z(n3978) );
  AND U3639 ( .A(n276), .B(n3991), .Z(n3993) );
  XNOR U3640 ( .A(n3994), .B(n3992), .Z(n3991) );
  IV U3641 ( .A(n3989), .Z(n3994) );
  XOR U3642 ( .A(n3995), .B(n3996), .Z(n3989) );
  AND U3643 ( .A(n279), .B(n3988), .Z(n3996) );
  XNOR U3644 ( .A(n3986), .B(n3995), .Z(n3988) );
  XNOR U3645 ( .A(n3997), .B(n3998), .Z(n3986) );
  AND U3646 ( .A(n283), .B(n3999), .Z(n3998) );
  XOR U3647 ( .A(p_input[261]), .B(n3997), .Z(n3999) );
  XNOR U3648 ( .A(n4000), .B(n4001), .Z(n3997) );
  AND U3649 ( .A(n287), .B(n4002), .Z(n4001) );
  XOR U3650 ( .A(n4003), .B(n4004), .Z(n3995) );
  AND U3651 ( .A(n291), .B(n4005), .Z(n4004) );
  XOR U3652 ( .A(n4006), .B(n4007), .Z(n3992) );
  AND U3653 ( .A(n295), .B(n4005), .Z(n4007) );
  XNOR U3654 ( .A(n4008), .B(n4006), .Z(n4005) );
  IV U3655 ( .A(n4003), .Z(n4008) );
  XOR U3656 ( .A(n4009), .B(n4010), .Z(n4003) );
  AND U3657 ( .A(n298), .B(n4002), .Z(n4010) );
  XNOR U3658 ( .A(n4000), .B(n4009), .Z(n4002) );
  XNOR U3659 ( .A(n4011), .B(n4012), .Z(n4000) );
  AND U3660 ( .A(n302), .B(n4013), .Z(n4012) );
  XOR U3661 ( .A(p_input[293]), .B(n4011), .Z(n4013) );
  XNOR U3662 ( .A(n4014), .B(n4015), .Z(n4011) );
  AND U3663 ( .A(n306), .B(n4016), .Z(n4015) );
  XOR U3664 ( .A(n4017), .B(n4018), .Z(n4009) );
  AND U3665 ( .A(n310), .B(n4019), .Z(n4018) );
  XOR U3666 ( .A(n4020), .B(n4021), .Z(n4006) );
  AND U3667 ( .A(n314), .B(n4019), .Z(n4021) );
  XNOR U3668 ( .A(n4022), .B(n4020), .Z(n4019) );
  IV U3669 ( .A(n4017), .Z(n4022) );
  XOR U3670 ( .A(n4023), .B(n4024), .Z(n4017) );
  AND U3671 ( .A(n317), .B(n4016), .Z(n4024) );
  XNOR U3672 ( .A(n4014), .B(n4023), .Z(n4016) );
  XNOR U3673 ( .A(n4025), .B(n4026), .Z(n4014) );
  AND U3674 ( .A(n321), .B(n4027), .Z(n4026) );
  XOR U3675 ( .A(p_input[325]), .B(n4025), .Z(n4027) );
  XNOR U3676 ( .A(n4028), .B(n4029), .Z(n4025) );
  AND U3677 ( .A(n325), .B(n4030), .Z(n4029) );
  XOR U3678 ( .A(n4031), .B(n4032), .Z(n4023) );
  AND U3679 ( .A(n329), .B(n4033), .Z(n4032) );
  XOR U3680 ( .A(n4034), .B(n4035), .Z(n4020) );
  AND U3681 ( .A(n333), .B(n4033), .Z(n4035) );
  XNOR U3682 ( .A(n4036), .B(n4034), .Z(n4033) );
  IV U3683 ( .A(n4031), .Z(n4036) );
  XOR U3684 ( .A(n4037), .B(n4038), .Z(n4031) );
  AND U3685 ( .A(n336), .B(n4030), .Z(n4038) );
  XNOR U3686 ( .A(n4028), .B(n4037), .Z(n4030) );
  XNOR U3687 ( .A(n4039), .B(n4040), .Z(n4028) );
  AND U3688 ( .A(n340), .B(n4041), .Z(n4040) );
  XOR U3689 ( .A(p_input[357]), .B(n4039), .Z(n4041) );
  XNOR U3690 ( .A(n4042), .B(n4043), .Z(n4039) );
  AND U3691 ( .A(n344), .B(n4044), .Z(n4043) );
  XOR U3692 ( .A(n4045), .B(n4046), .Z(n4037) );
  AND U3693 ( .A(n348), .B(n4047), .Z(n4046) );
  XOR U3694 ( .A(n4048), .B(n4049), .Z(n4034) );
  AND U3695 ( .A(n352), .B(n4047), .Z(n4049) );
  XNOR U3696 ( .A(n4050), .B(n4048), .Z(n4047) );
  IV U3697 ( .A(n4045), .Z(n4050) );
  XOR U3698 ( .A(n4051), .B(n4052), .Z(n4045) );
  AND U3699 ( .A(n355), .B(n4044), .Z(n4052) );
  XNOR U3700 ( .A(n4042), .B(n4051), .Z(n4044) );
  XNOR U3701 ( .A(n4053), .B(n4054), .Z(n4042) );
  AND U3702 ( .A(n359), .B(n4055), .Z(n4054) );
  XOR U3703 ( .A(p_input[389]), .B(n4053), .Z(n4055) );
  XNOR U3704 ( .A(n4056), .B(n4057), .Z(n4053) );
  AND U3705 ( .A(n363), .B(n4058), .Z(n4057) );
  XOR U3706 ( .A(n4059), .B(n4060), .Z(n4051) );
  AND U3707 ( .A(n367), .B(n4061), .Z(n4060) );
  XOR U3708 ( .A(n4062), .B(n4063), .Z(n4048) );
  AND U3709 ( .A(n371), .B(n4061), .Z(n4063) );
  XNOR U3710 ( .A(n4064), .B(n4062), .Z(n4061) );
  IV U3711 ( .A(n4059), .Z(n4064) );
  XOR U3712 ( .A(n4065), .B(n4066), .Z(n4059) );
  AND U3713 ( .A(n374), .B(n4058), .Z(n4066) );
  XNOR U3714 ( .A(n4056), .B(n4065), .Z(n4058) );
  XNOR U3715 ( .A(n4067), .B(n4068), .Z(n4056) );
  AND U3716 ( .A(n378), .B(n4069), .Z(n4068) );
  XOR U3717 ( .A(p_input[421]), .B(n4067), .Z(n4069) );
  XNOR U3718 ( .A(n4070), .B(n4071), .Z(n4067) );
  AND U3719 ( .A(n382), .B(n4072), .Z(n4071) );
  XOR U3720 ( .A(n4073), .B(n4074), .Z(n4065) );
  AND U3721 ( .A(n386), .B(n4075), .Z(n4074) );
  XOR U3722 ( .A(n4076), .B(n4077), .Z(n4062) );
  AND U3723 ( .A(n390), .B(n4075), .Z(n4077) );
  XNOR U3724 ( .A(n4078), .B(n4076), .Z(n4075) );
  IV U3725 ( .A(n4073), .Z(n4078) );
  XOR U3726 ( .A(n4079), .B(n4080), .Z(n4073) );
  AND U3727 ( .A(n393), .B(n4072), .Z(n4080) );
  XNOR U3728 ( .A(n4070), .B(n4079), .Z(n4072) );
  XNOR U3729 ( .A(n4081), .B(n4082), .Z(n4070) );
  AND U3730 ( .A(n397), .B(n4083), .Z(n4082) );
  XOR U3731 ( .A(p_input[453]), .B(n4081), .Z(n4083) );
  XNOR U3732 ( .A(n4084), .B(n4085), .Z(n4081) );
  AND U3733 ( .A(n401), .B(n4086), .Z(n4085) );
  XOR U3734 ( .A(n4087), .B(n4088), .Z(n4079) );
  AND U3735 ( .A(n405), .B(n4089), .Z(n4088) );
  XOR U3736 ( .A(n4090), .B(n4091), .Z(n4076) );
  AND U3737 ( .A(n409), .B(n4089), .Z(n4091) );
  XNOR U3738 ( .A(n4092), .B(n4090), .Z(n4089) );
  IV U3739 ( .A(n4087), .Z(n4092) );
  XOR U3740 ( .A(n4093), .B(n4094), .Z(n4087) );
  AND U3741 ( .A(n412), .B(n4086), .Z(n4094) );
  XNOR U3742 ( .A(n4084), .B(n4093), .Z(n4086) );
  XNOR U3743 ( .A(n4095), .B(n4096), .Z(n4084) );
  AND U3744 ( .A(n416), .B(n4097), .Z(n4096) );
  XOR U3745 ( .A(p_input[485]), .B(n4095), .Z(n4097) );
  XNOR U3746 ( .A(n4098), .B(n4099), .Z(n4095) );
  AND U3747 ( .A(n420), .B(n4100), .Z(n4099) );
  XOR U3748 ( .A(n4101), .B(n4102), .Z(n4093) );
  AND U3749 ( .A(n424), .B(n4103), .Z(n4102) );
  XOR U3750 ( .A(n4104), .B(n4105), .Z(n4090) );
  AND U3751 ( .A(n428), .B(n4103), .Z(n4105) );
  XNOR U3752 ( .A(n4106), .B(n4104), .Z(n4103) );
  IV U3753 ( .A(n4101), .Z(n4106) );
  XOR U3754 ( .A(n4107), .B(n4108), .Z(n4101) );
  AND U3755 ( .A(n431), .B(n4100), .Z(n4108) );
  XNOR U3756 ( .A(n4098), .B(n4107), .Z(n4100) );
  XNOR U3757 ( .A(n4109), .B(n4110), .Z(n4098) );
  AND U3758 ( .A(n435), .B(n4111), .Z(n4110) );
  XOR U3759 ( .A(p_input[517]), .B(n4109), .Z(n4111) );
  XNOR U3760 ( .A(n4112), .B(n4113), .Z(n4109) );
  AND U3761 ( .A(n439), .B(n4114), .Z(n4113) );
  XOR U3762 ( .A(n4115), .B(n4116), .Z(n4107) );
  AND U3763 ( .A(n443), .B(n4117), .Z(n4116) );
  XOR U3764 ( .A(n4118), .B(n4119), .Z(n4104) );
  AND U3765 ( .A(n447), .B(n4117), .Z(n4119) );
  XNOR U3766 ( .A(n4120), .B(n4118), .Z(n4117) );
  IV U3767 ( .A(n4115), .Z(n4120) );
  XOR U3768 ( .A(n4121), .B(n4122), .Z(n4115) );
  AND U3769 ( .A(n450), .B(n4114), .Z(n4122) );
  XNOR U3770 ( .A(n4112), .B(n4121), .Z(n4114) );
  XNOR U3771 ( .A(n4123), .B(n4124), .Z(n4112) );
  AND U3772 ( .A(n454), .B(n4125), .Z(n4124) );
  XOR U3773 ( .A(p_input[549]), .B(n4123), .Z(n4125) );
  XNOR U3774 ( .A(n4126), .B(n4127), .Z(n4123) );
  AND U3775 ( .A(n458), .B(n4128), .Z(n4127) );
  XOR U3776 ( .A(n4129), .B(n4130), .Z(n4121) );
  AND U3777 ( .A(n462), .B(n4131), .Z(n4130) );
  XOR U3778 ( .A(n4132), .B(n4133), .Z(n4118) );
  AND U3779 ( .A(n466), .B(n4131), .Z(n4133) );
  XNOR U3780 ( .A(n4134), .B(n4132), .Z(n4131) );
  IV U3781 ( .A(n4129), .Z(n4134) );
  XOR U3782 ( .A(n4135), .B(n4136), .Z(n4129) );
  AND U3783 ( .A(n469), .B(n4128), .Z(n4136) );
  XNOR U3784 ( .A(n4126), .B(n4135), .Z(n4128) );
  XNOR U3785 ( .A(n4137), .B(n4138), .Z(n4126) );
  AND U3786 ( .A(n473), .B(n4139), .Z(n4138) );
  XOR U3787 ( .A(p_input[581]), .B(n4137), .Z(n4139) );
  XNOR U3788 ( .A(n4140), .B(n4141), .Z(n4137) );
  AND U3789 ( .A(n477), .B(n4142), .Z(n4141) );
  XOR U3790 ( .A(n4143), .B(n4144), .Z(n4135) );
  AND U3791 ( .A(n481), .B(n4145), .Z(n4144) );
  XOR U3792 ( .A(n4146), .B(n4147), .Z(n4132) );
  AND U3793 ( .A(n485), .B(n4145), .Z(n4147) );
  XNOR U3794 ( .A(n4148), .B(n4146), .Z(n4145) );
  IV U3795 ( .A(n4143), .Z(n4148) );
  XOR U3796 ( .A(n4149), .B(n4150), .Z(n4143) );
  AND U3797 ( .A(n488), .B(n4142), .Z(n4150) );
  XNOR U3798 ( .A(n4140), .B(n4149), .Z(n4142) );
  XNOR U3799 ( .A(n4151), .B(n4152), .Z(n4140) );
  AND U3800 ( .A(n492), .B(n4153), .Z(n4152) );
  XOR U3801 ( .A(p_input[613]), .B(n4151), .Z(n4153) );
  XNOR U3802 ( .A(n4154), .B(n4155), .Z(n4151) );
  AND U3803 ( .A(n496), .B(n4156), .Z(n4155) );
  XOR U3804 ( .A(n4157), .B(n4158), .Z(n4149) );
  AND U3805 ( .A(n500), .B(n4159), .Z(n4158) );
  XOR U3806 ( .A(n4160), .B(n4161), .Z(n4146) );
  AND U3807 ( .A(n504), .B(n4159), .Z(n4161) );
  XNOR U3808 ( .A(n4162), .B(n4160), .Z(n4159) );
  IV U3809 ( .A(n4157), .Z(n4162) );
  XOR U3810 ( .A(n4163), .B(n4164), .Z(n4157) );
  AND U3811 ( .A(n507), .B(n4156), .Z(n4164) );
  XNOR U3812 ( .A(n4154), .B(n4163), .Z(n4156) );
  XNOR U3813 ( .A(n4165), .B(n4166), .Z(n4154) );
  AND U3814 ( .A(n511), .B(n4167), .Z(n4166) );
  XOR U3815 ( .A(p_input[645]), .B(n4165), .Z(n4167) );
  XNOR U3816 ( .A(n4168), .B(n4169), .Z(n4165) );
  AND U3817 ( .A(n515), .B(n4170), .Z(n4169) );
  XOR U3818 ( .A(n4171), .B(n4172), .Z(n4163) );
  AND U3819 ( .A(n519), .B(n4173), .Z(n4172) );
  XOR U3820 ( .A(n4174), .B(n4175), .Z(n4160) );
  AND U3821 ( .A(n523), .B(n4173), .Z(n4175) );
  XNOR U3822 ( .A(n4176), .B(n4174), .Z(n4173) );
  IV U3823 ( .A(n4171), .Z(n4176) );
  XOR U3824 ( .A(n4177), .B(n4178), .Z(n4171) );
  AND U3825 ( .A(n526), .B(n4170), .Z(n4178) );
  XNOR U3826 ( .A(n4168), .B(n4177), .Z(n4170) );
  XNOR U3827 ( .A(n4179), .B(n4180), .Z(n4168) );
  AND U3828 ( .A(n530), .B(n4181), .Z(n4180) );
  XOR U3829 ( .A(p_input[677]), .B(n4179), .Z(n4181) );
  XNOR U3830 ( .A(n4182), .B(n4183), .Z(n4179) );
  AND U3831 ( .A(n534), .B(n4184), .Z(n4183) );
  XOR U3832 ( .A(n4185), .B(n4186), .Z(n4177) );
  AND U3833 ( .A(n538), .B(n4187), .Z(n4186) );
  XOR U3834 ( .A(n4188), .B(n4189), .Z(n4174) );
  AND U3835 ( .A(n542), .B(n4187), .Z(n4189) );
  XNOR U3836 ( .A(n4190), .B(n4188), .Z(n4187) );
  IV U3837 ( .A(n4185), .Z(n4190) );
  XOR U3838 ( .A(n4191), .B(n4192), .Z(n4185) );
  AND U3839 ( .A(n545), .B(n4184), .Z(n4192) );
  XNOR U3840 ( .A(n4182), .B(n4191), .Z(n4184) );
  XNOR U3841 ( .A(n4193), .B(n4194), .Z(n4182) );
  AND U3842 ( .A(n549), .B(n4195), .Z(n4194) );
  XOR U3843 ( .A(p_input[709]), .B(n4193), .Z(n4195) );
  XNOR U3844 ( .A(n4196), .B(n4197), .Z(n4193) );
  AND U3845 ( .A(n553), .B(n4198), .Z(n4197) );
  XOR U3846 ( .A(n4199), .B(n4200), .Z(n4191) );
  AND U3847 ( .A(n557), .B(n4201), .Z(n4200) );
  XOR U3848 ( .A(n4202), .B(n4203), .Z(n4188) );
  AND U3849 ( .A(n561), .B(n4201), .Z(n4203) );
  XNOR U3850 ( .A(n4204), .B(n4202), .Z(n4201) );
  IV U3851 ( .A(n4199), .Z(n4204) );
  XOR U3852 ( .A(n4205), .B(n4206), .Z(n4199) );
  AND U3853 ( .A(n564), .B(n4198), .Z(n4206) );
  XNOR U3854 ( .A(n4196), .B(n4205), .Z(n4198) );
  XNOR U3855 ( .A(n4207), .B(n4208), .Z(n4196) );
  AND U3856 ( .A(n568), .B(n4209), .Z(n4208) );
  XOR U3857 ( .A(p_input[741]), .B(n4207), .Z(n4209) );
  XNOR U3858 ( .A(n4210), .B(n4211), .Z(n4207) );
  AND U3859 ( .A(n572), .B(n4212), .Z(n4211) );
  XOR U3860 ( .A(n4213), .B(n4214), .Z(n4205) );
  AND U3861 ( .A(n576), .B(n4215), .Z(n4214) );
  XOR U3862 ( .A(n4216), .B(n4217), .Z(n4202) );
  AND U3863 ( .A(n580), .B(n4215), .Z(n4217) );
  XNOR U3864 ( .A(n4218), .B(n4216), .Z(n4215) );
  IV U3865 ( .A(n4213), .Z(n4218) );
  XOR U3866 ( .A(n4219), .B(n4220), .Z(n4213) );
  AND U3867 ( .A(n583), .B(n4212), .Z(n4220) );
  XNOR U3868 ( .A(n4210), .B(n4219), .Z(n4212) );
  XNOR U3869 ( .A(n4221), .B(n4222), .Z(n4210) );
  AND U3870 ( .A(n587), .B(n4223), .Z(n4222) );
  XOR U3871 ( .A(p_input[773]), .B(n4221), .Z(n4223) );
  XNOR U3872 ( .A(n4224), .B(n4225), .Z(n4221) );
  AND U3873 ( .A(n591), .B(n4226), .Z(n4225) );
  XOR U3874 ( .A(n4227), .B(n4228), .Z(n4219) );
  AND U3875 ( .A(n595), .B(n4229), .Z(n4228) );
  XOR U3876 ( .A(n4230), .B(n4231), .Z(n4216) );
  AND U3877 ( .A(n599), .B(n4229), .Z(n4231) );
  XNOR U3878 ( .A(n4232), .B(n4230), .Z(n4229) );
  IV U3879 ( .A(n4227), .Z(n4232) );
  XOR U3880 ( .A(n4233), .B(n4234), .Z(n4227) );
  AND U3881 ( .A(n602), .B(n4226), .Z(n4234) );
  XNOR U3882 ( .A(n4224), .B(n4233), .Z(n4226) );
  XNOR U3883 ( .A(n4235), .B(n4236), .Z(n4224) );
  AND U3884 ( .A(n606), .B(n4237), .Z(n4236) );
  XOR U3885 ( .A(p_input[805]), .B(n4235), .Z(n4237) );
  XNOR U3886 ( .A(n4238), .B(n4239), .Z(n4235) );
  AND U3887 ( .A(n610), .B(n4240), .Z(n4239) );
  XOR U3888 ( .A(n4241), .B(n4242), .Z(n4233) );
  AND U3889 ( .A(n614), .B(n4243), .Z(n4242) );
  XOR U3890 ( .A(n4244), .B(n4245), .Z(n4230) );
  AND U3891 ( .A(n618), .B(n4243), .Z(n4245) );
  XNOR U3892 ( .A(n4246), .B(n4244), .Z(n4243) );
  IV U3893 ( .A(n4241), .Z(n4246) );
  XOR U3894 ( .A(n4247), .B(n4248), .Z(n4241) );
  AND U3895 ( .A(n621), .B(n4240), .Z(n4248) );
  XNOR U3896 ( .A(n4238), .B(n4247), .Z(n4240) );
  XNOR U3897 ( .A(n4249), .B(n4250), .Z(n4238) );
  AND U3898 ( .A(n625), .B(n4251), .Z(n4250) );
  XOR U3899 ( .A(p_input[837]), .B(n4249), .Z(n4251) );
  XNOR U3900 ( .A(n4252), .B(n4253), .Z(n4249) );
  AND U3901 ( .A(n629), .B(n4254), .Z(n4253) );
  XOR U3902 ( .A(n4255), .B(n4256), .Z(n4247) );
  AND U3903 ( .A(n633), .B(n4257), .Z(n4256) );
  XOR U3904 ( .A(n4258), .B(n4259), .Z(n4244) );
  AND U3905 ( .A(n637), .B(n4257), .Z(n4259) );
  XNOR U3906 ( .A(n4260), .B(n4258), .Z(n4257) );
  IV U3907 ( .A(n4255), .Z(n4260) );
  XOR U3908 ( .A(n4261), .B(n4262), .Z(n4255) );
  AND U3909 ( .A(n640), .B(n4254), .Z(n4262) );
  XNOR U3910 ( .A(n4252), .B(n4261), .Z(n4254) );
  XNOR U3911 ( .A(n4263), .B(n4264), .Z(n4252) );
  AND U3912 ( .A(n644), .B(n4265), .Z(n4264) );
  XOR U3913 ( .A(p_input[869]), .B(n4263), .Z(n4265) );
  XNOR U3914 ( .A(n4266), .B(n4267), .Z(n4263) );
  AND U3915 ( .A(n648), .B(n4268), .Z(n4267) );
  XOR U3916 ( .A(n4269), .B(n4270), .Z(n4261) );
  AND U3917 ( .A(n652), .B(n4271), .Z(n4270) );
  XOR U3918 ( .A(n4272), .B(n4273), .Z(n4258) );
  AND U3919 ( .A(n656), .B(n4271), .Z(n4273) );
  XNOR U3920 ( .A(n4274), .B(n4272), .Z(n4271) );
  IV U3921 ( .A(n4269), .Z(n4274) );
  XOR U3922 ( .A(n4275), .B(n4276), .Z(n4269) );
  AND U3923 ( .A(n659), .B(n4268), .Z(n4276) );
  XNOR U3924 ( .A(n4266), .B(n4275), .Z(n4268) );
  XNOR U3925 ( .A(n4277), .B(n4278), .Z(n4266) );
  AND U3926 ( .A(n663), .B(n4279), .Z(n4278) );
  XOR U3927 ( .A(p_input[901]), .B(n4277), .Z(n4279) );
  XNOR U3928 ( .A(n4280), .B(n4281), .Z(n4277) );
  AND U3929 ( .A(n667), .B(n4282), .Z(n4281) );
  XOR U3930 ( .A(n4283), .B(n4284), .Z(n4275) );
  AND U3931 ( .A(n671), .B(n4285), .Z(n4284) );
  XOR U3932 ( .A(n4286), .B(n4287), .Z(n4272) );
  AND U3933 ( .A(n675), .B(n4285), .Z(n4287) );
  XNOR U3934 ( .A(n4288), .B(n4286), .Z(n4285) );
  IV U3935 ( .A(n4283), .Z(n4288) );
  XOR U3936 ( .A(n4289), .B(n4290), .Z(n4283) );
  AND U3937 ( .A(n678), .B(n4282), .Z(n4290) );
  XNOR U3938 ( .A(n4280), .B(n4289), .Z(n4282) );
  XNOR U3939 ( .A(n4291), .B(n4292), .Z(n4280) );
  AND U3940 ( .A(n682), .B(n4293), .Z(n4292) );
  XOR U3941 ( .A(p_input[933]), .B(n4291), .Z(n4293) );
  XNOR U3942 ( .A(n4294), .B(n4295), .Z(n4291) );
  AND U3943 ( .A(n686), .B(n4296), .Z(n4295) );
  XOR U3944 ( .A(n4297), .B(n4298), .Z(n4289) );
  AND U3945 ( .A(n690), .B(n4299), .Z(n4298) );
  XOR U3946 ( .A(n4300), .B(n4301), .Z(n4286) );
  AND U3947 ( .A(n694), .B(n4299), .Z(n4301) );
  XNOR U3948 ( .A(n4302), .B(n4300), .Z(n4299) );
  IV U3949 ( .A(n4297), .Z(n4302) );
  XOR U3950 ( .A(n4303), .B(n4304), .Z(n4297) );
  AND U3951 ( .A(n697), .B(n4296), .Z(n4304) );
  XNOR U3952 ( .A(n4294), .B(n4303), .Z(n4296) );
  XNOR U3953 ( .A(n4305), .B(n4306), .Z(n4294) );
  AND U3954 ( .A(n701), .B(n4307), .Z(n4306) );
  XOR U3955 ( .A(p_input[965]), .B(n4305), .Z(n4307) );
  XNOR U3956 ( .A(n4308), .B(n4309), .Z(n4305) );
  AND U3957 ( .A(n705), .B(n4310), .Z(n4309) );
  XOR U3958 ( .A(n4311), .B(n4312), .Z(n4303) );
  AND U3959 ( .A(n709), .B(n4313), .Z(n4312) );
  XOR U3960 ( .A(n4314), .B(n4315), .Z(n4300) );
  AND U3961 ( .A(n713), .B(n4313), .Z(n4315) );
  XNOR U3962 ( .A(n4316), .B(n4314), .Z(n4313) );
  IV U3963 ( .A(n4311), .Z(n4316) );
  XOR U3964 ( .A(n4317), .B(n4318), .Z(n4311) );
  AND U3965 ( .A(n716), .B(n4310), .Z(n4318) );
  XNOR U3966 ( .A(n4308), .B(n4317), .Z(n4310) );
  XNOR U3967 ( .A(n4319), .B(n4320), .Z(n4308) );
  AND U3968 ( .A(n720), .B(n4321), .Z(n4320) );
  XOR U3969 ( .A(p_input[997]), .B(n4319), .Z(n4321) );
  XNOR U3970 ( .A(n4322), .B(n4323), .Z(n4319) );
  AND U3971 ( .A(n724), .B(n4324), .Z(n4323) );
  XOR U3972 ( .A(n4325), .B(n4326), .Z(n4317) );
  AND U3973 ( .A(n728), .B(n4327), .Z(n4326) );
  XOR U3974 ( .A(n4328), .B(n4329), .Z(n4314) );
  AND U3975 ( .A(n732), .B(n4327), .Z(n4329) );
  XNOR U3976 ( .A(n4330), .B(n4328), .Z(n4327) );
  IV U3977 ( .A(n4325), .Z(n4330) );
  XOR U3978 ( .A(n4331), .B(n4332), .Z(n4325) );
  AND U3979 ( .A(n735), .B(n4324), .Z(n4332) );
  XNOR U3980 ( .A(n4322), .B(n4331), .Z(n4324) );
  XNOR U3981 ( .A(n4333), .B(n4334), .Z(n4322) );
  AND U3982 ( .A(n739), .B(n4335), .Z(n4334) );
  XOR U3983 ( .A(p_input[1029]), .B(n4333), .Z(n4335) );
  XNOR U3984 ( .A(n4336), .B(n4337), .Z(n4333) );
  AND U3985 ( .A(n743), .B(n4338), .Z(n4337) );
  XOR U3986 ( .A(n4339), .B(n4340), .Z(n4331) );
  AND U3987 ( .A(n747), .B(n4341), .Z(n4340) );
  XOR U3988 ( .A(n4342), .B(n4343), .Z(n4328) );
  AND U3989 ( .A(n751), .B(n4341), .Z(n4343) );
  XNOR U3990 ( .A(n4344), .B(n4342), .Z(n4341) );
  IV U3991 ( .A(n4339), .Z(n4344) );
  XOR U3992 ( .A(n4345), .B(n4346), .Z(n4339) );
  AND U3993 ( .A(n754), .B(n4338), .Z(n4346) );
  XNOR U3994 ( .A(n4336), .B(n4345), .Z(n4338) );
  XNOR U3995 ( .A(n4347), .B(n4348), .Z(n4336) );
  AND U3996 ( .A(n758), .B(n4349), .Z(n4348) );
  XOR U3997 ( .A(p_input[1061]), .B(n4347), .Z(n4349) );
  XNOR U3998 ( .A(n4350), .B(n4351), .Z(n4347) );
  AND U3999 ( .A(n762), .B(n4352), .Z(n4351) );
  XOR U4000 ( .A(n4353), .B(n4354), .Z(n4345) );
  AND U4001 ( .A(n766), .B(n4355), .Z(n4354) );
  XOR U4002 ( .A(n4356), .B(n4357), .Z(n4342) );
  AND U4003 ( .A(n770), .B(n4355), .Z(n4357) );
  XNOR U4004 ( .A(n4358), .B(n4356), .Z(n4355) );
  IV U4005 ( .A(n4353), .Z(n4358) );
  XOR U4006 ( .A(n4359), .B(n4360), .Z(n4353) );
  AND U4007 ( .A(n773), .B(n4352), .Z(n4360) );
  XNOR U4008 ( .A(n4350), .B(n4359), .Z(n4352) );
  XNOR U4009 ( .A(n4361), .B(n4362), .Z(n4350) );
  AND U4010 ( .A(n777), .B(n4363), .Z(n4362) );
  XOR U4011 ( .A(p_input[1093]), .B(n4361), .Z(n4363) );
  XNOR U4012 ( .A(n4364), .B(n4365), .Z(n4361) );
  AND U4013 ( .A(n781), .B(n4366), .Z(n4365) );
  XOR U4014 ( .A(n4367), .B(n4368), .Z(n4359) );
  AND U4015 ( .A(n785), .B(n4369), .Z(n4368) );
  XOR U4016 ( .A(n4370), .B(n4371), .Z(n4356) );
  AND U4017 ( .A(n789), .B(n4369), .Z(n4371) );
  XNOR U4018 ( .A(n4372), .B(n4370), .Z(n4369) );
  IV U4019 ( .A(n4367), .Z(n4372) );
  XOR U4020 ( .A(n4373), .B(n4374), .Z(n4367) );
  AND U4021 ( .A(n792), .B(n4366), .Z(n4374) );
  XNOR U4022 ( .A(n4364), .B(n4373), .Z(n4366) );
  XNOR U4023 ( .A(n4375), .B(n4376), .Z(n4364) );
  AND U4024 ( .A(n796), .B(n4377), .Z(n4376) );
  XOR U4025 ( .A(p_input[1125]), .B(n4375), .Z(n4377) );
  XNOR U4026 ( .A(n4378), .B(n4379), .Z(n4375) );
  AND U4027 ( .A(n800), .B(n4380), .Z(n4379) );
  XOR U4028 ( .A(n4381), .B(n4382), .Z(n4373) );
  AND U4029 ( .A(n804), .B(n4383), .Z(n4382) );
  XOR U4030 ( .A(n4384), .B(n4385), .Z(n4370) );
  AND U4031 ( .A(n808), .B(n4383), .Z(n4385) );
  XNOR U4032 ( .A(n4386), .B(n4384), .Z(n4383) );
  IV U4033 ( .A(n4381), .Z(n4386) );
  XOR U4034 ( .A(n4387), .B(n4388), .Z(n4381) );
  AND U4035 ( .A(n811), .B(n4380), .Z(n4388) );
  XNOR U4036 ( .A(n4378), .B(n4387), .Z(n4380) );
  XNOR U4037 ( .A(n4389), .B(n4390), .Z(n4378) );
  AND U4038 ( .A(n815), .B(n4391), .Z(n4390) );
  XOR U4039 ( .A(p_input[1157]), .B(n4389), .Z(n4391) );
  XNOR U4040 ( .A(n4392), .B(n4393), .Z(n4389) );
  AND U4041 ( .A(n819), .B(n4394), .Z(n4393) );
  XOR U4042 ( .A(n4395), .B(n4396), .Z(n4387) );
  AND U4043 ( .A(n823), .B(n4397), .Z(n4396) );
  XOR U4044 ( .A(n4398), .B(n4399), .Z(n4384) );
  AND U4045 ( .A(n827), .B(n4397), .Z(n4399) );
  XNOR U4046 ( .A(n4400), .B(n4398), .Z(n4397) );
  IV U4047 ( .A(n4395), .Z(n4400) );
  XOR U4048 ( .A(n4401), .B(n4402), .Z(n4395) );
  AND U4049 ( .A(n830), .B(n4394), .Z(n4402) );
  XNOR U4050 ( .A(n4392), .B(n4401), .Z(n4394) );
  XNOR U4051 ( .A(n4403), .B(n4404), .Z(n4392) );
  AND U4052 ( .A(n834), .B(n4405), .Z(n4404) );
  XOR U4053 ( .A(p_input[1189]), .B(n4403), .Z(n4405) );
  XNOR U4054 ( .A(n4406), .B(n4407), .Z(n4403) );
  AND U4055 ( .A(n838), .B(n4408), .Z(n4407) );
  XOR U4056 ( .A(n4409), .B(n4410), .Z(n4401) );
  AND U4057 ( .A(n842), .B(n4411), .Z(n4410) );
  XOR U4058 ( .A(n4412), .B(n4413), .Z(n4398) );
  AND U4059 ( .A(n846), .B(n4411), .Z(n4413) );
  XNOR U4060 ( .A(n4414), .B(n4412), .Z(n4411) );
  IV U4061 ( .A(n4409), .Z(n4414) );
  XOR U4062 ( .A(n4415), .B(n4416), .Z(n4409) );
  AND U4063 ( .A(n849), .B(n4408), .Z(n4416) );
  XNOR U4064 ( .A(n4406), .B(n4415), .Z(n4408) );
  XNOR U4065 ( .A(n4417), .B(n4418), .Z(n4406) );
  AND U4066 ( .A(n853), .B(n4419), .Z(n4418) );
  XOR U4067 ( .A(p_input[1221]), .B(n4417), .Z(n4419) );
  XNOR U4068 ( .A(n4420), .B(n4421), .Z(n4417) );
  AND U4069 ( .A(n857), .B(n4422), .Z(n4421) );
  XOR U4070 ( .A(n4423), .B(n4424), .Z(n4415) );
  AND U4071 ( .A(n861), .B(n4425), .Z(n4424) );
  XOR U4072 ( .A(n4426), .B(n4427), .Z(n4412) );
  AND U4073 ( .A(n865), .B(n4425), .Z(n4427) );
  XNOR U4074 ( .A(n4428), .B(n4426), .Z(n4425) );
  IV U4075 ( .A(n4423), .Z(n4428) );
  XOR U4076 ( .A(n4429), .B(n4430), .Z(n4423) );
  AND U4077 ( .A(n868), .B(n4422), .Z(n4430) );
  XNOR U4078 ( .A(n4420), .B(n4429), .Z(n4422) );
  XNOR U4079 ( .A(n4431), .B(n4432), .Z(n4420) );
  AND U4080 ( .A(n872), .B(n4433), .Z(n4432) );
  XOR U4081 ( .A(p_input[1253]), .B(n4431), .Z(n4433) );
  XNOR U4082 ( .A(n4434), .B(n4435), .Z(n4431) );
  AND U4083 ( .A(n876), .B(n4436), .Z(n4435) );
  XOR U4084 ( .A(n4437), .B(n4438), .Z(n4429) );
  AND U4085 ( .A(n880), .B(n4439), .Z(n4438) );
  XOR U4086 ( .A(n4440), .B(n4441), .Z(n4426) );
  AND U4087 ( .A(n884), .B(n4439), .Z(n4441) );
  XNOR U4088 ( .A(n4442), .B(n4440), .Z(n4439) );
  IV U4089 ( .A(n4437), .Z(n4442) );
  XOR U4090 ( .A(n4443), .B(n4444), .Z(n4437) );
  AND U4091 ( .A(n887), .B(n4436), .Z(n4444) );
  XNOR U4092 ( .A(n4434), .B(n4443), .Z(n4436) );
  XNOR U4093 ( .A(n4445), .B(n4446), .Z(n4434) );
  AND U4094 ( .A(n891), .B(n4447), .Z(n4446) );
  XOR U4095 ( .A(p_input[1285]), .B(n4445), .Z(n4447) );
  XNOR U4096 ( .A(n4448), .B(n4449), .Z(n4445) );
  AND U4097 ( .A(n895), .B(n4450), .Z(n4449) );
  XOR U4098 ( .A(n4451), .B(n4452), .Z(n4443) );
  AND U4099 ( .A(n899), .B(n4453), .Z(n4452) );
  XOR U4100 ( .A(n4454), .B(n4455), .Z(n4440) );
  AND U4101 ( .A(n903), .B(n4453), .Z(n4455) );
  XNOR U4102 ( .A(n4456), .B(n4454), .Z(n4453) );
  IV U4103 ( .A(n4451), .Z(n4456) );
  XOR U4104 ( .A(n4457), .B(n4458), .Z(n4451) );
  AND U4105 ( .A(n906), .B(n4450), .Z(n4458) );
  XNOR U4106 ( .A(n4448), .B(n4457), .Z(n4450) );
  XNOR U4107 ( .A(n4459), .B(n4460), .Z(n4448) );
  AND U4108 ( .A(n910), .B(n4461), .Z(n4460) );
  XOR U4109 ( .A(p_input[1317]), .B(n4459), .Z(n4461) );
  XNOR U4110 ( .A(n4462), .B(n4463), .Z(n4459) );
  AND U4111 ( .A(n914), .B(n4464), .Z(n4463) );
  XOR U4112 ( .A(n4465), .B(n4466), .Z(n4457) );
  AND U4113 ( .A(n918), .B(n4467), .Z(n4466) );
  XOR U4114 ( .A(n4468), .B(n4469), .Z(n4454) );
  AND U4115 ( .A(n922), .B(n4467), .Z(n4469) );
  XNOR U4116 ( .A(n4470), .B(n4468), .Z(n4467) );
  IV U4117 ( .A(n4465), .Z(n4470) );
  XOR U4118 ( .A(n4471), .B(n4472), .Z(n4465) );
  AND U4119 ( .A(n925), .B(n4464), .Z(n4472) );
  XNOR U4120 ( .A(n4462), .B(n4471), .Z(n4464) );
  XNOR U4121 ( .A(n4473), .B(n4474), .Z(n4462) );
  AND U4122 ( .A(n929), .B(n4475), .Z(n4474) );
  XOR U4123 ( .A(p_input[1349]), .B(n4473), .Z(n4475) );
  XNOR U4124 ( .A(n4476), .B(n4477), .Z(n4473) );
  AND U4125 ( .A(n933), .B(n4478), .Z(n4477) );
  XOR U4126 ( .A(n4479), .B(n4480), .Z(n4471) );
  AND U4127 ( .A(n937), .B(n4481), .Z(n4480) );
  XOR U4128 ( .A(n4482), .B(n4483), .Z(n4468) );
  AND U4129 ( .A(n941), .B(n4481), .Z(n4483) );
  XNOR U4130 ( .A(n4484), .B(n4482), .Z(n4481) );
  IV U4131 ( .A(n4479), .Z(n4484) );
  XOR U4132 ( .A(n4485), .B(n4486), .Z(n4479) );
  AND U4133 ( .A(n944), .B(n4478), .Z(n4486) );
  XNOR U4134 ( .A(n4476), .B(n4485), .Z(n4478) );
  XNOR U4135 ( .A(n4487), .B(n4488), .Z(n4476) );
  AND U4136 ( .A(n948), .B(n4489), .Z(n4488) );
  XOR U4137 ( .A(p_input[1381]), .B(n4487), .Z(n4489) );
  XNOR U4138 ( .A(n4490), .B(n4491), .Z(n4487) );
  AND U4139 ( .A(n952), .B(n4492), .Z(n4491) );
  XOR U4140 ( .A(n4493), .B(n4494), .Z(n4485) );
  AND U4141 ( .A(n956), .B(n4495), .Z(n4494) );
  XOR U4142 ( .A(n4496), .B(n4497), .Z(n4482) );
  AND U4143 ( .A(n960), .B(n4495), .Z(n4497) );
  XNOR U4144 ( .A(n4498), .B(n4496), .Z(n4495) );
  IV U4145 ( .A(n4493), .Z(n4498) );
  XOR U4146 ( .A(n4499), .B(n4500), .Z(n4493) );
  AND U4147 ( .A(n963), .B(n4492), .Z(n4500) );
  XNOR U4148 ( .A(n4490), .B(n4499), .Z(n4492) );
  XNOR U4149 ( .A(n4501), .B(n4502), .Z(n4490) );
  AND U4150 ( .A(n967), .B(n4503), .Z(n4502) );
  XOR U4151 ( .A(p_input[1413]), .B(n4501), .Z(n4503) );
  XNOR U4152 ( .A(n4504), .B(n4505), .Z(n4501) );
  AND U4153 ( .A(n971), .B(n4506), .Z(n4505) );
  XOR U4154 ( .A(n4507), .B(n4508), .Z(n4499) );
  AND U4155 ( .A(n975), .B(n4509), .Z(n4508) );
  XOR U4156 ( .A(n4510), .B(n4511), .Z(n4496) );
  AND U4157 ( .A(n979), .B(n4509), .Z(n4511) );
  XNOR U4158 ( .A(n4512), .B(n4510), .Z(n4509) );
  IV U4159 ( .A(n4507), .Z(n4512) );
  XOR U4160 ( .A(n4513), .B(n4514), .Z(n4507) );
  AND U4161 ( .A(n982), .B(n4506), .Z(n4514) );
  XNOR U4162 ( .A(n4504), .B(n4513), .Z(n4506) );
  XNOR U4163 ( .A(n4515), .B(n4516), .Z(n4504) );
  AND U4164 ( .A(n986), .B(n4517), .Z(n4516) );
  XOR U4165 ( .A(p_input[1445]), .B(n4515), .Z(n4517) );
  XNOR U4166 ( .A(n4518), .B(n4519), .Z(n4515) );
  AND U4167 ( .A(n990), .B(n4520), .Z(n4519) );
  XOR U4168 ( .A(n4521), .B(n4522), .Z(n4513) );
  AND U4169 ( .A(n994), .B(n4523), .Z(n4522) );
  XOR U4170 ( .A(n4524), .B(n4525), .Z(n4510) );
  AND U4171 ( .A(n998), .B(n4523), .Z(n4525) );
  XNOR U4172 ( .A(n4526), .B(n4524), .Z(n4523) );
  IV U4173 ( .A(n4521), .Z(n4526) );
  XOR U4174 ( .A(n4527), .B(n4528), .Z(n4521) );
  AND U4175 ( .A(n1001), .B(n4520), .Z(n4528) );
  XNOR U4176 ( .A(n4518), .B(n4527), .Z(n4520) );
  XNOR U4177 ( .A(n4529), .B(n4530), .Z(n4518) );
  AND U4178 ( .A(n1005), .B(n4531), .Z(n4530) );
  XOR U4179 ( .A(p_input[1477]), .B(n4529), .Z(n4531) );
  XNOR U4180 ( .A(n4532), .B(n4533), .Z(n4529) );
  AND U4181 ( .A(n1009), .B(n4534), .Z(n4533) );
  XOR U4182 ( .A(n4535), .B(n4536), .Z(n4527) );
  AND U4183 ( .A(n1013), .B(n4537), .Z(n4536) );
  XOR U4184 ( .A(n4538), .B(n4539), .Z(n4524) );
  AND U4185 ( .A(n1017), .B(n4537), .Z(n4539) );
  XNOR U4186 ( .A(n4540), .B(n4538), .Z(n4537) );
  IV U4187 ( .A(n4535), .Z(n4540) );
  XOR U4188 ( .A(n4541), .B(n4542), .Z(n4535) );
  AND U4189 ( .A(n1020), .B(n4534), .Z(n4542) );
  XNOR U4190 ( .A(n4532), .B(n4541), .Z(n4534) );
  XNOR U4191 ( .A(n4543), .B(n4544), .Z(n4532) );
  AND U4192 ( .A(n1024), .B(n4545), .Z(n4544) );
  XOR U4193 ( .A(p_input[1509]), .B(n4543), .Z(n4545) );
  XNOR U4194 ( .A(n4546), .B(n4547), .Z(n4543) );
  AND U4195 ( .A(n1028), .B(n4548), .Z(n4547) );
  XOR U4196 ( .A(n4549), .B(n4550), .Z(n4541) );
  AND U4197 ( .A(n1032), .B(n4551), .Z(n4550) );
  XOR U4198 ( .A(n4552), .B(n4553), .Z(n4538) );
  AND U4199 ( .A(n1036), .B(n4551), .Z(n4553) );
  XNOR U4200 ( .A(n4554), .B(n4552), .Z(n4551) );
  IV U4201 ( .A(n4549), .Z(n4554) );
  XOR U4202 ( .A(n4555), .B(n4556), .Z(n4549) );
  AND U4203 ( .A(n1039), .B(n4548), .Z(n4556) );
  XNOR U4204 ( .A(n4546), .B(n4555), .Z(n4548) );
  XNOR U4205 ( .A(n4557), .B(n4558), .Z(n4546) );
  AND U4206 ( .A(n1043), .B(n4559), .Z(n4558) );
  XOR U4207 ( .A(p_input[1541]), .B(n4557), .Z(n4559) );
  XNOR U4208 ( .A(n4560), .B(n4561), .Z(n4557) );
  AND U4209 ( .A(n1047), .B(n4562), .Z(n4561) );
  XOR U4210 ( .A(n4563), .B(n4564), .Z(n4555) );
  AND U4211 ( .A(n1051), .B(n4565), .Z(n4564) );
  XOR U4212 ( .A(n4566), .B(n4567), .Z(n4552) );
  AND U4213 ( .A(n1055), .B(n4565), .Z(n4567) );
  XNOR U4214 ( .A(n4568), .B(n4566), .Z(n4565) );
  IV U4215 ( .A(n4563), .Z(n4568) );
  XOR U4216 ( .A(n4569), .B(n4570), .Z(n4563) );
  AND U4217 ( .A(n1058), .B(n4562), .Z(n4570) );
  XNOR U4218 ( .A(n4560), .B(n4569), .Z(n4562) );
  XNOR U4219 ( .A(n4571), .B(n4572), .Z(n4560) );
  AND U4220 ( .A(n1062), .B(n4573), .Z(n4572) );
  XOR U4221 ( .A(p_input[1573]), .B(n4571), .Z(n4573) );
  XNOR U4222 ( .A(n4574), .B(n4575), .Z(n4571) );
  AND U4223 ( .A(n1066), .B(n4576), .Z(n4575) );
  XOR U4224 ( .A(n4577), .B(n4578), .Z(n4569) );
  AND U4225 ( .A(n1070), .B(n4579), .Z(n4578) );
  XOR U4226 ( .A(n4580), .B(n4581), .Z(n4566) );
  AND U4227 ( .A(n1074), .B(n4579), .Z(n4581) );
  XNOR U4228 ( .A(n4582), .B(n4580), .Z(n4579) );
  IV U4229 ( .A(n4577), .Z(n4582) );
  XOR U4230 ( .A(n4583), .B(n4584), .Z(n4577) );
  AND U4231 ( .A(n1077), .B(n4576), .Z(n4584) );
  XNOR U4232 ( .A(n4574), .B(n4583), .Z(n4576) );
  XNOR U4233 ( .A(n4585), .B(n4586), .Z(n4574) );
  AND U4234 ( .A(n1081), .B(n4587), .Z(n4586) );
  XOR U4235 ( .A(p_input[1605]), .B(n4585), .Z(n4587) );
  XNOR U4236 ( .A(n4588), .B(n4589), .Z(n4585) );
  AND U4237 ( .A(n1085), .B(n4590), .Z(n4589) );
  XOR U4238 ( .A(n4591), .B(n4592), .Z(n4583) );
  AND U4239 ( .A(n1089), .B(n4593), .Z(n4592) );
  XOR U4240 ( .A(n4594), .B(n4595), .Z(n4580) );
  AND U4241 ( .A(n1093), .B(n4593), .Z(n4595) );
  XNOR U4242 ( .A(n4596), .B(n4594), .Z(n4593) );
  IV U4243 ( .A(n4591), .Z(n4596) );
  XOR U4244 ( .A(n4597), .B(n4598), .Z(n4591) );
  AND U4245 ( .A(n1096), .B(n4590), .Z(n4598) );
  XNOR U4246 ( .A(n4588), .B(n4597), .Z(n4590) );
  XNOR U4247 ( .A(n4599), .B(n4600), .Z(n4588) );
  AND U4248 ( .A(n1100), .B(n4601), .Z(n4600) );
  XOR U4249 ( .A(p_input[1637]), .B(n4599), .Z(n4601) );
  XNOR U4250 ( .A(n4602), .B(n4603), .Z(n4599) );
  AND U4251 ( .A(n1104), .B(n4604), .Z(n4603) );
  XOR U4252 ( .A(n4605), .B(n4606), .Z(n4597) );
  AND U4253 ( .A(n1108), .B(n4607), .Z(n4606) );
  XOR U4254 ( .A(n4608), .B(n4609), .Z(n4594) );
  AND U4255 ( .A(n1112), .B(n4607), .Z(n4609) );
  XNOR U4256 ( .A(n4610), .B(n4608), .Z(n4607) );
  IV U4257 ( .A(n4605), .Z(n4610) );
  XOR U4258 ( .A(n4611), .B(n4612), .Z(n4605) );
  AND U4259 ( .A(n1115), .B(n4604), .Z(n4612) );
  XNOR U4260 ( .A(n4602), .B(n4611), .Z(n4604) );
  XNOR U4261 ( .A(n4613), .B(n4614), .Z(n4602) );
  AND U4262 ( .A(n1119), .B(n4615), .Z(n4614) );
  XOR U4263 ( .A(p_input[1669]), .B(n4613), .Z(n4615) );
  XNOR U4264 ( .A(n4616), .B(n4617), .Z(n4613) );
  AND U4265 ( .A(n1123), .B(n4618), .Z(n4617) );
  XOR U4266 ( .A(n4619), .B(n4620), .Z(n4611) );
  AND U4267 ( .A(n1127), .B(n4621), .Z(n4620) );
  XOR U4268 ( .A(n4622), .B(n4623), .Z(n4608) );
  AND U4269 ( .A(n1131), .B(n4621), .Z(n4623) );
  XNOR U4270 ( .A(n4624), .B(n4622), .Z(n4621) );
  IV U4271 ( .A(n4619), .Z(n4624) );
  XOR U4272 ( .A(n4625), .B(n4626), .Z(n4619) );
  AND U4273 ( .A(n1134), .B(n4618), .Z(n4626) );
  XNOR U4274 ( .A(n4616), .B(n4625), .Z(n4618) );
  XNOR U4275 ( .A(n4627), .B(n4628), .Z(n4616) );
  AND U4276 ( .A(n1138), .B(n4629), .Z(n4628) );
  XOR U4277 ( .A(p_input[1701]), .B(n4627), .Z(n4629) );
  XNOR U4278 ( .A(n4630), .B(n4631), .Z(n4627) );
  AND U4279 ( .A(n1142), .B(n4632), .Z(n4631) );
  XOR U4280 ( .A(n4633), .B(n4634), .Z(n4625) );
  AND U4281 ( .A(n1146), .B(n4635), .Z(n4634) );
  XOR U4282 ( .A(n4636), .B(n4637), .Z(n4622) );
  AND U4283 ( .A(n1150), .B(n4635), .Z(n4637) );
  XNOR U4284 ( .A(n4638), .B(n4636), .Z(n4635) );
  IV U4285 ( .A(n4633), .Z(n4638) );
  XOR U4286 ( .A(n4639), .B(n4640), .Z(n4633) );
  AND U4287 ( .A(n1153), .B(n4632), .Z(n4640) );
  XNOR U4288 ( .A(n4630), .B(n4639), .Z(n4632) );
  XNOR U4289 ( .A(n4641), .B(n4642), .Z(n4630) );
  AND U4290 ( .A(n1157), .B(n4643), .Z(n4642) );
  XOR U4291 ( .A(p_input[1733]), .B(n4641), .Z(n4643) );
  XNOR U4292 ( .A(n4644), .B(n4645), .Z(n4641) );
  AND U4293 ( .A(n1161), .B(n4646), .Z(n4645) );
  XOR U4294 ( .A(n4647), .B(n4648), .Z(n4639) );
  AND U4295 ( .A(n1165), .B(n4649), .Z(n4648) );
  XOR U4296 ( .A(n4650), .B(n4651), .Z(n4636) );
  AND U4297 ( .A(n1169), .B(n4649), .Z(n4651) );
  XNOR U4298 ( .A(n4652), .B(n4650), .Z(n4649) );
  IV U4299 ( .A(n4647), .Z(n4652) );
  XOR U4300 ( .A(n4653), .B(n4654), .Z(n4647) );
  AND U4301 ( .A(n1172), .B(n4646), .Z(n4654) );
  XNOR U4302 ( .A(n4644), .B(n4653), .Z(n4646) );
  XNOR U4303 ( .A(n4655), .B(n4656), .Z(n4644) );
  AND U4304 ( .A(n1176), .B(n4657), .Z(n4656) );
  XOR U4305 ( .A(p_input[1765]), .B(n4655), .Z(n4657) );
  XNOR U4306 ( .A(n4658), .B(n4659), .Z(n4655) );
  AND U4307 ( .A(n1180), .B(n4660), .Z(n4659) );
  XOR U4308 ( .A(n4661), .B(n4662), .Z(n4653) );
  AND U4309 ( .A(n1184), .B(n4663), .Z(n4662) );
  XOR U4310 ( .A(n4664), .B(n4665), .Z(n4650) );
  AND U4311 ( .A(n1188), .B(n4663), .Z(n4665) );
  XNOR U4312 ( .A(n4666), .B(n4664), .Z(n4663) );
  IV U4313 ( .A(n4661), .Z(n4666) );
  XOR U4314 ( .A(n4667), .B(n4668), .Z(n4661) );
  AND U4315 ( .A(n1191), .B(n4660), .Z(n4668) );
  XNOR U4316 ( .A(n4658), .B(n4667), .Z(n4660) );
  XNOR U4317 ( .A(n4669), .B(n4670), .Z(n4658) );
  AND U4318 ( .A(n1195), .B(n4671), .Z(n4670) );
  XOR U4319 ( .A(p_input[1797]), .B(n4669), .Z(n4671) );
  XNOR U4320 ( .A(n4672), .B(n4673), .Z(n4669) );
  AND U4321 ( .A(n1199), .B(n4674), .Z(n4673) );
  XOR U4322 ( .A(n4675), .B(n4676), .Z(n4667) );
  AND U4323 ( .A(n1203), .B(n4677), .Z(n4676) );
  XOR U4324 ( .A(n4678), .B(n4679), .Z(n4664) );
  AND U4325 ( .A(n1207), .B(n4677), .Z(n4679) );
  XNOR U4326 ( .A(n4680), .B(n4678), .Z(n4677) );
  IV U4327 ( .A(n4675), .Z(n4680) );
  XOR U4328 ( .A(n4681), .B(n4682), .Z(n4675) );
  AND U4329 ( .A(n1210), .B(n4674), .Z(n4682) );
  XNOR U4330 ( .A(n4672), .B(n4681), .Z(n4674) );
  XNOR U4331 ( .A(n4683), .B(n4684), .Z(n4672) );
  AND U4332 ( .A(n1214), .B(n4685), .Z(n4684) );
  XOR U4333 ( .A(p_input[1829]), .B(n4683), .Z(n4685) );
  XNOR U4334 ( .A(n4686), .B(n4687), .Z(n4683) );
  AND U4335 ( .A(n1218), .B(n4688), .Z(n4687) );
  XOR U4336 ( .A(n4689), .B(n4690), .Z(n4681) );
  AND U4337 ( .A(n1222), .B(n4691), .Z(n4690) );
  XOR U4338 ( .A(n4692), .B(n4693), .Z(n4678) );
  AND U4339 ( .A(n1226), .B(n4691), .Z(n4693) );
  XNOR U4340 ( .A(n4694), .B(n4692), .Z(n4691) );
  IV U4341 ( .A(n4689), .Z(n4694) );
  XOR U4342 ( .A(n4695), .B(n4696), .Z(n4689) );
  AND U4343 ( .A(n1229), .B(n4688), .Z(n4696) );
  XNOR U4344 ( .A(n4686), .B(n4695), .Z(n4688) );
  XNOR U4345 ( .A(n4697), .B(n4698), .Z(n4686) );
  AND U4346 ( .A(n1233), .B(n4699), .Z(n4698) );
  XOR U4347 ( .A(p_input[1861]), .B(n4697), .Z(n4699) );
  XNOR U4348 ( .A(n4700), .B(n4701), .Z(n4697) );
  AND U4349 ( .A(n1237), .B(n4702), .Z(n4701) );
  XOR U4350 ( .A(n4703), .B(n4704), .Z(n4695) );
  AND U4351 ( .A(n1241), .B(n4705), .Z(n4704) );
  XOR U4352 ( .A(n4706), .B(n4707), .Z(n4692) );
  AND U4353 ( .A(n1245), .B(n4705), .Z(n4707) );
  XNOR U4354 ( .A(n4708), .B(n4706), .Z(n4705) );
  IV U4355 ( .A(n4703), .Z(n4708) );
  XOR U4356 ( .A(n4709), .B(n4710), .Z(n4703) );
  AND U4357 ( .A(n1248), .B(n4702), .Z(n4710) );
  XNOR U4358 ( .A(n4700), .B(n4709), .Z(n4702) );
  XNOR U4359 ( .A(n4711), .B(n4712), .Z(n4700) );
  AND U4360 ( .A(n1252), .B(n4713), .Z(n4712) );
  XOR U4361 ( .A(p_input[1893]), .B(n4711), .Z(n4713) );
  XNOR U4362 ( .A(n4714), .B(n4715), .Z(n4711) );
  AND U4363 ( .A(n1256), .B(n4716), .Z(n4715) );
  XOR U4364 ( .A(n4717), .B(n4718), .Z(n4709) );
  AND U4365 ( .A(n1260), .B(n4719), .Z(n4718) );
  XOR U4366 ( .A(n4720), .B(n4721), .Z(n4706) );
  AND U4367 ( .A(n1264), .B(n4719), .Z(n4721) );
  XNOR U4368 ( .A(n4722), .B(n4720), .Z(n4719) );
  IV U4369 ( .A(n4717), .Z(n4722) );
  XOR U4370 ( .A(n4723), .B(n4724), .Z(n4717) );
  AND U4371 ( .A(n1267), .B(n4716), .Z(n4724) );
  XNOR U4372 ( .A(n4714), .B(n4723), .Z(n4716) );
  XNOR U4373 ( .A(n4725), .B(n4726), .Z(n4714) );
  AND U4374 ( .A(n1271), .B(n4727), .Z(n4726) );
  XOR U4375 ( .A(p_input[1925]), .B(n4725), .Z(n4727) );
  XOR U4376 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n4728), 
        .Z(n4725) );
  AND U4377 ( .A(n1274), .B(n4729), .Z(n4728) );
  XOR U4378 ( .A(n4730), .B(n4731), .Z(n4723) );
  AND U4379 ( .A(n1278), .B(n4732), .Z(n4731) );
  XOR U4380 ( .A(n4733), .B(n4734), .Z(n4720) );
  AND U4381 ( .A(n1282), .B(n4732), .Z(n4734) );
  XNOR U4382 ( .A(n4735), .B(n4733), .Z(n4732) );
  IV U4383 ( .A(n4730), .Z(n4735) );
  XOR U4384 ( .A(n4736), .B(n4737), .Z(n4730) );
  AND U4385 ( .A(n1285), .B(n4729), .Z(n4737) );
  XOR U4386 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n4736), 
        .Z(n4729) );
  XOR U4387 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(n4738), 
        .Z(n4736) );
  AND U4388 ( .A(n1287), .B(n4739), .Z(n4738) );
  XOR U4389 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n4740), .Z(n4733) );
  AND U4390 ( .A(n1290), .B(n4739), .Z(n4740) );
  XOR U4391 ( .A(n4741), .B(n4742), .Z(n4739) );
  IV U4392 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .Z(n4742) );
  IV U4393 ( .A(\knn_comb_/min_val_out[0][5] ), .Z(n4741) );
  XOR U4394 ( .A(n103), .B(n4743), .Z(o[36]) );
  AND U4395 ( .A(n122), .B(n4744), .Z(n103) );
  XOR U4396 ( .A(n104), .B(n4743), .Z(n4744) );
  XOR U4397 ( .A(n4745), .B(n63), .Z(n4743) );
  AND U4398 ( .A(n125), .B(n4746), .Z(n63) );
  XOR U4399 ( .A(n64), .B(n4745), .Z(n4746) );
  XOR U4400 ( .A(n4747), .B(n4748), .Z(n64) );
  AND U4401 ( .A(n130), .B(n4749), .Z(n4748) );
  XOR U4402 ( .A(p_input[4]), .B(n4747), .Z(n4749) );
  XNOR U4403 ( .A(n4750), .B(n4751), .Z(n4747) );
  AND U4404 ( .A(n134), .B(n4752), .Z(n4751) );
  XOR U4405 ( .A(n4753), .B(n4754), .Z(n4745) );
  AND U4406 ( .A(n138), .B(n4755), .Z(n4754) );
  XOR U4407 ( .A(n4756), .B(n4757), .Z(n104) );
  AND U4408 ( .A(n142), .B(n4755), .Z(n4757) );
  XNOR U4409 ( .A(n4758), .B(n4756), .Z(n4755) );
  IV U4410 ( .A(n4753), .Z(n4758) );
  XOR U4411 ( .A(n4759), .B(n4760), .Z(n4753) );
  AND U4412 ( .A(n146), .B(n4752), .Z(n4760) );
  XNOR U4413 ( .A(n4750), .B(n4759), .Z(n4752) );
  XNOR U4414 ( .A(n4761), .B(n4762), .Z(n4750) );
  AND U4415 ( .A(n150), .B(n4763), .Z(n4762) );
  XOR U4416 ( .A(p_input[36]), .B(n4761), .Z(n4763) );
  XNOR U4417 ( .A(n4764), .B(n4765), .Z(n4761) );
  AND U4418 ( .A(n154), .B(n4766), .Z(n4765) );
  XOR U4419 ( .A(n4767), .B(n4768), .Z(n4759) );
  AND U4420 ( .A(n158), .B(n4769), .Z(n4768) );
  XOR U4421 ( .A(n4770), .B(n4771), .Z(n4756) );
  AND U4422 ( .A(n162), .B(n4769), .Z(n4771) );
  XNOR U4423 ( .A(n4772), .B(n4770), .Z(n4769) );
  IV U4424 ( .A(n4767), .Z(n4772) );
  XOR U4425 ( .A(n4773), .B(n4774), .Z(n4767) );
  AND U4426 ( .A(n165), .B(n4766), .Z(n4774) );
  XNOR U4427 ( .A(n4764), .B(n4773), .Z(n4766) );
  XNOR U4428 ( .A(n4775), .B(n4776), .Z(n4764) );
  AND U4429 ( .A(n169), .B(n4777), .Z(n4776) );
  XOR U4430 ( .A(p_input[68]), .B(n4775), .Z(n4777) );
  XNOR U4431 ( .A(n4778), .B(n4779), .Z(n4775) );
  AND U4432 ( .A(n173), .B(n4780), .Z(n4779) );
  XOR U4433 ( .A(n4781), .B(n4782), .Z(n4773) );
  AND U4434 ( .A(n177), .B(n4783), .Z(n4782) );
  XOR U4435 ( .A(n4784), .B(n4785), .Z(n4770) );
  AND U4436 ( .A(n181), .B(n4783), .Z(n4785) );
  XNOR U4437 ( .A(n4786), .B(n4784), .Z(n4783) );
  IV U4438 ( .A(n4781), .Z(n4786) );
  XOR U4439 ( .A(n4787), .B(n4788), .Z(n4781) );
  AND U4440 ( .A(n184), .B(n4780), .Z(n4788) );
  XNOR U4441 ( .A(n4778), .B(n4787), .Z(n4780) );
  XNOR U4442 ( .A(n4789), .B(n4790), .Z(n4778) );
  AND U4443 ( .A(n188), .B(n4791), .Z(n4790) );
  XOR U4444 ( .A(p_input[100]), .B(n4789), .Z(n4791) );
  XNOR U4445 ( .A(n4792), .B(n4793), .Z(n4789) );
  AND U4446 ( .A(n192), .B(n4794), .Z(n4793) );
  XOR U4447 ( .A(n4795), .B(n4796), .Z(n4787) );
  AND U4448 ( .A(n196), .B(n4797), .Z(n4796) );
  XOR U4449 ( .A(n4798), .B(n4799), .Z(n4784) );
  AND U4450 ( .A(n200), .B(n4797), .Z(n4799) );
  XNOR U4451 ( .A(n4800), .B(n4798), .Z(n4797) );
  IV U4452 ( .A(n4795), .Z(n4800) );
  XOR U4453 ( .A(n4801), .B(n4802), .Z(n4795) );
  AND U4454 ( .A(n203), .B(n4794), .Z(n4802) );
  XNOR U4455 ( .A(n4792), .B(n4801), .Z(n4794) );
  XNOR U4456 ( .A(n4803), .B(n4804), .Z(n4792) );
  AND U4457 ( .A(n207), .B(n4805), .Z(n4804) );
  XOR U4458 ( .A(p_input[132]), .B(n4803), .Z(n4805) );
  XNOR U4459 ( .A(n4806), .B(n4807), .Z(n4803) );
  AND U4460 ( .A(n211), .B(n4808), .Z(n4807) );
  XOR U4461 ( .A(n4809), .B(n4810), .Z(n4801) );
  AND U4462 ( .A(n215), .B(n4811), .Z(n4810) );
  XOR U4463 ( .A(n4812), .B(n4813), .Z(n4798) );
  AND U4464 ( .A(n219), .B(n4811), .Z(n4813) );
  XNOR U4465 ( .A(n4814), .B(n4812), .Z(n4811) );
  IV U4466 ( .A(n4809), .Z(n4814) );
  XOR U4467 ( .A(n4815), .B(n4816), .Z(n4809) );
  AND U4468 ( .A(n222), .B(n4808), .Z(n4816) );
  XNOR U4469 ( .A(n4806), .B(n4815), .Z(n4808) );
  XNOR U4470 ( .A(n4817), .B(n4818), .Z(n4806) );
  AND U4471 ( .A(n226), .B(n4819), .Z(n4818) );
  XOR U4472 ( .A(p_input[164]), .B(n4817), .Z(n4819) );
  XNOR U4473 ( .A(n4820), .B(n4821), .Z(n4817) );
  AND U4474 ( .A(n230), .B(n4822), .Z(n4821) );
  XOR U4475 ( .A(n4823), .B(n4824), .Z(n4815) );
  AND U4476 ( .A(n234), .B(n4825), .Z(n4824) );
  XOR U4477 ( .A(n4826), .B(n4827), .Z(n4812) );
  AND U4478 ( .A(n238), .B(n4825), .Z(n4827) );
  XNOR U4479 ( .A(n4828), .B(n4826), .Z(n4825) );
  IV U4480 ( .A(n4823), .Z(n4828) );
  XOR U4481 ( .A(n4829), .B(n4830), .Z(n4823) );
  AND U4482 ( .A(n241), .B(n4822), .Z(n4830) );
  XNOR U4483 ( .A(n4820), .B(n4829), .Z(n4822) );
  XNOR U4484 ( .A(n4831), .B(n4832), .Z(n4820) );
  AND U4485 ( .A(n245), .B(n4833), .Z(n4832) );
  XOR U4486 ( .A(p_input[196]), .B(n4831), .Z(n4833) );
  XNOR U4487 ( .A(n4834), .B(n4835), .Z(n4831) );
  AND U4488 ( .A(n249), .B(n4836), .Z(n4835) );
  XOR U4489 ( .A(n4837), .B(n4838), .Z(n4829) );
  AND U4490 ( .A(n253), .B(n4839), .Z(n4838) );
  XOR U4491 ( .A(n4840), .B(n4841), .Z(n4826) );
  AND U4492 ( .A(n257), .B(n4839), .Z(n4841) );
  XNOR U4493 ( .A(n4842), .B(n4840), .Z(n4839) );
  IV U4494 ( .A(n4837), .Z(n4842) );
  XOR U4495 ( .A(n4843), .B(n4844), .Z(n4837) );
  AND U4496 ( .A(n260), .B(n4836), .Z(n4844) );
  XNOR U4497 ( .A(n4834), .B(n4843), .Z(n4836) );
  XNOR U4498 ( .A(n4845), .B(n4846), .Z(n4834) );
  AND U4499 ( .A(n264), .B(n4847), .Z(n4846) );
  XOR U4500 ( .A(p_input[228]), .B(n4845), .Z(n4847) );
  XNOR U4501 ( .A(n4848), .B(n4849), .Z(n4845) );
  AND U4502 ( .A(n268), .B(n4850), .Z(n4849) );
  XOR U4503 ( .A(n4851), .B(n4852), .Z(n4843) );
  AND U4504 ( .A(n272), .B(n4853), .Z(n4852) );
  XOR U4505 ( .A(n4854), .B(n4855), .Z(n4840) );
  AND U4506 ( .A(n276), .B(n4853), .Z(n4855) );
  XNOR U4507 ( .A(n4856), .B(n4854), .Z(n4853) );
  IV U4508 ( .A(n4851), .Z(n4856) );
  XOR U4509 ( .A(n4857), .B(n4858), .Z(n4851) );
  AND U4510 ( .A(n279), .B(n4850), .Z(n4858) );
  XNOR U4511 ( .A(n4848), .B(n4857), .Z(n4850) );
  XNOR U4512 ( .A(n4859), .B(n4860), .Z(n4848) );
  AND U4513 ( .A(n283), .B(n4861), .Z(n4860) );
  XOR U4514 ( .A(p_input[260]), .B(n4859), .Z(n4861) );
  XNOR U4515 ( .A(n4862), .B(n4863), .Z(n4859) );
  AND U4516 ( .A(n287), .B(n4864), .Z(n4863) );
  XOR U4517 ( .A(n4865), .B(n4866), .Z(n4857) );
  AND U4518 ( .A(n291), .B(n4867), .Z(n4866) );
  XOR U4519 ( .A(n4868), .B(n4869), .Z(n4854) );
  AND U4520 ( .A(n295), .B(n4867), .Z(n4869) );
  XNOR U4521 ( .A(n4870), .B(n4868), .Z(n4867) );
  IV U4522 ( .A(n4865), .Z(n4870) );
  XOR U4523 ( .A(n4871), .B(n4872), .Z(n4865) );
  AND U4524 ( .A(n298), .B(n4864), .Z(n4872) );
  XNOR U4525 ( .A(n4862), .B(n4871), .Z(n4864) );
  XNOR U4526 ( .A(n4873), .B(n4874), .Z(n4862) );
  AND U4527 ( .A(n302), .B(n4875), .Z(n4874) );
  XOR U4528 ( .A(p_input[292]), .B(n4873), .Z(n4875) );
  XNOR U4529 ( .A(n4876), .B(n4877), .Z(n4873) );
  AND U4530 ( .A(n306), .B(n4878), .Z(n4877) );
  XOR U4531 ( .A(n4879), .B(n4880), .Z(n4871) );
  AND U4532 ( .A(n310), .B(n4881), .Z(n4880) );
  XOR U4533 ( .A(n4882), .B(n4883), .Z(n4868) );
  AND U4534 ( .A(n314), .B(n4881), .Z(n4883) );
  XNOR U4535 ( .A(n4884), .B(n4882), .Z(n4881) );
  IV U4536 ( .A(n4879), .Z(n4884) );
  XOR U4537 ( .A(n4885), .B(n4886), .Z(n4879) );
  AND U4538 ( .A(n317), .B(n4878), .Z(n4886) );
  XNOR U4539 ( .A(n4876), .B(n4885), .Z(n4878) );
  XNOR U4540 ( .A(n4887), .B(n4888), .Z(n4876) );
  AND U4541 ( .A(n321), .B(n4889), .Z(n4888) );
  XOR U4542 ( .A(p_input[324]), .B(n4887), .Z(n4889) );
  XNOR U4543 ( .A(n4890), .B(n4891), .Z(n4887) );
  AND U4544 ( .A(n325), .B(n4892), .Z(n4891) );
  XOR U4545 ( .A(n4893), .B(n4894), .Z(n4885) );
  AND U4546 ( .A(n329), .B(n4895), .Z(n4894) );
  XOR U4547 ( .A(n4896), .B(n4897), .Z(n4882) );
  AND U4548 ( .A(n333), .B(n4895), .Z(n4897) );
  XNOR U4549 ( .A(n4898), .B(n4896), .Z(n4895) );
  IV U4550 ( .A(n4893), .Z(n4898) );
  XOR U4551 ( .A(n4899), .B(n4900), .Z(n4893) );
  AND U4552 ( .A(n336), .B(n4892), .Z(n4900) );
  XNOR U4553 ( .A(n4890), .B(n4899), .Z(n4892) );
  XNOR U4554 ( .A(n4901), .B(n4902), .Z(n4890) );
  AND U4555 ( .A(n340), .B(n4903), .Z(n4902) );
  XOR U4556 ( .A(p_input[356]), .B(n4901), .Z(n4903) );
  XNOR U4557 ( .A(n4904), .B(n4905), .Z(n4901) );
  AND U4558 ( .A(n344), .B(n4906), .Z(n4905) );
  XOR U4559 ( .A(n4907), .B(n4908), .Z(n4899) );
  AND U4560 ( .A(n348), .B(n4909), .Z(n4908) );
  XOR U4561 ( .A(n4910), .B(n4911), .Z(n4896) );
  AND U4562 ( .A(n352), .B(n4909), .Z(n4911) );
  XNOR U4563 ( .A(n4912), .B(n4910), .Z(n4909) );
  IV U4564 ( .A(n4907), .Z(n4912) );
  XOR U4565 ( .A(n4913), .B(n4914), .Z(n4907) );
  AND U4566 ( .A(n355), .B(n4906), .Z(n4914) );
  XNOR U4567 ( .A(n4904), .B(n4913), .Z(n4906) );
  XNOR U4568 ( .A(n4915), .B(n4916), .Z(n4904) );
  AND U4569 ( .A(n359), .B(n4917), .Z(n4916) );
  XOR U4570 ( .A(p_input[388]), .B(n4915), .Z(n4917) );
  XNOR U4571 ( .A(n4918), .B(n4919), .Z(n4915) );
  AND U4572 ( .A(n363), .B(n4920), .Z(n4919) );
  XOR U4573 ( .A(n4921), .B(n4922), .Z(n4913) );
  AND U4574 ( .A(n367), .B(n4923), .Z(n4922) );
  XOR U4575 ( .A(n4924), .B(n4925), .Z(n4910) );
  AND U4576 ( .A(n371), .B(n4923), .Z(n4925) );
  XNOR U4577 ( .A(n4926), .B(n4924), .Z(n4923) );
  IV U4578 ( .A(n4921), .Z(n4926) );
  XOR U4579 ( .A(n4927), .B(n4928), .Z(n4921) );
  AND U4580 ( .A(n374), .B(n4920), .Z(n4928) );
  XNOR U4581 ( .A(n4918), .B(n4927), .Z(n4920) );
  XNOR U4582 ( .A(n4929), .B(n4930), .Z(n4918) );
  AND U4583 ( .A(n378), .B(n4931), .Z(n4930) );
  XOR U4584 ( .A(p_input[420]), .B(n4929), .Z(n4931) );
  XNOR U4585 ( .A(n4932), .B(n4933), .Z(n4929) );
  AND U4586 ( .A(n382), .B(n4934), .Z(n4933) );
  XOR U4587 ( .A(n4935), .B(n4936), .Z(n4927) );
  AND U4588 ( .A(n386), .B(n4937), .Z(n4936) );
  XOR U4589 ( .A(n4938), .B(n4939), .Z(n4924) );
  AND U4590 ( .A(n390), .B(n4937), .Z(n4939) );
  XNOR U4591 ( .A(n4940), .B(n4938), .Z(n4937) );
  IV U4592 ( .A(n4935), .Z(n4940) );
  XOR U4593 ( .A(n4941), .B(n4942), .Z(n4935) );
  AND U4594 ( .A(n393), .B(n4934), .Z(n4942) );
  XNOR U4595 ( .A(n4932), .B(n4941), .Z(n4934) );
  XNOR U4596 ( .A(n4943), .B(n4944), .Z(n4932) );
  AND U4597 ( .A(n397), .B(n4945), .Z(n4944) );
  XOR U4598 ( .A(p_input[452]), .B(n4943), .Z(n4945) );
  XNOR U4599 ( .A(n4946), .B(n4947), .Z(n4943) );
  AND U4600 ( .A(n401), .B(n4948), .Z(n4947) );
  XOR U4601 ( .A(n4949), .B(n4950), .Z(n4941) );
  AND U4602 ( .A(n405), .B(n4951), .Z(n4950) );
  XOR U4603 ( .A(n4952), .B(n4953), .Z(n4938) );
  AND U4604 ( .A(n409), .B(n4951), .Z(n4953) );
  XNOR U4605 ( .A(n4954), .B(n4952), .Z(n4951) );
  IV U4606 ( .A(n4949), .Z(n4954) );
  XOR U4607 ( .A(n4955), .B(n4956), .Z(n4949) );
  AND U4608 ( .A(n412), .B(n4948), .Z(n4956) );
  XNOR U4609 ( .A(n4946), .B(n4955), .Z(n4948) );
  XNOR U4610 ( .A(n4957), .B(n4958), .Z(n4946) );
  AND U4611 ( .A(n416), .B(n4959), .Z(n4958) );
  XOR U4612 ( .A(p_input[484]), .B(n4957), .Z(n4959) );
  XNOR U4613 ( .A(n4960), .B(n4961), .Z(n4957) );
  AND U4614 ( .A(n420), .B(n4962), .Z(n4961) );
  XOR U4615 ( .A(n4963), .B(n4964), .Z(n4955) );
  AND U4616 ( .A(n424), .B(n4965), .Z(n4964) );
  XOR U4617 ( .A(n4966), .B(n4967), .Z(n4952) );
  AND U4618 ( .A(n428), .B(n4965), .Z(n4967) );
  XNOR U4619 ( .A(n4968), .B(n4966), .Z(n4965) );
  IV U4620 ( .A(n4963), .Z(n4968) );
  XOR U4621 ( .A(n4969), .B(n4970), .Z(n4963) );
  AND U4622 ( .A(n431), .B(n4962), .Z(n4970) );
  XNOR U4623 ( .A(n4960), .B(n4969), .Z(n4962) );
  XNOR U4624 ( .A(n4971), .B(n4972), .Z(n4960) );
  AND U4625 ( .A(n435), .B(n4973), .Z(n4972) );
  XOR U4626 ( .A(p_input[516]), .B(n4971), .Z(n4973) );
  XNOR U4627 ( .A(n4974), .B(n4975), .Z(n4971) );
  AND U4628 ( .A(n439), .B(n4976), .Z(n4975) );
  XOR U4629 ( .A(n4977), .B(n4978), .Z(n4969) );
  AND U4630 ( .A(n443), .B(n4979), .Z(n4978) );
  XOR U4631 ( .A(n4980), .B(n4981), .Z(n4966) );
  AND U4632 ( .A(n447), .B(n4979), .Z(n4981) );
  XNOR U4633 ( .A(n4982), .B(n4980), .Z(n4979) );
  IV U4634 ( .A(n4977), .Z(n4982) );
  XOR U4635 ( .A(n4983), .B(n4984), .Z(n4977) );
  AND U4636 ( .A(n450), .B(n4976), .Z(n4984) );
  XNOR U4637 ( .A(n4974), .B(n4983), .Z(n4976) );
  XNOR U4638 ( .A(n4985), .B(n4986), .Z(n4974) );
  AND U4639 ( .A(n454), .B(n4987), .Z(n4986) );
  XOR U4640 ( .A(p_input[548]), .B(n4985), .Z(n4987) );
  XNOR U4641 ( .A(n4988), .B(n4989), .Z(n4985) );
  AND U4642 ( .A(n458), .B(n4990), .Z(n4989) );
  XOR U4643 ( .A(n4991), .B(n4992), .Z(n4983) );
  AND U4644 ( .A(n462), .B(n4993), .Z(n4992) );
  XOR U4645 ( .A(n4994), .B(n4995), .Z(n4980) );
  AND U4646 ( .A(n466), .B(n4993), .Z(n4995) );
  XNOR U4647 ( .A(n4996), .B(n4994), .Z(n4993) );
  IV U4648 ( .A(n4991), .Z(n4996) );
  XOR U4649 ( .A(n4997), .B(n4998), .Z(n4991) );
  AND U4650 ( .A(n469), .B(n4990), .Z(n4998) );
  XNOR U4651 ( .A(n4988), .B(n4997), .Z(n4990) );
  XNOR U4652 ( .A(n4999), .B(n5000), .Z(n4988) );
  AND U4653 ( .A(n473), .B(n5001), .Z(n5000) );
  XOR U4654 ( .A(p_input[580]), .B(n4999), .Z(n5001) );
  XNOR U4655 ( .A(n5002), .B(n5003), .Z(n4999) );
  AND U4656 ( .A(n477), .B(n5004), .Z(n5003) );
  XOR U4657 ( .A(n5005), .B(n5006), .Z(n4997) );
  AND U4658 ( .A(n481), .B(n5007), .Z(n5006) );
  XOR U4659 ( .A(n5008), .B(n5009), .Z(n4994) );
  AND U4660 ( .A(n485), .B(n5007), .Z(n5009) );
  XNOR U4661 ( .A(n5010), .B(n5008), .Z(n5007) );
  IV U4662 ( .A(n5005), .Z(n5010) );
  XOR U4663 ( .A(n5011), .B(n5012), .Z(n5005) );
  AND U4664 ( .A(n488), .B(n5004), .Z(n5012) );
  XNOR U4665 ( .A(n5002), .B(n5011), .Z(n5004) );
  XNOR U4666 ( .A(n5013), .B(n5014), .Z(n5002) );
  AND U4667 ( .A(n492), .B(n5015), .Z(n5014) );
  XOR U4668 ( .A(p_input[612]), .B(n5013), .Z(n5015) );
  XNOR U4669 ( .A(n5016), .B(n5017), .Z(n5013) );
  AND U4670 ( .A(n496), .B(n5018), .Z(n5017) );
  XOR U4671 ( .A(n5019), .B(n5020), .Z(n5011) );
  AND U4672 ( .A(n500), .B(n5021), .Z(n5020) );
  XOR U4673 ( .A(n5022), .B(n5023), .Z(n5008) );
  AND U4674 ( .A(n504), .B(n5021), .Z(n5023) );
  XNOR U4675 ( .A(n5024), .B(n5022), .Z(n5021) );
  IV U4676 ( .A(n5019), .Z(n5024) );
  XOR U4677 ( .A(n5025), .B(n5026), .Z(n5019) );
  AND U4678 ( .A(n507), .B(n5018), .Z(n5026) );
  XNOR U4679 ( .A(n5016), .B(n5025), .Z(n5018) );
  XNOR U4680 ( .A(n5027), .B(n5028), .Z(n5016) );
  AND U4681 ( .A(n511), .B(n5029), .Z(n5028) );
  XOR U4682 ( .A(p_input[644]), .B(n5027), .Z(n5029) );
  XNOR U4683 ( .A(n5030), .B(n5031), .Z(n5027) );
  AND U4684 ( .A(n515), .B(n5032), .Z(n5031) );
  XOR U4685 ( .A(n5033), .B(n5034), .Z(n5025) );
  AND U4686 ( .A(n519), .B(n5035), .Z(n5034) );
  XOR U4687 ( .A(n5036), .B(n5037), .Z(n5022) );
  AND U4688 ( .A(n523), .B(n5035), .Z(n5037) );
  XNOR U4689 ( .A(n5038), .B(n5036), .Z(n5035) );
  IV U4690 ( .A(n5033), .Z(n5038) );
  XOR U4691 ( .A(n5039), .B(n5040), .Z(n5033) );
  AND U4692 ( .A(n526), .B(n5032), .Z(n5040) );
  XNOR U4693 ( .A(n5030), .B(n5039), .Z(n5032) );
  XNOR U4694 ( .A(n5041), .B(n5042), .Z(n5030) );
  AND U4695 ( .A(n530), .B(n5043), .Z(n5042) );
  XOR U4696 ( .A(p_input[676]), .B(n5041), .Z(n5043) );
  XNOR U4697 ( .A(n5044), .B(n5045), .Z(n5041) );
  AND U4698 ( .A(n534), .B(n5046), .Z(n5045) );
  XOR U4699 ( .A(n5047), .B(n5048), .Z(n5039) );
  AND U4700 ( .A(n538), .B(n5049), .Z(n5048) );
  XOR U4701 ( .A(n5050), .B(n5051), .Z(n5036) );
  AND U4702 ( .A(n542), .B(n5049), .Z(n5051) );
  XNOR U4703 ( .A(n5052), .B(n5050), .Z(n5049) );
  IV U4704 ( .A(n5047), .Z(n5052) );
  XOR U4705 ( .A(n5053), .B(n5054), .Z(n5047) );
  AND U4706 ( .A(n545), .B(n5046), .Z(n5054) );
  XNOR U4707 ( .A(n5044), .B(n5053), .Z(n5046) );
  XNOR U4708 ( .A(n5055), .B(n5056), .Z(n5044) );
  AND U4709 ( .A(n549), .B(n5057), .Z(n5056) );
  XOR U4710 ( .A(p_input[708]), .B(n5055), .Z(n5057) );
  XNOR U4711 ( .A(n5058), .B(n5059), .Z(n5055) );
  AND U4712 ( .A(n553), .B(n5060), .Z(n5059) );
  XOR U4713 ( .A(n5061), .B(n5062), .Z(n5053) );
  AND U4714 ( .A(n557), .B(n5063), .Z(n5062) );
  XOR U4715 ( .A(n5064), .B(n5065), .Z(n5050) );
  AND U4716 ( .A(n561), .B(n5063), .Z(n5065) );
  XNOR U4717 ( .A(n5066), .B(n5064), .Z(n5063) );
  IV U4718 ( .A(n5061), .Z(n5066) );
  XOR U4719 ( .A(n5067), .B(n5068), .Z(n5061) );
  AND U4720 ( .A(n564), .B(n5060), .Z(n5068) );
  XNOR U4721 ( .A(n5058), .B(n5067), .Z(n5060) );
  XNOR U4722 ( .A(n5069), .B(n5070), .Z(n5058) );
  AND U4723 ( .A(n568), .B(n5071), .Z(n5070) );
  XOR U4724 ( .A(p_input[740]), .B(n5069), .Z(n5071) );
  XNOR U4725 ( .A(n5072), .B(n5073), .Z(n5069) );
  AND U4726 ( .A(n572), .B(n5074), .Z(n5073) );
  XOR U4727 ( .A(n5075), .B(n5076), .Z(n5067) );
  AND U4728 ( .A(n576), .B(n5077), .Z(n5076) );
  XOR U4729 ( .A(n5078), .B(n5079), .Z(n5064) );
  AND U4730 ( .A(n580), .B(n5077), .Z(n5079) );
  XNOR U4731 ( .A(n5080), .B(n5078), .Z(n5077) );
  IV U4732 ( .A(n5075), .Z(n5080) );
  XOR U4733 ( .A(n5081), .B(n5082), .Z(n5075) );
  AND U4734 ( .A(n583), .B(n5074), .Z(n5082) );
  XNOR U4735 ( .A(n5072), .B(n5081), .Z(n5074) );
  XNOR U4736 ( .A(n5083), .B(n5084), .Z(n5072) );
  AND U4737 ( .A(n587), .B(n5085), .Z(n5084) );
  XOR U4738 ( .A(p_input[772]), .B(n5083), .Z(n5085) );
  XNOR U4739 ( .A(n5086), .B(n5087), .Z(n5083) );
  AND U4740 ( .A(n591), .B(n5088), .Z(n5087) );
  XOR U4741 ( .A(n5089), .B(n5090), .Z(n5081) );
  AND U4742 ( .A(n595), .B(n5091), .Z(n5090) );
  XOR U4743 ( .A(n5092), .B(n5093), .Z(n5078) );
  AND U4744 ( .A(n599), .B(n5091), .Z(n5093) );
  XNOR U4745 ( .A(n5094), .B(n5092), .Z(n5091) );
  IV U4746 ( .A(n5089), .Z(n5094) );
  XOR U4747 ( .A(n5095), .B(n5096), .Z(n5089) );
  AND U4748 ( .A(n602), .B(n5088), .Z(n5096) );
  XNOR U4749 ( .A(n5086), .B(n5095), .Z(n5088) );
  XNOR U4750 ( .A(n5097), .B(n5098), .Z(n5086) );
  AND U4751 ( .A(n606), .B(n5099), .Z(n5098) );
  XOR U4752 ( .A(p_input[804]), .B(n5097), .Z(n5099) );
  XNOR U4753 ( .A(n5100), .B(n5101), .Z(n5097) );
  AND U4754 ( .A(n610), .B(n5102), .Z(n5101) );
  XOR U4755 ( .A(n5103), .B(n5104), .Z(n5095) );
  AND U4756 ( .A(n614), .B(n5105), .Z(n5104) );
  XOR U4757 ( .A(n5106), .B(n5107), .Z(n5092) );
  AND U4758 ( .A(n618), .B(n5105), .Z(n5107) );
  XNOR U4759 ( .A(n5108), .B(n5106), .Z(n5105) );
  IV U4760 ( .A(n5103), .Z(n5108) );
  XOR U4761 ( .A(n5109), .B(n5110), .Z(n5103) );
  AND U4762 ( .A(n621), .B(n5102), .Z(n5110) );
  XNOR U4763 ( .A(n5100), .B(n5109), .Z(n5102) );
  XNOR U4764 ( .A(n5111), .B(n5112), .Z(n5100) );
  AND U4765 ( .A(n625), .B(n5113), .Z(n5112) );
  XOR U4766 ( .A(p_input[836]), .B(n5111), .Z(n5113) );
  XNOR U4767 ( .A(n5114), .B(n5115), .Z(n5111) );
  AND U4768 ( .A(n629), .B(n5116), .Z(n5115) );
  XOR U4769 ( .A(n5117), .B(n5118), .Z(n5109) );
  AND U4770 ( .A(n633), .B(n5119), .Z(n5118) );
  XOR U4771 ( .A(n5120), .B(n5121), .Z(n5106) );
  AND U4772 ( .A(n637), .B(n5119), .Z(n5121) );
  XNOR U4773 ( .A(n5122), .B(n5120), .Z(n5119) );
  IV U4774 ( .A(n5117), .Z(n5122) );
  XOR U4775 ( .A(n5123), .B(n5124), .Z(n5117) );
  AND U4776 ( .A(n640), .B(n5116), .Z(n5124) );
  XNOR U4777 ( .A(n5114), .B(n5123), .Z(n5116) );
  XNOR U4778 ( .A(n5125), .B(n5126), .Z(n5114) );
  AND U4779 ( .A(n644), .B(n5127), .Z(n5126) );
  XOR U4780 ( .A(p_input[868]), .B(n5125), .Z(n5127) );
  XNOR U4781 ( .A(n5128), .B(n5129), .Z(n5125) );
  AND U4782 ( .A(n648), .B(n5130), .Z(n5129) );
  XOR U4783 ( .A(n5131), .B(n5132), .Z(n5123) );
  AND U4784 ( .A(n652), .B(n5133), .Z(n5132) );
  XOR U4785 ( .A(n5134), .B(n5135), .Z(n5120) );
  AND U4786 ( .A(n656), .B(n5133), .Z(n5135) );
  XNOR U4787 ( .A(n5136), .B(n5134), .Z(n5133) );
  IV U4788 ( .A(n5131), .Z(n5136) );
  XOR U4789 ( .A(n5137), .B(n5138), .Z(n5131) );
  AND U4790 ( .A(n659), .B(n5130), .Z(n5138) );
  XNOR U4791 ( .A(n5128), .B(n5137), .Z(n5130) );
  XNOR U4792 ( .A(n5139), .B(n5140), .Z(n5128) );
  AND U4793 ( .A(n663), .B(n5141), .Z(n5140) );
  XOR U4794 ( .A(p_input[900]), .B(n5139), .Z(n5141) );
  XNOR U4795 ( .A(n5142), .B(n5143), .Z(n5139) );
  AND U4796 ( .A(n667), .B(n5144), .Z(n5143) );
  XOR U4797 ( .A(n5145), .B(n5146), .Z(n5137) );
  AND U4798 ( .A(n671), .B(n5147), .Z(n5146) );
  XOR U4799 ( .A(n5148), .B(n5149), .Z(n5134) );
  AND U4800 ( .A(n675), .B(n5147), .Z(n5149) );
  XNOR U4801 ( .A(n5150), .B(n5148), .Z(n5147) );
  IV U4802 ( .A(n5145), .Z(n5150) );
  XOR U4803 ( .A(n5151), .B(n5152), .Z(n5145) );
  AND U4804 ( .A(n678), .B(n5144), .Z(n5152) );
  XNOR U4805 ( .A(n5142), .B(n5151), .Z(n5144) );
  XNOR U4806 ( .A(n5153), .B(n5154), .Z(n5142) );
  AND U4807 ( .A(n682), .B(n5155), .Z(n5154) );
  XOR U4808 ( .A(p_input[932]), .B(n5153), .Z(n5155) );
  XNOR U4809 ( .A(n5156), .B(n5157), .Z(n5153) );
  AND U4810 ( .A(n686), .B(n5158), .Z(n5157) );
  XOR U4811 ( .A(n5159), .B(n5160), .Z(n5151) );
  AND U4812 ( .A(n690), .B(n5161), .Z(n5160) );
  XOR U4813 ( .A(n5162), .B(n5163), .Z(n5148) );
  AND U4814 ( .A(n694), .B(n5161), .Z(n5163) );
  XNOR U4815 ( .A(n5164), .B(n5162), .Z(n5161) );
  IV U4816 ( .A(n5159), .Z(n5164) );
  XOR U4817 ( .A(n5165), .B(n5166), .Z(n5159) );
  AND U4818 ( .A(n697), .B(n5158), .Z(n5166) );
  XNOR U4819 ( .A(n5156), .B(n5165), .Z(n5158) );
  XNOR U4820 ( .A(n5167), .B(n5168), .Z(n5156) );
  AND U4821 ( .A(n701), .B(n5169), .Z(n5168) );
  XOR U4822 ( .A(p_input[964]), .B(n5167), .Z(n5169) );
  XNOR U4823 ( .A(n5170), .B(n5171), .Z(n5167) );
  AND U4824 ( .A(n705), .B(n5172), .Z(n5171) );
  XOR U4825 ( .A(n5173), .B(n5174), .Z(n5165) );
  AND U4826 ( .A(n709), .B(n5175), .Z(n5174) );
  XOR U4827 ( .A(n5176), .B(n5177), .Z(n5162) );
  AND U4828 ( .A(n713), .B(n5175), .Z(n5177) );
  XNOR U4829 ( .A(n5178), .B(n5176), .Z(n5175) );
  IV U4830 ( .A(n5173), .Z(n5178) );
  XOR U4831 ( .A(n5179), .B(n5180), .Z(n5173) );
  AND U4832 ( .A(n716), .B(n5172), .Z(n5180) );
  XNOR U4833 ( .A(n5170), .B(n5179), .Z(n5172) );
  XNOR U4834 ( .A(n5181), .B(n5182), .Z(n5170) );
  AND U4835 ( .A(n720), .B(n5183), .Z(n5182) );
  XOR U4836 ( .A(p_input[996]), .B(n5181), .Z(n5183) );
  XNOR U4837 ( .A(n5184), .B(n5185), .Z(n5181) );
  AND U4838 ( .A(n724), .B(n5186), .Z(n5185) );
  XOR U4839 ( .A(n5187), .B(n5188), .Z(n5179) );
  AND U4840 ( .A(n728), .B(n5189), .Z(n5188) );
  XOR U4841 ( .A(n5190), .B(n5191), .Z(n5176) );
  AND U4842 ( .A(n732), .B(n5189), .Z(n5191) );
  XNOR U4843 ( .A(n5192), .B(n5190), .Z(n5189) );
  IV U4844 ( .A(n5187), .Z(n5192) );
  XOR U4845 ( .A(n5193), .B(n5194), .Z(n5187) );
  AND U4846 ( .A(n735), .B(n5186), .Z(n5194) );
  XNOR U4847 ( .A(n5184), .B(n5193), .Z(n5186) );
  XNOR U4848 ( .A(n5195), .B(n5196), .Z(n5184) );
  AND U4849 ( .A(n739), .B(n5197), .Z(n5196) );
  XOR U4850 ( .A(p_input[1028]), .B(n5195), .Z(n5197) );
  XNOR U4851 ( .A(n5198), .B(n5199), .Z(n5195) );
  AND U4852 ( .A(n743), .B(n5200), .Z(n5199) );
  XOR U4853 ( .A(n5201), .B(n5202), .Z(n5193) );
  AND U4854 ( .A(n747), .B(n5203), .Z(n5202) );
  XOR U4855 ( .A(n5204), .B(n5205), .Z(n5190) );
  AND U4856 ( .A(n751), .B(n5203), .Z(n5205) );
  XNOR U4857 ( .A(n5206), .B(n5204), .Z(n5203) );
  IV U4858 ( .A(n5201), .Z(n5206) );
  XOR U4859 ( .A(n5207), .B(n5208), .Z(n5201) );
  AND U4860 ( .A(n754), .B(n5200), .Z(n5208) );
  XNOR U4861 ( .A(n5198), .B(n5207), .Z(n5200) );
  XNOR U4862 ( .A(n5209), .B(n5210), .Z(n5198) );
  AND U4863 ( .A(n758), .B(n5211), .Z(n5210) );
  XOR U4864 ( .A(p_input[1060]), .B(n5209), .Z(n5211) );
  XNOR U4865 ( .A(n5212), .B(n5213), .Z(n5209) );
  AND U4866 ( .A(n762), .B(n5214), .Z(n5213) );
  XOR U4867 ( .A(n5215), .B(n5216), .Z(n5207) );
  AND U4868 ( .A(n766), .B(n5217), .Z(n5216) );
  XOR U4869 ( .A(n5218), .B(n5219), .Z(n5204) );
  AND U4870 ( .A(n770), .B(n5217), .Z(n5219) );
  XNOR U4871 ( .A(n5220), .B(n5218), .Z(n5217) );
  IV U4872 ( .A(n5215), .Z(n5220) );
  XOR U4873 ( .A(n5221), .B(n5222), .Z(n5215) );
  AND U4874 ( .A(n773), .B(n5214), .Z(n5222) );
  XNOR U4875 ( .A(n5212), .B(n5221), .Z(n5214) );
  XNOR U4876 ( .A(n5223), .B(n5224), .Z(n5212) );
  AND U4877 ( .A(n777), .B(n5225), .Z(n5224) );
  XOR U4878 ( .A(p_input[1092]), .B(n5223), .Z(n5225) );
  XNOR U4879 ( .A(n5226), .B(n5227), .Z(n5223) );
  AND U4880 ( .A(n781), .B(n5228), .Z(n5227) );
  XOR U4881 ( .A(n5229), .B(n5230), .Z(n5221) );
  AND U4882 ( .A(n785), .B(n5231), .Z(n5230) );
  XOR U4883 ( .A(n5232), .B(n5233), .Z(n5218) );
  AND U4884 ( .A(n789), .B(n5231), .Z(n5233) );
  XNOR U4885 ( .A(n5234), .B(n5232), .Z(n5231) );
  IV U4886 ( .A(n5229), .Z(n5234) );
  XOR U4887 ( .A(n5235), .B(n5236), .Z(n5229) );
  AND U4888 ( .A(n792), .B(n5228), .Z(n5236) );
  XNOR U4889 ( .A(n5226), .B(n5235), .Z(n5228) );
  XNOR U4890 ( .A(n5237), .B(n5238), .Z(n5226) );
  AND U4891 ( .A(n796), .B(n5239), .Z(n5238) );
  XOR U4892 ( .A(p_input[1124]), .B(n5237), .Z(n5239) );
  XNOR U4893 ( .A(n5240), .B(n5241), .Z(n5237) );
  AND U4894 ( .A(n800), .B(n5242), .Z(n5241) );
  XOR U4895 ( .A(n5243), .B(n5244), .Z(n5235) );
  AND U4896 ( .A(n804), .B(n5245), .Z(n5244) );
  XOR U4897 ( .A(n5246), .B(n5247), .Z(n5232) );
  AND U4898 ( .A(n808), .B(n5245), .Z(n5247) );
  XNOR U4899 ( .A(n5248), .B(n5246), .Z(n5245) );
  IV U4900 ( .A(n5243), .Z(n5248) );
  XOR U4901 ( .A(n5249), .B(n5250), .Z(n5243) );
  AND U4902 ( .A(n811), .B(n5242), .Z(n5250) );
  XNOR U4903 ( .A(n5240), .B(n5249), .Z(n5242) );
  XNOR U4904 ( .A(n5251), .B(n5252), .Z(n5240) );
  AND U4905 ( .A(n815), .B(n5253), .Z(n5252) );
  XOR U4906 ( .A(p_input[1156]), .B(n5251), .Z(n5253) );
  XNOR U4907 ( .A(n5254), .B(n5255), .Z(n5251) );
  AND U4908 ( .A(n819), .B(n5256), .Z(n5255) );
  XOR U4909 ( .A(n5257), .B(n5258), .Z(n5249) );
  AND U4910 ( .A(n823), .B(n5259), .Z(n5258) );
  XOR U4911 ( .A(n5260), .B(n5261), .Z(n5246) );
  AND U4912 ( .A(n827), .B(n5259), .Z(n5261) );
  XNOR U4913 ( .A(n5262), .B(n5260), .Z(n5259) );
  IV U4914 ( .A(n5257), .Z(n5262) );
  XOR U4915 ( .A(n5263), .B(n5264), .Z(n5257) );
  AND U4916 ( .A(n830), .B(n5256), .Z(n5264) );
  XNOR U4917 ( .A(n5254), .B(n5263), .Z(n5256) );
  XNOR U4918 ( .A(n5265), .B(n5266), .Z(n5254) );
  AND U4919 ( .A(n834), .B(n5267), .Z(n5266) );
  XOR U4920 ( .A(p_input[1188]), .B(n5265), .Z(n5267) );
  XNOR U4921 ( .A(n5268), .B(n5269), .Z(n5265) );
  AND U4922 ( .A(n838), .B(n5270), .Z(n5269) );
  XOR U4923 ( .A(n5271), .B(n5272), .Z(n5263) );
  AND U4924 ( .A(n842), .B(n5273), .Z(n5272) );
  XOR U4925 ( .A(n5274), .B(n5275), .Z(n5260) );
  AND U4926 ( .A(n846), .B(n5273), .Z(n5275) );
  XNOR U4927 ( .A(n5276), .B(n5274), .Z(n5273) );
  IV U4928 ( .A(n5271), .Z(n5276) );
  XOR U4929 ( .A(n5277), .B(n5278), .Z(n5271) );
  AND U4930 ( .A(n849), .B(n5270), .Z(n5278) );
  XNOR U4931 ( .A(n5268), .B(n5277), .Z(n5270) );
  XNOR U4932 ( .A(n5279), .B(n5280), .Z(n5268) );
  AND U4933 ( .A(n853), .B(n5281), .Z(n5280) );
  XOR U4934 ( .A(p_input[1220]), .B(n5279), .Z(n5281) );
  XNOR U4935 ( .A(n5282), .B(n5283), .Z(n5279) );
  AND U4936 ( .A(n857), .B(n5284), .Z(n5283) );
  XOR U4937 ( .A(n5285), .B(n5286), .Z(n5277) );
  AND U4938 ( .A(n861), .B(n5287), .Z(n5286) );
  XOR U4939 ( .A(n5288), .B(n5289), .Z(n5274) );
  AND U4940 ( .A(n865), .B(n5287), .Z(n5289) );
  XNOR U4941 ( .A(n5290), .B(n5288), .Z(n5287) );
  IV U4942 ( .A(n5285), .Z(n5290) );
  XOR U4943 ( .A(n5291), .B(n5292), .Z(n5285) );
  AND U4944 ( .A(n868), .B(n5284), .Z(n5292) );
  XNOR U4945 ( .A(n5282), .B(n5291), .Z(n5284) );
  XNOR U4946 ( .A(n5293), .B(n5294), .Z(n5282) );
  AND U4947 ( .A(n872), .B(n5295), .Z(n5294) );
  XOR U4948 ( .A(p_input[1252]), .B(n5293), .Z(n5295) );
  XNOR U4949 ( .A(n5296), .B(n5297), .Z(n5293) );
  AND U4950 ( .A(n876), .B(n5298), .Z(n5297) );
  XOR U4951 ( .A(n5299), .B(n5300), .Z(n5291) );
  AND U4952 ( .A(n880), .B(n5301), .Z(n5300) );
  XOR U4953 ( .A(n5302), .B(n5303), .Z(n5288) );
  AND U4954 ( .A(n884), .B(n5301), .Z(n5303) );
  XNOR U4955 ( .A(n5304), .B(n5302), .Z(n5301) );
  IV U4956 ( .A(n5299), .Z(n5304) );
  XOR U4957 ( .A(n5305), .B(n5306), .Z(n5299) );
  AND U4958 ( .A(n887), .B(n5298), .Z(n5306) );
  XNOR U4959 ( .A(n5296), .B(n5305), .Z(n5298) );
  XNOR U4960 ( .A(n5307), .B(n5308), .Z(n5296) );
  AND U4961 ( .A(n891), .B(n5309), .Z(n5308) );
  XOR U4962 ( .A(p_input[1284]), .B(n5307), .Z(n5309) );
  XNOR U4963 ( .A(n5310), .B(n5311), .Z(n5307) );
  AND U4964 ( .A(n895), .B(n5312), .Z(n5311) );
  XOR U4965 ( .A(n5313), .B(n5314), .Z(n5305) );
  AND U4966 ( .A(n899), .B(n5315), .Z(n5314) );
  XOR U4967 ( .A(n5316), .B(n5317), .Z(n5302) );
  AND U4968 ( .A(n903), .B(n5315), .Z(n5317) );
  XNOR U4969 ( .A(n5318), .B(n5316), .Z(n5315) );
  IV U4970 ( .A(n5313), .Z(n5318) );
  XOR U4971 ( .A(n5319), .B(n5320), .Z(n5313) );
  AND U4972 ( .A(n906), .B(n5312), .Z(n5320) );
  XNOR U4973 ( .A(n5310), .B(n5319), .Z(n5312) );
  XNOR U4974 ( .A(n5321), .B(n5322), .Z(n5310) );
  AND U4975 ( .A(n910), .B(n5323), .Z(n5322) );
  XOR U4976 ( .A(p_input[1316]), .B(n5321), .Z(n5323) );
  XNOR U4977 ( .A(n5324), .B(n5325), .Z(n5321) );
  AND U4978 ( .A(n914), .B(n5326), .Z(n5325) );
  XOR U4979 ( .A(n5327), .B(n5328), .Z(n5319) );
  AND U4980 ( .A(n918), .B(n5329), .Z(n5328) );
  XOR U4981 ( .A(n5330), .B(n5331), .Z(n5316) );
  AND U4982 ( .A(n922), .B(n5329), .Z(n5331) );
  XNOR U4983 ( .A(n5332), .B(n5330), .Z(n5329) );
  IV U4984 ( .A(n5327), .Z(n5332) );
  XOR U4985 ( .A(n5333), .B(n5334), .Z(n5327) );
  AND U4986 ( .A(n925), .B(n5326), .Z(n5334) );
  XNOR U4987 ( .A(n5324), .B(n5333), .Z(n5326) );
  XNOR U4988 ( .A(n5335), .B(n5336), .Z(n5324) );
  AND U4989 ( .A(n929), .B(n5337), .Z(n5336) );
  XOR U4990 ( .A(p_input[1348]), .B(n5335), .Z(n5337) );
  XNOR U4991 ( .A(n5338), .B(n5339), .Z(n5335) );
  AND U4992 ( .A(n933), .B(n5340), .Z(n5339) );
  XOR U4993 ( .A(n5341), .B(n5342), .Z(n5333) );
  AND U4994 ( .A(n937), .B(n5343), .Z(n5342) );
  XOR U4995 ( .A(n5344), .B(n5345), .Z(n5330) );
  AND U4996 ( .A(n941), .B(n5343), .Z(n5345) );
  XNOR U4997 ( .A(n5346), .B(n5344), .Z(n5343) );
  IV U4998 ( .A(n5341), .Z(n5346) );
  XOR U4999 ( .A(n5347), .B(n5348), .Z(n5341) );
  AND U5000 ( .A(n944), .B(n5340), .Z(n5348) );
  XNOR U5001 ( .A(n5338), .B(n5347), .Z(n5340) );
  XNOR U5002 ( .A(n5349), .B(n5350), .Z(n5338) );
  AND U5003 ( .A(n948), .B(n5351), .Z(n5350) );
  XOR U5004 ( .A(p_input[1380]), .B(n5349), .Z(n5351) );
  XNOR U5005 ( .A(n5352), .B(n5353), .Z(n5349) );
  AND U5006 ( .A(n952), .B(n5354), .Z(n5353) );
  XOR U5007 ( .A(n5355), .B(n5356), .Z(n5347) );
  AND U5008 ( .A(n956), .B(n5357), .Z(n5356) );
  XOR U5009 ( .A(n5358), .B(n5359), .Z(n5344) );
  AND U5010 ( .A(n960), .B(n5357), .Z(n5359) );
  XNOR U5011 ( .A(n5360), .B(n5358), .Z(n5357) );
  IV U5012 ( .A(n5355), .Z(n5360) );
  XOR U5013 ( .A(n5361), .B(n5362), .Z(n5355) );
  AND U5014 ( .A(n963), .B(n5354), .Z(n5362) );
  XNOR U5015 ( .A(n5352), .B(n5361), .Z(n5354) );
  XNOR U5016 ( .A(n5363), .B(n5364), .Z(n5352) );
  AND U5017 ( .A(n967), .B(n5365), .Z(n5364) );
  XOR U5018 ( .A(p_input[1412]), .B(n5363), .Z(n5365) );
  XNOR U5019 ( .A(n5366), .B(n5367), .Z(n5363) );
  AND U5020 ( .A(n971), .B(n5368), .Z(n5367) );
  XOR U5021 ( .A(n5369), .B(n5370), .Z(n5361) );
  AND U5022 ( .A(n975), .B(n5371), .Z(n5370) );
  XOR U5023 ( .A(n5372), .B(n5373), .Z(n5358) );
  AND U5024 ( .A(n979), .B(n5371), .Z(n5373) );
  XNOR U5025 ( .A(n5374), .B(n5372), .Z(n5371) );
  IV U5026 ( .A(n5369), .Z(n5374) );
  XOR U5027 ( .A(n5375), .B(n5376), .Z(n5369) );
  AND U5028 ( .A(n982), .B(n5368), .Z(n5376) );
  XNOR U5029 ( .A(n5366), .B(n5375), .Z(n5368) );
  XNOR U5030 ( .A(n5377), .B(n5378), .Z(n5366) );
  AND U5031 ( .A(n986), .B(n5379), .Z(n5378) );
  XOR U5032 ( .A(p_input[1444]), .B(n5377), .Z(n5379) );
  XNOR U5033 ( .A(n5380), .B(n5381), .Z(n5377) );
  AND U5034 ( .A(n990), .B(n5382), .Z(n5381) );
  XOR U5035 ( .A(n5383), .B(n5384), .Z(n5375) );
  AND U5036 ( .A(n994), .B(n5385), .Z(n5384) );
  XOR U5037 ( .A(n5386), .B(n5387), .Z(n5372) );
  AND U5038 ( .A(n998), .B(n5385), .Z(n5387) );
  XNOR U5039 ( .A(n5388), .B(n5386), .Z(n5385) );
  IV U5040 ( .A(n5383), .Z(n5388) );
  XOR U5041 ( .A(n5389), .B(n5390), .Z(n5383) );
  AND U5042 ( .A(n1001), .B(n5382), .Z(n5390) );
  XNOR U5043 ( .A(n5380), .B(n5389), .Z(n5382) );
  XNOR U5044 ( .A(n5391), .B(n5392), .Z(n5380) );
  AND U5045 ( .A(n1005), .B(n5393), .Z(n5392) );
  XOR U5046 ( .A(p_input[1476]), .B(n5391), .Z(n5393) );
  XNOR U5047 ( .A(n5394), .B(n5395), .Z(n5391) );
  AND U5048 ( .A(n1009), .B(n5396), .Z(n5395) );
  XOR U5049 ( .A(n5397), .B(n5398), .Z(n5389) );
  AND U5050 ( .A(n1013), .B(n5399), .Z(n5398) );
  XOR U5051 ( .A(n5400), .B(n5401), .Z(n5386) );
  AND U5052 ( .A(n1017), .B(n5399), .Z(n5401) );
  XNOR U5053 ( .A(n5402), .B(n5400), .Z(n5399) );
  IV U5054 ( .A(n5397), .Z(n5402) );
  XOR U5055 ( .A(n5403), .B(n5404), .Z(n5397) );
  AND U5056 ( .A(n1020), .B(n5396), .Z(n5404) );
  XNOR U5057 ( .A(n5394), .B(n5403), .Z(n5396) );
  XNOR U5058 ( .A(n5405), .B(n5406), .Z(n5394) );
  AND U5059 ( .A(n1024), .B(n5407), .Z(n5406) );
  XOR U5060 ( .A(p_input[1508]), .B(n5405), .Z(n5407) );
  XNOR U5061 ( .A(n5408), .B(n5409), .Z(n5405) );
  AND U5062 ( .A(n1028), .B(n5410), .Z(n5409) );
  XOR U5063 ( .A(n5411), .B(n5412), .Z(n5403) );
  AND U5064 ( .A(n1032), .B(n5413), .Z(n5412) );
  XOR U5065 ( .A(n5414), .B(n5415), .Z(n5400) );
  AND U5066 ( .A(n1036), .B(n5413), .Z(n5415) );
  XNOR U5067 ( .A(n5416), .B(n5414), .Z(n5413) );
  IV U5068 ( .A(n5411), .Z(n5416) );
  XOR U5069 ( .A(n5417), .B(n5418), .Z(n5411) );
  AND U5070 ( .A(n1039), .B(n5410), .Z(n5418) );
  XNOR U5071 ( .A(n5408), .B(n5417), .Z(n5410) );
  XNOR U5072 ( .A(n5419), .B(n5420), .Z(n5408) );
  AND U5073 ( .A(n1043), .B(n5421), .Z(n5420) );
  XOR U5074 ( .A(p_input[1540]), .B(n5419), .Z(n5421) );
  XNOR U5075 ( .A(n5422), .B(n5423), .Z(n5419) );
  AND U5076 ( .A(n1047), .B(n5424), .Z(n5423) );
  XOR U5077 ( .A(n5425), .B(n5426), .Z(n5417) );
  AND U5078 ( .A(n1051), .B(n5427), .Z(n5426) );
  XOR U5079 ( .A(n5428), .B(n5429), .Z(n5414) );
  AND U5080 ( .A(n1055), .B(n5427), .Z(n5429) );
  XNOR U5081 ( .A(n5430), .B(n5428), .Z(n5427) );
  IV U5082 ( .A(n5425), .Z(n5430) );
  XOR U5083 ( .A(n5431), .B(n5432), .Z(n5425) );
  AND U5084 ( .A(n1058), .B(n5424), .Z(n5432) );
  XNOR U5085 ( .A(n5422), .B(n5431), .Z(n5424) );
  XNOR U5086 ( .A(n5433), .B(n5434), .Z(n5422) );
  AND U5087 ( .A(n1062), .B(n5435), .Z(n5434) );
  XOR U5088 ( .A(p_input[1572]), .B(n5433), .Z(n5435) );
  XNOR U5089 ( .A(n5436), .B(n5437), .Z(n5433) );
  AND U5090 ( .A(n1066), .B(n5438), .Z(n5437) );
  XOR U5091 ( .A(n5439), .B(n5440), .Z(n5431) );
  AND U5092 ( .A(n1070), .B(n5441), .Z(n5440) );
  XOR U5093 ( .A(n5442), .B(n5443), .Z(n5428) );
  AND U5094 ( .A(n1074), .B(n5441), .Z(n5443) );
  XNOR U5095 ( .A(n5444), .B(n5442), .Z(n5441) );
  IV U5096 ( .A(n5439), .Z(n5444) );
  XOR U5097 ( .A(n5445), .B(n5446), .Z(n5439) );
  AND U5098 ( .A(n1077), .B(n5438), .Z(n5446) );
  XNOR U5099 ( .A(n5436), .B(n5445), .Z(n5438) );
  XNOR U5100 ( .A(n5447), .B(n5448), .Z(n5436) );
  AND U5101 ( .A(n1081), .B(n5449), .Z(n5448) );
  XOR U5102 ( .A(p_input[1604]), .B(n5447), .Z(n5449) );
  XNOR U5103 ( .A(n5450), .B(n5451), .Z(n5447) );
  AND U5104 ( .A(n1085), .B(n5452), .Z(n5451) );
  XOR U5105 ( .A(n5453), .B(n5454), .Z(n5445) );
  AND U5106 ( .A(n1089), .B(n5455), .Z(n5454) );
  XOR U5107 ( .A(n5456), .B(n5457), .Z(n5442) );
  AND U5108 ( .A(n1093), .B(n5455), .Z(n5457) );
  XNOR U5109 ( .A(n5458), .B(n5456), .Z(n5455) );
  IV U5110 ( .A(n5453), .Z(n5458) );
  XOR U5111 ( .A(n5459), .B(n5460), .Z(n5453) );
  AND U5112 ( .A(n1096), .B(n5452), .Z(n5460) );
  XNOR U5113 ( .A(n5450), .B(n5459), .Z(n5452) );
  XNOR U5114 ( .A(n5461), .B(n5462), .Z(n5450) );
  AND U5115 ( .A(n1100), .B(n5463), .Z(n5462) );
  XOR U5116 ( .A(p_input[1636]), .B(n5461), .Z(n5463) );
  XNOR U5117 ( .A(n5464), .B(n5465), .Z(n5461) );
  AND U5118 ( .A(n1104), .B(n5466), .Z(n5465) );
  XOR U5119 ( .A(n5467), .B(n5468), .Z(n5459) );
  AND U5120 ( .A(n1108), .B(n5469), .Z(n5468) );
  XOR U5121 ( .A(n5470), .B(n5471), .Z(n5456) );
  AND U5122 ( .A(n1112), .B(n5469), .Z(n5471) );
  XNOR U5123 ( .A(n5472), .B(n5470), .Z(n5469) );
  IV U5124 ( .A(n5467), .Z(n5472) );
  XOR U5125 ( .A(n5473), .B(n5474), .Z(n5467) );
  AND U5126 ( .A(n1115), .B(n5466), .Z(n5474) );
  XNOR U5127 ( .A(n5464), .B(n5473), .Z(n5466) );
  XNOR U5128 ( .A(n5475), .B(n5476), .Z(n5464) );
  AND U5129 ( .A(n1119), .B(n5477), .Z(n5476) );
  XOR U5130 ( .A(p_input[1668]), .B(n5475), .Z(n5477) );
  XNOR U5131 ( .A(n5478), .B(n5479), .Z(n5475) );
  AND U5132 ( .A(n1123), .B(n5480), .Z(n5479) );
  XOR U5133 ( .A(n5481), .B(n5482), .Z(n5473) );
  AND U5134 ( .A(n1127), .B(n5483), .Z(n5482) );
  XOR U5135 ( .A(n5484), .B(n5485), .Z(n5470) );
  AND U5136 ( .A(n1131), .B(n5483), .Z(n5485) );
  XNOR U5137 ( .A(n5486), .B(n5484), .Z(n5483) );
  IV U5138 ( .A(n5481), .Z(n5486) );
  XOR U5139 ( .A(n5487), .B(n5488), .Z(n5481) );
  AND U5140 ( .A(n1134), .B(n5480), .Z(n5488) );
  XNOR U5141 ( .A(n5478), .B(n5487), .Z(n5480) );
  XNOR U5142 ( .A(n5489), .B(n5490), .Z(n5478) );
  AND U5143 ( .A(n1138), .B(n5491), .Z(n5490) );
  XOR U5144 ( .A(p_input[1700]), .B(n5489), .Z(n5491) );
  XNOR U5145 ( .A(n5492), .B(n5493), .Z(n5489) );
  AND U5146 ( .A(n1142), .B(n5494), .Z(n5493) );
  XOR U5147 ( .A(n5495), .B(n5496), .Z(n5487) );
  AND U5148 ( .A(n1146), .B(n5497), .Z(n5496) );
  XOR U5149 ( .A(n5498), .B(n5499), .Z(n5484) );
  AND U5150 ( .A(n1150), .B(n5497), .Z(n5499) );
  XNOR U5151 ( .A(n5500), .B(n5498), .Z(n5497) );
  IV U5152 ( .A(n5495), .Z(n5500) );
  XOR U5153 ( .A(n5501), .B(n5502), .Z(n5495) );
  AND U5154 ( .A(n1153), .B(n5494), .Z(n5502) );
  XNOR U5155 ( .A(n5492), .B(n5501), .Z(n5494) );
  XNOR U5156 ( .A(n5503), .B(n5504), .Z(n5492) );
  AND U5157 ( .A(n1157), .B(n5505), .Z(n5504) );
  XOR U5158 ( .A(p_input[1732]), .B(n5503), .Z(n5505) );
  XNOR U5159 ( .A(n5506), .B(n5507), .Z(n5503) );
  AND U5160 ( .A(n1161), .B(n5508), .Z(n5507) );
  XOR U5161 ( .A(n5509), .B(n5510), .Z(n5501) );
  AND U5162 ( .A(n1165), .B(n5511), .Z(n5510) );
  XOR U5163 ( .A(n5512), .B(n5513), .Z(n5498) );
  AND U5164 ( .A(n1169), .B(n5511), .Z(n5513) );
  XNOR U5165 ( .A(n5514), .B(n5512), .Z(n5511) );
  IV U5166 ( .A(n5509), .Z(n5514) );
  XOR U5167 ( .A(n5515), .B(n5516), .Z(n5509) );
  AND U5168 ( .A(n1172), .B(n5508), .Z(n5516) );
  XNOR U5169 ( .A(n5506), .B(n5515), .Z(n5508) );
  XNOR U5170 ( .A(n5517), .B(n5518), .Z(n5506) );
  AND U5171 ( .A(n1176), .B(n5519), .Z(n5518) );
  XOR U5172 ( .A(p_input[1764]), .B(n5517), .Z(n5519) );
  XNOR U5173 ( .A(n5520), .B(n5521), .Z(n5517) );
  AND U5174 ( .A(n1180), .B(n5522), .Z(n5521) );
  XOR U5175 ( .A(n5523), .B(n5524), .Z(n5515) );
  AND U5176 ( .A(n1184), .B(n5525), .Z(n5524) );
  XOR U5177 ( .A(n5526), .B(n5527), .Z(n5512) );
  AND U5178 ( .A(n1188), .B(n5525), .Z(n5527) );
  XNOR U5179 ( .A(n5528), .B(n5526), .Z(n5525) );
  IV U5180 ( .A(n5523), .Z(n5528) );
  XOR U5181 ( .A(n5529), .B(n5530), .Z(n5523) );
  AND U5182 ( .A(n1191), .B(n5522), .Z(n5530) );
  XNOR U5183 ( .A(n5520), .B(n5529), .Z(n5522) );
  XNOR U5184 ( .A(n5531), .B(n5532), .Z(n5520) );
  AND U5185 ( .A(n1195), .B(n5533), .Z(n5532) );
  XOR U5186 ( .A(p_input[1796]), .B(n5531), .Z(n5533) );
  XNOR U5187 ( .A(n5534), .B(n5535), .Z(n5531) );
  AND U5188 ( .A(n1199), .B(n5536), .Z(n5535) );
  XOR U5189 ( .A(n5537), .B(n5538), .Z(n5529) );
  AND U5190 ( .A(n1203), .B(n5539), .Z(n5538) );
  XOR U5191 ( .A(n5540), .B(n5541), .Z(n5526) );
  AND U5192 ( .A(n1207), .B(n5539), .Z(n5541) );
  XNOR U5193 ( .A(n5542), .B(n5540), .Z(n5539) );
  IV U5194 ( .A(n5537), .Z(n5542) );
  XOR U5195 ( .A(n5543), .B(n5544), .Z(n5537) );
  AND U5196 ( .A(n1210), .B(n5536), .Z(n5544) );
  XNOR U5197 ( .A(n5534), .B(n5543), .Z(n5536) );
  XNOR U5198 ( .A(n5545), .B(n5546), .Z(n5534) );
  AND U5199 ( .A(n1214), .B(n5547), .Z(n5546) );
  XOR U5200 ( .A(p_input[1828]), .B(n5545), .Z(n5547) );
  XNOR U5201 ( .A(n5548), .B(n5549), .Z(n5545) );
  AND U5202 ( .A(n1218), .B(n5550), .Z(n5549) );
  XOR U5203 ( .A(n5551), .B(n5552), .Z(n5543) );
  AND U5204 ( .A(n1222), .B(n5553), .Z(n5552) );
  XOR U5205 ( .A(n5554), .B(n5555), .Z(n5540) );
  AND U5206 ( .A(n1226), .B(n5553), .Z(n5555) );
  XNOR U5207 ( .A(n5556), .B(n5554), .Z(n5553) );
  IV U5208 ( .A(n5551), .Z(n5556) );
  XOR U5209 ( .A(n5557), .B(n5558), .Z(n5551) );
  AND U5210 ( .A(n1229), .B(n5550), .Z(n5558) );
  XNOR U5211 ( .A(n5548), .B(n5557), .Z(n5550) );
  XNOR U5212 ( .A(n5559), .B(n5560), .Z(n5548) );
  AND U5213 ( .A(n1233), .B(n5561), .Z(n5560) );
  XOR U5214 ( .A(p_input[1860]), .B(n5559), .Z(n5561) );
  XNOR U5215 ( .A(n5562), .B(n5563), .Z(n5559) );
  AND U5216 ( .A(n1237), .B(n5564), .Z(n5563) );
  XOR U5217 ( .A(n5565), .B(n5566), .Z(n5557) );
  AND U5218 ( .A(n1241), .B(n5567), .Z(n5566) );
  XOR U5219 ( .A(n5568), .B(n5569), .Z(n5554) );
  AND U5220 ( .A(n1245), .B(n5567), .Z(n5569) );
  XNOR U5221 ( .A(n5570), .B(n5568), .Z(n5567) );
  IV U5222 ( .A(n5565), .Z(n5570) );
  XOR U5223 ( .A(n5571), .B(n5572), .Z(n5565) );
  AND U5224 ( .A(n1248), .B(n5564), .Z(n5572) );
  XNOR U5225 ( .A(n5562), .B(n5571), .Z(n5564) );
  XNOR U5226 ( .A(n5573), .B(n5574), .Z(n5562) );
  AND U5227 ( .A(n1252), .B(n5575), .Z(n5574) );
  XOR U5228 ( .A(p_input[1892]), .B(n5573), .Z(n5575) );
  XNOR U5229 ( .A(n5576), .B(n5577), .Z(n5573) );
  AND U5230 ( .A(n1256), .B(n5578), .Z(n5577) );
  XOR U5231 ( .A(n5579), .B(n5580), .Z(n5571) );
  AND U5232 ( .A(n1260), .B(n5581), .Z(n5580) );
  XOR U5233 ( .A(n5582), .B(n5583), .Z(n5568) );
  AND U5234 ( .A(n1264), .B(n5581), .Z(n5583) );
  XNOR U5235 ( .A(n5584), .B(n5582), .Z(n5581) );
  IV U5236 ( .A(n5579), .Z(n5584) );
  XOR U5237 ( .A(n5585), .B(n5586), .Z(n5579) );
  AND U5238 ( .A(n1267), .B(n5578), .Z(n5586) );
  XNOR U5239 ( .A(n5576), .B(n5585), .Z(n5578) );
  XNOR U5240 ( .A(n5587), .B(n5588), .Z(n5576) );
  AND U5241 ( .A(n1271), .B(n5589), .Z(n5588) );
  XOR U5242 ( .A(p_input[1924]), .B(n5587), .Z(n5589) );
  XOR U5243 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(n5590), 
        .Z(n5587) );
  AND U5244 ( .A(n1274), .B(n5591), .Z(n5590) );
  XOR U5245 ( .A(n5592), .B(n5593), .Z(n5585) );
  AND U5246 ( .A(n1278), .B(n5594), .Z(n5593) );
  XOR U5247 ( .A(n5595), .B(n5596), .Z(n5582) );
  AND U5248 ( .A(n1282), .B(n5594), .Z(n5596) );
  XNOR U5249 ( .A(n5597), .B(n5595), .Z(n5594) );
  IV U5250 ( .A(n5592), .Z(n5597) );
  XOR U5251 ( .A(n5598), .B(n5599), .Z(n5592) );
  AND U5252 ( .A(n1285), .B(n5591), .Z(n5599) );
  XOR U5253 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(n5598), 
        .Z(n5591) );
  XOR U5254 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(n5600), 
        .Z(n5598) );
  AND U5255 ( .A(n1287), .B(n5601), .Z(n5600) );
  XOR U5256 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n5602), .Z(n5595) );
  AND U5257 ( .A(n1290), .B(n5601), .Z(n5602) );
  XOR U5258 ( .A(\knn_comb_/min_val_out[0][4] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .Z(n5601) );
  XOR U5259 ( .A(n2156), .B(n5603), .Z(o[35]) );
  AND U5260 ( .A(n122), .B(n5604), .Z(n2156) );
  XOR U5261 ( .A(n2157), .B(n5603), .Z(n5604) );
  XOR U5262 ( .A(n5605), .B(n65), .Z(n5603) );
  AND U5263 ( .A(n125), .B(n5606), .Z(n65) );
  XOR U5264 ( .A(n66), .B(n5605), .Z(n5606) );
  XOR U5265 ( .A(n5607), .B(n5608), .Z(n66) );
  AND U5266 ( .A(n130), .B(n5609), .Z(n5608) );
  XOR U5267 ( .A(p_input[3]), .B(n5607), .Z(n5609) );
  XNOR U5268 ( .A(n5610), .B(n5611), .Z(n5607) );
  AND U5269 ( .A(n134), .B(n5612), .Z(n5611) );
  XOR U5270 ( .A(n5613), .B(n5614), .Z(n5605) );
  AND U5271 ( .A(n138), .B(n5615), .Z(n5614) );
  XOR U5272 ( .A(n5616), .B(n5617), .Z(n2157) );
  AND U5273 ( .A(n142), .B(n5615), .Z(n5617) );
  XNOR U5274 ( .A(n5618), .B(n5616), .Z(n5615) );
  IV U5275 ( .A(n5613), .Z(n5618) );
  XOR U5276 ( .A(n5619), .B(n5620), .Z(n5613) );
  AND U5277 ( .A(n146), .B(n5612), .Z(n5620) );
  XNOR U5278 ( .A(n5610), .B(n5619), .Z(n5612) );
  XNOR U5279 ( .A(n5621), .B(n5622), .Z(n5610) );
  AND U5280 ( .A(n150), .B(n5623), .Z(n5622) );
  XOR U5281 ( .A(p_input[35]), .B(n5621), .Z(n5623) );
  XNOR U5282 ( .A(n5624), .B(n5625), .Z(n5621) );
  AND U5283 ( .A(n154), .B(n5626), .Z(n5625) );
  XOR U5284 ( .A(n5627), .B(n5628), .Z(n5619) );
  AND U5285 ( .A(n158), .B(n5629), .Z(n5628) );
  XOR U5286 ( .A(n5630), .B(n5631), .Z(n5616) );
  AND U5287 ( .A(n162), .B(n5629), .Z(n5631) );
  XNOR U5288 ( .A(n5632), .B(n5630), .Z(n5629) );
  IV U5289 ( .A(n5627), .Z(n5632) );
  XOR U5290 ( .A(n5633), .B(n5634), .Z(n5627) );
  AND U5291 ( .A(n165), .B(n5626), .Z(n5634) );
  XNOR U5292 ( .A(n5624), .B(n5633), .Z(n5626) );
  XNOR U5293 ( .A(n5635), .B(n5636), .Z(n5624) );
  AND U5294 ( .A(n169), .B(n5637), .Z(n5636) );
  XOR U5295 ( .A(p_input[67]), .B(n5635), .Z(n5637) );
  XNOR U5296 ( .A(n5638), .B(n5639), .Z(n5635) );
  AND U5297 ( .A(n173), .B(n5640), .Z(n5639) );
  XOR U5298 ( .A(n5641), .B(n5642), .Z(n5633) );
  AND U5299 ( .A(n177), .B(n5643), .Z(n5642) );
  XOR U5300 ( .A(n5644), .B(n5645), .Z(n5630) );
  AND U5301 ( .A(n181), .B(n5643), .Z(n5645) );
  XNOR U5302 ( .A(n5646), .B(n5644), .Z(n5643) );
  IV U5303 ( .A(n5641), .Z(n5646) );
  XOR U5304 ( .A(n5647), .B(n5648), .Z(n5641) );
  AND U5305 ( .A(n184), .B(n5640), .Z(n5648) );
  XNOR U5306 ( .A(n5638), .B(n5647), .Z(n5640) );
  XNOR U5307 ( .A(n5649), .B(n5650), .Z(n5638) );
  AND U5308 ( .A(n188), .B(n5651), .Z(n5650) );
  XOR U5309 ( .A(p_input[99]), .B(n5649), .Z(n5651) );
  XNOR U5310 ( .A(n5652), .B(n5653), .Z(n5649) );
  AND U5311 ( .A(n192), .B(n5654), .Z(n5653) );
  XOR U5312 ( .A(n5655), .B(n5656), .Z(n5647) );
  AND U5313 ( .A(n196), .B(n5657), .Z(n5656) );
  XOR U5314 ( .A(n5658), .B(n5659), .Z(n5644) );
  AND U5315 ( .A(n200), .B(n5657), .Z(n5659) );
  XNOR U5316 ( .A(n5660), .B(n5658), .Z(n5657) );
  IV U5317 ( .A(n5655), .Z(n5660) );
  XOR U5318 ( .A(n5661), .B(n5662), .Z(n5655) );
  AND U5319 ( .A(n203), .B(n5654), .Z(n5662) );
  XNOR U5320 ( .A(n5652), .B(n5661), .Z(n5654) );
  XNOR U5321 ( .A(n5663), .B(n5664), .Z(n5652) );
  AND U5322 ( .A(n207), .B(n5665), .Z(n5664) );
  XOR U5323 ( .A(p_input[131]), .B(n5663), .Z(n5665) );
  XNOR U5324 ( .A(n5666), .B(n5667), .Z(n5663) );
  AND U5325 ( .A(n211), .B(n5668), .Z(n5667) );
  XOR U5326 ( .A(n5669), .B(n5670), .Z(n5661) );
  AND U5327 ( .A(n215), .B(n5671), .Z(n5670) );
  XOR U5328 ( .A(n5672), .B(n5673), .Z(n5658) );
  AND U5329 ( .A(n219), .B(n5671), .Z(n5673) );
  XNOR U5330 ( .A(n5674), .B(n5672), .Z(n5671) );
  IV U5331 ( .A(n5669), .Z(n5674) );
  XOR U5332 ( .A(n5675), .B(n5676), .Z(n5669) );
  AND U5333 ( .A(n222), .B(n5668), .Z(n5676) );
  XNOR U5334 ( .A(n5666), .B(n5675), .Z(n5668) );
  XNOR U5335 ( .A(n5677), .B(n5678), .Z(n5666) );
  AND U5336 ( .A(n226), .B(n5679), .Z(n5678) );
  XOR U5337 ( .A(p_input[163]), .B(n5677), .Z(n5679) );
  XNOR U5338 ( .A(n5680), .B(n5681), .Z(n5677) );
  AND U5339 ( .A(n230), .B(n5682), .Z(n5681) );
  XOR U5340 ( .A(n5683), .B(n5684), .Z(n5675) );
  AND U5341 ( .A(n234), .B(n5685), .Z(n5684) );
  XOR U5342 ( .A(n5686), .B(n5687), .Z(n5672) );
  AND U5343 ( .A(n238), .B(n5685), .Z(n5687) );
  XNOR U5344 ( .A(n5688), .B(n5686), .Z(n5685) );
  IV U5345 ( .A(n5683), .Z(n5688) );
  XOR U5346 ( .A(n5689), .B(n5690), .Z(n5683) );
  AND U5347 ( .A(n241), .B(n5682), .Z(n5690) );
  XNOR U5348 ( .A(n5680), .B(n5689), .Z(n5682) );
  XNOR U5349 ( .A(n5691), .B(n5692), .Z(n5680) );
  AND U5350 ( .A(n245), .B(n5693), .Z(n5692) );
  XOR U5351 ( .A(p_input[195]), .B(n5691), .Z(n5693) );
  XNOR U5352 ( .A(n5694), .B(n5695), .Z(n5691) );
  AND U5353 ( .A(n249), .B(n5696), .Z(n5695) );
  XOR U5354 ( .A(n5697), .B(n5698), .Z(n5689) );
  AND U5355 ( .A(n253), .B(n5699), .Z(n5698) );
  XOR U5356 ( .A(n5700), .B(n5701), .Z(n5686) );
  AND U5357 ( .A(n257), .B(n5699), .Z(n5701) );
  XNOR U5358 ( .A(n5702), .B(n5700), .Z(n5699) );
  IV U5359 ( .A(n5697), .Z(n5702) );
  XOR U5360 ( .A(n5703), .B(n5704), .Z(n5697) );
  AND U5361 ( .A(n260), .B(n5696), .Z(n5704) );
  XNOR U5362 ( .A(n5694), .B(n5703), .Z(n5696) );
  XNOR U5363 ( .A(n5705), .B(n5706), .Z(n5694) );
  AND U5364 ( .A(n264), .B(n5707), .Z(n5706) );
  XOR U5365 ( .A(p_input[227]), .B(n5705), .Z(n5707) );
  XNOR U5366 ( .A(n5708), .B(n5709), .Z(n5705) );
  AND U5367 ( .A(n268), .B(n5710), .Z(n5709) );
  XOR U5368 ( .A(n5711), .B(n5712), .Z(n5703) );
  AND U5369 ( .A(n272), .B(n5713), .Z(n5712) );
  XOR U5370 ( .A(n5714), .B(n5715), .Z(n5700) );
  AND U5371 ( .A(n276), .B(n5713), .Z(n5715) );
  XNOR U5372 ( .A(n5716), .B(n5714), .Z(n5713) );
  IV U5373 ( .A(n5711), .Z(n5716) );
  XOR U5374 ( .A(n5717), .B(n5718), .Z(n5711) );
  AND U5375 ( .A(n279), .B(n5710), .Z(n5718) );
  XNOR U5376 ( .A(n5708), .B(n5717), .Z(n5710) );
  XNOR U5377 ( .A(n5719), .B(n5720), .Z(n5708) );
  AND U5378 ( .A(n283), .B(n5721), .Z(n5720) );
  XOR U5379 ( .A(p_input[259]), .B(n5719), .Z(n5721) );
  XNOR U5380 ( .A(n5722), .B(n5723), .Z(n5719) );
  AND U5381 ( .A(n287), .B(n5724), .Z(n5723) );
  XOR U5382 ( .A(n5725), .B(n5726), .Z(n5717) );
  AND U5383 ( .A(n291), .B(n5727), .Z(n5726) );
  XOR U5384 ( .A(n5728), .B(n5729), .Z(n5714) );
  AND U5385 ( .A(n295), .B(n5727), .Z(n5729) );
  XNOR U5386 ( .A(n5730), .B(n5728), .Z(n5727) );
  IV U5387 ( .A(n5725), .Z(n5730) );
  XOR U5388 ( .A(n5731), .B(n5732), .Z(n5725) );
  AND U5389 ( .A(n298), .B(n5724), .Z(n5732) );
  XNOR U5390 ( .A(n5722), .B(n5731), .Z(n5724) );
  XNOR U5391 ( .A(n5733), .B(n5734), .Z(n5722) );
  AND U5392 ( .A(n302), .B(n5735), .Z(n5734) );
  XOR U5393 ( .A(p_input[291]), .B(n5733), .Z(n5735) );
  XNOR U5394 ( .A(n5736), .B(n5737), .Z(n5733) );
  AND U5395 ( .A(n306), .B(n5738), .Z(n5737) );
  XOR U5396 ( .A(n5739), .B(n5740), .Z(n5731) );
  AND U5397 ( .A(n310), .B(n5741), .Z(n5740) );
  XOR U5398 ( .A(n5742), .B(n5743), .Z(n5728) );
  AND U5399 ( .A(n314), .B(n5741), .Z(n5743) );
  XNOR U5400 ( .A(n5744), .B(n5742), .Z(n5741) );
  IV U5401 ( .A(n5739), .Z(n5744) );
  XOR U5402 ( .A(n5745), .B(n5746), .Z(n5739) );
  AND U5403 ( .A(n317), .B(n5738), .Z(n5746) );
  XNOR U5404 ( .A(n5736), .B(n5745), .Z(n5738) );
  XNOR U5405 ( .A(n5747), .B(n5748), .Z(n5736) );
  AND U5406 ( .A(n321), .B(n5749), .Z(n5748) );
  XOR U5407 ( .A(p_input[323]), .B(n5747), .Z(n5749) );
  XNOR U5408 ( .A(n5750), .B(n5751), .Z(n5747) );
  AND U5409 ( .A(n325), .B(n5752), .Z(n5751) );
  XOR U5410 ( .A(n5753), .B(n5754), .Z(n5745) );
  AND U5411 ( .A(n329), .B(n5755), .Z(n5754) );
  XOR U5412 ( .A(n5756), .B(n5757), .Z(n5742) );
  AND U5413 ( .A(n333), .B(n5755), .Z(n5757) );
  XNOR U5414 ( .A(n5758), .B(n5756), .Z(n5755) );
  IV U5415 ( .A(n5753), .Z(n5758) );
  XOR U5416 ( .A(n5759), .B(n5760), .Z(n5753) );
  AND U5417 ( .A(n336), .B(n5752), .Z(n5760) );
  XNOR U5418 ( .A(n5750), .B(n5759), .Z(n5752) );
  XNOR U5419 ( .A(n5761), .B(n5762), .Z(n5750) );
  AND U5420 ( .A(n340), .B(n5763), .Z(n5762) );
  XOR U5421 ( .A(p_input[355]), .B(n5761), .Z(n5763) );
  XNOR U5422 ( .A(n5764), .B(n5765), .Z(n5761) );
  AND U5423 ( .A(n344), .B(n5766), .Z(n5765) );
  XOR U5424 ( .A(n5767), .B(n5768), .Z(n5759) );
  AND U5425 ( .A(n348), .B(n5769), .Z(n5768) );
  XOR U5426 ( .A(n5770), .B(n5771), .Z(n5756) );
  AND U5427 ( .A(n352), .B(n5769), .Z(n5771) );
  XNOR U5428 ( .A(n5772), .B(n5770), .Z(n5769) );
  IV U5429 ( .A(n5767), .Z(n5772) );
  XOR U5430 ( .A(n5773), .B(n5774), .Z(n5767) );
  AND U5431 ( .A(n355), .B(n5766), .Z(n5774) );
  XNOR U5432 ( .A(n5764), .B(n5773), .Z(n5766) );
  XNOR U5433 ( .A(n5775), .B(n5776), .Z(n5764) );
  AND U5434 ( .A(n359), .B(n5777), .Z(n5776) );
  XOR U5435 ( .A(p_input[387]), .B(n5775), .Z(n5777) );
  XNOR U5436 ( .A(n5778), .B(n5779), .Z(n5775) );
  AND U5437 ( .A(n363), .B(n5780), .Z(n5779) );
  XOR U5438 ( .A(n5781), .B(n5782), .Z(n5773) );
  AND U5439 ( .A(n367), .B(n5783), .Z(n5782) );
  XOR U5440 ( .A(n5784), .B(n5785), .Z(n5770) );
  AND U5441 ( .A(n371), .B(n5783), .Z(n5785) );
  XNOR U5442 ( .A(n5786), .B(n5784), .Z(n5783) );
  IV U5443 ( .A(n5781), .Z(n5786) );
  XOR U5444 ( .A(n5787), .B(n5788), .Z(n5781) );
  AND U5445 ( .A(n374), .B(n5780), .Z(n5788) );
  XNOR U5446 ( .A(n5778), .B(n5787), .Z(n5780) );
  XNOR U5447 ( .A(n5789), .B(n5790), .Z(n5778) );
  AND U5448 ( .A(n378), .B(n5791), .Z(n5790) );
  XOR U5449 ( .A(p_input[419]), .B(n5789), .Z(n5791) );
  XNOR U5450 ( .A(n5792), .B(n5793), .Z(n5789) );
  AND U5451 ( .A(n382), .B(n5794), .Z(n5793) );
  XOR U5452 ( .A(n5795), .B(n5796), .Z(n5787) );
  AND U5453 ( .A(n386), .B(n5797), .Z(n5796) );
  XOR U5454 ( .A(n5798), .B(n5799), .Z(n5784) );
  AND U5455 ( .A(n390), .B(n5797), .Z(n5799) );
  XNOR U5456 ( .A(n5800), .B(n5798), .Z(n5797) );
  IV U5457 ( .A(n5795), .Z(n5800) );
  XOR U5458 ( .A(n5801), .B(n5802), .Z(n5795) );
  AND U5459 ( .A(n393), .B(n5794), .Z(n5802) );
  XNOR U5460 ( .A(n5792), .B(n5801), .Z(n5794) );
  XNOR U5461 ( .A(n5803), .B(n5804), .Z(n5792) );
  AND U5462 ( .A(n397), .B(n5805), .Z(n5804) );
  XOR U5463 ( .A(p_input[451]), .B(n5803), .Z(n5805) );
  XNOR U5464 ( .A(n5806), .B(n5807), .Z(n5803) );
  AND U5465 ( .A(n401), .B(n5808), .Z(n5807) );
  XOR U5466 ( .A(n5809), .B(n5810), .Z(n5801) );
  AND U5467 ( .A(n405), .B(n5811), .Z(n5810) );
  XOR U5468 ( .A(n5812), .B(n5813), .Z(n5798) );
  AND U5469 ( .A(n409), .B(n5811), .Z(n5813) );
  XNOR U5470 ( .A(n5814), .B(n5812), .Z(n5811) );
  IV U5471 ( .A(n5809), .Z(n5814) );
  XOR U5472 ( .A(n5815), .B(n5816), .Z(n5809) );
  AND U5473 ( .A(n412), .B(n5808), .Z(n5816) );
  XNOR U5474 ( .A(n5806), .B(n5815), .Z(n5808) );
  XNOR U5475 ( .A(n5817), .B(n5818), .Z(n5806) );
  AND U5476 ( .A(n416), .B(n5819), .Z(n5818) );
  XOR U5477 ( .A(p_input[483]), .B(n5817), .Z(n5819) );
  XNOR U5478 ( .A(n5820), .B(n5821), .Z(n5817) );
  AND U5479 ( .A(n420), .B(n5822), .Z(n5821) );
  XOR U5480 ( .A(n5823), .B(n5824), .Z(n5815) );
  AND U5481 ( .A(n424), .B(n5825), .Z(n5824) );
  XOR U5482 ( .A(n5826), .B(n5827), .Z(n5812) );
  AND U5483 ( .A(n428), .B(n5825), .Z(n5827) );
  XNOR U5484 ( .A(n5828), .B(n5826), .Z(n5825) );
  IV U5485 ( .A(n5823), .Z(n5828) );
  XOR U5486 ( .A(n5829), .B(n5830), .Z(n5823) );
  AND U5487 ( .A(n431), .B(n5822), .Z(n5830) );
  XNOR U5488 ( .A(n5820), .B(n5829), .Z(n5822) );
  XNOR U5489 ( .A(n5831), .B(n5832), .Z(n5820) );
  AND U5490 ( .A(n435), .B(n5833), .Z(n5832) );
  XOR U5491 ( .A(p_input[515]), .B(n5831), .Z(n5833) );
  XNOR U5492 ( .A(n5834), .B(n5835), .Z(n5831) );
  AND U5493 ( .A(n439), .B(n5836), .Z(n5835) );
  XOR U5494 ( .A(n5837), .B(n5838), .Z(n5829) );
  AND U5495 ( .A(n443), .B(n5839), .Z(n5838) );
  XOR U5496 ( .A(n5840), .B(n5841), .Z(n5826) );
  AND U5497 ( .A(n447), .B(n5839), .Z(n5841) );
  XNOR U5498 ( .A(n5842), .B(n5840), .Z(n5839) );
  IV U5499 ( .A(n5837), .Z(n5842) );
  XOR U5500 ( .A(n5843), .B(n5844), .Z(n5837) );
  AND U5501 ( .A(n450), .B(n5836), .Z(n5844) );
  XNOR U5502 ( .A(n5834), .B(n5843), .Z(n5836) );
  XNOR U5503 ( .A(n5845), .B(n5846), .Z(n5834) );
  AND U5504 ( .A(n454), .B(n5847), .Z(n5846) );
  XOR U5505 ( .A(p_input[547]), .B(n5845), .Z(n5847) );
  XNOR U5506 ( .A(n5848), .B(n5849), .Z(n5845) );
  AND U5507 ( .A(n458), .B(n5850), .Z(n5849) );
  XOR U5508 ( .A(n5851), .B(n5852), .Z(n5843) );
  AND U5509 ( .A(n462), .B(n5853), .Z(n5852) );
  XOR U5510 ( .A(n5854), .B(n5855), .Z(n5840) );
  AND U5511 ( .A(n466), .B(n5853), .Z(n5855) );
  XNOR U5512 ( .A(n5856), .B(n5854), .Z(n5853) );
  IV U5513 ( .A(n5851), .Z(n5856) );
  XOR U5514 ( .A(n5857), .B(n5858), .Z(n5851) );
  AND U5515 ( .A(n469), .B(n5850), .Z(n5858) );
  XNOR U5516 ( .A(n5848), .B(n5857), .Z(n5850) );
  XNOR U5517 ( .A(n5859), .B(n5860), .Z(n5848) );
  AND U5518 ( .A(n473), .B(n5861), .Z(n5860) );
  XOR U5519 ( .A(p_input[579]), .B(n5859), .Z(n5861) );
  XNOR U5520 ( .A(n5862), .B(n5863), .Z(n5859) );
  AND U5521 ( .A(n477), .B(n5864), .Z(n5863) );
  XOR U5522 ( .A(n5865), .B(n5866), .Z(n5857) );
  AND U5523 ( .A(n481), .B(n5867), .Z(n5866) );
  XOR U5524 ( .A(n5868), .B(n5869), .Z(n5854) );
  AND U5525 ( .A(n485), .B(n5867), .Z(n5869) );
  XNOR U5526 ( .A(n5870), .B(n5868), .Z(n5867) );
  IV U5527 ( .A(n5865), .Z(n5870) );
  XOR U5528 ( .A(n5871), .B(n5872), .Z(n5865) );
  AND U5529 ( .A(n488), .B(n5864), .Z(n5872) );
  XNOR U5530 ( .A(n5862), .B(n5871), .Z(n5864) );
  XNOR U5531 ( .A(n5873), .B(n5874), .Z(n5862) );
  AND U5532 ( .A(n492), .B(n5875), .Z(n5874) );
  XOR U5533 ( .A(p_input[611]), .B(n5873), .Z(n5875) );
  XNOR U5534 ( .A(n5876), .B(n5877), .Z(n5873) );
  AND U5535 ( .A(n496), .B(n5878), .Z(n5877) );
  XOR U5536 ( .A(n5879), .B(n5880), .Z(n5871) );
  AND U5537 ( .A(n500), .B(n5881), .Z(n5880) );
  XOR U5538 ( .A(n5882), .B(n5883), .Z(n5868) );
  AND U5539 ( .A(n504), .B(n5881), .Z(n5883) );
  XNOR U5540 ( .A(n5884), .B(n5882), .Z(n5881) );
  IV U5541 ( .A(n5879), .Z(n5884) );
  XOR U5542 ( .A(n5885), .B(n5886), .Z(n5879) );
  AND U5543 ( .A(n507), .B(n5878), .Z(n5886) );
  XNOR U5544 ( .A(n5876), .B(n5885), .Z(n5878) );
  XNOR U5545 ( .A(n5887), .B(n5888), .Z(n5876) );
  AND U5546 ( .A(n511), .B(n5889), .Z(n5888) );
  XOR U5547 ( .A(p_input[643]), .B(n5887), .Z(n5889) );
  XNOR U5548 ( .A(n5890), .B(n5891), .Z(n5887) );
  AND U5549 ( .A(n515), .B(n5892), .Z(n5891) );
  XOR U5550 ( .A(n5893), .B(n5894), .Z(n5885) );
  AND U5551 ( .A(n519), .B(n5895), .Z(n5894) );
  XOR U5552 ( .A(n5896), .B(n5897), .Z(n5882) );
  AND U5553 ( .A(n523), .B(n5895), .Z(n5897) );
  XNOR U5554 ( .A(n5898), .B(n5896), .Z(n5895) );
  IV U5555 ( .A(n5893), .Z(n5898) );
  XOR U5556 ( .A(n5899), .B(n5900), .Z(n5893) );
  AND U5557 ( .A(n526), .B(n5892), .Z(n5900) );
  XNOR U5558 ( .A(n5890), .B(n5899), .Z(n5892) );
  XNOR U5559 ( .A(n5901), .B(n5902), .Z(n5890) );
  AND U5560 ( .A(n530), .B(n5903), .Z(n5902) );
  XOR U5561 ( .A(p_input[675]), .B(n5901), .Z(n5903) );
  XNOR U5562 ( .A(n5904), .B(n5905), .Z(n5901) );
  AND U5563 ( .A(n534), .B(n5906), .Z(n5905) );
  XOR U5564 ( .A(n5907), .B(n5908), .Z(n5899) );
  AND U5565 ( .A(n538), .B(n5909), .Z(n5908) );
  XOR U5566 ( .A(n5910), .B(n5911), .Z(n5896) );
  AND U5567 ( .A(n542), .B(n5909), .Z(n5911) );
  XNOR U5568 ( .A(n5912), .B(n5910), .Z(n5909) );
  IV U5569 ( .A(n5907), .Z(n5912) );
  XOR U5570 ( .A(n5913), .B(n5914), .Z(n5907) );
  AND U5571 ( .A(n545), .B(n5906), .Z(n5914) );
  XNOR U5572 ( .A(n5904), .B(n5913), .Z(n5906) );
  XNOR U5573 ( .A(n5915), .B(n5916), .Z(n5904) );
  AND U5574 ( .A(n549), .B(n5917), .Z(n5916) );
  XOR U5575 ( .A(p_input[707]), .B(n5915), .Z(n5917) );
  XNOR U5576 ( .A(n5918), .B(n5919), .Z(n5915) );
  AND U5577 ( .A(n553), .B(n5920), .Z(n5919) );
  XOR U5578 ( .A(n5921), .B(n5922), .Z(n5913) );
  AND U5579 ( .A(n557), .B(n5923), .Z(n5922) );
  XOR U5580 ( .A(n5924), .B(n5925), .Z(n5910) );
  AND U5581 ( .A(n561), .B(n5923), .Z(n5925) );
  XNOR U5582 ( .A(n5926), .B(n5924), .Z(n5923) );
  IV U5583 ( .A(n5921), .Z(n5926) );
  XOR U5584 ( .A(n5927), .B(n5928), .Z(n5921) );
  AND U5585 ( .A(n564), .B(n5920), .Z(n5928) );
  XNOR U5586 ( .A(n5918), .B(n5927), .Z(n5920) );
  XNOR U5587 ( .A(n5929), .B(n5930), .Z(n5918) );
  AND U5588 ( .A(n568), .B(n5931), .Z(n5930) );
  XOR U5589 ( .A(p_input[739]), .B(n5929), .Z(n5931) );
  XNOR U5590 ( .A(n5932), .B(n5933), .Z(n5929) );
  AND U5591 ( .A(n572), .B(n5934), .Z(n5933) );
  XOR U5592 ( .A(n5935), .B(n5936), .Z(n5927) );
  AND U5593 ( .A(n576), .B(n5937), .Z(n5936) );
  XOR U5594 ( .A(n5938), .B(n5939), .Z(n5924) );
  AND U5595 ( .A(n580), .B(n5937), .Z(n5939) );
  XNOR U5596 ( .A(n5940), .B(n5938), .Z(n5937) );
  IV U5597 ( .A(n5935), .Z(n5940) );
  XOR U5598 ( .A(n5941), .B(n5942), .Z(n5935) );
  AND U5599 ( .A(n583), .B(n5934), .Z(n5942) );
  XNOR U5600 ( .A(n5932), .B(n5941), .Z(n5934) );
  XNOR U5601 ( .A(n5943), .B(n5944), .Z(n5932) );
  AND U5602 ( .A(n587), .B(n5945), .Z(n5944) );
  XOR U5603 ( .A(p_input[771]), .B(n5943), .Z(n5945) );
  XNOR U5604 ( .A(n5946), .B(n5947), .Z(n5943) );
  AND U5605 ( .A(n591), .B(n5948), .Z(n5947) );
  XOR U5606 ( .A(n5949), .B(n5950), .Z(n5941) );
  AND U5607 ( .A(n595), .B(n5951), .Z(n5950) );
  XOR U5608 ( .A(n5952), .B(n5953), .Z(n5938) );
  AND U5609 ( .A(n599), .B(n5951), .Z(n5953) );
  XNOR U5610 ( .A(n5954), .B(n5952), .Z(n5951) );
  IV U5611 ( .A(n5949), .Z(n5954) );
  XOR U5612 ( .A(n5955), .B(n5956), .Z(n5949) );
  AND U5613 ( .A(n602), .B(n5948), .Z(n5956) );
  XNOR U5614 ( .A(n5946), .B(n5955), .Z(n5948) );
  XNOR U5615 ( .A(n5957), .B(n5958), .Z(n5946) );
  AND U5616 ( .A(n606), .B(n5959), .Z(n5958) );
  XOR U5617 ( .A(p_input[803]), .B(n5957), .Z(n5959) );
  XNOR U5618 ( .A(n5960), .B(n5961), .Z(n5957) );
  AND U5619 ( .A(n610), .B(n5962), .Z(n5961) );
  XOR U5620 ( .A(n5963), .B(n5964), .Z(n5955) );
  AND U5621 ( .A(n614), .B(n5965), .Z(n5964) );
  XOR U5622 ( .A(n5966), .B(n5967), .Z(n5952) );
  AND U5623 ( .A(n618), .B(n5965), .Z(n5967) );
  XNOR U5624 ( .A(n5968), .B(n5966), .Z(n5965) );
  IV U5625 ( .A(n5963), .Z(n5968) );
  XOR U5626 ( .A(n5969), .B(n5970), .Z(n5963) );
  AND U5627 ( .A(n621), .B(n5962), .Z(n5970) );
  XNOR U5628 ( .A(n5960), .B(n5969), .Z(n5962) );
  XNOR U5629 ( .A(n5971), .B(n5972), .Z(n5960) );
  AND U5630 ( .A(n625), .B(n5973), .Z(n5972) );
  XOR U5631 ( .A(p_input[835]), .B(n5971), .Z(n5973) );
  XNOR U5632 ( .A(n5974), .B(n5975), .Z(n5971) );
  AND U5633 ( .A(n629), .B(n5976), .Z(n5975) );
  XOR U5634 ( .A(n5977), .B(n5978), .Z(n5969) );
  AND U5635 ( .A(n633), .B(n5979), .Z(n5978) );
  XOR U5636 ( .A(n5980), .B(n5981), .Z(n5966) );
  AND U5637 ( .A(n637), .B(n5979), .Z(n5981) );
  XNOR U5638 ( .A(n5982), .B(n5980), .Z(n5979) );
  IV U5639 ( .A(n5977), .Z(n5982) );
  XOR U5640 ( .A(n5983), .B(n5984), .Z(n5977) );
  AND U5641 ( .A(n640), .B(n5976), .Z(n5984) );
  XNOR U5642 ( .A(n5974), .B(n5983), .Z(n5976) );
  XNOR U5643 ( .A(n5985), .B(n5986), .Z(n5974) );
  AND U5644 ( .A(n644), .B(n5987), .Z(n5986) );
  XOR U5645 ( .A(p_input[867]), .B(n5985), .Z(n5987) );
  XNOR U5646 ( .A(n5988), .B(n5989), .Z(n5985) );
  AND U5647 ( .A(n648), .B(n5990), .Z(n5989) );
  XOR U5648 ( .A(n5991), .B(n5992), .Z(n5983) );
  AND U5649 ( .A(n652), .B(n5993), .Z(n5992) );
  XOR U5650 ( .A(n5994), .B(n5995), .Z(n5980) );
  AND U5651 ( .A(n656), .B(n5993), .Z(n5995) );
  XNOR U5652 ( .A(n5996), .B(n5994), .Z(n5993) );
  IV U5653 ( .A(n5991), .Z(n5996) );
  XOR U5654 ( .A(n5997), .B(n5998), .Z(n5991) );
  AND U5655 ( .A(n659), .B(n5990), .Z(n5998) );
  XNOR U5656 ( .A(n5988), .B(n5997), .Z(n5990) );
  XNOR U5657 ( .A(n5999), .B(n6000), .Z(n5988) );
  AND U5658 ( .A(n663), .B(n6001), .Z(n6000) );
  XOR U5659 ( .A(p_input[899]), .B(n5999), .Z(n6001) );
  XNOR U5660 ( .A(n6002), .B(n6003), .Z(n5999) );
  AND U5661 ( .A(n667), .B(n6004), .Z(n6003) );
  XOR U5662 ( .A(n6005), .B(n6006), .Z(n5997) );
  AND U5663 ( .A(n671), .B(n6007), .Z(n6006) );
  XOR U5664 ( .A(n6008), .B(n6009), .Z(n5994) );
  AND U5665 ( .A(n675), .B(n6007), .Z(n6009) );
  XNOR U5666 ( .A(n6010), .B(n6008), .Z(n6007) );
  IV U5667 ( .A(n6005), .Z(n6010) );
  XOR U5668 ( .A(n6011), .B(n6012), .Z(n6005) );
  AND U5669 ( .A(n678), .B(n6004), .Z(n6012) );
  XNOR U5670 ( .A(n6002), .B(n6011), .Z(n6004) );
  XNOR U5671 ( .A(n6013), .B(n6014), .Z(n6002) );
  AND U5672 ( .A(n682), .B(n6015), .Z(n6014) );
  XOR U5673 ( .A(p_input[931]), .B(n6013), .Z(n6015) );
  XNOR U5674 ( .A(n6016), .B(n6017), .Z(n6013) );
  AND U5675 ( .A(n686), .B(n6018), .Z(n6017) );
  XOR U5676 ( .A(n6019), .B(n6020), .Z(n6011) );
  AND U5677 ( .A(n690), .B(n6021), .Z(n6020) );
  XOR U5678 ( .A(n6022), .B(n6023), .Z(n6008) );
  AND U5679 ( .A(n694), .B(n6021), .Z(n6023) );
  XNOR U5680 ( .A(n6024), .B(n6022), .Z(n6021) );
  IV U5681 ( .A(n6019), .Z(n6024) );
  XOR U5682 ( .A(n6025), .B(n6026), .Z(n6019) );
  AND U5683 ( .A(n697), .B(n6018), .Z(n6026) );
  XNOR U5684 ( .A(n6016), .B(n6025), .Z(n6018) );
  XNOR U5685 ( .A(n6027), .B(n6028), .Z(n6016) );
  AND U5686 ( .A(n701), .B(n6029), .Z(n6028) );
  XOR U5687 ( .A(p_input[963]), .B(n6027), .Z(n6029) );
  XNOR U5688 ( .A(n6030), .B(n6031), .Z(n6027) );
  AND U5689 ( .A(n705), .B(n6032), .Z(n6031) );
  XOR U5690 ( .A(n6033), .B(n6034), .Z(n6025) );
  AND U5691 ( .A(n709), .B(n6035), .Z(n6034) );
  XOR U5692 ( .A(n6036), .B(n6037), .Z(n6022) );
  AND U5693 ( .A(n713), .B(n6035), .Z(n6037) );
  XNOR U5694 ( .A(n6038), .B(n6036), .Z(n6035) );
  IV U5695 ( .A(n6033), .Z(n6038) );
  XOR U5696 ( .A(n6039), .B(n6040), .Z(n6033) );
  AND U5697 ( .A(n716), .B(n6032), .Z(n6040) );
  XNOR U5698 ( .A(n6030), .B(n6039), .Z(n6032) );
  XNOR U5699 ( .A(n6041), .B(n6042), .Z(n6030) );
  AND U5700 ( .A(n720), .B(n6043), .Z(n6042) );
  XOR U5701 ( .A(p_input[995]), .B(n6041), .Z(n6043) );
  XNOR U5702 ( .A(n6044), .B(n6045), .Z(n6041) );
  AND U5703 ( .A(n724), .B(n6046), .Z(n6045) );
  XOR U5704 ( .A(n6047), .B(n6048), .Z(n6039) );
  AND U5705 ( .A(n728), .B(n6049), .Z(n6048) );
  XOR U5706 ( .A(n6050), .B(n6051), .Z(n6036) );
  AND U5707 ( .A(n732), .B(n6049), .Z(n6051) );
  XNOR U5708 ( .A(n6052), .B(n6050), .Z(n6049) );
  IV U5709 ( .A(n6047), .Z(n6052) );
  XOR U5710 ( .A(n6053), .B(n6054), .Z(n6047) );
  AND U5711 ( .A(n735), .B(n6046), .Z(n6054) );
  XNOR U5712 ( .A(n6044), .B(n6053), .Z(n6046) );
  XNOR U5713 ( .A(n6055), .B(n6056), .Z(n6044) );
  AND U5714 ( .A(n739), .B(n6057), .Z(n6056) );
  XOR U5715 ( .A(p_input[1027]), .B(n6055), .Z(n6057) );
  XNOR U5716 ( .A(n6058), .B(n6059), .Z(n6055) );
  AND U5717 ( .A(n743), .B(n6060), .Z(n6059) );
  XOR U5718 ( .A(n6061), .B(n6062), .Z(n6053) );
  AND U5719 ( .A(n747), .B(n6063), .Z(n6062) );
  XOR U5720 ( .A(n6064), .B(n6065), .Z(n6050) );
  AND U5721 ( .A(n751), .B(n6063), .Z(n6065) );
  XNOR U5722 ( .A(n6066), .B(n6064), .Z(n6063) );
  IV U5723 ( .A(n6061), .Z(n6066) );
  XOR U5724 ( .A(n6067), .B(n6068), .Z(n6061) );
  AND U5725 ( .A(n754), .B(n6060), .Z(n6068) );
  XNOR U5726 ( .A(n6058), .B(n6067), .Z(n6060) );
  XNOR U5727 ( .A(n6069), .B(n6070), .Z(n6058) );
  AND U5728 ( .A(n758), .B(n6071), .Z(n6070) );
  XOR U5729 ( .A(p_input[1059]), .B(n6069), .Z(n6071) );
  XNOR U5730 ( .A(n6072), .B(n6073), .Z(n6069) );
  AND U5731 ( .A(n762), .B(n6074), .Z(n6073) );
  XOR U5732 ( .A(n6075), .B(n6076), .Z(n6067) );
  AND U5733 ( .A(n766), .B(n6077), .Z(n6076) );
  XOR U5734 ( .A(n6078), .B(n6079), .Z(n6064) );
  AND U5735 ( .A(n770), .B(n6077), .Z(n6079) );
  XNOR U5736 ( .A(n6080), .B(n6078), .Z(n6077) );
  IV U5737 ( .A(n6075), .Z(n6080) );
  XOR U5738 ( .A(n6081), .B(n6082), .Z(n6075) );
  AND U5739 ( .A(n773), .B(n6074), .Z(n6082) );
  XNOR U5740 ( .A(n6072), .B(n6081), .Z(n6074) );
  XNOR U5741 ( .A(n6083), .B(n6084), .Z(n6072) );
  AND U5742 ( .A(n777), .B(n6085), .Z(n6084) );
  XOR U5743 ( .A(p_input[1091]), .B(n6083), .Z(n6085) );
  XNOR U5744 ( .A(n6086), .B(n6087), .Z(n6083) );
  AND U5745 ( .A(n781), .B(n6088), .Z(n6087) );
  XOR U5746 ( .A(n6089), .B(n6090), .Z(n6081) );
  AND U5747 ( .A(n785), .B(n6091), .Z(n6090) );
  XOR U5748 ( .A(n6092), .B(n6093), .Z(n6078) );
  AND U5749 ( .A(n789), .B(n6091), .Z(n6093) );
  XNOR U5750 ( .A(n6094), .B(n6092), .Z(n6091) );
  IV U5751 ( .A(n6089), .Z(n6094) );
  XOR U5752 ( .A(n6095), .B(n6096), .Z(n6089) );
  AND U5753 ( .A(n792), .B(n6088), .Z(n6096) );
  XNOR U5754 ( .A(n6086), .B(n6095), .Z(n6088) );
  XNOR U5755 ( .A(n6097), .B(n6098), .Z(n6086) );
  AND U5756 ( .A(n796), .B(n6099), .Z(n6098) );
  XOR U5757 ( .A(p_input[1123]), .B(n6097), .Z(n6099) );
  XNOR U5758 ( .A(n6100), .B(n6101), .Z(n6097) );
  AND U5759 ( .A(n800), .B(n6102), .Z(n6101) );
  XOR U5760 ( .A(n6103), .B(n6104), .Z(n6095) );
  AND U5761 ( .A(n804), .B(n6105), .Z(n6104) );
  XOR U5762 ( .A(n6106), .B(n6107), .Z(n6092) );
  AND U5763 ( .A(n808), .B(n6105), .Z(n6107) );
  XNOR U5764 ( .A(n6108), .B(n6106), .Z(n6105) );
  IV U5765 ( .A(n6103), .Z(n6108) );
  XOR U5766 ( .A(n6109), .B(n6110), .Z(n6103) );
  AND U5767 ( .A(n811), .B(n6102), .Z(n6110) );
  XNOR U5768 ( .A(n6100), .B(n6109), .Z(n6102) );
  XNOR U5769 ( .A(n6111), .B(n6112), .Z(n6100) );
  AND U5770 ( .A(n815), .B(n6113), .Z(n6112) );
  XOR U5771 ( .A(p_input[1155]), .B(n6111), .Z(n6113) );
  XNOR U5772 ( .A(n6114), .B(n6115), .Z(n6111) );
  AND U5773 ( .A(n819), .B(n6116), .Z(n6115) );
  XOR U5774 ( .A(n6117), .B(n6118), .Z(n6109) );
  AND U5775 ( .A(n823), .B(n6119), .Z(n6118) );
  XOR U5776 ( .A(n6120), .B(n6121), .Z(n6106) );
  AND U5777 ( .A(n827), .B(n6119), .Z(n6121) );
  XNOR U5778 ( .A(n6122), .B(n6120), .Z(n6119) );
  IV U5779 ( .A(n6117), .Z(n6122) );
  XOR U5780 ( .A(n6123), .B(n6124), .Z(n6117) );
  AND U5781 ( .A(n830), .B(n6116), .Z(n6124) );
  XNOR U5782 ( .A(n6114), .B(n6123), .Z(n6116) );
  XNOR U5783 ( .A(n6125), .B(n6126), .Z(n6114) );
  AND U5784 ( .A(n834), .B(n6127), .Z(n6126) );
  XOR U5785 ( .A(p_input[1187]), .B(n6125), .Z(n6127) );
  XNOR U5786 ( .A(n6128), .B(n6129), .Z(n6125) );
  AND U5787 ( .A(n838), .B(n6130), .Z(n6129) );
  XOR U5788 ( .A(n6131), .B(n6132), .Z(n6123) );
  AND U5789 ( .A(n842), .B(n6133), .Z(n6132) );
  XOR U5790 ( .A(n6134), .B(n6135), .Z(n6120) );
  AND U5791 ( .A(n846), .B(n6133), .Z(n6135) );
  XNOR U5792 ( .A(n6136), .B(n6134), .Z(n6133) );
  IV U5793 ( .A(n6131), .Z(n6136) );
  XOR U5794 ( .A(n6137), .B(n6138), .Z(n6131) );
  AND U5795 ( .A(n849), .B(n6130), .Z(n6138) );
  XNOR U5796 ( .A(n6128), .B(n6137), .Z(n6130) );
  XNOR U5797 ( .A(n6139), .B(n6140), .Z(n6128) );
  AND U5798 ( .A(n853), .B(n6141), .Z(n6140) );
  XOR U5799 ( .A(p_input[1219]), .B(n6139), .Z(n6141) );
  XNOR U5800 ( .A(n6142), .B(n6143), .Z(n6139) );
  AND U5801 ( .A(n857), .B(n6144), .Z(n6143) );
  XOR U5802 ( .A(n6145), .B(n6146), .Z(n6137) );
  AND U5803 ( .A(n861), .B(n6147), .Z(n6146) );
  XOR U5804 ( .A(n6148), .B(n6149), .Z(n6134) );
  AND U5805 ( .A(n865), .B(n6147), .Z(n6149) );
  XNOR U5806 ( .A(n6150), .B(n6148), .Z(n6147) );
  IV U5807 ( .A(n6145), .Z(n6150) );
  XOR U5808 ( .A(n6151), .B(n6152), .Z(n6145) );
  AND U5809 ( .A(n868), .B(n6144), .Z(n6152) );
  XNOR U5810 ( .A(n6142), .B(n6151), .Z(n6144) );
  XNOR U5811 ( .A(n6153), .B(n6154), .Z(n6142) );
  AND U5812 ( .A(n872), .B(n6155), .Z(n6154) );
  XOR U5813 ( .A(p_input[1251]), .B(n6153), .Z(n6155) );
  XNOR U5814 ( .A(n6156), .B(n6157), .Z(n6153) );
  AND U5815 ( .A(n876), .B(n6158), .Z(n6157) );
  XOR U5816 ( .A(n6159), .B(n6160), .Z(n6151) );
  AND U5817 ( .A(n880), .B(n6161), .Z(n6160) );
  XOR U5818 ( .A(n6162), .B(n6163), .Z(n6148) );
  AND U5819 ( .A(n884), .B(n6161), .Z(n6163) );
  XNOR U5820 ( .A(n6164), .B(n6162), .Z(n6161) );
  IV U5821 ( .A(n6159), .Z(n6164) );
  XOR U5822 ( .A(n6165), .B(n6166), .Z(n6159) );
  AND U5823 ( .A(n887), .B(n6158), .Z(n6166) );
  XNOR U5824 ( .A(n6156), .B(n6165), .Z(n6158) );
  XNOR U5825 ( .A(n6167), .B(n6168), .Z(n6156) );
  AND U5826 ( .A(n891), .B(n6169), .Z(n6168) );
  XOR U5827 ( .A(p_input[1283]), .B(n6167), .Z(n6169) );
  XNOR U5828 ( .A(n6170), .B(n6171), .Z(n6167) );
  AND U5829 ( .A(n895), .B(n6172), .Z(n6171) );
  XOR U5830 ( .A(n6173), .B(n6174), .Z(n6165) );
  AND U5831 ( .A(n899), .B(n6175), .Z(n6174) );
  XOR U5832 ( .A(n6176), .B(n6177), .Z(n6162) );
  AND U5833 ( .A(n903), .B(n6175), .Z(n6177) );
  XNOR U5834 ( .A(n6178), .B(n6176), .Z(n6175) );
  IV U5835 ( .A(n6173), .Z(n6178) );
  XOR U5836 ( .A(n6179), .B(n6180), .Z(n6173) );
  AND U5837 ( .A(n906), .B(n6172), .Z(n6180) );
  XNOR U5838 ( .A(n6170), .B(n6179), .Z(n6172) );
  XNOR U5839 ( .A(n6181), .B(n6182), .Z(n6170) );
  AND U5840 ( .A(n910), .B(n6183), .Z(n6182) );
  XOR U5841 ( .A(p_input[1315]), .B(n6181), .Z(n6183) );
  XNOR U5842 ( .A(n6184), .B(n6185), .Z(n6181) );
  AND U5843 ( .A(n914), .B(n6186), .Z(n6185) );
  XOR U5844 ( .A(n6187), .B(n6188), .Z(n6179) );
  AND U5845 ( .A(n918), .B(n6189), .Z(n6188) );
  XOR U5846 ( .A(n6190), .B(n6191), .Z(n6176) );
  AND U5847 ( .A(n922), .B(n6189), .Z(n6191) );
  XNOR U5848 ( .A(n6192), .B(n6190), .Z(n6189) );
  IV U5849 ( .A(n6187), .Z(n6192) );
  XOR U5850 ( .A(n6193), .B(n6194), .Z(n6187) );
  AND U5851 ( .A(n925), .B(n6186), .Z(n6194) );
  XNOR U5852 ( .A(n6184), .B(n6193), .Z(n6186) );
  XNOR U5853 ( .A(n6195), .B(n6196), .Z(n6184) );
  AND U5854 ( .A(n929), .B(n6197), .Z(n6196) );
  XOR U5855 ( .A(p_input[1347]), .B(n6195), .Z(n6197) );
  XNOR U5856 ( .A(n6198), .B(n6199), .Z(n6195) );
  AND U5857 ( .A(n933), .B(n6200), .Z(n6199) );
  XOR U5858 ( .A(n6201), .B(n6202), .Z(n6193) );
  AND U5859 ( .A(n937), .B(n6203), .Z(n6202) );
  XOR U5860 ( .A(n6204), .B(n6205), .Z(n6190) );
  AND U5861 ( .A(n941), .B(n6203), .Z(n6205) );
  XNOR U5862 ( .A(n6206), .B(n6204), .Z(n6203) );
  IV U5863 ( .A(n6201), .Z(n6206) );
  XOR U5864 ( .A(n6207), .B(n6208), .Z(n6201) );
  AND U5865 ( .A(n944), .B(n6200), .Z(n6208) );
  XNOR U5866 ( .A(n6198), .B(n6207), .Z(n6200) );
  XNOR U5867 ( .A(n6209), .B(n6210), .Z(n6198) );
  AND U5868 ( .A(n948), .B(n6211), .Z(n6210) );
  XOR U5869 ( .A(p_input[1379]), .B(n6209), .Z(n6211) );
  XNOR U5870 ( .A(n6212), .B(n6213), .Z(n6209) );
  AND U5871 ( .A(n952), .B(n6214), .Z(n6213) );
  XOR U5872 ( .A(n6215), .B(n6216), .Z(n6207) );
  AND U5873 ( .A(n956), .B(n6217), .Z(n6216) );
  XOR U5874 ( .A(n6218), .B(n6219), .Z(n6204) );
  AND U5875 ( .A(n960), .B(n6217), .Z(n6219) );
  XNOR U5876 ( .A(n6220), .B(n6218), .Z(n6217) );
  IV U5877 ( .A(n6215), .Z(n6220) );
  XOR U5878 ( .A(n6221), .B(n6222), .Z(n6215) );
  AND U5879 ( .A(n963), .B(n6214), .Z(n6222) );
  XNOR U5880 ( .A(n6212), .B(n6221), .Z(n6214) );
  XNOR U5881 ( .A(n6223), .B(n6224), .Z(n6212) );
  AND U5882 ( .A(n967), .B(n6225), .Z(n6224) );
  XOR U5883 ( .A(p_input[1411]), .B(n6223), .Z(n6225) );
  XNOR U5884 ( .A(n6226), .B(n6227), .Z(n6223) );
  AND U5885 ( .A(n971), .B(n6228), .Z(n6227) );
  XOR U5886 ( .A(n6229), .B(n6230), .Z(n6221) );
  AND U5887 ( .A(n975), .B(n6231), .Z(n6230) );
  XOR U5888 ( .A(n6232), .B(n6233), .Z(n6218) );
  AND U5889 ( .A(n979), .B(n6231), .Z(n6233) );
  XNOR U5890 ( .A(n6234), .B(n6232), .Z(n6231) );
  IV U5891 ( .A(n6229), .Z(n6234) );
  XOR U5892 ( .A(n6235), .B(n6236), .Z(n6229) );
  AND U5893 ( .A(n982), .B(n6228), .Z(n6236) );
  XNOR U5894 ( .A(n6226), .B(n6235), .Z(n6228) );
  XNOR U5895 ( .A(n6237), .B(n6238), .Z(n6226) );
  AND U5896 ( .A(n986), .B(n6239), .Z(n6238) );
  XOR U5897 ( .A(p_input[1443]), .B(n6237), .Z(n6239) );
  XNOR U5898 ( .A(n6240), .B(n6241), .Z(n6237) );
  AND U5899 ( .A(n990), .B(n6242), .Z(n6241) );
  XOR U5900 ( .A(n6243), .B(n6244), .Z(n6235) );
  AND U5901 ( .A(n994), .B(n6245), .Z(n6244) );
  XOR U5902 ( .A(n6246), .B(n6247), .Z(n6232) );
  AND U5903 ( .A(n998), .B(n6245), .Z(n6247) );
  XNOR U5904 ( .A(n6248), .B(n6246), .Z(n6245) );
  IV U5905 ( .A(n6243), .Z(n6248) );
  XOR U5906 ( .A(n6249), .B(n6250), .Z(n6243) );
  AND U5907 ( .A(n1001), .B(n6242), .Z(n6250) );
  XNOR U5908 ( .A(n6240), .B(n6249), .Z(n6242) );
  XNOR U5909 ( .A(n6251), .B(n6252), .Z(n6240) );
  AND U5910 ( .A(n1005), .B(n6253), .Z(n6252) );
  XOR U5911 ( .A(p_input[1475]), .B(n6251), .Z(n6253) );
  XNOR U5912 ( .A(n6254), .B(n6255), .Z(n6251) );
  AND U5913 ( .A(n1009), .B(n6256), .Z(n6255) );
  XOR U5914 ( .A(n6257), .B(n6258), .Z(n6249) );
  AND U5915 ( .A(n1013), .B(n6259), .Z(n6258) );
  XOR U5916 ( .A(n6260), .B(n6261), .Z(n6246) );
  AND U5917 ( .A(n1017), .B(n6259), .Z(n6261) );
  XNOR U5918 ( .A(n6262), .B(n6260), .Z(n6259) );
  IV U5919 ( .A(n6257), .Z(n6262) );
  XOR U5920 ( .A(n6263), .B(n6264), .Z(n6257) );
  AND U5921 ( .A(n1020), .B(n6256), .Z(n6264) );
  XNOR U5922 ( .A(n6254), .B(n6263), .Z(n6256) );
  XNOR U5923 ( .A(n6265), .B(n6266), .Z(n6254) );
  AND U5924 ( .A(n1024), .B(n6267), .Z(n6266) );
  XOR U5925 ( .A(p_input[1507]), .B(n6265), .Z(n6267) );
  XNOR U5926 ( .A(n6268), .B(n6269), .Z(n6265) );
  AND U5927 ( .A(n1028), .B(n6270), .Z(n6269) );
  XOR U5928 ( .A(n6271), .B(n6272), .Z(n6263) );
  AND U5929 ( .A(n1032), .B(n6273), .Z(n6272) );
  XOR U5930 ( .A(n6274), .B(n6275), .Z(n6260) );
  AND U5931 ( .A(n1036), .B(n6273), .Z(n6275) );
  XNOR U5932 ( .A(n6276), .B(n6274), .Z(n6273) );
  IV U5933 ( .A(n6271), .Z(n6276) );
  XOR U5934 ( .A(n6277), .B(n6278), .Z(n6271) );
  AND U5935 ( .A(n1039), .B(n6270), .Z(n6278) );
  XNOR U5936 ( .A(n6268), .B(n6277), .Z(n6270) );
  XNOR U5937 ( .A(n6279), .B(n6280), .Z(n6268) );
  AND U5938 ( .A(n1043), .B(n6281), .Z(n6280) );
  XOR U5939 ( .A(p_input[1539]), .B(n6279), .Z(n6281) );
  XNOR U5940 ( .A(n6282), .B(n6283), .Z(n6279) );
  AND U5941 ( .A(n1047), .B(n6284), .Z(n6283) );
  XOR U5942 ( .A(n6285), .B(n6286), .Z(n6277) );
  AND U5943 ( .A(n1051), .B(n6287), .Z(n6286) );
  XOR U5944 ( .A(n6288), .B(n6289), .Z(n6274) );
  AND U5945 ( .A(n1055), .B(n6287), .Z(n6289) );
  XNOR U5946 ( .A(n6290), .B(n6288), .Z(n6287) );
  IV U5947 ( .A(n6285), .Z(n6290) );
  XOR U5948 ( .A(n6291), .B(n6292), .Z(n6285) );
  AND U5949 ( .A(n1058), .B(n6284), .Z(n6292) );
  XNOR U5950 ( .A(n6282), .B(n6291), .Z(n6284) );
  XNOR U5951 ( .A(n6293), .B(n6294), .Z(n6282) );
  AND U5952 ( .A(n1062), .B(n6295), .Z(n6294) );
  XOR U5953 ( .A(p_input[1571]), .B(n6293), .Z(n6295) );
  XNOR U5954 ( .A(n6296), .B(n6297), .Z(n6293) );
  AND U5955 ( .A(n1066), .B(n6298), .Z(n6297) );
  XOR U5956 ( .A(n6299), .B(n6300), .Z(n6291) );
  AND U5957 ( .A(n1070), .B(n6301), .Z(n6300) );
  XOR U5958 ( .A(n6302), .B(n6303), .Z(n6288) );
  AND U5959 ( .A(n1074), .B(n6301), .Z(n6303) );
  XNOR U5960 ( .A(n6304), .B(n6302), .Z(n6301) );
  IV U5961 ( .A(n6299), .Z(n6304) );
  XOR U5962 ( .A(n6305), .B(n6306), .Z(n6299) );
  AND U5963 ( .A(n1077), .B(n6298), .Z(n6306) );
  XNOR U5964 ( .A(n6296), .B(n6305), .Z(n6298) );
  XNOR U5965 ( .A(n6307), .B(n6308), .Z(n6296) );
  AND U5966 ( .A(n1081), .B(n6309), .Z(n6308) );
  XOR U5967 ( .A(p_input[1603]), .B(n6307), .Z(n6309) );
  XNOR U5968 ( .A(n6310), .B(n6311), .Z(n6307) );
  AND U5969 ( .A(n1085), .B(n6312), .Z(n6311) );
  XOR U5970 ( .A(n6313), .B(n6314), .Z(n6305) );
  AND U5971 ( .A(n1089), .B(n6315), .Z(n6314) );
  XOR U5972 ( .A(n6316), .B(n6317), .Z(n6302) );
  AND U5973 ( .A(n1093), .B(n6315), .Z(n6317) );
  XNOR U5974 ( .A(n6318), .B(n6316), .Z(n6315) );
  IV U5975 ( .A(n6313), .Z(n6318) );
  XOR U5976 ( .A(n6319), .B(n6320), .Z(n6313) );
  AND U5977 ( .A(n1096), .B(n6312), .Z(n6320) );
  XNOR U5978 ( .A(n6310), .B(n6319), .Z(n6312) );
  XNOR U5979 ( .A(n6321), .B(n6322), .Z(n6310) );
  AND U5980 ( .A(n1100), .B(n6323), .Z(n6322) );
  XOR U5981 ( .A(p_input[1635]), .B(n6321), .Z(n6323) );
  XNOR U5982 ( .A(n6324), .B(n6325), .Z(n6321) );
  AND U5983 ( .A(n1104), .B(n6326), .Z(n6325) );
  XOR U5984 ( .A(n6327), .B(n6328), .Z(n6319) );
  AND U5985 ( .A(n1108), .B(n6329), .Z(n6328) );
  XOR U5986 ( .A(n6330), .B(n6331), .Z(n6316) );
  AND U5987 ( .A(n1112), .B(n6329), .Z(n6331) );
  XNOR U5988 ( .A(n6332), .B(n6330), .Z(n6329) );
  IV U5989 ( .A(n6327), .Z(n6332) );
  XOR U5990 ( .A(n6333), .B(n6334), .Z(n6327) );
  AND U5991 ( .A(n1115), .B(n6326), .Z(n6334) );
  XNOR U5992 ( .A(n6324), .B(n6333), .Z(n6326) );
  XNOR U5993 ( .A(n6335), .B(n6336), .Z(n6324) );
  AND U5994 ( .A(n1119), .B(n6337), .Z(n6336) );
  XOR U5995 ( .A(p_input[1667]), .B(n6335), .Z(n6337) );
  XNOR U5996 ( .A(n6338), .B(n6339), .Z(n6335) );
  AND U5997 ( .A(n1123), .B(n6340), .Z(n6339) );
  XOR U5998 ( .A(n6341), .B(n6342), .Z(n6333) );
  AND U5999 ( .A(n1127), .B(n6343), .Z(n6342) );
  XOR U6000 ( .A(n6344), .B(n6345), .Z(n6330) );
  AND U6001 ( .A(n1131), .B(n6343), .Z(n6345) );
  XNOR U6002 ( .A(n6346), .B(n6344), .Z(n6343) );
  IV U6003 ( .A(n6341), .Z(n6346) );
  XOR U6004 ( .A(n6347), .B(n6348), .Z(n6341) );
  AND U6005 ( .A(n1134), .B(n6340), .Z(n6348) );
  XNOR U6006 ( .A(n6338), .B(n6347), .Z(n6340) );
  XNOR U6007 ( .A(n6349), .B(n6350), .Z(n6338) );
  AND U6008 ( .A(n1138), .B(n6351), .Z(n6350) );
  XOR U6009 ( .A(p_input[1699]), .B(n6349), .Z(n6351) );
  XNOR U6010 ( .A(n6352), .B(n6353), .Z(n6349) );
  AND U6011 ( .A(n1142), .B(n6354), .Z(n6353) );
  XOR U6012 ( .A(n6355), .B(n6356), .Z(n6347) );
  AND U6013 ( .A(n1146), .B(n6357), .Z(n6356) );
  XOR U6014 ( .A(n6358), .B(n6359), .Z(n6344) );
  AND U6015 ( .A(n1150), .B(n6357), .Z(n6359) );
  XNOR U6016 ( .A(n6360), .B(n6358), .Z(n6357) );
  IV U6017 ( .A(n6355), .Z(n6360) );
  XOR U6018 ( .A(n6361), .B(n6362), .Z(n6355) );
  AND U6019 ( .A(n1153), .B(n6354), .Z(n6362) );
  XNOR U6020 ( .A(n6352), .B(n6361), .Z(n6354) );
  XNOR U6021 ( .A(n6363), .B(n6364), .Z(n6352) );
  AND U6022 ( .A(n1157), .B(n6365), .Z(n6364) );
  XOR U6023 ( .A(p_input[1731]), .B(n6363), .Z(n6365) );
  XNOR U6024 ( .A(n6366), .B(n6367), .Z(n6363) );
  AND U6025 ( .A(n1161), .B(n6368), .Z(n6367) );
  XOR U6026 ( .A(n6369), .B(n6370), .Z(n6361) );
  AND U6027 ( .A(n1165), .B(n6371), .Z(n6370) );
  XOR U6028 ( .A(n6372), .B(n6373), .Z(n6358) );
  AND U6029 ( .A(n1169), .B(n6371), .Z(n6373) );
  XNOR U6030 ( .A(n6374), .B(n6372), .Z(n6371) );
  IV U6031 ( .A(n6369), .Z(n6374) );
  XOR U6032 ( .A(n6375), .B(n6376), .Z(n6369) );
  AND U6033 ( .A(n1172), .B(n6368), .Z(n6376) );
  XNOR U6034 ( .A(n6366), .B(n6375), .Z(n6368) );
  XNOR U6035 ( .A(n6377), .B(n6378), .Z(n6366) );
  AND U6036 ( .A(n1176), .B(n6379), .Z(n6378) );
  XOR U6037 ( .A(p_input[1763]), .B(n6377), .Z(n6379) );
  XNOR U6038 ( .A(n6380), .B(n6381), .Z(n6377) );
  AND U6039 ( .A(n1180), .B(n6382), .Z(n6381) );
  XOR U6040 ( .A(n6383), .B(n6384), .Z(n6375) );
  AND U6041 ( .A(n1184), .B(n6385), .Z(n6384) );
  XOR U6042 ( .A(n6386), .B(n6387), .Z(n6372) );
  AND U6043 ( .A(n1188), .B(n6385), .Z(n6387) );
  XNOR U6044 ( .A(n6388), .B(n6386), .Z(n6385) );
  IV U6045 ( .A(n6383), .Z(n6388) );
  XOR U6046 ( .A(n6389), .B(n6390), .Z(n6383) );
  AND U6047 ( .A(n1191), .B(n6382), .Z(n6390) );
  XNOR U6048 ( .A(n6380), .B(n6389), .Z(n6382) );
  XNOR U6049 ( .A(n6391), .B(n6392), .Z(n6380) );
  AND U6050 ( .A(n1195), .B(n6393), .Z(n6392) );
  XOR U6051 ( .A(p_input[1795]), .B(n6391), .Z(n6393) );
  XNOR U6052 ( .A(n6394), .B(n6395), .Z(n6391) );
  AND U6053 ( .A(n1199), .B(n6396), .Z(n6395) );
  XOR U6054 ( .A(n6397), .B(n6398), .Z(n6389) );
  AND U6055 ( .A(n1203), .B(n6399), .Z(n6398) );
  XOR U6056 ( .A(n6400), .B(n6401), .Z(n6386) );
  AND U6057 ( .A(n1207), .B(n6399), .Z(n6401) );
  XNOR U6058 ( .A(n6402), .B(n6400), .Z(n6399) );
  IV U6059 ( .A(n6397), .Z(n6402) );
  XOR U6060 ( .A(n6403), .B(n6404), .Z(n6397) );
  AND U6061 ( .A(n1210), .B(n6396), .Z(n6404) );
  XNOR U6062 ( .A(n6394), .B(n6403), .Z(n6396) );
  XNOR U6063 ( .A(n6405), .B(n6406), .Z(n6394) );
  AND U6064 ( .A(n1214), .B(n6407), .Z(n6406) );
  XOR U6065 ( .A(p_input[1827]), .B(n6405), .Z(n6407) );
  XNOR U6066 ( .A(n6408), .B(n6409), .Z(n6405) );
  AND U6067 ( .A(n1218), .B(n6410), .Z(n6409) );
  XOR U6068 ( .A(n6411), .B(n6412), .Z(n6403) );
  AND U6069 ( .A(n1222), .B(n6413), .Z(n6412) );
  XOR U6070 ( .A(n6414), .B(n6415), .Z(n6400) );
  AND U6071 ( .A(n1226), .B(n6413), .Z(n6415) );
  XNOR U6072 ( .A(n6416), .B(n6414), .Z(n6413) );
  IV U6073 ( .A(n6411), .Z(n6416) );
  XOR U6074 ( .A(n6417), .B(n6418), .Z(n6411) );
  AND U6075 ( .A(n1229), .B(n6410), .Z(n6418) );
  XNOR U6076 ( .A(n6408), .B(n6417), .Z(n6410) );
  XNOR U6077 ( .A(n6419), .B(n6420), .Z(n6408) );
  AND U6078 ( .A(n1233), .B(n6421), .Z(n6420) );
  XOR U6079 ( .A(p_input[1859]), .B(n6419), .Z(n6421) );
  XNOR U6080 ( .A(n6422), .B(n6423), .Z(n6419) );
  AND U6081 ( .A(n1237), .B(n6424), .Z(n6423) );
  XOR U6082 ( .A(n6425), .B(n6426), .Z(n6417) );
  AND U6083 ( .A(n1241), .B(n6427), .Z(n6426) );
  XOR U6084 ( .A(n6428), .B(n6429), .Z(n6414) );
  AND U6085 ( .A(n1245), .B(n6427), .Z(n6429) );
  XNOR U6086 ( .A(n6430), .B(n6428), .Z(n6427) );
  IV U6087 ( .A(n6425), .Z(n6430) );
  XOR U6088 ( .A(n6431), .B(n6432), .Z(n6425) );
  AND U6089 ( .A(n1248), .B(n6424), .Z(n6432) );
  XNOR U6090 ( .A(n6422), .B(n6431), .Z(n6424) );
  XNOR U6091 ( .A(n6433), .B(n6434), .Z(n6422) );
  AND U6092 ( .A(n1252), .B(n6435), .Z(n6434) );
  XOR U6093 ( .A(p_input[1891]), .B(n6433), .Z(n6435) );
  XNOR U6094 ( .A(n6436), .B(n6437), .Z(n6433) );
  AND U6095 ( .A(n1256), .B(n6438), .Z(n6437) );
  XOR U6096 ( .A(n6439), .B(n6440), .Z(n6431) );
  AND U6097 ( .A(n1260), .B(n6441), .Z(n6440) );
  XOR U6098 ( .A(n6442), .B(n6443), .Z(n6428) );
  AND U6099 ( .A(n1264), .B(n6441), .Z(n6443) );
  XNOR U6100 ( .A(n6444), .B(n6442), .Z(n6441) );
  IV U6101 ( .A(n6439), .Z(n6444) );
  XOR U6102 ( .A(n6445), .B(n6446), .Z(n6439) );
  AND U6103 ( .A(n1267), .B(n6438), .Z(n6446) );
  XNOR U6104 ( .A(n6436), .B(n6445), .Z(n6438) );
  XNOR U6105 ( .A(n6447), .B(n6448), .Z(n6436) );
  AND U6106 ( .A(n1271), .B(n6449), .Z(n6448) );
  XOR U6107 ( .A(p_input[1923]), .B(n6447), .Z(n6449) );
  XOR U6108 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(n6450), 
        .Z(n6447) );
  AND U6109 ( .A(n1274), .B(n6451), .Z(n6450) );
  XOR U6110 ( .A(n6452), .B(n6453), .Z(n6445) );
  AND U6111 ( .A(n1278), .B(n6454), .Z(n6453) );
  XOR U6112 ( .A(n6455), .B(n6456), .Z(n6442) );
  AND U6113 ( .A(n1282), .B(n6454), .Z(n6456) );
  XNOR U6114 ( .A(n6457), .B(n6455), .Z(n6454) );
  IV U6115 ( .A(n6452), .Z(n6457) );
  XOR U6116 ( .A(n6458), .B(n6459), .Z(n6452) );
  AND U6117 ( .A(n1285), .B(n6451), .Z(n6459) );
  XOR U6118 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(n6458), 
        .Z(n6451) );
  XOR U6119 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .B(n6460), 
        .Z(n6458) );
  AND U6120 ( .A(n1287), .B(n6461), .Z(n6460) );
  XOR U6121 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n6462), .Z(n6455) );
  AND U6122 ( .A(n1290), .B(n6461), .Z(n6462) );
  XOR U6123 ( .A(\knn_comb_/min_val_out[0][3] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .Z(n6461) );
  XOR U6124 ( .A(n6463), .B(n6464), .Z(o[34]) );
  XOR U6125 ( .A(n6465), .B(n6466), .Z(o[33]) );
  XOR U6126 ( .A(n6467), .B(n6468), .Z(o[32]) );
  XOR U6127 ( .A(n73), .B(n6469), .Z(o[31]) );
  AND U6128 ( .A(n122), .B(n6470), .Z(n73) );
  XOR U6129 ( .A(n74), .B(n6469), .Z(n6470) );
  XOR U6130 ( .A(n6471), .B(n6472), .Z(n6469) );
  AND U6131 ( .A(n142), .B(n6473), .Z(n6472) );
  XOR U6132 ( .A(n6474), .B(n3), .Z(n74) );
  AND U6133 ( .A(n125), .B(n6475), .Z(n3) );
  XOR U6134 ( .A(n4), .B(n6474), .Z(n6475) );
  XOR U6135 ( .A(n6476), .B(n6477), .Z(n4) );
  AND U6136 ( .A(n130), .B(n6478), .Z(n6477) );
  XOR U6137 ( .A(p_input[31]), .B(n6476), .Z(n6478) );
  XNOR U6138 ( .A(n6479), .B(n6480), .Z(n6476) );
  AND U6139 ( .A(n134), .B(n6481), .Z(n6480) );
  XOR U6140 ( .A(n6482), .B(n6483), .Z(n6474) );
  AND U6141 ( .A(n138), .B(n6473), .Z(n6483) );
  XNOR U6142 ( .A(n6484), .B(n6471), .Z(n6473) );
  XOR U6143 ( .A(n6485), .B(n6486), .Z(n6471) );
  AND U6144 ( .A(n162), .B(n6487), .Z(n6486) );
  IV U6145 ( .A(n6482), .Z(n6484) );
  XOR U6146 ( .A(n6488), .B(n6489), .Z(n6482) );
  AND U6147 ( .A(n146), .B(n6481), .Z(n6489) );
  XNOR U6148 ( .A(n6479), .B(n6488), .Z(n6481) );
  XNOR U6149 ( .A(n6490), .B(n6491), .Z(n6479) );
  AND U6150 ( .A(n150), .B(n6492), .Z(n6491) );
  XOR U6151 ( .A(p_input[63]), .B(n6490), .Z(n6492) );
  XNOR U6152 ( .A(n6493), .B(n6494), .Z(n6490) );
  AND U6153 ( .A(n154), .B(n6495), .Z(n6494) );
  XOR U6154 ( .A(n6496), .B(n6497), .Z(n6488) );
  AND U6155 ( .A(n158), .B(n6487), .Z(n6497) );
  XNOR U6156 ( .A(n6498), .B(n6485), .Z(n6487) );
  XOR U6157 ( .A(n6499), .B(n6500), .Z(n6485) );
  AND U6158 ( .A(n181), .B(n6501), .Z(n6500) );
  IV U6159 ( .A(n6496), .Z(n6498) );
  XOR U6160 ( .A(n6502), .B(n6503), .Z(n6496) );
  AND U6161 ( .A(n165), .B(n6495), .Z(n6503) );
  XNOR U6162 ( .A(n6493), .B(n6502), .Z(n6495) );
  XNOR U6163 ( .A(n6504), .B(n6505), .Z(n6493) );
  AND U6164 ( .A(n169), .B(n6506), .Z(n6505) );
  XOR U6165 ( .A(p_input[95]), .B(n6504), .Z(n6506) );
  XNOR U6166 ( .A(n6507), .B(n6508), .Z(n6504) );
  AND U6167 ( .A(n173), .B(n6509), .Z(n6508) );
  XOR U6168 ( .A(n6510), .B(n6511), .Z(n6502) );
  AND U6169 ( .A(n177), .B(n6501), .Z(n6511) );
  XNOR U6170 ( .A(n6512), .B(n6499), .Z(n6501) );
  XOR U6171 ( .A(n6513), .B(n6514), .Z(n6499) );
  AND U6172 ( .A(n200), .B(n6515), .Z(n6514) );
  IV U6173 ( .A(n6510), .Z(n6512) );
  XOR U6174 ( .A(n6516), .B(n6517), .Z(n6510) );
  AND U6175 ( .A(n184), .B(n6509), .Z(n6517) );
  XNOR U6176 ( .A(n6507), .B(n6516), .Z(n6509) );
  XNOR U6177 ( .A(n6518), .B(n6519), .Z(n6507) );
  AND U6178 ( .A(n188), .B(n6520), .Z(n6519) );
  XOR U6179 ( .A(p_input[127]), .B(n6518), .Z(n6520) );
  XNOR U6180 ( .A(n6521), .B(n6522), .Z(n6518) );
  AND U6181 ( .A(n192), .B(n6523), .Z(n6522) );
  XOR U6182 ( .A(n6524), .B(n6525), .Z(n6516) );
  AND U6183 ( .A(n196), .B(n6515), .Z(n6525) );
  XNOR U6184 ( .A(n6526), .B(n6513), .Z(n6515) );
  XOR U6185 ( .A(n6527), .B(n6528), .Z(n6513) );
  AND U6186 ( .A(n219), .B(n6529), .Z(n6528) );
  IV U6187 ( .A(n6524), .Z(n6526) );
  XOR U6188 ( .A(n6530), .B(n6531), .Z(n6524) );
  AND U6189 ( .A(n203), .B(n6523), .Z(n6531) );
  XNOR U6190 ( .A(n6521), .B(n6530), .Z(n6523) );
  XNOR U6191 ( .A(n6532), .B(n6533), .Z(n6521) );
  AND U6192 ( .A(n207), .B(n6534), .Z(n6533) );
  XOR U6193 ( .A(p_input[159]), .B(n6532), .Z(n6534) );
  XNOR U6194 ( .A(n6535), .B(n6536), .Z(n6532) );
  AND U6195 ( .A(n211), .B(n6537), .Z(n6536) );
  XOR U6196 ( .A(n6538), .B(n6539), .Z(n6530) );
  AND U6197 ( .A(n215), .B(n6529), .Z(n6539) );
  XNOR U6198 ( .A(n6540), .B(n6527), .Z(n6529) );
  XOR U6199 ( .A(n6541), .B(n6542), .Z(n6527) );
  AND U6200 ( .A(n238), .B(n6543), .Z(n6542) );
  IV U6201 ( .A(n6538), .Z(n6540) );
  XOR U6202 ( .A(n6544), .B(n6545), .Z(n6538) );
  AND U6203 ( .A(n222), .B(n6537), .Z(n6545) );
  XNOR U6204 ( .A(n6535), .B(n6544), .Z(n6537) );
  XNOR U6205 ( .A(n6546), .B(n6547), .Z(n6535) );
  AND U6206 ( .A(n226), .B(n6548), .Z(n6547) );
  XOR U6207 ( .A(p_input[191]), .B(n6546), .Z(n6548) );
  XNOR U6208 ( .A(n6549), .B(n6550), .Z(n6546) );
  AND U6209 ( .A(n230), .B(n6551), .Z(n6550) );
  XOR U6210 ( .A(n6552), .B(n6553), .Z(n6544) );
  AND U6211 ( .A(n234), .B(n6543), .Z(n6553) );
  XNOR U6212 ( .A(n6554), .B(n6541), .Z(n6543) );
  XOR U6213 ( .A(n6555), .B(n6556), .Z(n6541) );
  AND U6214 ( .A(n257), .B(n6557), .Z(n6556) );
  IV U6215 ( .A(n6552), .Z(n6554) );
  XOR U6216 ( .A(n6558), .B(n6559), .Z(n6552) );
  AND U6217 ( .A(n241), .B(n6551), .Z(n6559) );
  XNOR U6218 ( .A(n6549), .B(n6558), .Z(n6551) );
  XNOR U6219 ( .A(n6560), .B(n6561), .Z(n6549) );
  AND U6220 ( .A(n245), .B(n6562), .Z(n6561) );
  XOR U6221 ( .A(p_input[223]), .B(n6560), .Z(n6562) );
  XNOR U6222 ( .A(n6563), .B(n6564), .Z(n6560) );
  AND U6223 ( .A(n249), .B(n6565), .Z(n6564) );
  XOR U6224 ( .A(n6566), .B(n6567), .Z(n6558) );
  AND U6225 ( .A(n253), .B(n6557), .Z(n6567) );
  XNOR U6226 ( .A(n6568), .B(n6555), .Z(n6557) );
  XOR U6227 ( .A(n6569), .B(n6570), .Z(n6555) );
  AND U6228 ( .A(n276), .B(n6571), .Z(n6570) );
  IV U6229 ( .A(n6566), .Z(n6568) );
  XOR U6230 ( .A(n6572), .B(n6573), .Z(n6566) );
  AND U6231 ( .A(n260), .B(n6565), .Z(n6573) );
  XNOR U6232 ( .A(n6563), .B(n6572), .Z(n6565) );
  XNOR U6233 ( .A(n6574), .B(n6575), .Z(n6563) );
  AND U6234 ( .A(n264), .B(n6576), .Z(n6575) );
  XOR U6235 ( .A(p_input[255]), .B(n6574), .Z(n6576) );
  XNOR U6236 ( .A(n6577), .B(n6578), .Z(n6574) );
  AND U6237 ( .A(n268), .B(n6579), .Z(n6578) );
  XOR U6238 ( .A(n6580), .B(n6581), .Z(n6572) );
  AND U6239 ( .A(n272), .B(n6571), .Z(n6581) );
  XNOR U6240 ( .A(n6582), .B(n6569), .Z(n6571) );
  XOR U6241 ( .A(n6583), .B(n6584), .Z(n6569) );
  AND U6242 ( .A(n295), .B(n6585), .Z(n6584) );
  IV U6243 ( .A(n6580), .Z(n6582) );
  XOR U6244 ( .A(n6586), .B(n6587), .Z(n6580) );
  AND U6245 ( .A(n279), .B(n6579), .Z(n6587) );
  XNOR U6246 ( .A(n6577), .B(n6586), .Z(n6579) );
  XNOR U6247 ( .A(n6588), .B(n6589), .Z(n6577) );
  AND U6248 ( .A(n283), .B(n6590), .Z(n6589) );
  XOR U6249 ( .A(p_input[287]), .B(n6588), .Z(n6590) );
  XNOR U6250 ( .A(n6591), .B(n6592), .Z(n6588) );
  AND U6251 ( .A(n287), .B(n6593), .Z(n6592) );
  XOR U6252 ( .A(n6594), .B(n6595), .Z(n6586) );
  AND U6253 ( .A(n291), .B(n6585), .Z(n6595) );
  XNOR U6254 ( .A(n6596), .B(n6583), .Z(n6585) );
  XOR U6255 ( .A(n6597), .B(n6598), .Z(n6583) );
  AND U6256 ( .A(n314), .B(n6599), .Z(n6598) );
  IV U6257 ( .A(n6594), .Z(n6596) );
  XOR U6258 ( .A(n6600), .B(n6601), .Z(n6594) );
  AND U6259 ( .A(n298), .B(n6593), .Z(n6601) );
  XNOR U6260 ( .A(n6591), .B(n6600), .Z(n6593) );
  XNOR U6261 ( .A(n6602), .B(n6603), .Z(n6591) );
  AND U6262 ( .A(n302), .B(n6604), .Z(n6603) );
  XOR U6263 ( .A(p_input[319]), .B(n6602), .Z(n6604) );
  XNOR U6264 ( .A(n6605), .B(n6606), .Z(n6602) );
  AND U6265 ( .A(n306), .B(n6607), .Z(n6606) );
  XOR U6266 ( .A(n6608), .B(n6609), .Z(n6600) );
  AND U6267 ( .A(n310), .B(n6599), .Z(n6609) );
  XNOR U6268 ( .A(n6610), .B(n6597), .Z(n6599) );
  XOR U6269 ( .A(n6611), .B(n6612), .Z(n6597) );
  AND U6270 ( .A(n333), .B(n6613), .Z(n6612) );
  IV U6271 ( .A(n6608), .Z(n6610) );
  XOR U6272 ( .A(n6614), .B(n6615), .Z(n6608) );
  AND U6273 ( .A(n317), .B(n6607), .Z(n6615) );
  XNOR U6274 ( .A(n6605), .B(n6614), .Z(n6607) );
  XNOR U6275 ( .A(n6616), .B(n6617), .Z(n6605) );
  AND U6276 ( .A(n321), .B(n6618), .Z(n6617) );
  XOR U6277 ( .A(p_input[351]), .B(n6616), .Z(n6618) );
  XNOR U6278 ( .A(n6619), .B(n6620), .Z(n6616) );
  AND U6279 ( .A(n325), .B(n6621), .Z(n6620) );
  XOR U6280 ( .A(n6622), .B(n6623), .Z(n6614) );
  AND U6281 ( .A(n329), .B(n6613), .Z(n6623) );
  XNOR U6282 ( .A(n6624), .B(n6611), .Z(n6613) );
  XOR U6283 ( .A(n6625), .B(n6626), .Z(n6611) );
  AND U6284 ( .A(n352), .B(n6627), .Z(n6626) );
  IV U6285 ( .A(n6622), .Z(n6624) );
  XOR U6286 ( .A(n6628), .B(n6629), .Z(n6622) );
  AND U6287 ( .A(n336), .B(n6621), .Z(n6629) );
  XNOR U6288 ( .A(n6619), .B(n6628), .Z(n6621) );
  XNOR U6289 ( .A(n6630), .B(n6631), .Z(n6619) );
  AND U6290 ( .A(n340), .B(n6632), .Z(n6631) );
  XOR U6291 ( .A(p_input[383]), .B(n6630), .Z(n6632) );
  XNOR U6292 ( .A(n6633), .B(n6634), .Z(n6630) );
  AND U6293 ( .A(n344), .B(n6635), .Z(n6634) );
  XOR U6294 ( .A(n6636), .B(n6637), .Z(n6628) );
  AND U6295 ( .A(n348), .B(n6627), .Z(n6637) );
  XNOR U6296 ( .A(n6638), .B(n6625), .Z(n6627) );
  XOR U6297 ( .A(n6639), .B(n6640), .Z(n6625) );
  AND U6298 ( .A(n371), .B(n6641), .Z(n6640) );
  IV U6299 ( .A(n6636), .Z(n6638) );
  XOR U6300 ( .A(n6642), .B(n6643), .Z(n6636) );
  AND U6301 ( .A(n355), .B(n6635), .Z(n6643) );
  XNOR U6302 ( .A(n6633), .B(n6642), .Z(n6635) );
  XNOR U6303 ( .A(n6644), .B(n6645), .Z(n6633) );
  AND U6304 ( .A(n359), .B(n6646), .Z(n6645) );
  XOR U6305 ( .A(p_input[415]), .B(n6644), .Z(n6646) );
  XNOR U6306 ( .A(n6647), .B(n6648), .Z(n6644) );
  AND U6307 ( .A(n363), .B(n6649), .Z(n6648) );
  XOR U6308 ( .A(n6650), .B(n6651), .Z(n6642) );
  AND U6309 ( .A(n367), .B(n6641), .Z(n6651) );
  XNOR U6310 ( .A(n6652), .B(n6639), .Z(n6641) );
  XOR U6311 ( .A(n6653), .B(n6654), .Z(n6639) );
  AND U6312 ( .A(n390), .B(n6655), .Z(n6654) );
  IV U6313 ( .A(n6650), .Z(n6652) );
  XOR U6314 ( .A(n6656), .B(n6657), .Z(n6650) );
  AND U6315 ( .A(n374), .B(n6649), .Z(n6657) );
  XNOR U6316 ( .A(n6647), .B(n6656), .Z(n6649) );
  XNOR U6317 ( .A(n6658), .B(n6659), .Z(n6647) );
  AND U6318 ( .A(n378), .B(n6660), .Z(n6659) );
  XOR U6319 ( .A(p_input[447]), .B(n6658), .Z(n6660) );
  XNOR U6320 ( .A(n6661), .B(n6662), .Z(n6658) );
  AND U6321 ( .A(n382), .B(n6663), .Z(n6662) );
  XOR U6322 ( .A(n6664), .B(n6665), .Z(n6656) );
  AND U6323 ( .A(n386), .B(n6655), .Z(n6665) );
  XNOR U6324 ( .A(n6666), .B(n6653), .Z(n6655) );
  XOR U6325 ( .A(n6667), .B(n6668), .Z(n6653) );
  AND U6326 ( .A(n409), .B(n6669), .Z(n6668) );
  IV U6327 ( .A(n6664), .Z(n6666) );
  XOR U6328 ( .A(n6670), .B(n6671), .Z(n6664) );
  AND U6329 ( .A(n393), .B(n6663), .Z(n6671) );
  XNOR U6330 ( .A(n6661), .B(n6670), .Z(n6663) );
  XNOR U6331 ( .A(n6672), .B(n6673), .Z(n6661) );
  AND U6332 ( .A(n397), .B(n6674), .Z(n6673) );
  XOR U6333 ( .A(p_input[479]), .B(n6672), .Z(n6674) );
  XNOR U6334 ( .A(n6675), .B(n6676), .Z(n6672) );
  AND U6335 ( .A(n401), .B(n6677), .Z(n6676) );
  XOR U6336 ( .A(n6678), .B(n6679), .Z(n6670) );
  AND U6337 ( .A(n405), .B(n6669), .Z(n6679) );
  XNOR U6338 ( .A(n6680), .B(n6667), .Z(n6669) );
  XOR U6339 ( .A(n6681), .B(n6682), .Z(n6667) );
  AND U6340 ( .A(n428), .B(n6683), .Z(n6682) );
  IV U6341 ( .A(n6678), .Z(n6680) );
  XOR U6342 ( .A(n6684), .B(n6685), .Z(n6678) );
  AND U6343 ( .A(n412), .B(n6677), .Z(n6685) );
  XNOR U6344 ( .A(n6675), .B(n6684), .Z(n6677) );
  XNOR U6345 ( .A(n6686), .B(n6687), .Z(n6675) );
  AND U6346 ( .A(n416), .B(n6688), .Z(n6687) );
  XOR U6347 ( .A(p_input[511]), .B(n6686), .Z(n6688) );
  XNOR U6348 ( .A(n6689), .B(n6690), .Z(n6686) );
  AND U6349 ( .A(n420), .B(n6691), .Z(n6690) );
  XOR U6350 ( .A(n6692), .B(n6693), .Z(n6684) );
  AND U6351 ( .A(n424), .B(n6683), .Z(n6693) );
  XNOR U6352 ( .A(n6694), .B(n6681), .Z(n6683) );
  XOR U6353 ( .A(n6695), .B(n6696), .Z(n6681) );
  AND U6354 ( .A(n447), .B(n6697), .Z(n6696) );
  IV U6355 ( .A(n6692), .Z(n6694) );
  XOR U6356 ( .A(n6698), .B(n6699), .Z(n6692) );
  AND U6357 ( .A(n431), .B(n6691), .Z(n6699) );
  XNOR U6358 ( .A(n6689), .B(n6698), .Z(n6691) );
  XNOR U6359 ( .A(n6700), .B(n6701), .Z(n6689) );
  AND U6360 ( .A(n435), .B(n6702), .Z(n6701) );
  XOR U6361 ( .A(p_input[543]), .B(n6700), .Z(n6702) );
  XNOR U6362 ( .A(n6703), .B(n6704), .Z(n6700) );
  AND U6363 ( .A(n439), .B(n6705), .Z(n6704) );
  XOR U6364 ( .A(n6706), .B(n6707), .Z(n6698) );
  AND U6365 ( .A(n443), .B(n6697), .Z(n6707) );
  XNOR U6366 ( .A(n6708), .B(n6695), .Z(n6697) );
  XOR U6367 ( .A(n6709), .B(n6710), .Z(n6695) );
  AND U6368 ( .A(n466), .B(n6711), .Z(n6710) );
  IV U6369 ( .A(n6706), .Z(n6708) );
  XOR U6370 ( .A(n6712), .B(n6713), .Z(n6706) );
  AND U6371 ( .A(n450), .B(n6705), .Z(n6713) );
  XNOR U6372 ( .A(n6703), .B(n6712), .Z(n6705) );
  XNOR U6373 ( .A(n6714), .B(n6715), .Z(n6703) );
  AND U6374 ( .A(n454), .B(n6716), .Z(n6715) );
  XOR U6375 ( .A(p_input[575]), .B(n6714), .Z(n6716) );
  XNOR U6376 ( .A(n6717), .B(n6718), .Z(n6714) );
  AND U6377 ( .A(n458), .B(n6719), .Z(n6718) );
  XOR U6378 ( .A(n6720), .B(n6721), .Z(n6712) );
  AND U6379 ( .A(n462), .B(n6711), .Z(n6721) );
  XNOR U6380 ( .A(n6722), .B(n6709), .Z(n6711) );
  XOR U6381 ( .A(n6723), .B(n6724), .Z(n6709) );
  AND U6382 ( .A(n485), .B(n6725), .Z(n6724) );
  IV U6383 ( .A(n6720), .Z(n6722) );
  XOR U6384 ( .A(n6726), .B(n6727), .Z(n6720) );
  AND U6385 ( .A(n469), .B(n6719), .Z(n6727) );
  XNOR U6386 ( .A(n6717), .B(n6726), .Z(n6719) );
  XNOR U6387 ( .A(n6728), .B(n6729), .Z(n6717) );
  AND U6388 ( .A(n473), .B(n6730), .Z(n6729) );
  XOR U6389 ( .A(p_input[607]), .B(n6728), .Z(n6730) );
  XNOR U6390 ( .A(n6731), .B(n6732), .Z(n6728) );
  AND U6391 ( .A(n477), .B(n6733), .Z(n6732) );
  XOR U6392 ( .A(n6734), .B(n6735), .Z(n6726) );
  AND U6393 ( .A(n481), .B(n6725), .Z(n6735) );
  XNOR U6394 ( .A(n6736), .B(n6723), .Z(n6725) );
  XOR U6395 ( .A(n6737), .B(n6738), .Z(n6723) );
  AND U6396 ( .A(n504), .B(n6739), .Z(n6738) );
  IV U6397 ( .A(n6734), .Z(n6736) );
  XOR U6398 ( .A(n6740), .B(n6741), .Z(n6734) );
  AND U6399 ( .A(n488), .B(n6733), .Z(n6741) );
  XNOR U6400 ( .A(n6731), .B(n6740), .Z(n6733) );
  XNOR U6401 ( .A(n6742), .B(n6743), .Z(n6731) );
  AND U6402 ( .A(n492), .B(n6744), .Z(n6743) );
  XOR U6403 ( .A(p_input[639]), .B(n6742), .Z(n6744) );
  XNOR U6404 ( .A(n6745), .B(n6746), .Z(n6742) );
  AND U6405 ( .A(n496), .B(n6747), .Z(n6746) );
  XOR U6406 ( .A(n6748), .B(n6749), .Z(n6740) );
  AND U6407 ( .A(n500), .B(n6739), .Z(n6749) );
  XNOR U6408 ( .A(n6750), .B(n6737), .Z(n6739) );
  XOR U6409 ( .A(n6751), .B(n6752), .Z(n6737) );
  AND U6410 ( .A(n523), .B(n6753), .Z(n6752) );
  IV U6411 ( .A(n6748), .Z(n6750) );
  XOR U6412 ( .A(n6754), .B(n6755), .Z(n6748) );
  AND U6413 ( .A(n507), .B(n6747), .Z(n6755) );
  XNOR U6414 ( .A(n6745), .B(n6754), .Z(n6747) );
  XNOR U6415 ( .A(n6756), .B(n6757), .Z(n6745) );
  AND U6416 ( .A(n511), .B(n6758), .Z(n6757) );
  XOR U6417 ( .A(p_input[671]), .B(n6756), .Z(n6758) );
  XNOR U6418 ( .A(n6759), .B(n6760), .Z(n6756) );
  AND U6419 ( .A(n515), .B(n6761), .Z(n6760) );
  XOR U6420 ( .A(n6762), .B(n6763), .Z(n6754) );
  AND U6421 ( .A(n519), .B(n6753), .Z(n6763) );
  XNOR U6422 ( .A(n6764), .B(n6751), .Z(n6753) );
  XOR U6423 ( .A(n6765), .B(n6766), .Z(n6751) );
  AND U6424 ( .A(n542), .B(n6767), .Z(n6766) );
  IV U6425 ( .A(n6762), .Z(n6764) );
  XOR U6426 ( .A(n6768), .B(n6769), .Z(n6762) );
  AND U6427 ( .A(n526), .B(n6761), .Z(n6769) );
  XNOR U6428 ( .A(n6759), .B(n6768), .Z(n6761) );
  XNOR U6429 ( .A(n6770), .B(n6771), .Z(n6759) );
  AND U6430 ( .A(n530), .B(n6772), .Z(n6771) );
  XOR U6431 ( .A(p_input[703]), .B(n6770), .Z(n6772) );
  XNOR U6432 ( .A(n6773), .B(n6774), .Z(n6770) );
  AND U6433 ( .A(n534), .B(n6775), .Z(n6774) );
  XOR U6434 ( .A(n6776), .B(n6777), .Z(n6768) );
  AND U6435 ( .A(n538), .B(n6767), .Z(n6777) );
  XNOR U6436 ( .A(n6778), .B(n6765), .Z(n6767) );
  XOR U6437 ( .A(n6779), .B(n6780), .Z(n6765) );
  AND U6438 ( .A(n561), .B(n6781), .Z(n6780) );
  IV U6439 ( .A(n6776), .Z(n6778) );
  XOR U6440 ( .A(n6782), .B(n6783), .Z(n6776) );
  AND U6441 ( .A(n545), .B(n6775), .Z(n6783) );
  XNOR U6442 ( .A(n6773), .B(n6782), .Z(n6775) );
  XNOR U6443 ( .A(n6784), .B(n6785), .Z(n6773) );
  AND U6444 ( .A(n549), .B(n6786), .Z(n6785) );
  XOR U6445 ( .A(p_input[735]), .B(n6784), .Z(n6786) );
  XNOR U6446 ( .A(n6787), .B(n6788), .Z(n6784) );
  AND U6447 ( .A(n553), .B(n6789), .Z(n6788) );
  XOR U6448 ( .A(n6790), .B(n6791), .Z(n6782) );
  AND U6449 ( .A(n557), .B(n6781), .Z(n6791) );
  XNOR U6450 ( .A(n6792), .B(n6779), .Z(n6781) );
  XOR U6451 ( .A(n6793), .B(n6794), .Z(n6779) );
  AND U6452 ( .A(n580), .B(n6795), .Z(n6794) );
  IV U6453 ( .A(n6790), .Z(n6792) );
  XOR U6454 ( .A(n6796), .B(n6797), .Z(n6790) );
  AND U6455 ( .A(n564), .B(n6789), .Z(n6797) );
  XNOR U6456 ( .A(n6787), .B(n6796), .Z(n6789) );
  XNOR U6457 ( .A(n6798), .B(n6799), .Z(n6787) );
  AND U6458 ( .A(n568), .B(n6800), .Z(n6799) );
  XOR U6459 ( .A(p_input[767]), .B(n6798), .Z(n6800) );
  XNOR U6460 ( .A(n6801), .B(n6802), .Z(n6798) );
  AND U6461 ( .A(n572), .B(n6803), .Z(n6802) );
  XOR U6462 ( .A(n6804), .B(n6805), .Z(n6796) );
  AND U6463 ( .A(n576), .B(n6795), .Z(n6805) );
  XNOR U6464 ( .A(n6806), .B(n6793), .Z(n6795) );
  XOR U6465 ( .A(n6807), .B(n6808), .Z(n6793) );
  AND U6466 ( .A(n599), .B(n6809), .Z(n6808) );
  IV U6467 ( .A(n6804), .Z(n6806) );
  XOR U6468 ( .A(n6810), .B(n6811), .Z(n6804) );
  AND U6469 ( .A(n583), .B(n6803), .Z(n6811) );
  XNOR U6470 ( .A(n6801), .B(n6810), .Z(n6803) );
  XNOR U6471 ( .A(n6812), .B(n6813), .Z(n6801) );
  AND U6472 ( .A(n587), .B(n6814), .Z(n6813) );
  XOR U6473 ( .A(p_input[799]), .B(n6812), .Z(n6814) );
  XNOR U6474 ( .A(n6815), .B(n6816), .Z(n6812) );
  AND U6475 ( .A(n591), .B(n6817), .Z(n6816) );
  XOR U6476 ( .A(n6818), .B(n6819), .Z(n6810) );
  AND U6477 ( .A(n595), .B(n6809), .Z(n6819) );
  XNOR U6478 ( .A(n6820), .B(n6807), .Z(n6809) );
  XOR U6479 ( .A(n6821), .B(n6822), .Z(n6807) );
  AND U6480 ( .A(n618), .B(n6823), .Z(n6822) );
  IV U6481 ( .A(n6818), .Z(n6820) );
  XOR U6482 ( .A(n6824), .B(n6825), .Z(n6818) );
  AND U6483 ( .A(n602), .B(n6817), .Z(n6825) );
  XNOR U6484 ( .A(n6815), .B(n6824), .Z(n6817) );
  XNOR U6485 ( .A(n6826), .B(n6827), .Z(n6815) );
  AND U6486 ( .A(n606), .B(n6828), .Z(n6827) );
  XOR U6487 ( .A(p_input[831]), .B(n6826), .Z(n6828) );
  XNOR U6488 ( .A(n6829), .B(n6830), .Z(n6826) );
  AND U6489 ( .A(n610), .B(n6831), .Z(n6830) );
  XOR U6490 ( .A(n6832), .B(n6833), .Z(n6824) );
  AND U6491 ( .A(n614), .B(n6823), .Z(n6833) );
  XNOR U6492 ( .A(n6834), .B(n6821), .Z(n6823) );
  XOR U6493 ( .A(n6835), .B(n6836), .Z(n6821) );
  AND U6494 ( .A(n637), .B(n6837), .Z(n6836) );
  IV U6495 ( .A(n6832), .Z(n6834) );
  XOR U6496 ( .A(n6838), .B(n6839), .Z(n6832) );
  AND U6497 ( .A(n621), .B(n6831), .Z(n6839) );
  XNOR U6498 ( .A(n6829), .B(n6838), .Z(n6831) );
  XNOR U6499 ( .A(n6840), .B(n6841), .Z(n6829) );
  AND U6500 ( .A(n625), .B(n6842), .Z(n6841) );
  XOR U6501 ( .A(p_input[863]), .B(n6840), .Z(n6842) );
  XNOR U6502 ( .A(n6843), .B(n6844), .Z(n6840) );
  AND U6503 ( .A(n629), .B(n6845), .Z(n6844) );
  XOR U6504 ( .A(n6846), .B(n6847), .Z(n6838) );
  AND U6505 ( .A(n633), .B(n6837), .Z(n6847) );
  XNOR U6506 ( .A(n6848), .B(n6835), .Z(n6837) );
  XOR U6507 ( .A(n6849), .B(n6850), .Z(n6835) );
  AND U6508 ( .A(n656), .B(n6851), .Z(n6850) );
  IV U6509 ( .A(n6846), .Z(n6848) );
  XOR U6510 ( .A(n6852), .B(n6853), .Z(n6846) );
  AND U6511 ( .A(n640), .B(n6845), .Z(n6853) );
  XNOR U6512 ( .A(n6843), .B(n6852), .Z(n6845) );
  XNOR U6513 ( .A(n6854), .B(n6855), .Z(n6843) );
  AND U6514 ( .A(n644), .B(n6856), .Z(n6855) );
  XOR U6515 ( .A(p_input[895]), .B(n6854), .Z(n6856) );
  XNOR U6516 ( .A(n6857), .B(n6858), .Z(n6854) );
  AND U6517 ( .A(n648), .B(n6859), .Z(n6858) );
  XOR U6518 ( .A(n6860), .B(n6861), .Z(n6852) );
  AND U6519 ( .A(n652), .B(n6851), .Z(n6861) );
  XNOR U6520 ( .A(n6862), .B(n6849), .Z(n6851) );
  XOR U6521 ( .A(n6863), .B(n6864), .Z(n6849) );
  AND U6522 ( .A(n675), .B(n6865), .Z(n6864) );
  IV U6523 ( .A(n6860), .Z(n6862) );
  XOR U6524 ( .A(n6866), .B(n6867), .Z(n6860) );
  AND U6525 ( .A(n659), .B(n6859), .Z(n6867) );
  XNOR U6526 ( .A(n6857), .B(n6866), .Z(n6859) );
  XNOR U6527 ( .A(n6868), .B(n6869), .Z(n6857) );
  AND U6528 ( .A(n663), .B(n6870), .Z(n6869) );
  XOR U6529 ( .A(p_input[927]), .B(n6868), .Z(n6870) );
  XNOR U6530 ( .A(n6871), .B(n6872), .Z(n6868) );
  AND U6531 ( .A(n667), .B(n6873), .Z(n6872) );
  XOR U6532 ( .A(n6874), .B(n6875), .Z(n6866) );
  AND U6533 ( .A(n671), .B(n6865), .Z(n6875) );
  XNOR U6534 ( .A(n6876), .B(n6863), .Z(n6865) );
  XOR U6535 ( .A(n6877), .B(n6878), .Z(n6863) );
  AND U6536 ( .A(n694), .B(n6879), .Z(n6878) );
  IV U6537 ( .A(n6874), .Z(n6876) );
  XOR U6538 ( .A(n6880), .B(n6881), .Z(n6874) );
  AND U6539 ( .A(n678), .B(n6873), .Z(n6881) );
  XNOR U6540 ( .A(n6871), .B(n6880), .Z(n6873) );
  XNOR U6541 ( .A(n6882), .B(n6883), .Z(n6871) );
  AND U6542 ( .A(n682), .B(n6884), .Z(n6883) );
  XOR U6543 ( .A(p_input[959]), .B(n6882), .Z(n6884) );
  XNOR U6544 ( .A(n6885), .B(n6886), .Z(n6882) );
  AND U6545 ( .A(n686), .B(n6887), .Z(n6886) );
  XOR U6546 ( .A(n6888), .B(n6889), .Z(n6880) );
  AND U6547 ( .A(n690), .B(n6879), .Z(n6889) );
  XNOR U6548 ( .A(n6890), .B(n6877), .Z(n6879) );
  XOR U6549 ( .A(n6891), .B(n6892), .Z(n6877) );
  AND U6550 ( .A(n713), .B(n6893), .Z(n6892) );
  IV U6551 ( .A(n6888), .Z(n6890) );
  XOR U6552 ( .A(n6894), .B(n6895), .Z(n6888) );
  AND U6553 ( .A(n697), .B(n6887), .Z(n6895) );
  XNOR U6554 ( .A(n6885), .B(n6894), .Z(n6887) );
  XNOR U6555 ( .A(n6896), .B(n6897), .Z(n6885) );
  AND U6556 ( .A(n701), .B(n6898), .Z(n6897) );
  XOR U6557 ( .A(p_input[991]), .B(n6896), .Z(n6898) );
  XNOR U6558 ( .A(n6899), .B(n6900), .Z(n6896) );
  AND U6559 ( .A(n705), .B(n6901), .Z(n6900) );
  XOR U6560 ( .A(n6902), .B(n6903), .Z(n6894) );
  AND U6561 ( .A(n709), .B(n6893), .Z(n6903) );
  XNOR U6562 ( .A(n6904), .B(n6891), .Z(n6893) );
  XOR U6563 ( .A(n6905), .B(n6906), .Z(n6891) );
  AND U6564 ( .A(n732), .B(n6907), .Z(n6906) );
  IV U6565 ( .A(n6902), .Z(n6904) );
  XOR U6566 ( .A(n6908), .B(n6909), .Z(n6902) );
  AND U6567 ( .A(n716), .B(n6901), .Z(n6909) );
  XNOR U6568 ( .A(n6899), .B(n6908), .Z(n6901) );
  XNOR U6569 ( .A(n6910), .B(n6911), .Z(n6899) );
  AND U6570 ( .A(n720), .B(n6912), .Z(n6911) );
  XOR U6571 ( .A(p_input[1023]), .B(n6910), .Z(n6912) );
  XNOR U6572 ( .A(n6913), .B(n6914), .Z(n6910) );
  AND U6573 ( .A(n724), .B(n6915), .Z(n6914) );
  XOR U6574 ( .A(n6916), .B(n6917), .Z(n6908) );
  AND U6575 ( .A(n728), .B(n6907), .Z(n6917) );
  XNOR U6576 ( .A(n6918), .B(n6905), .Z(n6907) );
  XOR U6577 ( .A(n6919), .B(n6920), .Z(n6905) );
  AND U6578 ( .A(n751), .B(n6921), .Z(n6920) );
  IV U6579 ( .A(n6916), .Z(n6918) );
  XOR U6580 ( .A(n6922), .B(n6923), .Z(n6916) );
  AND U6581 ( .A(n735), .B(n6915), .Z(n6923) );
  XNOR U6582 ( .A(n6913), .B(n6922), .Z(n6915) );
  XNOR U6583 ( .A(n6924), .B(n6925), .Z(n6913) );
  AND U6584 ( .A(n739), .B(n6926), .Z(n6925) );
  XOR U6585 ( .A(p_input[1055]), .B(n6924), .Z(n6926) );
  XNOR U6586 ( .A(n6927), .B(n6928), .Z(n6924) );
  AND U6587 ( .A(n743), .B(n6929), .Z(n6928) );
  XOR U6588 ( .A(n6930), .B(n6931), .Z(n6922) );
  AND U6589 ( .A(n747), .B(n6921), .Z(n6931) );
  XNOR U6590 ( .A(n6932), .B(n6919), .Z(n6921) );
  XOR U6591 ( .A(n6933), .B(n6934), .Z(n6919) );
  AND U6592 ( .A(n770), .B(n6935), .Z(n6934) );
  IV U6593 ( .A(n6930), .Z(n6932) );
  XOR U6594 ( .A(n6936), .B(n6937), .Z(n6930) );
  AND U6595 ( .A(n754), .B(n6929), .Z(n6937) );
  XNOR U6596 ( .A(n6927), .B(n6936), .Z(n6929) );
  XNOR U6597 ( .A(n6938), .B(n6939), .Z(n6927) );
  AND U6598 ( .A(n758), .B(n6940), .Z(n6939) );
  XOR U6599 ( .A(p_input[1087]), .B(n6938), .Z(n6940) );
  XNOR U6600 ( .A(n6941), .B(n6942), .Z(n6938) );
  AND U6601 ( .A(n762), .B(n6943), .Z(n6942) );
  XOR U6602 ( .A(n6944), .B(n6945), .Z(n6936) );
  AND U6603 ( .A(n766), .B(n6935), .Z(n6945) );
  XNOR U6604 ( .A(n6946), .B(n6933), .Z(n6935) );
  XOR U6605 ( .A(n6947), .B(n6948), .Z(n6933) );
  AND U6606 ( .A(n789), .B(n6949), .Z(n6948) );
  IV U6607 ( .A(n6944), .Z(n6946) );
  XOR U6608 ( .A(n6950), .B(n6951), .Z(n6944) );
  AND U6609 ( .A(n773), .B(n6943), .Z(n6951) );
  XNOR U6610 ( .A(n6941), .B(n6950), .Z(n6943) );
  XNOR U6611 ( .A(n6952), .B(n6953), .Z(n6941) );
  AND U6612 ( .A(n777), .B(n6954), .Z(n6953) );
  XOR U6613 ( .A(p_input[1119]), .B(n6952), .Z(n6954) );
  XNOR U6614 ( .A(n6955), .B(n6956), .Z(n6952) );
  AND U6615 ( .A(n781), .B(n6957), .Z(n6956) );
  XOR U6616 ( .A(n6958), .B(n6959), .Z(n6950) );
  AND U6617 ( .A(n785), .B(n6949), .Z(n6959) );
  XNOR U6618 ( .A(n6960), .B(n6947), .Z(n6949) );
  XOR U6619 ( .A(n6961), .B(n6962), .Z(n6947) );
  AND U6620 ( .A(n808), .B(n6963), .Z(n6962) );
  IV U6621 ( .A(n6958), .Z(n6960) );
  XOR U6622 ( .A(n6964), .B(n6965), .Z(n6958) );
  AND U6623 ( .A(n792), .B(n6957), .Z(n6965) );
  XNOR U6624 ( .A(n6955), .B(n6964), .Z(n6957) );
  XNOR U6625 ( .A(n6966), .B(n6967), .Z(n6955) );
  AND U6626 ( .A(n796), .B(n6968), .Z(n6967) );
  XOR U6627 ( .A(p_input[1151]), .B(n6966), .Z(n6968) );
  XNOR U6628 ( .A(n6969), .B(n6970), .Z(n6966) );
  AND U6629 ( .A(n800), .B(n6971), .Z(n6970) );
  XOR U6630 ( .A(n6972), .B(n6973), .Z(n6964) );
  AND U6631 ( .A(n804), .B(n6963), .Z(n6973) );
  XNOR U6632 ( .A(n6974), .B(n6961), .Z(n6963) );
  XOR U6633 ( .A(n6975), .B(n6976), .Z(n6961) );
  AND U6634 ( .A(n827), .B(n6977), .Z(n6976) );
  IV U6635 ( .A(n6972), .Z(n6974) );
  XOR U6636 ( .A(n6978), .B(n6979), .Z(n6972) );
  AND U6637 ( .A(n811), .B(n6971), .Z(n6979) );
  XNOR U6638 ( .A(n6969), .B(n6978), .Z(n6971) );
  XNOR U6639 ( .A(n6980), .B(n6981), .Z(n6969) );
  AND U6640 ( .A(n815), .B(n6982), .Z(n6981) );
  XOR U6641 ( .A(p_input[1183]), .B(n6980), .Z(n6982) );
  XNOR U6642 ( .A(n6983), .B(n6984), .Z(n6980) );
  AND U6643 ( .A(n819), .B(n6985), .Z(n6984) );
  XOR U6644 ( .A(n6986), .B(n6987), .Z(n6978) );
  AND U6645 ( .A(n823), .B(n6977), .Z(n6987) );
  XNOR U6646 ( .A(n6988), .B(n6975), .Z(n6977) );
  XOR U6647 ( .A(n6989), .B(n6990), .Z(n6975) );
  AND U6648 ( .A(n846), .B(n6991), .Z(n6990) );
  IV U6649 ( .A(n6986), .Z(n6988) );
  XOR U6650 ( .A(n6992), .B(n6993), .Z(n6986) );
  AND U6651 ( .A(n830), .B(n6985), .Z(n6993) );
  XNOR U6652 ( .A(n6983), .B(n6992), .Z(n6985) );
  XNOR U6653 ( .A(n6994), .B(n6995), .Z(n6983) );
  AND U6654 ( .A(n834), .B(n6996), .Z(n6995) );
  XOR U6655 ( .A(p_input[1215]), .B(n6994), .Z(n6996) );
  XNOR U6656 ( .A(n6997), .B(n6998), .Z(n6994) );
  AND U6657 ( .A(n838), .B(n6999), .Z(n6998) );
  XOR U6658 ( .A(n7000), .B(n7001), .Z(n6992) );
  AND U6659 ( .A(n842), .B(n6991), .Z(n7001) );
  XNOR U6660 ( .A(n7002), .B(n6989), .Z(n6991) );
  XOR U6661 ( .A(n7003), .B(n7004), .Z(n6989) );
  AND U6662 ( .A(n865), .B(n7005), .Z(n7004) );
  IV U6663 ( .A(n7000), .Z(n7002) );
  XOR U6664 ( .A(n7006), .B(n7007), .Z(n7000) );
  AND U6665 ( .A(n849), .B(n6999), .Z(n7007) );
  XNOR U6666 ( .A(n6997), .B(n7006), .Z(n6999) );
  XNOR U6667 ( .A(n7008), .B(n7009), .Z(n6997) );
  AND U6668 ( .A(n853), .B(n7010), .Z(n7009) );
  XOR U6669 ( .A(p_input[1247]), .B(n7008), .Z(n7010) );
  XNOR U6670 ( .A(n7011), .B(n7012), .Z(n7008) );
  AND U6671 ( .A(n857), .B(n7013), .Z(n7012) );
  XOR U6672 ( .A(n7014), .B(n7015), .Z(n7006) );
  AND U6673 ( .A(n861), .B(n7005), .Z(n7015) );
  XNOR U6674 ( .A(n7016), .B(n7003), .Z(n7005) );
  XOR U6675 ( .A(n7017), .B(n7018), .Z(n7003) );
  AND U6676 ( .A(n884), .B(n7019), .Z(n7018) );
  IV U6677 ( .A(n7014), .Z(n7016) );
  XOR U6678 ( .A(n7020), .B(n7021), .Z(n7014) );
  AND U6679 ( .A(n868), .B(n7013), .Z(n7021) );
  XNOR U6680 ( .A(n7011), .B(n7020), .Z(n7013) );
  XNOR U6681 ( .A(n7022), .B(n7023), .Z(n7011) );
  AND U6682 ( .A(n872), .B(n7024), .Z(n7023) );
  XOR U6683 ( .A(p_input[1279]), .B(n7022), .Z(n7024) );
  XNOR U6684 ( .A(n7025), .B(n7026), .Z(n7022) );
  AND U6685 ( .A(n876), .B(n7027), .Z(n7026) );
  XOR U6686 ( .A(n7028), .B(n7029), .Z(n7020) );
  AND U6687 ( .A(n880), .B(n7019), .Z(n7029) );
  XNOR U6688 ( .A(n7030), .B(n7017), .Z(n7019) );
  XOR U6689 ( .A(n7031), .B(n7032), .Z(n7017) );
  AND U6690 ( .A(n903), .B(n7033), .Z(n7032) );
  IV U6691 ( .A(n7028), .Z(n7030) );
  XOR U6692 ( .A(n7034), .B(n7035), .Z(n7028) );
  AND U6693 ( .A(n887), .B(n7027), .Z(n7035) );
  XNOR U6694 ( .A(n7025), .B(n7034), .Z(n7027) );
  XNOR U6695 ( .A(n7036), .B(n7037), .Z(n7025) );
  AND U6696 ( .A(n891), .B(n7038), .Z(n7037) );
  XOR U6697 ( .A(p_input[1311]), .B(n7036), .Z(n7038) );
  XNOR U6698 ( .A(n7039), .B(n7040), .Z(n7036) );
  AND U6699 ( .A(n895), .B(n7041), .Z(n7040) );
  XOR U6700 ( .A(n7042), .B(n7043), .Z(n7034) );
  AND U6701 ( .A(n899), .B(n7033), .Z(n7043) );
  XNOR U6702 ( .A(n7044), .B(n7031), .Z(n7033) );
  XOR U6703 ( .A(n7045), .B(n7046), .Z(n7031) );
  AND U6704 ( .A(n922), .B(n7047), .Z(n7046) );
  IV U6705 ( .A(n7042), .Z(n7044) );
  XOR U6706 ( .A(n7048), .B(n7049), .Z(n7042) );
  AND U6707 ( .A(n906), .B(n7041), .Z(n7049) );
  XNOR U6708 ( .A(n7039), .B(n7048), .Z(n7041) );
  XNOR U6709 ( .A(n7050), .B(n7051), .Z(n7039) );
  AND U6710 ( .A(n910), .B(n7052), .Z(n7051) );
  XOR U6711 ( .A(p_input[1343]), .B(n7050), .Z(n7052) );
  XNOR U6712 ( .A(n7053), .B(n7054), .Z(n7050) );
  AND U6713 ( .A(n914), .B(n7055), .Z(n7054) );
  XOR U6714 ( .A(n7056), .B(n7057), .Z(n7048) );
  AND U6715 ( .A(n918), .B(n7047), .Z(n7057) );
  XNOR U6716 ( .A(n7058), .B(n7045), .Z(n7047) );
  XOR U6717 ( .A(n7059), .B(n7060), .Z(n7045) );
  AND U6718 ( .A(n941), .B(n7061), .Z(n7060) );
  IV U6719 ( .A(n7056), .Z(n7058) );
  XOR U6720 ( .A(n7062), .B(n7063), .Z(n7056) );
  AND U6721 ( .A(n925), .B(n7055), .Z(n7063) );
  XNOR U6722 ( .A(n7053), .B(n7062), .Z(n7055) );
  XNOR U6723 ( .A(n7064), .B(n7065), .Z(n7053) );
  AND U6724 ( .A(n929), .B(n7066), .Z(n7065) );
  XOR U6725 ( .A(p_input[1375]), .B(n7064), .Z(n7066) );
  XNOR U6726 ( .A(n7067), .B(n7068), .Z(n7064) );
  AND U6727 ( .A(n933), .B(n7069), .Z(n7068) );
  XOR U6728 ( .A(n7070), .B(n7071), .Z(n7062) );
  AND U6729 ( .A(n937), .B(n7061), .Z(n7071) );
  XNOR U6730 ( .A(n7072), .B(n7059), .Z(n7061) );
  XOR U6731 ( .A(n7073), .B(n7074), .Z(n7059) );
  AND U6732 ( .A(n960), .B(n7075), .Z(n7074) );
  IV U6733 ( .A(n7070), .Z(n7072) );
  XOR U6734 ( .A(n7076), .B(n7077), .Z(n7070) );
  AND U6735 ( .A(n944), .B(n7069), .Z(n7077) );
  XNOR U6736 ( .A(n7067), .B(n7076), .Z(n7069) );
  XNOR U6737 ( .A(n7078), .B(n7079), .Z(n7067) );
  AND U6738 ( .A(n948), .B(n7080), .Z(n7079) );
  XOR U6739 ( .A(p_input[1407]), .B(n7078), .Z(n7080) );
  XNOR U6740 ( .A(n7081), .B(n7082), .Z(n7078) );
  AND U6741 ( .A(n952), .B(n7083), .Z(n7082) );
  XOR U6742 ( .A(n7084), .B(n7085), .Z(n7076) );
  AND U6743 ( .A(n956), .B(n7075), .Z(n7085) );
  XNOR U6744 ( .A(n7086), .B(n7073), .Z(n7075) );
  XOR U6745 ( .A(n7087), .B(n7088), .Z(n7073) );
  AND U6746 ( .A(n979), .B(n7089), .Z(n7088) );
  IV U6747 ( .A(n7084), .Z(n7086) );
  XOR U6748 ( .A(n7090), .B(n7091), .Z(n7084) );
  AND U6749 ( .A(n963), .B(n7083), .Z(n7091) );
  XNOR U6750 ( .A(n7081), .B(n7090), .Z(n7083) );
  XNOR U6751 ( .A(n7092), .B(n7093), .Z(n7081) );
  AND U6752 ( .A(n967), .B(n7094), .Z(n7093) );
  XOR U6753 ( .A(p_input[1439]), .B(n7092), .Z(n7094) );
  XNOR U6754 ( .A(n7095), .B(n7096), .Z(n7092) );
  AND U6755 ( .A(n971), .B(n7097), .Z(n7096) );
  XOR U6756 ( .A(n7098), .B(n7099), .Z(n7090) );
  AND U6757 ( .A(n975), .B(n7089), .Z(n7099) );
  XNOR U6758 ( .A(n7100), .B(n7087), .Z(n7089) );
  XOR U6759 ( .A(n7101), .B(n7102), .Z(n7087) );
  AND U6760 ( .A(n998), .B(n7103), .Z(n7102) );
  IV U6761 ( .A(n7098), .Z(n7100) );
  XOR U6762 ( .A(n7104), .B(n7105), .Z(n7098) );
  AND U6763 ( .A(n982), .B(n7097), .Z(n7105) );
  XNOR U6764 ( .A(n7095), .B(n7104), .Z(n7097) );
  XNOR U6765 ( .A(n7106), .B(n7107), .Z(n7095) );
  AND U6766 ( .A(n986), .B(n7108), .Z(n7107) );
  XOR U6767 ( .A(p_input[1471]), .B(n7106), .Z(n7108) );
  XNOR U6768 ( .A(n7109), .B(n7110), .Z(n7106) );
  AND U6769 ( .A(n990), .B(n7111), .Z(n7110) );
  XOR U6770 ( .A(n7112), .B(n7113), .Z(n7104) );
  AND U6771 ( .A(n994), .B(n7103), .Z(n7113) );
  XNOR U6772 ( .A(n7114), .B(n7101), .Z(n7103) );
  XOR U6773 ( .A(n7115), .B(n7116), .Z(n7101) );
  AND U6774 ( .A(n1017), .B(n7117), .Z(n7116) );
  IV U6775 ( .A(n7112), .Z(n7114) );
  XOR U6776 ( .A(n7118), .B(n7119), .Z(n7112) );
  AND U6777 ( .A(n1001), .B(n7111), .Z(n7119) );
  XNOR U6778 ( .A(n7109), .B(n7118), .Z(n7111) );
  XNOR U6779 ( .A(n7120), .B(n7121), .Z(n7109) );
  AND U6780 ( .A(n1005), .B(n7122), .Z(n7121) );
  XOR U6781 ( .A(p_input[1503]), .B(n7120), .Z(n7122) );
  XNOR U6782 ( .A(n7123), .B(n7124), .Z(n7120) );
  AND U6783 ( .A(n1009), .B(n7125), .Z(n7124) );
  XOR U6784 ( .A(n7126), .B(n7127), .Z(n7118) );
  AND U6785 ( .A(n1013), .B(n7117), .Z(n7127) );
  XNOR U6786 ( .A(n7128), .B(n7115), .Z(n7117) );
  XOR U6787 ( .A(n7129), .B(n7130), .Z(n7115) );
  AND U6788 ( .A(n1036), .B(n7131), .Z(n7130) );
  IV U6789 ( .A(n7126), .Z(n7128) );
  XOR U6790 ( .A(n7132), .B(n7133), .Z(n7126) );
  AND U6791 ( .A(n1020), .B(n7125), .Z(n7133) );
  XNOR U6792 ( .A(n7123), .B(n7132), .Z(n7125) );
  XNOR U6793 ( .A(n7134), .B(n7135), .Z(n7123) );
  AND U6794 ( .A(n1024), .B(n7136), .Z(n7135) );
  XOR U6795 ( .A(p_input[1535]), .B(n7134), .Z(n7136) );
  XNOR U6796 ( .A(n7137), .B(n7138), .Z(n7134) );
  AND U6797 ( .A(n1028), .B(n7139), .Z(n7138) );
  XOR U6798 ( .A(n7140), .B(n7141), .Z(n7132) );
  AND U6799 ( .A(n1032), .B(n7131), .Z(n7141) );
  XNOR U6800 ( .A(n7142), .B(n7129), .Z(n7131) );
  XOR U6801 ( .A(n7143), .B(n7144), .Z(n7129) );
  AND U6802 ( .A(n1055), .B(n7145), .Z(n7144) );
  IV U6803 ( .A(n7140), .Z(n7142) );
  XOR U6804 ( .A(n7146), .B(n7147), .Z(n7140) );
  AND U6805 ( .A(n1039), .B(n7139), .Z(n7147) );
  XNOR U6806 ( .A(n7137), .B(n7146), .Z(n7139) );
  XNOR U6807 ( .A(n7148), .B(n7149), .Z(n7137) );
  AND U6808 ( .A(n1043), .B(n7150), .Z(n7149) );
  XOR U6809 ( .A(p_input[1567]), .B(n7148), .Z(n7150) );
  XNOR U6810 ( .A(n7151), .B(n7152), .Z(n7148) );
  AND U6811 ( .A(n1047), .B(n7153), .Z(n7152) );
  XOR U6812 ( .A(n7154), .B(n7155), .Z(n7146) );
  AND U6813 ( .A(n1051), .B(n7145), .Z(n7155) );
  XNOR U6814 ( .A(n7156), .B(n7143), .Z(n7145) );
  XOR U6815 ( .A(n7157), .B(n7158), .Z(n7143) );
  AND U6816 ( .A(n1074), .B(n7159), .Z(n7158) );
  IV U6817 ( .A(n7154), .Z(n7156) );
  XOR U6818 ( .A(n7160), .B(n7161), .Z(n7154) );
  AND U6819 ( .A(n1058), .B(n7153), .Z(n7161) );
  XNOR U6820 ( .A(n7151), .B(n7160), .Z(n7153) );
  XNOR U6821 ( .A(n7162), .B(n7163), .Z(n7151) );
  AND U6822 ( .A(n1062), .B(n7164), .Z(n7163) );
  XOR U6823 ( .A(p_input[1599]), .B(n7162), .Z(n7164) );
  XNOR U6824 ( .A(n7165), .B(n7166), .Z(n7162) );
  AND U6825 ( .A(n1066), .B(n7167), .Z(n7166) );
  XOR U6826 ( .A(n7168), .B(n7169), .Z(n7160) );
  AND U6827 ( .A(n1070), .B(n7159), .Z(n7169) );
  XNOR U6828 ( .A(n7170), .B(n7157), .Z(n7159) );
  XOR U6829 ( .A(n7171), .B(n7172), .Z(n7157) );
  AND U6830 ( .A(n1093), .B(n7173), .Z(n7172) );
  IV U6831 ( .A(n7168), .Z(n7170) );
  XOR U6832 ( .A(n7174), .B(n7175), .Z(n7168) );
  AND U6833 ( .A(n1077), .B(n7167), .Z(n7175) );
  XNOR U6834 ( .A(n7165), .B(n7174), .Z(n7167) );
  XNOR U6835 ( .A(n7176), .B(n7177), .Z(n7165) );
  AND U6836 ( .A(n1081), .B(n7178), .Z(n7177) );
  XOR U6837 ( .A(p_input[1631]), .B(n7176), .Z(n7178) );
  XNOR U6838 ( .A(n7179), .B(n7180), .Z(n7176) );
  AND U6839 ( .A(n1085), .B(n7181), .Z(n7180) );
  XOR U6840 ( .A(n7182), .B(n7183), .Z(n7174) );
  AND U6841 ( .A(n1089), .B(n7173), .Z(n7183) );
  XNOR U6842 ( .A(n7184), .B(n7171), .Z(n7173) );
  XOR U6843 ( .A(n7185), .B(n7186), .Z(n7171) );
  AND U6844 ( .A(n1112), .B(n7187), .Z(n7186) );
  IV U6845 ( .A(n7182), .Z(n7184) );
  XOR U6846 ( .A(n7188), .B(n7189), .Z(n7182) );
  AND U6847 ( .A(n1096), .B(n7181), .Z(n7189) );
  XNOR U6848 ( .A(n7179), .B(n7188), .Z(n7181) );
  XNOR U6849 ( .A(n7190), .B(n7191), .Z(n7179) );
  AND U6850 ( .A(n1100), .B(n7192), .Z(n7191) );
  XOR U6851 ( .A(p_input[1663]), .B(n7190), .Z(n7192) );
  XNOR U6852 ( .A(n7193), .B(n7194), .Z(n7190) );
  AND U6853 ( .A(n1104), .B(n7195), .Z(n7194) );
  XOR U6854 ( .A(n7196), .B(n7197), .Z(n7188) );
  AND U6855 ( .A(n1108), .B(n7187), .Z(n7197) );
  XNOR U6856 ( .A(n7198), .B(n7185), .Z(n7187) );
  XOR U6857 ( .A(n7199), .B(n7200), .Z(n7185) );
  AND U6858 ( .A(n1131), .B(n7201), .Z(n7200) );
  IV U6859 ( .A(n7196), .Z(n7198) );
  XOR U6860 ( .A(n7202), .B(n7203), .Z(n7196) );
  AND U6861 ( .A(n1115), .B(n7195), .Z(n7203) );
  XNOR U6862 ( .A(n7193), .B(n7202), .Z(n7195) );
  XNOR U6863 ( .A(n7204), .B(n7205), .Z(n7193) );
  AND U6864 ( .A(n1119), .B(n7206), .Z(n7205) );
  XOR U6865 ( .A(p_input[1695]), .B(n7204), .Z(n7206) );
  XNOR U6866 ( .A(n7207), .B(n7208), .Z(n7204) );
  AND U6867 ( .A(n1123), .B(n7209), .Z(n7208) );
  XOR U6868 ( .A(n7210), .B(n7211), .Z(n7202) );
  AND U6869 ( .A(n1127), .B(n7201), .Z(n7211) );
  XNOR U6870 ( .A(n7212), .B(n7199), .Z(n7201) );
  XOR U6871 ( .A(n7213), .B(n7214), .Z(n7199) );
  AND U6872 ( .A(n1150), .B(n7215), .Z(n7214) );
  IV U6873 ( .A(n7210), .Z(n7212) );
  XOR U6874 ( .A(n7216), .B(n7217), .Z(n7210) );
  AND U6875 ( .A(n1134), .B(n7209), .Z(n7217) );
  XNOR U6876 ( .A(n7207), .B(n7216), .Z(n7209) );
  XNOR U6877 ( .A(n7218), .B(n7219), .Z(n7207) );
  AND U6878 ( .A(n1138), .B(n7220), .Z(n7219) );
  XOR U6879 ( .A(p_input[1727]), .B(n7218), .Z(n7220) );
  XNOR U6880 ( .A(n7221), .B(n7222), .Z(n7218) );
  AND U6881 ( .A(n1142), .B(n7223), .Z(n7222) );
  XOR U6882 ( .A(n7224), .B(n7225), .Z(n7216) );
  AND U6883 ( .A(n1146), .B(n7215), .Z(n7225) );
  XNOR U6884 ( .A(n7226), .B(n7213), .Z(n7215) );
  XOR U6885 ( .A(n7227), .B(n7228), .Z(n7213) );
  AND U6886 ( .A(n1169), .B(n7229), .Z(n7228) );
  IV U6887 ( .A(n7224), .Z(n7226) );
  XOR U6888 ( .A(n7230), .B(n7231), .Z(n7224) );
  AND U6889 ( .A(n1153), .B(n7223), .Z(n7231) );
  XNOR U6890 ( .A(n7221), .B(n7230), .Z(n7223) );
  XNOR U6891 ( .A(n7232), .B(n7233), .Z(n7221) );
  AND U6892 ( .A(n1157), .B(n7234), .Z(n7233) );
  XOR U6893 ( .A(p_input[1759]), .B(n7232), .Z(n7234) );
  XNOR U6894 ( .A(n7235), .B(n7236), .Z(n7232) );
  AND U6895 ( .A(n1161), .B(n7237), .Z(n7236) );
  XOR U6896 ( .A(n7238), .B(n7239), .Z(n7230) );
  AND U6897 ( .A(n1165), .B(n7229), .Z(n7239) );
  XNOR U6898 ( .A(n7240), .B(n7227), .Z(n7229) );
  XOR U6899 ( .A(n7241), .B(n7242), .Z(n7227) );
  AND U6900 ( .A(n1188), .B(n7243), .Z(n7242) );
  IV U6901 ( .A(n7238), .Z(n7240) );
  XOR U6902 ( .A(n7244), .B(n7245), .Z(n7238) );
  AND U6903 ( .A(n1172), .B(n7237), .Z(n7245) );
  XNOR U6904 ( .A(n7235), .B(n7244), .Z(n7237) );
  XNOR U6905 ( .A(n7246), .B(n7247), .Z(n7235) );
  AND U6906 ( .A(n1176), .B(n7248), .Z(n7247) );
  XOR U6907 ( .A(p_input[1791]), .B(n7246), .Z(n7248) );
  XNOR U6908 ( .A(n7249), .B(n7250), .Z(n7246) );
  AND U6909 ( .A(n1180), .B(n7251), .Z(n7250) );
  XOR U6910 ( .A(n7252), .B(n7253), .Z(n7244) );
  AND U6911 ( .A(n1184), .B(n7243), .Z(n7253) );
  XNOR U6912 ( .A(n7254), .B(n7241), .Z(n7243) );
  XOR U6913 ( .A(n7255), .B(n7256), .Z(n7241) );
  AND U6914 ( .A(n1207), .B(n7257), .Z(n7256) );
  IV U6915 ( .A(n7252), .Z(n7254) );
  XOR U6916 ( .A(n7258), .B(n7259), .Z(n7252) );
  AND U6917 ( .A(n1191), .B(n7251), .Z(n7259) );
  XNOR U6918 ( .A(n7249), .B(n7258), .Z(n7251) );
  XNOR U6919 ( .A(n7260), .B(n7261), .Z(n7249) );
  AND U6920 ( .A(n1195), .B(n7262), .Z(n7261) );
  XOR U6921 ( .A(p_input[1823]), .B(n7260), .Z(n7262) );
  XNOR U6922 ( .A(n7263), .B(n7264), .Z(n7260) );
  AND U6923 ( .A(n1199), .B(n7265), .Z(n7264) );
  XOR U6924 ( .A(n7266), .B(n7267), .Z(n7258) );
  AND U6925 ( .A(n1203), .B(n7257), .Z(n7267) );
  XNOR U6926 ( .A(n7268), .B(n7255), .Z(n7257) );
  XOR U6927 ( .A(n7269), .B(n7270), .Z(n7255) );
  AND U6928 ( .A(n1226), .B(n7271), .Z(n7270) );
  IV U6929 ( .A(n7266), .Z(n7268) );
  XOR U6930 ( .A(n7272), .B(n7273), .Z(n7266) );
  AND U6931 ( .A(n1210), .B(n7265), .Z(n7273) );
  XNOR U6932 ( .A(n7263), .B(n7272), .Z(n7265) );
  XNOR U6933 ( .A(n7274), .B(n7275), .Z(n7263) );
  AND U6934 ( .A(n1214), .B(n7276), .Z(n7275) );
  XOR U6935 ( .A(p_input[1855]), .B(n7274), .Z(n7276) );
  XNOR U6936 ( .A(n7277), .B(n7278), .Z(n7274) );
  AND U6937 ( .A(n1218), .B(n7279), .Z(n7278) );
  XOR U6938 ( .A(n7280), .B(n7281), .Z(n7272) );
  AND U6939 ( .A(n1222), .B(n7271), .Z(n7281) );
  XNOR U6940 ( .A(n7282), .B(n7269), .Z(n7271) );
  XOR U6941 ( .A(n7283), .B(n7284), .Z(n7269) );
  AND U6942 ( .A(n1245), .B(n7285), .Z(n7284) );
  IV U6943 ( .A(n7280), .Z(n7282) );
  XOR U6944 ( .A(n7286), .B(n7287), .Z(n7280) );
  AND U6945 ( .A(n1229), .B(n7279), .Z(n7287) );
  XNOR U6946 ( .A(n7277), .B(n7286), .Z(n7279) );
  XNOR U6947 ( .A(n7288), .B(n7289), .Z(n7277) );
  AND U6948 ( .A(n1233), .B(n7290), .Z(n7289) );
  XOR U6949 ( .A(p_input[1887]), .B(n7288), .Z(n7290) );
  XNOR U6950 ( .A(n7291), .B(n7292), .Z(n7288) );
  AND U6951 ( .A(n1237), .B(n7293), .Z(n7292) );
  XOR U6952 ( .A(n7294), .B(n7295), .Z(n7286) );
  AND U6953 ( .A(n1241), .B(n7285), .Z(n7295) );
  XNOR U6954 ( .A(n7296), .B(n7283), .Z(n7285) );
  XOR U6955 ( .A(n7297), .B(n7298), .Z(n7283) );
  AND U6956 ( .A(n1264), .B(n7299), .Z(n7298) );
  IV U6957 ( .A(n7294), .Z(n7296) );
  XOR U6958 ( .A(n7300), .B(n7301), .Z(n7294) );
  AND U6959 ( .A(n1248), .B(n7293), .Z(n7301) );
  XNOR U6960 ( .A(n7291), .B(n7300), .Z(n7293) );
  XNOR U6961 ( .A(n7302), .B(n7303), .Z(n7291) );
  AND U6962 ( .A(n1252), .B(n7304), .Z(n7303) );
  XOR U6963 ( .A(p_input[1919]), .B(n7302), .Z(n7304) );
  XNOR U6964 ( .A(n7305), .B(n7306), .Z(n7302) );
  AND U6965 ( .A(n1256), .B(n7307), .Z(n7306) );
  XOR U6966 ( .A(n7308), .B(n7309), .Z(n7300) );
  AND U6967 ( .A(n1260), .B(n7299), .Z(n7309) );
  XNOR U6968 ( .A(n7310), .B(n7297), .Z(n7299) );
  XOR U6969 ( .A(n7311), .B(n7312), .Z(n7297) );
  AND U6970 ( .A(n1282), .B(n7313), .Z(n7312) );
  IV U6971 ( .A(n7308), .Z(n7310) );
  XOR U6972 ( .A(n7314), .B(n7315), .Z(n7308) );
  AND U6973 ( .A(n1267), .B(n7307), .Z(n7315) );
  XNOR U6974 ( .A(n7305), .B(n7314), .Z(n7307) );
  XNOR U6975 ( .A(n7316), .B(n7317), .Z(n7305) );
  AND U6976 ( .A(n1271), .B(n7318), .Z(n7317) );
  XOR U6977 ( .A(p_input[1951]), .B(n7316), .Z(n7318) );
  XOR U6978 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][31] ), .B(n7319), 
        .Z(n7316) );
  AND U6979 ( .A(n1274), .B(n7320), .Z(n7319) );
  XOR U6980 ( .A(n7321), .B(n7322), .Z(n7314) );
  AND U6981 ( .A(n1278), .B(n7313), .Z(n7322) );
  XNOR U6982 ( .A(n7323), .B(n7311), .Z(n7313) );
  XOR U6983 ( .A(\knn_comb_/min_val_out[0][31] ), .B(n7324), .Z(n7311) );
  AND U6984 ( .A(n1290), .B(n7325), .Z(n7324) );
  IV U6985 ( .A(n7321), .Z(n7323) );
  XOR U6986 ( .A(n7326), .B(n7327), .Z(n7321) );
  AND U6987 ( .A(n1285), .B(n7320), .Z(n7327) );
  XOR U6988 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][31] ), .B(n7326), 
        .Z(n7320) );
  XOR U6989 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .B(n7328), 
        .Z(n7326) );
  AND U6990 ( .A(n1287), .B(n7325), .Z(n7328) );
  XOR U6991 ( .A(n7329), .B(n7330), .Z(n7325) );
  IV U6992 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .Z(n7330) );
  IV U6993 ( .A(\knn_comb_/min_val_out[0][31] ), .Z(n7329) );
  XOR U6994 ( .A(n75), .B(n7331), .Z(o[30]) );
  AND U6995 ( .A(n122), .B(n7332), .Z(n75) );
  XOR U6996 ( .A(n76), .B(n7331), .Z(n7332) );
  XOR U6997 ( .A(n7333), .B(n7334), .Z(n7331) );
  AND U6998 ( .A(n142), .B(n7335), .Z(n7334) );
  XOR U6999 ( .A(n7336), .B(n5), .Z(n76) );
  AND U7000 ( .A(n125), .B(n7337), .Z(n5) );
  XOR U7001 ( .A(n6), .B(n7336), .Z(n7337) );
  XOR U7002 ( .A(n7338), .B(n7339), .Z(n6) );
  AND U7003 ( .A(n130), .B(n7340), .Z(n7339) );
  XOR U7004 ( .A(p_input[30]), .B(n7338), .Z(n7340) );
  XNOR U7005 ( .A(n7341), .B(n7342), .Z(n7338) );
  AND U7006 ( .A(n134), .B(n7343), .Z(n7342) );
  XOR U7007 ( .A(n7344), .B(n7345), .Z(n7336) );
  AND U7008 ( .A(n138), .B(n7335), .Z(n7345) );
  XNOR U7009 ( .A(n7346), .B(n7333), .Z(n7335) );
  XOR U7010 ( .A(n7347), .B(n7348), .Z(n7333) );
  AND U7011 ( .A(n162), .B(n7349), .Z(n7348) );
  IV U7012 ( .A(n7344), .Z(n7346) );
  XOR U7013 ( .A(n7350), .B(n7351), .Z(n7344) );
  AND U7014 ( .A(n146), .B(n7343), .Z(n7351) );
  XNOR U7015 ( .A(n7341), .B(n7350), .Z(n7343) );
  XNOR U7016 ( .A(n7352), .B(n7353), .Z(n7341) );
  AND U7017 ( .A(n150), .B(n7354), .Z(n7353) );
  XOR U7018 ( .A(p_input[62]), .B(n7352), .Z(n7354) );
  XNOR U7019 ( .A(n7355), .B(n7356), .Z(n7352) );
  AND U7020 ( .A(n154), .B(n7357), .Z(n7356) );
  XOR U7021 ( .A(n7358), .B(n7359), .Z(n7350) );
  AND U7022 ( .A(n158), .B(n7349), .Z(n7359) );
  XNOR U7023 ( .A(n7360), .B(n7347), .Z(n7349) );
  XOR U7024 ( .A(n7361), .B(n7362), .Z(n7347) );
  AND U7025 ( .A(n181), .B(n7363), .Z(n7362) );
  IV U7026 ( .A(n7358), .Z(n7360) );
  XOR U7027 ( .A(n7364), .B(n7365), .Z(n7358) );
  AND U7028 ( .A(n165), .B(n7357), .Z(n7365) );
  XNOR U7029 ( .A(n7355), .B(n7364), .Z(n7357) );
  XNOR U7030 ( .A(n7366), .B(n7367), .Z(n7355) );
  AND U7031 ( .A(n169), .B(n7368), .Z(n7367) );
  XOR U7032 ( .A(p_input[94]), .B(n7366), .Z(n7368) );
  XNOR U7033 ( .A(n7369), .B(n7370), .Z(n7366) );
  AND U7034 ( .A(n173), .B(n7371), .Z(n7370) );
  XOR U7035 ( .A(n7372), .B(n7373), .Z(n7364) );
  AND U7036 ( .A(n177), .B(n7363), .Z(n7373) );
  XNOR U7037 ( .A(n7374), .B(n7361), .Z(n7363) );
  XOR U7038 ( .A(n7375), .B(n7376), .Z(n7361) );
  AND U7039 ( .A(n200), .B(n7377), .Z(n7376) );
  IV U7040 ( .A(n7372), .Z(n7374) );
  XOR U7041 ( .A(n7378), .B(n7379), .Z(n7372) );
  AND U7042 ( .A(n184), .B(n7371), .Z(n7379) );
  XNOR U7043 ( .A(n7369), .B(n7378), .Z(n7371) );
  XNOR U7044 ( .A(n7380), .B(n7381), .Z(n7369) );
  AND U7045 ( .A(n188), .B(n7382), .Z(n7381) );
  XOR U7046 ( .A(p_input[126]), .B(n7380), .Z(n7382) );
  XNOR U7047 ( .A(n7383), .B(n7384), .Z(n7380) );
  AND U7048 ( .A(n192), .B(n7385), .Z(n7384) );
  XOR U7049 ( .A(n7386), .B(n7387), .Z(n7378) );
  AND U7050 ( .A(n196), .B(n7377), .Z(n7387) );
  XNOR U7051 ( .A(n7388), .B(n7375), .Z(n7377) );
  XOR U7052 ( .A(n7389), .B(n7390), .Z(n7375) );
  AND U7053 ( .A(n219), .B(n7391), .Z(n7390) );
  IV U7054 ( .A(n7386), .Z(n7388) );
  XOR U7055 ( .A(n7392), .B(n7393), .Z(n7386) );
  AND U7056 ( .A(n203), .B(n7385), .Z(n7393) );
  XNOR U7057 ( .A(n7383), .B(n7392), .Z(n7385) );
  XNOR U7058 ( .A(n7394), .B(n7395), .Z(n7383) );
  AND U7059 ( .A(n207), .B(n7396), .Z(n7395) );
  XOR U7060 ( .A(p_input[158]), .B(n7394), .Z(n7396) );
  XNOR U7061 ( .A(n7397), .B(n7398), .Z(n7394) );
  AND U7062 ( .A(n211), .B(n7399), .Z(n7398) );
  XOR U7063 ( .A(n7400), .B(n7401), .Z(n7392) );
  AND U7064 ( .A(n215), .B(n7391), .Z(n7401) );
  XNOR U7065 ( .A(n7402), .B(n7389), .Z(n7391) );
  XOR U7066 ( .A(n7403), .B(n7404), .Z(n7389) );
  AND U7067 ( .A(n238), .B(n7405), .Z(n7404) );
  IV U7068 ( .A(n7400), .Z(n7402) );
  XOR U7069 ( .A(n7406), .B(n7407), .Z(n7400) );
  AND U7070 ( .A(n222), .B(n7399), .Z(n7407) );
  XNOR U7071 ( .A(n7397), .B(n7406), .Z(n7399) );
  XNOR U7072 ( .A(n7408), .B(n7409), .Z(n7397) );
  AND U7073 ( .A(n226), .B(n7410), .Z(n7409) );
  XOR U7074 ( .A(p_input[190]), .B(n7408), .Z(n7410) );
  XNOR U7075 ( .A(n7411), .B(n7412), .Z(n7408) );
  AND U7076 ( .A(n230), .B(n7413), .Z(n7412) );
  XOR U7077 ( .A(n7414), .B(n7415), .Z(n7406) );
  AND U7078 ( .A(n234), .B(n7405), .Z(n7415) );
  XNOR U7079 ( .A(n7416), .B(n7403), .Z(n7405) );
  XOR U7080 ( .A(n7417), .B(n7418), .Z(n7403) );
  AND U7081 ( .A(n257), .B(n7419), .Z(n7418) );
  IV U7082 ( .A(n7414), .Z(n7416) );
  XOR U7083 ( .A(n7420), .B(n7421), .Z(n7414) );
  AND U7084 ( .A(n241), .B(n7413), .Z(n7421) );
  XNOR U7085 ( .A(n7411), .B(n7420), .Z(n7413) );
  XNOR U7086 ( .A(n7422), .B(n7423), .Z(n7411) );
  AND U7087 ( .A(n245), .B(n7424), .Z(n7423) );
  XOR U7088 ( .A(p_input[222]), .B(n7422), .Z(n7424) );
  XNOR U7089 ( .A(n7425), .B(n7426), .Z(n7422) );
  AND U7090 ( .A(n249), .B(n7427), .Z(n7426) );
  XOR U7091 ( .A(n7428), .B(n7429), .Z(n7420) );
  AND U7092 ( .A(n253), .B(n7419), .Z(n7429) );
  XNOR U7093 ( .A(n7430), .B(n7417), .Z(n7419) );
  XOR U7094 ( .A(n7431), .B(n7432), .Z(n7417) );
  AND U7095 ( .A(n276), .B(n7433), .Z(n7432) );
  IV U7096 ( .A(n7428), .Z(n7430) );
  XOR U7097 ( .A(n7434), .B(n7435), .Z(n7428) );
  AND U7098 ( .A(n260), .B(n7427), .Z(n7435) );
  XNOR U7099 ( .A(n7425), .B(n7434), .Z(n7427) );
  XNOR U7100 ( .A(n7436), .B(n7437), .Z(n7425) );
  AND U7101 ( .A(n264), .B(n7438), .Z(n7437) );
  XOR U7102 ( .A(p_input[254]), .B(n7436), .Z(n7438) );
  XNOR U7103 ( .A(n7439), .B(n7440), .Z(n7436) );
  AND U7104 ( .A(n268), .B(n7441), .Z(n7440) );
  XOR U7105 ( .A(n7442), .B(n7443), .Z(n7434) );
  AND U7106 ( .A(n272), .B(n7433), .Z(n7443) );
  XNOR U7107 ( .A(n7444), .B(n7431), .Z(n7433) );
  XOR U7108 ( .A(n7445), .B(n7446), .Z(n7431) );
  AND U7109 ( .A(n295), .B(n7447), .Z(n7446) );
  IV U7110 ( .A(n7442), .Z(n7444) );
  XOR U7111 ( .A(n7448), .B(n7449), .Z(n7442) );
  AND U7112 ( .A(n279), .B(n7441), .Z(n7449) );
  XNOR U7113 ( .A(n7439), .B(n7448), .Z(n7441) );
  XNOR U7114 ( .A(n7450), .B(n7451), .Z(n7439) );
  AND U7115 ( .A(n283), .B(n7452), .Z(n7451) );
  XOR U7116 ( .A(p_input[286]), .B(n7450), .Z(n7452) );
  XNOR U7117 ( .A(n7453), .B(n7454), .Z(n7450) );
  AND U7118 ( .A(n287), .B(n7455), .Z(n7454) );
  XOR U7119 ( .A(n7456), .B(n7457), .Z(n7448) );
  AND U7120 ( .A(n291), .B(n7447), .Z(n7457) );
  XNOR U7121 ( .A(n7458), .B(n7445), .Z(n7447) );
  XOR U7122 ( .A(n7459), .B(n7460), .Z(n7445) );
  AND U7123 ( .A(n314), .B(n7461), .Z(n7460) );
  IV U7124 ( .A(n7456), .Z(n7458) );
  XOR U7125 ( .A(n7462), .B(n7463), .Z(n7456) );
  AND U7126 ( .A(n298), .B(n7455), .Z(n7463) );
  XNOR U7127 ( .A(n7453), .B(n7462), .Z(n7455) );
  XNOR U7128 ( .A(n7464), .B(n7465), .Z(n7453) );
  AND U7129 ( .A(n302), .B(n7466), .Z(n7465) );
  XOR U7130 ( .A(p_input[318]), .B(n7464), .Z(n7466) );
  XNOR U7131 ( .A(n7467), .B(n7468), .Z(n7464) );
  AND U7132 ( .A(n306), .B(n7469), .Z(n7468) );
  XOR U7133 ( .A(n7470), .B(n7471), .Z(n7462) );
  AND U7134 ( .A(n310), .B(n7461), .Z(n7471) );
  XNOR U7135 ( .A(n7472), .B(n7459), .Z(n7461) );
  XOR U7136 ( .A(n7473), .B(n7474), .Z(n7459) );
  AND U7137 ( .A(n333), .B(n7475), .Z(n7474) );
  IV U7138 ( .A(n7470), .Z(n7472) );
  XOR U7139 ( .A(n7476), .B(n7477), .Z(n7470) );
  AND U7140 ( .A(n317), .B(n7469), .Z(n7477) );
  XNOR U7141 ( .A(n7467), .B(n7476), .Z(n7469) );
  XNOR U7142 ( .A(n7478), .B(n7479), .Z(n7467) );
  AND U7143 ( .A(n321), .B(n7480), .Z(n7479) );
  XOR U7144 ( .A(p_input[350]), .B(n7478), .Z(n7480) );
  XNOR U7145 ( .A(n7481), .B(n7482), .Z(n7478) );
  AND U7146 ( .A(n325), .B(n7483), .Z(n7482) );
  XOR U7147 ( .A(n7484), .B(n7485), .Z(n7476) );
  AND U7148 ( .A(n329), .B(n7475), .Z(n7485) );
  XNOR U7149 ( .A(n7486), .B(n7473), .Z(n7475) );
  XOR U7150 ( .A(n7487), .B(n7488), .Z(n7473) );
  AND U7151 ( .A(n352), .B(n7489), .Z(n7488) );
  IV U7152 ( .A(n7484), .Z(n7486) );
  XOR U7153 ( .A(n7490), .B(n7491), .Z(n7484) );
  AND U7154 ( .A(n336), .B(n7483), .Z(n7491) );
  XNOR U7155 ( .A(n7481), .B(n7490), .Z(n7483) );
  XNOR U7156 ( .A(n7492), .B(n7493), .Z(n7481) );
  AND U7157 ( .A(n340), .B(n7494), .Z(n7493) );
  XOR U7158 ( .A(p_input[382]), .B(n7492), .Z(n7494) );
  XNOR U7159 ( .A(n7495), .B(n7496), .Z(n7492) );
  AND U7160 ( .A(n344), .B(n7497), .Z(n7496) );
  XOR U7161 ( .A(n7498), .B(n7499), .Z(n7490) );
  AND U7162 ( .A(n348), .B(n7489), .Z(n7499) );
  XNOR U7163 ( .A(n7500), .B(n7487), .Z(n7489) );
  XOR U7164 ( .A(n7501), .B(n7502), .Z(n7487) );
  AND U7165 ( .A(n371), .B(n7503), .Z(n7502) );
  IV U7166 ( .A(n7498), .Z(n7500) );
  XOR U7167 ( .A(n7504), .B(n7505), .Z(n7498) );
  AND U7168 ( .A(n355), .B(n7497), .Z(n7505) );
  XNOR U7169 ( .A(n7495), .B(n7504), .Z(n7497) );
  XNOR U7170 ( .A(n7506), .B(n7507), .Z(n7495) );
  AND U7171 ( .A(n359), .B(n7508), .Z(n7507) );
  XOR U7172 ( .A(p_input[414]), .B(n7506), .Z(n7508) );
  XNOR U7173 ( .A(n7509), .B(n7510), .Z(n7506) );
  AND U7174 ( .A(n363), .B(n7511), .Z(n7510) );
  XOR U7175 ( .A(n7512), .B(n7513), .Z(n7504) );
  AND U7176 ( .A(n367), .B(n7503), .Z(n7513) );
  XNOR U7177 ( .A(n7514), .B(n7501), .Z(n7503) );
  XOR U7178 ( .A(n7515), .B(n7516), .Z(n7501) );
  AND U7179 ( .A(n390), .B(n7517), .Z(n7516) );
  IV U7180 ( .A(n7512), .Z(n7514) );
  XOR U7181 ( .A(n7518), .B(n7519), .Z(n7512) );
  AND U7182 ( .A(n374), .B(n7511), .Z(n7519) );
  XNOR U7183 ( .A(n7509), .B(n7518), .Z(n7511) );
  XNOR U7184 ( .A(n7520), .B(n7521), .Z(n7509) );
  AND U7185 ( .A(n378), .B(n7522), .Z(n7521) );
  XOR U7186 ( .A(p_input[446]), .B(n7520), .Z(n7522) );
  XNOR U7187 ( .A(n7523), .B(n7524), .Z(n7520) );
  AND U7188 ( .A(n382), .B(n7525), .Z(n7524) );
  XOR U7189 ( .A(n7526), .B(n7527), .Z(n7518) );
  AND U7190 ( .A(n386), .B(n7517), .Z(n7527) );
  XNOR U7191 ( .A(n7528), .B(n7515), .Z(n7517) );
  XOR U7192 ( .A(n7529), .B(n7530), .Z(n7515) );
  AND U7193 ( .A(n409), .B(n7531), .Z(n7530) );
  IV U7194 ( .A(n7526), .Z(n7528) );
  XOR U7195 ( .A(n7532), .B(n7533), .Z(n7526) );
  AND U7196 ( .A(n393), .B(n7525), .Z(n7533) );
  XNOR U7197 ( .A(n7523), .B(n7532), .Z(n7525) );
  XNOR U7198 ( .A(n7534), .B(n7535), .Z(n7523) );
  AND U7199 ( .A(n397), .B(n7536), .Z(n7535) );
  XOR U7200 ( .A(p_input[478]), .B(n7534), .Z(n7536) );
  XNOR U7201 ( .A(n7537), .B(n7538), .Z(n7534) );
  AND U7202 ( .A(n401), .B(n7539), .Z(n7538) );
  XOR U7203 ( .A(n7540), .B(n7541), .Z(n7532) );
  AND U7204 ( .A(n405), .B(n7531), .Z(n7541) );
  XNOR U7205 ( .A(n7542), .B(n7529), .Z(n7531) );
  XOR U7206 ( .A(n7543), .B(n7544), .Z(n7529) );
  AND U7207 ( .A(n428), .B(n7545), .Z(n7544) );
  IV U7208 ( .A(n7540), .Z(n7542) );
  XOR U7209 ( .A(n7546), .B(n7547), .Z(n7540) );
  AND U7210 ( .A(n412), .B(n7539), .Z(n7547) );
  XNOR U7211 ( .A(n7537), .B(n7546), .Z(n7539) );
  XNOR U7212 ( .A(n7548), .B(n7549), .Z(n7537) );
  AND U7213 ( .A(n416), .B(n7550), .Z(n7549) );
  XOR U7214 ( .A(p_input[510]), .B(n7548), .Z(n7550) );
  XNOR U7215 ( .A(n7551), .B(n7552), .Z(n7548) );
  AND U7216 ( .A(n420), .B(n7553), .Z(n7552) );
  XOR U7217 ( .A(n7554), .B(n7555), .Z(n7546) );
  AND U7218 ( .A(n424), .B(n7545), .Z(n7555) );
  XNOR U7219 ( .A(n7556), .B(n7543), .Z(n7545) );
  XOR U7220 ( .A(n7557), .B(n7558), .Z(n7543) );
  AND U7221 ( .A(n447), .B(n7559), .Z(n7558) );
  IV U7222 ( .A(n7554), .Z(n7556) );
  XOR U7223 ( .A(n7560), .B(n7561), .Z(n7554) );
  AND U7224 ( .A(n431), .B(n7553), .Z(n7561) );
  XNOR U7225 ( .A(n7551), .B(n7560), .Z(n7553) );
  XNOR U7226 ( .A(n7562), .B(n7563), .Z(n7551) );
  AND U7227 ( .A(n435), .B(n7564), .Z(n7563) );
  XOR U7228 ( .A(p_input[542]), .B(n7562), .Z(n7564) );
  XNOR U7229 ( .A(n7565), .B(n7566), .Z(n7562) );
  AND U7230 ( .A(n439), .B(n7567), .Z(n7566) );
  XOR U7231 ( .A(n7568), .B(n7569), .Z(n7560) );
  AND U7232 ( .A(n443), .B(n7559), .Z(n7569) );
  XNOR U7233 ( .A(n7570), .B(n7557), .Z(n7559) );
  XOR U7234 ( .A(n7571), .B(n7572), .Z(n7557) );
  AND U7235 ( .A(n466), .B(n7573), .Z(n7572) );
  IV U7236 ( .A(n7568), .Z(n7570) );
  XOR U7237 ( .A(n7574), .B(n7575), .Z(n7568) );
  AND U7238 ( .A(n450), .B(n7567), .Z(n7575) );
  XNOR U7239 ( .A(n7565), .B(n7574), .Z(n7567) );
  XNOR U7240 ( .A(n7576), .B(n7577), .Z(n7565) );
  AND U7241 ( .A(n454), .B(n7578), .Z(n7577) );
  XOR U7242 ( .A(p_input[574]), .B(n7576), .Z(n7578) );
  XNOR U7243 ( .A(n7579), .B(n7580), .Z(n7576) );
  AND U7244 ( .A(n458), .B(n7581), .Z(n7580) );
  XOR U7245 ( .A(n7582), .B(n7583), .Z(n7574) );
  AND U7246 ( .A(n462), .B(n7573), .Z(n7583) );
  XNOR U7247 ( .A(n7584), .B(n7571), .Z(n7573) );
  XOR U7248 ( .A(n7585), .B(n7586), .Z(n7571) );
  AND U7249 ( .A(n485), .B(n7587), .Z(n7586) );
  IV U7250 ( .A(n7582), .Z(n7584) );
  XOR U7251 ( .A(n7588), .B(n7589), .Z(n7582) );
  AND U7252 ( .A(n469), .B(n7581), .Z(n7589) );
  XNOR U7253 ( .A(n7579), .B(n7588), .Z(n7581) );
  XNOR U7254 ( .A(n7590), .B(n7591), .Z(n7579) );
  AND U7255 ( .A(n473), .B(n7592), .Z(n7591) );
  XOR U7256 ( .A(p_input[606]), .B(n7590), .Z(n7592) );
  XNOR U7257 ( .A(n7593), .B(n7594), .Z(n7590) );
  AND U7258 ( .A(n477), .B(n7595), .Z(n7594) );
  XOR U7259 ( .A(n7596), .B(n7597), .Z(n7588) );
  AND U7260 ( .A(n481), .B(n7587), .Z(n7597) );
  XNOR U7261 ( .A(n7598), .B(n7585), .Z(n7587) );
  XOR U7262 ( .A(n7599), .B(n7600), .Z(n7585) );
  AND U7263 ( .A(n504), .B(n7601), .Z(n7600) );
  IV U7264 ( .A(n7596), .Z(n7598) );
  XOR U7265 ( .A(n7602), .B(n7603), .Z(n7596) );
  AND U7266 ( .A(n488), .B(n7595), .Z(n7603) );
  XNOR U7267 ( .A(n7593), .B(n7602), .Z(n7595) );
  XNOR U7268 ( .A(n7604), .B(n7605), .Z(n7593) );
  AND U7269 ( .A(n492), .B(n7606), .Z(n7605) );
  XOR U7270 ( .A(p_input[638]), .B(n7604), .Z(n7606) );
  XNOR U7271 ( .A(n7607), .B(n7608), .Z(n7604) );
  AND U7272 ( .A(n496), .B(n7609), .Z(n7608) );
  XOR U7273 ( .A(n7610), .B(n7611), .Z(n7602) );
  AND U7274 ( .A(n500), .B(n7601), .Z(n7611) );
  XNOR U7275 ( .A(n7612), .B(n7599), .Z(n7601) );
  XOR U7276 ( .A(n7613), .B(n7614), .Z(n7599) );
  AND U7277 ( .A(n523), .B(n7615), .Z(n7614) );
  IV U7278 ( .A(n7610), .Z(n7612) );
  XOR U7279 ( .A(n7616), .B(n7617), .Z(n7610) );
  AND U7280 ( .A(n507), .B(n7609), .Z(n7617) );
  XNOR U7281 ( .A(n7607), .B(n7616), .Z(n7609) );
  XNOR U7282 ( .A(n7618), .B(n7619), .Z(n7607) );
  AND U7283 ( .A(n511), .B(n7620), .Z(n7619) );
  XOR U7284 ( .A(p_input[670]), .B(n7618), .Z(n7620) );
  XNOR U7285 ( .A(n7621), .B(n7622), .Z(n7618) );
  AND U7286 ( .A(n515), .B(n7623), .Z(n7622) );
  XOR U7287 ( .A(n7624), .B(n7625), .Z(n7616) );
  AND U7288 ( .A(n519), .B(n7615), .Z(n7625) );
  XNOR U7289 ( .A(n7626), .B(n7613), .Z(n7615) );
  XOR U7290 ( .A(n7627), .B(n7628), .Z(n7613) );
  AND U7291 ( .A(n542), .B(n7629), .Z(n7628) );
  IV U7292 ( .A(n7624), .Z(n7626) );
  XOR U7293 ( .A(n7630), .B(n7631), .Z(n7624) );
  AND U7294 ( .A(n526), .B(n7623), .Z(n7631) );
  XNOR U7295 ( .A(n7621), .B(n7630), .Z(n7623) );
  XNOR U7296 ( .A(n7632), .B(n7633), .Z(n7621) );
  AND U7297 ( .A(n530), .B(n7634), .Z(n7633) );
  XOR U7298 ( .A(p_input[702]), .B(n7632), .Z(n7634) );
  XNOR U7299 ( .A(n7635), .B(n7636), .Z(n7632) );
  AND U7300 ( .A(n534), .B(n7637), .Z(n7636) );
  XOR U7301 ( .A(n7638), .B(n7639), .Z(n7630) );
  AND U7302 ( .A(n538), .B(n7629), .Z(n7639) );
  XNOR U7303 ( .A(n7640), .B(n7627), .Z(n7629) );
  XOR U7304 ( .A(n7641), .B(n7642), .Z(n7627) );
  AND U7305 ( .A(n561), .B(n7643), .Z(n7642) );
  IV U7306 ( .A(n7638), .Z(n7640) );
  XOR U7307 ( .A(n7644), .B(n7645), .Z(n7638) );
  AND U7308 ( .A(n545), .B(n7637), .Z(n7645) );
  XNOR U7309 ( .A(n7635), .B(n7644), .Z(n7637) );
  XNOR U7310 ( .A(n7646), .B(n7647), .Z(n7635) );
  AND U7311 ( .A(n549), .B(n7648), .Z(n7647) );
  XOR U7312 ( .A(p_input[734]), .B(n7646), .Z(n7648) );
  XNOR U7313 ( .A(n7649), .B(n7650), .Z(n7646) );
  AND U7314 ( .A(n553), .B(n7651), .Z(n7650) );
  XOR U7315 ( .A(n7652), .B(n7653), .Z(n7644) );
  AND U7316 ( .A(n557), .B(n7643), .Z(n7653) );
  XNOR U7317 ( .A(n7654), .B(n7641), .Z(n7643) );
  XOR U7318 ( .A(n7655), .B(n7656), .Z(n7641) );
  AND U7319 ( .A(n580), .B(n7657), .Z(n7656) );
  IV U7320 ( .A(n7652), .Z(n7654) );
  XOR U7321 ( .A(n7658), .B(n7659), .Z(n7652) );
  AND U7322 ( .A(n564), .B(n7651), .Z(n7659) );
  XNOR U7323 ( .A(n7649), .B(n7658), .Z(n7651) );
  XNOR U7324 ( .A(n7660), .B(n7661), .Z(n7649) );
  AND U7325 ( .A(n568), .B(n7662), .Z(n7661) );
  XOR U7326 ( .A(p_input[766]), .B(n7660), .Z(n7662) );
  XNOR U7327 ( .A(n7663), .B(n7664), .Z(n7660) );
  AND U7328 ( .A(n572), .B(n7665), .Z(n7664) );
  XOR U7329 ( .A(n7666), .B(n7667), .Z(n7658) );
  AND U7330 ( .A(n576), .B(n7657), .Z(n7667) );
  XNOR U7331 ( .A(n7668), .B(n7655), .Z(n7657) );
  XOR U7332 ( .A(n7669), .B(n7670), .Z(n7655) );
  AND U7333 ( .A(n599), .B(n7671), .Z(n7670) );
  IV U7334 ( .A(n7666), .Z(n7668) );
  XOR U7335 ( .A(n7672), .B(n7673), .Z(n7666) );
  AND U7336 ( .A(n583), .B(n7665), .Z(n7673) );
  XNOR U7337 ( .A(n7663), .B(n7672), .Z(n7665) );
  XNOR U7338 ( .A(n7674), .B(n7675), .Z(n7663) );
  AND U7339 ( .A(n587), .B(n7676), .Z(n7675) );
  XOR U7340 ( .A(p_input[798]), .B(n7674), .Z(n7676) );
  XNOR U7341 ( .A(n7677), .B(n7678), .Z(n7674) );
  AND U7342 ( .A(n591), .B(n7679), .Z(n7678) );
  XOR U7343 ( .A(n7680), .B(n7681), .Z(n7672) );
  AND U7344 ( .A(n595), .B(n7671), .Z(n7681) );
  XNOR U7345 ( .A(n7682), .B(n7669), .Z(n7671) );
  XOR U7346 ( .A(n7683), .B(n7684), .Z(n7669) );
  AND U7347 ( .A(n618), .B(n7685), .Z(n7684) );
  IV U7348 ( .A(n7680), .Z(n7682) );
  XOR U7349 ( .A(n7686), .B(n7687), .Z(n7680) );
  AND U7350 ( .A(n602), .B(n7679), .Z(n7687) );
  XNOR U7351 ( .A(n7677), .B(n7686), .Z(n7679) );
  XNOR U7352 ( .A(n7688), .B(n7689), .Z(n7677) );
  AND U7353 ( .A(n606), .B(n7690), .Z(n7689) );
  XOR U7354 ( .A(p_input[830]), .B(n7688), .Z(n7690) );
  XNOR U7355 ( .A(n7691), .B(n7692), .Z(n7688) );
  AND U7356 ( .A(n610), .B(n7693), .Z(n7692) );
  XOR U7357 ( .A(n7694), .B(n7695), .Z(n7686) );
  AND U7358 ( .A(n614), .B(n7685), .Z(n7695) );
  XNOR U7359 ( .A(n7696), .B(n7683), .Z(n7685) );
  XOR U7360 ( .A(n7697), .B(n7698), .Z(n7683) );
  AND U7361 ( .A(n637), .B(n7699), .Z(n7698) );
  IV U7362 ( .A(n7694), .Z(n7696) );
  XOR U7363 ( .A(n7700), .B(n7701), .Z(n7694) );
  AND U7364 ( .A(n621), .B(n7693), .Z(n7701) );
  XNOR U7365 ( .A(n7691), .B(n7700), .Z(n7693) );
  XNOR U7366 ( .A(n7702), .B(n7703), .Z(n7691) );
  AND U7367 ( .A(n625), .B(n7704), .Z(n7703) );
  XOR U7368 ( .A(p_input[862]), .B(n7702), .Z(n7704) );
  XNOR U7369 ( .A(n7705), .B(n7706), .Z(n7702) );
  AND U7370 ( .A(n629), .B(n7707), .Z(n7706) );
  XOR U7371 ( .A(n7708), .B(n7709), .Z(n7700) );
  AND U7372 ( .A(n633), .B(n7699), .Z(n7709) );
  XNOR U7373 ( .A(n7710), .B(n7697), .Z(n7699) );
  XOR U7374 ( .A(n7711), .B(n7712), .Z(n7697) );
  AND U7375 ( .A(n656), .B(n7713), .Z(n7712) );
  IV U7376 ( .A(n7708), .Z(n7710) );
  XOR U7377 ( .A(n7714), .B(n7715), .Z(n7708) );
  AND U7378 ( .A(n640), .B(n7707), .Z(n7715) );
  XNOR U7379 ( .A(n7705), .B(n7714), .Z(n7707) );
  XNOR U7380 ( .A(n7716), .B(n7717), .Z(n7705) );
  AND U7381 ( .A(n644), .B(n7718), .Z(n7717) );
  XOR U7382 ( .A(p_input[894]), .B(n7716), .Z(n7718) );
  XNOR U7383 ( .A(n7719), .B(n7720), .Z(n7716) );
  AND U7384 ( .A(n648), .B(n7721), .Z(n7720) );
  XOR U7385 ( .A(n7722), .B(n7723), .Z(n7714) );
  AND U7386 ( .A(n652), .B(n7713), .Z(n7723) );
  XNOR U7387 ( .A(n7724), .B(n7711), .Z(n7713) );
  XOR U7388 ( .A(n7725), .B(n7726), .Z(n7711) );
  AND U7389 ( .A(n675), .B(n7727), .Z(n7726) );
  IV U7390 ( .A(n7722), .Z(n7724) );
  XOR U7391 ( .A(n7728), .B(n7729), .Z(n7722) );
  AND U7392 ( .A(n659), .B(n7721), .Z(n7729) );
  XNOR U7393 ( .A(n7719), .B(n7728), .Z(n7721) );
  XNOR U7394 ( .A(n7730), .B(n7731), .Z(n7719) );
  AND U7395 ( .A(n663), .B(n7732), .Z(n7731) );
  XOR U7396 ( .A(p_input[926]), .B(n7730), .Z(n7732) );
  XNOR U7397 ( .A(n7733), .B(n7734), .Z(n7730) );
  AND U7398 ( .A(n667), .B(n7735), .Z(n7734) );
  XOR U7399 ( .A(n7736), .B(n7737), .Z(n7728) );
  AND U7400 ( .A(n671), .B(n7727), .Z(n7737) );
  XNOR U7401 ( .A(n7738), .B(n7725), .Z(n7727) );
  XOR U7402 ( .A(n7739), .B(n7740), .Z(n7725) );
  AND U7403 ( .A(n694), .B(n7741), .Z(n7740) );
  IV U7404 ( .A(n7736), .Z(n7738) );
  XOR U7405 ( .A(n7742), .B(n7743), .Z(n7736) );
  AND U7406 ( .A(n678), .B(n7735), .Z(n7743) );
  XNOR U7407 ( .A(n7733), .B(n7742), .Z(n7735) );
  XNOR U7408 ( .A(n7744), .B(n7745), .Z(n7733) );
  AND U7409 ( .A(n682), .B(n7746), .Z(n7745) );
  XOR U7410 ( .A(p_input[958]), .B(n7744), .Z(n7746) );
  XNOR U7411 ( .A(n7747), .B(n7748), .Z(n7744) );
  AND U7412 ( .A(n686), .B(n7749), .Z(n7748) );
  XOR U7413 ( .A(n7750), .B(n7751), .Z(n7742) );
  AND U7414 ( .A(n690), .B(n7741), .Z(n7751) );
  XNOR U7415 ( .A(n7752), .B(n7739), .Z(n7741) );
  XOR U7416 ( .A(n7753), .B(n7754), .Z(n7739) );
  AND U7417 ( .A(n713), .B(n7755), .Z(n7754) );
  IV U7418 ( .A(n7750), .Z(n7752) );
  XOR U7419 ( .A(n7756), .B(n7757), .Z(n7750) );
  AND U7420 ( .A(n697), .B(n7749), .Z(n7757) );
  XNOR U7421 ( .A(n7747), .B(n7756), .Z(n7749) );
  XNOR U7422 ( .A(n7758), .B(n7759), .Z(n7747) );
  AND U7423 ( .A(n701), .B(n7760), .Z(n7759) );
  XOR U7424 ( .A(p_input[990]), .B(n7758), .Z(n7760) );
  XNOR U7425 ( .A(n7761), .B(n7762), .Z(n7758) );
  AND U7426 ( .A(n705), .B(n7763), .Z(n7762) );
  XOR U7427 ( .A(n7764), .B(n7765), .Z(n7756) );
  AND U7428 ( .A(n709), .B(n7755), .Z(n7765) );
  XNOR U7429 ( .A(n7766), .B(n7753), .Z(n7755) );
  XOR U7430 ( .A(n7767), .B(n7768), .Z(n7753) );
  AND U7431 ( .A(n732), .B(n7769), .Z(n7768) );
  IV U7432 ( .A(n7764), .Z(n7766) );
  XOR U7433 ( .A(n7770), .B(n7771), .Z(n7764) );
  AND U7434 ( .A(n716), .B(n7763), .Z(n7771) );
  XNOR U7435 ( .A(n7761), .B(n7770), .Z(n7763) );
  XNOR U7436 ( .A(n7772), .B(n7773), .Z(n7761) );
  AND U7437 ( .A(n720), .B(n7774), .Z(n7773) );
  XOR U7438 ( .A(p_input[1022]), .B(n7772), .Z(n7774) );
  XNOR U7439 ( .A(n7775), .B(n7776), .Z(n7772) );
  AND U7440 ( .A(n724), .B(n7777), .Z(n7776) );
  XOR U7441 ( .A(n7778), .B(n7779), .Z(n7770) );
  AND U7442 ( .A(n728), .B(n7769), .Z(n7779) );
  XNOR U7443 ( .A(n7780), .B(n7767), .Z(n7769) );
  XOR U7444 ( .A(n7781), .B(n7782), .Z(n7767) );
  AND U7445 ( .A(n751), .B(n7783), .Z(n7782) );
  IV U7446 ( .A(n7778), .Z(n7780) );
  XOR U7447 ( .A(n7784), .B(n7785), .Z(n7778) );
  AND U7448 ( .A(n735), .B(n7777), .Z(n7785) );
  XNOR U7449 ( .A(n7775), .B(n7784), .Z(n7777) );
  XNOR U7450 ( .A(n7786), .B(n7787), .Z(n7775) );
  AND U7451 ( .A(n739), .B(n7788), .Z(n7787) );
  XOR U7452 ( .A(p_input[1054]), .B(n7786), .Z(n7788) );
  XNOR U7453 ( .A(n7789), .B(n7790), .Z(n7786) );
  AND U7454 ( .A(n743), .B(n7791), .Z(n7790) );
  XOR U7455 ( .A(n7792), .B(n7793), .Z(n7784) );
  AND U7456 ( .A(n747), .B(n7783), .Z(n7793) );
  XNOR U7457 ( .A(n7794), .B(n7781), .Z(n7783) );
  XOR U7458 ( .A(n7795), .B(n7796), .Z(n7781) );
  AND U7459 ( .A(n770), .B(n7797), .Z(n7796) );
  IV U7460 ( .A(n7792), .Z(n7794) );
  XOR U7461 ( .A(n7798), .B(n7799), .Z(n7792) );
  AND U7462 ( .A(n754), .B(n7791), .Z(n7799) );
  XNOR U7463 ( .A(n7789), .B(n7798), .Z(n7791) );
  XNOR U7464 ( .A(n7800), .B(n7801), .Z(n7789) );
  AND U7465 ( .A(n758), .B(n7802), .Z(n7801) );
  XOR U7466 ( .A(p_input[1086]), .B(n7800), .Z(n7802) );
  XNOR U7467 ( .A(n7803), .B(n7804), .Z(n7800) );
  AND U7468 ( .A(n762), .B(n7805), .Z(n7804) );
  XOR U7469 ( .A(n7806), .B(n7807), .Z(n7798) );
  AND U7470 ( .A(n766), .B(n7797), .Z(n7807) );
  XNOR U7471 ( .A(n7808), .B(n7795), .Z(n7797) );
  XOR U7472 ( .A(n7809), .B(n7810), .Z(n7795) );
  AND U7473 ( .A(n789), .B(n7811), .Z(n7810) );
  IV U7474 ( .A(n7806), .Z(n7808) );
  XOR U7475 ( .A(n7812), .B(n7813), .Z(n7806) );
  AND U7476 ( .A(n773), .B(n7805), .Z(n7813) );
  XNOR U7477 ( .A(n7803), .B(n7812), .Z(n7805) );
  XNOR U7478 ( .A(n7814), .B(n7815), .Z(n7803) );
  AND U7479 ( .A(n777), .B(n7816), .Z(n7815) );
  XOR U7480 ( .A(p_input[1118]), .B(n7814), .Z(n7816) );
  XNOR U7481 ( .A(n7817), .B(n7818), .Z(n7814) );
  AND U7482 ( .A(n781), .B(n7819), .Z(n7818) );
  XOR U7483 ( .A(n7820), .B(n7821), .Z(n7812) );
  AND U7484 ( .A(n785), .B(n7811), .Z(n7821) );
  XNOR U7485 ( .A(n7822), .B(n7809), .Z(n7811) );
  XOR U7486 ( .A(n7823), .B(n7824), .Z(n7809) );
  AND U7487 ( .A(n808), .B(n7825), .Z(n7824) );
  IV U7488 ( .A(n7820), .Z(n7822) );
  XOR U7489 ( .A(n7826), .B(n7827), .Z(n7820) );
  AND U7490 ( .A(n792), .B(n7819), .Z(n7827) );
  XNOR U7491 ( .A(n7817), .B(n7826), .Z(n7819) );
  XNOR U7492 ( .A(n7828), .B(n7829), .Z(n7817) );
  AND U7493 ( .A(n796), .B(n7830), .Z(n7829) );
  XOR U7494 ( .A(p_input[1150]), .B(n7828), .Z(n7830) );
  XNOR U7495 ( .A(n7831), .B(n7832), .Z(n7828) );
  AND U7496 ( .A(n800), .B(n7833), .Z(n7832) );
  XOR U7497 ( .A(n7834), .B(n7835), .Z(n7826) );
  AND U7498 ( .A(n804), .B(n7825), .Z(n7835) );
  XNOR U7499 ( .A(n7836), .B(n7823), .Z(n7825) );
  XOR U7500 ( .A(n7837), .B(n7838), .Z(n7823) );
  AND U7501 ( .A(n827), .B(n7839), .Z(n7838) );
  IV U7502 ( .A(n7834), .Z(n7836) );
  XOR U7503 ( .A(n7840), .B(n7841), .Z(n7834) );
  AND U7504 ( .A(n811), .B(n7833), .Z(n7841) );
  XNOR U7505 ( .A(n7831), .B(n7840), .Z(n7833) );
  XNOR U7506 ( .A(n7842), .B(n7843), .Z(n7831) );
  AND U7507 ( .A(n815), .B(n7844), .Z(n7843) );
  XOR U7508 ( .A(p_input[1182]), .B(n7842), .Z(n7844) );
  XNOR U7509 ( .A(n7845), .B(n7846), .Z(n7842) );
  AND U7510 ( .A(n819), .B(n7847), .Z(n7846) );
  XOR U7511 ( .A(n7848), .B(n7849), .Z(n7840) );
  AND U7512 ( .A(n823), .B(n7839), .Z(n7849) );
  XNOR U7513 ( .A(n7850), .B(n7837), .Z(n7839) );
  XOR U7514 ( .A(n7851), .B(n7852), .Z(n7837) );
  AND U7515 ( .A(n846), .B(n7853), .Z(n7852) );
  IV U7516 ( .A(n7848), .Z(n7850) );
  XOR U7517 ( .A(n7854), .B(n7855), .Z(n7848) );
  AND U7518 ( .A(n830), .B(n7847), .Z(n7855) );
  XNOR U7519 ( .A(n7845), .B(n7854), .Z(n7847) );
  XNOR U7520 ( .A(n7856), .B(n7857), .Z(n7845) );
  AND U7521 ( .A(n834), .B(n7858), .Z(n7857) );
  XOR U7522 ( .A(p_input[1214]), .B(n7856), .Z(n7858) );
  XNOR U7523 ( .A(n7859), .B(n7860), .Z(n7856) );
  AND U7524 ( .A(n838), .B(n7861), .Z(n7860) );
  XOR U7525 ( .A(n7862), .B(n7863), .Z(n7854) );
  AND U7526 ( .A(n842), .B(n7853), .Z(n7863) );
  XNOR U7527 ( .A(n7864), .B(n7851), .Z(n7853) );
  XOR U7528 ( .A(n7865), .B(n7866), .Z(n7851) );
  AND U7529 ( .A(n865), .B(n7867), .Z(n7866) );
  IV U7530 ( .A(n7862), .Z(n7864) );
  XOR U7531 ( .A(n7868), .B(n7869), .Z(n7862) );
  AND U7532 ( .A(n849), .B(n7861), .Z(n7869) );
  XNOR U7533 ( .A(n7859), .B(n7868), .Z(n7861) );
  XNOR U7534 ( .A(n7870), .B(n7871), .Z(n7859) );
  AND U7535 ( .A(n853), .B(n7872), .Z(n7871) );
  XOR U7536 ( .A(p_input[1246]), .B(n7870), .Z(n7872) );
  XNOR U7537 ( .A(n7873), .B(n7874), .Z(n7870) );
  AND U7538 ( .A(n857), .B(n7875), .Z(n7874) );
  XOR U7539 ( .A(n7876), .B(n7877), .Z(n7868) );
  AND U7540 ( .A(n861), .B(n7867), .Z(n7877) );
  XNOR U7541 ( .A(n7878), .B(n7865), .Z(n7867) );
  XOR U7542 ( .A(n7879), .B(n7880), .Z(n7865) );
  AND U7543 ( .A(n884), .B(n7881), .Z(n7880) );
  IV U7544 ( .A(n7876), .Z(n7878) );
  XOR U7545 ( .A(n7882), .B(n7883), .Z(n7876) );
  AND U7546 ( .A(n868), .B(n7875), .Z(n7883) );
  XNOR U7547 ( .A(n7873), .B(n7882), .Z(n7875) );
  XNOR U7548 ( .A(n7884), .B(n7885), .Z(n7873) );
  AND U7549 ( .A(n872), .B(n7886), .Z(n7885) );
  XOR U7550 ( .A(p_input[1278]), .B(n7884), .Z(n7886) );
  XNOR U7551 ( .A(n7887), .B(n7888), .Z(n7884) );
  AND U7552 ( .A(n876), .B(n7889), .Z(n7888) );
  XOR U7553 ( .A(n7890), .B(n7891), .Z(n7882) );
  AND U7554 ( .A(n880), .B(n7881), .Z(n7891) );
  XNOR U7555 ( .A(n7892), .B(n7879), .Z(n7881) );
  XOR U7556 ( .A(n7893), .B(n7894), .Z(n7879) );
  AND U7557 ( .A(n903), .B(n7895), .Z(n7894) );
  IV U7558 ( .A(n7890), .Z(n7892) );
  XOR U7559 ( .A(n7896), .B(n7897), .Z(n7890) );
  AND U7560 ( .A(n887), .B(n7889), .Z(n7897) );
  XNOR U7561 ( .A(n7887), .B(n7896), .Z(n7889) );
  XNOR U7562 ( .A(n7898), .B(n7899), .Z(n7887) );
  AND U7563 ( .A(n891), .B(n7900), .Z(n7899) );
  XOR U7564 ( .A(p_input[1310]), .B(n7898), .Z(n7900) );
  XNOR U7565 ( .A(n7901), .B(n7902), .Z(n7898) );
  AND U7566 ( .A(n895), .B(n7903), .Z(n7902) );
  XOR U7567 ( .A(n7904), .B(n7905), .Z(n7896) );
  AND U7568 ( .A(n899), .B(n7895), .Z(n7905) );
  XNOR U7569 ( .A(n7906), .B(n7893), .Z(n7895) );
  XOR U7570 ( .A(n7907), .B(n7908), .Z(n7893) );
  AND U7571 ( .A(n922), .B(n7909), .Z(n7908) );
  IV U7572 ( .A(n7904), .Z(n7906) );
  XOR U7573 ( .A(n7910), .B(n7911), .Z(n7904) );
  AND U7574 ( .A(n906), .B(n7903), .Z(n7911) );
  XNOR U7575 ( .A(n7901), .B(n7910), .Z(n7903) );
  XNOR U7576 ( .A(n7912), .B(n7913), .Z(n7901) );
  AND U7577 ( .A(n910), .B(n7914), .Z(n7913) );
  XOR U7578 ( .A(p_input[1342]), .B(n7912), .Z(n7914) );
  XNOR U7579 ( .A(n7915), .B(n7916), .Z(n7912) );
  AND U7580 ( .A(n914), .B(n7917), .Z(n7916) );
  XOR U7581 ( .A(n7918), .B(n7919), .Z(n7910) );
  AND U7582 ( .A(n918), .B(n7909), .Z(n7919) );
  XNOR U7583 ( .A(n7920), .B(n7907), .Z(n7909) );
  XOR U7584 ( .A(n7921), .B(n7922), .Z(n7907) );
  AND U7585 ( .A(n941), .B(n7923), .Z(n7922) );
  IV U7586 ( .A(n7918), .Z(n7920) );
  XOR U7587 ( .A(n7924), .B(n7925), .Z(n7918) );
  AND U7588 ( .A(n925), .B(n7917), .Z(n7925) );
  XNOR U7589 ( .A(n7915), .B(n7924), .Z(n7917) );
  XNOR U7590 ( .A(n7926), .B(n7927), .Z(n7915) );
  AND U7591 ( .A(n929), .B(n7928), .Z(n7927) );
  XOR U7592 ( .A(p_input[1374]), .B(n7926), .Z(n7928) );
  XNOR U7593 ( .A(n7929), .B(n7930), .Z(n7926) );
  AND U7594 ( .A(n933), .B(n7931), .Z(n7930) );
  XOR U7595 ( .A(n7932), .B(n7933), .Z(n7924) );
  AND U7596 ( .A(n937), .B(n7923), .Z(n7933) );
  XNOR U7597 ( .A(n7934), .B(n7921), .Z(n7923) );
  XOR U7598 ( .A(n7935), .B(n7936), .Z(n7921) );
  AND U7599 ( .A(n960), .B(n7937), .Z(n7936) );
  IV U7600 ( .A(n7932), .Z(n7934) );
  XOR U7601 ( .A(n7938), .B(n7939), .Z(n7932) );
  AND U7602 ( .A(n944), .B(n7931), .Z(n7939) );
  XNOR U7603 ( .A(n7929), .B(n7938), .Z(n7931) );
  XNOR U7604 ( .A(n7940), .B(n7941), .Z(n7929) );
  AND U7605 ( .A(n948), .B(n7942), .Z(n7941) );
  XOR U7606 ( .A(p_input[1406]), .B(n7940), .Z(n7942) );
  XNOR U7607 ( .A(n7943), .B(n7944), .Z(n7940) );
  AND U7608 ( .A(n952), .B(n7945), .Z(n7944) );
  XOR U7609 ( .A(n7946), .B(n7947), .Z(n7938) );
  AND U7610 ( .A(n956), .B(n7937), .Z(n7947) );
  XNOR U7611 ( .A(n7948), .B(n7935), .Z(n7937) );
  XOR U7612 ( .A(n7949), .B(n7950), .Z(n7935) );
  AND U7613 ( .A(n979), .B(n7951), .Z(n7950) );
  IV U7614 ( .A(n7946), .Z(n7948) );
  XOR U7615 ( .A(n7952), .B(n7953), .Z(n7946) );
  AND U7616 ( .A(n963), .B(n7945), .Z(n7953) );
  XNOR U7617 ( .A(n7943), .B(n7952), .Z(n7945) );
  XNOR U7618 ( .A(n7954), .B(n7955), .Z(n7943) );
  AND U7619 ( .A(n967), .B(n7956), .Z(n7955) );
  XOR U7620 ( .A(p_input[1438]), .B(n7954), .Z(n7956) );
  XNOR U7621 ( .A(n7957), .B(n7958), .Z(n7954) );
  AND U7622 ( .A(n971), .B(n7959), .Z(n7958) );
  XOR U7623 ( .A(n7960), .B(n7961), .Z(n7952) );
  AND U7624 ( .A(n975), .B(n7951), .Z(n7961) );
  XNOR U7625 ( .A(n7962), .B(n7949), .Z(n7951) );
  XOR U7626 ( .A(n7963), .B(n7964), .Z(n7949) );
  AND U7627 ( .A(n998), .B(n7965), .Z(n7964) );
  IV U7628 ( .A(n7960), .Z(n7962) );
  XOR U7629 ( .A(n7966), .B(n7967), .Z(n7960) );
  AND U7630 ( .A(n982), .B(n7959), .Z(n7967) );
  XNOR U7631 ( .A(n7957), .B(n7966), .Z(n7959) );
  XNOR U7632 ( .A(n7968), .B(n7969), .Z(n7957) );
  AND U7633 ( .A(n986), .B(n7970), .Z(n7969) );
  XOR U7634 ( .A(p_input[1470]), .B(n7968), .Z(n7970) );
  XNOR U7635 ( .A(n7971), .B(n7972), .Z(n7968) );
  AND U7636 ( .A(n990), .B(n7973), .Z(n7972) );
  XOR U7637 ( .A(n7974), .B(n7975), .Z(n7966) );
  AND U7638 ( .A(n994), .B(n7965), .Z(n7975) );
  XNOR U7639 ( .A(n7976), .B(n7963), .Z(n7965) );
  XOR U7640 ( .A(n7977), .B(n7978), .Z(n7963) );
  AND U7641 ( .A(n1017), .B(n7979), .Z(n7978) );
  IV U7642 ( .A(n7974), .Z(n7976) );
  XOR U7643 ( .A(n7980), .B(n7981), .Z(n7974) );
  AND U7644 ( .A(n1001), .B(n7973), .Z(n7981) );
  XNOR U7645 ( .A(n7971), .B(n7980), .Z(n7973) );
  XNOR U7646 ( .A(n7982), .B(n7983), .Z(n7971) );
  AND U7647 ( .A(n1005), .B(n7984), .Z(n7983) );
  XOR U7648 ( .A(p_input[1502]), .B(n7982), .Z(n7984) );
  XNOR U7649 ( .A(n7985), .B(n7986), .Z(n7982) );
  AND U7650 ( .A(n1009), .B(n7987), .Z(n7986) );
  XOR U7651 ( .A(n7988), .B(n7989), .Z(n7980) );
  AND U7652 ( .A(n1013), .B(n7979), .Z(n7989) );
  XNOR U7653 ( .A(n7990), .B(n7977), .Z(n7979) );
  XOR U7654 ( .A(n7991), .B(n7992), .Z(n7977) );
  AND U7655 ( .A(n1036), .B(n7993), .Z(n7992) );
  IV U7656 ( .A(n7988), .Z(n7990) );
  XOR U7657 ( .A(n7994), .B(n7995), .Z(n7988) );
  AND U7658 ( .A(n1020), .B(n7987), .Z(n7995) );
  XNOR U7659 ( .A(n7985), .B(n7994), .Z(n7987) );
  XNOR U7660 ( .A(n7996), .B(n7997), .Z(n7985) );
  AND U7661 ( .A(n1024), .B(n7998), .Z(n7997) );
  XOR U7662 ( .A(p_input[1534]), .B(n7996), .Z(n7998) );
  XNOR U7663 ( .A(n7999), .B(n8000), .Z(n7996) );
  AND U7664 ( .A(n1028), .B(n8001), .Z(n8000) );
  XOR U7665 ( .A(n8002), .B(n8003), .Z(n7994) );
  AND U7666 ( .A(n1032), .B(n7993), .Z(n8003) );
  XNOR U7667 ( .A(n8004), .B(n7991), .Z(n7993) );
  XOR U7668 ( .A(n8005), .B(n8006), .Z(n7991) );
  AND U7669 ( .A(n1055), .B(n8007), .Z(n8006) );
  IV U7670 ( .A(n8002), .Z(n8004) );
  XOR U7671 ( .A(n8008), .B(n8009), .Z(n8002) );
  AND U7672 ( .A(n1039), .B(n8001), .Z(n8009) );
  XNOR U7673 ( .A(n7999), .B(n8008), .Z(n8001) );
  XNOR U7674 ( .A(n8010), .B(n8011), .Z(n7999) );
  AND U7675 ( .A(n1043), .B(n8012), .Z(n8011) );
  XOR U7676 ( .A(p_input[1566]), .B(n8010), .Z(n8012) );
  XNOR U7677 ( .A(n8013), .B(n8014), .Z(n8010) );
  AND U7678 ( .A(n1047), .B(n8015), .Z(n8014) );
  XOR U7679 ( .A(n8016), .B(n8017), .Z(n8008) );
  AND U7680 ( .A(n1051), .B(n8007), .Z(n8017) );
  XNOR U7681 ( .A(n8018), .B(n8005), .Z(n8007) );
  XOR U7682 ( .A(n8019), .B(n8020), .Z(n8005) );
  AND U7683 ( .A(n1074), .B(n8021), .Z(n8020) );
  IV U7684 ( .A(n8016), .Z(n8018) );
  XOR U7685 ( .A(n8022), .B(n8023), .Z(n8016) );
  AND U7686 ( .A(n1058), .B(n8015), .Z(n8023) );
  XNOR U7687 ( .A(n8013), .B(n8022), .Z(n8015) );
  XNOR U7688 ( .A(n8024), .B(n8025), .Z(n8013) );
  AND U7689 ( .A(n1062), .B(n8026), .Z(n8025) );
  XOR U7690 ( .A(p_input[1598]), .B(n8024), .Z(n8026) );
  XNOR U7691 ( .A(n8027), .B(n8028), .Z(n8024) );
  AND U7692 ( .A(n1066), .B(n8029), .Z(n8028) );
  XOR U7693 ( .A(n8030), .B(n8031), .Z(n8022) );
  AND U7694 ( .A(n1070), .B(n8021), .Z(n8031) );
  XNOR U7695 ( .A(n8032), .B(n8019), .Z(n8021) );
  XOR U7696 ( .A(n8033), .B(n8034), .Z(n8019) );
  AND U7697 ( .A(n1093), .B(n8035), .Z(n8034) );
  IV U7698 ( .A(n8030), .Z(n8032) );
  XOR U7699 ( .A(n8036), .B(n8037), .Z(n8030) );
  AND U7700 ( .A(n1077), .B(n8029), .Z(n8037) );
  XNOR U7701 ( .A(n8027), .B(n8036), .Z(n8029) );
  XNOR U7702 ( .A(n8038), .B(n8039), .Z(n8027) );
  AND U7703 ( .A(n1081), .B(n8040), .Z(n8039) );
  XOR U7704 ( .A(p_input[1630]), .B(n8038), .Z(n8040) );
  XNOR U7705 ( .A(n8041), .B(n8042), .Z(n8038) );
  AND U7706 ( .A(n1085), .B(n8043), .Z(n8042) );
  XOR U7707 ( .A(n8044), .B(n8045), .Z(n8036) );
  AND U7708 ( .A(n1089), .B(n8035), .Z(n8045) );
  XNOR U7709 ( .A(n8046), .B(n8033), .Z(n8035) );
  XOR U7710 ( .A(n8047), .B(n8048), .Z(n8033) );
  AND U7711 ( .A(n1112), .B(n8049), .Z(n8048) );
  IV U7712 ( .A(n8044), .Z(n8046) );
  XOR U7713 ( .A(n8050), .B(n8051), .Z(n8044) );
  AND U7714 ( .A(n1096), .B(n8043), .Z(n8051) );
  XNOR U7715 ( .A(n8041), .B(n8050), .Z(n8043) );
  XNOR U7716 ( .A(n8052), .B(n8053), .Z(n8041) );
  AND U7717 ( .A(n1100), .B(n8054), .Z(n8053) );
  XOR U7718 ( .A(p_input[1662]), .B(n8052), .Z(n8054) );
  XNOR U7719 ( .A(n8055), .B(n8056), .Z(n8052) );
  AND U7720 ( .A(n1104), .B(n8057), .Z(n8056) );
  XOR U7721 ( .A(n8058), .B(n8059), .Z(n8050) );
  AND U7722 ( .A(n1108), .B(n8049), .Z(n8059) );
  XNOR U7723 ( .A(n8060), .B(n8047), .Z(n8049) );
  XOR U7724 ( .A(n8061), .B(n8062), .Z(n8047) );
  AND U7725 ( .A(n1131), .B(n8063), .Z(n8062) );
  IV U7726 ( .A(n8058), .Z(n8060) );
  XOR U7727 ( .A(n8064), .B(n8065), .Z(n8058) );
  AND U7728 ( .A(n1115), .B(n8057), .Z(n8065) );
  XNOR U7729 ( .A(n8055), .B(n8064), .Z(n8057) );
  XNOR U7730 ( .A(n8066), .B(n8067), .Z(n8055) );
  AND U7731 ( .A(n1119), .B(n8068), .Z(n8067) );
  XOR U7732 ( .A(p_input[1694]), .B(n8066), .Z(n8068) );
  XNOR U7733 ( .A(n8069), .B(n8070), .Z(n8066) );
  AND U7734 ( .A(n1123), .B(n8071), .Z(n8070) );
  XOR U7735 ( .A(n8072), .B(n8073), .Z(n8064) );
  AND U7736 ( .A(n1127), .B(n8063), .Z(n8073) );
  XNOR U7737 ( .A(n8074), .B(n8061), .Z(n8063) );
  XOR U7738 ( .A(n8075), .B(n8076), .Z(n8061) );
  AND U7739 ( .A(n1150), .B(n8077), .Z(n8076) );
  IV U7740 ( .A(n8072), .Z(n8074) );
  XOR U7741 ( .A(n8078), .B(n8079), .Z(n8072) );
  AND U7742 ( .A(n1134), .B(n8071), .Z(n8079) );
  XNOR U7743 ( .A(n8069), .B(n8078), .Z(n8071) );
  XNOR U7744 ( .A(n8080), .B(n8081), .Z(n8069) );
  AND U7745 ( .A(n1138), .B(n8082), .Z(n8081) );
  XOR U7746 ( .A(p_input[1726]), .B(n8080), .Z(n8082) );
  XNOR U7747 ( .A(n8083), .B(n8084), .Z(n8080) );
  AND U7748 ( .A(n1142), .B(n8085), .Z(n8084) );
  XOR U7749 ( .A(n8086), .B(n8087), .Z(n8078) );
  AND U7750 ( .A(n1146), .B(n8077), .Z(n8087) );
  XNOR U7751 ( .A(n8088), .B(n8075), .Z(n8077) );
  XOR U7752 ( .A(n8089), .B(n8090), .Z(n8075) );
  AND U7753 ( .A(n1169), .B(n8091), .Z(n8090) );
  IV U7754 ( .A(n8086), .Z(n8088) );
  XOR U7755 ( .A(n8092), .B(n8093), .Z(n8086) );
  AND U7756 ( .A(n1153), .B(n8085), .Z(n8093) );
  XNOR U7757 ( .A(n8083), .B(n8092), .Z(n8085) );
  XNOR U7758 ( .A(n8094), .B(n8095), .Z(n8083) );
  AND U7759 ( .A(n1157), .B(n8096), .Z(n8095) );
  XOR U7760 ( .A(p_input[1758]), .B(n8094), .Z(n8096) );
  XNOR U7761 ( .A(n8097), .B(n8098), .Z(n8094) );
  AND U7762 ( .A(n1161), .B(n8099), .Z(n8098) );
  XOR U7763 ( .A(n8100), .B(n8101), .Z(n8092) );
  AND U7764 ( .A(n1165), .B(n8091), .Z(n8101) );
  XNOR U7765 ( .A(n8102), .B(n8089), .Z(n8091) );
  XOR U7766 ( .A(n8103), .B(n8104), .Z(n8089) );
  AND U7767 ( .A(n1188), .B(n8105), .Z(n8104) );
  IV U7768 ( .A(n8100), .Z(n8102) );
  XOR U7769 ( .A(n8106), .B(n8107), .Z(n8100) );
  AND U7770 ( .A(n1172), .B(n8099), .Z(n8107) );
  XNOR U7771 ( .A(n8097), .B(n8106), .Z(n8099) );
  XNOR U7772 ( .A(n8108), .B(n8109), .Z(n8097) );
  AND U7773 ( .A(n1176), .B(n8110), .Z(n8109) );
  XOR U7774 ( .A(p_input[1790]), .B(n8108), .Z(n8110) );
  XNOR U7775 ( .A(n8111), .B(n8112), .Z(n8108) );
  AND U7776 ( .A(n1180), .B(n8113), .Z(n8112) );
  XOR U7777 ( .A(n8114), .B(n8115), .Z(n8106) );
  AND U7778 ( .A(n1184), .B(n8105), .Z(n8115) );
  XNOR U7779 ( .A(n8116), .B(n8103), .Z(n8105) );
  XOR U7780 ( .A(n8117), .B(n8118), .Z(n8103) );
  AND U7781 ( .A(n1207), .B(n8119), .Z(n8118) );
  IV U7782 ( .A(n8114), .Z(n8116) );
  XOR U7783 ( .A(n8120), .B(n8121), .Z(n8114) );
  AND U7784 ( .A(n1191), .B(n8113), .Z(n8121) );
  XNOR U7785 ( .A(n8111), .B(n8120), .Z(n8113) );
  XNOR U7786 ( .A(n8122), .B(n8123), .Z(n8111) );
  AND U7787 ( .A(n1195), .B(n8124), .Z(n8123) );
  XOR U7788 ( .A(p_input[1822]), .B(n8122), .Z(n8124) );
  XNOR U7789 ( .A(n8125), .B(n8126), .Z(n8122) );
  AND U7790 ( .A(n1199), .B(n8127), .Z(n8126) );
  XOR U7791 ( .A(n8128), .B(n8129), .Z(n8120) );
  AND U7792 ( .A(n1203), .B(n8119), .Z(n8129) );
  XNOR U7793 ( .A(n8130), .B(n8117), .Z(n8119) );
  XOR U7794 ( .A(n8131), .B(n8132), .Z(n8117) );
  AND U7795 ( .A(n1226), .B(n8133), .Z(n8132) );
  IV U7796 ( .A(n8128), .Z(n8130) );
  XOR U7797 ( .A(n8134), .B(n8135), .Z(n8128) );
  AND U7798 ( .A(n1210), .B(n8127), .Z(n8135) );
  XNOR U7799 ( .A(n8125), .B(n8134), .Z(n8127) );
  XNOR U7800 ( .A(n8136), .B(n8137), .Z(n8125) );
  AND U7801 ( .A(n1214), .B(n8138), .Z(n8137) );
  XOR U7802 ( .A(p_input[1854]), .B(n8136), .Z(n8138) );
  XNOR U7803 ( .A(n8139), .B(n8140), .Z(n8136) );
  AND U7804 ( .A(n1218), .B(n8141), .Z(n8140) );
  XOR U7805 ( .A(n8142), .B(n8143), .Z(n8134) );
  AND U7806 ( .A(n1222), .B(n8133), .Z(n8143) );
  XNOR U7807 ( .A(n8144), .B(n8131), .Z(n8133) );
  XOR U7808 ( .A(n8145), .B(n8146), .Z(n8131) );
  AND U7809 ( .A(n1245), .B(n8147), .Z(n8146) );
  IV U7810 ( .A(n8142), .Z(n8144) );
  XOR U7811 ( .A(n8148), .B(n8149), .Z(n8142) );
  AND U7812 ( .A(n1229), .B(n8141), .Z(n8149) );
  XNOR U7813 ( .A(n8139), .B(n8148), .Z(n8141) );
  XNOR U7814 ( .A(n8150), .B(n8151), .Z(n8139) );
  AND U7815 ( .A(n1233), .B(n8152), .Z(n8151) );
  XOR U7816 ( .A(p_input[1886]), .B(n8150), .Z(n8152) );
  XNOR U7817 ( .A(n8153), .B(n8154), .Z(n8150) );
  AND U7818 ( .A(n1237), .B(n8155), .Z(n8154) );
  XOR U7819 ( .A(n8156), .B(n8157), .Z(n8148) );
  AND U7820 ( .A(n1241), .B(n8147), .Z(n8157) );
  XNOR U7821 ( .A(n8158), .B(n8145), .Z(n8147) );
  XOR U7822 ( .A(n8159), .B(n8160), .Z(n8145) );
  AND U7823 ( .A(n1264), .B(n8161), .Z(n8160) );
  IV U7824 ( .A(n8156), .Z(n8158) );
  XOR U7825 ( .A(n8162), .B(n8163), .Z(n8156) );
  AND U7826 ( .A(n1248), .B(n8155), .Z(n8163) );
  XNOR U7827 ( .A(n8153), .B(n8162), .Z(n8155) );
  XNOR U7828 ( .A(n8164), .B(n8165), .Z(n8153) );
  AND U7829 ( .A(n1252), .B(n8166), .Z(n8165) );
  XOR U7830 ( .A(p_input[1918]), .B(n8164), .Z(n8166) );
  XNOR U7831 ( .A(n8167), .B(n8168), .Z(n8164) );
  AND U7832 ( .A(n1256), .B(n8169), .Z(n8168) );
  XOR U7833 ( .A(n8170), .B(n8171), .Z(n8162) );
  AND U7834 ( .A(n1260), .B(n8161), .Z(n8171) );
  XNOR U7835 ( .A(n8172), .B(n8159), .Z(n8161) );
  XOR U7836 ( .A(n8173), .B(n8174), .Z(n8159) );
  AND U7837 ( .A(n1282), .B(n8175), .Z(n8174) );
  IV U7838 ( .A(n8170), .Z(n8172) );
  XOR U7839 ( .A(n8176), .B(n8177), .Z(n8170) );
  AND U7840 ( .A(n1267), .B(n8169), .Z(n8177) );
  XNOR U7841 ( .A(n8167), .B(n8176), .Z(n8169) );
  XNOR U7842 ( .A(n8178), .B(n8179), .Z(n8167) );
  AND U7843 ( .A(n1271), .B(n8180), .Z(n8179) );
  XOR U7844 ( .A(p_input[1950]), .B(n8178), .Z(n8180) );
  XOR U7845 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][30] ), .B(n8181), 
        .Z(n8178) );
  AND U7846 ( .A(n1274), .B(n8182), .Z(n8181) );
  XOR U7847 ( .A(n8183), .B(n8184), .Z(n8176) );
  AND U7848 ( .A(n1278), .B(n8175), .Z(n8184) );
  XNOR U7849 ( .A(n8185), .B(n8173), .Z(n8175) );
  XOR U7850 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n8186), .Z(n8173) );
  AND U7851 ( .A(n1290), .B(n8187), .Z(n8186) );
  IV U7852 ( .A(n8183), .Z(n8185) );
  XOR U7853 ( .A(n8188), .B(n8189), .Z(n8183) );
  AND U7854 ( .A(n1285), .B(n8182), .Z(n8189) );
  XOR U7855 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][30] ), .B(n8188), 
        .Z(n8182) );
  XOR U7856 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .B(n8190), 
        .Z(n8188) );
  AND U7857 ( .A(n1287), .B(n8187), .Z(n8190) );
  XOR U7858 ( .A(n8191), .B(n8192), .Z(n8187) );
  IV U7859 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .Z(n8192) );
  IV U7860 ( .A(\knn_comb_/min_val_out[0][30] ), .Z(n8191) );
  XOR U7861 ( .A(n6463), .B(n8193), .Z(o[2]) );
  AND U7862 ( .A(n122), .B(n8194), .Z(n6463) );
  XOR U7863 ( .A(n6464), .B(n8193), .Z(n8194) );
  XOR U7864 ( .A(n8195), .B(n8196), .Z(n8193) );
  AND U7865 ( .A(n142), .B(n8197), .Z(n8196) );
  XOR U7866 ( .A(n8198), .B(n67), .Z(n6464) );
  AND U7867 ( .A(n125), .B(n8199), .Z(n67) );
  XOR U7868 ( .A(n68), .B(n8198), .Z(n8199) );
  XOR U7869 ( .A(n8200), .B(n8201), .Z(n68) );
  AND U7870 ( .A(n130), .B(n8202), .Z(n8201) );
  XOR U7871 ( .A(p_input[2]), .B(n8200), .Z(n8202) );
  XNOR U7872 ( .A(n8203), .B(n8204), .Z(n8200) );
  AND U7873 ( .A(n134), .B(n8205), .Z(n8204) );
  XOR U7874 ( .A(n8206), .B(n8207), .Z(n8198) );
  AND U7875 ( .A(n138), .B(n8197), .Z(n8207) );
  XNOR U7876 ( .A(n8208), .B(n8195), .Z(n8197) );
  XOR U7877 ( .A(n8209), .B(n8210), .Z(n8195) );
  AND U7878 ( .A(n162), .B(n8211), .Z(n8210) );
  IV U7879 ( .A(n8206), .Z(n8208) );
  XOR U7880 ( .A(n8212), .B(n8213), .Z(n8206) );
  AND U7881 ( .A(n146), .B(n8205), .Z(n8213) );
  XNOR U7882 ( .A(n8203), .B(n8212), .Z(n8205) );
  XNOR U7883 ( .A(n8214), .B(n8215), .Z(n8203) );
  AND U7884 ( .A(n150), .B(n8216), .Z(n8215) );
  XOR U7885 ( .A(p_input[34]), .B(n8214), .Z(n8216) );
  XNOR U7886 ( .A(n8217), .B(n8218), .Z(n8214) );
  AND U7887 ( .A(n154), .B(n8219), .Z(n8218) );
  XOR U7888 ( .A(n8220), .B(n8221), .Z(n8212) );
  AND U7889 ( .A(n158), .B(n8211), .Z(n8221) );
  XNOR U7890 ( .A(n8222), .B(n8209), .Z(n8211) );
  XOR U7891 ( .A(n8223), .B(n8224), .Z(n8209) );
  AND U7892 ( .A(n181), .B(n8225), .Z(n8224) );
  IV U7893 ( .A(n8220), .Z(n8222) );
  XOR U7894 ( .A(n8226), .B(n8227), .Z(n8220) );
  AND U7895 ( .A(n165), .B(n8219), .Z(n8227) );
  XNOR U7896 ( .A(n8217), .B(n8226), .Z(n8219) );
  XNOR U7897 ( .A(n8228), .B(n8229), .Z(n8217) );
  AND U7898 ( .A(n169), .B(n8230), .Z(n8229) );
  XOR U7899 ( .A(p_input[66]), .B(n8228), .Z(n8230) );
  XNOR U7900 ( .A(n8231), .B(n8232), .Z(n8228) );
  AND U7901 ( .A(n173), .B(n8233), .Z(n8232) );
  XOR U7902 ( .A(n8234), .B(n8235), .Z(n8226) );
  AND U7903 ( .A(n177), .B(n8225), .Z(n8235) );
  XNOR U7904 ( .A(n8236), .B(n8223), .Z(n8225) );
  XOR U7905 ( .A(n8237), .B(n8238), .Z(n8223) );
  AND U7906 ( .A(n200), .B(n8239), .Z(n8238) );
  IV U7907 ( .A(n8234), .Z(n8236) );
  XOR U7908 ( .A(n8240), .B(n8241), .Z(n8234) );
  AND U7909 ( .A(n184), .B(n8233), .Z(n8241) );
  XNOR U7910 ( .A(n8231), .B(n8240), .Z(n8233) );
  XNOR U7911 ( .A(n8242), .B(n8243), .Z(n8231) );
  AND U7912 ( .A(n188), .B(n8244), .Z(n8243) );
  XOR U7913 ( .A(p_input[98]), .B(n8242), .Z(n8244) );
  XNOR U7914 ( .A(n8245), .B(n8246), .Z(n8242) );
  AND U7915 ( .A(n192), .B(n8247), .Z(n8246) );
  XOR U7916 ( .A(n8248), .B(n8249), .Z(n8240) );
  AND U7917 ( .A(n196), .B(n8239), .Z(n8249) );
  XNOR U7918 ( .A(n8250), .B(n8237), .Z(n8239) );
  XOR U7919 ( .A(n8251), .B(n8252), .Z(n8237) );
  AND U7920 ( .A(n219), .B(n8253), .Z(n8252) );
  IV U7921 ( .A(n8248), .Z(n8250) );
  XOR U7922 ( .A(n8254), .B(n8255), .Z(n8248) );
  AND U7923 ( .A(n203), .B(n8247), .Z(n8255) );
  XNOR U7924 ( .A(n8245), .B(n8254), .Z(n8247) );
  XNOR U7925 ( .A(n8256), .B(n8257), .Z(n8245) );
  AND U7926 ( .A(n207), .B(n8258), .Z(n8257) );
  XOR U7927 ( .A(p_input[130]), .B(n8256), .Z(n8258) );
  XNOR U7928 ( .A(n8259), .B(n8260), .Z(n8256) );
  AND U7929 ( .A(n211), .B(n8261), .Z(n8260) );
  XOR U7930 ( .A(n8262), .B(n8263), .Z(n8254) );
  AND U7931 ( .A(n215), .B(n8253), .Z(n8263) );
  XNOR U7932 ( .A(n8264), .B(n8251), .Z(n8253) );
  XOR U7933 ( .A(n8265), .B(n8266), .Z(n8251) );
  AND U7934 ( .A(n238), .B(n8267), .Z(n8266) );
  IV U7935 ( .A(n8262), .Z(n8264) );
  XOR U7936 ( .A(n8268), .B(n8269), .Z(n8262) );
  AND U7937 ( .A(n222), .B(n8261), .Z(n8269) );
  XNOR U7938 ( .A(n8259), .B(n8268), .Z(n8261) );
  XNOR U7939 ( .A(n8270), .B(n8271), .Z(n8259) );
  AND U7940 ( .A(n226), .B(n8272), .Z(n8271) );
  XOR U7941 ( .A(p_input[162]), .B(n8270), .Z(n8272) );
  XNOR U7942 ( .A(n8273), .B(n8274), .Z(n8270) );
  AND U7943 ( .A(n230), .B(n8275), .Z(n8274) );
  XOR U7944 ( .A(n8276), .B(n8277), .Z(n8268) );
  AND U7945 ( .A(n234), .B(n8267), .Z(n8277) );
  XNOR U7946 ( .A(n8278), .B(n8265), .Z(n8267) );
  XOR U7947 ( .A(n8279), .B(n8280), .Z(n8265) );
  AND U7948 ( .A(n257), .B(n8281), .Z(n8280) );
  IV U7949 ( .A(n8276), .Z(n8278) );
  XOR U7950 ( .A(n8282), .B(n8283), .Z(n8276) );
  AND U7951 ( .A(n241), .B(n8275), .Z(n8283) );
  XNOR U7952 ( .A(n8273), .B(n8282), .Z(n8275) );
  XNOR U7953 ( .A(n8284), .B(n8285), .Z(n8273) );
  AND U7954 ( .A(n245), .B(n8286), .Z(n8285) );
  XOR U7955 ( .A(p_input[194]), .B(n8284), .Z(n8286) );
  XNOR U7956 ( .A(n8287), .B(n8288), .Z(n8284) );
  AND U7957 ( .A(n249), .B(n8289), .Z(n8288) );
  XOR U7958 ( .A(n8290), .B(n8291), .Z(n8282) );
  AND U7959 ( .A(n253), .B(n8281), .Z(n8291) );
  XNOR U7960 ( .A(n8292), .B(n8279), .Z(n8281) );
  XOR U7961 ( .A(n8293), .B(n8294), .Z(n8279) );
  AND U7962 ( .A(n276), .B(n8295), .Z(n8294) );
  IV U7963 ( .A(n8290), .Z(n8292) );
  XOR U7964 ( .A(n8296), .B(n8297), .Z(n8290) );
  AND U7965 ( .A(n260), .B(n8289), .Z(n8297) );
  XNOR U7966 ( .A(n8287), .B(n8296), .Z(n8289) );
  XNOR U7967 ( .A(n8298), .B(n8299), .Z(n8287) );
  AND U7968 ( .A(n264), .B(n8300), .Z(n8299) );
  XOR U7969 ( .A(p_input[226]), .B(n8298), .Z(n8300) );
  XNOR U7970 ( .A(n8301), .B(n8302), .Z(n8298) );
  AND U7971 ( .A(n268), .B(n8303), .Z(n8302) );
  XOR U7972 ( .A(n8304), .B(n8305), .Z(n8296) );
  AND U7973 ( .A(n272), .B(n8295), .Z(n8305) );
  XNOR U7974 ( .A(n8306), .B(n8293), .Z(n8295) );
  XOR U7975 ( .A(n8307), .B(n8308), .Z(n8293) );
  AND U7976 ( .A(n295), .B(n8309), .Z(n8308) );
  IV U7977 ( .A(n8304), .Z(n8306) );
  XOR U7978 ( .A(n8310), .B(n8311), .Z(n8304) );
  AND U7979 ( .A(n279), .B(n8303), .Z(n8311) );
  XNOR U7980 ( .A(n8301), .B(n8310), .Z(n8303) );
  XNOR U7981 ( .A(n8312), .B(n8313), .Z(n8301) );
  AND U7982 ( .A(n283), .B(n8314), .Z(n8313) );
  XOR U7983 ( .A(p_input[258]), .B(n8312), .Z(n8314) );
  XNOR U7984 ( .A(n8315), .B(n8316), .Z(n8312) );
  AND U7985 ( .A(n287), .B(n8317), .Z(n8316) );
  XOR U7986 ( .A(n8318), .B(n8319), .Z(n8310) );
  AND U7987 ( .A(n291), .B(n8309), .Z(n8319) );
  XNOR U7988 ( .A(n8320), .B(n8307), .Z(n8309) );
  XOR U7989 ( .A(n8321), .B(n8322), .Z(n8307) );
  AND U7990 ( .A(n314), .B(n8323), .Z(n8322) );
  IV U7991 ( .A(n8318), .Z(n8320) );
  XOR U7992 ( .A(n8324), .B(n8325), .Z(n8318) );
  AND U7993 ( .A(n298), .B(n8317), .Z(n8325) );
  XNOR U7994 ( .A(n8315), .B(n8324), .Z(n8317) );
  XNOR U7995 ( .A(n8326), .B(n8327), .Z(n8315) );
  AND U7996 ( .A(n302), .B(n8328), .Z(n8327) );
  XOR U7997 ( .A(p_input[290]), .B(n8326), .Z(n8328) );
  XNOR U7998 ( .A(n8329), .B(n8330), .Z(n8326) );
  AND U7999 ( .A(n306), .B(n8331), .Z(n8330) );
  XOR U8000 ( .A(n8332), .B(n8333), .Z(n8324) );
  AND U8001 ( .A(n310), .B(n8323), .Z(n8333) );
  XNOR U8002 ( .A(n8334), .B(n8321), .Z(n8323) );
  XOR U8003 ( .A(n8335), .B(n8336), .Z(n8321) );
  AND U8004 ( .A(n333), .B(n8337), .Z(n8336) );
  IV U8005 ( .A(n8332), .Z(n8334) );
  XOR U8006 ( .A(n8338), .B(n8339), .Z(n8332) );
  AND U8007 ( .A(n317), .B(n8331), .Z(n8339) );
  XNOR U8008 ( .A(n8329), .B(n8338), .Z(n8331) );
  XNOR U8009 ( .A(n8340), .B(n8341), .Z(n8329) );
  AND U8010 ( .A(n321), .B(n8342), .Z(n8341) );
  XOR U8011 ( .A(p_input[322]), .B(n8340), .Z(n8342) );
  XNOR U8012 ( .A(n8343), .B(n8344), .Z(n8340) );
  AND U8013 ( .A(n325), .B(n8345), .Z(n8344) );
  XOR U8014 ( .A(n8346), .B(n8347), .Z(n8338) );
  AND U8015 ( .A(n329), .B(n8337), .Z(n8347) );
  XNOR U8016 ( .A(n8348), .B(n8335), .Z(n8337) );
  XOR U8017 ( .A(n8349), .B(n8350), .Z(n8335) );
  AND U8018 ( .A(n352), .B(n8351), .Z(n8350) );
  IV U8019 ( .A(n8346), .Z(n8348) );
  XOR U8020 ( .A(n8352), .B(n8353), .Z(n8346) );
  AND U8021 ( .A(n336), .B(n8345), .Z(n8353) );
  XNOR U8022 ( .A(n8343), .B(n8352), .Z(n8345) );
  XNOR U8023 ( .A(n8354), .B(n8355), .Z(n8343) );
  AND U8024 ( .A(n340), .B(n8356), .Z(n8355) );
  XOR U8025 ( .A(p_input[354]), .B(n8354), .Z(n8356) );
  XNOR U8026 ( .A(n8357), .B(n8358), .Z(n8354) );
  AND U8027 ( .A(n344), .B(n8359), .Z(n8358) );
  XOR U8028 ( .A(n8360), .B(n8361), .Z(n8352) );
  AND U8029 ( .A(n348), .B(n8351), .Z(n8361) );
  XNOR U8030 ( .A(n8362), .B(n8349), .Z(n8351) );
  XOR U8031 ( .A(n8363), .B(n8364), .Z(n8349) );
  AND U8032 ( .A(n371), .B(n8365), .Z(n8364) );
  IV U8033 ( .A(n8360), .Z(n8362) );
  XOR U8034 ( .A(n8366), .B(n8367), .Z(n8360) );
  AND U8035 ( .A(n355), .B(n8359), .Z(n8367) );
  XNOR U8036 ( .A(n8357), .B(n8366), .Z(n8359) );
  XNOR U8037 ( .A(n8368), .B(n8369), .Z(n8357) );
  AND U8038 ( .A(n359), .B(n8370), .Z(n8369) );
  XOR U8039 ( .A(p_input[386]), .B(n8368), .Z(n8370) );
  XNOR U8040 ( .A(n8371), .B(n8372), .Z(n8368) );
  AND U8041 ( .A(n363), .B(n8373), .Z(n8372) );
  XOR U8042 ( .A(n8374), .B(n8375), .Z(n8366) );
  AND U8043 ( .A(n367), .B(n8365), .Z(n8375) );
  XNOR U8044 ( .A(n8376), .B(n8363), .Z(n8365) );
  XOR U8045 ( .A(n8377), .B(n8378), .Z(n8363) );
  AND U8046 ( .A(n390), .B(n8379), .Z(n8378) );
  IV U8047 ( .A(n8374), .Z(n8376) );
  XOR U8048 ( .A(n8380), .B(n8381), .Z(n8374) );
  AND U8049 ( .A(n374), .B(n8373), .Z(n8381) );
  XNOR U8050 ( .A(n8371), .B(n8380), .Z(n8373) );
  XNOR U8051 ( .A(n8382), .B(n8383), .Z(n8371) );
  AND U8052 ( .A(n378), .B(n8384), .Z(n8383) );
  XOR U8053 ( .A(p_input[418]), .B(n8382), .Z(n8384) );
  XNOR U8054 ( .A(n8385), .B(n8386), .Z(n8382) );
  AND U8055 ( .A(n382), .B(n8387), .Z(n8386) );
  XOR U8056 ( .A(n8388), .B(n8389), .Z(n8380) );
  AND U8057 ( .A(n386), .B(n8379), .Z(n8389) );
  XNOR U8058 ( .A(n8390), .B(n8377), .Z(n8379) );
  XOR U8059 ( .A(n8391), .B(n8392), .Z(n8377) );
  AND U8060 ( .A(n409), .B(n8393), .Z(n8392) );
  IV U8061 ( .A(n8388), .Z(n8390) );
  XOR U8062 ( .A(n8394), .B(n8395), .Z(n8388) );
  AND U8063 ( .A(n393), .B(n8387), .Z(n8395) );
  XNOR U8064 ( .A(n8385), .B(n8394), .Z(n8387) );
  XNOR U8065 ( .A(n8396), .B(n8397), .Z(n8385) );
  AND U8066 ( .A(n397), .B(n8398), .Z(n8397) );
  XOR U8067 ( .A(p_input[450]), .B(n8396), .Z(n8398) );
  XNOR U8068 ( .A(n8399), .B(n8400), .Z(n8396) );
  AND U8069 ( .A(n401), .B(n8401), .Z(n8400) );
  XOR U8070 ( .A(n8402), .B(n8403), .Z(n8394) );
  AND U8071 ( .A(n405), .B(n8393), .Z(n8403) );
  XNOR U8072 ( .A(n8404), .B(n8391), .Z(n8393) );
  XOR U8073 ( .A(n8405), .B(n8406), .Z(n8391) );
  AND U8074 ( .A(n428), .B(n8407), .Z(n8406) );
  IV U8075 ( .A(n8402), .Z(n8404) );
  XOR U8076 ( .A(n8408), .B(n8409), .Z(n8402) );
  AND U8077 ( .A(n412), .B(n8401), .Z(n8409) );
  XNOR U8078 ( .A(n8399), .B(n8408), .Z(n8401) );
  XNOR U8079 ( .A(n8410), .B(n8411), .Z(n8399) );
  AND U8080 ( .A(n416), .B(n8412), .Z(n8411) );
  XOR U8081 ( .A(p_input[482]), .B(n8410), .Z(n8412) );
  XNOR U8082 ( .A(n8413), .B(n8414), .Z(n8410) );
  AND U8083 ( .A(n420), .B(n8415), .Z(n8414) );
  XOR U8084 ( .A(n8416), .B(n8417), .Z(n8408) );
  AND U8085 ( .A(n424), .B(n8407), .Z(n8417) );
  XNOR U8086 ( .A(n8418), .B(n8405), .Z(n8407) );
  XOR U8087 ( .A(n8419), .B(n8420), .Z(n8405) );
  AND U8088 ( .A(n447), .B(n8421), .Z(n8420) );
  IV U8089 ( .A(n8416), .Z(n8418) );
  XOR U8090 ( .A(n8422), .B(n8423), .Z(n8416) );
  AND U8091 ( .A(n431), .B(n8415), .Z(n8423) );
  XNOR U8092 ( .A(n8413), .B(n8422), .Z(n8415) );
  XNOR U8093 ( .A(n8424), .B(n8425), .Z(n8413) );
  AND U8094 ( .A(n435), .B(n8426), .Z(n8425) );
  XOR U8095 ( .A(p_input[514]), .B(n8424), .Z(n8426) );
  XNOR U8096 ( .A(n8427), .B(n8428), .Z(n8424) );
  AND U8097 ( .A(n439), .B(n8429), .Z(n8428) );
  XOR U8098 ( .A(n8430), .B(n8431), .Z(n8422) );
  AND U8099 ( .A(n443), .B(n8421), .Z(n8431) );
  XNOR U8100 ( .A(n8432), .B(n8419), .Z(n8421) );
  XOR U8101 ( .A(n8433), .B(n8434), .Z(n8419) );
  AND U8102 ( .A(n466), .B(n8435), .Z(n8434) );
  IV U8103 ( .A(n8430), .Z(n8432) );
  XOR U8104 ( .A(n8436), .B(n8437), .Z(n8430) );
  AND U8105 ( .A(n450), .B(n8429), .Z(n8437) );
  XNOR U8106 ( .A(n8427), .B(n8436), .Z(n8429) );
  XNOR U8107 ( .A(n8438), .B(n8439), .Z(n8427) );
  AND U8108 ( .A(n454), .B(n8440), .Z(n8439) );
  XOR U8109 ( .A(p_input[546]), .B(n8438), .Z(n8440) );
  XNOR U8110 ( .A(n8441), .B(n8442), .Z(n8438) );
  AND U8111 ( .A(n458), .B(n8443), .Z(n8442) );
  XOR U8112 ( .A(n8444), .B(n8445), .Z(n8436) );
  AND U8113 ( .A(n462), .B(n8435), .Z(n8445) );
  XNOR U8114 ( .A(n8446), .B(n8433), .Z(n8435) );
  XOR U8115 ( .A(n8447), .B(n8448), .Z(n8433) );
  AND U8116 ( .A(n485), .B(n8449), .Z(n8448) );
  IV U8117 ( .A(n8444), .Z(n8446) );
  XOR U8118 ( .A(n8450), .B(n8451), .Z(n8444) );
  AND U8119 ( .A(n469), .B(n8443), .Z(n8451) );
  XNOR U8120 ( .A(n8441), .B(n8450), .Z(n8443) );
  XNOR U8121 ( .A(n8452), .B(n8453), .Z(n8441) );
  AND U8122 ( .A(n473), .B(n8454), .Z(n8453) );
  XOR U8123 ( .A(p_input[578]), .B(n8452), .Z(n8454) );
  XNOR U8124 ( .A(n8455), .B(n8456), .Z(n8452) );
  AND U8125 ( .A(n477), .B(n8457), .Z(n8456) );
  XOR U8126 ( .A(n8458), .B(n8459), .Z(n8450) );
  AND U8127 ( .A(n481), .B(n8449), .Z(n8459) );
  XNOR U8128 ( .A(n8460), .B(n8447), .Z(n8449) );
  XOR U8129 ( .A(n8461), .B(n8462), .Z(n8447) );
  AND U8130 ( .A(n504), .B(n8463), .Z(n8462) );
  IV U8131 ( .A(n8458), .Z(n8460) );
  XOR U8132 ( .A(n8464), .B(n8465), .Z(n8458) );
  AND U8133 ( .A(n488), .B(n8457), .Z(n8465) );
  XNOR U8134 ( .A(n8455), .B(n8464), .Z(n8457) );
  XNOR U8135 ( .A(n8466), .B(n8467), .Z(n8455) );
  AND U8136 ( .A(n492), .B(n8468), .Z(n8467) );
  XOR U8137 ( .A(p_input[610]), .B(n8466), .Z(n8468) );
  XNOR U8138 ( .A(n8469), .B(n8470), .Z(n8466) );
  AND U8139 ( .A(n496), .B(n8471), .Z(n8470) );
  XOR U8140 ( .A(n8472), .B(n8473), .Z(n8464) );
  AND U8141 ( .A(n500), .B(n8463), .Z(n8473) );
  XNOR U8142 ( .A(n8474), .B(n8461), .Z(n8463) );
  XOR U8143 ( .A(n8475), .B(n8476), .Z(n8461) );
  AND U8144 ( .A(n523), .B(n8477), .Z(n8476) );
  IV U8145 ( .A(n8472), .Z(n8474) );
  XOR U8146 ( .A(n8478), .B(n8479), .Z(n8472) );
  AND U8147 ( .A(n507), .B(n8471), .Z(n8479) );
  XNOR U8148 ( .A(n8469), .B(n8478), .Z(n8471) );
  XNOR U8149 ( .A(n8480), .B(n8481), .Z(n8469) );
  AND U8150 ( .A(n511), .B(n8482), .Z(n8481) );
  XOR U8151 ( .A(p_input[642]), .B(n8480), .Z(n8482) );
  XNOR U8152 ( .A(n8483), .B(n8484), .Z(n8480) );
  AND U8153 ( .A(n515), .B(n8485), .Z(n8484) );
  XOR U8154 ( .A(n8486), .B(n8487), .Z(n8478) );
  AND U8155 ( .A(n519), .B(n8477), .Z(n8487) );
  XNOR U8156 ( .A(n8488), .B(n8475), .Z(n8477) );
  XOR U8157 ( .A(n8489), .B(n8490), .Z(n8475) );
  AND U8158 ( .A(n542), .B(n8491), .Z(n8490) );
  IV U8159 ( .A(n8486), .Z(n8488) );
  XOR U8160 ( .A(n8492), .B(n8493), .Z(n8486) );
  AND U8161 ( .A(n526), .B(n8485), .Z(n8493) );
  XNOR U8162 ( .A(n8483), .B(n8492), .Z(n8485) );
  XNOR U8163 ( .A(n8494), .B(n8495), .Z(n8483) );
  AND U8164 ( .A(n530), .B(n8496), .Z(n8495) );
  XOR U8165 ( .A(p_input[674]), .B(n8494), .Z(n8496) );
  XNOR U8166 ( .A(n8497), .B(n8498), .Z(n8494) );
  AND U8167 ( .A(n534), .B(n8499), .Z(n8498) );
  XOR U8168 ( .A(n8500), .B(n8501), .Z(n8492) );
  AND U8169 ( .A(n538), .B(n8491), .Z(n8501) );
  XNOR U8170 ( .A(n8502), .B(n8489), .Z(n8491) );
  XOR U8171 ( .A(n8503), .B(n8504), .Z(n8489) );
  AND U8172 ( .A(n561), .B(n8505), .Z(n8504) );
  IV U8173 ( .A(n8500), .Z(n8502) );
  XOR U8174 ( .A(n8506), .B(n8507), .Z(n8500) );
  AND U8175 ( .A(n545), .B(n8499), .Z(n8507) );
  XNOR U8176 ( .A(n8497), .B(n8506), .Z(n8499) );
  XNOR U8177 ( .A(n8508), .B(n8509), .Z(n8497) );
  AND U8178 ( .A(n549), .B(n8510), .Z(n8509) );
  XOR U8179 ( .A(p_input[706]), .B(n8508), .Z(n8510) );
  XNOR U8180 ( .A(n8511), .B(n8512), .Z(n8508) );
  AND U8181 ( .A(n553), .B(n8513), .Z(n8512) );
  XOR U8182 ( .A(n8514), .B(n8515), .Z(n8506) );
  AND U8183 ( .A(n557), .B(n8505), .Z(n8515) );
  XNOR U8184 ( .A(n8516), .B(n8503), .Z(n8505) );
  XOR U8185 ( .A(n8517), .B(n8518), .Z(n8503) );
  AND U8186 ( .A(n580), .B(n8519), .Z(n8518) );
  IV U8187 ( .A(n8514), .Z(n8516) );
  XOR U8188 ( .A(n8520), .B(n8521), .Z(n8514) );
  AND U8189 ( .A(n564), .B(n8513), .Z(n8521) );
  XNOR U8190 ( .A(n8511), .B(n8520), .Z(n8513) );
  XNOR U8191 ( .A(n8522), .B(n8523), .Z(n8511) );
  AND U8192 ( .A(n568), .B(n8524), .Z(n8523) );
  XOR U8193 ( .A(p_input[738]), .B(n8522), .Z(n8524) );
  XNOR U8194 ( .A(n8525), .B(n8526), .Z(n8522) );
  AND U8195 ( .A(n572), .B(n8527), .Z(n8526) );
  XOR U8196 ( .A(n8528), .B(n8529), .Z(n8520) );
  AND U8197 ( .A(n576), .B(n8519), .Z(n8529) );
  XNOR U8198 ( .A(n8530), .B(n8517), .Z(n8519) );
  XOR U8199 ( .A(n8531), .B(n8532), .Z(n8517) );
  AND U8200 ( .A(n599), .B(n8533), .Z(n8532) );
  IV U8201 ( .A(n8528), .Z(n8530) );
  XOR U8202 ( .A(n8534), .B(n8535), .Z(n8528) );
  AND U8203 ( .A(n583), .B(n8527), .Z(n8535) );
  XNOR U8204 ( .A(n8525), .B(n8534), .Z(n8527) );
  XNOR U8205 ( .A(n8536), .B(n8537), .Z(n8525) );
  AND U8206 ( .A(n587), .B(n8538), .Z(n8537) );
  XOR U8207 ( .A(p_input[770]), .B(n8536), .Z(n8538) );
  XNOR U8208 ( .A(n8539), .B(n8540), .Z(n8536) );
  AND U8209 ( .A(n591), .B(n8541), .Z(n8540) );
  XOR U8210 ( .A(n8542), .B(n8543), .Z(n8534) );
  AND U8211 ( .A(n595), .B(n8533), .Z(n8543) );
  XNOR U8212 ( .A(n8544), .B(n8531), .Z(n8533) );
  XOR U8213 ( .A(n8545), .B(n8546), .Z(n8531) );
  AND U8214 ( .A(n618), .B(n8547), .Z(n8546) );
  IV U8215 ( .A(n8542), .Z(n8544) );
  XOR U8216 ( .A(n8548), .B(n8549), .Z(n8542) );
  AND U8217 ( .A(n602), .B(n8541), .Z(n8549) );
  XNOR U8218 ( .A(n8539), .B(n8548), .Z(n8541) );
  XNOR U8219 ( .A(n8550), .B(n8551), .Z(n8539) );
  AND U8220 ( .A(n606), .B(n8552), .Z(n8551) );
  XOR U8221 ( .A(p_input[802]), .B(n8550), .Z(n8552) );
  XNOR U8222 ( .A(n8553), .B(n8554), .Z(n8550) );
  AND U8223 ( .A(n610), .B(n8555), .Z(n8554) );
  XOR U8224 ( .A(n8556), .B(n8557), .Z(n8548) );
  AND U8225 ( .A(n614), .B(n8547), .Z(n8557) );
  XNOR U8226 ( .A(n8558), .B(n8545), .Z(n8547) );
  XOR U8227 ( .A(n8559), .B(n8560), .Z(n8545) );
  AND U8228 ( .A(n637), .B(n8561), .Z(n8560) );
  IV U8229 ( .A(n8556), .Z(n8558) );
  XOR U8230 ( .A(n8562), .B(n8563), .Z(n8556) );
  AND U8231 ( .A(n621), .B(n8555), .Z(n8563) );
  XNOR U8232 ( .A(n8553), .B(n8562), .Z(n8555) );
  XNOR U8233 ( .A(n8564), .B(n8565), .Z(n8553) );
  AND U8234 ( .A(n625), .B(n8566), .Z(n8565) );
  XOR U8235 ( .A(p_input[834]), .B(n8564), .Z(n8566) );
  XNOR U8236 ( .A(n8567), .B(n8568), .Z(n8564) );
  AND U8237 ( .A(n629), .B(n8569), .Z(n8568) );
  XOR U8238 ( .A(n8570), .B(n8571), .Z(n8562) );
  AND U8239 ( .A(n633), .B(n8561), .Z(n8571) );
  XNOR U8240 ( .A(n8572), .B(n8559), .Z(n8561) );
  XOR U8241 ( .A(n8573), .B(n8574), .Z(n8559) );
  AND U8242 ( .A(n656), .B(n8575), .Z(n8574) );
  IV U8243 ( .A(n8570), .Z(n8572) );
  XOR U8244 ( .A(n8576), .B(n8577), .Z(n8570) );
  AND U8245 ( .A(n640), .B(n8569), .Z(n8577) );
  XNOR U8246 ( .A(n8567), .B(n8576), .Z(n8569) );
  XNOR U8247 ( .A(n8578), .B(n8579), .Z(n8567) );
  AND U8248 ( .A(n644), .B(n8580), .Z(n8579) );
  XOR U8249 ( .A(p_input[866]), .B(n8578), .Z(n8580) );
  XNOR U8250 ( .A(n8581), .B(n8582), .Z(n8578) );
  AND U8251 ( .A(n648), .B(n8583), .Z(n8582) );
  XOR U8252 ( .A(n8584), .B(n8585), .Z(n8576) );
  AND U8253 ( .A(n652), .B(n8575), .Z(n8585) );
  XNOR U8254 ( .A(n8586), .B(n8573), .Z(n8575) );
  XOR U8255 ( .A(n8587), .B(n8588), .Z(n8573) );
  AND U8256 ( .A(n675), .B(n8589), .Z(n8588) );
  IV U8257 ( .A(n8584), .Z(n8586) );
  XOR U8258 ( .A(n8590), .B(n8591), .Z(n8584) );
  AND U8259 ( .A(n659), .B(n8583), .Z(n8591) );
  XNOR U8260 ( .A(n8581), .B(n8590), .Z(n8583) );
  XNOR U8261 ( .A(n8592), .B(n8593), .Z(n8581) );
  AND U8262 ( .A(n663), .B(n8594), .Z(n8593) );
  XOR U8263 ( .A(p_input[898]), .B(n8592), .Z(n8594) );
  XNOR U8264 ( .A(n8595), .B(n8596), .Z(n8592) );
  AND U8265 ( .A(n667), .B(n8597), .Z(n8596) );
  XOR U8266 ( .A(n8598), .B(n8599), .Z(n8590) );
  AND U8267 ( .A(n671), .B(n8589), .Z(n8599) );
  XNOR U8268 ( .A(n8600), .B(n8587), .Z(n8589) );
  XOR U8269 ( .A(n8601), .B(n8602), .Z(n8587) );
  AND U8270 ( .A(n694), .B(n8603), .Z(n8602) );
  IV U8271 ( .A(n8598), .Z(n8600) );
  XOR U8272 ( .A(n8604), .B(n8605), .Z(n8598) );
  AND U8273 ( .A(n678), .B(n8597), .Z(n8605) );
  XNOR U8274 ( .A(n8595), .B(n8604), .Z(n8597) );
  XNOR U8275 ( .A(n8606), .B(n8607), .Z(n8595) );
  AND U8276 ( .A(n682), .B(n8608), .Z(n8607) );
  XOR U8277 ( .A(p_input[930]), .B(n8606), .Z(n8608) );
  XNOR U8278 ( .A(n8609), .B(n8610), .Z(n8606) );
  AND U8279 ( .A(n686), .B(n8611), .Z(n8610) );
  XOR U8280 ( .A(n8612), .B(n8613), .Z(n8604) );
  AND U8281 ( .A(n690), .B(n8603), .Z(n8613) );
  XNOR U8282 ( .A(n8614), .B(n8601), .Z(n8603) );
  XOR U8283 ( .A(n8615), .B(n8616), .Z(n8601) );
  AND U8284 ( .A(n713), .B(n8617), .Z(n8616) );
  IV U8285 ( .A(n8612), .Z(n8614) );
  XOR U8286 ( .A(n8618), .B(n8619), .Z(n8612) );
  AND U8287 ( .A(n697), .B(n8611), .Z(n8619) );
  XNOR U8288 ( .A(n8609), .B(n8618), .Z(n8611) );
  XNOR U8289 ( .A(n8620), .B(n8621), .Z(n8609) );
  AND U8290 ( .A(n701), .B(n8622), .Z(n8621) );
  XOR U8291 ( .A(p_input[962]), .B(n8620), .Z(n8622) );
  XNOR U8292 ( .A(n8623), .B(n8624), .Z(n8620) );
  AND U8293 ( .A(n705), .B(n8625), .Z(n8624) );
  XOR U8294 ( .A(n8626), .B(n8627), .Z(n8618) );
  AND U8295 ( .A(n709), .B(n8617), .Z(n8627) );
  XNOR U8296 ( .A(n8628), .B(n8615), .Z(n8617) );
  XOR U8297 ( .A(n8629), .B(n8630), .Z(n8615) );
  AND U8298 ( .A(n732), .B(n8631), .Z(n8630) );
  IV U8299 ( .A(n8626), .Z(n8628) );
  XOR U8300 ( .A(n8632), .B(n8633), .Z(n8626) );
  AND U8301 ( .A(n716), .B(n8625), .Z(n8633) );
  XNOR U8302 ( .A(n8623), .B(n8632), .Z(n8625) );
  XNOR U8303 ( .A(n8634), .B(n8635), .Z(n8623) );
  AND U8304 ( .A(n720), .B(n8636), .Z(n8635) );
  XOR U8305 ( .A(p_input[994]), .B(n8634), .Z(n8636) );
  XNOR U8306 ( .A(n8637), .B(n8638), .Z(n8634) );
  AND U8307 ( .A(n724), .B(n8639), .Z(n8638) );
  XOR U8308 ( .A(n8640), .B(n8641), .Z(n8632) );
  AND U8309 ( .A(n728), .B(n8631), .Z(n8641) );
  XNOR U8310 ( .A(n8642), .B(n8629), .Z(n8631) );
  XOR U8311 ( .A(n8643), .B(n8644), .Z(n8629) );
  AND U8312 ( .A(n751), .B(n8645), .Z(n8644) );
  IV U8313 ( .A(n8640), .Z(n8642) );
  XOR U8314 ( .A(n8646), .B(n8647), .Z(n8640) );
  AND U8315 ( .A(n735), .B(n8639), .Z(n8647) );
  XNOR U8316 ( .A(n8637), .B(n8646), .Z(n8639) );
  XNOR U8317 ( .A(n8648), .B(n8649), .Z(n8637) );
  AND U8318 ( .A(n739), .B(n8650), .Z(n8649) );
  XOR U8319 ( .A(p_input[1026]), .B(n8648), .Z(n8650) );
  XNOR U8320 ( .A(n8651), .B(n8652), .Z(n8648) );
  AND U8321 ( .A(n743), .B(n8653), .Z(n8652) );
  XOR U8322 ( .A(n8654), .B(n8655), .Z(n8646) );
  AND U8323 ( .A(n747), .B(n8645), .Z(n8655) );
  XNOR U8324 ( .A(n8656), .B(n8643), .Z(n8645) );
  XOR U8325 ( .A(n8657), .B(n8658), .Z(n8643) );
  AND U8326 ( .A(n770), .B(n8659), .Z(n8658) );
  IV U8327 ( .A(n8654), .Z(n8656) );
  XOR U8328 ( .A(n8660), .B(n8661), .Z(n8654) );
  AND U8329 ( .A(n754), .B(n8653), .Z(n8661) );
  XNOR U8330 ( .A(n8651), .B(n8660), .Z(n8653) );
  XNOR U8331 ( .A(n8662), .B(n8663), .Z(n8651) );
  AND U8332 ( .A(n758), .B(n8664), .Z(n8663) );
  XOR U8333 ( .A(p_input[1058]), .B(n8662), .Z(n8664) );
  XNOR U8334 ( .A(n8665), .B(n8666), .Z(n8662) );
  AND U8335 ( .A(n762), .B(n8667), .Z(n8666) );
  XOR U8336 ( .A(n8668), .B(n8669), .Z(n8660) );
  AND U8337 ( .A(n766), .B(n8659), .Z(n8669) );
  XNOR U8338 ( .A(n8670), .B(n8657), .Z(n8659) );
  XOR U8339 ( .A(n8671), .B(n8672), .Z(n8657) );
  AND U8340 ( .A(n789), .B(n8673), .Z(n8672) );
  IV U8341 ( .A(n8668), .Z(n8670) );
  XOR U8342 ( .A(n8674), .B(n8675), .Z(n8668) );
  AND U8343 ( .A(n773), .B(n8667), .Z(n8675) );
  XNOR U8344 ( .A(n8665), .B(n8674), .Z(n8667) );
  XNOR U8345 ( .A(n8676), .B(n8677), .Z(n8665) );
  AND U8346 ( .A(n777), .B(n8678), .Z(n8677) );
  XOR U8347 ( .A(p_input[1090]), .B(n8676), .Z(n8678) );
  XNOR U8348 ( .A(n8679), .B(n8680), .Z(n8676) );
  AND U8349 ( .A(n781), .B(n8681), .Z(n8680) );
  XOR U8350 ( .A(n8682), .B(n8683), .Z(n8674) );
  AND U8351 ( .A(n785), .B(n8673), .Z(n8683) );
  XNOR U8352 ( .A(n8684), .B(n8671), .Z(n8673) );
  XOR U8353 ( .A(n8685), .B(n8686), .Z(n8671) );
  AND U8354 ( .A(n808), .B(n8687), .Z(n8686) );
  IV U8355 ( .A(n8682), .Z(n8684) );
  XOR U8356 ( .A(n8688), .B(n8689), .Z(n8682) );
  AND U8357 ( .A(n792), .B(n8681), .Z(n8689) );
  XNOR U8358 ( .A(n8679), .B(n8688), .Z(n8681) );
  XNOR U8359 ( .A(n8690), .B(n8691), .Z(n8679) );
  AND U8360 ( .A(n796), .B(n8692), .Z(n8691) );
  XOR U8361 ( .A(p_input[1122]), .B(n8690), .Z(n8692) );
  XNOR U8362 ( .A(n8693), .B(n8694), .Z(n8690) );
  AND U8363 ( .A(n800), .B(n8695), .Z(n8694) );
  XOR U8364 ( .A(n8696), .B(n8697), .Z(n8688) );
  AND U8365 ( .A(n804), .B(n8687), .Z(n8697) );
  XNOR U8366 ( .A(n8698), .B(n8685), .Z(n8687) );
  XOR U8367 ( .A(n8699), .B(n8700), .Z(n8685) );
  AND U8368 ( .A(n827), .B(n8701), .Z(n8700) );
  IV U8369 ( .A(n8696), .Z(n8698) );
  XOR U8370 ( .A(n8702), .B(n8703), .Z(n8696) );
  AND U8371 ( .A(n811), .B(n8695), .Z(n8703) );
  XNOR U8372 ( .A(n8693), .B(n8702), .Z(n8695) );
  XNOR U8373 ( .A(n8704), .B(n8705), .Z(n8693) );
  AND U8374 ( .A(n815), .B(n8706), .Z(n8705) );
  XOR U8375 ( .A(p_input[1154]), .B(n8704), .Z(n8706) );
  XNOR U8376 ( .A(n8707), .B(n8708), .Z(n8704) );
  AND U8377 ( .A(n819), .B(n8709), .Z(n8708) );
  XOR U8378 ( .A(n8710), .B(n8711), .Z(n8702) );
  AND U8379 ( .A(n823), .B(n8701), .Z(n8711) );
  XNOR U8380 ( .A(n8712), .B(n8699), .Z(n8701) );
  XOR U8381 ( .A(n8713), .B(n8714), .Z(n8699) );
  AND U8382 ( .A(n846), .B(n8715), .Z(n8714) );
  IV U8383 ( .A(n8710), .Z(n8712) );
  XOR U8384 ( .A(n8716), .B(n8717), .Z(n8710) );
  AND U8385 ( .A(n830), .B(n8709), .Z(n8717) );
  XNOR U8386 ( .A(n8707), .B(n8716), .Z(n8709) );
  XNOR U8387 ( .A(n8718), .B(n8719), .Z(n8707) );
  AND U8388 ( .A(n834), .B(n8720), .Z(n8719) );
  XOR U8389 ( .A(p_input[1186]), .B(n8718), .Z(n8720) );
  XNOR U8390 ( .A(n8721), .B(n8722), .Z(n8718) );
  AND U8391 ( .A(n838), .B(n8723), .Z(n8722) );
  XOR U8392 ( .A(n8724), .B(n8725), .Z(n8716) );
  AND U8393 ( .A(n842), .B(n8715), .Z(n8725) );
  XNOR U8394 ( .A(n8726), .B(n8713), .Z(n8715) );
  XOR U8395 ( .A(n8727), .B(n8728), .Z(n8713) );
  AND U8396 ( .A(n865), .B(n8729), .Z(n8728) );
  IV U8397 ( .A(n8724), .Z(n8726) );
  XOR U8398 ( .A(n8730), .B(n8731), .Z(n8724) );
  AND U8399 ( .A(n849), .B(n8723), .Z(n8731) );
  XNOR U8400 ( .A(n8721), .B(n8730), .Z(n8723) );
  XNOR U8401 ( .A(n8732), .B(n8733), .Z(n8721) );
  AND U8402 ( .A(n853), .B(n8734), .Z(n8733) );
  XOR U8403 ( .A(p_input[1218]), .B(n8732), .Z(n8734) );
  XNOR U8404 ( .A(n8735), .B(n8736), .Z(n8732) );
  AND U8405 ( .A(n857), .B(n8737), .Z(n8736) );
  XOR U8406 ( .A(n8738), .B(n8739), .Z(n8730) );
  AND U8407 ( .A(n861), .B(n8729), .Z(n8739) );
  XNOR U8408 ( .A(n8740), .B(n8727), .Z(n8729) );
  XOR U8409 ( .A(n8741), .B(n8742), .Z(n8727) );
  AND U8410 ( .A(n884), .B(n8743), .Z(n8742) );
  IV U8411 ( .A(n8738), .Z(n8740) );
  XOR U8412 ( .A(n8744), .B(n8745), .Z(n8738) );
  AND U8413 ( .A(n868), .B(n8737), .Z(n8745) );
  XNOR U8414 ( .A(n8735), .B(n8744), .Z(n8737) );
  XNOR U8415 ( .A(n8746), .B(n8747), .Z(n8735) );
  AND U8416 ( .A(n872), .B(n8748), .Z(n8747) );
  XOR U8417 ( .A(p_input[1250]), .B(n8746), .Z(n8748) );
  XNOR U8418 ( .A(n8749), .B(n8750), .Z(n8746) );
  AND U8419 ( .A(n876), .B(n8751), .Z(n8750) );
  XOR U8420 ( .A(n8752), .B(n8753), .Z(n8744) );
  AND U8421 ( .A(n880), .B(n8743), .Z(n8753) );
  XNOR U8422 ( .A(n8754), .B(n8741), .Z(n8743) );
  XOR U8423 ( .A(n8755), .B(n8756), .Z(n8741) );
  AND U8424 ( .A(n903), .B(n8757), .Z(n8756) );
  IV U8425 ( .A(n8752), .Z(n8754) );
  XOR U8426 ( .A(n8758), .B(n8759), .Z(n8752) );
  AND U8427 ( .A(n887), .B(n8751), .Z(n8759) );
  XNOR U8428 ( .A(n8749), .B(n8758), .Z(n8751) );
  XNOR U8429 ( .A(n8760), .B(n8761), .Z(n8749) );
  AND U8430 ( .A(n891), .B(n8762), .Z(n8761) );
  XOR U8431 ( .A(p_input[1282]), .B(n8760), .Z(n8762) );
  XNOR U8432 ( .A(n8763), .B(n8764), .Z(n8760) );
  AND U8433 ( .A(n895), .B(n8765), .Z(n8764) );
  XOR U8434 ( .A(n8766), .B(n8767), .Z(n8758) );
  AND U8435 ( .A(n899), .B(n8757), .Z(n8767) );
  XNOR U8436 ( .A(n8768), .B(n8755), .Z(n8757) );
  XOR U8437 ( .A(n8769), .B(n8770), .Z(n8755) );
  AND U8438 ( .A(n922), .B(n8771), .Z(n8770) );
  IV U8439 ( .A(n8766), .Z(n8768) );
  XOR U8440 ( .A(n8772), .B(n8773), .Z(n8766) );
  AND U8441 ( .A(n906), .B(n8765), .Z(n8773) );
  XNOR U8442 ( .A(n8763), .B(n8772), .Z(n8765) );
  XNOR U8443 ( .A(n8774), .B(n8775), .Z(n8763) );
  AND U8444 ( .A(n910), .B(n8776), .Z(n8775) );
  XOR U8445 ( .A(p_input[1314]), .B(n8774), .Z(n8776) );
  XNOR U8446 ( .A(n8777), .B(n8778), .Z(n8774) );
  AND U8447 ( .A(n914), .B(n8779), .Z(n8778) );
  XOR U8448 ( .A(n8780), .B(n8781), .Z(n8772) );
  AND U8449 ( .A(n918), .B(n8771), .Z(n8781) );
  XNOR U8450 ( .A(n8782), .B(n8769), .Z(n8771) );
  XOR U8451 ( .A(n8783), .B(n8784), .Z(n8769) );
  AND U8452 ( .A(n941), .B(n8785), .Z(n8784) );
  IV U8453 ( .A(n8780), .Z(n8782) );
  XOR U8454 ( .A(n8786), .B(n8787), .Z(n8780) );
  AND U8455 ( .A(n925), .B(n8779), .Z(n8787) );
  XNOR U8456 ( .A(n8777), .B(n8786), .Z(n8779) );
  XNOR U8457 ( .A(n8788), .B(n8789), .Z(n8777) );
  AND U8458 ( .A(n929), .B(n8790), .Z(n8789) );
  XOR U8459 ( .A(p_input[1346]), .B(n8788), .Z(n8790) );
  XNOR U8460 ( .A(n8791), .B(n8792), .Z(n8788) );
  AND U8461 ( .A(n933), .B(n8793), .Z(n8792) );
  XOR U8462 ( .A(n8794), .B(n8795), .Z(n8786) );
  AND U8463 ( .A(n937), .B(n8785), .Z(n8795) );
  XNOR U8464 ( .A(n8796), .B(n8783), .Z(n8785) );
  XOR U8465 ( .A(n8797), .B(n8798), .Z(n8783) );
  AND U8466 ( .A(n960), .B(n8799), .Z(n8798) );
  IV U8467 ( .A(n8794), .Z(n8796) );
  XOR U8468 ( .A(n8800), .B(n8801), .Z(n8794) );
  AND U8469 ( .A(n944), .B(n8793), .Z(n8801) );
  XNOR U8470 ( .A(n8791), .B(n8800), .Z(n8793) );
  XNOR U8471 ( .A(n8802), .B(n8803), .Z(n8791) );
  AND U8472 ( .A(n948), .B(n8804), .Z(n8803) );
  XOR U8473 ( .A(p_input[1378]), .B(n8802), .Z(n8804) );
  XNOR U8474 ( .A(n8805), .B(n8806), .Z(n8802) );
  AND U8475 ( .A(n952), .B(n8807), .Z(n8806) );
  XOR U8476 ( .A(n8808), .B(n8809), .Z(n8800) );
  AND U8477 ( .A(n956), .B(n8799), .Z(n8809) );
  XNOR U8478 ( .A(n8810), .B(n8797), .Z(n8799) );
  XOR U8479 ( .A(n8811), .B(n8812), .Z(n8797) );
  AND U8480 ( .A(n979), .B(n8813), .Z(n8812) );
  IV U8481 ( .A(n8808), .Z(n8810) );
  XOR U8482 ( .A(n8814), .B(n8815), .Z(n8808) );
  AND U8483 ( .A(n963), .B(n8807), .Z(n8815) );
  XNOR U8484 ( .A(n8805), .B(n8814), .Z(n8807) );
  XNOR U8485 ( .A(n8816), .B(n8817), .Z(n8805) );
  AND U8486 ( .A(n967), .B(n8818), .Z(n8817) );
  XOR U8487 ( .A(p_input[1410]), .B(n8816), .Z(n8818) );
  XNOR U8488 ( .A(n8819), .B(n8820), .Z(n8816) );
  AND U8489 ( .A(n971), .B(n8821), .Z(n8820) );
  XOR U8490 ( .A(n8822), .B(n8823), .Z(n8814) );
  AND U8491 ( .A(n975), .B(n8813), .Z(n8823) );
  XNOR U8492 ( .A(n8824), .B(n8811), .Z(n8813) );
  XOR U8493 ( .A(n8825), .B(n8826), .Z(n8811) );
  AND U8494 ( .A(n998), .B(n8827), .Z(n8826) );
  IV U8495 ( .A(n8822), .Z(n8824) );
  XOR U8496 ( .A(n8828), .B(n8829), .Z(n8822) );
  AND U8497 ( .A(n982), .B(n8821), .Z(n8829) );
  XNOR U8498 ( .A(n8819), .B(n8828), .Z(n8821) );
  XNOR U8499 ( .A(n8830), .B(n8831), .Z(n8819) );
  AND U8500 ( .A(n986), .B(n8832), .Z(n8831) );
  XOR U8501 ( .A(p_input[1442]), .B(n8830), .Z(n8832) );
  XNOR U8502 ( .A(n8833), .B(n8834), .Z(n8830) );
  AND U8503 ( .A(n990), .B(n8835), .Z(n8834) );
  XOR U8504 ( .A(n8836), .B(n8837), .Z(n8828) );
  AND U8505 ( .A(n994), .B(n8827), .Z(n8837) );
  XNOR U8506 ( .A(n8838), .B(n8825), .Z(n8827) );
  XOR U8507 ( .A(n8839), .B(n8840), .Z(n8825) );
  AND U8508 ( .A(n1017), .B(n8841), .Z(n8840) );
  IV U8509 ( .A(n8836), .Z(n8838) );
  XOR U8510 ( .A(n8842), .B(n8843), .Z(n8836) );
  AND U8511 ( .A(n1001), .B(n8835), .Z(n8843) );
  XNOR U8512 ( .A(n8833), .B(n8842), .Z(n8835) );
  XNOR U8513 ( .A(n8844), .B(n8845), .Z(n8833) );
  AND U8514 ( .A(n1005), .B(n8846), .Z(n8845) );
  XOR U8515 ( .A(p_input[1474]), .B(n8844), .Z(n8846) );
  XNOR U8516 ( .A(n8847), .B(n8848), .Z(n8844) );
  AND U8517 ( .A(n1009), .B(n8849), .Z(n8848) );
  XOR U8518 ( .A(n8850), .B(n8851), .Z(n8842) );
  AND U8519 ( .A(n1013), .B(n8841), .Z(n8851) );
  XNOR U8520 ( .A(n8852), .B(n8839), .Z(n8841) );
  XOR U8521 ( .A(n8853), .B(n8854), .Z(n8839) );
  AND U8522 ( .A(n1036), .B(n8855), .Z(n8854) );
  IV U8523 ( .A(n8850), .Z(n8852) );
  XOR U8524 ( .A(n8856), .B(n8857), .Z(n8850) );
  AND U8525 ( .A(n1020), .B(n8849), .Z(n8857) );
  XNOR U8526 ( .A(n8847), .B(n8856), .Z(n8849) );
  XNOR U8527 ( .A(n8858), .B(n8859), .Z(n8847) );
  AND U8528 ( .A(n1024), .B(n8860), .Z(n8859) );
  XOR U8529 ( .A(p_input[1506]), .B(n8858), .Z(n8860) );
  XNOR U8530 ( .A(n8861), .B(n8862), .Z(n8858) );
  AND U8531 ( .A(n1028), .B(n8863), .Z(n8862) );
  XOR U8532 ( .A(n8864), .B(n8865), .Z(n8856) );
  AND U8533 ( .A(n1032), .B(n8855), .Z(n8865) );
  XNOR U8534 ( .A(n8866), .B(n8853), .Z(n8855) );
  XOR U8535 ( .A(n8867), .B(n8868), .Z(n8853) );
  AND U8536 ( .A(n1055), .B(n8869), .Z(n8868) );
  IV U8537 ( .A(n8864), .Z(n8866) );
  XOR U8538 ( .A(n8870), .B(n8871), .Z(n8864) );
  AND U8539 ( .A(n1039), .B(n8863), .Z(n8871) );
  XNOR U8540 ( .A(n8861), .B(n8870), .Z(n8863) );
  XNOR U8541 ( .A(n8872), .B(n8873), .Z(n8861) );
  AND U8542 ( .A(n1043), .B(n8874), .Z(n8873) );
  XOR U8543 ( .A(p_input[1538]), .B(n8872), .Z(n8874) );
  XNOR U8544 ( .A(n8875), .B(n8876), .Z(n8872) );
  AND U8545 ( .A(n1047), .B(n8877), .Z(n8876) );
  XOR U8546 ( .A(n8878), .B(n8879), .Z(n8870) );
  AND U8547 ( .A(n1051), .B(n8869), .Z(n8879) );
  XNOR U8548 ( .A(n8880), .B(n8867), .Z(n8869) );
  XOR U8549 ( .A(n8881), .B(n8882), .Z(n8867) );
  AND U8550 ( .A(n1074), .B(n8883), .Z(n8882) );
  IV U8551 ( .A(n8878), .Z(n8880) );
  XOR U8552 ( .A(n8884), .B(n8885), .Z(n8878) );
  AND U8553 ( .A(n1058), .B(n8877), .Z(n8885) );
  XNOR U8554 ( .A(n8875), .B(n8884), .Z(n8877) );
  XNOR U8555 ( .A(n8886), .B(n8887), .Z(n8875) );
  AND U8556 ( .A(n1062), .B(n8888), .Z(n8887) );
  XOR U8557 ( .A(p_input[1570]), .B(n8886), .Z(n8888) );
  XNOR U8558 ( .A(n8889), .B(n8890), .Z(n8886) );
  AND U8559 ( .A(n1066), .B(n8891), .Z(n8890) );
  XOR U8560 ( .A(n8892), .B(n8893), .Z(n8884) );
  AND U8561 ( .A(n1070), .B(n8883), .Z(n8893) );
  XNOR U8562 ( .A(n8894), .B(n8881), .Z(n8883) );
  XOR U8563 ( .A(n8895), .B(n8896), .Z(n8881) );
  AND U8564 ( .A(n1093), .B(n8897), .Z(n8896) );
  IV U8565 ( .A(n8892), .Z(n8894) );
  XOR U8566 ( .A(n8898), .B(n8899), .Z(n8892) );
  AND U8567 ( .A(n1077), .B(n8891), .Z(n8899) );
  XNOR U8568 ( .A(n8889), .B(n8898), .Z(n8891) );
  XNOR U8569 ( .A(n8900), .B(n8901), .Z(n8889) );
  AND U8570 ( .A(n1081), .B(n8902), .Z(n8901) );
  XOR U8571 ( .A(p_input[1602]), .B(n8900), .Z(n8902) );
  XNOR U8572 ( .A(n8903), .B(n8904), .Z(n8900) );
  AND U8573 ( .A(n1085), .B(n8905), .Z(n8904) );
  XOR U8574 ( .A(n8906), .B(n8907), .Z(n8898) );
  AND U8575 ( .A(n1089), .B(n8897), .Z(n8907) );
  XNOR U8576 ( .A(n8908), .B(n8895), .Z(n8897) );
  XOR U8577 ( .A(n8909), .B(n8910), .Z(n8895) );
  AND U8578 ( .A(n1112), .B(n8911), .Z(n8910) );
  IV U8579 ( .A(n8906), .Z(n8908) );
  XOR U8580 ( .A(n8912), .B(n8913), .Z(n8906) );
  AND U8581 ( .A(n1096), .B(n8905), .Z(n8913) );
  XNOR U8582 ( .A(n8903), .B(n8912), .Z(n8905) );
  XNOR U8583 ( .A(n8914), .B(n8915), .Z(n8903) );
  AND U8584 ( .A(n1100), .B(n8916), .Z(n8915) );
  XOR U8585 ( .A(p_input[1634]), .B(n8914), .Z(n8916) );
  XNOR U8586 ( .A(n8917), .B(n8918), .Z(n8914) );
  AND U8587 ( .A(n1104), .B(n8919), .Z(n8918) );
  XOR U8588 ( .A(n8920), .B(n8921), .Z(n8912) );
  AND U8589 ( .A(n1108), .B(n8911), .Z(n8921) );
  XNOR U8590 ( .A(n8922), .B(n8909), .Z(n8911) );
  XOR U8591 ( .A(n8923), .B(n8924), .Z(n8909) );
  AND U8592 ( .A(n1131), .B(n8925), .Z(n8924) );
  IV U8593 ( .A(n8920), .Z(n8922) );
  XOR U8594 ( .A(n8926), .B(n8927), .Z(n8920) );
  AND U8595 ( .A(n1115), .B(n8919), .Z(n8927) );
  XNOR U8596 ( .A(n8917), .B(n8926), .Z(n8919) );
  XNOR U8597 ( .A(n8928), .B(n8929), .Z(n8917) );
  AND U8598 ( .A(n1119), .B(n8930), .Z(n8929) );
  XOR U8599 ( .A(p_input[1666]), .B(n8928), .Z(n8930) );
  XNOR U8600 ( .A(n8931), .B(n8932), .Z(n8928) );
  AND U8601 ( .A(n1123), .B(n8933), .Z(n8932) );
  XOR U8602 ( .A(n8934), .B(n8935), .Z(n8926) );
  AND U8603 ( .A(n1127), .B(n8925), .Z(n8935) );
  XNOR U8604 ( .A(n8936), .B(n8923), .Z(n8925) );
  XOR U8605 ( .A(n8937), .B(n8938), .Z(n8923) );
  AND U8606 ( .A(n1150), .B(n8939), .Z(n8938) );
  IV U8607 ( .A(n8934), .Z(n8936) );
  XOR U8608 ( .A(n8940), .B(n8941), .Z(n8934) );
  AND U8609 ( .A(n1134), .B(n8933), .Z(n8941) );
  XNOR U8610 ( .A(n8931), .B(n8940), .Z(n8933) );
  XNOR U8611 ( .A(n8942), .B(n8943), .Z(n8931) );
  AND U8612 ( .A(n1138), .B(n8944), .Z(n8943) );
  XOR U8613 ( .A(p_input[1698]), .B(n8942), .Z(n8944) );
  XNOR U8614 ( .A(n8945), .B(n8946), .Z(n8942) );
  AND U8615 ( .A(n1142), .B(n8947), .Z(n8946) );
  XOR U8616 ( .A(n8948), .B(n8949), .Z(n8940) );
  AND U8617 ( .A(n1146), .B(n8939), .Z(n8949) );
  XNOR U8618 ( .A(n8950), .B(n8937), .Z(n8939) );
  XOR U8619 ( .A(n8951), .B(n8952), .Z(n8937) );
  AND U8620 ( .A(n1169), .B(n8953), .Z(n8952) );
  IV U8621 ( .A(n8948), .Z(n8950) );
  XOR U8622 ( .A(n8954), .B(n8955), .Z(n8948) );
  AND U8623 ( .A(n1153), .B(n8947), .Z(n8955) );
  XNOR U8624 ( .A(n8945), .B(n8954), .Z(n8947) );
  XNOR U8625 ( .A(n8956), .B(n8957), .Z(n8945) );
  AND U8626 ( .A(n1157), .B(n8958), .Z(n8957) );
  XOR U8627 ( .A(p_input[1730]), .B(n8956), .Z(n8958) );
  XNOR U8628 ( .A(n8959), .B(n8960), .Z(n8956) );
  AND U8629 ( .A(n1161), .B(n8961), .Z(n8960) );
  XOR U8630 ( .A(n8962), .B(n8963), .Z(n8954) );
  AND U8631 ( .A(n1165), .B(n8953), .Z(n8963) );
  XNOR U8632 ( .A(n8964), .B(n8951), .Z(n8953) );
  XOR U8633 ( .A(n8965), .B(n8966), .Z(n8951) );
  AND U8634 ( .A(n1188), .B(n8967), .Z(n8966) );
  IV U8635 ( .A(n8962), .Z(n8964) );
  XOR U8636 ( .A(n8968), .B(n8969), .Z(n8962) );
  AND U8637 ( .A(n1172), .B(n8961), .Z(n8969) );
  XNOR U8638 ( .A(n8959), .B(n8968), .Z(n8961) );
  XNOR U8639 ( .A(n8970), .B(n8971), .Z(n8959) );
  AND U8640 ( .A(n1176), .B(n8972), .Z(n8971) );
  XOR U8641 ( .A(p_input[1762]), .B(n8970), .Z(n8972) );
  XNOR U8642 ( .A(n8973), .B(n8974), .Z(n8970) );
  AND U8643 ( .A(n1180), .B(n8975), .Z(n8974) );
  XOR U8644 ( .A(n8976), .B(n8977), .Z(n8968) );
  AND U8645 ( .A(n1184), .B(n8967), .Z(n8977) );
  XNOR U8646 ( .A(n8978), .B(n8965), .Z(n8967) );
  XOR U8647 ( .A(n8979), .B(n8980), .Z(n8965) );
  AND U8648 ( .A(n1207), .B(n8981), .Z(n8980) );
  IV U8649 ( .A(n8976), .Z(n8978) );
  XOR U8650 ( .A(n8982), .B(n8983), .Z(n8976) );
  AND U8651 ( .A(n1191), .B(n8975), .Z(n8983) );
  XNOR U8652 ( .A(n8973), .B(n8982), .Z(n8975) );
  XNOR U8653 ( .A(n8984), .B(n8985), .Z(n8973) );
  AND U8654 ( .A(n1195), .B(n8986), .Z(n8985) );
  XOR U8655 ( .A(p_input[1794]), .B(n8984), .Z(n8986) );
  XNOR U8656 ( .A(n8987), .B(n8988), .Z(n8984) );
  AND U8657 ( .A(n1199), .B(n8989), .Z(n8988) );
  XOR U8658 ( .A(n8990), .B(n8991), .Z(n8982) );
  AND U8659 ( .A(n1203), .B(n8981), .Z(n8991) );
  XNOR U8660 ( .A(n8992), .B(n8979), .Z(n8981) );
  XOR U8661 ( .A(n8993), .B(n8994), .Z(n8979) );
  AND U8662 ( .A(n1226), .B(n8995), .Z(n8994) );
  IV U8663 ( .A(n8990), .Z(n8992) );
  XOR U8664 ( .A(n8996), .B(n8997), .Z(n8990) );
  AND U8665 ( .A(n1210), .B(n8989), .Z(n8997) );
  XNOR U8666 ( .A(n8987), .B(n8996), .Z(n8989) );
  XNOR U8667 ( .A(n8998), .B(n8999), .Z(n8987) );
  AND U8668 ( .A(n1214), .B(n9000), .Z(n8999) );
  XOR U8669 ( .A(p_input[1826]), .B(n8998), .Z(n9000) );
  XNOR U8670 ( .A(n9001), .B(n9002), .Z(n8998) );
  AND U8671 ( .A(n1218), .B(n9003), .Z(n9002) );
  XOR U8672 ( .A(n9004), .B(n9005), .Z(n8996) );
  AND U8673 ( .A(n1222), .B(n8995), .Z(n9005) );
  XNOR U8674 ( .A(n9006), .B(n8993), .Z(n8995) );
  XOR U8675 ( .A(n9007), .B(n9008), .Z(n8993) );
  AND U8676 ( .A(n1245), .B(n9009), .Z(n9008) );
  IV U8677 ( .A(n9004), .Z(n9006) );
  XOR U8678 ( .A(n9010), .B(n9011), .Z(n9004) );
  AND U8679 ( .A(n1229), .B(n9003), .Z(n9011) );
  XNOR U8680 ( .A(n9001), .B(n9010), .Z(n9003) );
  XNOR U8681 ( .A(n9012), .B(n9013), .Z(n9001) );
  AND U8682 ( .A(n1233), .B(n9014), .Z(n9013) );
  XOR U8683 ( .A(p_input[1858]), .B(n9012), .Z(n9014) );
  XNOR U8684 ( .A(n9015), .B(n9016), .Z(n9012) );
  AND U8685 ( .A(n1237), .B(n9017), .Z(n9016) );
  XOR U8686 ( .A(n9018), .B(n9019), .Z(n9010) );
  AND U8687 ( .A(n1241), .B(n9009), .Z(n9019) );
  XNOR U8688 ( .A(n9020), .B(n9007), .Z(n9009) );
  XOR U8689 ( .A(n9021), .B(n9022), .Z(n9007) );
  AND U8690 ( .A(n1264), .B(n9023), .Z(n9022) );
  IV U8691 ( .A(n9018), .Z(n9020) );
  XOR U8692 ( .A(n9024), .B(n9025), .Z(n9018) );
  AND U8693 ( .A(n1248), .B(n9017), .Z(n9025) );
  XNOR U8694 ( .A(n9015), .B(n9024), .Z(n9017) );
  XNOR U8695 ( .A(n9026), .B(n9027), .Z(n9015) );
  AND U8696 ( .A(n1252), .B(n9028), .Z(n9027) );
  XOR U8697 ( .A(p_input[1890]), .B(n9026), .Z(n9028) );
  XNOR U8698 ( .A(n9029), .B(n9030), .Z(n9026) );
  AND U8699 ( .A(n1256), .B(n9031), .Z(n9030) );
  XOR U8700 ( .A(n9032), .B(n9033), .Z(n9024) );
  AND U8701 ( .A(n1260), .B(n9023), .Z(n9033) );
  XNOR U8702 ( .A(n9034), .B(n9021), .Z(n9023) );
  XOR U8703 ( .A(n9035), .B(n9036), .Z(n9021) );
  AND U8704 ( .A(n1282), .B(n9037), .Z(n9036) );
  IV U8705 ( .A(n9032), .Z(n9034) );
  XOR U8706 ( .A(n9038), .B(n9039), .Z(n9032) );
  AND U8707 ( .A(n1267), .B(n9031), .Z(n9039) );
  XNOR U8708 ( .A(n9029), .B(n9038), .Z(n9031) );
  XNOR U8709 ( .A(n9040), .B(n9041), .Z(n9029) );
  AND U8710 ( .A(n1271), .B(n9042), .Z(n9041) );
  XOR U8711 ( .A(p_input[1922]), .B(n9040), .Z(n9042) );
  XOR U8712 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n9043), 
        .Z(n9040) );
  AND U8713 ( .A(n1274), .B(n9044), .Z(n9043) );
  XOR U8714 ( .A(n9045), .B(n9046), .Z(n9038) );
  AND U8715 ( .A(n1278), .B(n9037), .Z(n9046) );
  XNOR U8716 ( .A(n9047), .B(n9035), .Z(n9037) );
  XOR U8717 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n9048), .Z(n9035) );
  AND U8718 ( .A(n1290), .B(n9049), .Z(n9048) );
  IV U8719 ( .A(n9045), .Z(n9047) );
  XOR U8720 ( .A(n9050), .B(n9051), .Z(n9045) );
  AND U8721 ( .A(n1285), .B(n9044), .Z(n9051) );
  XOR U8722 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n9050), 
        .Z(n9044) );
  XOR U8723 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .B(n9052), 
        .Z(n9050) );
  AND U8724 ( .A(n1287), .B(n9049), .Z(n9052) );
  XOR U8725 ( .A(\knn_comb_/min_val_out[0][2] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n9049) );
  XOR U8726 ( .A(n77), .B(n9053), .Z(o[29]) );
  AND U8727 ( .A(n122), .B(n9054), .Z(n77) );
  XOR U8728 ( .A(n78), .B(n9053), .Z(n9054) );
  XOR U8729 ( .A(n9055), .B(n9056), .Z(n9053) );
  AND U8730 ( .A(n142), .B(n9057), .Z(n9056) );
  XOR U8731 ( .A(n9058), .B(n7), .Z(n78) );
  AND U8732 ( .A(n125), .B(n9059), .Z(n7) );
  XOR U8733 ( .A(n8), .B(n9058), .Z(n9059) );
  XOR U8734 ( .A(n9060), .B(n9061), .Z(n8) );
  AND U8735 ( .A(n130), .B(n9062), .Z(n9061) );
  XOR U8736 ( .A(p_input[29]), .B(n9060), .Z(n9062) );
  XNOR U8737 ( .A(n9063), .B(n9064), .Z(n9060) );
  AND U8738 ( .A(n134), .B(n9065), .Z(n9064) );
  XOR U8739 ( .A(n9066), .B(n9067), .Z(n9058) );
  AND U8740 ( .A(n138), .B(n9057), .Z(n9067) );
  XNOR U8741 ( .A(n9068), .B(n9055), .Z(n9057) );
  XOR U8742 ( .A(n9069), .B(n9070), .Z(n9055) );
  AND U8743 ( .A(n162), .B(n9071), .Z(n9070) );
  IV U8744 ( .A(n9066), .Z(n9068) );
  XOR U8745 ( .A(n9072), .B(n9073), .Z(n9066) );
  AND U8746 ( .A(n146), .B(n9065), .Z(n9073) );
  XNOR U8747 ( .A(n9063), .B(n9072), .Z(n9065) );
  XNOR U8748 ( .A(n9074), .B(n9075), .Z(n9063) );
  AND U8749 ( .A(n150), .B(n9076), .Z(n9075) );
  XOR U8750 ( .A(p_input[61]), .B(n9074), .Z(n9076) );
  XNOR U8751 ( .A(n9077), .B(n9078), .Z(n9074) );
  AND U8752 ( .A(n154), .B(n9079), .Z(n9078) );
  XOR U8753 ( .A(n9080), .B(n9081), .Z(n9072) );
  AND U8754 ( .A(n158), .B(n9071), .Z(n9081) );
  XNOR U8755 ( .A(n9082), .B(n9069), .Z(n9071) );
  XOR U8756 ( .A(n9083), .B(n9084), .Z(n9069) );
  AND U8757 ( .A(n181), .B(n9085), .Z(n9084) );
  IV U8758 ( .A(n9080), .Z(n9082) );
  XOR U8759 ( .A(n9086), .B(n9087), .Z(n9080) );
  AND U8760 ( .A(n165), .B(n9079), .Z(n9087) );
  XNOR U8761 ( .A(n9077), .B(n9086), .Z(n9079) );
  XNOR U8762 ( .A(n9088), .B(n9089), .Z(n9077) );
  AND U8763 ( .A(n169), .B(n9090), .Z(n9089) );
  XOR U8764 ( .A(p_input[93]), .B(n9088), .Z(n9090) );
  XNOR U8765 ( .A(n9091), .B(n9092), .Z(n9088) );
  AND U8766 ( .A(n173), .B(n9093), .Z(n9092) );
  XOR U8767 ( .A(n9094), .B(n9095), .Z(n9086) );
  AND U8768 ( .A(n177), .B(n9085), .Z(n9095) );
  XNOR U8769 ( .A(n9096), .B(n9083), .Z(n9085) );
  XOR U8770 ( .A(n9097), .B(n9098), .Z(n9083) );
  AND U8771 ( .A(n200), .B(n9099), .Z(n9098) );
  IV U8772 ( .A(n9094), .Z(n9096) );
  XOR U8773 ( .A(n9100), .B(n9101), .Z(n9094) );
  AND U8774 ( .A(n184), .B(n9093), .Z(n9101) );
  XNOR U8775 ( .A(n9091), .B(n9100), .Z(n9093) );
  XNOR U8776 ( .A(n9102), .B(n9103), .Z(n9091) );
  AND U8777 ( .A(n188), .B(n9104), .Z(n9103) );
  XOR U8778 ( .A(p_input[125]), .B(n9102), .Z(n9104) );
  XNOR U8779 ( .A(n9105), .B(n9106), .Z(n9102) );
  AND U8780 ( .A(n192), .B(n9107), .Z(n9106) );
  XOR U8781 ( .A(n9108), .B(n9109), .Z(n9100) );
  AND U8782 ( .A(n196), .B(n9099), .Z(n9109) );
  XNOR U8783 ( .A(n9110), .B(n9097), .Z(n9099) );
  XOR U8784 ( .A(n9111), .B(n9112), .Z(n9097) );
  AND U8785 ( .A(n219), .B(n9113), .Z(n9112) );
  IV U8786 ( .A(n9108), .Z(n9110) );
  XOR U8787 ( .A(n9114), .B(n9115), .Z(n9108) );
  AND U8788 ( .A(n203), .B(n9107), .Z(n9115) );
  XNOR U8789 ( .A(n9105), .B(n9114), .Z(n9107) );
  XNOR U8790 ( .A(n9116), .B(n9117), .Z(n9105) );
  AND U8791 ( .A(n207), .B(n9118), .Z(n9117) );
  XOR U8792 ( .A(p_input[157]), .B(n9116), .Z(n9118) );
  XNOR U8793 ( .A(n9119), .B(n9120), .Z(n9116) );
  AND U8794 ( .A(n211), .B(n9121), .Z(n9120) );
  XOR U8795 ( .A(n9122), .B(n9123), .Z(n9114) );
  AND U8796 ( .A(n215), .B(n9113), .Z(n9123) );
  XNOR U8797 ( .A(n9124), .B(n9111), .Z(n9113) );
  XOR U8798 ( .A(n9125), .B(n9126), .Z(n9111) );
  AND U8799 ( .A(n238), .B(n9127), .Z(n9126) );
  IV U8800 ( .A(n9122), .Z(n9124) );
  XOR U8801 ( .A(n9128), .B(n9129), .Z(n9122) );
  AND U8802 ( .A(n222), .B(n9121), .Z(n9129) );
  XNOR U8803 ( .A(n9119), .B(n9128), .Z(n9121) );
  XNOR U8804 ( .A(n9130), .B(n9131), .Z(n9119) );
  AND U8805 ( .A(n226), .B(n9132), .Z(n9131) );
  XOR U8806 ( .A(p_input[189]), .B(n9130), .Z(n9132) );
  XNOR U8807 ( .A(n9133), .B(n9134), .Z(n9130) );
  AND U8808 ( .A(n230), .B(n9135), .Z(n9134) );
  XOR U8809 ( .A(n9136), .B(n9137), .Z(n9128) );
  AND U8810 ( .A(n234), .B(n9127), .Z(n9137) );
  XNOR U8811 ( .A(n9138), .B(n9125), .Z(n9127) );
  XOR U8812 ( .A(n9139), .B(n9140), .Z(n9125) );
  AND U8813 ( .A(n257), .B(n9141), .Z(n9140) );
  IV U8814 ( .A(n9136), .Z(n9138) );
  XOR U8815 ( .A(n9142), .B(n9143), .Z(n9136) );
  AND U8816 ( .A(n241), .B(n9135), .Z(n9143) );
  XNOR U8817 ( .A(n9133), .B(n9142), .Z(n9135) );
  XNOR U8818 ( .A(n9144), .B(n9145), .Z(n9133) );
  AND U8819 ( .A(n245), .B(n9146), .Z(n9145) );
  XOR U8820 ( .A(p_input[221]), .B(n9144), .Z(n9146) );
  XNOR U8821 ( .A(n9147), .B(n9148), .Z(n9144) );
  AND U8822 ( .A(n249), .B(n9149), .Z(n9148) );
  XOR U8823 ( .A(n9150), .B(n9151), .Z(n9142) );
  AND U8824 ( .A(n253), .B(n9141), .Z(n9151) );
  XNOR U8825 ( .A(n9152), .B(n9139), .Z(n9141) );
  XOR U8826 ( .A(n9153), .B(n9154), .Z(n9139) );
  AND U8827 ( .A(n276), .B(n9155), .Z(n9154) );
  IV U8828 ( .A(n9150), .Z(n9152) );
  XOR U8829 ( .A(n9156), .B(n9157), .Z(n9150) );
  AND U8830 ( .A(n260), .B(n9149), .Z(n9157) );
  XNOR U8831 ( .A(n9147), .B(n9156), .Z(n9149) );
  XNOR U8832 ( .A(n9158), .B(n9159), .Z(n9147) );
  AND U8833 ( .A(n264), .B(n9160), .Z(n9159) );
  XOR U8834 ( .A(p_input[253]), .B(n9158), .Z(n9160) );
  XNOR U8835 ( .A(n9161), .B(n9162), .Z(n9158) );
  AND U8836 ( .A(n268), .B(n9163), .Z(n9162) );
  XOR U8837 ( .A(n9164), .B(n9165), .Z(n9156) );
  AND U8838 ( .A(n272), .B(n9155), .Z(n9165) );
  XNOR U8839 ( .A(n9166), .B(n9153), .Z(n9155) );
  XOR U8840 ( .A(n9167), .B(n9168), .Z(n9153) );
  AND U8841 ( .A(n295), .B(n9169), .Z(n9168) );
  IV U8842 ( .A(n9164), .Z(n9166) );
  XOR U8843 ( .A(n9170), .B(n9171), .Z(n9164) );
  AND U8844 ( .A(n279), .B(n9163), .Z(n9171) );
  XNOR U8845 ( .A(n9161), .B(n9170), .Z(n9163) );
  XNOR U8846 ( .A(n9172), .B(n9173), .Z(n9161) );
  AND U8847 ( .A(n283), .B(n9174), .Z(n9173) );
  XOR U8848 ( .A(p_input[285]), .B(n9172), .Z(n9174) );
  XNOR U8849 ( .A(n9175), .B(n9176), .Z(n9172) );
  AND U8850 ( .A(n287), .B(n9177), .Z(n9176) );
  XOR U8851 ( .A(n9178), .B(n9179), .Z(n9170) );
  AND U8852 ( .A(n291), .B(n9169), .Z(n9179) );
  XNOR U8853 ( .A(n9180), .B(n9167), .Z(n9169) );
  XOR U8854 ( .A(n9181), .B(n9182), .Z(n9167) );
  AND U8855 ( .A(n314), .B(n9183), .Z(n9182) );
  IV U8856 ( .A(n9178), .Z(n9180) );
  XOR U8857 ( .A(n9184), .B(n9185), .Z(n9178) );
  AND U8858 ( .A(n298), .B(n9177), .Z(n9185) );
  XNOR U8859 ( .A(n9175), .B(n9184), .Z(n9177) );
  XNOR U8860 ( .A(n9186), .B(n9187), .Z(n9175) );
  AND U8861 ( .A(n302), .B(n9188), .Z(n9187) );
  XOR U8862 ( .A(p_input[317]), .B(n9186), .Z(n9188) );
  XNOR U8863 ( .A(n9189), .B(n9190), .Z(n9186) );
  AND U8864 ( .A(n306), .B(n9191), .Z(n9190) );
  XOR U8865 ( .A(n9192), .B(n9193), .Z(n9184) );
  AND U8866 ( .A(n310), .B(n9183), .Z(n9193) );
  XNOR U8867 ( .A(n9194), .B(n9181), .Z(n9183) );
  XOR U8868 ( .A(n9195), .B(n9196), .Z(n9181) );
  AND U8869 ( .A(n333), .B(n9197), .Z(n9196) );
  IV U8870 ( .A(n9192), .Z(n9194) );
  XOR U8871 ( .A(n9198), .B(n9199), .Z(n9192) );
  AND U8872 ( .A(n317), .B(n9191), .Z(n9199) );
  XNOR U8873 ( .A(n9189), .B(n9198), .Z(n9191) );
  XNOR U8874 ( .A(n9200), .B(n9201), .Z(n9189) );
  AND U8875 ( .A(n321), .B(n9202), .Z(n9201) );
  XOR U8876 ( .A(p_input[349]), .B(n9200), .Z(n9202) );
  XNOR U8877 ( .A(n9203), .B(n9204), .Z(n9200) );
  AND U8878 ( .A(n325), .B(n9205), .Z(n9204) );
  XOR U8879 ( .A(n9206), .B(n9207), .Z(n9198) );
  AND U8880 ( .A(n329), .B(n9197), .Z(n9207) );
  XNOR U8881 ( .A(n9208), .B(n9195), .Z(n9197) );
  XOR U8882 ( .A(n9209), .B(n9210), .Z(n9195) );
  AND U8883 ( .A(n352), .B(n9211), .Z(n9210) );
  IV U8884 ( .A(n9206), .Z(n9208) );
  XOR U8885 ( .A(n9212), .B(n9213), .Z(n9206) );
  AND U8886 ( .A(n336), .B(n9205), .Z(n9213) );
  XNOR U8887 ( .A(n9203), .B(n9212), .Z(n9205) );
  XNOR U8888 ( .A(n9214), .B(n9215), .Z(n9203) );
  AND U8889 ( .A(n340), .B(n9216), .Z(n9215) );
  XOR U8890 ( .A(p_input[381]), .B(n9214), .Z(n9216) );
  XNOR U8891 ( .A(n9217), .B(n9218), .Z(n9214) );
  AND U8892 ( .A(n344), .B(n9219), .Z(n9218) );
  XOR U8893 ( .A(n9220), .B(n9221), .Z(n9212) );
  AND U8894 ( .A(n348), .B(n9211), .Z(n9221) );
  XNOR U8895 ( .A(n9222), .B(n9209), .Z(n9211) );
  XOR U8896 ( .A(n9223), .B(n9224), .Z(n9209) );
  AND U8897 ( .A(n371), .B(n9225), .Z(n9224) );
  IV U8898 ( .A(n9220), .Z(n9222) );
  XOR U8899 ( .A(n9226), .B(n9227), .Z(n9220) );
  AND U8900 ( .A(n355), .B(n9219), .Z(n9227) );
  XNOR U8901 ( .A(n9217), .B(n9226), .Z(n9219) );
  XNOR U8902 ( .A(n9228), .B(n9229), .Z(n9217) );
  AND U8903 ( .A(n359), .B(n9230), .Z(n9229) );
  XOR U8904 ( .A(p_input[413]), .B(n9228), .Z(n9230) );
  XNOR U8905 ( .A(n9231), .B(n9232), .Z(n9228) );
  AND U8906 ( .A(n363), .B(n9233), .Z(n9232) );
  XOR U8907 ( .A(n9234), .B(n9235), .Z(n9226) );
  AND U8908 ( .A(n367), .B(n9225), .Z(n9235) );
  XNOR U8909 ( .A(n9236), .B(n9223), .Z(n9225) );
  XOR U8910 ( .A(n9237), .B(n9238), .Z(n9223) );
  AND U8911 ( .A(n390), .B(n9239), .Z(n9238) );
  IV U8912 ( .A(n9234), .Z(n9236) );
  XOR U8913 ( .A(n9240), .B(n9241), .Z(n9234) );
  AND U8914 ( .A(n374), .B(n9233), .Z(n9241) );
  XNOR U8915 ( .A(n9231), .B(n9240), .Z(n9233) );
  XNOR U8916 ( .A(n9242), .B(n9243), .Z(n9231) );
  AND U8917 ( .A(n378), .B(n9244), .Z(n9243) );
  XOR U8918 ( .A(p_input[445]), .B(n9242), .Z(n9244) );
  XNOR U8919 ( .A(n9245), .B(n9246), .Z(n9242) );
  AND U8920 ( .A(n382), .B(n9247), .Z(n9246) );
  XOR U8921 ( .A(n9248), .B(n9249), .Z(n9240) );
  AND U8922 ( .A(n386), .B(n9239), .Z(n9249) );
  XNOR U8923 ( .A(n9250), .B(n9237), .Z(n9239) );
  XOR U8924 ( .A(n9251), .B(n9252), .Z(n9237) );
  AND U8925 ( .A(n409), .B(n9253), .Z(n9252) );
  IV U8926 ( .A(n9248), .Z(n9250) );
  XOR U8927 ( .A(n9254), .B(n9255), .Z(n9248) );
  AND U8928 ( .A(n393), .B(n9247), .Z(n9255) );
  XNOR U8929 ( .A(n9245), .B(n9254), .Z(n9247) );
  XNOR U8930 ( .A(n9256), .B(n9257), .Z(n9245) );
  AND U8931 ( .A(n397), .B(n9258), .Z(n9257) );
  XOR U8932 ( .A(p_input[477]), .B(n9256), .Z(n9258) );
  XNOR U8933 ( .A(n9259), .B(n9260), .Z(n9256) );
  AND U8934 ( .A(n401), .B(n9261), .Z(n9260) );
  XOR U8935 ( .A(n9262), .B(n9263), .Z(n9254) );
  AND U8936 ( .A(n405), .B(n9253), .Z(n9263) );
  XNOR U8937 ( .A(n9264), .B(n9251), .Z(n9253) );
  XOR U8938 ( .A(n9265), .B(n9266), .Z(n9251) );
  AND U8939 ( .A(n428), .B(n9267), .Z(n9266) );
  IV U8940 ( .A(n9262), .Z(n9264) );
  XOR U8941 ( .A(n9268), .B(n9269), .Z(n9262) );
  AND U8942 ( .A(n412), .B(n9261), .Z(n9269) );
  XNOR U8943 ( .A(n9259), .B(n9268), .Z(n9261) );
  XNOR U8944 ( .A(n9270), .B(n9271), .Z(n9259) );
  AND U8945 ( .A(n416), .B(n9272), .Z(n9271) );
  XOR U8946 ( .A(p_input[509]), .B(n9270), .Z(n9272) );
  XNOR U8947 ( .A(n9273), .B(n9274), .Z(n9270) );
  AND U8948 ( .A(n420), .B(n9275), .Z(n9274) );
  XOR U8949 ( .A(n9276), .B(n9277), .Z(n9268) );
  AND U8950 ( .A(n424), .B(n9267), .Z(n9277) );
  XNOR U8951 ( .A(n9278), .B(n9265), .Z(n9267) );
  XOR U8952 ( .A(n9279), .B(n9280), .Z(n9265) );
  AND U8953 ( .A(n447), .B(n9281), .Z(n9280) );
  IV U8954 ( .A(n9276), .Z(n9278) );
  XOR U8955 ( .A(n9282), .B(n9283), .Z(n9276) );
  AND U8956 ( .A(n431), .B(n9275), .Z(n9283) );
  XNOR U8957 ( .A(n9273), .B(n9282), .Z(n9275) );
  XNOR U8958 ( .A(n9284), .B(n9285), .Z(n9273) );
  AND U8959 ( .A(n435), .B(n9286), .Z(n9285) );
  XOR U8960 ( .A(p_input[541]), .B(n9284), .Z(n9286) );
  XNOR U8961 ( .A(n9287), .B(n9288), .Z(n9284) );
  AND U8962 ( .A(n439), .B(n9289), .Z(n9288) );
  XOR U8963 ( .A(n9290), .B(n9291), .Z(n9282) );
  AND U8964 ( .A(n443), .B(n9281), .Z(n9291) );
  XNOR U8965 ( .A(n9292), .B(n9279), .Z(n9281) );
  XOR U8966 ( .A(n9293), .B(n9294), .Z(n9279) );
  AND U8967 ( .A(n466), .B(n9295), .Z(n9294) );
  IV U8968 ( .A(n9290), .Z(n9292) );
  XOR U8969 ( .A(n9296), .B(n9297), .Z(n9290) );
  AND U8970 ( .A(n450), .B(n9289), .Z(n9297) );
  XNOR U8971 ( .A(n9287), .B(n9296), .Z(n9289) );
  XNOR U8972 ( .A(n9298), .B(n9299), .Z(n9287) );
  AND U8973 ( .A(n454), .B(n9300), .Z(n9299) );
  XOR U8974 ( .A(p_input[573]), .B(n9298), .Z(n9300) );
  XNOR U8975 ( .A(n9301), .B(n9302), .Z(n9298) );
  AND U8976 ( .A(n458), .B(n9303), .Z(n9302) );
  XOR U8977 ( .A(n9304), .B(n9305), .Z(n9296) );
  AND U8978 ( .A(n462), .B(n9295), .Z(n9305) );
  XNOR U8979 ( .A(n9306), .B(n9293), .Z(n9295) );
  XOR U8980 ( .A(n9307), .B(n9308), .Z(n9293) );
  AND U8981 ( .A(n485), .B(n9309), .Z(n9308) );
  IV U8982 ( .A(n9304), .Z(n9306) );
  XOR U8983 ( .A(n9310), .B(n9311), .Z(n9304) );
  AND U8984 ( .A(n469), .B(n9303), .Z(n9311) );
  XNOR U8985 ( .A(n9301), .B(n9310), .Z(n9303) );
  XNOR U8986 ( .A(n9312), .B(n9313), .Z(n9301) );
  AND U8987 ( .A(n473), .B(n9314), .Z(n9313) );
  XOR U8988 ( .A(p_input[605]), .B(n9312), .Z(n9314) );
  XNOR U8989 ( .A(n9315), .B(n9316), .Z(n9312) );
  AND U8990 ( .A(n477), .B(n9317), .Z(n9316) );
  XOR U8991 ( .A(n9318), .B(n9319), .Z(n9310) );
  AND U8992 ( .A(n481), .B(n9309), .Z(n9319) );
  XNOR U8993 ( .A(n9320), .B(n9307), .Z(n9309) );
  XOR U8994 ( .A(n9321), .B(n9322), .Z(n9307) );
  AND U8995 ( .A(n504), .B(n9323), .Z(n9322) );
  IV U8996 ( .A(n9318), .Z(n9320) );
  XOR U8997 ( .A(n9324), .B(n9325), .Z(n9318) );
  AND U8998 ( .A(n488), .B(n9317), .Z(n9325) );
  XNOR U8999 ( .A(n9315), .B(n9324), .Z(n9317) );
  XNOR U9000 ( .A(n9326), .B(n9327), .Z(n9315) );
  AND U9001 ( .A(n492), .B(n9328), .Z(n9327) );
  XOR U9002 ( .A(p_input[637]), .B(n9326), .Z(n9328) );
  XNOR U9003 ( .A(n9329), .B(n9330), .Z(n9326) );
  AND U9004 ( .A(n496), .B(n9331), .Z(n9330) );
  XOR U9005 ( .A(n9332), .B(n9333), .Z(n9324) );
  AND U9006 ( .A(n500), .B(n9323), .Z(n9333) );
  XNOR U9007 ( .A(n9334), .B(n9321), .Z(n9323) );
  XOR U9008 ( .A(n9335), .B(n9336), .Z(n9321) );
  AND U9009 ( .A(n523), .B(n9337), .Z(n9336) );
  IV U9010 ( .A(n9332), .Z(n9334) );
  XOR U9011 ( .A(n9338), .B(n9339), .Z(n9332) );
  AND U9012 ( .A(n507), .B(n9331), .Z(n9339) );
  XNOR U9013 ( .A(n9329), .B(n9338), .Z(n9331) );
  XNOR U9014 ( .A(n9340), .B(n9341), .Z(n9329) );
  AND U9015 ( .A(n511), .B(n9342), .Z(n9341) );
  XOR U9016 ( .A(p_input[669]), .B(n9340), .Z(n9342) );
  XNOR U9017 ( .A(n9343), .B(n9344), .Z(n9340) );
  AND U9018 ( .A(n515), .B(n9345), .Z(n9344) );
  XOR U9019 ( .A(n9346), .B(n9347), .Z(n9338) );
  AND U9020 ( .A(n519), .B(n9337), .Z(n9347) );
  XNOR U9021 ( .A(n9348), .B(n9335), .Z(n9337) );
  XOR U9022 ( .A(n9349), .B(n9350), .Z(n9335) );
  AND U9023 ( .A(n542), .B(n9351), .Z(n9350) );
  IV U9024 ( .A(n9346), .Z(n9348) );
  XOR U9025 ( .A(n9352), .B(n9353), .Z(n9346) );
  AND U9026 ( .A(n526), .B(n9345), .Z(n9353) );
  XNOR U9027 ( .A(n9343), .B(n9352), .Z(n9345) );
  XNOR U9028 ( .A(n9354), .B(n9355), .Z(n9343) );
  AND U9029 ( .A(n530), .B(n9356), .Z(n9355) );
  XOR U9030 ( .A(p_input[701]), .B(n9354), .Z(n9356) );
  XNOR U9031 ( .A(n9357), .B(n9358), .Z(n9354) );
  AND U9032 ( .A(n534), .B(n9359), .Z(n9358) );
  XOR U9033 ( .A(n9360), .B(n9361), .Z(n9352) );
  AND U9034 ( .A(n538), .B(n9351), .Z(n9361) );
  XNOR U9035 ( .A(n9362), .B(n9349), .Z(n9351) );
  XOR U9036 ( .A(n9363), .B(n9364), .Z(n9349) );
  AND U9037 ( .A(n561), .B(n9365), .Z(n9364) );
  IV U9038 ( .A(n9360), .Z(n9362) );
  XOR U9039 ( .A(n9366), .B(n9367), .Z(n9360) );
  AND U9040 ( .A(n545), .B(n9359), .Z(n9367) );
  XNOR U9041 ( .A(n9357), .B(n9366), .Z(n9359) );
  XNOR U9042 ( .A(n9368), .B(n9369), .Z(n9357) );
  AND U9043 ( .A(n549), .B(n9370), .Z(n9369) );
  XOR U9044 ( .A(p_input[733]), .B(n9368), .Z(n9370) );
  XNOR U9045 ( .A(n9371), .B(n9372), .Z(n9368) );
  AND U9046 ( .A(n553), .B(n9373), .Z(n9372) );
  XOR U9047 ( .A(n9374), .B(n9375), .Z(n9366) );
  AND U9048 ( .A(n557), .B(n9365), .Z(n9375) );
  XNOR U9049 ( .A(n9376), .B(n9363), .Z(n9365) );
  XOR U9050 ( .A(n9377), .B(n9378), .Z(n9363) );
  AND U9051 ( .A(n580), .B(n9379), .Z(n9378) );
  IV U9052 ( .A(n9374), .Z(n9376) );
  XOR U9053 ( .A(n9380), .B(n9381), .Z(n9374) );
  AND U9054 ( .A(n564), .B(n9373), .Z(n9381) );
  XNOR U9055 ( .A(n9371), .B(n9380), .Z(n9373) );
  XNOR U9056 ( .A(n9382), .B(n9383), .Z(n9371) );
  AND U9057 ( .A(n568), .B(n9384), .Z(n9383) );
  XOR U9058 ( .A(p_input[765]), .B(n9382), .Z(n9384) );
  XNOR U9059 ( .A(n9385), .B(n9386), .Z(n9382) );
  AND U9060 ( .A(n572), .B(n9387), .Z(n9386) );
  XOR U9061 ( .A(n9388), .B(n9389), .Z(n9380) );
  AND U9062 ( .A(n576), .B(n9379), .Z(n9389) );
  XNOR U9063 ( .A(n9390), .B(n9377), .Z(n9379) );
  XOR U9064 ( .A(n9391), .B(n9392), .Z(n9377) );
  AND U9065 ( .A(n599), .B(n9393), .Z(n9392) );
  IV U9066 ( .A(n9388), .Z(n9390) );
  XOR U9067 ( .A(n9394), .B(n9395), .Z(n9388) );
  AND U9068 ( .A(n583), .B(n9387), .Z(n9395) );
  XNOR U9069 ( .A(n9385), .B(n9394), .Z(n9387) );
  XNOR U9070 ( .A(n9396), .B(n9397), .Z(n9385) );
  AND U9071 ( .A(n587), .B(n9398), .Z(n9397) );
  XOR U9072 ( .A(p_input[797]), .B(n9396), .Z(n9398) );
  XNOR U9073 ( .A(n9399), .B(n9400), .Z(n9396) );
  AND U9074 ( .A(n591), .B(n9401), .Z(n9400) );
  XOR U9075 ( .A(n9402), .B(n9403), .Z(n9394) );
  AND U9076 ( .A(n595), .B(n9393), .Z(n9403) );
  XNOR U9077 ( .A(n9404), .B(n9391), .Z(n9393) );
  XOR U9078 ( .A(n9405), .B(n9406), .Z(n9391) );
  AND U9079 ( .A(n618), .B(n9407), .Z(n9406) );
  IV U9080 ( .A(n9402), .Z(n9404) );
  XOR U9081 ( .A(n9408), .B(n9409), .Z(n9402) );
  AND U9082 ( .A(n602), .B(n9401), .Z(n9409) );
  XNOR U9083 ( .A(n9399), .B(n9408), .Z(n9401) );
  XNOR U9084 ( .A(n9410), .B(n9411), .Z(n9399) );
  AND U9085 ( .A(n606), .B(n9412), .Z(n9411) );
  XOR U9086 ( .A(p_input[829]), .B(n9410), .Z(n9412) );
  XNOR U9087 ( .A(n9413), .B(n9414), .Z(n9410) );
  AND U9088 ( .A(n610), .B(n9415), .Z(n9414) );
  XOR U9089 ( .A(n9416), .B(n9417), .Z(n9408) );
  AND U9090 ( .A(n614), .B(n9407), .Z(n9417) );
  XNOR U9091 ( .A(n9418), .B(n9405), .Z(n9407) );
  XOR U9092 ( .A(n9419), .B(n9420), .Z(n9405) );
  AND U9093 ( .A(n637), .B(n9421), .Z(n9420) );
  IV U9094 ( .A(n9416), .Z(n9418) );
  XOR U9095 ( .A(n9422), .B(n9423), .Z(n9416) );
  AND U9096 ( .A(n621), .B(n9415), .Z(n9423) );
  XNOR U9097 ( .A(n9413), .B(n9422), .Z(n9415) );
  XNOR U9098 ( .A(n9424), .B(n9425), .Z(n9413) );
  AND U9099 ( .A(n625), .B(n9426), .Z(n9425) );
  XOR U9100 ( .A(p_input[861]), .B(n9424), .Z(n9426) );
  XNOR U9101 ( .A(n9427), .B(n9428), .Z(n9424) );
  AND U9102 ( .A(n629), .B(n9429), .Z(n9428) );
  XOR U9103 ( .A(n9430), .B(n9431), .Z(n9422) );
  AND U9104 ( .A(n633), .B(n9421), .Z(n9431) );
  XNOR U9105 ( .A(n9432), .B(n9419), .Z(n9421) );
  XOR U9106 ( .A(n9433), .B(n9434), .Z(n9419) );
  AND U9107 ( .A(n656), .B(n9435), .Z(n9434) );
  IV U9108 ( .A(n9430), .Z(n9432) );
  XOR U9109 ( .A(n9436), .B(n9437), .Z(n9430) );
  AND U9110 ( .A(n640), .B(n9429), .Z(n9437) );
  XNOR U9111 ( .A(n9427), .B(n9436), .Z(n9429) );
  XNOR U9112 ( .A(n9438), .B(n9439), .Z(n9427) );
  AND U9113 ( .A(n644), .B(n9440), .Z(n9439) );
  XOR U9114 ( .A(p_input[893]), .B(n9438), .Z(n9440) );
  XNOR U9115 ( .A(n9441), .B(n9442), .Z(n9438) );
  AND U9116 ( .A(n648), .B(n9443), .Z(n9442) );
  XOR U9117 ( .A(n9444), .B(n9445), .Z(n9436) );
  AND U9118 ( .A(n652), .B(n9435), .Z(n9445) );
  XNOR U9119 ( .A(n9446), .B(n9433), .Z(n9435) );
  XOR U9120 ( .A(n9447), .B(n9448), .Z(n9433) );
  AND U9121 ( .A(n675), .B(n9449), .Z(n9448) );
  IV U9122 ( .A(n9444), .Z(n9446) );
  XOR U9123 ( .A(n9450), .B(n9451), .Z(n9444) );
  AND U9124 ( .A(n659), .B(n9443), .Z(n9451) );
  XNOR U9125 ( .A(n9441), .B(n9450), .Z(n9443) );
  XNOR U9126 ( .A(n9452), .B(n9453), .Z(n9441) );
  AND U9127 ( .A(n663), .B(n9454), .Z(n9453) );
  XOR U9128 ( .A(p_input[925]), .B(n9452), .Z(n9454) );
  XNOR U9129 ( .A(n9455), .B(n9456), .Z(n9452) );
  AND U9130 ( .A(n667), .B(n9457), .Z(n9456) );
  XOR U9131 ( .A(n9458), .B(n9459), .Z(n9450) );
  AND U9132 ( .A(n671), .B(n9449), .Z(n9459) );
  XNOR U9133 ( .A(n9460), .B(n9447), .Z(n9449) );
  XOR U9134 ( .A(n9461), .B(n9462), .Z(n9447) );
  AND U9135 ( .A(n694), .B(n9463), .Z(n9462) );
  IV U9136 ( .A(n9458), .Z(n9460) );
  XOR U9137 ( .A(n9464), .B(n9465), .Z(n9458) );
  AND U9138 ( .A(n678), .B(n9457), .Z(n9465) );
  XNOR U9139 ( .A(n9455), .B(n9464), .Z(n9457) );
  XNOR U9140 ( .A(n9466), .B(n9467), .Z(n9455) );
  AND U9141 ( .A(n682), .B(n9468), .Z(n9467) );
  XOR U9142 ( .A(p_input[957]), .B(n9466), .Z(n9468) );
  XNOR U9143 ( .A(n9469), .B(n9470), .Z(n9466) );
  AND U9144 ( .A(n686), .B(n9471), .Z(n9470) );
  XOR U9145 ( .A(n9472), .B(n9473), .Z(n9464) );
  AND U9146 ( .A(n690), .B(n9463), .Z(n9473) );
  XNOR U9147 ( .A(n9474), .B(n9461), .Z(n9463) );
  XOR U9148 ( .A(n9475), .B(n9476), .Z(n9461) );
  AND U9149 ( .A(n713), .B(n9477), .Z(n9476) );
  IV U9150 ( .A(n9472), .Z(n9474) );
  XOR U9151 ( .A(n9478), .B(n9479), .Z(n9472) );
  AND U9152 ( .A(n697), .B(n9471), .Z(n9479) );
  XNOR U9153 ( .A(n9469), .B(n9478), .Z(n9471) );
  XNOR U9154 ( .A(n9480), .B(n9481), .Z(n9469) );
  AND U9155 ( .A(n701), .B(n9482), .Z(n9481) );
  XOR U9156 ( .A(p_input[989]), .B(n9480), .Z(n9482) );
  XNOR U9157 ( .A(n9483), .B(n9484), .Z(n9480) );
  AND U9158 ( .A(n705), .B(n9485), .Z(n9484) );
  XOR U9159 ( .A(n9486), .B(n9487), .Z(n9478) );
  AND U9160 ( .A(n709), .B(n9477), .Z(n9487) );
  XNOR U9161 ( .A(n9488), .B(n9475), .Z(n9477) );
  XOR U9162 ( .A(n9489), .B(n9490), .Z(n9475) );
  AND U9163 ( .A(n732), .B(n9491), .Z(n9490) );
  IV U9164 ( .A(n9486), .Z(n9488) );
  XOR U9165 ( .A(n9492), .B(n9493), .Z(n9486) );
  AND U9166 ( .A(n716), .B(n9485), .Z(n9493) );
  XNOR U9167 ( .A(n9483), .B(n9492), .Z(n9485) );
  XNOR U9168 ( .A(n9494), .B(n9495), .Z(n9483) );
  AND U9169 ( .A(n720), .B(n9496), .Z(n9495) );
  XOR U9170 ( .A(p_input[1021]), .B(n9494), .Z(n9496) );
  XNOR U9171 ( .A(n9497), .B(n9498), .Z(n9494) );
  AND U9172 ( .A(n724), .B(n9499), .Z(n9498) );
  XOR U9173 ( .A(n9500), .B(n9501), .Z(n9492) );
  AND U9174 ( .A(n728), .B(n9491), .Z(n9501) );
  XNOR U9175 ( .A(n9502), .B(n9489), .Z(n9491) );
  XOR U9176 ( .A(n9503), .B(n9504), .Z(n9489) );
  AND U9177 ( .A(n751), .B(n9505), .Z(n9504) );
  IV U9178 ( .A(n9500), .Z(n9502) );
  XOR U9179 ( .A(n9506), .B(n9507), .Z(n9500) );
  AND U9180 ( .A(n735), .B(n9499), .Z(n9507) );
  XNOR U9181 ( .A(n9497), .B(n9506), .Z(n9499) );
  XNOR U9182 ( .A(n9508), .B(n9509), .Z(n9497) );
  AND U9183 ( .A(n739), .B(n9510), .Z(n9509) );
  XOR U9184 ( .A(p_input[1053]), .B(n9508), .Z(n9510) );
  XNOR U9185 ( .A(n9511), .B(n9512), .Z(n9508) );
  AND U9186 ( .A(n743), .B(n9513), .Z(n9512) );
  XOR U9187 ( .A(n9514), .B(n9515), .Z(n9506) );
  AND U9188 ( .A(n747), .B(n9505), .Z(n9515) );
  XNOR U9189 ( .A(n9516), .B(n9503), .Z(n9505) );
  XOR U9190 ( .A(n9517), .B(n9518), .Z(n9503) );
  AND U9191 ( .A(n770), .B(n9519), .Z(n9518) );
  IV U9192 ( .A(n9514), .Z(n9516) );
  XOR U9193 ( .A(n9520), .B(n9521), .Z(n9514) );
  AND U9194 ( .A(n754), .B(n9513), .Z(n9521) );
  XNOR U9195 ( .A(n9511), .B(n9520), .Z(n9513) );
  XNOR U9196 ( .A(n9522), .B(n9523), .Z(n9511) );
  AND U9197 ( .A(n758), .B(n9524), .Z(n9523) );
  XOR U9198 ( .A(p_input[1085]), .B(n9522), .Z(n9524) );
  XNOR U9199 ( .A(n9525), .B(n9526), .Z(n9522) );
  AND U9200 ( .A(n762), .B(n9527), .Z(n9526) );
  XOR U9201 ( .A(n9528), .B(n9529), .Z(n9520) );
  AND U9202 ( .A(n766), .B(n9519), .Z(n9529) );
  XNOR U9203 ( .A(n9530), .B(n9517), .Z(n9519) );
  XOR U9204 ( .A(n9531), .B(n9532), .Z(n9517) );
  AND U9205 ( .A(n789), .B(n9533), .Z(n9532) );
  IV U9206 ( .A(n9528), .Z(n9530) );
  XOR U9207 ( .A(n9534), .B(n9535), .Z(n9528) );
  AND U9208 ( .A(n773), .B(n9527), .Z(n9535) );
  XNOR U9209 ( .A(n9525), .B(n9534), .Z(n9527) );
  XNOR U9210 ( .A(n9536), .B(n9537), .Z(n9525) );
  AND U9211 ( .A(n777), .B(n9538), .Z(n9537) );
  XOR U9212 ( .A(p_input[1117]), .B(n9536), .Z(n9538) );
  XNOR U9213 ( .A(n9539), .B(n9540), .Z(n9536) );
  AND U9214 ( .A(n781), .B(n9541), .Z(n9540) );
  XOR U9215 ( .A(n9542), .B(n9543), .Z(n9534) );
  AND U9216 ( .A(n785), .B(n9533), .Z(n9543) );
  XNOR U9217 ( .A(n9544), .B(n9531), .Z(n9533) );
  XOR U9218 ( .A(n9545), .B(n9546), .Z(n9531) );
  AND U9219 ( .A(n808), .B(n9547), .Z(n9546) );
  IV U9220 ( .A(n9542), .Z(n9544) );
  XOR U9221 ( .A(n9548), .B(n9549), .Z(n9542) );
  AND U9222 ( .A(n792), .B(n9541), .Z(n9549) );
  XNOR U9223 ( .A(n9539), .B(n9548), .Z(n9541) );
  XNOR U9224 ( .A(n9550), .B(n9551), .Z(n9539) );
  AND U9225 ( .A(n796), .B(n9552), .Z(n9551) );
  XOR U9226 ( .A(p_input[1149]), .B(n9550), .Z(n9552) );
  XNOR U9227 ( .A(n9553), .B(n9554), .Z(n9550) );
  AND U9228 ( .A(n800), .B(n9555), .Z(n9554) );
  XOR U9229 ( .A(n9556), .B(n9557), .Z(n9548) );
  AND U9230 ( .A(n804), .B(n9547), .Z(n9557) );
  XNOR U9231 ( .A(n9558), .B(n9545), .Z(n9547) );
  XOR U9232 ( .A(n9559), .B(n9560), .Z(n9545) );
  AND U9233 ( .A(n827), .B(n9561), .Z(n9560) );
  IV U9234 ( .A(n9556), .Z(n9558) );
  XOR U9235 ( .A(n9562), .B(n9563), .Z(n9556) );
  AND U9236 ( .A(n811), .B(n9555), .Z(n9563) );
  XNOR U9237 ( .A(n9553), .B(n9562), .Z(n9555) );
  XNOR U9238 ( .A(n9564), .B(n9565), .Z(n9553) );
  AND U9239 ( .A(n815), .B(n9566), .Z(n9565) );
  XOR U9240 ( .A(p_input[1181]), .B(n9564), .Z(n9566) );
  XNOR U9241 ( .A(n9567), .B(n9568), .Z(n9564) );
  AND U9242 ( .A(n819), .B(n9569), .Z(n9568) );
  XOR U9243 ( .A(n9570), .B(n9571), .Z(n9562) );
  AND U9244 ( .A(n823), .B(n9561), .Z(n9571) );
  XNOR U9245 ( .A(n9572), .B(n9559), .Z(n9561) );
  XOR U9246 ( .A(n9573), .B(n9574), .Z(n9559) );
  AND U9247 ( .A(n846), .B(n9575), .Z(n9574) );
  IV U9248 ( .A(n9570), .Z(n9572) );
  XOR U9249 ( .A(n9576), .B(n9577), .Z(n9570) );
  AND U9250 ( .A(n830), .B(n9569), .Z(n9577) );
  XNOR U9251 ( .A(n9567), .B(n9576), .Z(n9569) );
  XNOR U9252 ( .A(n9578), .B(n9579), .Z(n9567) );
  AND U9253 ( .A(n834), .B(n9580), .Z(n9579) );
  XOR U9254 ( .A(p_input[1213]), .B(n9578), .Z(n9580) );
  XNOR U9255 ( .A(n9581), .B(n9582), .Z(n9578) );
  AND U9256 ( .A(n838), .B(n9583), .Z(n9582) );
  XOR U9257 ( .A(n9584), .B(n9585), .Z(n9576) );
  AND U9258 ( .A(n842), .B(n9575), .Z(n9585) );
  XNOR U9259 ( .A(n9586), .B(n9573), .Z(n9575) );
  XOR U9260 ( .A(n9587), .B(n9588), .Z(n9573) );
  AND U9261 ( .A(n865), .B(n9589), .Z(n9588) );
  IV U9262 ( .A(n9584), .Z(n9586) );
  XOR U9263 ( .A(n9590), .B(n9591), .Z(n9584) );
  AND U9264 ( .A(n849), .B(n9583), .Z(n9591) );
  XNOR U9265 ( .A(n9581), .B(n9590), .Z(n9583) );
  XNOR U9266 ( .A(n9592), .B(n9593), .Z(n9581) );
  AND U9267 ( .A(n853), .B(n9594), .Z(n9593) );
  XOR U9268 ( .A(p_input[1245]), .B(n9592), .Z(n9594) );
  XNOR U9269 ( .A(n9595), .B(n9596), .Z(n9592) );
  AND U9270 ( .A(n857), .B(n9597), .Z(n9596) );
  XOR U9271 ( .A(n9598), .B(n9599), .Z(n9590) );
  AND U9272 ( .A(n861), .B(n9589), .Z(n9599) );
  XNOR U9273 ( .A(n9600), .B(n9587), .Z(n9589) );
  XOR U9274 ( .A(n9601), .B(n9602), .Z(n9587) );
  AND U9275 ( .A(n884), .B(n9603), .Z(n9602) );
  IV U9276 ( .A(n9598), .Z(n9600) );
  XOR U9277 ( .A(n9604), .B(n9605), .Z(n9598) );
  AND U9278 ( .A(n868), .B(n9597), .Z(n9605) );
  XNOR U9279 ( .A(n9595), .B(n9604), .Z(n9597) );
  XNOR U9280 ( .A(n9606), .B(n9607), .Z(n9595) );
  AND U9281 ( .A(n872), .B(n9608), .Z(n9607) );
  XOR U9282 ( .A(p_input[1277]), .B(n9606), .Z(n9608) );
  XNOR U9283 ( .A(n9609), .B(n9610), .Z(n9606) );
  AND U9284 ( .A(n876), .B(n9611), .Z(n9610) );
  XOR U9285 ( .A(n9612), .B(n9613), .Z(n9604) );
  AND U9286 ( .A(n880), .B(n9603), .Z(n9613) );
  XNOR U9287 ( .A(n9614), .B(n9601), .Z(n9603) );
  XOR U9288 ( .A(n9615), .B(n9616), .Z(n9601) );
  AND U9289 ( .A(n903), .B(n9617), .Z(n9616) );
  IV U9290 ( .A(n9612), .Z(n9614) );
  XOR U9291 ( .A(n9618), .B(n9619), .Z(n9612) );
  AND U9292 ( .A(n887), .B(n9611), .Z(n9619) );
  XNOR U9293 ( .A(n9609), .B(n9618), .Z(n9611) );
  XNOR U9294 ( .A(n9620), .B(n9621), .Z(n9609) );
  AND U9295 ( .A(n891), .B(n9622), .Z(n9621) );
  XOR U9296 ( .A(p_input[1309]), .B(n9620), .Z(n9622) );
  XNOR U9297 ( .A(n9623), .B(n9624), .Z(n9620) );
  AND U9298 ( .A(n895), .B(n9625), .Z(n9624) );
  XOR U9299 ( .A(n9626), .B(n9627), .Z(n9618) );
  AND U9300 ( .A(n899), .B(n9617), .Z(n9627) );
  XNOR U9301 ( .A(n9628), .B(n9615), .Z(n9617) );
  XOR U9302 ( .A(n9629), .B(n9630), .Z(n9615) );
  AND U9303 ( .A(n922), .B(n9631), .Z(n9630) );
  IV U9304 ( .A(n9626), .Z(n9628) );
  XOR U9305 ( .A(n9632), .B(n9633), .Z(n9626) );
  AND U9306 ( .A(n906), .B(n9625), .Z(n9633) );
  XNOR U9307 ( .A(n9623), .B(n9632), .Z(n9625) );
  XNOR U9308 ( .A(n9634), .B(n9635), .Z(n9623) );
  AND U9309 ( .A(n910), .B(n9636), .Z(n9635) );
  XOR U9310 ( .A(p_input[1341]), .B(n9634), .Z(n9636) );
  XNOR U9311 ( .A(n9637), .B(n9638), .Z(n9634) );
  AND U9312 ( .A(n914), .B(n9639), .Z(n9638) );
  XOR U9313 ( .A(n9640), .B(n9641), .Z(n9632) );
  AND U9314 ( .A(n918), .B(n9631), .Z(n9641) );
  XNOR U9315 ( .A(n9642), .B(n9629), .Z(n9631) );
  XOR U9316 ( .A(n9643), .B(n9644), .Z(n9629) );
  AND U9317 ( .A(n941), .B(n9645), .Z(n9644) );
  IV U9318 ( .A(n9640), .Z(n9642) );
  XOR U9319 ( .A(n9646), .B(n9647), .Z(n9640) );
  AND U9320 ( .A(n925), .B(n9639), .Z(n9647) );
  XNOR U9321 ( .A(n9637), .B(n9646), .Z(n9639) );
  XNOR U9322 ( .A(n9648), .B(n9649), .Z(n9637) );
  AND U9323 ( .A(n929), .B(n9650), .Z(n9649) );
  XOR U9324 ( .A(p_input[1373]), .B(n9648), .Z(n9650) );
  XNOR U9325 ( .A(n9651), .B(n9652), .Z(n9648) );
  AND U9326 ( .A(n933), .B(n9653), .Z(n9652) );
  XOR U9327 ( .A(n9654), .B(n9655), .Z(n9646) );
  AND U9328 ( .A(n937), .B(n9645), .Z(n9655) );
  XNOR U9329 ( .A(n9656), .B(n9643), .Z(n9645) );
  XOR U9330 ( .A(n9657), .B(n9658), .Z(n9643) );
  AND U9331 ( .A(n960), .B(n9659), .Z(n9658) );
  IV U9332 ( .A(n9654), .Z(n9656) );
  XOR U9333 ( .A(n9660), .B(n9661), .Z(n9654) );
  AND U9334 ( .A(n944), .B(n9653), .Z(n9661) );
  XNOR U9335 ( .A(n9651), .B(n9660), .Z(n9653) );
  XNOR U9336 ( .A(n9662), .B(n9663), .Z(n9651) );
  AND U9337 ( .A(n948), .B(n9664), .Z(n9663) );
  XOR U9338 ( .A(p_input[1405]), .B(n9662), .Z(n9664) );
  XNOR U9339 ( .A(n9665), .B(n9666), .Z(n9662) );
  AND U9340 ( .A(n952), .B(n9667), .Z(n9666) );
  XOR U9341 ( .A(n9668), .B(n9669), .Z(n9660) );
  AND U9342 ( .A(n956), .B(n9659), .Z(n9669) );
  XNOR U9343 ( .A(n9670), .B(n9657), .Z(n9659) );
  XOR U9344 ( .A(n9671), .B(n9672), .Z(n9657) );
  AND U9345 ( .A(n979), .B(n9673), .Z(n9672) );
  IV U9346 ( .A(n9668), .Z(n9670) );
  XOR U9347 ( .A(n9674), .B(n9675), .Z(n9668) );
  AND U9348 ( .A(n963), .B(n9667), .Z(n9675) );
  XNOR U9349 ( .A(n9665), .B(n9674), .Z(n9667) );
  XNOR U9350 ( .A(n9676), .B(n9677), .Z(n9665) );
  AND U9351 ( .A(n967), .B(n9678), .Z(n9677) );
  XOR U9352 ( .A(p_input[1437]), .B(n9676), .Z(n9678) );
  XNOR U9353 ( .A(n9679), .B(n9680), .Z(n9676) );
  AND U9354 ( .A(n971), .B(n9681), .Z(n9680) );
  XOR U9355 ( .A(n9682), .B(n9683), .Z(n9674) );
  AND U9356 ( .A(n975), .B(n9673), .Z(n9683) );
  XNOR U9357 ( .A(n9684), .B(n9671), .Z(n9673) );
  XOR U9358 ( .A(n9685), .B(n9686), .Z(n9671) );
  AND U9359 ( .A(n998), .B(n9687), .Z(n9686) );
  IV U9360 ( .A(n9682), .Z(n9684) );
  XOR U9361 ( .A(n9688), .B(n9689), .Z(n9682) );
  AND U9362 ( .A(n982), .B(n9681), .Z(n9689) );
  XNOR U9363 ( .A(n9679), .B(n9688), .Z(n9681) );
  XNOR U9364 ( .A(n9690), .B(n9691), .Z(n9679) );
  AND U9365 ( .A(n986), .B(n9692), .Z(n9691) );
  XOR U9366 ( .A(p_input[1469]), .B(n9690), .Z(n9692) );
  XNOR U9367 ( .A(n9693), .B(n9694), .Z(n9690) );
  AND U9368 ( .A(n990), .B(n9695), .Z(n9694) );
  XOR U9369 ( .A(n9696), .B(n9697), .Z(n9688) );
  AND U9370 ( .A(n994), .B(n9687), .Z(n9697) );
  XNOR U9371 ( .A(n9698), .B(n9685), .Z(n9687) );
  XOR U9372 ( .A(n9699), .B(n9700), .Z(n9685) );
  AND U9373 ( .A(n1017), .B(n9701), .Z(n9700) );
  IV U9374 ( .A(n9696), .Z(n9698) );
  XOR U9375 ( .A(n9702), .B(n9703), .Z(n9696) );
  AND U9376 ( .A(n1001), .B(n9695), .Z(n9703) );
  XNOR U9377 ( .A(n9693), .B(n9702), .Z(n9695) );
  XNOR U9378 ( .A(n9704), .B(n9705), .Z(n9693) );
  AND U9379 ( .A(n1005), .B(n9706), .Z(n9705) );
  XOR U9380 ( .A(p_input[1501]), .B(n9704), .Z(n9706) );
  XNOR U9381 ( .A(n9707), .B(n9708), .Z(n9704) );
  AND U9382 ( .A(n1009), .B(n9709), .Z(n9708) );
  XOR U9383 ( .A(n9710), .B(n9711), .Z(n9702) );
  AND U9384 ( .A(n1013), .B(n9701), .Z(n9711) );
  XNOR U9385 ( .A(n9712), .B(n9699), .Z(n9701) );
  XOR U9386 ( .A(n9713), .B(n9714), .Z(n9699) );
  AND U9387 ( .A(n1036), .B(n9715), .Z(n9714) );
  IV U9388 ( .A(n9710), .Z(n9712) );
  XOR U9389 ( .A(n9716), .B(n9717), .Z(n9710) );
  AND U9390 ( .A(n1020), .B(n9709), .Z(n9717) );
  XNOR U9391 ( .A(n9707), .B(n9716), .Z(n9709) );
  XNOR U9392 ( .A(n9718), .B(n9719), .Z(n9707) );
  AND U9393 ( .A(n1024), .B(n9720), .Z(n9719) );
  XOR U9394 ( .A(p_input[1533]), .B(n9718), .Z(n9720) );
  XNOR U9395 ( .A(n9721), .B(n9722), .Z(n9718) );
  AND U9396 ( .A(n1028), .B(n9723), .Z(n9722) );
  XOR U9397 ( .A(n9724), .B(n9725), .Z(n9716) );
  AND U9398 ( .A(n1032), .B(n9715), .Z(n9725) );
  XNOR U9399 ( .A(n9726), .B(n9713), .Z(n9715) );
  XOR U9400 ( .A(n9727), .B(n9728), .Z(n9713) );
  AND U9401 ( .A(n1055), .B(n9729), .Z(n9728) );
  IV U9402 ( .A(n9724), .Z(n9726) );
  XOR U9403 ( .A(n9730), .B(n9731), .Z(n9724) );
  AND U9404 ( .A(n1039), .B(n9723), .Z(n9731) );
  XNOR U9405 ( .A(n9721), .B(n9730), .Z(n9723) );
  XNOR U9406 ( .A(n9732), .B(n9733), .Z(n9721) );
  AND U9407 ( .A(n1043), .B(n9734), .Z(n9733) );
  XOR U9408 ( .A(p_input[1565]), .B(n9732), .Z(n9734) );
  XNOR U9409 ( .A(n9735), .B(n9736), .Z(n9732) );
  AND U9410 ( .A(n1047), .B(n9737), .Z(n9736) );
  XOR U9411 ( .A(n9738), .B(n9739), .Z(n9730) );
  AND U9412 ( .A(n1051), .B(n9729), .Z(n9739) );
  XNOR U9413 ( .A(n9740), .B(n9727), .Z(n9729) );
  XOR U9414 ( .A(n9741), .B(n9742), .Z(n9727) );
  AND U9415 ( .A(n1074), .B(n9743), .Z(n9742) );
  IV U9416 ( .A(n9738), .Z(n9740) );
  XOR U9417 ( .A(n9744), .B(n9745), .Z(n9738) );
  AND U9418 ( .A(n1058), .B(n9737), .Z(n9745) );
  XNOR U9419 ( .A(n9735), .B(n9744), .Z(n9737) );
  XNOR U9420 ( .A(n9746), .B(n9747), .Z(n9735) );
  AND U9421 ( .A(n1062), .B(n9748), .Z(n9747) );
  XOR U9422 ( .A(p_input[1597]), .B(n9746), .Z(n9748) );
  XNOR U9423 ( .A(n9749), .B(n9750), .Z(n9746) );
  AND U9424 ( .A(n1066), .B(n9751), .Z(n9750) );
  XOR U9425 ( .A(n9752), .B(n9753), .Z(n9744) );
  AND U9426 ( .A(n1070), .B(n9743), .Z(n9753) );
  XNOR U9427 ( .A(n9754), .B(n9741), .Z(n9743) );
  XOR U9428 ( .A(n9755), .B(n9756), .Z(n9741) );
  AND U9429 ( .A(n1093), .B(n9757), .Z(n9756) );
  IV U9430 ( .A(n9752), .Z(n9754) );
  XOR U9431 ( .A(n9758), .B(n9759), .Z(n9752) );
  AND U9432 ( .A(n1077), .B(n9751), .Z(n9759) );
  XNOR U9433 ( .A(n9749), .B(n9758), .Z(n9751) );
  XNOR U9434 ( .A(n9760), .B(n9761), .Z(n9749) );
  AND U9435 ( .A(n1081), .B(n9762), .Z(n9761) );
  XOR U9436 ( .A(p_input[1629]), .B(n9760), .Z(n9762) );
  XNOR U9437 ( .A(n9763), .B(n9764), .Z(n9760) );
  AND U9438 ( .A(n1085), .B(n9765), .Z(n9764) );
  XOR U9439 ( .A(n9766), .B(n9767), .Z(n9758) );
  AND U9440 ( .A(n1089), .B(n9757), .Z(n9767) );
  XNOR U9441 ( .A(n9768), .B(n9755), .Z(n9757) );
  XOR U9442 ( .A(n9769), .B(n9770), .Z(n9755) );
  AND U9443 ( .A(n1112), .B(n9771), .Z(n9770) );
  IV U9444 ( .A(n9766), .Z(n9768) );
  XOR U9445 ( .A(n9772), .B(n9773), .Z(n9766) );
  AND U9446 ( .A(n1096), .B(n9765), .Z(n9773) );
  XNOR U9447 ( .A(n9763), .B(n9772), .Z(n9765) );
  XNOR U9448 ( .A(n9774), .B(n9775), .Z(n9763) );
  AND U9449 ( .A(n1100), .B(n9776), .Z(n9775) );
  XOR U9450 ( .A(p_input[1661]), .B(n9774), .Z(n9776) );
  XNOR U9451 ( .A(n9777), .B(n9778), .Z(n9774) );
  AND U9452 ( .A(n1104), .B(n9779), .Z(n9778) );
  XOR U9453 ( .A(n9780), .B(n9781), .Z(n9772) );
  AND U9454 ( .A(n1108), .B(n9771), .Z(n9781) );
  XNOR U9455 ( .A(n9782), .B(n9769), .Z(n9771) );
  XOR U9456 ( .A(n9783), .B(n9784), .Z(n9769) );
  AND U9457 ( .A(n1131), .B(n9785), .Z(n9784) );
  IV U9458 ( .A(n9780), .Z(n9782) );
  XOR U9459 ( .A(n9786), .B(n9787), .Z(n9780) );
  AND U9460 ( .A(n1115), .B(n9779), .Z(n9787) );
  XNOR U9461 ( .A(n9777), .B(n9786), .Z(n9779) );
  XNOR U9462 ( .A(n9788), .B(n9789), .Z(n9777) );
  AND U9463 ( .A(n1119), .B(n9790), .Z(n9789) );
  XOR U9464 ( .A(p_input[1693]), .B(n9788), .Z(n9790) );
  XNOR U9465 ( .A(n9791), .B(n9792), .Z(n9788) );
  AND U9466 ( .A(n1123), .B(n9793), .Z(n9792) );
  XOR U9467 ( .A(n9794), .B(n9795), .Z(n9786) );
  AND U9468 ( .A(n1127), .B(n9785), .Z(n9795) );
  XNOR U9469 ( .A(n9796), .B(n9783), .Z(n9785) );
  XOR U9470 ( .A(n9797), .B(n9798), .Z(n9783) );
  AND U9471 ( .A(n1150), .B(n9799), .Z(n9798) );
  IV U9472 ( .A(n9794), .Z(n9796) );
  XOR U9473 ( .A(n9800), .B(n9801), .Z(n9794) );
  AND U9474 ( .A(n1134), .B(n9793), .Z(n9801) );
  XNOR U9475 ( .A(n9791), .B(n9800), .Z(n9793) );
  XNOR U9476 ( .A(n9802), .B(n9803), .Z(n9791) );
  AND U9477 ( .A(n1138), .B(n9804), .Z(n9803) );
  XOR U9478 ( .A(p_input[1725]), .B(n9802), .Z(n9804) );
  XNOR U9479 ( .A(n9805), .B(n9806), .Z(n9802) );
  AND U9480 ( .A(n1142), .B(n9807), .Z(n9806) );
  XOR U9481 ( .A(n9808), .B(n9809), .Z(n9800) );
  AND U9482 ( .A(n1146), .B(n9799), .Z(n9809) );
  XNOR U9483 ( .A(n9810), .B(n9797), .Z(n9799) );
  XOR U9484 ( .A(n9811), .B(n9812), .Z(n9797) );
  AND U9485 ( .A(n1169), .B(n9813), .Z(n9812) );
  IV U9486 ( .A(n9808), .Z(n9810) );
  XOR U9487 ( .A(n9814), .B(n9815), .Z(n9808) );
  AND U9488 ( .A(n1153), .B(n9807), .Z(n9815) );
  XNOR U9489 ( .A(n9805), .B(n9814), .Z(n9807) );
  XNOR U9490 ( .A(n9816), .B(n9817), .Z(n9805) );
  AND U9491 ( .A(n1157), .B(n9818), .Z(n9817) );
  XOR U9492 ( .A(p_input[1757]), .B(n9816), .Z(n9818) );
  XNOR U9493 ( .A(n9819), .B(n9820), .Z(n9816) );
  AND U9494 ( .A(n1161), .B(n9821), .Z(n9820) );
  XOR U9495 ( .A(n9822), .B(n9823), .Z(n9814) );
  AND U9496 ( .A(n1165), .B(n9813), .Z(n9823) );
  XNOR U9497 ( .A(n9824), .B(n9811), .Z(n9813) );
  XOR U9498 ( .A(n9825), .B(n9826), .Z(n9811) );
  AND U9499 ( .A(n1188), .B(n9827), .Z(n9826) );
  IV U9500 ( .A(n9822), .Z(n9824) );
  XOR U9501 ( .A(n9828), .B(n9829), .Z(n9822) );
  AND U9502 ( .A(n1172), .B(n9821), .Z(n9829) );
  XNOR U9503 ( .A(n9819), .B(n9828), .Z(n9821) );
  XNOR U9504 ( .A(n9830), .B(n9831), .Z(n9819) );
  AND U9505 ( .A(n1176), .B(n9832), .Z(n9831) );
  XOR U9506 ( .A(p_input[1789]), .B(n9830), .Z(n9832) );
  XNOR U9507 ( .A(n9833), .B(n9834), .Z(n9830) );
  AND U9508 ( .A(n1180), .B(n9835), .Z(n9834) );
  XOR U9509 ( .A(n9836), .B(n9837), .Z(n9828) );
  AND U9510 ( .A(n1184), .B(n9827), .Z(n9837) );
  XNOR U9511 ( .A(n9838), .B(n9825), .Z(n9827) );
  XOR U9512 ( .A(n9839), .B(n9840), .Z(n9825) );
  AND U9513 ( .A(n1207), .B(n9841), .Z(n9840) );
  IV U9514 ( .A(n9836), .Z(n9838) );
  XOR U9515 ( .A(n9842), .B(n9843), .Z(n9836) );
  AND U9516 ( .A(n1191), .B(n9835), .Z(n9843) );
  XNOR U9517 ( .A(n9833), .B(n9842), .Z(n9835) );
  XNOR U9518 ( .A(n9844), .B(n9845), .Z(n9833) );
  AND U9519 ( .A(n1195), .B(n9846), .Z(n9845) );
  XOR U9520 ( .A(p_input[1821]), .B(n9844), .Z(n9846) );
  XNOR U9521 ( .A(n9847), .B(n9848), .Z(n9844) );
  AND U9522 ( .A(n1199), .B(n9849), .Z(n9848) );
  XOR U9523 ( .A(n9850), .B(n9851), .Z(n9842) );
  AND U9524 ( .A(n1203), .B(n9841), .Z(n9851) );
  XNOR U9525 ( .A(n9852), .B(n9839), .Z(n9841) );
  XOR U9526 ( .A(n9853), .B(n9854), .Z(n9839) );
  AND U9527 ( .A(n1226), .B(n9855), .Z(n9854) );
  IV U9528 ( .A(n9850), .Z(n9852) );
  XOR U9529 ( .A(n9856), .B(n9857), .Z(n9850) );
  AND U9530 ( .A(n1210), .B(n9849), .Z(n9857) );
  XNOR U9531 ( .A(n9847), .B(n9856), .Z(n9849) );
  XNOR U9532 ( .A(n9858), .B(n9859), .Z(n9847) );
  AND U9533 ( .A(n1214), .B(n9860), .Z(n9859) );
  XOR U9534 ( .A(p_input[1853]), .B(n9858), .Z(n9860) );
  XNOR U9535 ( .A(n9861), .B(n9862), .Z(n9858) );
  AND U9536 ( .A(n1218), .B(n9863), .Z(n9862) );
  XOR U9537 ( .A(n9864), .B(n9865), .Z(n9856) );
  AND U9538 ( .A(n1222), .B(n9855), .Z(n9865) );
  XNOR U9539 ( .A(n9866), .B(n9853), .Z(n9855) );
  XOR U9540 ( .A(n9867), .B(n9868), .Z(n9853) );
  AND U9541 ( .A(n1245), .B(n9869), .Z(n9868) );
  IV U9542 ( .A(n9864), .Z(n9866) );
  XOR U9543 ( .A(n9870), .B(n9871), .Z(n9864) );
  AND U9544 ( .A(n1229), .B(n9863), .Z(n9871) );
  XNOR U9545 ( .A(n9861), .B(n9870), .Z(n9863) );
  XNOR U9546 ( .A(n9872), .B(n9873), .Z(n9861) );
  AND U9547 ( .A(n1233), .B(n9874), .Z(n9873) );
  XOR U9548 ( .A(p_input[1885]), .B(n9872), .Z(n9874) );
  XNOR U9549 ( .A(n9875), .B(n9876), .Z(n9872) );
  AND U9550 ( .A(n1237), .B(n9877), .Z(n9876) );
  XOR U9551 ( .A(n9878), .B(n9879), .Z(n9870) );
  AND U9552 ( .A(n1241), .B(n9869), .Z(n9879) );
  XNOR U9553 ( .A(n9880), .B(n9867), .Z(n9869) );
  XOR U9554 ( .A(n9881), .B(n9882), .Z(n9867) );
  AND U9555 ( .A(n1264), .B(n9883), .Z(n9882) );
  IV U9556 ( .A(n9878), .Z(n9880) );
  XOR U9557 ( .A(n9884), .B(n9885), .Z(n9878) );
  AND U9558 ( .A(n1248), .B(n9877), .Z(n9885) );
  XNOR U9559 ( .A(n9875), .B(n9884), .Z(n9877) );
  XNOR U9560 ( .A(n9886), .B(n9887), .Z(n9875) );
  AND U9561 ( .A(n1252), .B(n9888), .Z(n9887) );
  XOR U9562 ( .A(p_input[1917]), .B(n9886), .Z(n9888) );
  XNOR U9563 ( .A(n9889), .B(n9890), .Z(n9886) );
  AND U9564 ( .A(n1256), .B(n9891), .Z(n9890) );
  XOR U9565 ( .A(n9892), .B(n9893), .Z(n9884) );
  AND U9566 ( .A(n1260), .B(n9883), .Z(n9893) );
  XNOR U9567 ( .A(n9894), .B(n9881), .Z(n9883) );
  XOR U9568 ( .A(n9895), .B(n9896), .Z(n9881) );
  AND U9569 ( .A(n1282), .B(n9897), .Z(n9896) );
  IV U9570 ( .A(n9892), .Z(n9894) );
  XOR U9571 ( .A(n9898), .B(n9899), .Z(n9892) );
  AND U9572 ( .A(n1267), .B(n9891), .Z(n9899) );
  XNOR U9573 ( .A(n9889), .B(n9898), .Z(n9891) );
  XNOR U9574 ( .A(n9900), .B(n9901), .Z(n9889) );
  AND U9575 ( .A(n1271), .B(n9902), .Z(n9901) );
  XOR U9576 ( .A(p_input[1949]), .B(n9900), .Z(n9902) );
  XOR U9577 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][29] ), .B(n9903), 
        .Z(n9900) );
  AND U9578 ( .A(n1274), .B(n9904), .Z(n9903) );
  XOR U9579 ( .A(n9905), .B(n9906), .Z(n9898) );
  AND U9580 ( .A(n1278), .B(n9897), .Z(n9906) );
  XNOR U9581 ( .A(n9907), .B(n9895), .Z(n9897) );
  XOR U9582 ( .A(\knn_comb_/min_val_out[0][29] ), .B(n9908), .Z(n9895) );
  AND U9583 ( .A(n1290), .B(n9909), .Z(n9908) );
  IV U9584 ( .A(n9905), .Z(n9907) );
  XOR U9585 ( .A(n9910), .B(n9911), .Z(n9905) );
  AND U9586 ( .A(n1285), .B(n9904), .Z(n9911) );
  XOR U9587 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][29] ), .B(n9910), 
        .Z(n9904) );
  XOR U9588 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .B(n9912), 
        .Z(n9910) );
  AND U9589 ( .A(n1287), .B(n9909), .Z(n9912) );
  XOR U9590 ( .A(\knn_comb_/min_val_out[0][29] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .Z(n9909) );
  XOR U9591 ( .A(n79), .B(n9913), .Z(o[28]) );
  AND U9592 ( .A(n122), .B(n9914), .Z(n79) );
  XOR U9593 ( .A(n80), .B(n9913), .Z(n9914) );
  XOR U9594 ( .A(n9915), .B(n9916), .Z(n9913) );
  AND U9595 ( .A(n142), .B(n9917), .Z(n9916) );
  XOR U9596 ( .A(n9918), .B(n9), .Z(n80) );
  AND U9597 ( .A(n125), .B(n9919), .Z(n9) );
  XOR U9598 ( .A(n10), .B(n9918), .Z(n9919) );
  XOR U9599 ( .A(n9920), .B(n9921), .Z(n10) );
  AND U9600 ( .A(n130), .B(n9922), .Z(n9921) );
  XOR U9601 ( .A(p_input[28]), .B(n9920), .Z(n9922) );
  XNOR U9602 ( .A(n9923), .B(n9924), .Z(n9920) );
  AND U9603 ( .A(n134), .B(n9925), .Z(n9924) );
  XOR U9604 ( .A(n9926), .B(n9927), .Z(n9918) );
  AND U9605 ( .A(n138), .B(n9917), .Z(n9927) );
  XNOR U9606 ( .A(n9928), .B(n9915), .Z(n9917) );
  XOR U9607 ( .A(n9929), .B(n9930), .Z(n9915) );
  AND U9608 ( .A(n162), .B(n9931), .Z(n9930) );
  IV U9609 ( .A(n9926), .Z(n9928) );
  XOR U9610 ( .A(n9932), .B(n9933), .Z(n9926) );
  AND U9611 ( .A(n146), .B(n9925), .Z(n9933) );
  XNOR U9612 ( .A(n9923), .B(n9932), .Z(n9925) );
  XNOR U9613 ( .A(n9934), .B(n9935), .Z(n9923) );
  AND U9614 ( .A(n150), .B(n9936), .Z(n9935) );
  XOR U9615 ( .A(p_input[60]), .B(n9934), .Z(n9936) );
  XNOR U9616 ( .A(n9937), .B(n9938), .Z(n9934) );
  AND U9617 ( .A(n154), .B(n9939), .Z(n9938) );
  XOR U9618 ( .A(n9940), .B(n9941), .Z(n9932) );
  AND U9619 ( .A(n158), .B(n9931), .Z(n9941) );
  XNOR U9620 ( .A(n9942), .B(n9929), .Z(n9931) );
  XOR U9621 ( .A(n9943), .B(n9944), .Z(n9929) );
  AND U9622 ( .A(n181), .B(n9945), .Z(n9944) );
  IV U9623 ( .A(n9940), .Z(n9942) );
  XOR U9624 ( .A(n9946), .B(n9947), .Z(n9940) );
  AND U9625 ( .A(n165), .B(n9939), .Z(n9947) );
  XNOR U9626 ( .A(n9937), .B(n9946), .Z(n9939) );
  XNOR U9627 ( .A(n9948), .B(n9949), .Z(n9937) );
  AND U9628 ( .A(n169), .B(n9950), .Z(n9949) );
  XOR U9629 ( .A(p_input[92]), .B(n9948), .Z(n9950) );
  XNOR U9630 ( .A(n9951), .B(n9952), .Z(n9948) );
  AND U9631 ( .A(n173), .B(n9953), .Z(n9952) );
  XOR U9632 ( .A(n9954), .B(n9955), .Z(n9946) );
  AND U9633 ( .A(n177), .B(n9945), .Z(n9955) );
  XNOR U9634 ( .A(n9956), .B(n9943), .Z(n9945) );
  XOR U9635 ( .A(n9957), .B(n9958), .Z(n9943) );
  AND U9636 ( .A(n200), .B(n9959), .Z(n9958) );
  IV U9637 ( .A(n9954), .Z(n9956) );
  XOR U9638 ( .A(n9960), .B(n9961), .Z(n9954) );
  AND U9639 ( .A(n184), .B(n9953), .Z(n9961) );
  XNOR U9640 ( .A(n9951), .B(n9960), .Z(n9953) );
  XNOR U9641 ( .A(n9962), .B(n9963), .Z(n9951) );
  AND U9642 ( .A(n188), .B(n9964), .Z(n9963) );
  XOR U9643 ( .A(p_input[124]), .B(n9962), .Z(n9964) );
  XNOR U9644 ( .A(n9965), .B(n9966), .Z(n9962) );
  AND U9645 ( .A(n192), .B(n9967), .Z(n9966) );
  XOR U9646 ( .A(n9968), .B(n9969), .Z(n9960) );
  AND U9647 ( .A(n196), .B(n9959), .Z(n9969) );
  XNOR U9648 ( .A(n9970), .B(n9957), .Z(n9959) );
  XOR U9649 ( .A(n9971), .B(n9972), .Z(n9957) );
  AND U9650 ( .A(n219), .B(n9973), .Z(n9972) );
  IV U9651 ( .A(n9968), .Z(n9970) );
  XOR U9652 ( .A(n9974), .B(n9975), .Z(n9968) );
  AND U9653 ( .A(n203), .B(n9967), .Z(n9975) );
  XNOR U9654 ( .A(n9965), .B(n9974), .Z(n9967) );
  XNOR U9655 ( .A(n9976), .B(n9977), .Z(n9965) );
  AND U9656 ( .A(n207), .B(n9978), .Z(n9977) );
  XOR U9657 ( .A(p_input[156]), .B(n9976), .Z(n9978) );
  XNOR U9658 ( .A(n9979), .B(n9980), .Z(n9976) );
  AND U9659 ( .A(n211), .B(n9981), .Z(n9980) );
  XOR U9660 ( .A(n9982), .B(n9983), .Z(n9974) );
  AND U9661 ( .A(n215), .B(n9973), .Z(n9983) );
  XNOR U9662 ( .A(n9984), .B(n9971), .Z(n9973) );
  XOR U9663 ( .A(n9985), .B(n9986), .Z(n9971) );
  AND U9664 ( .A(n238), .B(n9987), .Z(n9986) );
  IV U9665 ( .A(n9982), .Z(n9984) );
  XOR U9666 ( .A(n9988), .B(n9989), .Z(n9982) );
  AND U9667 ( .A(n222), .B(n9981), .Z(n9989) );
  XNOR U9668 ( .A(n9979), .B(n9988), .Z(n9981) );
  XNOR U9669 ( .A(n9990), .B(n9991), .Z(n9979) );
  AND U9670 ( .A(n226), .B(n9992), .Z(n9991) );
  XOR U9671 ( .A(p_input[188]), .B(n9990), .Z(n9992) );
  XNOR U9672 ( .A(n9993), .B(n9994), .Z(n9990) );
  AND U9673 ( .A(n230), .B(n9995), .Z(n9994) );
  XOR U9674 ( .A(n9996), .B(n9997), .Z(n9988) );
  AND U9675 ( .A(n234), .B(n9987), .Z(n9997) );
  XNOR U9676 ( .A(n9998), .B(n9985), .Z(n9987) );
  XOR U9677 ( .A(n9999), .B(n10000), .Z(n9985) );
  AND U9678 ( .A(n257), .B(n10001), .Z(n10000) );
  IV U9679 ( .A(n9996), .Z(n9998) );
  XOR U9680 ( .A(n10002), .B(n10003), .Z(n9996) );
  AND U9681 ( .A(n241), .B(n9995), .Z(n10003) );
  XNOR U9682 ( .A(n9993), .B(n10002), .Z(n9995) );
  XNOR U9683 ( .A(n10004), .B(n10005), .Z(n9993) );
  AND U9684 ( .A(n245), .B(n10006), .Z(n10005) );
  XOR U9685 ( .A(p_input[220]), .B(n10004), .Z(n10006) );
  XNOR U9686 ( .A(n10007), .B(n10008), .Z(n10004) );
  AND U9687 ( .A(n249), .B(n10009), .Z(n10008) );
  XOR U9688 ( .A(n10010), .B(n10011), .Z(n10002) );
  AND U9689 ( .A(n253), .B(n10001), .Z(n10011) );
  XNOR U9690 ( .A(n10012), .B(n9999), .Z(n10001) );
  XOR U9691 ( .A(n10013), .B(n10014), .Z(n9999) );
  AND U9692 ( .A(n276), .B(n10015), .Z(n10014) );
  IV U9693 ( .A(n10010), .Z(n10012) );
  XOR U9694 ( .A(n10016), .B(n10017), .Z(n10010) );
  AND U9695 ( .A(n260), .B(n10009), .Z(n10017) );
  XNOR U9696 ( .A(n10007), .B(n10016), .Z(n10009) );
  XNOR U9697 ( .A(n10018), .B(n10019), .Z(n10007) );
  AND U9698 ( .A(n264), .B(n10020), .Z(n10019) );
  XOR U9699 ( .A(p_input[252]), .B(n10018), .Z(n10020) );
  XNOR U9700 ( .A(n10021), .B(n10022), .Z(n10018) );
  AND U9701 ( .A(n268), .B(n10023), .Z(n10022) );
  XOR U9702 ( .A(n10024), .B(n10025), .Z(n10016) );
  AND U9703 ( .A(n272), .B(n10015), .Z(n10025) );
  XNOR U9704 ( .A(n10026), .B(n10013), .Z(n10015) );
  XOR U9705 ( .A(n10027), .B(n10028), .Z(n10013) );
  AND U9706 ( .A(n295), .B(n10029), .Z(n10028) );
  IV U9707 ( .A(n10024), .Z(n10026) );
  XOR U9708 ( .A(n10030), .B(n10031), .Z(n10024) );
  AND U9709 ( .A(n279), .B(n10023), .Z(n10031) );
  XNOR U9710 ( .A(n10021), .B(n10030), .Z(n10023) );
  XNOR U9711 ( .A(n10032), .B(n10033), .Z(n10021) );
  AND U9712 ( .A(n283), .B(n10034), .Z(n10033) );
  XOR U9713 ( .A(p_input[284]), .B(n10032), .Z(n10034) );
  XNOR U9714 ( .A(n10035), .B(n10036), .Z(n10032) );
  AND U9715 ( .A(n287), .B(n10037), .Z(n10036) );
  XOR U9716 ( .A(n10038), .B(n10039), .Z(n10030) );
  AND U9717 ( .A(n291), .B(n10029), .Z(n10039) );
  XNOR U9718 ( .A(n10040), .B(n10027), .Z(n10029) );
  XOR U9719 ( .A(n10041), .B(n10042), .Z(n10027) );
  AND U9720 ( .A(n314), .B(n10043), .Z(n10042) );
  IV U9721 ( .A(n10038), .Z(n10040) );
  XOR U9722 ( .A(n10044), .B(n10045), .Z(n10038) );
  AND U9723 ( .A(n298), .B(n10037), .Z(n10045) );
  XNOR U9724 ( .A(n10035), .B(n10044), .Z(n10037) );
  XNOR U9725 ( .A(n10046), .B(n10047), .Z(n10035) );
  AND U9726 ( .A(n302), .B(n10048), .Z(n10047) );
  XOR U9727 ( .A(p_input[316]), .B(n10046), .Z(n10048) );
  XNOR U9728 ( .A(n10049), .B(n10050), .Z(n10046) );
  AND U9729 ( .A(n306), .B(n10051), .Z(n10050) );
  XOR U9730 ( .A(n10052), .B(n10053), .Z(n10044) );
  AND U9731 ( .A(n310), .B(n10043), .Z(n10053) );
  XNOR U9732 ( .A(n10054), .B(n10041), .Z(n10043) );
  XOR U9733 ( .A(n10055), .B(n10056), .Z(n10041) );
  AND U9734 ( .A(n333), .B(n10057), .Z(n10056) );
  IV U9735 ( .A(n10052), .Z(n10054) );
  XOR U9736 ( .A(n10058), .B(n10059), .Z(n10052) );
  AND U9737 ( .A(n317), .B(n10051), .Z(n10059) );
  XNOR U9738 ( .A(n10049), .B(n10058), .Z(n10051) );
  XNOR U9739 ( .A(n10060), .B(n10061), .Z(n10049) );
  AND U9740 ( .A(n321), .B(n10062), .Z(n10061) );
  XOR U9741 ( .A(p_input[348]), .B(n10060), .Z(n10062) );
  XNOR U9742 ( .A(n10063), .B(n10064), .Z(n10060) );
  AND U9743 ( .A(n325), .B(n10065), .Z(n10064) );
  XOR U9744 ( .A(n10066), .B(n10067), .Z(n10058) );
  AND U9745 ( .A(n329), .B(n10057), .Z(n10067) );
  XNOR U9746 ( .A(n10068), .B(n10055), .Z(n10057) );
  XOR U9747 ( .A(n10069), .B(n10070), .Z(n10055) );
  AND U9748 ( .A(n352), .B(n10071), .Z(n10070) );
  IV U9749 ( .A(n10066), .Z(n10068) );
  XOR U9750 ( .A(n10072), .B(n10073), .Z(n10066) );
  AND U9751 ( .A(n336), .B(n10065), .Z(n10073) );
  XNOR U9752 ( .A(n10063), .B(n10072), .Z(n10065) );
  XNOR U9753 ( .A(n10074), .B(n10075), .Z(n10063) );
  AND U9754 ( .A(n340), .B(n10076), .Z(n10075) );
  XOR U9755 ( .A(p_input[380]), .B(n10074), .Z(n10076) );
  XNOR U9756 ( .A(n10077), .B(n10078), .Z(n10074) );
  AND U9757 ( .A(n344), .B(n10079), .Z(n10078) );
  XOR U9758 ( .A(n10080), .B(n10081), .Z(n10072) );
  AND U9759 ( .A(n348), .B(n10071), .Z(n10081) );
  XNOR U9760 ( .A(n10082), .B(n10069), .Z(n10071) );
  XOR U9761 ( .A(n10083), .B(n10084), .Z(n10069) );
  AND U9762 ( .A(n371), .B(n10085), .Z(n10084) );
  IV U9763 ( .A(n10080), .Z(n10082) );
  XOR U9764 ( .A(n10086), .B(n10087), .Z(n10080) );
  AND U9765 ( .A(n355), .B(n10079), .Z(n10087) );
  XNOR U9766 ( .A(n10077), .B(n10086), .Z(n10079) );
  XNOR U9767 ( .A(n10088), .B(n10089), .Z(n10077) );
  AND U9768 ( .A(n359), .B(n10090), .Z(n10089) );
  XOR U9769 ( .A(p_input[412]), .B(n10088), .Z(n10090) );
  XNOR U9770 ( .A(n10091), .B(n10092), .Z(n10088) );
  AND U9771 ( .A(n363), .B(n10093), .Z(n10092) );
  XOR U9772 ( .A(n10094), .B(n10095), .Z(n10086) );
  AND U9773 ( .A(n367), .B(n10085), .Z(n10095) );
  XNOR U9774 ( .A(n10096), .B(n10083), .Z(n10085) );
  XOR U9775 ( .A(n10097), .B(n10098), .Z(n10083) );
  AND U9776 ( .A(n390), .B(n10099), .Z(n10098) );
  IV U9777 ( .A(n10094), .Z(n10096) );
  XOR U9778 ( .A(n10100), .B(n10101), .Z(n10094) );
  AND U9779 ( .A(n374), .B(n10093), .Z(n10101) );
  XNOR U9780 ( .A(n10091), .B(n10100), .Z(n10093) );
  XNOR U9781 ( .A(n10102), .B(n10103), .Z(n10091) );
  AND U9782 ( .A(n378), .B(n10104), .Z(n10103) );
  XOR U9783 ( .A(p_input[444]), .B(n10102), .Z(n10104) );
  XNOR U9784 ( .A(n10105), .B(n10106), .Z(n10102) );
  AND U9785 ( .A(n382), .B(n10107), .Z(n10106) );
  XOR U9786 ( .A(n10108), .B(n10109), .Z(n10100) );
  AND U9787 ( .A(n386), .B(n10099), .Z(n10109) );
  XNOR U9788 ( .A(n10110), .B(n10097), .Z(n10099) );
  XOR U9789 ( .A(n10111), .B(n10112), .Z(n10097) );
  AND U9790 ( .A(n409), .B(n10113), .Z(n10112) );
  IV U9791 ( .A(n10108), .Z(n10110) );
  XOR U9792 ( .A(n10114), .B(n10115), .Z(n10108) );
  AND U9793 ( .A(n393), .B(n10107), .Z(n10115) );
  XNOR U9794 ( .A(n10105), .B(n10114), .Z(n10107) );
  XNOR U9795 ( .A(n10116), .B(n10117), .Z(n10105) );
  AND U9796 ( .A(n397), .B(n10118), .Z(n10117) );
  XOR U9797 ( .A(p_input[476]), .B(n10116), .Z(n10118) );
  XNOR U9798 ( .A(n10119), .B(n10120), .Z(n10116) );
  AND U9799 ( .A(n401), .B(n10121), .Z(n10120) );
  XOR U9800 ( .A(n10122), .B(n10123), .Z(n10114) );
  AND U9801 ( .A(n405), .B(n10113), .Z(n10123) );
  XNOR U9802 ( .A(n10124), .B(n10111), .Z(n10113) );
  XOR U9803 ( .A(n10125), .B(n10126), .Z(n10111) );
  AND U9804 ( .A(n428), .B(n10127), .Z(n10126) );
  IV U9805 ( .A(n10122), .Z(n10124) );
  XOR U9806 ( .A(n10128), .B(n10129), .Z(n10122) );
  AND U9807 ( .A(n412), .B(n10121), .Z(n10129) );
  XNOR U9808 ( .A(n10119), .B(n10128), .Z(n10121) );
  XNOR U9809 ( .A(n10130), .B(n10131), .Z(n10119) );
  AND U9810 ( .A(n416), .B(n10132), .Z(n10131) );
  XOR U9811 ( .A(p_input[508]), .B(n10130), .Z(n10132) );
  XNOR U9812 ( .A(n10133), .B(n10134), .Z(n10130) );
  AND U9813 ( .A(n420), .B(n10135), .Z(n10134) );
  XOR U9814 ( .A(n10136), .B(n10137), .Z(n10128) );
  AND U9815 ( .A(n424), .B(n10127), .Z(n10137) );
  XNOR U9816 ( .A(n10138), .B(n10125), .Z(n10127) );
  XOR U9817 ( .A(n10139), .B(n10140), .Z(n10125) );
  AND U9818 ( .A(n447), .B(n10141), .Z(n10140) );
  IV U9819 ( .A(n10136), .Z(n10138) );
  XOR U9820 ( .A(n10142), .B(n10143), .Z(n10136) );
  AND U9821 ( .A(n431), .B(n10135), .Z(n10143) );
  XNOR U9822 ( .A(n10133), .B(n10142), .Z(n10135) );
  XNOR U9823 ( .A(n10144), .B(n10145), .Z(n10133) );
  AND U9824 ( .A(n435), .B(n10146), .Z(n10145) );
  XOR U9825 ( .A(p_input[540]), .B(n10144), .Z(n10146) );
  XNOR U9826 ( .A(n10147), .B(n10148), .Z(n10144) );
  AND U9827 ( .A(n439), .B(n10149), .Z(n10148) );
  XOR U9828 ( .A(n10150), .B(n10151), .Z(n10142) );
  AND U9829 ( .A(n443), .B(n10141), .Z(n10151) );
  XNOR U9830 ( .A(n10152), .B(n10139), .Z(n10141) );
  XOR U9831 ( .A(n10153), .B(n10154), .Z(n10139) );
  AND U9832 ( .A(n466), .B(n10155), .Z(n10154) );
  IV U9833 ( .A(n10150), .Z(n10152) );
  XOR U9834 ( .A(n10156), .B(n10157), .Z(n10150) );
  AND U9835 ( .A(n450), .B(n10149), .Z(n10157) );
  XNOR U9836 ( .A(n10147), .B(n10156), .Z(n10149) );
  XNOR U9837 ( .A(n10158), .B(n10159), .Z(n10147) );
  AND U9838 ( .A(n454), .B(n10160), .Z(n10159) );
  XOR U9839 ( .A(p_input[572]), .B(n10158), .Z(n10160) );
  XNOR U9840 ( .A(n10161), .B(n10162), .Z(n10158) );
  AND U9841 ( .A(n458), .B(n10163), .Z(n10162) );
  XOR U9842 ( .A(n10164), .B(n10165), .Z(n10156) );
  AND U9843 ( .A(n462), .B(n10155), .Z(n10165) );
  XNOR U9844 ( .A(n10166), .B(n10153), .Z(n10155) );
  XOR U9845 ( .A(n10167), .B(n10168), .Z(n10153) );
  AND U9846 ( .A(n485), .B(n10169), .Z(n10168) );
  IV U9847 ( .A(n10164), .Z(n10166) );
  XOR U9848 ( .A(n10170), .B(n10171), .Z(n10164) );
  AND U9849 ( .A(n469), .B(n10163), .Z(n10171) );
  XNOR U9850 ( .A(n10161), .B(n10170), .Z(n10163) );
  XNOR U9851 ( .A(n10172), .B(n10173), .Z(n10161) );
  AND U9852 ( .A(n473), .B(n10174), .Z(n10173) );
  XOR U9853 ( .A(p_input[604]), .B(n10172), .Z(n10174) );
  XNOR U9854 ( .A(n10175), .B(n10176), .Z(n10172) );
  AND U9855 ( .A(n477), .B(n10177), .Z(n10176) );
  XOR U9856 ( .A(n10178), .B(n10179), .Z(n10170) );
  AND U9857 ( .A(n481), .B(n10169), .Z(n10179) );
  XNOR U9858 ( .A(n10180), .B(n10167), .Z(n10169) );
  XOR U9859 ( .A(n10181), .B(n10182), .Z(n10167) );
  AND U9860 ( .A(n504), .B(n10183), .Z(n10182) );
  IV U9861 ( .A(n10178), .Z(n10180) );
  XOR U9862 ( .A(n10184), .B(n10185), .Z(n10178) );
  AND U9863 ( .A(n488), .B(n10177), .Z(n10185) );
  XNOR U9864 ( .A(n10175), .B(n10184), .Z(n10177) );
  XNOR U9865 ( .A(n10186), .B(n10187), .Z(n10175) );
  AND U9866 ( .A(n492), .B(n10188), .Z(n10187) );
  XOR U9867 ( .A(p_input[636]), .B(n10186), .Z(n10188) );
  XNOR U9868 ( .A(n10189), .B(n10190), .Z(n10186) );
  AND U9869 ( .A(n496), .B(n10191), .Z(n10190) );
  XOR U9870 ( .A(n10192), .B(n10193), .Z(n10184) );
  AND U9871 ( .A(n500), .B(n10183), .Z(n10193) );
  XNOR U9872 ( .A(n10194), .B(n10181), .Z(n10183) );
  XOR U9873 ( .A(n10195), .B(n10196), .Z(n10181) );
  AND U9874 ( .A(n523), .B(n10197), .Z(n10196) );
  IV U9875 ( .A(n10192), .Z(n10194) );
  XOR U9876 ( .A(n10198), .B(n10199), .Z(n10192) );
  AND U9877 ( .A(n507), .B(n10191), .Z(n10199) );
  XNOR U9878 ( .A(n10189), .B(n10198), .Z(n10191) );
  XNOR U9879 ( .A(n10200), .B(n10201), .Z(n10189) );
  AND U9880 ( .A(n511), .B(n10202), .Z(n10201) );
  XOR U9881 ( .A(p_input[668]), .B(n10200), .Z(n10202) );
  XNOR U9882 ( .A(n10203), .B(n10204), .Z(n10200) );
  AND U9883 ( .A(n515), .B(n10205), .Z(n10204) );
  XOR U9884 ( .A(n10206), .B(n10207), .Z(n10198) );
  AND U9885 ( .A(n519), .B(n10197), .Z(n10207) );
  XNOR U9886 ( .A(n10208), .B(n10195), .Z(n10197) );
  XOR U9887 ( .A(n10209), .B(n10210), .Z(n10195) );
  AND U9888 ( .A(n542), .B(n10211), .Z(n10210) );
  IV U9889 ( .A(n10206), .Z(n10208) );
  XOR U9890 ( .A(n10212), .B(n10213), .Z(n10206) );
  AND U9891 ( .A(n526), .B(n10205), .Z(n10213) );
  XNOR U9892 ( .A(n10203), .B(n10212), .Z(n10205) );
  XNOR U9893 ( .A(n10214), .B(n10215), .Z(n10203) );
  AND U9894 ( .A(n530), .B(n10216), .Z(n10215) );
  XOR U9895 ( .A(p_input[700]), .B(n10214), .Z(n10216) );
  XNOR U9896 ( .A(n10217), .B(n10218), .Z(n10214) );
  AND U9897 ( .A(n534), .B(n10219), .Z(n10218) );
  XOR U9898 ( .A(n10220), .B(n10221), .Z(n10212) );
  AND U9899 ( .A(n538), .B(n10211), .Z(n10221) );
  XNOR U9900 ( .A(n10222), .B(n10209), .Z(n10211) );
  XOR U9901 ( .A(n10223), .B(n10224), .Z(n10209) );
  AND U9902 ( .A(n561), .B(n10225), .Z(n10224) );
  IV U9903 ( .A(n10220), .Z(n10222) );
  XOR U9904 ( .A(n10226), .B(n10227), .Z(n10220) );
  AND U9905 ( .A(n545), .B(n10219), .Z(n10227) );
  XNOR U9906 ( .A(n10217), .B(n10226), .Z(n10219) );
  XNOR U9907 ( .A(n10228), .B(n10229), .Z(n10217) );
  AND U9908 ( .A(n549), .B(n10230), .Z(n10229) );
  XOR U9909 ( .A(p_input[732]), .B(n10228), .Z(n10230) );
  XNOR U9910 ( .A(n10231), .B(n10232), .Z(n10228) );
  AND U9911 ( .A(n553), .B(n10233), .Z(n10232) );
  XOR U9912 ( .A(n10234), .B(n10235), .Z(n10226) );
  AND U9913 ( .A(n557), .B(n10225), .Z(n10235) );
  XNOR U9914 ( .A(n10236), .B(n10223), .Z(n10225) );
  XOR U9915 ( .A(n10237), .B(n10238), .Z(n10223) );
  AND U9916 ( .A(n580), .B(n10239), .Z(n10238) );
  IV U9917 ( .A(n10234), .Z(n10236) );
  XOR U9918 ( .A(n10240), .B(n10241), .Z(n10234) );
  AND U9919 ( .A(n564), .B(n10233), .Z(n10241) );
  XNOR U9920 ( .A(n10231), .B(n10240), .Z(n10233) );
  XNOR U9921 ( .A(n10242), .B(n10243), .Z(n10231) );
  AND U9922 ( .A(n568), .B(n10244), .Z(n10243) );
  XOR U9923 ( .A(p_input[764]), .B(n10242), .Z(n10244) );
  XNOR U9924 ( .A(n10245), .B(n10246), .Z(n10242) );
  AND U9925 ( .A(n572), .B(n10247), .Z(n10246) );
  XOR U9926 ( .A(n10248), .B(n10249), .Z(n10240) );
  AND U9927 ( .A(n576), .B(n10239), .Z(n10249) );
  XNOR U9928 ( .A(n10250), .B(n10237), .Z(n10239) );
  XOR U9929 ( .A(n10251), .B(n10252), .Z(n10237) );
  AND U9930 ( .A(n599), .B(n10253), .Z(n10252) );
  IV U9931 ( .A(n10248), .Z(n10250) );
  XOR U9932 ( .A(n10254), .B(n10255), .Z(n10248) );
  AND U9933 ( .A(n583), .B(n10247), .Z(n10255) );
  XNOR U9934 ( .A(n10245), .B(n10254), .Z(n10247) );
  XNOR U9935 ( .A(n10256), .B(n10257), .Z(n10245) );
  AND U9936 ( .A(n587), .B(n10258), .Z(n10257) );
  XOR U9937 ( .A(p_input[796]), .B(n10256), .Z(n10258) );
  XNOR U9938 ( .A(n10259), .B(n10260), .Z(n10256) );
  AND U9939 ( .A(n591), .B(n10261), .Z(n10260) );
  XOR U9940 ( .A(n10262), .B(n10263), .Z(n10254) );
  AND U9941 ( .A(n595), .B(n10253), .Z(n10263) );
  XNOR U9942 ( .A(n10264), .B(n10251), .Z(n10253) );
  XOR U9943 ( .A(n10265), .B(n10266), .Z(n10251) );
  AND U9944 ( .A(n618), .B(n10267), .Z(n10266) );
  IV U9945 ( .A(n10262), .Z(n10264) );
  XOR U9946 ( .A(n10268), .B(n10269), .Z(n10262) );
  AND U9947 ( .A(n602), .B(n10261), .Z(n10269) );
  XNOR U9948 ( .A(n10259), .B(n10268), .Z(n10261) );
  XNOR U9949 ( .A(n10270), .B(n10271), .Z(n10259) );
  AND U9950 ( .A(n606), .B(n10272), .Z(n10271) );
  XOR U9951 ( .A(p_input[828]), .B(n10270), .Z(n10272) );
  XNOR U9952 ( .A(n10273), .B(n10274), .Z(n10270) );
  AND U9953 ( .A(n610), .B(n10275), .Z(n10274) );
  XOR U9954 ( .A(n10276), .B(n10277), .Z(n10268) );
  AND U9955 ( .A(n614), .B(n10267), .Z(n10277) );
  XNOR U9956 ( .A(n10278), .B(n10265), .Z(n10267) );
  XOR U9957 ( .A(n10279), .B(n10280), .Z(n10265) );
  AND U9958 ( .A(n637), .B(n10281), .Z(n10280) );
  IV U9959 ( .A(n10276), .Z(n10278) );
  XOR U9960 ( .A(n10282), .B(n10283), .Z(n10276) );
  AND U9961 ( .A(n621), .B(n10275), .Z(n10283) );
  XNOR U9962 ( .A(n10273), .B(n10282), .Z(n10275) );
  XNOR U9963 ( .A(n10284), .B(n10285), .Z(n10273) );
  AND U9964 ( .A(n625), .B(n10286), .Z(n10285) );
  XOR U9965 ( .A(p_input[860]), .B(n10284), .Z(n10286) );
  XNOR U9966 ( .A(n10287), .B(n10288), .Z(n10284) );
  AND U9967 ( .A(n629), .B(n10289), .Z(n10288) );
  XOR U9968 ( .A(n10290), .B(n10291), .Z(n10282) );
  AND U9969 ( .A(n633), .B(n10281), .Z(n10291) );
  XNOR U9970 ( .A(n10292), .B(n10279), .Z(n10281) );
  XOR U9971 ( .A(n10293), .B(n10294), .Z(n10279) );
  AND U9972 ( .A(n656), .B(n10295), .Z(n10294) );
  IV U9973 ( .A(n10290), .Z(n10292) );
  XOR U9974 ( .A(n10296), .B(n10297), .Z(n10290) );
  AND U9975 ( .A(n640), .B(n10289), .Z(n10297) );
  XNOR U9976 ( .A(n10287), .B(n10296), .Z(n10289) );
  XNOR U9977 ( .A(n10298), .B(n10299), .Z(n10287) );
  AND U9978 ( .A(n644), .B(n10300), .Z(n10299) );
  XOR U9979 ( .A(p_input[892]), .B(n10298), .Z(n10300) );
  XNOR U9980 ( .A(n10301), .B(n10302), .Z(n10298) );
  AND U9981 ( .A(n648), .B(n10303), .Z(n10302) );
  XOR U9982 ( .A(n10304), .B(n10305), .Z(n10296) );
  AND U9983 ( .A(n652), .B(n10295), .Z(n10305) );
  XNOR U9984 ( .A(n10306), .B(n10293), .Z(n10295) );
  XOR U9985 ( .A(n10307), .B(n10308), .Z(n10293) );
  AND U9986 ( .A(n675), .B(n10309), .Z(n10308) );
  IV U9987 ( .A(n10304), .Z(n10306) );
  XOR U9988 ( .A(n10310), .B(n10311), .Z(n10304) );
  AND U9989 ( .A(n659), .B(n10303), .Z(n10311) );
  XNOR U9990 ( .A(n10301), .B(n10310), .Z(n10303) );
  XNOR U9991 ( .A(n10312), .B(n10313), .Z(n10301) );
  AND U9992 ( .A(n663), .B(n10314), .Z(n10313) );
  XOR U9993 ( .A(p_input[924]), .B(n10312), .Z(n10314) );
  XNOR U9994 ( .A(n10315), .B(n10316), .Z(n10312) );
  AND U9995 ( .A(n667), .B(n10317), .Z(n10316) );
  XOR U9996 ( .A(n10318), .B(n10319), .Z(n10310) );
  AND U9997 ( .A(n671), .B(n10309), .Z(n10319) );
  XNOR U9998 ( .A(n10320), .B(n10307), .Z(n10309) );
  XOR U9999 ( .A(n10321), .B(n10322), .Z(n10307) );
  AND U10000 ( .A(n694), .B(n10323), .Z(n10322) );
  IV U10001 ( .A(n10318), .Z(n10320) );
  XOR U10002 ( .A(n10324), .B(n10325), .Z(n10318) );
  AND U10003 ( .A(n678), .B(n10317), .Z(n10325) );
  XNOR U10004 ( .A(n10315), .B(n10324), .Z(n10317) );
  XNOR U10005 ( .A(n10326), .B(n10327), .Z(n10315) );
  AND U10006 ( .A(n682), .B(n10328), .Z(n10327) );
  XOR U10007 ( .A(p_input[956]), .B(n10326), .Z(n10328) );
  XNOR U10008 ( .A(n10329), .B(n10330), .Z(n10326) );
  AND U10009 ( .A(n686), .B(n10331), .Z(n10330) );
  XOR U10010 ( .A(n10332), .B(n10333), .Z(n10324) );
  AND U10011 ( .A(n690), .B(n10323), .Z(n10333) );
  XNOR U10012 ( .A(n10334), .B(n10321), .Z(n10323) );
  XOR U10013 ( .A(n10335), .B(n10336), .Z(n10321) );
  AND U10014 ( .A(n713), .B(n10337), .Z(n10336) );
  IV U10015 ( .A(n10332), .Z(n10334) );
  XOR U10016 ( .A(n10338), .B(n10339), .Z(n10332) );
  AND U10017 ( .A(n697), .B(n10331), .Z(n10339) );
  XNOR U10018 ( .A(n10329), .B(n10338), .Z(n10331) );
  XNOR U10019 ( .A(n10340), .B(n10341), .Z(n10329) );
  AND U10020 ( .A(n701), .B(n10342), .Z(n10341) );
  XOR U10021 ( .A(p_input[988]), .B(n10340), .Z(n10342) );
  XNOR U10022 ( .A(n10343), .B(n10344), .Z(n10340) );
  AND U10023 ( .A(n705), .B(n10345), .Z(n10344) );
  XOR U10024 ( .A(n10346), .B(n10347), .Z(n10338) );
  AND U10025 ( .A(n709), .B(n10337), .Z(n10347) );
  XNOR U10026 ( .A(n10348), .B(n10335), .Z(n10337) );
  XOR U10027 ( .A(n10349), .B(n10350), .Z(n10335) );
  AND U10028 ( .A(n732), .B(n10351), .Z(n10350) );
  IV U10029 ( .A(n10346), .Z(n10348) );
  XOR U10030 ( .A(n10352), .B(n10353), .Z(n10346) );
  AND U10031 ( .A(n716), .B(n10345), .Z(n10353) );
  XNOR U10032 ( .A(n10343), .B(n10352), .Z(n10345) );
  XNOR U10033 ( .A(n10354), .B(n10355), .Z(n10343) );
  AND U10034 ( .A(n720), .B(n10356), .Z(n10355) );
  XOR U10035 ( .A(p_input[1020]), .B(n10354), .Z(n10356) );
  XNOR U10036 ( .A(n10357), .B(n10358), .Z(n10354) );
  AND U10037 ( .A(n724), .B(n10359), .Z(n10358) );
  XOR U10038 ( .A(n10360), .B(n10361), .Z(n10352) );
  AND U10039 ( .A(n728), .B(n10351), .Z(n10361) );
  XNOR U10040 ( .A(n10362), .B(n10349), .Z(n10351) );
  XOR U10041 ( .A(n10363), .B(n10364), .Z(n10349) );
  AND U10042 ( .A(n751), .B(n10365), .Z(n10364) );
  IV U10043 ( .A(n10360), .Z(n10362) );
  XOR U10044 ( .A(n10366), .B(n10367), .Z(n10360) );
  AND U10045 ( .A(n735), .B(n10359), .Z(n10367) );
  XNOR U10046 ( .A(n10357), .B(n10366), .Z(n10359) );
  XNOR U10047 ( .A(n10368), .B(n10369), .Z(n10357) );
  AND U10048 ( .A(n739), .B(n10370), .Z(n10369) );
  XOR U10049 ( .A(p_input[1052]), .B(n10368), .Z(n10370) );
  XNOR U10050 ( .A(n10371), .B(n10372), .Z(n10368) );
  AND U10051 ( .A(n743), .B(n10373), .Z(n10372) );
  XOR U10052 ( .A(n10374), .B(n10375), .Z(n10366) );
  AND U10053 ( .A(n747), .B(n10365), .Z(n10375) );
  XNOR U10054 ( .A(n10376), .B(n10363), .Z(n10365) );
  XOR U10055 ( .A(n10377), .B(n10378), .Z(n10363) );
  AND U10056 ( .A(n770), .B(n10379), .Z(n10378) );
  IV U10057 ( .A(n10374), .Z(n10376) );
  XOR U10058 ( .A(n10380), .B(n10381), .Z(n10374) );
  AND U10059 ( .A(n754), .B(n10373), .Z(n10381) );
  XNOR U10060 ( .A(n10371), .B(n10380), .Z(n10373) );
  XNOR U10061 ( .A(n10382), .B(n10383), .Z(n10371) );
  AND U10062 ( .A(n758), .B(n10384), .Z(n10383) );
  XOR U10063 ( .A(p_input[1084]), .B(n10382), .Z(n10384) );
  XNOR U10064 ( .A(n10385), .B(n10386), .Z(n10382) );
  AND U10065 ( .A(n762), .B(n10387), .Z(n10386) );
  XOR U10066 ( .A(n10388), .B(n10389), .Z(n10380) );
  AND U10067 ( .A(n766), .B(n10379), .Z(n10389) );
  XNOR U10068 ( .A(n10390), .B(n10377), .Z(n10379) );
  XOR U10069 ( .A(n10391), .B(n10392), .Z(n10377) );
  AND U10070 ( .A(n789), .B(n10393), .Z(n10392) );
  IV U10071 ( .A(n10388), .Z(n10390) );
  XOR U10072 ( .A(n10394), .B(n10395), .Z(n10388) );
  AND U10073 ( .A(n773), .B(n10387), .Z(n10395) );
  XNOR U10074 ( .A(n10385), .B(n10394), .Z(n10387) );
  XNOR U10075 ( .A(n10396), .B(n10397), .Z(n10385) );
  AND U10076 ( .A(n777), .B(n10398), .Z(n10397) );
  XOR U10077 ( .A(p_input[1116]), .B(n10396), .Z(n10398) );
  XNOR U10078 ( .A(n10399), .B(n10400), .Z(n10396) );
  AND U10079 ( .A(n781), .B(n10401), .Z(n10400) );
  XOR U10080 ( .A(n10402), .B(n10403), .Z(n10394) );
  AND U10081 ( .A(n785), .B(n10393), .Z(n10403) );
  XNOR U10082 ( .A(n10404), .B(n10391), .Z(n10393) );
  XOR U10083 ( .A(n10405), .B(n10406), .Z(n10391) );
  AND U10084 ( .A(n808), .B(n10407), .Z(n10406) );
  IV U10085 ( .A(n10402), .Z(n10404) );
  XOR U10086 ( .A(n10408), .B(n10409), .Z(n10402) );
  AND U10087 ( .A(n792), .B(n10401), .Z(n10409) );
  XNOR U10088 ( .A(n10399), .B(n10408), .Z(n10401) );
  XNOR U10089 ( .A(n10410), .B(n10411), .Z(n10399) );
  AND U10090 ( .A(n796), .B(n10412), .Z(n10411) );
  XOR U10091 ( .A(p_input[1148]), .B(n10410), .Z(n10412) );
  XNOR U10092 ( .A(n10413), .B(n10414), .Z(n10410) );
  AND U10093 ( .A(n800), .B(n10415), .Z(n10414) );
  XOR U10094 ( .A(n10416), .B(n10417), .Z(n10408) );
  AND U10095 ( .A(n804), .B(n10407), .Z(n10417) );
  XNOR U10096 ( .A(n10418), .B(n10405), .Z(n10407) );
  XOR U10097 ( .A(n10419), .B(n10420), .Z(n10405) );
  AND U10098 ( .A(n827), .B(n10421), .Z(n10420) );
  IV U10099 ( .A(n10416), .Z(n10418) );
  XOR U10100 ( .A(n10422), .B(n10423), .Z(n10416) );
  AND U10101 ( .A(n811), .B(n10415), .Z(n10423) );
  XNOR U10102 ( .A(n10413), .B(n10422), .Z(n10415) );
  XNOR U10103 ( .A(n10424), .B(n10425), .Z(n10413) );
  AND U10104 ( .A(n815), .B(n10426), .Z(n10425) );
  XOR U10105 ( .A(p_input[1180]), .B(n10424), .Z(n10426) );
  XNOR U10106 ( .A(n10427), .B(n10428), .Z(n10424) );
  AND U10107 ( .A(n819), .B(n10429), .Z(n10428) );
  XOR U10108 ( .A(n10430), .B(n10431), .Z(n10422) );
  AND U10109 ( .A(n823), .B(n10421), .Z(n10431) );
  XNOR U10110 ( .A(n10432), .B(n10419), .Z(n10421) );
  XOR U10111 ( .A(n10433), .B(n10434), .Z(n10419) );
  AND U10112 ( .A(n846), .B(n10435), .Z(n10434) );
  IV U10113 ( .A(n10430), .Z(n10432) );
  XOR U10114 ( .A(n10436), .B(n10437), .Z(n10430) );
  AND U10115 ( .A(n830), .B(n10429), .Z(n10437) );
  XNOR U10116 ( .A(n10427), .B(n10436), .Z(n10429) );
  XNOR U10117 ( .A(n10438), .B(n10439), .Z(n10427) );
  AND U10118 ( .A(n834), .B(n10440), .Z(n10439) );
  XOR U10119 ( .A(p_input[1212]), .B(n10438), .Z(n10440) );
  XNOR U10120 ( .A(n10441), .B(n10442), .Z(n10438) );
  AND U10121 ( .A(n838), .B(n10443), .Z(n10442) );
  XOR U10122 ( .A(n10444), .B(n10445), .Z(n10436) );
  AND U10123 ( .A(n842), .B(n10435), .Z(n10445) );
  XNOR U10124 ( .A(n10446), .B(n10433), .Z(n10435) );
  XOR U10125 ( .A(n10447), .B(n10448), .Z(n10433) );
  AND U10126 ( .A(n865), .B(n10449), .Z(n10448) );
  IV U10127 ( .A(n10444), .Z(n10446) );
  XOR U10128 ( .A(n10450), .B(n10451), .Z(n10444) );
  AND U10129 ( .A(n849), .B(n10443), .Z(n10451) );
  XNOR U10130 ( .A(n10441), .B(n10450), .Z(n10443) );
  XNOR U10131 ( .A(n10452), .B(n10453), .Z(n10441) );
  AND U10132 ( .A(n853), .B(n10454), .Z(n10453) );
  XOR U10133 ( .A(p_input[1244]), .B(n10452), .Z(n10454) );
  XNOR U10134 ( .A(n10455), .B(n10456), .Z(n10452) );
  AND U10135 ( .A(n857), .B(n10457), .Z(n10456) );
  XOR U10136 ( .A(n10458), .B(n10459), .Z(n10450) );
  AND U10137 ( .A(n861), .B(n10449), .Z(n10459) );
  XNOR U10138 ( .A(n10460), .B(n10447), .Z(n10449) );
  XOR U10139 ( .A(n10461), .B(n10462), .Z(n10447) );
  AND U10140 ( .A(n884), .B(n10463), .Z(n10462) );
  IV U10141 ( .A(n10458), .Z(n10460) );
  XOR U10142 ( .A(n10464), .B(n10465), .Z(n10458) );
  AND U10143 ( .A(n868), .B(n10457), .Z(n10465) );
  XNOR U10144 ( .A(n10455), .B(n10464), .Z(n10457) );
  XNOR U10145 ( .A(n10466), .B(n10467), .Z(n10455) );
  AND U10146 ( .A(n872), .B(n10468), .Z(n10467) );
  XOR U10147 ( .A(p_input[1276]), .B(n10466), .Z(n10468) );
  XNOR U10148 ( .A(n10469), .B(n10470), .Z(n10466) );
  AND U10149 ( .A(n876), .B(n10471), .Z(n10470) );
  XOR U10150 ( .A(n10472), .B(n10473), .Z(n10464) );
  AND U10151 ( .A(n880), .B(n10463), .Z(n10473) );
  XNOR U10152 ( .A(n10474), .B(n10461), .Z(n10463) );
  XOR U10153 ( .A(n10475), .B(n10476), .Z(n10461) );
  AND U10154 ( .A(n903), .B(n10477), .Z(n10476) );
  IV U10155 ( .A(n10472), .Z(n10474) );
  XOR U10156 ( .A(n10478), .B(n10479), .Z(n10472) );
  AND U10157 ( .A(n887), .B(n10471), .Z(n10479) );
  XNOR U10158 ( .A(n10469), .B(n10478), .Z(n10471) );
  XNOR U10159 ( .A(n10480), .B(n10481), .Z(n10469) );
  AND U10160 ( .A(n891), .B(n10482), .Z(n10481) );
  XOR U10161 ( .A(p_input[1308]), .B(n10480), .Z(n10482) );
  XNOR U10162 ( .A(n10483), .B(n10484), .Z(n10480) );
  AND U10163 ( .A(n895), .B(n10485), .Z(n10484) );
  XOR U10164 ( .A(n10486), .B(n10487), .Z(n10478) );
  AND U10165 ( .A(n899), .B(n10477), .Z(n10487) );
  XNOR U10166 ( .A(n10488), .B(n10475), .Z(n10477) );
  XOR U10167 ( .A(n10489), .B(n10490), .Z(n10475) );
  AND U10168 ( .A(n922), .B(n10491), .Z(n10490) );
  IV U10169 ( .A(n10486), .Z(n10488) );
  XOR U10170 ( .A(n10492), .B(n10493), .Z(n10486) );
  AND U10171 ( .A(n906), .B(n10485), .Z(n10493) );
  XNOR U10172 ( .A(n10483), .B(n10492), .Z(n10485) );
  XNOR U10173 ( .A(n10494), .B(n10495), .Z(n10483) );
  AND U10174 ( .A(n910), .B(n10496), .Z(n10495) );
  XOR U10175 ( .A(p_input[1340]), .B(n10494), .Z(n10496) );
  XNOR U10176 ( .A(n10497), .B(n10498), .Z(n10494) );
  AND U10177 ( .A(n914), .B(n10499), .Z(n10498) );
  XOR U10178 ( .A(n10500), .B(n10501), .Z(n10492) );
  AND U10179 ( .A(n918), .B(n10491), .Z(n10501) );
  XNOR U10180 ( .A(n10502), .B(n10489), .Z(n10491) );
  XOR U10181 ( .A(n10503), .B(n10504), .Z(n10489) );
  AND U10182 ( .A(n941), .B(n10505), .Z(n10504) );
  IV U10183 ( .A(n10500), .Z(n10502) );
  XOR U10184 ( .A(n10506), .B(n10507), .Z(n10500) );
  AND U10185 ( .A(n925), .B(n10499), .Z(n10507) );
  XNOR U10186 ( .A(n10497), .B(n10506), .Z(n10499) );
  XNOR U10187 ( .A(n10508), .B(n10509), .Z(n10497) );
  AND U10188 ( .A(n929), .B(n10510), .Z(n10509) );
  XOR U10189 ( .A(p_input[1372]), .B(n10508), .Z(n10510) );
  XNOR U10190 ( .A(n10511), .B(n10512), .Z(n10508) );
  AND U10191 ( .A(n933), .B(n10513), .Z(n10512) );
  XOR U10192 ( .A(n10514), .B(n10515), .Z(n10506) );
  AND U10193 ( .A(n937), .B(n10505), .Z(n10515) );
  XNOR U10194 ( .A(n10516), .B(n10503), .Z(n10505) );
  XOR U10195 ( .A(n10517), .B(n10518), .Z(n10503) );
  AND U10196 ( .A(n960), .B(n10519), .Z(n10518) );
  IV U10197 ( .A(n10514), .Z(n10516) );
  XOR U10198 ( .A(n10520), .B(n10521), .Z(n10514) );
  AND U10199 ( .A(n944), .B(n10513), .Z(n10521) );
  XNOR U10200 ( .A(n10511), .B(n10520), .Z(n10513) );
  XNOR U10201 ( .A(n10522), .B(n10523), .Z(n10511) );
  AND U10202 ( .A(n948), .B(n10524), .Z(n10523) );
  XOR U10203 ( .A(p_input[1404]), .B(n10522), .Z(n10524) );
  XNOR U10204 ( .A(n10525), .B(n10526), .Z(n10522) );
  AND U10205 ( .A(n952), .B(n10527), .Z(n10526) );
  XOR U10206 ( .A(n10528), .B(n10529), .Z(n10520) );
  AND U10207 ( .A(n956), .B(n10519), .Z(n10529) );
  XNOR U10208 ( .A(n10530), .B(n10517), .Z(n10519) );
  XOR U10209 ( .A(n10531), .B(n10532), .Z(n10517) );
  AND U10210 ( .A(n979), .B(n10533), .Z(n10532) );
  IV U10211 ( .A(n10528), .Z(n10530) );
  XOR U10212 ( .A(n10534), .B(n10535), .Z(n10528) );
  AND U10213 ( .A(n963), .B(n10527), .Z(n10535) );
  XNOR U10214 ( .A(n10525), .B(n10534), .Z(n10527) );
  XNOR U10215 ( .A(n10536), .B(n10537), .Z(n10525) );
  AND U10216 ( .A(n967), .B(n10538), .Z(n10537) );
  XOR U10217 ( .A(p_input[1436]), .B(n10536), .Z(n10538) );
  XNOR U10218 ( .A(n10539), .B(n10540), .Z(n10536) );
  AND U10219 ( .A(n971), .B(n10541), .Z(n10540) );
  XOR U10220 ( .A(n10542), .B(n10543), .Z(n10534) );
  AND U10221 ( .A(n975), .B(n10533), .Z(n10543) );
  XNOR U10222 ( .A(n10544), .B(n10531), .Z(n10533) );
  XOR U10223 ( .A(n10545), .B(n10546), .Z(n10531) );
  AND U10224 ( .A(n998), .B(n10547), .Z(n10546) );
  IV U10225 ( .A(n10542), .Z(n10544) );
  XOR U10226 ( .A(n10548), .B(n10549), .Z(n10542) );
  AND U10227 ( .A(n982), .B(n10541), .Z(n10549) );
  XNOR U10228 ( .A(n10539), .B(n10548), .Z(n10541) );
  XNOR U10229 ( .A(n10550), .B(n10551), .Z(n10539) );
  AND U10230 ( .A(n986), .B(n10552), .Z(n10551) );
  XOR U10231 ( .A(p_input[1468]), .B(n10550), .Z(n10552) );
  XNOR U10232 ( .A(n10553), .B(n10554), .Z(n10550) );
  AND U10233 ( .A(n990), .B(n10555), .Z(n10554) );
  XOR U10234 ( .A(n10556), .B(n10557), .Z(n10548) );
  AND U10235 ( .A(n994), .B(n10547), .Z(n10557) );
  XNOR U10236 ( .A(n10558), .B(n10545), .Z(n10547) );
  XOR U10237 ( .A(n10559), .B(n10560), .Z(n10545) );
  AND U10238 ( .A(n1017), .B(n10561), .Z(n10560) );
  IV U10239 ( .A(n10556), .Z(n10558) );
  XOR U10240 ( .A(n10562), .B(n10563), .Z(n10556) );
  AND U10241 ( .A(n1001), .B(n10555), .Z(n10563) );
  XNOR U10242 ( .A(n10553), .B(n10562), .Z(n10555) );
  XNOR U10243 ( .A(n10564), .B(n10565), .Z(n10553) );
  AND U10244 ( .A(n1005), .B(n10566), .Z(n10565) );
  XOR U10245 ( .A(p_input[1500]), .B(n10564), .Z(n10566) );
  XNOR U10246 ( .A(n10567), .B(n10568), .Z(n10564) );
  AND U10247 ( .A(n1009), .B(n10569), .Z(n10568) );
  XOR U10248 ( .A(n10570), .B(n10571), .Z(n10562) );
  AND U10249 ( .A(n1013), .B(n10561), .Z(n10571) );
  XNOR U10250 ( .A(n10572), .B(n10559), .Z(n10561) );
  XOR U10251 ( .A(n10573), .B(n10574), .Z(n10559) );
  AND U10252 ( .A(n1036), .B(n10575), .Z(n10574) );
  IV U10253 ( .A(n10570), .Z(n10572) );
  XOR U10254 ( .A(n10576), .B(n10577), .Z(n10570) );
  AND U10255 ( .A(n1020), .B(n10569), .Z(n10577) );
  XNOR U10256 ( .A(n10567), .B(n10576), .Z(n10569) );
  XNOR U10257 ( .A(n10578), .B(n10579), .Z(n10567) );
  AND U10258 ( .A(n1024), .B(n10580), .Z(n10579) );
  XOR U10259 ( .A(p_input[1532]), .B(n10578), .Z(n10580) );
  XNOR U10260 ( .A(n10581), .B(n10582), .Z(n10578) );
  AND U10261 ( .A(n1028), .B(n10583), .Z(n10582) );
  XOR U10262 ( .A(n10584), .B(n10585), .Z(n10576) );
  AND U10263 ( .A(n1032), .B(n10575), .Z(n10585) );
  XNOR U10264 ( .A(n10586), .B(n10573), .Z(n10575) );
  XOR U10265 ( .A(n10587), .B(n10588), .Z(n10573) );
  AND U10266 ( .A(n1055), .B(n10589), .Z(n10588) );
  IV U10267 ( .A(n10584), .Z(n10586) );
  XOR U10268 ( .A(n10590), .B(n10591), .Z(n10584) );
  AND U10269 ( .A(n1039), .B(n10583), .Z(n10591) );
  XNOR U10270 ( .A(n10581), .B(n10590), .Z(n10583) );
  XNOR U10271 ( .A(n10592), .B(n10593), .Z(n10581) );
  AND U10272 ( .A(n1043), .B(n10594), .Z(n10593) );
  XOR U10273 ( .A(p_input[1564]), .B(n10592), .Z(n10594) );
  XNOR U10274 ( .A(n10595), .B(n10596), .Z(n10592) );
  AND U10275 ( .A(n1047), .B(n10597), .Z(n10596) );
  XOR U10276 ( .A(n10598), .B(n10599), .Z(n10590) );
  AND U10277 ( .A(n1051), .B(n10589), .Z(n10599) );
  XNOR U10278 ( .A(n10600), .B(n10587), .Z(n10589) );
  XOR U10279 ( .A(n10601), .B(n10602), .Z(n10587) );
  AND U10280 ( .A(n1074), .B(n10603), .Z(n10602) );
  IV U10281 ( .A(n10598), .Z(n10600) );
  XOR U10282 ( .A(n10604), .B(n10605), .Z(n10598) );
  AND U10283 ( .A(n1058), .B(n10597), .Z(n10605) );
  XNOR U10284 ( .A(n10595), .B(n10604), .Z(n10597) );
  XNOR U10285 ( .A(n10606), .B(n10607), .Z(n10595) );
  AND U10286 ( .A(n1062), .B(n10608), .Z(n10607) );
  XOR U10287 ( .A(p_input[1596]), .B(n10606), .Z(n10608) );
  XNOR U10288 ( .A(n10609), .B(n10610), .Z(n10606) );
  AND U10289 ( .A(n1066), .B(n10611), .Z(n10610) );
  XOR U10290 ( .A(n10612), .B(n10613), .Z(n10604) );
  AND U10291 ( .A(n1070), .B(n10603), .Z(n10613) );
  XNOR U10292 ( .A(n10614), .B(n10601), .Z(n10603) );
  XOR U10293 ( .A(n10615), .B(n10616), .Z(n10601) );
  AND U10294 ( .A(n1093), .B(n10617), .Z(n10616) );
  IV U10295 ( .A(n10612), .Z(n10614) );
  XOR U10296 ( .A(n10618), .B(n10619), .Z(n10612) );
  AND U10297 ( .A(n1077), .B(n10611), .Z(n10619) );
  XNOR U10298 ( .A(n10609), .B(n10618), .Z(n10611) );
  XNOR U10299 ( .A(n10620), .B(n10621), .Z(n10609) );
  AND U10300 ( .A(n1081), .B(n10622), .Z(n10621) );
  XOR U10301 ( .A(p_input[1628]), .B(n10620), .Z(n10622) );
  XNOR U10302 ( .A(n10623), .B(n10624), .Z(n10620) );
  AND U10303 ( .A(n1085), .B(n10625), .Z(n10624) );
  XOR U10304 ( .A(n10626), .B(n10627), .Z(n10618) );
  AND U10305 ( .A(n1089), .B(n10617), .Z(n10627) );
  XNOR U10306 ( .A(n10628), .B(n10615), .Z(n10617) );
  XOR U10307 ( .A(n10629), .B(n10630), .Z(n10615) );
  AND U10308 ( .A(n1112), .B(n10631), .Z(n10630) );
  IV U10309 ( .A(n10626), .Z(n10628) );
  XOR U10310 ( .A(n10632), .B(n10633), .Z(n10626) );
  AND U10311 ( .A(n1096), .B(n10625), .Z(n10633) );
  XNOR U10312 ( .A(n10623), .B(n10632), .Z(n10625) );
  XNOR U10313 ( .A(n10634), .B(n10635), .Z(n10623) );
  AND U10314 ( .A(n1100), .B(n10636), .Z(n10635) );
  XOR U10315 ( .A(p_input[1660]), .B(n10634), .Z(n10636) );
  XNOR U10316 ( .A(n10637), .B(n10638), .Z(n10634) );
  AND U10317 ( .A(n1104), .B(n10639), .Z(n10638) );
  XOR U10318 ( .A(n10640), .B(n10641), .Z(n10632) );
  AND U10319 ( .A(n1108), .B(n10631), .Z(n10641) );
  XNOR U10320 ( .A(n10642), .B(n10629), .Z(n10631) );
  XOR U10321 ( .A(n10643), .B(n10644), .Z(n10629) );
  AND U10322 ( .A(n1131), .B(n10645), .Z(n10644) );
  IV U10323 ( .A(n10640), .Z(n10642) );
  XOR U10324 ( .A(n10646), .B(n10647), .Z(n10640) );
  AND U10325 ( .A(n1115), .B(n10639), .Z(n10647) );
  XNOR U10326 ( .A(n10637), .B(n10646), .Z(n10639) );
  XNOR U10327 ( .A(n10648), .B(n10649), .Z(n10637) );
  AND U10328 ( .A(n1119), .B(n10650), .Z(n10649) );
  XOR U10329 ( .A(p_input[1692]), .B(n10648), .Z(n10650) );
  XNOR U10330 ( .A(n10651), .B(n10652), .Z(n10648) );
  AND U10331 ( .A(n1123), .B(n10653), .Z(n10652) );
  XOR U10332 ( .A(n10654), .B(n10655), .Z(n10646) );
  AND U10333 ( .A(n1127), .B(n10645), .Z(n10655) );
  XNOR U10334 ( .A(n10656), .B(n10643), .Z(n10645) );
  XOR U10335 ( .A(n10657), .B(n10658), .Z(n10643) );
  AND U10336 ( .A(n1150), .B(n10659), .Z(n10658) );
  IV U10337 ( .A(n10654), .Z(n10656) );
  XOR U10338 ( .A(n10660), .B(n10661), .Z(n10654) );
  AND U10339 ( .A(n1134), .B(n10653), .Z(n10661) );
  XNOR U10340 ( .A(n10651), .B(n10660), .Z(n10653) );
  XNOR U10341 ( .A(n10662), .B(n10663), .Z(n10651) );
  AND U10342 ( .A(n1138), .B(n10664), .Z(n10663) );
  XOR U10343 ( .A(p_input[1724]), .B(n10662), .Z(n10664) );
  XNOR U10344 ( .A(n10665), .B(n10666), .Z(n10662) );
  AND U10345 ( .A(n1142), .B(n10667), .Z(n10666) );
  XOR U10346 ( .A(n10668), .B(n10669), .Z(n10660) );
  AND U10347 ( .A(n1146), .B(n10659), .Z(n10669) );
  XNOR U10348 ( .A(n10670), .B(n10657), .Z(n10659) );
  XOR U10349 ( .A(n10671), .B(n10672), .Z(n10657) );
  AND U10350 ( .A(n1169), .B(n10673), .Z(n10672) );
  IV U10351 ( .A(n10668), .Z(n10670) );
  XOR U10352 ( .A(n10674), .B(n10675), .Z(n10668) );
  AND U10353 ( .A(n1153), .B(n10667), .Z(n10675) );
  XNOR U10354 ( .A(n10665), .B(n10674), .Z(n10667) );
  XNOR U10355 ( .A(n10676), .B(n10677), .Z(n10665) );
  AND U10356 ( .A(n1157), .B(n10678), .Z(n10677) );
  XOR U10357 ( .A(p_input[1756]), .B(n10676), .Z(n10678) );
  XNOR U10358 ( .A(n10679), .B(n10680), .Z(n10676) );
  AND U10359 ( .A(n1161), .B(n10681), .Z(n10680) );
  XOR U10360 ( .A(n10682), .B(n10683), .Z(n10674) );
  AND U10361 ( .A(n1165), .B(n10673), .Z(n10683) );
  XNOR U10362 ( .A(n10684), .B(n10671), .Z(n10673) );
  XOR U10363 ( .A(n10685), .B(n10686), .Z(n10671) );
  AND U10364 ( .A(n1188), .B(n10687), .Z(n10686) );
  IV U10365 ( .A(n10682), .Z(n10684) );
  XOR U10366 ( .A(n10688), .B(n10689), .Z(n10682) );
  AND U10367 ( .A(n1172), .B(n10681), .Z(n10689) );
  XNOR U10368 ( .A(n10679), .B(n10688), .Z(n10681) );
  XNOR U10369 ( .A(n10690), .B(n10691), .Z(n10679) );
  AND U10370 ( .A(n1176), .B(n10692), .Z(n10691) );
  XOR U10371 ( .A(p_input[1788]), .B(n10690), .Z(n10692) );
  XNOR U10372 ( .A(n10693), .B(n10694), .Z(n10690) );
  AND U10373 ( .A(n1180), .B(n10695), .Z(n10694) );
  XOR U10374 ( .A(n10696), .B(n10697), .Z(n10688) );
  AND U10375 ( .A(n1184), .B(n10687), .Z(n10697) );
  XNOR U10376 ( .A(n10698), .B(n10685), .Z(n10687) );
  XOR U10377 ( .A(n10699), .B(n10700), .Z(n10685) );
  AND U10378 ( .A(n1207), .B(n10701), .Z(n10700) );
  IV U10379 ( .A(n10696), .Z(n10698) );
  XOR U10380 ( .A(n10702), .B(n10703), .Z(n10696) );
  AND U10381 ( .A(n1191), .B(n10695), .Z(n10703) );
  XNOR U10382 ( .A(n10693), .B(n10702), .Z(n10695) );
  XNOR U10383 ( .A(n10704), .B(n10705), .Z(n10693) );
  AND U10384 ( .A(n1195), .B(n10706), .Z(n10705) );
  XOR U10385 ( .A(p_input[1820]), .B(n10704), .Z(n10706) );
  XNOR U10386 ( .A(n10707), .B(n10708), .Z(n10704) );
  AND U10387 ( .A(n1199), .B(n10709), .Z(n10708) );
  XOR U10388 ( .A(n10710), .B(n10711), .Z(n10702) );
  AND U10389 ( .A(n1203), .B(n10701), .Z(n10711) );
  XNOR U10390 ( .A(n10712), .B(n10699), .Z(n10701) );
  XOR U10391 ( .A(n10713), .B(n10714), .Z(n10699) );
  AND U10392 ( .A(n1226), .B(n10715), .Z(n10714) );
  IV U10393 ( .A(n10710), .Z(n10712) );
  XOR U10394 ( .A(n10716), .B(n10717), .Z(n10710) );
  AND U10395 ( .A(n1210), .B(n10709), .Z(n10717) );
  XNOR U10396 ( .A(n10707), .B(n10716), .Z(n10709) );
  XNOR U10397 ( .A(n10718), .B(n10719), .Z(n10707) );
  AND U10398 ( .A(n1214), .B(n10720), .Z(n10719) );
  XOR U10399 ( .A(p_input[1852]), .B(n10718), .Z(n10720) );
  XNOR U10400 ( .A(n10721), .B(n10722), .Z(n10718) );
  AND U10401 ( .A(n1218), .B(n10723), .Z(n10722) );
  XOR U10402 ( .A(n10724), .B(n10725), .Z(n10716) );
  AND U10403 ( .A(n1222), .B(n10715), .Z(n10725) );
  XNOR U10404 ( .A(n10726), .B(n10713), .Z(n10715) );
  XOR U10405 ( .A(n10727), .B(n10728), .Z(n10713) );
  AND U10406 ( .A(n1245), .B(n10729), .Z(n10728) );
  IV U10407 ( .A(n10724), .Z(n10726) );
  XOR U10408 ( .A(n10730), .B(n10731), .Z(n10724) );
  AND U10409 ( .A(n1229), .B(n10723), .Z(n10731) );
  XNOR U10410 ( .A(n10721), .B(n10730), .Z(n10723) );
  XNOR U10411 ( .A(n10732), .B(n10733), .Z(n10721) );
  AND U10412 ( .A(n1233), .B(n10734), .Z(n10733) );
  XOR U10413 ( .A(p_input[1884]), .B(n10732), .Z(n10734) );
  XNOR U10414 ( .A(n10735), .B(n10736), .Z(n10732) );
  AND U10415 ( .A(n1237), .B(n10737), .Z(n10736) );
  XOR U10416 ( .A(n10738), .B(n10739), .Z(n10730) );
  AND U10417 ( .A(n1241), .B(n10729), .Z(n10739) );
  XNOR U10418 ( .A(n10740), .B(n10727), .Z(n10729) );
  XOR U10419 ( .A(n10741), .B(n10742), .Z(n10727) );
  AND U10420 ( .A(n1264), .B(n10743), .Z(n10742) );
  IV U10421 ( .A(n10738), .Z(n10740) );
  XOR U10422 ( .A(n10744), .B(n10745), .Z(n10738) );
  AND U10423 ( .A(n1248), .B(n10737), .Z(n10745) );
  XNOR U10424 ( .A(n10735), .B(n10744), .Z(n10737) );
  XNOR U10425 ( .A(n10746), .B(n10747), .Z(n10735) );
  AND U10426 ( .A(n1252), .B(n10748), .Z(n10747) );
  XOR U10427 ( .A(p_input[1916]), .B(n10746), .Z(n10748) );
  XNOR U10428 ( .A(n10749), .B(n10750), .Z(n10746) );
  AND U10429 ( .A(n1256), .B(n10751), .Z(n10750) );
  XOR U10430 ( .A(n10752), .B(n10753), .Z(n10744) );
  AND U10431 ( .A(n1260), .B(n10743), .Z(n10753) );
  XNOR U10432 ( .A(n10754), .B(n10741), .Z(n10743) );
  XOR U10433 ( .A(n10755), .B(n10756), .Z(n10741) );
  AND U10434 ( .A(n1282), .B(n10757), .Z(n10756) );
  IV U10435 ( .A(n10752), .Z(n10754) );
  XOR U10436 ( .A(n10758), .B(n10759), .Z(n10752) );
  AND U10437 ( .A(n1267), .B(n10751), .Z(n10759) );
  XNOR U10438 ( .A(n10749), .B(n10758), .Z(n10751) );
  XNOR U10439 ( .A(n10760), .B(n10761), .Z(n10749) );
  AND U10440 ( .A(n1271), .B(n10762), .Z(n10761) );
  XOR U10441 ( .A(p_input[1948]), .B(n10760), .Z(n10762) );
  XOR U10442 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][28] ), .B(n10763), 
        .Z(n10760) );
  AND U10443 ( .A(n1274), .B(n10764), .Z(n10763) );
  XOR U10444 ( .A(n10765), .B(n10766), .Z(n10758) );
  AND U10445 ( .A(n1278), .B(n10757), .Z(n10766) );
  XNOR U10446 ( .A(n10767), .B(n10755), .Z(n10757) );
  XOR U10447 ( .A(\knn_comb_/min_val_out[0][28] ), .B(n10768), .Z(n10755) );
  AND U10448 ( .A(n1290), .B(n10769), .Z(n10768) );
  IV U10449 ( .A(n10765), .Z(n10767) );
  XOR U10450 ( .A(n10770), .B(n10771), .Z(n10765) );
  AND U10451 ( .A(n1285), .B(n10764), .Z(n10771) );
  XOR U10452 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][28] ), .B(n10770), 
        .Z(n10764) );
  XOR U10453 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .B(n10772), 
        .Z(n10770) );
  AND U10454 ( .A(n1287), .B(n10769), .Z(n10772) );
  XOR U10455 ( .A(\knn_comb_/min_val_out[0][28] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .Z(n10769) );
  XOR U10456 ( .A(n83), .B(n10773), .Z(o[27]) );
  AND U10457 ( .A(n122), .B(n10774), .Z(n83) );
  XOR U10458 ( .A(n84), .B(n10773), .Z(n10774) );
  XOR U10459 ( .A(n10775), .B(n10776), .Z(n10773) );
  AND U10460 ( .A(n142), .B(n10777), .Z(n10776) );
  XOR U10461 ( .A(n10778), .B(n11), .Z(n84) );
  AND U10462 ( .A(n125), .B(n10779), .Z(n11) );
  XOR U10463 ( .A(n12), .B(n10778), .Z(n10779) );
  XOR U10464 ( .A(n10780), .B(n10781), .Z(n12) );
  AND U10465 ( .A(n130), .B(n10782), .Z(n10781) );
  XOR U10466 ( .A(p_input[27]), .B(n10780), .Z(n10782) );
  XNOR U10467 ( .A(n10783), .B(n10784), .Z(n10780) );
  AND U10468 ( .A(n134), .B(n10785), .Z(n10784) );
  XOR U10469 ( .A(n10786), .B(n10787), .Z(n10778) );
  AND U10470 ( .A(n138), .B(n10777), .Z(n10787) );
  XNOR U10471 ( .A(n10788), .B(n10775), .Z(n10777) );
  XOR U10472 ( .A(n10789), .B(n10790), .Z(n10775) );
  AND U10473 ( .A(n162), .B(n10791), .Z(n10790) );
  IV U10474 ( .A(n10786), .Z(n10788) );
  XOR U10475 ( .A(n10792), .B(n10793), .Z(n10786) );
  AND U10476 ( .A(n146), .B(n10785), .Z(n10793) );
  XNOR U10477 ( .A(n10783), .B(n10792), .Z(n10785) );
  XNOR U10478 ( .A(n10794), .B(n10795), .Z(n10783) );
  AND U10479 ( .A(n150), .B(n10796), .Z(n10795) );
  XOR U10480 ( .A(p_input[59]), .B(n10794), .Z(n10796) );
  XNOR U10481 ( .A(n10797), .B(n10798), .Z(n10794) );
  AND U10482 ( .A(n154), .B(n10799), .Z(n10798) );
  XOR U10483 ( .A(n10800), .B(n10801), .Z(n10792) );
  AND U10484 ( .A(n158), .B(n10791), .Z(n10801) );
  XNOR U10485 ( .A(n10802), .B(n10789), .Z(n10791) );
  XOR U10486 ( .A(n10803), .B(n10804), .Z(n10789) );
  AND U10487 ( .A(n181), .B(n10805), .Z(n10804) );
  IV U10488 ( .A(n10800), .Z(n10802) );
  XOR U10489 ( .A(n10806), .B(n10807), .Z(n10800) );
  AND U10490 ( .A(n165), .B(n10799), .Z(n10807) );
  XNOR U10491 ( .A(n10797), .B(n10806), .Z(n10799) );
  XNOR U10492 ( .A(n10808), .B(n10809), .Z(n10797) );
  AND U10493 ( .A(n169), .B(n10810), .Z(n10809) );
  XOR U10494 ( .A(p_input[91]), .B(n10808), .Z(n10810) );
  XNOR U10495 ( .A(n10811), .B(n10812), .Z(n10808) );
  AND U10496 ( .A(n173), .B(n10813), .Z(n10812) );
  XOR U10497 ( .A(n10814), .B(n10815), .Z(n10806) );
  AND U10498 ( .A(n177), .B(n10805), .Z(n10815) );
  XNOR U10499 ( .A(n10816), .B(n10803), .Z(n10805) );
  XOR U10500 ( .A(n10817), .B(n10818), .Z(n10803) );
  AND U10501 ( .A(n200), .B(n10819), .Z(n10818) );
  IV U10502 ( .A(n10814), .Z(n10816) );
  XOR U10503 ( .A(n10820), .B(n10821), .Z(n10814) );
  AND U10504 ( .A(n184), .B(n10813), .Z(n10821) );
  XNOR U10505 ( .A(n10811), .B(n10820), .Z(n10813) );
  XNOR U10506 ( .A(n10822), .B(n10823), .Z(n10811) );
  AND U10507 ( .A(n188), .B(n10824), .Z(n10823) );
  XOR U10508 ( .A(p_input[123]), .B(n10822), .Z(n10824) );
  XNOR U10509 ( .A(n10825), .B(n10826), .Z(n10822) );
  AND U10510 ( .A(n192), .B(n10827), .Z(n10826) );
  XOR U10511 ( .A(n10828), .B(n10829), .Z(n10820) );
  AND U10512 ( .A(n196), .B(n10819), .Z(n10829) );
  XNOR U10513 ( .A(n10830), .B(n10817), .Z(n10819) );
  XOR U10514 ( .A(n10831), .B(n10832), .Z(n10817) );
  AND U10515 ( .A(n219), .B(n10833), .Z(n10832) );
  IV U10516 ( .A(n10828), .Z(n10830) );
  XOR U10517 ( .A(n10834), .B(n10835), .Z(n10828) );
  AND U10518 ( .A(n203), .B(n10827), .Z(n10835) );
  XNOR U10519 ( .A(n10825), .B(n10834), .Z(n10827) );
  XNOR U10520 ( .A(n10836), .B(n10837), .Z(n10825) );
  AND U10521 ( .A(n207), .B(n10838), .Z(n10837) );
  XOR U10522 ( .A(p_input[155]), .B(n10836), .Z(n10838) );
  XNOR U10523 ( .A(n10839), .B(n10840), .Z(n10836) );
  AND U10524 ( .A(n211), .B(n10841), .Z(n10840) );
  XOR U10525 ( .A(n10842), .B(n10843), .Z(n10834) );
  AND U10526 ( .A(n215), .B(n10833), .Z(n10843) );
  XNOR U10527 ( .A(n10844), .B(n10831), .Z(n10833) );
  XOR U10528 ( .A(n10845), .B(n10846), .Z(n10831) );
  AND U10529 ( .A(n238), .B(n10847), .Z(n10846) );
  IV U10530 ( .A(n10842), .Z(n10844) );
  XOR U10531 ( .A(n10848), .B(n10849), .Z(n10842) );
  AND U10532 ( .A(n222), .B(n10841), .Z(n10849) );
  XNOR U10533 ( .A(n10839), .B(n10848), .Z(n10841) );
  XNOR U10534 ( .A(n10850), .B(n10851), .Z(n10839) );
  AND U10535 ( .A(n226), .B(n10852), .Z(n10851) );
  XOR U10536 ( .A(p_input[187]), .B(n10850), .Z(n10852) );
  XNOR U10537 ( .A(n10853), .B(n10854), .Z(n10850) );
  AND U10538 ( .A(n230), .B(n10855), .Z(n10854) );
  XOR U10539 ( .A(n10856), .B(n10857), .Z(n10848) );
  AND U10540 ( .A(n234), .B(n10847), .Z(n10857) );
  XNOR U10541 ( .A(n10858), .B(n10845), .Z(n10847) );
  XOR U10542 ( .A(n10859), .B(n10860), .Z(n10845) );
  AND U10543 ( .A(n257), .B(n10861), .Z(n10860) );
  IV U10544 ( .A(n10856), .Z(n10858) );
  XOR U10545 ( .A(n10862), .B(n10863), .Z(n10856) );
  AND U10546 ( .A(n241), .B(n10855), .Z(n10863) );
  XNOR U10547 ( .A(n10853), .B(n10862), .Z(n10855) );
  XNOR U10548 ( .A(n10864), .B(n10865), .Z(n10853) );
  AND U10549 ( .A(n245), .B(n10866), .Z(n10865) );
  XOR U10550 ( .A(p_input[219]), .B(n10864), .Z(n10866) );
  XNOR U10551 ( .A(n10867), .B(n10868), .Z(n10864) );
  AND U10552 ( .A(n249), .B(n10869), .Z(n10868) );
  XOR U10553 ( .A(n10870), .B(n10871), .Z(n10862) );
  AND U10554 ( .A(n253), .B(n10861), .Z(n10871) );
  XNOR U10555 ( .A(n10872), .B(n10859), .Z(n10861) );
  XOR U10556 ( .A(n10873), .B(n10874), .Z(n10859) );
  AND U10557 ( .A(n276), .B(n10875), .Z(n10874) );
  IV U10558 ( .A(n10870), .Z(n10872) );
  XOR U10559 ( .A(n10876), .B(n10877), .Z(n10870) );
  AND U10560 ( .A(n260), .B(n10869), .Z(n10877) );
  XNOR U10561 ( .A(n10867), .B(n10876), .Z(n10869) );
  XNOR U10562 ( .A(n10878), .B(n10879), .Z(n10867) );
  AND U10563 ( .A(n264), .B(n10880), .Z(n10879) );
  XOR U10564 ( .A(p_input[251]), .B(n10878), .Z(n10880) );
  XNOR U10565 ( .A(n10881), .B(n10882), .Z(n10878) );
  AND U10566 ( .A(n268), .B(n10883), .Z(n10882) );
  XOR U10567 ( .A(n10884), .B(n10885), .Z(n10876) );
  AND U10568 ( .A(n272), .B(n10875), .Z(n10885) );
  XNOR U10569 ( .A(n10886), .B(n10873), .Z(n10875) );
  XOR U10570 ( .A(n10887), .B(n10888), .Z(n10873) );
  AND U10571 ( .A(n295), .B(n10889), .Z(n10888) );
  IV U10572 ( .A(n10884), .Z(n10886) );
  XOR U10573 ( .A(n10890), .B(n10891), .Z(n10884) );
  AND U10574 ( .A(n279), .B(n10883), .Z(n10891) );
  XNOR U10575 ( .A(n10881), .B(n10890), .Z(n10883) );
  XNOR U10576 ( .A(n10892), .B(n10893), .Z(n10881) );
  AND U10577 ( .A(n283), .B(n10894), .Z(n10893) );
  XOR U10578 ( .A(p_input[283]), .B(n10892), .Z(n10894) );
  XNOR U10579 ( .A(n10895), .B(n10896), .Z(n10892) );
  AND U10580 ( .A(n287), .B(n10897), .Z(n10896) );
  XOR U10581 ( .A(n10898), .B(n10899), .Z(n10890) );
  AND U10582 ( .A(n291), .B(n10889), .Z(n10899) );
  XNOR U10583 ( .A(n10900), .B(n10887), .Z(n10889) );
  XOR U10584 ( .A(n10901), .B(n10902), .Z(n10887) );
  AND U10585 ( .A(n314), .B(n10903), .Z(n10902) );
  IV U10586 ( .A(n10898), .Z(n10900) );
  XOR U10587 ( .A(n10904), .B(n10905), .Z(n10898) );
  AND U10588 ( .A(n298), .B(n10897), .Z(n10905) );
  XNOR U10589 ( .A(n10895), .B(n10904), .Z(n10897) );
  XNOR U10590 ( .A(n10906), .B(n10907), .Z(n10895) );
  AND U10591 ( .A(n302), .B(n10908), .Z(n10907) );
  XOR U10592 ( .A(p_input[315]), .B(n10906), .Z(n10908) );
  XNOR U10593 ( .A(n10909), .B(n10910), .Z(n10906) );
  AND U10594 ( .A(n306), .B(n10911), .Z(n10910) );
  XOR U10595 ( .A(n10912), .B(n10913), .Z(n10904) );
  AND U10596 ( .A(n310), .B(n10903), .Z(n10913) );
  XNOR U10597 ( .A(n10914), .B(n10901), .Z(n10903) );
  XOR U10598 ( .A(n10915), .B(n10916), .Z(n10901) );
  AND U10599 ( .A(n333), .B(n10917), .Z(n10916) );
  IV U10600 ( .A(n10912), .Z(n10914) );
  XOR U10601 ( .A(n10918), .B(n10919), .Z(n10912) );
  AND U10602 ( .A(n317), .B(n10911), .Z(n10919) );
  XNOR U10603 ( .A(n10909), .B(n10918), .Z(n10911) );
  XNOR U10604 ( .A(n10920), .B(n10921), .Z(n10909) );
  AND U10605 ( .A(n321), .B(n10922), .Z(n10921) );
  XOR U10606 ( .A(p_input[347]), .B(n10920), .Z(n10922) );
  XNOR U10607 ( .A(n10923), .B(n10924), .Z(n10920) );
  AND U10608 ( .A(n325), .B(n10925), .Z(n10924) );
  XOR U10609 ( .A(n10926), .B(n10927), .Z(n10918) );
  AND U10610 ( .A(n329), .B(n10917), .Z(n10927) );
  XNOR U10611 ( .A(n10928), .B(n10915), .Z(n10917) );
  XOR U10612 ( .A(n10929), .B(n10930), .Z(n10915) );
  AND U10613 ( .A(n352), .B(n10931), .Z(n10930) );
  IV U10614 ( .A(n10926), .Z(n10928) );
  XOR U10615 ( .A(n10932), .B(n10933), .Z(n10926) );
  AND U10616 ( .A(n336), .B(n10925), .Z(n10933) );
  XNOR U10617 ( .A(n10923), .B(n10932), .Z(n10925) );
  XNOR U10618 ( .A(n10934), .B(n10935), .Z(n10923) );
  AND U10619 ( .A(n340), .B(n10936), .Z(n10935) );
  XOR U10620 ( .A(p_input[379]), .B(n10934), .Z(n10936) );
  XNOR U10621 ( .A(n10937), .B(n10938), .Z(n10934) );
  AND U10622 ( .A(n344), .B(n10939), .Z(n10938) );
  XOR U10623 ( .A(n10940), .B(n10941), .Z(n10932) );
  AND U10624 ( .A(n348), .B(n10931), .Z(n10941) );
  XNOR U10625 ( .A(n10942), .B(n10929), .Z(n10931) );
  XOR U10626 ( .A(n10943), .B(n10944), .Z(n10929) );
  AND U10627 ( .A(n371), .B(n10945), .Z(n10944) );
  IV U10628 ( .A(n10940), .Z(n10942) );
  XOR U10629 ( .A(n10946), .B(n10947), .Z(n10940) );
  AND U10630 ( .A(n355), .B(n10939), .Z(n10947) );
  XNOR U10631 ( .A(n10937), .B(n10946), .Z(n10939) );
  XNOR U10632 ( .A(n10948), .B(n10949), .Z(n10937) );
  AND U10633 ( .A(n359), .B(n10950), .Z(n10949) );
  XOR U10634 ( .A(p_input[411]), .B(n10948), .Z(n10950) );
  XNOR U10635 ( .A(n10951), .B(n10952), .Z(n10948) );
  AND U10636 ( .A(n363), .B(n10953), .Z(n10952) );
  XOR U10637 ( .A(n10954), .B(n10955), .Z(n10946) );
  AND U10638 ( .A(n367), .B(n10945), .Z(n10955) );
  XNOR U10639 ( .A(n10956), .B(n10943), .Z(n10945) );
  XOR U10640 ( .A(n10957), .B(n10958), .Z(n10943) );
  AND U10641 ( .A(n390), .B(n10959), .Z(n10958) );
  IV U10642 ( .A(n10954), .Z(n10956) );
  XOR U10643 ( .A(n10960), .B(n10961), .Z(n10954) );
  AND U10644 ( .A(n374), .B(n10953), .Z(n10961) );
  XNOR U10645 ( .A(n10951), .B(n10960), .Z(n10953) );
  XNOR U10646 ( .A(n10962), .B(n10963), .Z(n10951) );
  AND U10647 ( .A(n378), .B(n10964), .Z(n10963) );
  XOR U10648 ( .A(p_input[443]), .B(n10962), .Z(n10964) );
  XNOR U10649 ( .A(n10965), .B(n10966), .Z(n10962) );
  AND U10650 ( .A(n382), .B(n10967), .Z(n10966) );
  XOR U10651 ( .A(n10968), .B(n10969), .Z(n10960) );
  AND U10652 ( .A(n386), .B(n10959), .Z(n10969) );
  XNOR U10653 ( .A(n10970), .B(n10957), .Z(n10959) );
  XOR U10654 ( .A(n10971), .B(n10972), .Z(n10957) );
  AND U10655 ( .A(n409), .B(n10973), .Z(n10972) );
  IV U10656 ( .A(n10968), .Z(n10970) );
  XOR U10657 ( .A(n10974), .B(n10975), .Z(n10968) );
  AND U10658 ( .A(n393), .B(n10967), .Z(n10975) );
  XNOR U10659 ( .A(n10965), .B(n10974), .Z(n10967) );
  XNOR U10660 ( .A(n10976), .B(n10977), .Z(n10965) );
  AND U10661 ( .A(n397), .B(n10978), .Z(n10977) );
  XOR U10662 ( .A(p_input[475]), .B(n10976), .Z(n10978) );
  XNOR U10663 ( .A(n10979), .B(n10980), .Z(n10976) );
  AND U10664 ( .A(n401), .B(n10981), .Z(n10980) );
  XOR U10665 ( .A(n10982), .B(n10983), .Z(n10974) );
  AND U10666 ( .A(n405), .B(n10973), .Z(n10983) );
  XNOR U10667 ( .A(n10984), .B(n10971), .Z(n10973) );
  XOR U10668 ( .A(n10985), .B(n10986), .Z(n10971) );
  AND U10669 ( .A(n428), .B(n10987), .Z(n10986) );
  IV U10670 ( .A(n10982), .Z(n10984) );
  XOR U10671 ( .A(n10988), .B(n10989), .Z(n10982) );
  AND U10672 ( .A(n412), .B(n10981), .Z(n10989) );
  XNOR U10673 ( .A(n10979), .B(n10988), .Z(n10981) );
  XNOR U10674 ( .A(n10990), .B(n10991), .Z(n10979) );
  AND U10675 ( .A(n416), .B(n10992), .Z(n10991) );
  XOR U10676 ( .A(p_input[507]), .B(n10990), .Z(n10992) );
  XNOR U10677 ( .A(n10993), .B(n10994), .Z(n10990) );
  AND U10678 ( .A(n420), .B(n10995), .Z(n10994) );
  XOR U10679 ( .A(n10996), .B(n10997), .Z(n10988) );
  AND U10680 ( .A(n424), .B(n10987), .Z(n10997) );
  XNOR U10681 ( .A(n10998), .B(n10985), .Z(n10987) );
  XOR U10682 ( .A(n10999), .B(n11000), .Z(n10985) );
  AND U10683 ( .A(n447), .B(n11001), .Z(n11000) );
  IV U10684 ( .A(n10996), .Z(n10998) );
  XOR U10685 ( .A(n11002), .B(n11003), .Z(n10996) );
  AND U10686 ( .A(n431), .B(n10995), .Z(n11003) );
  XNOR U10687 ( .A(n10993), .B(n11002), .Z(n10995) );
  XNOR U10688 ( .A(n11004), .B(n11005), .Z(n10993) );
  AND U10689 ( .A(n435), .B(n11006), .Z(n11005) );
  XOR U10690 ( .A(p_input[539]), .B(n11004), .Z(n11006) );
  XNOR U10691 ( .A(n11007), .B(n11008), .Z(n11004) );
  AND U10692 ( .A(n439), .B(n11009), .Z(n11008) );
  XOR U10693 ( .A(n11010), .B(n11011), .Z(n11002) );
  AND U10694 ( .A(n443), .B(n11001), .Z(n11011) );
  XNOR U10695 ( .A(n11012), .B(n10999), .Z(n11001) );
  XOR U10696 ( .A(n11013), .B(n11014), .Z(n10999) );
  AND U10697 ( .A(n466), .B(n11015), .Z(n11014) );
  IV U10698 ( .A(n11010), .Z(n11012) );
  XOR U10699 ( .A(n11016), .B(n11017), .Z(n11010) );
  AND U10700 ( .A(n450), .B(n11009), .Z(n11017) );
  XNOR U10701 ( .A(n11007), .B(n11016), .Z(n11009) );
  XNOR U10702 ( .A(n11018), .B(n11019), .Z(n11007) );
  AND U10703 ( .A(n454), .B(n11020), .Z(n11019) );
  XOR U10704 ( .A(p_input[571]), .B(n11018), .Z(n11020) );
  XNOR U10705 ( .A(n11021), .B(n11022), .Z(n11018) );
  AND U10706 ( .A(n458), .B(n11023), .Z(n11022) );
  XOR U10707 ( .A(n11024), .B(n11025), .Z(n11016) );
  AND U10708 ( .A(n462), .B(n11015), .Z(n11025) );
  XNOR U10709 ( .A(n11026), .B(n11013), .Z(n11015) );
  XOR U10710 ( .A(n11027), .B(n11028), .Z(n11013) );
  AND U10711 ( .A(n485), .B(n11029), .Z(n11028) );
  IV U10712 ( .A(n11024), .Z(n11026) );
  XOR U10713 ( .A(n11030), .B(n11031), .Z(n11024) );
  AND U10714 ( .A(n469), .B(n11023), .Z(n11031) );
  XNOR U10715 ( .A(n11021), .B(n11030), .Z(n11023) );
  XNOR U10716 ( .A(n11032), .B(n11033), .Z(n11021) );
  AND U10717 ( .A(n473), .B(n11034), .Z(n11033) );
  XOR U10718 ( .A(p_input[603]), .B(n11032), .Z(n11034) );
  XNOR U10719 ( .A(n11035), .B(n11036), .Z(n11032) );
  AND U10720 ( .A(n477), .B(n11037), .Z(n11036) );
  XOR U10721 ( .A(n11038), .B(n11039), .Z(n11030) );
  AND U10722 ( .A(n481), .B(n11029), .Z(n11039) );
  XNOR U10723 ( .A(n11040), .B(n11027), .Z(n11029) );
  XOR U10724 ( .A(n11041), .B(n11042), .Z(n11027) );
  AND U10725 ( .A(n504), .B(n11043), .Z(n11042) );
  IV U10726 ( .A(n11038), .Z(n11040) );
  XOR U10727 ( .A(n11044), .B(n11045), .Z(n11038) );
  AND U10728 ( .A(n488), .B(n11037), .Z(n11045) );
  XNOR U10729 ( .A(n11035), .B(n11044), .Z(n11037) );
  XNOR U10730 ( .A(n11046), .B(n11047), .Z(n11035) );
  AND U10731 ( .A(n492), .B(n11048), .Z(n11047) );
  XOR U10732 ( .A(p_input[635]), .B(n11046), .Z(n11048) );
  XNOR U10733 ( .A(n11049), .B(n11050), .Z(n11046) );
  AND U10734 ( .A(n496), .B(n11051), .Z(n11050) );
  XOR U10735 ( .A(n11052), .B(n11053), .Z(n11044) );
  AND U10736 ( .A(n500), .B(n11043), .Z(n11053) );
  XNOR U10737 ( .A(n11054), .B(n11041), .Z(n11043) );
  XOR U10738 ( .A(n11055), .B(n11056), .Z(n11041) );
  AND U10739 ( .A(n523), .B(n11057), .Z(n11056) );
  IV U10740 ( .A(n11052), .Z(n11054) );
  XOR U10741 ( .A(n11058), .B(n11059), .Z(n11052) );
  AND U10742 ( .A(n507), .B(n11051), .Z(n11059) );
  XNOR U10743 ( .A(n11049), .B(n11058), .Z(n11051) );
  XNOR U10744 ( .A(n11060), .B(n11061), .Z(n11049) );
  AND U10745 ( .A(n511), .B(n11062), .Z(n11061) );
  XOR U10746 ( .A(p_input[667]), .B(n11060), .Z(n11062) );
  XNOR U10747 ( .A(n11063), .B(n11064), .Z(n11060) );
  AND U10748 ( .A(n515), .B(n11065), .Z(n11064) );
  XOR U10749 ( .A(n11066), .B(n11067), .Z(n11058) );
  AND U10750 ( .A(n519), .B(n11057), .Z(n11067) );
  XNOR U10751 ( .A(n11068), .B(n11055), .Z(n11057) );
  XOR U10752 ( .A(n11069), .B(n11070), .Z(n11055) );
  AND U10753 ( .A(n542), .B(n11071), .Z(n11070) );
  IV U10754 ( .A(n11066), .Z(n11068) );
  XOR U10755 ( .A(n11072), .B(n11073), .Z(n11066) );
  AND U10756 ( .A(n526), .B(n11065), .Z(n11073) );
  XNOR U10757 ( .A(n11063), .B(n11072), .Z(n11065) );
  XNOR U10758 ( .A(n11074), .B(n11075), .Z(n11063) );
  AND U10759 ( .A(n530), .B(n11076), .Z(n11075) );
  XOR U10760 ( .A(p_input[699]), .B(n11074), .Z(n11076) );
  XNOR U10761 ( .A(n11077), .B(n11078), .Z(n11074) );
  AND U10762 ( .A(n534), .B(n11079), .Z(n11078) );
  XOR U10763 ( .A(n11080), .B(n11081), .Z(n11072) );
  AND U10764 ( .A(n538), .B(n11071), .Z(n11081) );
  XNOR U10765 ( .A(n11082), .B(n11069), .Z(n11071) );
  XOR U10766 ( .A(n11083), .B(n11084), .Z(n11069) );
  AND U10767 ( .A(n561), .B(n11085), .Z(n11084) );
  IV U10768 ( .A(n11080), .Z(n11082) );
  XOR U10769 ( .A(n11086), .B(n11087), .Z(n11080) );
  AND U10770 ( .A(n545), .B(n11079), .Z(n11087) );
  XNOR U10771 ( .A(n11077), .B(n11086), .Z(n11079) );
  XNOR U10772 ( .A(n11088), .B(n11089), .Z(n11077) );
  AND U10773 ( .A(n549), .B(n11090), .Z(n11089) );
  XOR U10774 ( .A(p_input[731]), .B(n11088), .Z(n11090) );
  XNOR U10775 ( .A(n11091), .B(n11092), .Z(n11088) );
  AND U10776 ( .A(n553), .B(n11093), .Z(n11092) );
  XOR U10777 ( .A(n11094), .B(n11095), .Z(n11086) );
  AND U10778 ( .A(n557), .B(n11085), .Z(n11095) );
  XNOR U10779 ( .A(n11096), .B(n11083), .Z(n11085) );
  XOR U10780 ( .A(n11097), .B(n11098), .Z(n11083) );
  AND U10781 ( .A(n580), .B(n11099), .Z(n11098) );
  IV U10782 ( .A(n11094), .Z(n11096) );
  XOR U10783 ( .A(n11100), .B(n11101), .Z(n11094) );
  AND U10784 ( .A(n564), .B(n11093), .Z(n11101) );
  XNOR U10785 ( .A(n11091), .B(n11100), .Z(n11093) );
  XNOR U10786 ( .A(n11102), .B(n11103), .Z(n11091) );
  AND U10787 ( .A(n568), .B(n11104), .Z(n11103) );
  XOR U10788 ( .A(p_input[763]), .B(n11102), .Z(n11104) );
  XNOR U10789 ( .A(n11105), .B(n11106), .Z(n11102) );
  AND U10790 ( .A(n572), .B(n11107), .Z(n11106) );
  XOR U10791 ( .A(n11108), .B(n11109), .Z(n11100) );
  AND U10792 ( .A(n576), .B(n11099), .Z(n11109) );
  XNOR U10793 ( .A(n11110), .B(n11097), .Z(n11099) );
  XOR U10794 ( .A(n11111), .B(n11112), .Z(n11097) );
  AND U10795 ( .A(n599), .B(n11113), .Z(n11112) );
  IV U10796 ( .A(n11108), .Z(n11110) );
  XOR U10797 ( .A(n11114), .B(n11115), .Z(n11108) );
  AND U10798 ( .A(n583), .B(n11107), .Z(n11115) );
  XNOR U10799 ( .A(n11105), .B(n11114), .Z(n11107) );
  XNOR U10800 ( .A(n11116), .B(n11117), .Z(n11105) );
  AND U10801 ( .A(n587), .B(n11118), .Z(n11117) );
  XOR U10802 ( .A(p_input[795]), .B(n11116), .Z(n11118) );
  XNOR U10803 ( .A(n11119), .B(n11120), .Z(n11116) );
  AND U10804 ( .A(n591), .B(n11121), .Z(n11120) );
  XOR U10805 ( .A(n11122), .B(n11123), .Z(n11114) );
  AND U10806 ( .A(n595), .B(n11113), .Z(n11123) );
  XNOR U10807 ( .A(n11124), .B(n11111), .Z(n11113) );
  XOR U10808 ( .A(n11125), .B(n11126), .Z(n11111) );
  AND U10809 ( .A(n618), .B(n11127), .Z(n11126) );
  IV U10810 ( .A(n11122), .Z(n11124) );
  XOR U10811 ( .A(n11128), .B(n11129), .Z(n11122) );
  AND U10812 ( .A(n602), .B(n11121), .Z(n11129) );
  XNOR U10813 ( .A(n11119), .B(n11128), .Z(n11121) );
  XNOR U10814 ( .A(n11130), .B(n11131), .Z(n11119) );
  AND U10815 ( .A(n606), .B(n11132), .Z(n11131) );
  XOR U10816 ( .A(p_input[827]), .B(n11130), .Z(n11132) );
  XNOR U10817 ( .A(n11133), .B(n11134), .Z(n11130) );
  AND U10818 ( .A(n610), .B(n11135), .Z(n11134) );
  XOR U10819 ( .A(n11136), .B(n11137), .Z(n11128) );
  AND U10820 ( .A(n614), .B(n11127), .Z(n11137) );
  XNOR U10821 ( .A(n11138), .B(n11125), .Z(n11127) );
  XOR U10822 ( .A(n11139), .B(n11140), .Z(n11125) );
  AND U10823 ( .A(n637), .B(n11141), .Z(n11140) );
  IV U10824 ( .A(n11136), .Z(n11138) );
  XOR U10825 ( .A(n11142), .B(n11143), .Z(n11136) );
  AND U10826 ( .A(n621), .B(n11135), .Z(n11143) );
  XNOR U10827 ( .A(n11133), .B(n11142), .Z(n11135) );
  XNOR U10828 ( .A(n11144), .B(n11145), .Z(n11133) );
  AND U10829 ( .A(n625), .B(n11146), .Z(n11145) );
  XOR U10830 ( .A(p_input[859]), .B(n11144), .Z(n11146) );
  XNOR U10831 ( .A(n11147), .B(n11148), .Z(n11144) );
  AND U10832 ( .A(n629), .B(n11149), .Z(n11148) );
  XOR U10833 ( .A(n11150), .B(n11151), .Z(n11142) );
  AND U10834 ( .A(n633), .B(n11141), .Z(n11151) );
  XNOR U10835 ( .A(n11152), .B(n11139), .Z(n11141) );
  XOR U10836 ( .A(n11153), .B(n11154), .Z(n11139) );
  AND U10837 ( .A(n656), .B(n11155), .Z(n11154) );
  IV U10838 ( .A(n11150), .Z(n11152) );
  XOR U10839 ( .A(n11156), .B(n11157), .Z(n11150) );
  AND U10840 ( .A(n640), .B(n11149), .Z(n11157) );
  XNOR U10841 ( .A(n11147), .B(n11156), .Z(n11149) );
  XNOR U10842 ( .A(n11158), .B(n11159), .Z(n11147) );
  AND U10843 ( .A(n644), .B(n11160), .Z(n11159) );
  XOR U10844 ( .A(p_input[891]), .B(n11158), .Z(n11160) );
  XNOR U10845 ( .A(n11161), .B(n11162), .Z(n11158) );
  AND U10846 ( .A(n648), .B(n11163), .Z(n11162) );
  XOR U10847 ( .A(n11164), .B(n11165), .Z(n11156) );
  AND U10848 ( .A(n652), .B(n11155), .Z(n11165) );
  XNOR U10849 ( .A(n11166), .B(n11153), .Z(n11155) );
  XOR U10850 ( .A(n11167), .B(n11168), .Z(n11153) );
  AND U10851 ( .A(n675), .B(n11169), .Z(n11168) );
  IV U10852 ( .A(n11164), .Z(n11166) );
  XOR U10853 ( .A(n11170), .B(n11171), .Z(n11164) );
  AND U10854 ( .A(n659), .B(n11163), .Z(n11171) );
  XNOR U10855 ( .A(n11161), .B(n11170), .Z(n11163) );
  XNOR U10856 ( .A(n11172), .B(n11173), .Z(n11161) );
  AND U10857 ( .A(n663), .B(n11174), .Z(n11173) );
  XOR U10858 ( .A(p_input[923]), .B(n11172), .Z(n11174) );
  XNOR U10859 ( .A(n11175), .B(n11176), .Z(n11172) );
  AND U10860 ( .A(n667), .B(n11177), .Z(n11176) );
  XOR U10861 ( .A(n11178), .B(n11179), .Z(n11170) );
  AND U10862 ( .A(n671), .B(n11169), .Z(n11179) );
  XNOR U10863 ( .A(n11180), .B(n11167), .Z(n11169) );
  XOR U10864 ( .A(n11181), .B(n11182), .Z(n11167) );
  AND U10865 ( .A(n694), .B(n11183), .Z(n11182) );
  IV U10866 ( .A(n11178), .Z(n11180) );
  XOR U10867 ( .A(n11184), .B(n11185), .Z(n11178) );
  AND U10868 ( .A(n678), .B(n11177), .Z(n11185) );
  XNOR U10869 ( .A(n11175), .B(n11184), .Z(n11177) );
  XNOR U10870 ( .A(n11186), .B(n11187), .Z(n11175) );
  AND U10871 ( .A(n682), .B(n11188), .Z(n11187) );
  XOR U10872 ( .A(p_input[955]), .B(n11186), .Z(n11188) );
  XNOR U10873 ( .A(n11189), .B(n11190), .Z(n11186) );
  AND U10874 ( .A(n686), .B(n11191), .Z(n11190) );
  XOR U10875 ( .A(n11192), .B(n11193), .Z(n11184) );
  AND U10876 ( .A(n690), .B(n11183), .Z(n11193) );
  XNOR U10877 ( .A(n11194), .B(n11181), .Z(n11183) );
  XOR U10878 ( .A(n11195), .B(n11196), .Z(n11181) );
  AND U10879 ( .A(n713), .B(n11197), .Z(n11196) );
  IV U10880 ( .A(n11192), .Z(n11194) );
  XOR U10881 ( .A(n11198), .B(n11199), .Z(n11192) );
  AND U10882 ( .A(n697), .B(n11191), .Z(n11199) );
  XNOR U10883 ( .A(n11189), .B(n11198), .Z(n11191) );
  XNOR U10884 ( .A(n11200), .B(n11201), .Z(n11189) );
  AND U10885 ( .A(n701), .B(n11202), .Z(n11201) );
  XOR U10886 ( .A(p_input[987]), .B(n11200), .Z(n11202) );
  XNOR U10887 ( .A(n11203), .B(n11204), .Z(n11200) );
  AND U10888 ( .A(n705), .B(n11205), .Z(n11204) );
  XOR U10889 ( .A(n11206), .B(n11207), .Z(n11198) );
  AND U10890 ( .A(n709), .B(n11197), .Z(n11207) );
  XNOR U10891 ( .A(n11208), .B(n11195), .Z(n11197) );
  XOR U10892 ( .A(n11209), .B(n11210), .Z(n11195) );
  AND U10893 ( .A(n732), .B(n11211), .Z(n11210) );
  IV U10894 ( .A(n11206), .Z(n11208) );
  XOR U10895 ( .A(n11212), .B(n11213), .Z(n11206) );
  AND U10896 ( .A(n716), .B(n11205), .Z(n11213) );
  XNOR U10897 ( .A(n11203), .B(n11212), .Z(n11205) );
  XNOR U10898 ( .A(n11214), .B(n11215), .Z(n11203) );
  AND U10899 ( .A(n720), .B(n11216), .Z(n11215) );
  XOR U10900 ( .A(p_input[1019]), .B(n11214), .Z(n11216) );
  XNOR U10901 ( .A(n11217), .B(n11218), .Z(n11214) );
  AND U10902 ( .A(n724), .B(n11219), .Z(n11218) );
  XOR U10903 ( .A(n11220), .B(n11221), .Z(n11212) );
  AND U10904 ( .A(n728), .B(n11211), .Z(n11221) );
  XNOR U10905 ( .A(n11222), .B(n11209), .Z(n11211) );
  XOR U10906 ( .A(n11223), .B(n11224), .Z(n11209) );
  AND U10907 ( .A(n751), .B(n11225), .Z(n11224) );
  IV U10908 ( .A(n11220), .Z(n11222) );
  XOR U10909 ( .A(n11226), .B(n11227), .Z(n11220) );
  AND U10910 ( .A(n735), .B(n11219), .Z(n11227) );
  XNOR U10911 ( .A(n11217), .B(n11226), .Z(n11219) );
  XNOR U10912 ( .A(n11228), .B(n11229), .Z(n11217) );
  AND U10913 ( .A(n739), .B(n11230), .Z(n11229) );
  XOR U10914 ( .A(p_input[1051]), .B(n11228), .Z(n11230) );
  XNOR U10915 ( .A(n11231), .B(n11232), .Z(n11228) );
  AND U10916 ( .A(n743), .B(n11233), .Z(n11232) );
  XOR U10917 ( .A(n11234), .B(n11235), .Z(n11226) );
  AND U10918 ( .A(n747), .B(n11225), .Z(n11235) );
  XNOR U10919 ( .A(n11236), .B(n11223), .Z(n11225) );
  XOR U10920 ( .A(n11237), .B(n11238), .Z(n11223) );
  AND U10921 ( .A(n770), .B(n11239), .Z(n11238) );
  IV U10922 ( .A(n11234), .Z(n11236) );
  XOR U10923 ( .A(n11240), .B(n11241), .Z(n11234) );
  AND U10924 ( .A(n754), .B(n11233), .Z(n11241) );
  XNOR U10925 ( .A(n11231), .B(n11240), .Z(n11233) );
  XNOR U10926 ( .A(n11242), .B(n11243), .Z(n11231) );
  AND U10927 ( .A(n758), .B(n11244), .Z(n11243) );
  XOR U10928 ( .A(p_input[1083]), .B(n11242), .Z(n11244) );
  XNOR U10929 ( .A(n11245), .B(n11246), .Z(n11242) );
  AND U10930 ( .A(n762), .B(n11247), .Z(n11246) );
  XOR U10931 ( .A(n11248), .B(n11249), .Z(n11240) );
  AND U10932 ( .A(n766), .B(n11239), .Z(n11249) );
  XNOR U10933 ( .A(n11250), .B(n11237), .Z(n11239) );
  XOR U10934 ( .A(n11251), .B(n11252), .Z(n11237) );
  AND U10935 ( .A(n789), .B(n11253), .Z(n11252) );
  IV U10936 ( .A(n11248), .Z(n11250) );
  XOR U10937 ( .A(n11254), .B(n11255), .Z(n11248) );
  AND U10938 ( .A(n773), .B(n11247), .Z(n11255) );
  XNOR U10939 ( .A(n11245), .B(n11254), .Z(n11247) );
  XNOR U10940 ( .A(n11256), .B(n11257), .Z(n11245) );
  AND U10941 ( .A(n777), .B(n11258), .Z(n11257) );
  XOR U10942 ( .A(p_input[1115]), .B(n11256), .Z(n11258) );
  XNOR U10943 ( .A(n11259), .B(n11260), .Z(n11256) );
  AND U10944 ( .A(n781), .B(n11261), .Z(n11260) );
  XOR U10945 ( .A(n11262), .B(n11263), .Z(n11254) );
  AND U10946 ( .A(n785), .B(n11253), .Z(n11263) );
  XNOR U10947 ( .A(n11264), .B(n11251), .Z(n11253) );
  XOR U10948 ( .A(n11265), .B(n11266), .Z(n11251) );
  AND U10949 ( .A(n808), .B(n11267), .Z(n11266) );
  IV U10950 ( .A(n11262), .Z(n11264) );
  XOR U10951 ( .A(n11268), .B(n11269), .Z(n11262) );
  AND U10952 ( .A(n792), .B(n11261), .Z(n11269) );
  XNOR U10953 ( .A(n11259), .B(n11268), .Z(n11261) );
  XNOR U10954 ( .A(n11270), .B(n11271), .Z(n11259) );
  AND U10955 ( .A(n796), .B(n11272), .Z(n11271) );
  XOR U10956 ( .A(p_input[1147]), .B(n11270), .Z(n11272) );
  XNOR U10957 ( .A(n11273), .B(n11274), .Z(n11270) );
  AND U10958 ( .A(n800), .B(n11275), .Z(n11274) );
  XOR U10959 ( .A(n11276), .B(n11277), .Z(n11268) );
  AND U10960 ( .A(n804), .B(n11267), .Z(n11277) );
  XNOR U10961 ( .A(n11278), .B(n11265), .Z(n11267) );
  XOR U10962 ( .A(n11279), .B(n11280), .Z(n11265) );
  AND U10963 ( .A(n827), .B(n11281), .Z(n11280) );
  IV U10964 ( .A(n11276), .Z(n11278) );
  XOR U10965 ( .A(n11282), .B(n11283), .Z(n11276) );
  AND U10966 ( .A(n811), .B(n11275), .Z(n11283) );
  XNOR U10967 ( .A(n11273), .B(n11282), .Z(n11275) );
  XNOR U10968 ( .A(n11284), .B(n11285), .Z(n11273) );
  AND U10969 ( .A(n815), .B(n11286), .Z(n11285) );
  XOR U10970 ( .A(p_input[1179]), .B(n11284), .Z(n11286) );
  XNOR U10971 ( .A(n11287), .B(n11288), .Z(n11284) );
  AND U10972 ( .A(n819), .B(n11289), .Z(n11288) );
  XOR U10973 ( .A(n11290), .B(n11291), .Z(n11282) );
  AND U10974 ( .A(n823), .B(n11281), .Z(n11291) );
  XNOR U10975 ( .A(n11292), .B(n11279), .Z(n11281) );
  XOR U10976 ( .A(n11293), .B(n11294), .Z(n11279) );
  AND U10977 ( .A(n846), .B(n11295), .Z(n11294) );
  IV U10978 ( .A(n11290), .Z(n11292) );
  XOR U10979 ( .A(n11296), .B(n11297), .Z(n11290) );
  AND U10980 ( .A(n830), .B(n11289), .Z(n11297) );
  XNOR U10981 ( .A(n11287), .B(n11296), .Z(n11289) );
  XNOR U10982 ( .A(n11298), .B(n11299), .Z(n11287) );
  AND U10983 ( .A(n834), .B(n11300), .Z(n11299) );
  XOR U10984 ( .A(p_input[1211]), .B(n11298), .Z(n11300) );
  XNOR U10985 ( .A(n11301), .B(n11302), .Z(n11298) );
  AND U10986 ( .A(n838), .B(n11303), .Z(n11302) );
  XOR U10987 ( .A(n11304), .B(n11305), .Z(n11296) );
  AND U10988 ( .A(n842), .B(n11295), .Z(n11305) );
  XNOR U10989 ( .A(n11306), .B(n11293), .Z(n11295) );
  XOR U10990 ( .A(n11307), .B(n11308), .Z(n11293) );
  AND U10991 ( .A(n865), .B(n11309), .Z(n11308) );
  IV U10992 ( .A(n11304), .Z(n11306) );
  XOR U10993 ( .A(n11310), .B(n11311), .Z(n11304) );
  AND U10994 ( .A(n849), .B(n11303), .Z(n11311) );
  XNOR U10995 ( .A(n11301), .B(n11310), .Z(n11303) );
  XNOR U10996 ( .A(n11312), .B(n11313), .Z(n11301) );
  AND U10997 ( .A(n853), .B(n11314), .Z(n11313) );
  XOR U10998 ( .A(p_input[1243]), .B(n11312), .Z(n11314) );
  XNOR U10999 ( .A(n11315), .B(n11316), .Z(n11312) );
  AND U11000 ( .A(n857), .B(n11317), .Z(n11316) );
  XOR U11001 ( .A(n11318), .B(n11319), .Z(n11310) );
  AND U11002 ( .A(n861), .B(n11309), .Z(n11319) );
  XNOR U11003 ( .A(n11320), .B(n11307), .Z(n11309) );
  XOR U11004 ( .A(n11321), .B(n11322), .Z(n11307) );
  AND U11005 ( .A(n884), .B(n11323), .Z(n11322) );
  IV U11006 ( .A(n11318), .Z(n11320) );
  XOR U11007 ( .A(n11324), .B(n11325), .Z(n11318) );
  AND U11008 ( .A(n868), .B(n11317), .Z(n11325) );
  XNOR U11009 ( .A(n11315), .B(n11324), .Z(n11317) );
  XNOR U11010 ( .A(n11326), .B(n11327), .Z(n11315) );
  AND U11011 ( .A(n872), .B(n11328), .Z(n11327) );
  XOR U11012 ( .A(p_input[1275]), .B(n11326), .Z(n11328) );
  XNOR U11013 ( .A(n11329), .B(n11330), .Z(n11326) );
  AND U11014 ( .A(n876), .B(n11331), .Z(n11330) );
  XOR U11015 ( .A(n11332), .B(n11333), .Z(n11324) );
  AND U11016 ( .A(n880), .B(n11323), .Z(n11333) );
  XNOR U11017 ( .A(n11334), .B(n11321), .Z(n11323) );
  XOR U11018 ( .A(n11335), .B(n11336), .Z(n11321) );
  AND U11019 ( .A(n903), .B(n11337), .Z(n11336) );
  IV U11020 ( .A(n11332), .Z(n11334) );
  XOR U11021 ( .A(n11338), .B(n11339), .Z(n11332) );
  AND U11022 ( .A(n887), .B(n11331), .Z(n11339) );
  XNOR U11023 ( .A(n11329), .B(n11338), .Z(n11331) );
  XNOR U11024 ( .A(n11340), .B(n11341), .Z(n11329) );
  AND U11025 ( .A(n891), .B(n11342), .Z(n11341) );
  XOR U11026 ( .A(p_input[1307]), .B(n11340), .Z(n11342) );
  XNOR U11027 ( .A(n11343), .B(n11344), .Z(n11340) );
  AND U11028 ( .A(n895), .B(n11345), .Z(n11344) );
  XOR U11029 ( .A(n11346), .B(n11347), .Z(n11338) );
  AND U11030 ( .A(n899), .B(n11337), .Z(n11347) );
  XNOR U11031 ( .A(n11348), .B(n11335), .Z(n11337) );
  XOR U11032 ( .A(n11349), .B(n11350), .Z(n11335) );
  AND U11033 ( .A(n922), .B(n11351), .Z(n11350) );
  IV U11034 ( .A(n11346), .Z(n11348) );
  XOR U11035 ( .A(n11352), .B(n11353), .Z(n11346) );
  AND U11036 ( .A(n906), .B(n11345), .Z(n11353) );
  XNOR U11037 ( .A(n11343), .B(n11352), .Z(n11345) );
  XNOR U11038 ( .A(n11354), .B(n11355), .Z(n11343) );
  AND U11039 ( .A(n910), .B(n11356), .Z(n11355) );
  XOR U11040 ( .A(p_input[1339]), .B(n11354), .Z(n11356) );
  XNOR U11041 ( .A(n11357), .B(n11358), .Z(n11354) );
  AND U11042 ( .A(n914), .B(n11359), .Z(n11358) );
  XOR U11043 ( .A(n11360), .B(n11361), .Z(n11352) );
  AND U11044 ( .A(n918), .B(n11351), .Z(n11361) );
  XNOR U11045 ( .A(n11362), .B(n11349), .Z(n11351) );
  XOR U11046 ( .A(n11363), .B(n11364), .Z(n11349) );
  AND U11047 ( .A(n941), .B(n11365), .Z(n11364) );
  IV U11048 ( .A(n11360), .Z(n11362) );
  XOR U11049 ( .A(n11366), .B(n11367), .Z(n11360) );
  AND U11050 ( .A(n925), .B(n11359), .Z(n11367) );
  XNOR U11051 ( .A(n11357), .B(n11366), .Z(n11359) );
  XNOR U11052 ( .A(n11368), .B(n11369), .Z(n11357) );
  AND U11053 ( .A(n929), .B(n11370), .Z(n11369) );
  XOR U11054 ( .A(p_input[1371]), .B(n11368), .Z(n11370) );
  XNOR U11055 ( .A(n11371), .B(n11372), .Z(n11368) );
  AND U11056 ( .A(n933), .B(n11373), .Z(n11372) );
  XOR U11057 ( .A(n11374), .B(n11375), .Z(n11366) );
  AND U11058 ( .A(n937), .B(n11365), .Z(n11375) );
  XNOR U11059 ( .A(n11376), .B(n11363), .Z(n11365) );
  XOR U11060 ( .A(n11377), .B(n11378), .Z(n11363) );
  AND U11061 ( .A(n960), .B(n11379), .Z(n11378) );
  IV U11062 ( .A(n11374), .Z(n11376) );
  XOR U11063 ( .A(n11380), .B(n11381), .Z(n11374) );
  AND U11064 ( .A(n944), .B(n11373), .Z(n11381) );
  XNOR U11065 ( .A(n11371), .B(n11380), .Z(n11373) );
  XNOR U11066 ( .A(n11382), .B(n11383), .Z(n11371) );
  AND U11067 ( .A(n948), .B(n11384), .Z(n11383) );
  XOR U11068 ( .A(p_input[1403]), .B(n11382), .Z(n11384) );
  XNOR U11069 ( .A(n11385), .B(n11386), .Z(n11382) );
  AND U11070 ( .A(n952), .B(n11387), .Z(n11386) );
  XOR U11071 ( .A(n11388), .B(n11389), .Z(n11380) );
  AND U11072 ( .A(n956), .B(n11379), .Z(n11389) );
  XNOR U11073 ( .A(n11390), .B(n11377), .Z(n11379) );
  XOR U11074 ( .A(n11391), .B(n11392), .Z(n11377) );
  AND U11075 ( .A(n979), .B(n11393), .Z(n11392) );
  IV U11076 ( .A(n11388), .Z(n11390) );
  XOR U11077 ( .A(n11394), .B(n11395), .Z(n11388) );
  AND U11078 ( .A(n963), .B(n11387), .Z(n11395) );
  XNOR U11079 ( .A(n11385), .B(n11394), .Z(n11387) );
  XNOR U11080 ( .A(n11396), .B(n11397), .Z(n11385) );
  AND U11081 ( .A(n967), .B(n11398), .Z(n11397) );
  XOR U11082 ( .A(p_input[1435]), .B(n11396), .Z(n11398) );
  XNOR U11083 ( .A(n11399), .B(n11400), .Z(n11396) );
  AND U11084 ( .A(n971), .B(n11401), .Z(n11400) );
  XOR U11085 ( .A(n11402), .B(n11403), .Z(n11394) );
  AND U11086 ( .A(n975), .B(n11393), .Z(n11403) );
  XNOR U11087 ( .A(n11404), .B(n11391), .Z(n11393) );
  XOR U11088 ( .A(n11405), .B(n11406), .Z(n11391) );
  AND U11089 ( .A(n998), .B(n11407), .Z(n11406) );
  IV U11090 ( .A(n11402), .Z(n11404) );
  XOR U11091 ( .A(n11408), .B(n11409), .Z(n11402) );
  AND U11092 ( .A(n982), .B(n11401), .Z(n11409) );
  XNOR U11093 ( .A(n11399), .B(n11408), .Z(n11401) );
  XNOR U11094 ( .A(n11410), .B(n11411), .Z(n11399) );
  AND U11095 ( .A(n986), .B(n11412), .Z(n11411) );
  XOR U11096 ( .A(p_input[1467]), .B(n11410), .Z(n11412) );
  XNOR U11097 ( .A(n11413), .B(n11414), .Z(n11410) );
  AND U11098 ( .A(n990), .B(n11415), .Z(n11414) );
  XOR U11099 ( .A(n11416), .B(n11417), .Z(n11408) );
  AND U11100 ( .A(n994), .B(n11407), .Z(n11417) );
  XNOR U11101 ( .A(n11418), .B(n11405), .Z(n11407) );
  XOR U11102 ( .A(n11419), .B(n11420), .Z(n11405) );
  AND U11103 ( .A(n1017), .B(n11421), .Z(n11420) );
  IV U11104 ( .A(n11416), .Z(n11418) );
  XOR U11105 ( .A(n11422), .B(n11423), .Z(n11416) );
  AND U11106 ( .A(n1001), .B(n11415), .Z(n11423) );
  XNOR U11107 ( .A(n11413), .B(n11422), .Z(n11415) );
  XNOR U11108 ( .A(n11424), .B(n11425), .Z(n11413) );
  AND U11109 ( .A(n1005), .B(n11426), .Z(n11425) );
  XOR U11110 ( .A(p_input[1499]), .B(n11424), .Z(n11426) );
  XNOR U11111 ( .A(n11427), .B(n11428), .Z(n11424) );
  AND U11112 ( .A(n1009), .B(n11429), .Z(n11428) );
  XOR U11113 ( .A(n11430), .B(n11431), .Z(n11422) );
  AND U11114 ( .A(n1013), .B(n11421), .Z(n11431) );
  XNOR U11115 ( .A(n11432), .B(n11419), .Z(n11421) );
  XOR U11116 ( .A(n11433), .B(n11434), .Z(n11419) );
  AND U11117 ( .A(n1036), .B(n11435), .Z(n11434) );
  IV U11118 ( .A(n11430), .Z(n11432) );
  XOR U11119 ( .A(n11436), .B(n11437), .Z(n11430) );
  AND U11120 ( .A(n1020), .B(n11429), .Z(n11437) );
  XNOR U11121 ( .A(n11427), .B(n11436), .Z(n11429) );
  XNOR U11122 ( .A(n11438), .B(n11439), .Z(n11427) );
  AND U11123 ( .A(n1024), .B(n11440), .Z(n11439) );
  XOR U11124 ( .A(p_input[1531]), .B(n11438), .Z(n11440) );
  XNOR U11125 ( .A(n11441), .B(n11442), .Z(n11438) );
  AND U11126 ( .A(n1028), .B(n11443), .Z(n11442) );
  XOR U11127 ( .A(n11444), .B(n11445), .Z(n11436) );
  AND U11128 ( .A(n1032), .B(n11435), .Z(n11445) );
  XNOR U11129 ( .A(n11446), .B(n11433), .Z(n11435) );
  XOR U11130 ( .A(n11447), .B(n11448), .Z(n11433) );
  AND U11131 ( .A(n1055), .B(n11449), .Z(n11448) );
  IV U11132 ( .A(n11444), .Z(n11446) );
  XOR U11133 ( .A(n11450), .B(n11451), .Z(n11444) );
  AND U11134 ( .A(n1039), .B(n11443), .Z(n11451) );
  XNOR U11135 ( .A(n11441), .B(n11450), .Z(n11443) );
  XNOR U11136 ( .A(n11452), .B(n11453), .Z(n11441) );
  AND U11137 ( .A(n1043), .B(n11454), .Z(n11453) );
  XOR U11138 ( .A(p_input[1563]), .B(n11452), .Z(n11454) );
  XNOR U11139 ( .A(n11455), .B(n11456), .Z(n11452) );
  AND U11140 ( .A(n1047), .B(n11457), .Z(n11456) );
  XOR U11141 ( .A(n11458), .B(n11459), .Z(n11450) );
  AND U11142 ( .A(n1051), .B(n11449), .Z(n11459) );
  XNOR U11143 ( .A(n11460), .B(n11447), .Z(n11449) );
  XOR U11144 ( .A(n11461), .B(n11462), .Z(n11447) );
  AND U11145 ( .A(n1074), .B(n11463), .Z(n11462) );
  IV U11146 ( .A(n11458), .Z(n11460) );
  XOR U11147 ( .A(n11464), .B(n11465), .Z(n11458) );
  AND U11148 ( .A(n1058), .B(n11457), .Z(n11465) );
  XNOR U11149 ( .A(n11455), .B(n11464), .Z(n11457) );
  XNOR U11150 ( .A(n11466), .B(n11467), .Z(n11455) );
  AND U11151 ( .A(n1062), .B(n11468), .Z(n11467) );
  XOR U11152 ( .A(p_input[1595]), .B(n11466), .Z(n11468) );
  XNOR U11153 ( .A(n11469), .B(n11470), .Z(n11466) );
  AND U11154 ( .A(n1066), .B(n11471), .Z(n11470) );
  XOR U11155 ( .A(n11472), .B(n11473), .Z(n11464) );
  AND U11156 ( .A(n1070), .B(n11463), .Z(n11473) );
  XNOR U11157 ( .A(n11474), .B(n11461), .Z(n11463) );
  XOR U11158 ( .A(n11475), .B(n11476), .Z(n11461) );
  AND U11159 ( .A(n1093), .B(n11477), .Z(n11476) );
  IV U11160 ( .A(n11472), .Z(n11474) );
  XOR U11161 ( .A(n11478), .B(n11479), .Z(n11472) );
  AND U11162 ( .A(n1077), .B(n11471), .Z(n11479) );
  XNOR U11163 ( .A(n11469), .B(n11478), .Z(n11471) );
  XNOR U11164 ( .A(n11480), .B(n11481), .Z(n11469) );
  AND U11165 ( .A(n1081), .B(n11482), .Z(n11481) );
  XOR U11166 ( .A(p_input[1627]), .B(n11480), .Z(n11482) );
  XNOR U11167 ( .A(n11483), .B(n11484), .Z(n11480) );
  AND U11168 ( .A(n1085), .B(n11485), .Z(n11484) );
  XOR U11169 ( .A(n11486), .B(n11487), .Z(n11478) );
  AND U11170 ( .A(n1089), .B(n11477), .Z(n11487) );
  XNOR U11171 ( .A(n11488), .B(n11475), .Z(n11477) );
  XOR U11172 ( .A(n11489), .B(n11490), .Z(n11475) );
  AND U11173 ( .A(n1112), .B(n11491), .Z(n11490) );
  IV U11174 ( .A(n11486), .Z(n11488) );
  XOR U11175 ( .A(n11492), .B(n11493), .Z(n11486) );
  AND U11176 ( .A(n1096), .B(n11485), .Z(n11493) );
  XNOR U11177 ( .A(n11483), .B(n11492), .Z(n11485) );
  XNOR U11178 ( .A(n11494), .B(n11495), .Z(n11483) );
  AND U11179 ( .A(n1100), .B(n11496), .Z(n11495) );
  XOR U11180 ( .A(p_input[1659]), .B(n11494), .Z(n11496) );
  XNOR U11181 ( .A(n11497), .B(n11498), .Z(n11494) );
  AND U11182 ( .A(n1104), .B(n11499), .Z(n11498) );
  XOR U11183 ( .A(n11500), .B(n11501), .Z(n11492) );
  AND U11184 ( .A(n1108), .B(n11491), .Z(n11501) );
  XNOR U11185 ( .A(n11502), .B(n11489), .Z(n11491) );
  XOR U11186 ( .A(n11503), .B(n11504), .Z(n11489) );
  AND U11187 ( .A(n1131), .B(n11505), .Z(n11504) );
  IV U11188 ( .A(n11500), .Z(n11502) );
  XOR U11189 ( .A(n11506), .B(n11507), .Z(n11500) );
  AND U11190 ( .A(n1115), .B(n11499), .Z(n11507) );
  XNOR U11191 ( .A(n11497), .B(n11506), .Z(n11499) );
  XNOR U11192 ( .A(n11508), .B(n11509), .Z(n11497) );
  AND U11193 ( .A(n1119), .B(n11510), .Z(n11509) );
  XOR U11194 ( .A(p_input[1691]), .B(n11508), .Z(n11510) );
  XNOR U11195 ( .A(n11511), .B(n11512), .Z(n11508) );
  AND U11196 ( .A(n1123), .B(n11513), .Z(n11512) );
  XOR U11197 ( .A(n11514), .B(n11515), .Z(n11506) );
  AND U11198 ( .A(n1127), .B(n11505), .Z(n11515) );
  XNOR U11199 ( .A(n11516), .B(n11503), .Z(n11505) );
  XOR U11200 ( .A(n11517), .B(n11518), .Z(n11503) );
  AND U11201 ( .A(n1150), .B(n11519), .Z(n11518) );
  IV U11202 ( .A(n11514), .Z(n11516) );
  XOR U11203 ( .A(n11520), .B(n11521), .Z(n11514) );
  AND U11204 ( .A(n1134), .B(n11513), .Z(n11521) );
  XNOR U11205 ( .A(n11511), .B(n11520), .Z(n11513) );
  XNOR U11206 ( .A(n11522), .B(n11523), .Z(n11511) );
  AND U11207 ( .A(n1138), .B(n11524), .Z(n11523) );
  XOR U11208 ( .A(p_input[1723]), .B(n11522), .Z(n11524) );
  XNOR U11209 ( .A(n11525), .B(n11526), .Z(n11522) );
  AND U11210 ( .A(n1142), .B(n11527), .Z(n11526) );
  XOR U11211 ( .A(n11528), .B(n11529), .Z(n11520) );
  AND U11212 ( .A(n1146), .B(n11519), .Z(n11529) );
  XNOR U11213 ( .A(n11530), .B(n11517), .Z(n11519) );
  XOR U11214 ( .A(n11531), .B(n11532), .Z(n11517) );
  AND U11215 ( .A(n1169), .B(n11533), .Z(n11532) );
  IV U11216 ( .A(n11528), .Z(n11530) );
  XOR U11217 ( .A(n11534), .B(n11535), .Z(n11528) );
  AND U11218 ( .A(n1153), .B(n11527), .Z(n11535) );
  XNOR U11219 ( .A(n11525), .B(n11534), .Z(n11527) );
  XNOR U11220 ( .A(n11536), .B(n11537), .Z(n11525) );
  AND U11221 ( .A(n1157), .B(n11538), .Z(n11537) );
  XOR U11222 ( .A(p_input[1755]), .B(n11536), .Z(n11538) );
  XNOR U11223 ( .A(n11539), .B(n11540), .Z(n11536) );
  AND U11224 ( .A(n1161), .B(n11541), .Z(n11540) );
  XOR U11225 ( .A(n11542), .B(n11543), .Z(n11534) );
  AND U11226 ( .A(n1165), .B(n11533), .Z(n11543) );
  XNOR U11227 ( .A(n11544), .B(n11531), .Z(n11533) );
  XOR U11228 ( .A(n11545), .B(n11546), .Z(n11531) );
  AND U11229 ( .A(n1188), .B(n11547), .Z(n11546) );
  IV U11230 ( .A(n11542), .Z(n11544) );
  XOR U11231 ( .A(n11548), .B(n11549), .Z(n11542) );
  AND U11232 ( .A(n1172), .B(n11541), .Z(n11549) );
  XNOR U11233 ( .A(n11539), .B(n11548), .Z(n11541) );
  XNOR U11234 ( .A(n11550), .B(n11551), .Z(n11539) );
  AND U11235 ( .A(n1176), .B(n11552), .Z(n11551) );
  XOR U11236 ( .A(p_input[1787]), .B(n11550), .Z(n11552) );
  XNOR U11237 ( .A(n11553), .B(n11554), .Z(n11550) );
  AND U11238 ( .A(n1180), .B(n11555), .Z(n11554) );
  XOR U11239 ( .A(n11556), .B(n11557), .Z(n11548) );
  AND U11240 ( .A(n1184), .B(n11547), .Z(n11557) );
  XNOR U11241 ( .A(n11558), .B(n11545), .Z(n11547) );
  XOR U11242 ( .A(n11559), .B(n11560), .Z(n11545) );
  AND U11243 ( .A(n1207), .B(n11561), .Z(n11560) );
  IV U11244 ( .A(n11556), .Z(n11558) );
  XOR U11245 ( .A(n11562), .B(n11563), .Z(n11556) );
  AND U11246 ( .A(n1191), .B(n11555), .Z(n11563) );
  XNOR U11247 ( .A(n11553), .B(n11562), .Z(n11555) );
  XNOR U11248 ( .A(n11564), .B(n11565), .Z(n11553) );
  AND U11249 ( .A(n1195), .B(n11566), .Z(n11565) );
  XOR U11250 ( .A(p_input[1819]), .B(n11564), .Z(n11566) );
  XNOR U11251 ( .A(n11567), .B(n11568), .Z(n11564) );
  AND U11252 ( .A(n1199), .B(n11569), .Z(n11568) );
  XOR U11253 ( .A(n11570), .B(n11571), .Z(n11562) );
  AND U11254 ( .A(n1203), .B(n11561), .Z(n11571) );
  XNOR U11255 ( .A(n11572), .B(n11559), .Z(n11561) );
  XOR U11256 ( .A(n11573), .B(n11574), .Z(n11559) );
  AND U11257 ( .A(n1226), .B(n11575), .Z(n11574) );
  IV U11258 ( .A(n11570), .Z(n11572) );
  XOR U11259 ( .A(n11576), .B(n11577), .Z(n11570) );
  AND U11260 ( .A(n1210), .B(n11569), .Z(n11577) );
  XNOR U11261 ( .A(n11567), .B(n11576), .Z(n11569) );
  XNOR U11262 ( .A(n11578), .B(n11579), .Z(n11567) );
  AND U11263 ( .A(n1214), .B(n11580), .Z(n11579) );
  XOR U11264 ( .A(p_input[1851]), .B(n11578), .Z(n11580) );
  XNOR U11265 ( .A(n11581), .B(n11582), .Z(n11578) );
  AND U11266 ( .A(n1218), .B(n11583), .Z(n11582) );
  XOR U11267 ( .A(n11584), .B(n11585), .Z(n11576) );
  AND U11268 ( .A(n1222), .B(n11575), .Z(n11585) );
  XNOR U11269 ( .A(n11586), .B(n11573), .Z(n11575) );
  XOR U11270 ( .A(n11587), .B(n11588), .Z(n11573) );
  AND U11271 ( .A(n1245), .B(n11589), .Z(n11588) );
  IV U11272 ( .A(n11584), .Z(n11586) );
  XOR U11273 ( .A(n11590), .B(n11591), .Z(n11584) );
  AND U11274 ( .A(n1229), .B(n11583), .Z(n11591) );
  XNOR U11275 ( .A(n11581), .B(n11590), .Z(n11583) );
  XNOR U11276 ( .A(n11592), .B(n11593), .Z(n11581) );
  AND U11277 ( .A(n1233), .B(n11594), .Z(n11593) );
  XOR U11278 ( .A(p_input[1883]), .B(n11592), .Z(n11594) );
  XNOR U11279 ( .A(n11595), .B(n11596), .Z(n11592) );
  AND U11280 ( .A(n1237), .B(n11597), .Z(n11596) );
  XOR U11281 ( .A(n11598), .B(n11599), .Z(n11590) );
  AND U11282 ( .A(n1241), .B(n11589), .Z(n11599) );
  XNOR U11283 ( .A(n11600), .B(n11587), .Z(n11589) );
  XOR U11284 ( .A(n11601), .B(n11602), .Z(n11587) );
  AND U11285 ( .A(n1264), .B(n11603), .Z(n11602) );
  IV U11286 ( .A(n11598), .Z(n11600) );
  XOR U11287 ( .A(n11604), .B(n11605), .Z(n11598) );
  AND U11288 ( .A(n1248), .B(n11597), .Z(n11605) );
  XNOR U11289 ( .A(n11595), .B(n11604), .Z(n11597) );
  XNOR U11290 ( .A(n11606), .B(n11607), .Z(n11595) );
  AND U11291 ( .A(n1252), .B(n11608), .Z(n11607) );
  XOR U11292 ( .A(p_input[1915]), .B(n11606), .Z(n11608) );
  XNOR U11293 ( .A(n11609), .B(n11610), .Z(n11606) );
  AND U11294 ( .A(n1256), .B(n11611), .Z(n11610) );
  XOR U11295 ( .A(n11612), .B(n11613), .Z(n11604) );
  AND U11296 ( .A(n1260), .B(n11603), .Z(n11613) );
  XNOR U11297 ( .A(n11614), .B(n11601), .Z(n11603) );
  XOR U11298 ( .A(n11615), .B(n11616), .Z(n11601) );
  AND U11299 ( .A(n1282), .B(n11617), .Z(n11616) );
  IV U11300 ( .A(n11612), .Z(n11614) );
  XOR U11301 ( .A(n11618), .B(n11619), .Z(n11612) );
  AND U11302 ( .A(n1267), .B(n11611), .Z(n11619) );
  XNOR U11303 ( .A(n11609), .B(n11618), .Z(n11611) );
  XNOR U11304 ( .A(n11620), .B(n11621), .Z(n11609) );
  AND U11305 ( .A(n1271), .B(n11622), .Z(n11621) );
  XOR U11306 ( .A(p_input[1947]), .B(n11620), .Z(n11622) );
  XOR U11307 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][27] ), .B(n11623), 
        .Z(n11620) );
  AND U11308 ( .A(n1274), .B(n11624), .Z(n11623) );
  XOR U11309 ( .A(n11625), .B(n11626), .Z(n11618) );
  AND U11310 ( .A(n1278), .B(n11617), .Z(n11626) );
  XNOR U11311 ( .A(n11627), .B(n11615), .Z(n11617) );
  XOR U11312 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n11628), .Z(n11615) );
  AND U11313 ( .A(n1290), .B(n11629), .Z(n11628) );
  IV U11314 ( .A(n11625), .Z(n11627) );
  XOR U11315 ( .A(n11630), .B(n11631), .Z(n11625) );
  AND U11316 ( .A(n1285), .B(n11624), .Z(n11631) );
  XOR U11317 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][27] ), .B(n11630), 
        .Z(n11624) );
  XOR U11318 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .B(n11632), 
        .Z(n11630) );
  AND U11319 ( .A(n1287), .B(n11629), .Z(n11632) );
  XOR U11320 ( .A(n11633), .B(n11634), .Z(n11629) );
  IV U11321 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .Z(n11634)
         );
  IV U11322 ( .A(\knn_comb_/min_val_out[0][27] ), .Z(n11633) );
  XOR U11323 ( .A(n85), .B(n11635), .Z(o[26]) );
  AND U11324 ( .A(n122), .B(n11636), .Z(n85) );
  XOR U11325 ( .A(n86), .B(n11635), .Z(n11636) );
  XOR U11326 ( .A(n11637), .B(n11638), .Z(n11635) );
  AND U11327 ( .A(n142), .B(n11639), .Z(n11638) );
  XOR U11328 ( .A(n11640), .B(n13), .Z(n86) );
  AND U11329 ( .A(n125), .B(n11641), .Z(n13) );
  XOR U11330 ( .A(n14), .B(n11640), .Z(n11641) );
  XOR U11331 ( .A(n11642), .B(n11643), .Z(n14) );
  AND U11332 ( .A(n130), .B(n11644), .Z(n11643) );
  XOR U11333 ( .A(p_input[26]), .B(n11642), .Z(n11644) );
  XNOR U11334 ( .A(n11645), .B(n11646), .Z(n11642) );
  AND U11335 ( .A(n134), .B(n11647), .Z(n11646) );
  XOR U11336 ( .A(n11648), .B(n11649), .Z(n11640) );
  AND U11337 ( .A(n138), .B(n11639), .Z(n11649) );
  XNOR U11338 ( .A(n11650), .B(n11637), .Z(n11639) );
  XOR U11339 ( .A(n11651), .B(n11652), .Z(n11637) );
  AND U11340 ( .A(n162), .B(n11653), .Z(n11652) );
  IV U11341 ( .A(n11648), .Z(n11650) );
  XOR U11342 ( .A(n11654), .B(n11655), .Z(n11648) );
  AND U11343 ( .A(n146), .B(n11647), .Z(n11655) );
  XNOR U11344 ( .A(n11645), .B(n11654), .Z(n11647) );
  XNOR U11345 ( .A(n11656), .B(n11657), .Z(n11645) );
  AND U11346 ( .A(n150), .B(n11658), .Z(n11657) );
  XOR U11347 ( .A(p_input[58]), .B(n11656), .Z(n11658) );
  XNOR U11348 ( .A(n11659), .B(n11660), .Z(n11656) );
  AND U11349 ( .A(n154), .B(n11661), .Z(n11660) );
  XOR U11350 ( .A(n11662), .B(n11663), .Z(n11654) );
  AND U11351 ( .A(n158), .B(n11653), .Z(n11663) );
  XNOR U11352 ( .A(n11664), .B(n11651), .Z(n11653) );
  XOR U11353 ( .A(n11665), .B(n11666), .Z(n11651) );
  AND U11354 ( .A(n181), .B(n11667), .Z(n11666) );
  IV U11355 ( .A(n11662), .Z(n11664) );
  XOR U11356 ( .A(n11668), .B(n11669), .Z(n11662) );
  AND U11357 ( .A(n165), .B(n11661), .Z(n11669) );
  XNOR U11358 ( .A(n11659), .B(n11668), .Z(n11661) );
  XNOR U11359 ( .A(n11670), .B(n11671), .Z(n11659) );
  AND U11360 ( .A(n169), .B(n11672), .Z(n11671) );
  XOR U11361 ( .A(p_input[90]), .B(n11670), .Z(n11672) );
  XNOR U11362 ( .A(n11673), .B(n11674), .Z(n11670) );
  AND U11363 ( .A(n173), .B(n11675), .Z(n11674) );
  XOR U11364 ( .A(n11676), .B(n11677), .Z(n11668) );
  AND U11365 ( .A(n177), .B(n11667), .Z(n11677) );
  XNOR U11366 ( .A(n11678), .B(n11665), .Z(n11667) );
  XOR U11367 ( .A(n11679), .B(n11680), .Z(n11665) );
  AND U11368 ( .A(n200), .B(n11681), .Z(n11680) );
  IV U11369 ( .A(n11676), .Z(n11678) );
  XOR U11370 ( .A(n11682), .B(n11683), .Z(n11676) );
  AND U11371 ( .A(n184), .B(n11675), .Z(n11683) );
  XNOR U11372 ( .A(n11673), .B(n11682), .Z(n11675) );
  XNOR U11373 ( .A(n11684), .B(n11685), .Z(n11673) );
  AND U11374 ( .A(n188), .B(n11686), .Z(n11685) );
  XOR U11375 ( .A(p_input[122]), .B(n11684), .Z(n11686) );
  XNOR U11376 ( .A(n11687), .B(n11688), .Z(n11684) );
  AND U11377 ( .A(n192), .B(n11689), .Z(n11688) );
  XOR U11378 ( .A(n11690), .B(n11691), .Z(n11682) );
  AND U11379 ( .A(n196), .B(n11681), .Z(n11691) );
  XNOR U11380 ( .A(n11692), .B(n11679), .Z(n11681) );
  XOR U11381 ( .A(n11693), .B(n11694), .Z(n11679) );
  AND U11382 ( .A(n219), .B(n11695), .Z(n11694) );
  IV U11383 ( .A(n11690), .Z(n11692) );
  XOR U11384 ( .A(n11696), .B(n11697), .Z(n11690) );
  AND U11385 ( .A(n203), .B(n11689), .Z(n11697) );
  XNOR U11386 ( .A(n11687), .B(n11696), .Z(n11689) );
  XNOR U11387 ( .A(n11698), .B(n11699), .Z(n11687) );
  AND U11388 ( .A(n207), .B(n11700), .Z(n11699) );
  XOR U11389 ( .A(p_input[154]), .B(n11698), .Z(n11700) );
  XNOR U11390 ( .A(n11701), .B(n11702), .Z(n11698) );
  AND U11391 ( .A(n211), .B(n11703), .Z(n11702) );
  XOR U11392 ( .A(n11704), .B(n11705), .Z(n11696) );
  AND U11393 ( .A(n215), .B(n11695), .Z(n11705) );
  XNOR U11394 ( .A(n11706), .B(n11693), .Z(n11695) );
  XOR U11395 ( .A(n11707), .B(n11708), .Z(n11693) );
  AND U11396 ( .A(n238), .B(n11709), .Z(n11708) );
  IV U11397 ( .A(n11704), .Z(n11706) );
  XOR U11398 ( .A(n11710), .B(n11711), .Z(n11704) );
  AND U11399 ( .A(n222), .B(n11703), .Z(n11711) );
  XNOR U11400 ( .A(n11701), .B(n11710), .Z(n11703) );
  XNOR U11401 ( .A(n11712), .B(n11713), .Z(n11701) );
  AND U11402 ( .A(n226), .B(n11714), .Z(n11713) );
  XOR U11403 ( .A(p_input[186]), .B(n11712), .Z(n11714) );
  XNOR U11404 ( .A(n11715), .B(n11716), .Z(n11712) );
  AND U11405 ( .A(n230), .B(n11717), .Z(n11716) );
  XOR U11406 ( .A(n11718), .B(n11719), .Z(n11710) );
  AND U11407 ( .A(n234), .B(n11709), .Z(n11719) );
  XNOR U11408 ( .A(n11720), .B(n11707), .Z(n11709) );
  XOR U11409 ( .A(n11721), .B(n11722), .Z(n11707) );
  AND U11410 ( .A(n257), .B(n11723), .Z(n11722) );
  IV U11411 ( .A(n11718), .Z(n11720) );
  XOR U11412 ( .A(n11724), .B(n11725), .Z(n11718) );
  AND U11413 ( .A(n241), .B(n11717), .Z(n11725) );
  XNOR U11414 ( .A(n11715), .B(n11724), .Z(n11717) );
  XNOR U11415 ( .A(n11726), .B(n11727), .Z(n11715) );
  AND U11416 ( .A(n245), .B(n11728), .Z(n11727) );
  XOR U11417 ( .A(p_input[218]), .B(n11726), .Z(n11728) );
  XNOR U11418 ( .A(n11729), .B(n11730), .Z(n11726) );
  AND U11419 ( .A(n249), .B(n11731), .Z(n11730) );
  XOR U11420 ( .A(n11732), .B(n11733), .Z(n11724) );
  AND U11421 ( .A(n253), .B(n11723), .Z(n11733) );
  XNOR U11422 ( .A(n11734), .B(n11721), .Z(n11723) );
  XOR U11423 ( .A(n11735), .B(n11736), .Z(n11721) );
  AND U11424 ( .A(n276), .B(n11737), .Z(n11736) );
  IV U11425 ( .A(n11732), .Z(n11734) );
  XOR U11426 ( .A(n11738), .B(n11739), .Z(n11732) );
  AND U11427 ( .A(n260), .B(n11731), .Z(n11739) );
  XNOR U11428 ( .A(n11729), .B(n11738), .Z(n11731) );
  XNOR U11429 ( .A(n11740), .B(n11741), .Z(n11729) );
  AND U11430 ( .A(n264), .B(n11742), .Z(n11741) );
  XOR U11431 ( .A(p_input[250]), .B(n11740), .Z(n11742) );
  XNOR U11432 ( .A(n11743), .B(n11744), .Z(n11740) );
  AND U11433 ( .A(n268), .B(n11745), .Z(n11744) );
  XOR U11434 ( .A(n11746), .B(n11747), .Z(n11738) );
  AND U11435 ( .A(n272), .B(n11737), .Z(n11747) );
  XNOR U11436 ( .A(n11748), .B(n11735), .Z(n11737) );
  XOR U11437 ( .A(n11749), .B(n11750), .Z(n11735) );
  AND U11438 ( .A(n295), .B(n11751), .Z(n11750) );
  IV U11439 ( .A(n11746), .Z(n11748) );
  XOR U11440 ( .A(n11752), .B(n11753), .Z(n11746) );
  AND U11441 ( .A(n279), .B(n11745), .Z(n11753) );
  XNOR U11442 ( .A(n11743), .B(n11752), .Z(n11745) );
  XNOR U11443 ( .A(n11754), .B(n11755), .Z(n11743) );
  AND U11444 ( .A(n283), .B(n11756), .Z(n11755) );
  XOR U11445 ( .A(p_input[282]), .B(n11754), .Z(n11756) );
  XNOR U11446 ( .A(n11757), .B(n11758), .Z(n11754) );
  AND U11447 ( .A(n287), .B(n11759), .Z(n11758) );
  XOR U11448 ( .A(n11760), .B(n11761), .Z(n11752) );
  AND U11449 ( .A(n291), .B(n11751), .Z(n11761) );
  XNOR U11450 ( .A(n11762), .B(n11749), .Z(n11751) );
  XOR U11451 ( .A(n11763), .B(n11764), .Z(n11749) );
  AND U11452 ( .A(n314), .B(n11765), .Z(n11764) );
  IV U11453 ( .A(n11760), .Z(n11762) );
  XOR U11454 ( .A(n11766), .B(n11767), .Z(n11760) );
  AND U11455 ( .A(n298), .B(n11759), .Z(n11767) );
  XNOR U11456 ( .A(n11757), .B(n11766), .Z(n11759) );
  XNOR U11457 ( .A(n11768), .B(n11769), .Z(n11757) );
  AND U11458 ( .A(n302), .B(n11770), .Z(n11769) );
  XOR U11459 ( .A(p_input[314]), .B(n11768), .Z(n11770) );
  XNOR U11460 ( .A(n11771), .B(n11772), .Z(n11768) );
  AND U11461 ( .A(n306), .B(n11773), .Z(n11772) );
  XOR U11462 ( .A(n11774), .B(n11775), .Z(n11766) );
  AND U11463 ( .A(n310), .B(n11765), .Z(n11775) );
  XNOR U11464 ( .A(n11776), .B(n11763), .Z(n11765) );
  XOR U11465 ( .A(n11777), .B(n11778), .Z(n11763) );
  AND U11466 ( .A(n333), .B(n11779), .Z(n11778) );
  IV U11467 ( .A(n11774), .Z(n11776) );
  XOR U11468 ( .A(n11780), .B(n11781), .Z(n11774) );
  AND U11469 ( .A(n317), .B(n11773), .Z(n11781) );
  XNOR U11470 ( .A(n11771), .B(n11780), .Z(n11773) );
  XNOR U11471 ( .A(n11782), .B(n11783), .Z(n11771) );
  AND U11472 ( .A(n321), .B(n11784), .Z(n11783) );
  XOR U11473 ( .A(p_input[346]), .B(n11782), .Z(n11784) );
  XNOR U11474 ( .A(n11785), .B(n11786), .Z(n11782) );
  AND U11475 ( .A(n325), .B(n11787), .Z(n11786) );
  XOR U11476 ( .A(n11788), .B(n11789), .Z(n11780) );
  AND U11477 ( .A(n329), .B(n11779), .Z(n11789) );
  XNOR U11478 ( .A(n11790), .B(n11777), .Z(n11779) );
  XOR U11479 ( .A(n11791), .B(n11792), .Z(n11777) );
  AND U11480 ( .A(n352), .B(n11793), .Z(n11792) );
  IV U11481 ( .A(n11788), .Z(n11790) );
  XOR U11482 ( .A(n11794), .B(n11795), .Z(n11788) );
  AND U11483 ( .A(n336), .B(n11787), .Z(n11795) );
  XNOR U11484 ( .A(n11785), .B(n11794), .Z(n11787) );
  XNOR U11485 ( .A(n11796), .B(n11797), .Z(n11785) );
  AND U11486 ( .A(n340), .B(n11798), .Z(n11797) );
  XOR U11487 ( .A(p_input[378]), .B(n11796), .Z(n11798) );
  XNOR U11488 ( .A(n11799), .B(n11800), .Z(n11796) );
  AND U11489 ( .A(n344), .B(n11801), .Z(n11800) );
  XOR U11490 ( .A(n11802), .B(n11803), .Z(n11794) );
  AND U11491 ( .A(n348), .B(n11793), .Z(n11803) );
  XNOR U11492 ( .A(n11804), .B(n11791), .Z(n11793) );
  XOR U11493 ( .A(n11805), .B(n11806), .Z(n11791) );
  AND U11494 ( .A(n371), .B(n11807), .Z(n11806) );
  IV U11495 ( .A(n11802), .Z(n11804) );
  XOR U11496 ( .A(n11808), .B(n11809), .Z(n11802) );
  AND U11497 ( .A(n355), .B(n11801), .Z(n11809) );
  XNOR U11498 ( .A(n11799), .B(n11808), .Z(n11801) );
  XNOR U11499 ( .A(n11810), .B(n11811), .Z(n11799) );
  AND U11500 ( .A(n359), .B(n11812), .Z(n11811) );
  XOR U11501 ( .A(p_input[410]), .B(n11810), .Z(n11812) );
  XNOR U11502 ( .A(n11813), .B(n11814), .Z(n11810) );
  AND U11503 ( .A(n363), .B(n11815), .Z(n11814) );
  XOR U11504 ( .A(n11816), .B(n11817), .Z(n11808) );
  AND U11505 ( .A(n367), .B(n11807), .Z(n11817) );
  XNOR U11506 ( .A(n11818), .B(n11805), .Z(n11807) );
  XOR U11507 ( .A(n11819), .B(n11820), .Z(n11805) );
  AND U11508 ( .A(n390), .B(n11821), .Z(n11820) );
  IV U11509 ( .A(n11816), .Z(n11818) );
  XOR U11510 ( .A(n11822), .B(n11823), .Z(n11816) );
  AND U11511 ( .A(n374), .B(n11815), .Z(n11823) );
  XNOR U11512 ( .A(n11813), .B(n11822), .Z(n11815) );
  XNOR U11513 ( .A(n11824), .B(n11825), .Z(n11813) );
  AND U11514 ( .A(n378), .B(n11826), .Z(n11825) );
  XOR U11515 ( .A(p_input[442]), .B(n11824), .Z(n11826) );
  XNOR U11516 ( .A(n11827), .B(n11828), .Z(n11824) );
  AND U11517 ( .A(n382), .B(n11829), .Z(n11828) );
  XOR U11518 ( .A(n11830), .B(n11831), .Z(n11822) );
  AND U11519 ( .A(n386), .B(n11821), .Z(n11831) );
  XNOR U11520 ( .A(n11832), .B(n11819), .Z(n11821) );
  XOR U11521 ( .A(n11833), .B(n11834), .Z(n11819) );
  AND U11522 ( .A(n409), .B(n11835), .Z(n11834) );
  IV U11523 ( .A(n11830), .Z(n11832) );
  XOR U11524 ( .A(n11836), .B(n11837), .Z(n11830) );
  AND U11525 ( .A(n393), .B(n11829), .Z(n11837) );
  XNOR U11526 ( .A(n11827), .B(n11836), .Z(n11829) );
  XNOR U11527 ( .A(n11838), .B(n11839), .Z(n11827) );
  AND U11528 ( .A(n397), .B(n11840), .Z(n11839) );
  XOR U11529 ( .A(p_input[474]), .B(n11838), .Z(n11840) );
  XNOR U11530 ( .A(n11841), .B(n11842), .Z(n11838) );
  AND U11531 ( .A(n401), .B(n11843), .Z(n11842) );
  XOR U11532 ( .A(n11844), .B(n11845), .Z(n11836) );
  AND U11533 ( .A(n405), .B(n11835), .Z(n11845) );
  XNOR U11534 ( .A(n11846), .B(n11833), .Z(n11835) );
  XOR U11535 ( .A(n11847), .B(n11848), .Z(n11833) );
  AND U11536 ( .A(n428), .B(n11849), .Z(n11848) );
  IV U11537 ( .A(n11844), .Z(n11846) );
  XOR U11538 ( .A(n11850), .B(n11851), .Z(n11844) );
  AND U11539 ( .A(n412), .B(n11843), .Z(n11851) );
  XNOR U11540 ( .A(n11841), .B(n11850), .Z(n11843) );
  XNOR U11541 ( .A(n11852), .B(n11853), .Z(n11841) );
  AND U11542 ( .A(n416), .B(n11854), .Z(n11853) );
  XOR U11543 ( .A(p_input[506]), .B(n11852), .Z(n11854) );
  XNOR U11544 ( .A(n11855), .B(n11856), .Z(n11852) );
  AND U11545 ( .A(n420), .B(n11857), .Z(n11856) );
  XOR U11546 ( .A(n11858), .B(n11859), .Z(n11850) );
  AND U11547 ( .A(n424), .B(n11849), .Z(n11859) );
  XNOR U11548 ( .A(n11860), .B(n11847), .Z(n11849) );
  XOR U11549 ( .A(n11861), .B(n11862), .Z(n11847) );
  AND U11550 ( .A(n447), .B(n11863), .Z(n11862) );
  IV U11551 ( .A(n11858), .Z(n11860) );
  XOR U11552 ( .A(n11864), .B(n11865), .Z(n11858) );
  AND U11553 ( .A(n431), .B(n11857), .Z(n11865) );
  XNOR U11554 ( .A(n11855), .B(n11864), .Z(n11857) );
  XNOR U11555 ( .A(n11866), .B(n11867), .Z(n11855) );
  AND U11556 ( .A(n435), .B(n11868), .Z(n11867) );
  XOR U11557 ( .A(p_input[538]), .B(n11866), .Z(n11868) );
  XNOR U11558 ( .A(n11869), .B(n11870), .Z(n11866) );
  AND U11559 ( .A(n439), .B(n11871), .Z(n11870) );
  XOR U11560 ( .A(n11872), .B(n11873), .Z(n11864) );
  AND U11561 ( .A(n443), .B(n11863), .Z(n11873) );
  XNOR U11562 ( .A(n11874), .B(n11861), .Z(n11863) );
  XOR U11563 ( .A(n11875), .B(n11876), .Z(n11861) );
  AND U11564 ( .A(n466), .B(n11877), .Z(n11876) );
  IV U11565 ( .A(n11872), .Z(n11874) );
  XOR U11566 ( .A(n11878), .B(n11879), .Z(n11872) );
  AND U11567 ( .A(n450), .B(n11871), .Z(n11879) );
  XNOR U11568 ( .A(n11869), .B(n11878), .Z(n11871) );
  XNOR U11569 ( .A(n11880), .B(n11881), .Z(n11869) );
  AND U11570 ( .A(n454), .B(n11882), .Z(n11881) );
  XOR U11571 ( .A(p_input[570]), .B(n11880), .Z(n11882) );
  XNOR U11572 ( .A(n11883), .B(n11884), .Z(n11880) );
  AND U11573 ( .A(n458), .B(n11885), .Z(n11884) );
  XOR U11574 ( .A(n11886), .B(n11887), .Z(n11878) );
  AND U11575 ( .A(n462), .B(n11877), .Z(n11887) );
  XNOR U11576 ( .A(n11888), .B(n11875), .Z(n11877) );
  XOR U11577 ( .A(n11889), .B(n11890), .Z(n11875) );
  AND U11578 ( .A(n485), .B(n11891), .Z(n11890) );
  IV U11579 ( .A(n11886), .Z(n11888) );
  XOR U11580 ( .A(n11892), .B(n11893), .Z(n11886) );
  AND U11581 ( .A(n469), .B(n11885), .Z(n11893) );
  XNOR U11582 ( .A(n11883), .B(n11892), .Z(n11885) );
  XNOR U11583 ( .A(n11894), .B(n11895), .Z(n11883) );
  AND U11584 ( .A(n473), .B(n11896), .Z(n11895) );
  XOR U11585 ( .A(p_input[602]), .B(n11894), .Z(n11896) );
  XNOR U11586 ( .A(n11897), .B(n11898), .Z(n11894) );
  AND U11587 ( .A(n477), .B(n11899), .Z(n11898) );
  XOR U11588 ( .A(n11900), .B(n11901), .Z(n11892) );
  AND U11589 ( .A(n481), .B(n11891), .Z(n11901) );
  XNOR U11590 ( .A(n11902), .B(n11889), .Z(n11891) );
  XOR U11591 ( .A(n11903), .B(n11904), .Z(n11889) );
  AND U11592 ( .A(n504), .B(n11905), .Z(n11904) );
  IV U11593 ( .A(n11900), .Z(n11902) );
  XOR U11594 ( .A(n11906), .B(n11907), .Z(n11900) );
  AND U11595 ( .A(n488), .B(n11899), .Z(n11907) );
  XNOR U11596 ( .A(n11897), .B(n11906), .Z(n11899) );
  XNOR U11597 ( .A(n11908), .B(n11909), .Z(n11897) );
  AND U11598 ( .A(n492), .B(n11910), .Z(n11909) );
  XOR U11599 ( .A(p_input[634]), .B(n11908), .Z(n11910) );
  XNOR U11600 ( .A(n11911), .B(n11912), .Z(n11908) );
  AND U11601 ( .A(n496), .B(n11913), .Z(n11912) );
  XOR U11602 ( .A(n11914), .B(n11915), .Z(n11906) );
  AND U11603 ( .A(n500), .B(n11905), .Z(n11915) );
  XNOR U11604 ( .A(n11916), .B(n11903), .Z(n11905) );
  XOR U11605 ( .A(n11917), .B(n11918), .Z(n11903) );
  AND U11606 ( .A(n523), .B(n11919), .Z(n11918) );
  IV U11607 ( .A(n11914), .Z(n11916) );
  XOR U11608 ( .A(n11920), .B(n11921), .Z(n11914) );
  AND U11609 ( .A(n507), .B(n11913), .Z(n11921) );
  XNOR U11610 ( .A(n11911), .B(n11920), .Z(n11913) );
  XNOR U11611 ( .A(n11922), .B(n11923), .Z(n11911) );
  AND U11612 ( .A(n511), .B(n11924), .Z(n11923) );
  XOR U11613 ( .A(p_input[666]), .B(n11922), .Z(n11924) );
  XNOR U11614 ( .A(n11925), .B(n11926), .Z(n11922) );
  AND U11615 ( .A(n515), .B(n11927), .Z(n11926) );
  XOR U11616 ( .A(n11928), .B(n11929), .Z(n11920) );
  AND U11617 ( .A(n519), .B(n11919), .Z(n11929) );
  XNOR U11618 ( .A(n11930), .B(n11917), .Z(n11919) );
  XOR U11619 ( .A(n11931), .B(n11932), .Z(n11917) );
  AND U11620 ( .A(n542), .B(n11933), .Z(n11932) );
  IV U11621 ( .A(n11928), .Z(n11930) );
  XOR U11622 ( .A(n11934), .B(n11935), .Z(n11928) );
  AND U11623 ( .A(n526), .B(n11927), .Z(n11935) );
  XNOR U11624 ( .A(n11925), .B(n11934), .Z(n11927) );
  XNOR U11625 ( .A(n11936), .B(n11937), .Z(n11925) );
  AND U11626 ( .A(n530), .B(n11938), .Z(n11937) );
  XOR U11627 ( .A(p_input[698]), .B(n11936), .Z(n11938) );
  XNOR U11628 ( .A(n11939), .B(n11940), .Z(n11936) );
  AND U11629 ( .A(n534), .B(n11941), .Z(n11940) );
  XOR U11630 ( .A(n11942), .B(n11943), .Z(n11934) );
  AND U11631 ( .A(n538), .B(n11933), .Z(n11943) );
  XNOR U11632 ( .A(n11944), .B(n11931), .Z(n11933) );
  XOR U11633 ( .A(n11945), .B(n11946), .Z(n11931) );
  AND U11634 ( .A(n561), .B(n11947), .Z(n11946) );
  IV U11635 ( .A(n11942), .Z(n11944) );
  XOR U11636 ( .A(n11948), .B(n11949), .Z(n11942) );
  AND U11637 ( .A(n545), .B(n11941), .Z(n11949) );
  XNOR U11638 ( .A(n11939), .B(n11948), .Z(n11941) );
  XNOR U11639 ( .A(n11950), .B(n11951), .Z(n11939) );
  AND U11640 ( .A(n549), .B(n11952), .Z(n11951) );
  XOR U11641 ( .A(p_input[730]), .B(n11950), .Z(n11952) );
  XNOR U11642 ( .A(n11953), .B(n11954), .Z(n11950) );
  AND U11643 ( .A(n553), .B(n11955), .Z(n11954) );
  XOR U11644 ( .A(n11956), .B(n11957), .Z(n11948) );
  AND U11645 ( .A(n557), .B(n11947), .Z(n11957) );
  XNOR U11646 ( .A(n11958), .B(n11945), .Z(n11947) );
  XOR U11647 ( .A(n11959), .B(n11960), .Z(n11945) );
  AND U11648 ( .A(n580), .B(n11961), .Z(n11960) );
  IV U11649 ( .A(n11956), .Z(n11958) );
  XOR U11650 ( .A(n11962), .B(n11963), .Z(n11956) );
  AND U11651 ( .A(n564), .B(n11955), .Z(n11963) );
  XNOR U11652 ( .A(n11953), .B(n11962), .Z(n11955) );
  XNOR U11653 ( .A(n11964), .B(n11965), .Z(n11953) );
  AND U11654 ( .A(n568), .B(n11966), .Z(n11965) );
  XOR U11655 ( .A(p_input[762]), .B(n11964), .Z(n11966) );
  XNOR U11656 ( .A(n11967), .B(n11968), .Z(n11964) );
  AND U11657 ( .A(n572), .B(n11969), .Z(n11968) );
  XOR U11658 ( .A(n11970), .B(n11971), .Z(n11962) );
  AND U11659 ( .A(n576), .B(n11961), .Z(n11971) );
  XNOR U11660 ( .A(n11972), .B(n11959), .Z(n11961) );
  XOR U11661 ( .A(n11973), .B(n11974), .Z(n11959) );
  AND U11662 ( .A(n599), .B(n11975), .Z(n11974) );
  IV U11663 ( .A(n11970), .Z(n11972) );
  XOR U11664 ( .A(n11976), .B(n11977), .Z(n11970) );
  AND U11665 ( .A(n583), .B(n11969), .Z(n11977) );
  XNOR U11666 ( .A(n11967), .B(n11976), .Z(n11969) );
  XNOR U11667 ( .A(n11978), .B(n11979), .Z(n11967) );
  AND U11668 ( .A(n587), .B(n11980), .Z(n11979) );
  XOR U11669 ( .A(p_input[794]), .B(n11978), .Z(n11980) );
  XNOR U11670 ( .A(n11981), .B(n11982), .Z(n11978) );
  AND U11671 ( .A(n591), .B(n11983), .Z(n11982) );
  XOR U11672 ( .A(n11984), .B(n11985), .Z(n11976) );
  AND U11673 ( .A(n595), .B(n11975), .Z(n11985) );
  XNOR U11674 ( .A(n11986), .B(n11973), .Z(n11975) );
  XOR U11675 ( .A(n11987), .B(n11988), .Z(n11973) );
  AND U11676 ( .A(n618), .B(n11989), .Z(n11988) );
  IV U11677 ( .A(n11984), .Z(n11986) );
  XOR U11678 ( .A(n11990), .B(n11991), .Z(n11984) );
  AND U11679 ( .A(n602), .B(n11983), .Z(n11991) );
  XNOR U11680 ( .A(n11981), .B(n11990), .Z(n11983) );
  XNOR U11681 ( .A(n11992), .B(n11993), .Z(n11981) );
  AND U11682 ( .A(n606), .B(n11994), .Z(n11993) );
  XOR U11683 ( .A(p_input[826]), .B(n11992), .Z(n11994) );
  XNOR U11684 ( .A(n11995), .B(n11996), .Z(n11992) );
  AND U11685 ( .A(n610), .B(n11997), .Z(n11996) );
  XOR U11686 ( .A(n11998), .B(n11999), .Z(n11990) );
  AND U11687 ( .A(n614), .B(n11989), .Z(n11999) );
  XNOR U11688 ( .A(n12000), .B(n11987), .Z(n11989) );
  XOR U11689 ( .A(n12001), .B(n12002), .Z(n11987) );
  AND U11690 ( .A(n637), .B(n12003), .Z(n12002) );
  IV U11691 ( .A(n11998), .Z(n12000) );
  XOR U11692 ( .A(n12004), .B(n12005), .Z(n11998) );
  AND U11693 ( .A(n621), .B(n11997), .Z(n12005) );
  XNOR U11694 ( .A(n11995), .B(n12004), .Z(n11997) );
  XNOR U11695 ( .A(n12006), .B(n12007), .Z(n11995) );
  AND U11696 ( .A(n625), .B(n12008), .Z(n12007) );
  XOR U11697 ( .A(p_input[858]), .B(n12006), .Z(n12008) );
  XNOR U11698 ( .A(n12009), .B(n12010), .Z(n12006) );
  AND U11699 ( .A(n629), .B(n12011), .Z(n12010) );
  XOR U11700 ( .A(n12012), .B(n12013), .Z(n12004) );
  AND U11701 ( .A(n633), .B(n12003), .Z(n12013) );
  XNOR U11702 ( .A(n12014), .B(n12001), .Z(n12003) );
  XOR U11703 ( .A(n12015), .B(n12016), .Z(n12001) );
  AND U11704 ( .A(n656), .B(n12017), .Z(n12016) );
  IV U11705 ( .A(n12012), .Z(n12014) );
  XOR U11706 ( .A(n12018), .B(n12019), .Z(n12012) );
  AND U11707 ( .A(n640), .B(n12011), .Z(n12019) );
  XNOR U11708 ( .A(n12009), .B(n12018), .Z(n12011) );
  XNOR U11709 ( .A(n12020), .B(n12021), .Z(n12009) );
  AND U11710 ( .A(n644), .B(n12022), .Z(n12021) );
  XOR U11711 ( .A(p_input[890]), .B(n12020), .Z(n12022) );
  XNOR U11712 ( .A(n12023), .B(n12024), .Z(n12020) );
  AND U11713 ( .A(n648), .B(n12025), .Z(n12024) );
  XOR U11714 ( .A(n12026), .B(n12027), .Z(n12018) );
  AND U11715 ( .A(n652), .B(n12017), .Z(n12027) );
  XNOR U11716 ( .A(n12028), .B(n12015), .Z(n12017) );
  XOR U11717 ( .A(n12029), .B(n12030), .Z(n12015) );
  AND U11718 ( .A(n675), .B(n12031), .Z(n12030) );
  IV U11719 ( .A(n12026), .Z(n12028) );
  XOR U11720 ( .A(n12032), .B(n12033), .Z(n12026) );
  AND U11721 ( .A(n659), .B(n12025), .Z(n12033) );
  XNOR U11722 ( .A(n12023), .B(n12032), .Z(n12025) );
  XNOR U11723 ( .A(n12034), .B(n12035), .Z(n12023) );
  AND U11724 ( .A(n663), .B(n12036), .Z(n12035) );
  XOR U11725 ( .A(p_input[922]), .B(n12034), .Z(n12036) );
  XNOR U11726 ( .A(n12037), .B(n12038), .Z(n12034) );
  AND U11727 ( .A(n667), .B(n12039), .Z(n12038) );
  XOR U11728 ( .A(n12040), .B(n12041), .Z(n12032) );
  AND U11729 ( .A(n671), .B(n12031), .Z(n12041) );
  XNOR U11730 ( .A(n12042), .B(n12029), .Z(n12031) );
  XOR U11731 ( .A(n12043), .B(n12044), .Z(n12029) );
  AND U11732 ( .A(n694), .B(n12045), .Z(n12044) );
  IV U11733 ( .A(n12040), .Z(n12042) );
  XOR U11734 ( .A(n12046), .B(n12047), .Z(n12040) );
  AND U11735 ( .A(n678), .B(n12039), .Z(n12047) );
  XNOR U11736 ( .A(n12037), .B(n12046), .Z(n12039) );
  XNOR U11737 ( .A(n12048), .B(n12049), .Z(n12037) );
  AND U11738 ( .A(n682), .B(n12050), .Z(n12049) );
  XOR U11739 ( .A(p_input[954]), .B(n12048), .Z(n12050) );
  XNOR U11740 ( .A(n12051), .B(n12052), .Z(n12048) );
  AND U11741 ( .A(n686), .B(n12053), .Z(n12052) );
  XOR U11742 ( .A(n12054), .B(n12055), .Z(n12046) );
  AND U11743 ( .A(n690), .B(n12045), .Z(n12055) );
  XNOR U11744 ( .A(n12056), .B(n12043), .Z(n12045) );
  XOR U11745 ( .A(n12057), .B(n12058), .Z(n12043) );
  AND U11746 ( .A(n713), .B(n12059), .Z(n12058) );
  IV U11747 ( .A(n12054), .Z(n12056) );
  XOR U11748 ( .A(n12060), .B(n12061), .Z(n12054) );
  AND U11749 ( .A(n697), .B(n12053), .Z(n12061) );
  XNOR U11750 ( .A(n12051), .B(n12060), .Z(n12053) );
  XNOR U11751 ( .A(n12062), .B(n12063), .Z(n12051) );
  AND U11752 ( .A(n701), .B(n12064), .Z(n12063) );
  XOR U11753 ( .A(p_input[986]), .B(n12062), .Z(n12064) );
  XNOR U11754 ( .A(n12065), .B(n12066), .Z(n12062) );
  AND U11755 ( .A(n705), .B(n12067), .Z(n12066) );
  XOR U11756 ( .A(n12068), .B(n12069), .Z(n12060) );
  AND U11757 ( .A(n709), .B(n12059), .Z(n12069) );
  XNOR U11758 ( .A(n12070), .B(n12057), .Z(n12059) );
  XOR U11759 ( .A(n12071), .B(n12072), .Z(n12057) );
  AND U11760 ( .A(n732), .B(n12073), .Z(n12072) );
  IV U11761 ( .A(n12068), .Z(n12070) );
  XOR U11762 ( .A(n12074), .B(n12075), .Z(n12068) );
  AND U11763 ( .A(n716), .B(n12067), .Z(n12075) );
  XNOR U11764 ( .A(n12065), .B(n12074), .Z(n12067) );
  XNOR U11765 ( .A(n12076), .B(n12077), .Z(n12065) );
  AND U11766 ( .A(n720), .B(n12078), .Z(n12077) );
  XOR U11767 ( .A(p_input[1018]), .B(n12076), .Z(n12078) );
  XNOR U11768 ( .A(n12079), .B(n12080), .Z(n12076) );
  AND U11769 ( .A(n724), .B(n12081), .Z(n12080) );
  XOR U11770 ( .A(n12082), .B(n12083), .Z(n12074) );
  AND U11771 ( .A(n728), .B(n12073), .Z(n12083) );
  XNOR U11772 ( .A(n12084), .B(n12071), .Z(n12073) );
  XOR U11773 ( .A(n12085), .B(n12086), .Z(n12071) );
  AND U11774 ( .A(n751), .B(n12087), .Z(n12086) );
  IV U11775 ( .A(n12082), .Z(n12084) );
  XOR U11776 ( .A(n12088), .B(n12089), .Z(n12082) );
  AND U11777 ( .A(n735), .B(n12081), .Z(n12089) );
  XNOR U11778 ( .A(n12079), .B(n12088), .Z(n12081) );
  XNOR U11779 ( .A(n12090), .B(n12091), .Z(n12079) );
  AND U11780 ( .A(n739), .B(n12092), .Z(n12091) );
  XOR U11781 ( .A(p_input[1050]), .B(n12090), .Z(n12092) );
  XNOR U11782 ( .A(n12093), .B(n12094), .Z(n12090) );
  AND U11783 ( .A(n743), .B(n12095), .Z(n12094) );
  XOR U11784 ( .A(n12096), .B(n12097), .Z(n12088) );
  AND U11785 ( .A(n747), .B(n12087), .Z(n12097) );
  XNOR U11786 ( .A(n12098), .B(n12085), .Z(n12087) );
  XOR U11787 ( .A(n12099), .B(n12100), .Z(n12085) );
  AND U11788 ( .A(n770), .B(n12101), .Z(n12100) );
  IV U11789 ( .A(n12096), .Z(n12098) );
  XOR U11790 ( .A(n12102), .B(n12103), .Z(n12096) );
  AND U11791 ( .A(n754), .B(n12095), .Z(n12103) );
  XNOR U11792 ( .A(n12093), .B(n12102), .Z(n12095) );
  XNOR U11793 ( .A(n12104), .B(n12105), .Z(n12093) );
  AND U11794 ( .A(n758), .B(n12106), .Z(n12105) );
  XOR U11795 ( .A(p_input[1082]), .B(n12104), .Z(n12106) );
  XNOR U11796 ( .A(n12107), .B(n12108), .Z(n12104) );
  AND U11797 ( .A(n762), .B(n12109), .Z(n12108) );
  XOR U11798 ( .A(n12110), .B(n12111), .Z(n12102) );
  AND U11799 ( .A(n766), .B(n12101), .Z(n12111) );
  XNOR U11800 ( .A(n12112), .B(n12099), .Z(n12101) );
  XOR U11801 ( .A(n12113), .B(n12114), .Z(n12099) );
  AND U11802 ( .A(n789), .B(n12115), .Z(n12114) );
  IV U11803 ( .A(n12110), .Z(n12112) );
  XOR U11804 ( .A(n12116), .B(n12117), .Z(n12110) );
  AND U11805 ( .A(n773), .B(n12109), .Z(n12117) );
  XNOR U11806 ( .A(n12107), .B(n12116), .Z(n12109) );
  XNOR U11807 ( .A(n12118), .B(n12119), .Z(n12107) );
  AND U11808 ( .A(n777), .B(n12120), .Z(n12119) );
  XOR U11809 ( .A(p_input[1114]), .B(n12118), .Z(n12120) );
  XNOR U11810 ( .A(n12121), .B(n12122), .Z(n12118) );
  AND U11811 ( .A(n781), .B(n12123), .Z(n12122) );
  XOR U11812 ( .A(n12124), .B(n12125), .Z(n12116) );
  AND U11813 ( .A(n785), .B(n12115), .Z(n12125) );
  XNOR U11814 ( .A(n12126), .B(n12113), .Z(n12115) );
  XOR U11815 ( .A(n12127), .B(n12128), .Z(n12113) );
  AND U11816 ( .A(n808), .B(n12129), .Z(n12128) );
  IV U11817 ( .A(n12124), .Z(n12126) );
  XOR U11818 ( .A(n12130), .B(n12131), .Z(n12124) );
  AND U11819 ( .A(n792), .B(n12123), .Z(n12131) );
  XNOR U11820 ( .A(n12121), .B(n12130), .Z(n12123) );
  XNOR U11821 ( .A(n12132), .B(n12133), .Z(n12121) );
  AND U11822 ( .A(n796), .B(n12134), .Z(n12133) );
  XOR U11823 ( .A(p_input[1146]), .B(n12132), .Z(n12134) );
  XNOR U11824 ( .A(n12135), .B(n12136), .Z(n12132) );
  AND U11825 ( .A(n800), .B(n12137), .Z(n12136) );
  XOR U11826 ( .A(n12138), .B(n12139), .Z(n12130) );
  AND U11827 ( .A(n804), .B(n12129), .Z(n12139) );
  XNOR U11828 ( .A(n12140), .B(n12127), .Z(n12129) );
  XOR U11829 ( .A(n12141), .B(n12142), .Z(n12127) );
  AND U11830 ( .A(n827), .B(n12143), .Z(n12142) );
  IV U11831 ( .A(n12138), .Z(n12140) );
  XOR U11832 ( .A(n12144), .B(n12145), .Z(n12138) );
  AND U11833 ( .A(n811), .B(n12137), .Z(n12145) );
  XNOR U11834 ( .A(n12135), .B(n12144), .Z(n12137) );
  XNOR U11835 ( .A(n12146), .B(n12147), .Z(n12135) );
  AND U11836 ( .A(n815), .B(n12148), .Z(n12147) );
  XOR U11837 ( .A(p_input[1178]), .B(n12146), .Z(n12148) );
  XNOR U11838 ( .A(n12149), .B(n12150), .Z(n12146) );
  AND U11839 ( .A(n819), .B(n12151), .Z(n12150) );
  XOR U11840 ( .A(n12152), .B(n12153), .Z(n12144) );
  AND U11841 ( .A(n823), .B(n12143), .Z(n12153) );
  XNOR U11842 ( .A(n12154), .B(n12141), .Z(n12143) );
  XOR U11843 ( .A(n12155), .B(n12156), .Z(n12141) );
  AND U11844 ( .A(n846), .B(n12157), .Z(n12156) );
  IV U11845 ( .A(n12152), .Z(n12154) );
  XOR U11846 ( .A(n12158), .B(n12159), .Z(n12152) );
  AND U11847 ( .A(n830), .B(n12151), .Z(n12159) );
  XNOR U11848 ( .A(n12149), .B(n12158), .Z(n12151) );
  XNOR U11849 ( .A(n12160), .B(n12161), .Z(n12149) );
  AND U11850 ( .A(n834), .B(n12162), .Z(n12161) );
  XOR U11851 ( .A(p_input[1210]), .B(n12160), .Z(n12162) );
  XNOR U11852 ( .A(n12163), .B(n12164), .Z(n12160) );
  AND U11853 ( .A(n838), .B(n12165), .Z(n12164) );
  XOR U11854 ( .A(n12166), .B(n12167), .Z(n12158) );
  AND U11855 ( .A(n842), .B(n12157), .Z(n12167) );
  XNOR U11856 ( .A(n12168), .B(n12155), .Z(n12157) );
  XOR U11857 ( .A(n12169), .B(n12170), .Z(n12155) );
  AND U11858 ( .A(n865), .B(n12171), .Z(n12170) );
  IV U11859 ( .A(n12166), .Z(n12168) );
  XOR U11860 ( .A(n12172), .B(n12173), .Z(n12166) );
  AND U11861 ( .A(n849), .B(n12165), .Z(n12173) );
  XNOR U11862 ( .A(n12163), .B(n12172), .Z(n12165) );
  XNOR U11863 ( .A(n12174), .B(n12175), .Z(n12163) );
  AND U11864 ( .A(n853), .B(n12176), .Z(n12175) );
  XOR U11865 ( .A(p_input[1242]), .B(n12174), .Z(n12176) );
  XNOR U11866 ( .A(n12177), .B(n12178), .Z(n12174) );
  AND U11867 ( .A(n857), .B(n12179), .Z(n12178) );
  XOR U11868 ( .A(n12180), .B(n12181), .Z(n12172) );
  AND U11869 ( .A(n861), .B(n12171), .Z(n12181) );
  XNOR U11870 ( .A(n12182), .B(n12169), .Z(n12171) );
  XOR U11871 ( .A(n12183), .B(n12184), .Z(n12169) );
  AND U11872 ( .A(n884), .B(n12185), .Z(n12184) );
  IV U11873 ( .A(n12180), .Z(n12182) );
  XOR U11874 ( .A(n12186), .B(n12187), .Z(n12180) );
  AND U11875 ( .A(n868), .B(n12179), .Z(n12187) );
  XNOR U11876 ( .A(n12177), .B(n12186), .Z(n12179) );
  XNOR U11877 ( .A(n12188), .B(n12189), .Z(n12177) );
  AND U11878 ( .A(n872), .B(n12190), .Z(n12189) );
  XOR U11879 ( .A(p_input[1274]), .B(n12188), .Z(n12190) );
  XNOR U11880 ( .A(n12191), .B(n12192), .Z(n12188) );
  AND U11881 ( .A(n876), .B(n12193), .Z(n12192) );
  XOR U11882 ( .A(n12194), .B(n12195), .Z(n12186) );
  AND U11883 ( .A(n880), .B(n12185), .Z(n12195) );
  XNOR U11884 ( .A(n12196), .B(n12183), .Z(n12185) );
  XOR U11885 ( .A(n12197), .B(n12198), .Z(n12183) );
  AND U11886 ( .A(n903), .B(n12199), .Z(n12198) );
  IV U11887 ( .A(n12194), .Z(n12196) );
  XOR U11888 ( .A(n12200), .B(n12201), .Z(n12194) );
  AND U11889 ( .A(n887), .B(n12193), .Z(n12201) );
  XNOR U11890 ( .A(n12191), .B(n12200), .Z(n12193) );
  XNOR U11891 ( .A(n12202), .B(n12203), .Z(n12191) );
  AND U11892 ( .A(n891), .B(n12204), .Z(n12203) );
  XOR U11893 ( .A(p_input[1306]), .B(n12202), .Z(n12204) );
  XNOR U11894 ( .A(n12205), .B(n12206), .Z(n12202) );
  AND U11895 ( .A(n895), .B(n12207), .Z(n12206) );
  XOR U11896 ( .A(n12208), .B(n12209), .Z(n12200) );
  AND U11897 ( .A(n899), .B(n12199), .Z(n12209) );
  XNOR U11898 ( .A(n12210), .B(n12197), .Z(n12199) );
  XOR U11899 ( .A(n12211), .B(n12212), .Z(n12197) );
  AND U11900 ( .A(n922), .B(n12213), .Z(n12212) );
  IV U11901 ( .A(n12208), .Z(n12210) );
  XOR U11902 ( .A(n12214), .B(n12215), .Z(n12208) );
  AND U11903 ( .A(n906), .B(n12207), .Z(n12215) );
  XNOR U11904 ( .A(n12205), .B(n12214), .Z(n12207) );
  XNOR U11905 ( .A(n12216), .B(n12217), .Z(n12205) );
  AND U11906 ( .A(n910), .B(n12218), .Z(n12217) );
  XOR U11907 ( .A(p_input[1338]), .B(n12216), .Z(n12218) );
  XNOR U11908 ( .A(n12219), .B(n12220), .Z(n12216) );
  AND U11909 ( .A(n914), .B(n12221), .Z(n12220) );
  XOR U11910 ( .A(n12222), .B(n12223), .Z(n12214) );
  AND U11911 ( .A(n918), .B(n12213), .Z(n12223) );
  XNOR U11912 ( .A(n12224), .B(n12211), .Z(n12213) );
  XOR U11913 ( .A(n12225), .B(n12226), .Z(n12211) );
  AND U11914 ( .A(n941), .B(n12227), .Z(n12226) );
  IV U11915 ( .A(n12222), .Z(n12224) );
  XOR U11916 ( .A(n12228), .B(n12229), .Z(n12222) );
  AND U11917 ( .A(n925), .B(n12221), .Z(n12229) );
  XNOR U11918 ( .A(n12219), .B(n12228), .Z(n12221) );
  XNOR U11919 ( .A(n12230), .B(n12231), .Z(n12219) );
  AND U11920 ( .A(n929), .B(n12232), .Z(n12231) );
  XOR U11921 ( .A(p_input[1370]), .B(n12230), .Z(n12232) );
  XNOR U11922 ( .A(n12233), .B(n12234), .Z(n12230) );
  AND U11923 ( .A(n933), .B(n12235), .Z(n12234) );
  XOR U11924 ( .A(n12236), .B(n12237), .Z(n12228) );
  AND U11925 ( .A(n937), .B(n12227), .Z(n12237) );
  XNOR U11926 ( .A(n12238), .B(n12225), .Z(n12227) );
  XOR U11927 ( .A(n12239), .B(n12240), .Z(n12225) );
  AND U11928 ( .A(n960), .B(n12241), .Z(n12240) );
  IV U11929 ( .A(n12236), .Z(n12238) );
  XOR U11930 ( .A(n12242), .B(n12243), .Z(n12236) );
  AND U11931 ( .A(n944), .B(n12235), .Z(n12243) );
  XNOR U11932 ( .A(n12233), .B(n12242), .Z(n12235) );
  XNOR U11933 ( .A(n12244), .B(n12245), .Z(n12233) );
  AND U11934 ( .A(n948), .B(n12246), .Z(n12245) );
  XOR U11935 ( .A(p_input[1402]), .B(n12244), .Z(n12246) );
  XNOR U11936 ( .A(n12247), .B(n12248), .Z(n12244) );
  AND U11937 ( .A(n952), .B(n12249), .Z(n12248) );
  XOR U11938 ( .A(n12250), .B(n12251), .Z(n12242) );
  AND U11939 ( .A(n956), .B(n12241), .Z(n12251) );
  XNOR U11940 ( .A(n12252), .B(n12239), .Z(n12241) );
  XOR U11941 ( .A(n12253), .B(n12254), .Z(n12239) );
  AND U11942 ( .A(n979), .B(n12255), .Z(n12254) );
  IV U11943 ( .A(n12250), .Z(n12252) );
  XOR U11944 ( .A(n12256), .B(n12257), .Z(n12250) );
  AND U11945 ( .A(n963), .B(n12249), .Z(n12257) );
  XNOR U11946 ( .A(n12247), .B(n12256), .Z(n12249) );
  XNOR U11947 ( .A(n12258), .B(n12259), .Z(n12247) );
  AND U11948 ( .A(n967), .B(n12260), .Z(n12259) );
  XOR U11949 ( .A(p_input[1434]), .B(n12258), .Z(n12260) );
  XNOR U11950 ( .A(n12261), .B(n12262), .Z(n12258) );
  AND U11951 ( .A(n971), .B(n12263), .Z(n12262) );
  XOR U11952 ( .A(n12264), .B(n12265), .Z(n12256) );
  AND U11953 ( .A(n975), .B(n12255), .Z(n12265) );
  XNOR U11954 ( .A(n12266), .B(n12253), .Z(n12255) );
  XOR U11955 ( .A(n12267), .B(n12268), .Z(n12253) );
  AND U11956 ( .A(n998), .B(n12269), .Z(n12268) );
  IV U11957 ( .A(n12264), .Z(n12266) );
  XOR U11958 ( .A(n12270), .B(n12271), .Z(n12264) );
  AND U11959 ( .A(n982), .B(n12263), .Z(n12271) );
  XNOR U11960 ( .A(n12261), .B(n12270), .Z(n12263) );
  XNOR U11961 ( .A(n12272), .B(n12273), .Z(n12261) );
  AND U11962 ( .A(n986), .B(n12274), .Z(n12273) );
  XOR U11963 ( .A(p_input[1466]), .B(n12272), .Z(n12274) );
  XNOR U11964 ( .A(n12275), .B(n12276), .Z(n12272) );
  AND U11965 ( .A(n990), .B(n12277), .Z(n12276) );
  XOR U11966 ( .A(n12278), .B(n12279), .Z(n12270) );
  AND U11967 ( .A(n994), .B(n12269), .Z(n12279) );
  XNOR U11968 ( .A(n12280), .B(n12267), .Z(n12269) );
  XOR U11969 ( .A(n12281), .B(n12282), .Z(n12267) );
  AND U11970 ( .A(n1017), .B(n12283), .Z(n12282) );
  IV U11971 ( .A(n12278), .Z(n12280) );
  XOR U11972 ( .A(n12284), .B(n12285), .Z(n12278) );
  AND U11973 ( .A(n1001), .B(n12277), .Z(n12285) );
  XNOR U11974 ( .A(n12275), .B(n12284), .Z(n12277) );
  XNOR U11975 ( .A(n12286), .B(n12287), .Z(n12275) );
  AND U11976 ( .A(n1005), .B(n12288), .Z(n12287) );
  XOR U11977 ( .A(p_input[1498]), .B(n12286), .Z(n12288) );
  XNOR U11978 ( .A(n12289), .B(n12290), .Z(n12286) );
  AND U11979 ( .A(n1009), .B(n12291), .Z(n12290) );
  XOR U11980 ( .A(n12292), .B(n12293), .Z(n12284) );
  AND U11981 ( .A(n1013), .B(n12283), .Z(n12293) );
  XNOR U11982 ( .A(n12294), .B(n12281), .Z(n12283) );
  XOR U11983 ( .A(n12295), .B(n12296), .Z(n12281) );
  AND U11984 ( .A(n1036), .B(n12297), .Z(n12296) );
  IV U11985 ( .A(n12292), .Z(n12294) );
  XOR U11986 ( .A(n12298), .B(n12299), .Z(n12292) );
  AND U11987 ( .A(n1020), .B(n12291), .Z(n12299) );
  XNOR U11988 ( .A(n12289), .B(n12298), .Z(n12291) );
  XNOR U11989 ( .A(n12300), .B(n12301), .Z(n12289) );
  AND U11990 ( .A(n1024), .B(n12302), .Z(n12301) );
  XOR U11991 ( .A(p_input[1530]), .B(n12300), .Z(n12302) );
  XNOR U11992 ( .A(n12303), .B(n12304), .Z(n12300) );
  AND U11993 ( .A(n1028), .B(n12305), .Z(n12304) );
  XOR U11994 ( .A(n12306), .B(n12307), .Z(n12298) );
  AND U11995 ( .A(n1032), .B(n12297), .Z(n12307) );
  XNOR U11996 ( .A(n12308), .B(n12295), .Z(n12297) );
  XOR U11997 ( .A(n12309), .B(n12310), .Z(n12295) );
  AND U11998 ( .A(n1055), .B(n12311), .Z(n12310) );
  IV U11999 ( .A(n12306), .Z(n12308) );
  XOR U12000 ( .A(n12312), .B(n12313), .Z(n12306) );
  AND U12001 ( .A(n1039), .B(n12305), .Z(n12313) );
  XNOR U12002 ( .A(n12303), .B(n12312), .Z(n12305) );
  XNOR U12003 ( .A(n12314), .B(n12315), .Z(n12303) );
  AND U12004 ( .A(n1043), .B(n12316), .Z(n12315) );
  XOR U12005 ( .A(p_input[1562]), .B(n12314), .Z(n12316) );
  XNOR U12006 ( .A(n12317), .B(n12318), .Z(n12314) );
  AND U12007 ( .A(n1047), .B(n12319), .Z(n12318) );
  XOR U12008 ( .A(n12320), .B(n12321), .Z(n12312) );
  AND U12009 ( .A(n1051), .B(n12311), .Z(n12321) );
  XNOR U12010 ( .A(n12322), .B(n12309), .Z(n12311) );
  XOR U12011 ( .A(n12323), .B(n12324), .Z(n12309) );
  AND U12012 ( .A(n1074), .B(n12325), .Z(n12324) );
  IV U12013 ( .A(n12320), .Z(n12322) );
  XOR U12014 ( .A(n12326), .B(n12327), .Z(n12320) );
  AND U12015 ( .A(n1058), .B(n12319), .Z(n12327) );
  XNOR U12016 ( .A(n12317), .B(n12326), .Z(n12319) );
  XNOR U12017 ( .A(n12328), .B(n12329), .Z(n12317) );
  AND U12018 ( .A(n1062), .B(n12330), .Z(n12329) );
  XOR U12019 ( .A(p_input[1594]), .B(n12328), .Z(n12330) );
  XNOR U12020 ( .A(n12331), .B(n12332), .Z(n12328) );
  AND U12021 ( .A(n1066), .B(n12333), .Z(n12332) );
  XOR U12022 ( .A(n12334), .B(n12335), .Z(n12326) );
  AND U12023 ( .A(n1070), .B(n12325), .Z(n12335) );
  XNOR U12024 ( .A(n12336), .B(n12323), .Z(n12325) );
  XOR U12025 ( .A(n12337), .B(n12338), .Z(n12323) );
  AND U12026 ( .A(n1093), .B(n12339), .Z(n12338) );
  IV U12027 ( .A(n12334), .Z(n12336) );
  XOR U12028 ( .A(n12340), .B(n12341), .Z(n12334) );
  AND U12029 ( .A(n1077), .B(n12333), .Z(n12341) );
  XNOR U12030 ( .A(n12331), .B(n12340), .Z(n12333) );
  XNOR U12031 ( .A(n12342), .B(n12343), .Z(n12331) );
  AND U12032 ( .A(n1081), .B(n12344), .Z(n12343) );
  XOR U12033 ( .A(p_input[1626]), .B(n12342), .Z(n12344) );
  XNOR U12034 ( .A(n12345), .B(n12346), .Z(n12342) );
  AND U12035 ( .A(n1085), .B(n12347), .Z(n12346) );
  XOR U12036 ( .A(n12348), .B(n12349), .Z(n12340) );
  AND U12037 ( .A(n1089), .B(n12339), .Z(n12349) );
  XNOR U12038 ( .A(n12350), .B(n12337), .Z(n12339) );
  XOR U12039 ( .A(n12351), .B(n12352), .Z(n12337) );
  AND U12040 ( .A(n1112), .B(n12353), .Z(n12352) );
  IV U12041 ( .A(n12348), .Z(n12350) );
  XOR U12042 ( .A(n12354), .B(n12355), .Z(n12348) );
  AND U12043 ( .A(n1096), .B(n12347), .Z(n12355) );
  XNOR U12044 ( .A(n12345), .B(n12354), .Z(n12347) );
  XNOR U12045 ( .A(n12356), .B(n12357), .Z(n12345) );
  AND U12046 ( .A(n1100), .B(n12358), .Z(n12357) );
  XOR U12047 ( .A(p_input[1658]), .B(n12356), .Z(n12358) );
  XNOR U12048 ( .A(n12359), .B(n12360), .Z(n12356) );
  AND U12049 ( .A(n1104), .B(n12361), .Z(n12360) );
  XOR U12050 ( .A(n12362), .B(n12363), .Z(n12354) );
  AND U12051 ( .A(n1108), .B(n12353), .Z(n12363) );
  XNOR U12052 ( .A(n12364), .B(n12351), .Z(n12353) );
  XOR U12053 ( .A(n12365), .B(n12366), .Z(n12351) );
  AND U12054 ( .A(n1131), .B(n12367), .Z(n12366) );
  IV U12055 ( .A(n12362), .Z(n12364) );
  XOR U12056 ( .A(n12368), .B(n12369), .Z(n12362) );
  AND U12057 ( .A(n1115), .B(n12361), .Z(n12369) );
  XNOR U12058 ( .A(n12359), .B(n12368), .Z(n12361) );
  XNOR U12059 ( .A(n12370), .B(n12371), .Z(n12359) );
  AND U12060 ( .A(n1119), .B(n12372), .Z(n12371) );
  XOR U12061 ( .A(p_input[1690]), .B(n12370), .Z(n12372) );
  XNOR U12062 ( .A(n12373), .B(n12374), .Z(n12370) );
  AND U12063 ( .A(n1123), .B(n12375), .Z(n12374) );
  XOR U12064 ( .A(n12376), .B(n12377), .Z(n12368) );
  AND U12065 ( .A(n1127), .B(n12367), .Z(n12377) );
  XNOR U12066 ( .A(n12378), .B(n12365), .Z(n12367) );
  XOR U12067 ( .A(n12379), .B(n12380), .Z(n12365) );
  AND U12068 ( .A(n1150), .B(n12381), .Z(n12380) );
  IV U12069 ( .A(n12376), .Z(n12378) );
  XOR U12070 ( .A(n12382), .B(n12383), .Z(n12376) );
  AND U12071 ( .A(n1134), .B(n12375), .Z(n12383) );
  XNOR U12072 ( .A(n12373), .B(n12382), .Z(n12375) );
  XNOR U12073 ( .A(n12384), .B(n12385), .Z(n12373) );
  AND U12074 ( .A(n1138), .B(n12386), .Z(n12385) );
  XOR U12075 ( .A(p_input[1722]), .B(n12384), .Z(n12386) );
  XNOR U12076 ( .A(n12387), .B(n12388), .Z(n12384) );
  AND U12077 ( .A(n1142), .B(n12389), .Z(n12388) );
  XOR U12078 ( .A(n12390), .B(n12391), .Z(n12382) );
  AND U12079 ( .A(n1146), .B(n12381), .Z(n12391) );
  XNOR U12080 ( .A(n12392), .B(n12379), .Z(n12381) );
  XOR U12081 ( .A(n12393), .B(n12394), .Z(n12379) );
  AND U12082 ( .A(n1169), .B(n12395), .Z(n12394) );
  IV U12083 ( .A(n12390), .Z(n12392) );
  XOR U12084 ( .A(n12396), .B(n12397), .Z(n12390) );
  AND U12085 ( .A(n1153), .B(n12389), .Z(n12397) );
  XNOR U12086 ( .A(n12387), .B(n12396), .Z(n12389) );
  XNOR U12087 ( .A(n12398), .B(n12399), .Z(n12387) );
  AND U12088 ( .A(n1157), .B(n12400), .Z(n12399) );
  XOR U12089 ( .A(p_input[1754]), .B(n12398), .Z(n12400) );
  XNOR U12090 ( .A(n12401), .B(n12402), .Z(n12398) );
  AND U12091 ( .A(n1161), .B(n12403), .Z(n12402) );
  XOR U12092 ( .A(n12404), .B(n12405), .Z(n12396) );
  AND U12093 ( .A(n1165), .B(n12395), .Z(n12405) );
  XNOR U12094 ( .A(n12406), .B(n12393), .Z(n12395) );
  XOR U12095 ( .A(n12407), .B(n12408), .Z(n12393) );
  AND U12096 ( .A(n1188), .B(n12409), .Z(n12408) );
  IV U12097 ( .A(n12404), .Z(n12406) );
  XOR U12098 ( .A(n12410), .B(n12411), .Z(n12404) );
  AND U12099 ( .A(n1172), .B(n12403), .Z(n12411) );
  XNOR U12100 ( .A(n12401), .B(n12410), .Z(n12403) );
  XNOR U12101 ( .A(n12412), .B(n12413), .Z(n12401) );
  AND U12102 ( .A(n1176), .B(n12414), .Z(n12413) );
  XOR U12103 ( .A(p_input[1786]), .B(n12412), .Z(n12414) );
  XNOR U12104 ( .A(n12415), .B(n12416), .Z(n12412) );
  AND U12105 ( .A(n1180), .B(n12417), .Z(n12416) );
  XOR U12106 ( .A(n12418), .B(n12419), .Z(n12410) );
  AND U12107 ( .A(n1184), .B(n12409), .Z(n12419) );
  XNOR U12108 ( .A(n12420), .B(n12407), .Z(n12409) );
  XOR U12109 ( .A(n12421), .B(n12422), .Z(n12407) );
  AND U12110 ( .A(n1207), .B(n12423), .Z(n12422) );
  IV U12111 ( .A(n12418), .Z(n12420) );
  XOR U12112 ( .A(n12424), .B(n12425), .Z(n12418) );
  AND U12113 ( .A(n1191), .B(n12417), .Z(n12425) );
  XNOR U12114 ( .A(n12415), .B(n12424), .Z(n12417) );
  XNOR U12115 ( .A(n12426), .B(n12427), .Z(n12415) );
  AND U12116 ( .A(n1195), .B(n12428), .Z(n12427) );
  XOR U12117 ( .A(p_input[1818]), .B(n12426), .Z(n12428) );
  XNOR U12118 ( .A(n12429), .B(n12430), .Z(n12426) );
  AND U12119 ( .A(n1199), .B(n12431), .Z(n12430) );
  XOR U12120 ( .A(n12432), .B(n12433), .Z(n12424) );
  AND U12121 ( .A(n1203), .B(n12423), .Z(n12433) );
  XNOR U12122 ( .A(n12434), .B(n12421), .Z(n12423) );
  XOR U12123 ( .A(n12435), .B(n12436), .Z(n12421) );
  AND U12124 ( .A(n1226), .B(n12437), .Z(n12436) );
  IV U12125 ( .A(n12432), .Z(n12434) );
  XOR U12126 ( .A(n12438), .B(n12439), .Z(n12432) );
  AND U12127 ( .A(n1210), .B(n12431), .Z(n12439) );
  XNOR U12128 ( .A(n12429), .B(n12438), .Z(n12431) );
  XNOR U12129 ( .A(n12440), .B(n12441), .Z(n12429) );
  AND U12130 ( .A(n1214), .B(n12442), .Z(n12441) );
  XOR U12131 ( .A(p_input[1850]), .B(n12440), .Z(n12442) );
  XNOR U12132 ( .A(n12443), .B(n12444), .Z(n12440) );
  AND U12133 ( .A(n1218), .B(n12445), .Z(n12444) );
  XOR U12134 ( .A(n12446), .B(n12447), .Z(n12438) );
  AND U12135 ( .A(n1222), .B(n12437), .Z(n12447) );
  XNOR U12136 ( .A(n12448), .B(n12435), .Z(n12437) );
  XOR U12137 ( .A(n12449), .B(n12450), .Z(n12435) );
  AND U12138 ( .A(n1245), .B(n12451), .Z(n12450) );
  IV U12139 ( .A(n12446), .Z(n12448) );
  XOR U12140 ( .A(n12452), .B(n12453), .Z(n12446) );
  AND U12141 ( .A(n1229), .B(n12445), .Z(n12453) );
  XNOR U12142 ( .A(n12443), .B(n12452), .Z(n12445) );
  XNOR U12143 ( .A(n12454), .B(n12455), .Z(n12443) );
  AND U12144 ( .A(n1233), .B(n12456), .Z(n12455) );
  XOR U12145 ( .A(p_input[1882]), .B(n12454), .Z(n12456) );
  XNOR U12146 ( .A(n12457), .B(n12458), .Z(n12454) );
  AND U12147 ( .A(n1237), .B(n12459), .Z(n12458) );
  XOR U12148 ( .A(n12460), .B(n12461), .Z(n12452) );
  AND U12149 ( .A(n1241), .B(n12451), .Z(n12461) );
  XNOR U12150 ( .A(n12462), .B(n12449), .Z(n12451) );
  XOR U12151 ( .A(n12463), .B(n12464), .Z(n12449) );
  AND U12152 ( .A(n1264), .B(n12465), .Z(n12464) );
  IV U12153 ( .A(n12460), .Z(n12462) );
  XOR U12154 ( .A(n12466), .B(n12467), .Z(n12460) );
  AND U12155 ( .A(n1248), .B(n12459), .Z(n12467) );
  XNOR U12156 ( .A(n12457), .B(n12466), .Z(n12459) );
  XNOR U12157 ( .A(n12468), .B(n12469), .Z(n12457) );
  AND U12158 ( .A(n1252), .B(n12470), .Z(n12469) );
  XOR U12159 ( .A(p_input[1914]), .B(n12468), .Z(n12470) );
  XNOR U12160 ( .A(n12471), .B(n12472), .Z(n12468) );
  AND U12161 ( .A(n1256), .B(n12473), .Z(n12472) );
  XOR U12162 ( .A(n12474), .B(n12475), .Z(n12466) );
  AND U12163 ( .A(n1260), .B(n12465), .Z(n12475) );
  XNOR U12164 ( .A(n12476), .B(n12463), .Z(n12465) );
  XOR U12165 ( .A(n12477), .B(n12478), .Z(n12463) );
  AND U12166 ( .A(n1282), .B(n12479), .Z(n12478) );
  IV U12167 ( .A(n12474), .Z(n12476) );
  XOR U12168 ( .A(n12480), .B(n12481), .Z(n12474) );
  AND U12169 ( .A(n1267), .B(n12473), .Z(n12481) );
  XNOR U12170 ( .A(n12471), .B(n12480), .Z(n12473) );
  XNOR U12171 ( .A(n12482), .B(n12483), .Z(n12471) );
  AND U12172 ( .A(n1271), .B(n12484), .Z(n12483) );
  XOR U12173 ( .A(p_input[1946]), .B(n12482), .Z(n12484) );
  XOR U12174 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][26] ), .B(n12485), 
        .Z(n12482) );
  AND U12175 ( .A(n1274), .B(n12486), .Z(n12485) );
  XOR U12176 ( .A(n12487), .B(n12488), .Z(n12480) );
  AND U12177 ( .A(n1278), .B(n12479), .Z(n12488) );
  XNOR U12178 ( .A(n12489), .B(n12477), .Z(n12479) );
  XOR U12179 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n12490), .Z(n12477) );
  AND U12180 ( .A(n1290), .B(n12491), .Z(n12490) );
  IV U12181 ( .A(n12487), .Z(n12489) );
  XOR U12182 ( .A(n12492), .B(n12493), .Z(n12487) );
  AND U12183 ( .A(n1285), .B(n12486), .Z(n12493) );
  XOR U12184 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][26] ), .B(n12492), 
        .Z(n12486) );
  XOR U12185 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .B(n12494), 
        .Z(n12492) );
  AND U12186 ( .A(n1287), .B(n12491), .Z(n12494) );
  XOR U12187 ( .A(\knn_comb_/min_val_out[0][26] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .Z(n12491) );
  XOR U12188 ( .A(n87), .B(n12495), .Z(o[25]) );
  AND U12189 ( .A(n122), .B(n12496), .Z(n87) );
  XOR U12190 ( .A(n88), .B(n12495), .Z(n12496) );
  XOR U12191 ( .A(n12497), .B(n12498), .Z(n12495) );
  AND U12192 ( .A(n142), .B(n12499), .Z(n12498) );
  XOR U12193 ( .A(n12500), .B(n17), .Z(n88) );
  AND U12194 ( .A(n125), .B(n12501), .Z(n17) );
  XOR U12195 ( .A(n18), .B(n12500), .Z(n12501) );
  XOR U12196 ( .A(n12502), .B(n12503), .Z(n18) );
  AND U12197 ( .A(n130), .B(n12504), .Z(n12503) );
  XOR U12198 ( .A(p_input[25]), .B(n12502), .Z(n12504) );
  XNOR U12199 ( .A(n12505), .B(n12506), .Z(n12502) );
  AND U12200 ( .A(n134), .B(n12507), .Z(n12506) );
  XOR U12201 ( .A(n12508), .B(n12509), .Z(n12500) );
  AND U12202 ( .A(n138), .B(n12499), .Z(n12509) );
  XNOR U12203 ( .A(n12510), .B(n12497), .Z(n12499) );
  XOR U12204 ( .A(n12511), .B(n12512), .Z(n12497) );
  AND U12205 ( .A(n162), .B(n12513), .Z(n12512) );
  IV U12206 ( .A(n12508), .Z(n12510) );
  XOR U12207 ( .A(n12514), .B(n12515), .Z(n12508) );
  AND U12208 ( .A(n146), .B(n12507), .Z(n12515) );
  XNOR U12209 ( .A(n12505), .B(n12514), .Z(n12507) );
  XNOR U12210 ( .A(n12516), .B(n12517), .Z(n12505) );
  AND U12211 ( .A(n150), .B(n12518), .Z(n12517) );
  XOR U12212 ( .A(p_input[57]), .B(n12516), .Z(n12518) );
  XNOR U12213 ( .A(n12519), .B(n12520), .Z(n12516) );
  AND U12214 ( .A(n154), .B(n12521), .Z(n12520) );
  XOR U12215 ( .A(n12522), .B(n12523), .Z(n12514) );
  AND U12216 ( .A(n158), .B(n12513), .Z(n12523) );
  XNOR U12217 ( .A(n12524), .B(n12511), .Z(n12513) );
  XOR U12218 ( .A(n12525), .B(n12526), .Z(n12511) );
  AND U12219 ( .A(n181), .B(n12527), .Z(n12526) );
  IV U12220 ( .A(n12522), .Z(n12524) );
  XOR U12221 ( .A(n12528), .B(n12529), .Z(n12522) );
  AND U12222 ( .A(n165), .B(n12521), .Z(n12529) );
  XNOR U12223 ( .A(n12519), .B(n12528), .Z(n12521) );
  XNOR U12224 ( .A(n12530), .B(n12531), .Z(n12519) );
  AND U12225 ( .A(n169), .B(n12532), .Z(n12531) );
  XOR U12226 ( .A(p_input[89]), .B(n12530), .Z(n12532) );
  XNOR U12227 ( .A(n12533), .B(n12534), .Z(n12530) );
  AND U12228 ( .A(n173), .B(n12535), .Z(n12534) );
  XOR U12229 ( .A(n12536), .B(n12537), .Z(n12528) );
  AND U12230 ( .A(n177), .B(n12527), .Z(n12537) );
  XNOR U12231 ( .A(n12538), .B(n12525), .Z(n12527) );
  XOR U12232 ( .A(n12539), .B(n12540), .Z(n12525) );
  AND U12233 ( .A(n200), .B(n12541), .Z(n12540) );
  IV U12234 ( .A(n12536), .Z(n12538) );
  XOR U12235 ( .A(n12542), .B(n12543), .Z(n12536) );
  AND U12236 ( .A(n184), .B(n12535), .Z(n12543) );
  XNOR U12237 ( .A(n12533), .B(n12542), .Z(n12535) );
  XNOR U12238 ( .A(n12544), .B(n12545), .Z(n12533) );
  AND U12239 ( .A(n188), .B(n12546), .Z(n12545) );
  XOR U12240 ( .A(p_input[121]), .B(n12544), .Z(n12546) );
  XNOR U12241 ( .A(n12547), .B(n12548), .Z(n12544) );
  AND U12242 ( .A(n192), .B(n12549), .Z(n12548) );
  XOR U12243 ( .A(n12550), .B(n12551), .Z(n12542) );
  AND U12244 ( .A(n196), .B(n12541), .Z(n12551) );
  XNOR U12245 ( .A(n12552), .B(n12539), .Z(n12541) );
  XOR U12246 ( .A(n12553), .B(n12554), .Z(n12539) );
  AND U12247 ( .A(n219), .B(n12555), .Z(n12554) );
  IV U12248 ( .A(n12550), .Z(n12552) );
  XOR U12249 ( .A(n12556), .B(n12557), .Z(n12550) );
  AND U12250 ( .A(n203), .B(n12549), .Z(n12557) );
  XNOR U12251 ( .A(n12547), .B(n12556), .Z(n12549) );
  XNOR U12252 ( .A(n12558), .B(n12559), .Z(n12547) );
  AND U12253 ( .A(n207), .B(n12560), .Z(n12559) );
  XOR U12254 ( .A(p_input[153]), .B(n12558), .Z(n12560) );
  XNOR U12255 ( .A(n12561), .B(n12562), .Z(n12558) );
  AND U12256 ( .A(n211), .B(n12563), .Z(n12562) );
  XOR U12257 ( .A(n12564), .B(n12565), .Z(n12556) );
  AND U12258 ( .A(n215), .B(n12555), .Z(n12565) );
  XNOR U12259 ( .A(n12566), .B(n12553), .Z(n12555) );
  XOR U12260 ( .A(n12567), .B(n12568), .Z(n12553) );
  AND U12261 ( .A(n238), .B(n12569), .Z(n12568) );
  IV U12262 ( .A(n12564), .Z(n12566) );
  XOR U12263 ( .A(n12570), .B(n12571), .Z(n12564) );
  AND U12264 ( .A(n222), .B(n12563), .Z(n12571) );
  XNOR U12265 ( .A(n12561), .B(n12570), .Z(n12563) );
  XNOR U12266 ( .A(n12572), .B(n12573), .Z(n12561) );
  AND U12267 ( .A(n226), .B(n12574), .Z(n12573) );
  XOR U12268 ( .A(p_input[185]), .B(n12572), .Z(n12574) );
  XNOR U12269 ( .A(n12575), .B(n12576), .Z(n12572) );
  AND U12270 ( .A(n230), .B(n12577), .Z(n12576) );
  XOR U12271 ( .A(n12578), .B(n12579), .Z(n12570) );
  AND U12272 ( .A(n234), .B(n12569), .Z(n12579) );
  XNOR U12273 ( .A(n12580), .B(n12567), .Z(n12569) );
  XOR U12274 ( .A(n12581), .B(n12582), .Z(n12567) );
  AND U12275 ( .A(n257), .B(n12583), .Z(n12582) );
  IV U12276 ( .A(n12578), .Z(n12580) );
  XOR U12277 ( .A(n12584), .B(n12585), .Z(n12578) );
  AND U12278 ( .A(n241), .B(n12577), .Z(n12585) );
  XNOR U12279 ( .A(n12575), .B(n12584), .Z(n12577) );
  XNOR U12280 ( .A(n12586), .B(n12587), .Z(n12575) );
  AND U12281 ( .A(n245), .B(n12588), .Z(n12587) );
  XOR U12282 ( .A(p_input[217]), .B(n12586), .Z(n12588) );
  XNOR U12283 ( .A(n12589), .B(n12590), .Z(n12586) );
  AND U12284 ( .A(n249), .B(n12591), .Z(n12590) );
  XOR U12285 ( .A(n12592), .B(n12593), .Z(n12584) );
  AND U12286 ( .A(n253), .B(n12583), .Z(n12593) );
  XNOR U12287 ( .A(n12594), .B(n12581), .Z(n12583) );
  XOR U12288 ( .A(n12595), .B(n12596), .Z(n12581) );
  AND U12289 ( .A(n276), .B(n12597), .Z(n12596) );
  IV U12290 ( .A(n12592), .Z(n12594) );
  XOR U12291 ( .A(n12598), .B(n12599), .Z(n12592) );
  AND U12292 ( .A(n260), .B(n12591), .Z(n12599) );
  XNOR U12293 ( .A(n12589), .B(n12598), .Z(n12591) );
  XNOR U12294 ( .A(n12600), .B(n12601), .Z(n12589) );
  AND U12295 ( .A(n264), .B(n12602), .Z(n12601) );
  XOR U12296 ( .A(p_input[249]), .B(n12600), .Z(n12602) );
  XNOR U12297 ( .A(n12603), .B(n12604), .Z(n12600) );
  AND U12298 ( .A(n268), .B(n12605), .Z(n12604) );
  XOR U12299 ( .A(n12606), .B(n12607), .Z(n12598) );
  AND U12300 ( .A(n272), .B(n12597), .Z(n12607) );
  XNOR U12301 ( .A(n12608), .B(n12595), .Z(n12597) );
  XOR U12302 ( .A(n12609), .B(n12610), .Z(n12595) );
  AND U12303 ( .A(n295), .B(n12611), .Z(n12610) );
  IV U12304 ( .A(n12606), .Z(n12608) );
  XOR U12305 ( .A(n12612), .B(n12613), .Z(n12606) );
  AND U12306 ( .A(n279), .B(n12605), .Z(n12613) );
  XNOR U12307 ( .A(n12603), .B(n12612), .Z(n12605) );
  XNOR U12308 ( .A(n12614), .B(n12615), .Z(n12603) );
  AND U12309 ( .A(n283), .B(n12616), .Z(n12615) );
  XOR U12310 ( .A(p_input[281]), .B(n12614), .Z(n12616) );
  XNOR U12311 ( .A(n12617), .B(n12618), .Z(n12614) );
  AND U12312 ( .A(n287), .B(n12619), .Z(n12618) );
  XOR U12313 ( .A(n12620), .B(n12621), .Z(n12612) );
  AND U12314 ( .A(n291), .B(n12611), .Z(n12621) );
  XNOR U12315 ( .A(n12622), .B(n12609), .Z(n12611) );
  XOR U12316 ( .A(n12623), .B(n12624), .Z(n12609) );
  AND U12317 ( .A(n314), .B(n12625), .Z(n12624) );
  IV U12318 ( .A(n12620), .Z(n12622) );
  XOR U12319 ( .A(n12626), .B(n12627), .Z(n12620) );
  AND U12320 ( .A(n298), .B(n12619), .Z(n12627) );
  XNOR U12321 ( .A(n12617), .B(n12626), .Z(n12619) );
  XNOR U12322 ( .A(n12628), .B(n12629), .Z(n12617) );
  AND U12323 ( .A(n302), .B(n12630), .Z(n12629) );
  XOR U12324 ( .A(p_input[313]), .B(n12628), .Z(n12630) );
  XNOR U12325 ( .A(n12631), .B(n12632), .Z(n12628) );
  AND U12326 ( .A(n306), .B(n12633), .Z(n12632) );
  XOR U12327 ( .A(n12634), .B(n12635), .Z(n12626) );
  AND U12328 ( .A(n310), .B(n12625), .Z(n12635) );
  XNOR U12329 ( .A(n12636), .B(n12623), .Z(n12625) );
  XOR U12330 ( .A(n12637), .B(n12638), .Z(n12623) );
  AND U12331 ( .A(n333), .B(n12639), .Z(n12638) );
  IV U12332 ( .A(n12634), .Z(n12636) );
  XOR U12333 ( .A(n12640), .B(n12641), .Z(n12634) );
  AND U12334 ( .A(n317), .B(n12633), .Z(n12641) );
  XNOR U12335 ( .A(n12631), .B(n12640), .Z(n12633) );
  XNOR U12336 ( .A(n12642), .B(n12643), .Z(n12631) );
  AND U12337 ( .A(n321), .B(n12644), .Z(n12643) );
  XOR U12338 ( .A(p_input[345]), .B(n12642), .Z(n12644) );
  XNOR U12339 ( .A(n12645), .B(n12646), .Z(n12642) );
  AND U12340 ( .A(n325), .B(n12647), .Z(n12646) );
  XOR U12341 ( .A(n12648), .B(n12649), .Z(n12640) );
  AND U12342 ( .A(n329), .B(n12639), .Z(n12649) );
  XNOR U12343 ( .A(n12650), .B(n12637), .Z(n12639) );
  XOR U12344 ( .A(n12651), .B(n12652), .Z(n12637) );
  AND U12345 ( .A(n352), .B(n12653), .Z(n12652) );
  IV U12346 ( .A(n12648), .Z(n12650) );
  XOR U12347 ( .A(n12654), .B(n12655), .Z(n12648) );
  AND U12348 ( .A(n336), .B(n12647), .Z(n12655) );
  XNOR U12349 ( .A(n12645), .B(n12654), .Z(n12647) );
  XNOR U12350 ( .A(n12656), .B(n12657), .Z(n12645) );
  AND U12351 ( .A(n340), .B(n12658), .Z(n12657) );
  XOR U12352 ( .A(p_input[377]), .B(n12656), .Z(n12658) );
  XNOR U12353 ( .A(n12659), .B(n12660), .Z(n12656) );
  AND U12354 ( .A(n344), .B(n12661), .Z(n12660) );
  XOR U12355 ( .A(n12662), .B(n12663), .Z(n12654) );
  AND U12356 ( .A(n348), .B(n12653), .Z(n12663) );
  XNOR U12357 ( .A(n12664), .B(n12651), .Z(n12653) );
  XOR U12358 ( .A(n12665), .B(n12666), .Z(n12651) );
  AND U12359 ( .A(n371), .B(n12667), .Z(n12666) );
  IV U12360 ( .A(n12662), .Z(n12664) );
  XOR U12361 ( .A(n12668), .B(n12669), .Z(n12662) );
  AND U12362 ( .A(n355), .B(n12661), .Z(n12669) );
  XNOR U12363 ( .A(n12659), .B(n12668), .Z(n12661) );
  XNOR U12364 ( .A(n12670), .B(n12671), .Z(n12659) );
  AND U12365 ( .A(n359), .B(n12672), .Z(n12671) );
  XOR U12366 ( .A(p_input[409]), .B(n12670), .Z(n12672) );
  XNOR U12367 ( .A(n12673), .B(n12674), .Z(n12670) );
  AND U12368 ( .A(n363), .B(n12675), .Z(n12674) );
  XOR U12369 ( .A(n12676), .B(n12677), .Z(n12668) );
  AND U12370 ( .A(n367), .B(n12667), .Z(n12677) );
  XNOR U12371 ( .A(n12678), .B(n12665), .Z(n12667) );
  XOR U12372 ( .A(n12679), .B(n12680), .Z(n12665) );
  AND U12373 ( .A(n390), .B(n12681), .Z(n12680) );
  IV U12374 ( .A(n12676), .Z(n12678) );
  XOR U12375 ( .A(n12682), .B(n12683), .Z(n12676) );
  AND U12376 ( .A(n374), .B(n12675), .Z(n12683) );
  XNOR U12377 ( .A(n12673), .B(n12682), .Z(n12675) );
  XNOR U12378 ( .A(n12684), .B(n12685), .Z(n12673) );
  AND U12379 ( .A(n378), .B(n12686), .Z(n12685) );
  XOR U12380 ( .A(p_input[441]), .B(n12684), .Z(n12686) );
  XNOR U12381 ( .A(n12687), .B(n12688), .Z(n12684) );
  AND U12382 ( .A(n382), .B(n12689), .Z(n12688) );
  XOR U12383 ( .A(n12690), .B(n12691), .Z(n12682) );
  AND U12384 ( .A(n386), .B(n12681), .Z(n12691) );
  XNOR U12385 ( .A(n12692), .B(n12679), .Z(n12681) );
  XOR U12386 ( .A(n12693), .B(n12694), .Z(n12679) );
  AND U12387 ( .A(n409), .B(n12695), .Z(n12694) );
  IV U12388 ( .A(n12690), .Z(n12692) );
  XOR U12389 ( .A(n12696), .B(n12697), .Z(n12690) );
  AND U12390 ( .A(n393), .B(n12689), .Z(n12697) );
  XNOR U12391 ( .A(n12687), .B(n12696), .Z(n12689) );
  XNOR U12392 ( .A(n12698), .B(n12699), .Z(n12687) );
  AND U12393 ( .A(n397), .B(n12700), .Z(n12699) );
  XOR U12394 ( .A(p_input[473]), .B(n12698), .Z(n12700) );
  XNOR U12395 ( .A(n12701), .B(n12702), .Z(n12698) );
  AND U12396 ( .A(n401), .B(n12703), .Z(n12702) );
  XOR U12397 ( .A(n12704), .B(n12705), .Z(n12696) );
  AND U12398 ( .A(n405), .B(n12695), .Z(n12705) );
  XNOR U12399 ( .A(n12706), .B(n12693), .Z(n12695) );
  XOR U12400 ( .A(n12707), .B(n12708), .Z(n12693) );
  AND U12401 ( .A(n428), .B(n12709), .Z(n12708) );
  IV U12402 ( .A(n12704), .Z(n12706) );
  XOR U12403 ( .A(n12710), .B(n12711), .Z(n12704) );
  AND U12404 ( .A(n412), .B(n12703), .Z(n12711) );
  XNOR U12405 ( .A(n12701), .B(n12710), .Z(n12703) );
  XNOR U12406 ( .A(n12712), .B(n12713), .Z(n12701) );
  AND U12407 ( .A(n416), .B(n12714), .Z(n12713) );
  XOR U12408 ( .A(p_input[505]), .B(n12712), .Z(n12714) );
  XNOR U12409 ( .A(n12715), .B(n12716), .Z(n12712) );
  AND U12410 ( .A(n420), .B(n12717), .Z(n12716) );
  XOR U12411 ( .A(n12718), .B(n12719), .Z(n12710) );
  AND U12412 ( .A(n424), .B(n12709), .Z(n12719) );
  XNOR U12413 ( .A(n12720), .B(n12707), .Z(n12709) );
  XOR U12414 ( .A(n12721), .B(n12722), .Z(n12707) );
  AND U12415 ( .A(n447), .B(n12723), .Z(n12722) );
  IV U12416 ( .A(n12718), .Z(n12720) );
  XOR U12417 ( .A(n12724), .B(n12725), .Z(n12718) );
  AND U12418 ( .A(n431), .B(n12717), .Z(n12725) );
  XNOR U12419 ( .A(n12715), .B(n12724), .Z(n12717) );
  XNOR U12420 ( .A(n12726), .B(n12727), .Z(n12715) );
  AND U12421 ( .A(n435), .B(n12728), .Z(n12727) );
  XOR U12422 ( .A(p_input[537]), .B(n12726), .Z(n12728) );
  XNOR U12423 ( .A(n12729), .B(n12730), .Z(n12726) );
  AND U12424 ( .A(n439), .B(n12731), .Z(n12730) );
  XOR U12425 ( .A(n12732), .B(n12733), .Z(n12724) );
  AND U12426 ( .A(n443), .B(n12723), .Z(n12733) );
  XNOR U12427 ( .A(n12734), .B(n12721), .Z(n12723) );
  XOR U12428 ( .A(n12735), .B(n12736), .Z(n12721) );
  AND U12429 ( .A(n466), .B(n12737), .Z(n12736) );
  IV U12430 ( .A(n12732), .Z(n12734) );
  XOR U12431 ( .A(n12738), .B(n12739), .Z(n12732) );
  AND U12432 ( .A(n450), .B(n12731), .Z(n12739) );
  XNOR U12433 ( .A(n12729), .B(n12738), .Z(n12731) );
  XNOR U12434 ( .A(n12740), .B(n12741), .Z(n12729) );
  AND U12435 ( .A(n454), .B(n12742), .Z(n12741) );
  XOR U12436 ( .A(p_input[569]), .B(n12740), .Z(n12742) );
  XNOR U12437 ( .A(n12743), .B(n12744), .Z(n12740) );
  AND U12438 ( .A(n458), .B(n12745), .Z(n12744) );
  XOR U12439 ( .A(n12746), .B(n12747), .Z(n12738) );
  AND U12440 ( .A(n462), .B(n12737), .Z(n12747) );
  XNOR U12441 ( .A(n12748), .B(n12735), .Z(n12737) );
  XOR U12442 ( .A(n12749), .B(n12750), .Z(n12735) );
  AND U12443 ( .A(n485), .B(n12751), .Z(n12750) );
  IV U12444 ( .A(n12746), .Z(n12748) );
  XOR U12445 ( .A(n12752), .B(n12753), .Z(n12746) );
  AND U12446 ( .A(n469), .B(n12745), .Z(n12753) );
  XNOR U12447 ( .A(n12743), .B(n12752), .Z(n12745) );
  XNOR U12448 ( .A(n12754), .B(n12755), .Z(n12743) );
  AND U12449 ( .A(n473), .B(n12756), .Z(n12755) );
  XOR U12450 ( .A(p_input[601]), .B(n12754), .Z(n12756) );
  XNOR U12451 ( .A(n12757), .B(n12758), .Z(n12754) );
  AND U12452 ( .A(n477), .B(n12759), .Z(n12758) );
  XOR U12453 ( .A(n12760), .B(n12761), .Z(n12752) );
  AND U12454 ( .A(n481), .B(n12751), .Z(n12761) );
  XNOR U12455 ( .A(n12762), .B(n12749), .Z(n12751) );
  XOR U12456 ( .A(n12763), .B(n12764), .Z(n12749) );
  AND U12457 ( .A(n504), .B(n12765), .Z(n12764) );
  IV U12458 ( .A(n12760), .Z(n12762) );
  XOR U12459 ( .A(n12766), .B(n12767), .Z(n12760) );
  AND U12460 ( .A(n488), .B(n12759), .Z(n12767) );
  XNOR U12461 ( .A(n12757), .B(n12766), .Z(n12759) );
  XNOR U12462 ( .A(n12768), .B(n12769), .Z(n12757) );
  AND U12463 ( .A(n492), .B(n12770), .Z(n12769) );
  XOR U12464 ( .A(p_input[633]), .B(n12768), .Z(n12770) );
  XNOR U12465 ( .A(n12771), .B(n12772), .Z(n12768) );
  AND U12466 ( .A(n496), .B(n12773), .Z(n12772) );
  XOR U12467 ( .A(n12774), .B(n12775), .Z(n12766) );
  AND U12468 ( .A(n500), .B(n12765), .Z(n12775) );
  XNOR U12469 ( .A(n12776), .B(n12763), .Z(n12765) );
  XOR U12470 ( .A(n12777), .B(n12778), .Z(n12763) );
  AND U12471 ( .A(n523), .B(n12779), .Z(n12778) );
  IV U12472 ( .A(n12774), .Z(n12776) );
  XOR U12473 ( .A(n12780), .B(n12781), .Z(n12774) );
  AND U12474 ( .A(n507), .B(n12773), .Z(n12781) );
  XNOR U12475 ( .A(n12771), .B(n12780), .Z(n12773) );
  XNOR U12476 ( .A(n12782), .B(n12783), .Z(n12771) );
  AND U12477 ( .A(n511), .B(n12784), .Z(n12783) );
  XOR U12478 ( .A(p_input[665]), .B(n12782), .Z(n12784) );
  XNOR U12479 ( .A(n12785), .B(n12786), .Z(n12782) );
  AND U12480 ( .A(n515), .B(n12787), .Z(n12786) );
  XOR U12481 ( .A(n12788), .B(n12789), .Z(n12780) );
  AND U12482 ( .A(n519), .B(n12779), .Z(n12789) );
  XNOR U12483 ( .A(n12790), .B(n12777), .Z(n12779) );
  XOR U12484 ( .A(n12791), .B(n12792), .Z(n12777) );
  AND U12485 ( .A(n542), .B(n12793), .Z(n12792) );
  IV U12486 ( .A(n12788), .Z(n12790) );
  XOR U12487 ( .A(n12794), .B(n12795), .Z(n12788) );
  AND U12488 ( .A(n526), .B(n12787), .Z(n12795) );
  XNOR U12489 ( .A(n12785), .B(n12794), .Z(n12787) );
  XNOR U12490 ( .A(n12796), .B(n12797), .Z(n12785) );
  AND U12491 ( .A(n530), .B(n12798), .Z(n12797) );
  XOR U12492 ( .A(p_input[697]), .B(n12796), .Z(n12798) );
  XNOR U12493 ( .A(n12799), .B(n12800), .Z(n12796) );
  AND U12494 ( .A(n534), .B(n12801), .Z(n12800) );
  XOR U12495 ( .A(n12802), .B(n12803), .Z(n12794) );
  AND U12496 ( .A(n538), .B(n12793), .Z(n12803) );
  XNOR U12497 ( .A(n12804), .B(n12791), .Z(n12793) );
  XOR U12498 ( .A(n12805), .B(n12806), .Z(n12791) );
  AND U12499 ( .A(n561), .B(n12807), .Z(n12806) );
  IV U12500 ( .A(n12802), .Z(n12804) );
  XOR U12501 ( .A(n12808), .B(n12809), .Z(n12802) );
  AND U12502 ( .A(n545), .B(n12801), .Z(n12809) );
  XNOR U12503 ( .A(n12799), .B(n12808), .Z(n12801) );
  XNOR U12504 ( .A(n12810), .B(n12811), .Z(n12799) );
  AND U12505 ( .A(n549), .B(n12812), .Z(n12811) );
  XOR U12506 ( .A(p_input[729]), .B(n12810), .Z(n12812) );
  XNOR U12507 ( .A(n12813), .B(n12814), .Z(n12810) );
  AND U12508 ( .A(n553), .B(n12815), .Z(n12814) );
  XOR U12509 ( .A(n12816), .B(n12817), .Z(n12808) );
  AND U12510 ( .A(n557), .B(n12807), .Z(n12817) );
  XNOR U12511 ( .A(n12818), .B(n12805), .Z(n12807) );
  XOR U12512 ( .A(n12819), .B(n12820), .Z(n12805) );
  AND U12513 ( .A(n580), .B(n12821), .Z(n12820) );
  IV U12514 ( .A(n12816), .Z(n12818) );
  XOR U12515 ( .A(n12822), .B(n12823), .Z(n12816) );
  AND U12516 ( .A(n564), .B(n12815), .Z(n12823) );
  XNOR U12517 ( .A(n12813), .B(n12822), .Z(n12815) );
  XNOR U12518 ( .A(n12824), .B(n12825), .Z(n12813) );
  AND U12519 ( .A(n568), .B(n12826), .Z(n12825) );
  XOR U12520 ( .A(p_input[761]), .B(n12824), .Z(n12826) );
  XNOR U12521 ( .A(n12827), .B(n12828), .Z(n12824) );
  AND U12522 ( .A(n572), .B(n12829), .Z(n12828) );
  XOR U12523 ( .A(n12830), .B(n12831), .Z(n12822) );
  AND U12524 ( .A(n576), .B(n12821), .Z(n12831) );
  XNOR U12525 ( .A(n12832), .B(n12819), .Z(n12821) );
  XOR U12526 ( .A(n12833), .B(n12834), .Z(n12819) );
  AND U12527 ( .A(n599), .B(n12835), .Z(n12834) );
  IV U12528 ( .A(n12830), .Z(n12832) );
  XOR U12529 ( .A(n12836), .B(n12837), .Z(n12830) );
  AND U12530 ( .A(n583), .B(n12829), .Z(n12837) );
  XNOR U12531 ( .A(n12827), .B(n12836), .Z(n12829) );
  XNOR U12532 ( .A(n12838), .B(n12839), .Z(n12827) );
  AND U12533 ( .A(n587), .B(n12840), .Z(n12839) );
  XOR U12534 ( .A(p_input[793]), .B(n12838), .Z(n12840) );
  XNOR U12535 ( .A(n12841), .B(n12842), .Z(n12838) );
  AND U12536 ( .A(n591), .B(n12843), .Z(n12842) );
  XOR U12537 ( .A(n12844), .B(n12845), .Z(n12836) );
  AND U12538 ( .A(n595), .B(n12835), .Z(n12845) );
  XNOR U12539 ( .A(n12846), .B(n12833), .Z(n12835) );
  XOR U12540 ( .A(n12847), .B(n12848), .Z(n12833) );
  AND U12541 ( .A(n618), .B(n12849), .Z(n12848) );
  IV U12542 ( .A(n12844), .Z(n12846) );
  XOR U12543 ( .A(n12850), .B(n12851), .Z(n12844) );
  AND U12544 ( .A(n602), .B(n12843), .Z(n12851) );
  XNOR U12545 ( .A(n12841), .B(n12850), .Z(n12843) );
  XNOR U12546 ( .A(n12852), .B(n12853), .Z(n12841) );
  AND U12547 ( .A(n606), .B(n12854), .Z(n12853) );
  XOR U12548 ( .A(p_input[825]), .B(n12852), .Z(n12854) );
  XNOR U12549 ( .A(n12855), .B(n12856), .Z(n12852) );
  AND U12550 ( .A(n610), .B(n12857), .Z(n12856) );
  XOR U12551 ( .A(n12858), .B(n12859), .Z(n12850) );
  AND U12552 ( .A(n614), .B(n12849), .Z(n12859) );
  XNOR U12553 ( .A(n12860), .B(n12847), .Z(n12849) );
  XOR U12554 ( .A(n12861), .B(n12862), .Z(n12847) );
  AND U12555 ( .A(n637), .B(n12863), .Z(n12862) );
  IV U12556 ( .A(n12858), .Z(n12860) );
  XOR U12557 ( .A(n12864), .B(n12865), .Z(n12858) );
  AND U12558 ( .A(n621), .B(n12857), .Z(n12865) );
  XNOR U12559 ( .A(n12855), .B(n12864), .Z(n12857) );
  XNOR U12560 ( .A(n12866), .B(n12867), .Z(n12855) );
  AND U12561 ( .A(n625), .B(n12868), .Z(n12867) );
  XOR U12562 ( .A(p_input[857]), .B(n12866), .Z(n12868) );
  XNOR U12563 ( .A(n12869), .B(n12870), .Z(n12866) );
  AND U12564 ( .A(n629), .B(n12871), .Z(n12870) );
  XOR U12565 ( .A(n12872), .B(n12873), .Z(n12864) );
  AND U12566 ( .A(n633), .B(n12863), .Z(n12873) );
  XNOR U12567 ( .A(n12874), .B(n12861), .Z(n12863) );
  XOR U12568 ( .A(n12875), .B(n12876), .Z(n12861) );
  AND U12569 ( .A(n656), .B(n12877), .Z(n12876) );
  IV U12570 ( .A(n12872), .Z(n12874) );
  XOR U12571 ( .A(n12878), .B(n12879), .Z(n12872) );
  AND U12572 ( .A(n640), .B(n12871), .Z(n12879) );
  XNOR U12573 ( .A(n12869), .B(n12878), .Z(n12871) );
  XNOR U12574 ( .A(n12880), .B(n12881), .Z(n12869) );
  AND U12575 ( .A(n644), .B(n12882), .Z(n12881) );
  XOR U12576 ( .A(p_input[889]), .B(n12880), .Z(n12882) );
  XNOR U12577 ( .A(n12883), .B(n12884), .Z(n12880) );
  AND U12578 ( .A(n648), .B(n12885), .Z(n12884) );
  XOR U12579 ( .A(n12886), .B(n12887), .Z(n12878) );
  AND U12580 ( .A(n652), .B(n12877), .Z(n12887) );
  XNOR U12581 ( .A(n12888), .B(n12875), .Z(n12877) );
  XOR U12582 ( .A(n12889), .B(n12890), .Z(n12875) );
  AND U12583 ( .A(n675), .B(n12891), .Z(n12890) );
  IV U12584 ( .A(n12886), .Z(n12888) );
  XOR U12585 ( .A(n12892), .B(n12893), .Z(n12886) );
  AND U12586 ( .A(n659), .B(n12885), .Z(n12893) );
  XNOR U12587 ( .A(n12883), .B(n12892), .Z(n12885) );
  XNOR U12588 ( .A(n12894), .B(n12895), .Z(n12883) );
  AND U12589 ( .A(n663), .B(n12896), .Z(n12895) );
  XOR U12590 ( .A(p_input[921]), .B(n12894), .Z(n12896) );
  XNOR U12591 ( .A(n12897), .B(n12898), .Z(n12894) );
  AND U12592 ( .A(n667), .B(n12899), .Z(n12898) );
  XOR U12593 ( .A(n12900), .B(n12901), .Z(n12892) );
  AND U12594 ( .A(n671), .B(n12891), .Z(n12901) );
  XNOR U12595 ( .A(n12902), .B(n12889), .Z(n12891) );
  XOR U12596 ( .A(n12903), .B(n12904), .Z(n12889) );
  AND U12597 ( .A(n694), .B(n12905), .Z(n12904) );
  IV U12598 ( .A(n12900), .Z(n12902) );
  XOR U12599 ( .A(n12906), .B(n12907), .Z(n12900) );
  AND U12600 ( .A(n678), .B(n12899), .Z(n12907) );
  XNOR U12601 ( .A(n12897), .B(n12906), .Z(n12899) );
  XNOR U12602 ( .A(n12908), .B(n12909), .Z(n12897) );
  AND U12603 ( .A(n682), .B(n12910), .Z(n12909) );
  XOR U12604 ( .A(p_input[953]), .B(n12908), .Z(n12910) );
  XNOR U12605 ( .A(n12911), .B(n12912), .Z(n12908) );
  AND U12606 ( .A(n686), .B(n12913), .Z(n12912) );
  XOR U12607 ( .A(n12914), .B(n12915), .Z(n12906) );
  AND U12608 ( .A(n690), .B(n12905), .Z(n12915) );
  XNOR U12609 ( .A(n12916), .B(n12903), .Z(n12905) );
  XOR U12610 ( .A(n12917), .B(n12918), .Z(n12903) );
  AND U12611 ( .A(n713), .B(n12919), .Z(n12918) );
  IV U12612 ( .A(n12914), .Z(n12916) );
  XOR U12613 ( .A(n12920), .B(n12921), .Z(n12914) );
  AND U12614 ( .A(n697), .B(n12913), .Z(n12921) );
  XNOR U12615 ( .A(n12911), .B(n12920), .Z(n12913) );
  XNOR U12616 ( .A(n12922), .B(n12923), .Z(n12911) );
  AND U12617 ( .A(n701), .B(n12924), .Z(n12923) );
  XOR U12618 ( .A(p_input[985]), .B(n12922), .Z(n12924) );
  XNOR U12619 ( .A(n12925), .B(n12926), .Z(n12922) );
  AND U12620 ( .A(n705), .B(n12927), .Z(n12926) );
  XOR U12621 ( .A(n12928), .B(n12929), .Z(n12920) );
  AND U12622 ( .A(n709), .B(n12919), .Z(n12929) );
  XNOR U12623 ( .A(n12930), .B(n12917), .Z(n12919) );
  XOR U12624 ( .A(n12931), .B(n12932), .Z(n12917) );
  AND U12625 ( .A(n732), .B(n12933), .Z(n12932) );
  IV U12626 ( .A(n12928), .Z(n12930) );
  XOR U12627 ( .A(n12934), .B(n12935), .Z(n12928) );
  AND U12628 ( .A(n716), .B(n12927), .Z(n12935) );
  XNOR U12629 ( .A(n12925), .B(n12934), .Z(n12927) );
  XNOR U12630 ( .A(n12936), .B(n12937), .Z(n12925) );
  AND U12631 ( .A(n720), .B(n12938), .Z(n12937) );
  XOR U12632 ( .A(p_input[1017]), .B(n12936), .Z(n12938) );
  XNOR U12633 ( .A(n12939), .B(n12940), .Z(n12936) );
  AND U12634 ( .A(n724), .B(n12941), .Z(n12940) );
  XOR U12635 ( .A(n12942), .B(n12943), .Z(n12934) );
  AND U12636 ( .A(n728), .B(n12933), .Z(n12943) );
  XNOR U12637 ( .A(n12944), .B(n12931), .Z(n12933) );
  XOR U12638 ( .A(n12945), .B(n12946), .Z(n12931) );
  AND U12639 ( .A(n751), .B(n12947), .Z(n12946) );
  IV U12640 ( .A(n12942), .Z(n12944) );
  XOR U12641 ( .A(n12948), .B(n12949), .Z(n12942) );
  AND U12642 ( .A(n735), .B(n12941), .Z(n12949) );
  XNOR U12643 ( .A(n12939), .B(n12948), .Z(n12941) );
  XNOR U12644 ( .A(n12950), .B(n12951), .Z(n12939) );
  AND U12645 ( .A(n739), .B(n12952), .Z(n12951) );
  XOR U12646 ( .A(p_input[1049]), .B(n12950), .Z(n12952) );
  XNOR U12647 ( .A(n12953), .B(n12954), .Z(n12950) );
  AND U12648 ( .A(n743), .B(n12955), .Z(n12954) );
  XOR U12649 ( .A(n12956), .B(n12957), .Z(n12948) );
  AND U12650 ( .A(n747), .B(n12947), .Z(n12957) );
  XNOR U12651 ( .A(n12958), .B(n12945), .Z(n12947) );
  XOR U12652 ( .A(n12959), .B(n12960), .Z(n12945) );
  AND U12653 ( .A(n770), .B(n12961), .Z(n12960) );
  IV U12654 ( .A(n12956), .Z(n12958) );
  XOR U12655 ( .A(n12962), .B(n12963), .Z(n12956) );
  AND U12656 ( .A(n754), .B(n12955), .Z(n12963) );
  XNOR U12657 ( .A(n12953), .B(n12962), .Z(n12955) );
  XNOR U12658 ( .A(n12964), .B(n12965), .Z(n12953) );
  AND U12659 ( .A(n758), .B(n12966), .Z(n12965) );
  XOR U12660 ( .A(p_input[1081]), .B(n12964), .Z(n12966) );
  XNOR U12661 ( .A(n12967), .B(n12968), .Z(n12964) );
  AND U12662 ( .A(n762), .B(n12969), .Z(n12968) );
  XOR U12663 ( .A(n12970), .B(n12971), .Z(n12962) );
  AND U12664 ( .A(n766), .B(n12961), .Z(n12971) );
  XNOR U12665 ( .A(n12972), .B(n12959), .Z(n12961) );
  XOR U12666 ( .A(n12973), .B(n12974), .Z(n12959) );
  AND U12667 ( .A(n789), .B(n12975), .Z(n12974) );
  IV U12668 ( .A(n12970), .Z(n12972) );
  XOR U12669 ( .A(n12976), .B(n12977), .Z(n12970) );
  AND U12670 ( .A(n773), .B(n12969), .Z(n12977) );
  XNOR U12671 ( .A(n12967), .B(n12976), .Z(n12969) );
  XNOR U12672 ( .A(n12978), .B(n12979), .Z(n12967) );
  AND U12673 ( .A(n777), .B(n12980), .Z(n12979) );
  XOR U12674 ( .A(p_input[1113]), .B(n12978), .Z(n12980) );
  XNOR U12675 ( .A(n12981), .B(n12982), .Z(n12978) );
  AND U12676 ( .A(n781), .B(n12983), .Z(n12982) );
  XOR U12677 ( .A(n12984), .B(n12985), .Z(n12976) );
  AND U12678 ( .A(n785), .B(n12975), .Z(n12985) );
  XNOR U12679 ( .A(n12986), .B(n12973), .Z(n12975) );
  XOR U12680 ( .A(n12987), .B(n12988), .Z(n12973) );
  AND U12681 ( .A(n808), .B(n12989), .Z(n12988) );
  IV U12682 ( .A(n12984), .Z(n12986) );
  XOR U12683 ( .A(n12990), .B(n12991), .Z(n12984) );
  AND U12684 ( .A(n792), .B(n12983), .Z(n12991) );
  XNOR U12685 ( .A(n12981), .B(n12990), .Z(n12983) );
  XNOR U12686 ( .A(n12992), .B(n12993), .Z(n12981) );
  AND U12687 ( .A(n796), .B(n12994), .Z(n12993) );
  XOR U12688 ( .A(p_input[1145]), .B(n12992), .Z(n12994) );
  XNOR U12689 ( .A(n12995), .B(n12996), .Z(n12992) );
  AND U12690 ( .A(n800), .B(n12997), .Z(n12996) );
  XOR U12691 ( .A(n12998), .B(n12999), .Z(n12990) );
  AND U12692 ( .A(n804), .B(n12989), .Z(n12999) );
  XNOR U12693 ( .A(n13000), .B(n12987), .Z(n12989) );
  XOR U12694 ( .A(n13001), .B(n13002), .Z(n12987) );
  AND U12695 ( .A(n827), .B(n13003), .Z(n13002) );
  IV U12696 ( .A(n12998), .Z(n13000) );
  XOR U12697 ( .A(n13004), .B(n13005), .Z(n12998) );
  AND U12698 ( .A(n811), .B(n12997), .Z(n13005) );
  XNOR U12699 ( .A(n12995), .B(n13004), .Z(n12997) );
  XNOR U12700 ( .A(n13006), .B(n13007), .Z(n12995) );
  AND U12701 ( .A(n815), .B(n13008), .Z(n13007) );
  XOR U12702 ( .A(p_input[1177]), .B(n13006), .Z(n13008) );
  XNOR U12703 ( .A(n13009), .B(n13010), .Z(n13006) );
  AND U12704 ( .A(n819), .B(n13011), .Z(n13010) );
  XOR U12705 ( .A(n13012), .B(n13013), .Z(n13004) );
  AND U12706 ( .A(n823), .B(n13003), .Z(n13013) );
  XNOR U12707 ( .A(n13014), .B(n13001), .Z(n13003) );
  XOR U12708 ( .A(n13015), .B(n13016), .Z(n13001) );
  AND U12709 ( .A(n846), .B(n13017), .Z(n13016) );
  IV U12710 ( .A(n13012), .Z(n13014) );
  XOR U12711 ( .A(n13018), .B(n13019), .Z(n13012) );
  AND U12712 ( .A(n830), .B(n13011), .Z(n13019) );
  XNOR U12713 ( .A(n13009), .B(n13018), .Z(n13011) );
  XNOR U12714 ( .A(n13020), .B(n13021), .Z(n13009) );
  AND U12715 ( .A(n834), .B(n13022), .Z(n13021) );
  XOR U12716 ( .A(p_input[1209]), .B(n13020), .Z(n13022) );
  XNOR U12717 ( .A(n13023), .B(n13024), .Z(n13020) );
  AND U12718 ( .A(n838), .B(n13025), .Z(n13024) );
  XOR U12719 ( .A(n13026), .B(n13027), .Z(n13018) );
  AND U12720 ( .A(n842), .B(n13017), .Z(n13027) );
  XNOR U12721 ( .A(n13028), .B(n13015), .Z(n13017) );
  XOR U12722 ( .A(n13029), .B(n13030), .Z(n13015) );
  AND U12723 ( .A(n865), .B(n13031), .Z(n13030) );
  IV U12724 ( .A(n13026), .Z(n13028) );
  XOR U12725 ( .A(n13032), .B(n13033), .Z(n13026) );
  AND U12726 ( .A(n849), .B(n13025), .Z(n13033) );
  XNOR U12727 ( .A(n13023), .B(n13032), .Z(n13025) );
  XNOR U12728 ( .A(n13034), .B(n13035), .Z(n13023) );
  AND U12729 ( .A(n853), .B(n13036), .Z(n13035) );
  XOR U12730 ( .A(p_input[1241]), .B(n13034), .Z(n13036) );
  XNOR U12731 ( .A(n13037), .B(n13038), .Z(n13034) );
  AND U12732 ( .A(n857), .B(n13039), .Z(n13038) );
  XOR U12733 ( .A(n13040), .B(n13041), .Z(n13032) );
  AND U12734 ( .A(n861), .B(n13031), .Z(n13041) );
  XNOR U12735 ( .A(n13042), .B(n13029), .Z(n13031) );
  XOR U12736 ( .A(n13043), .B(n13044), .Z(n13029) );
  AND U12737 ( .A(n884), .B(n13045), .Z(n13044) );
  IV U12738 ( .A(n13040), .Z(n13042) );
  XOR U12739 ( .A(n13046), .B(n13047), .Z(n13040) );
  AND U12740 ( .A(n868), .B(n13039), .Z(n13047) );
  XNOR U12741 ( .A(n13037), .B(n13046), .Z(n13039) );
  XNOR U12742 ( .A(n13048), .B(n13049), .Z(n13037) );
  AND U12743 ( .A(n872), .B(n13050), .Z(n13049) );
  XOR U12744 ( .A(p_input[1273]), .B(n13048), .Z(n13050) );
  XNOR U12745 ( .A(n13051), .B(n13052), .Z(n13048) );
  AND U12746 ( .A(n876), .B(n13053), .Z(n13052) );
  XOR U12747 ( .A(n13054), .B(n13055), .Z(n13046) );
  AND U12748 ( .A(n880), .B(n13045), .Z(n13055) );
  XNOR U12749 ( .A(n13056), .B(n13043), .Z(n13045) );
  XOR U12750 ( .A(n13057), .B(n13058), .Z(n13043) );
  AND U12751 ( .A(n903), .B(n13059), .Z(n13058) );
  IV U12752 ( .A(n13054), .Z(n13056) );
  XOR U12753 ( .A(n13060), .B(n13061), .Z(n13054) );
  AND U12754 ( .A(n887), .B(n13053), .Z(n13061) );
  XNOR U12755 ( .A(n13051), .B(n13060), .Z(n13053) );
  XNOR U12756 ( .A(n13062), .B(n13063), .Z(n13051) );
  AND U12757 ( .A(n891), .B(n13064), .Z(n13063) );
  XOR U12758 ( .A(p_input[1305]), .B(n13062), .Z(n13064) );
  XNOR U12759 ( .A(n13065), .B(n13066), .Z(n13062) );
  AND U12760 ( .A(n895), .B(n13067), .Z(n13066) );
  XOR U12761 ( .A(n13068), .B(n13069), .Z(n13060) );
  AND U12762 ( .A(n899), .B(n13059), .Z(n13069) );
  XNOR U12763 ( .A(n13070), .B(n13057), .Z(n13059) );
  XOR U12764 ( .A(n13071), .B(n13072), .Z(n13057) );
  AND U12765 ( .A(n922), .B(n13073), .Z(n13072) );
  IV U12766 ( .A(n13068), .Z(n13070) );
  XOR U12767 ( .A(n13074), .B(n13075), .Z(n13068) );
  AND U12768 ( .A(n906), .B(n13067), .Z(n13075) );
  XNOR U12769 ( .A(n13065), .B(n13074), .Z(n13067) );
  XNOR U12770 ( .A(n13076), .B(n13077), .Z(n13065) );
  AND U12771 ( .A(n910), .B(n13078), .Z(n13077) );
  XOR U12772 ( .A(p_input[1337]), .B(n13076), .Z(n13078) );
  XNOR U12773 ( .A(n13079), .B(n13080), .Z(n13076) );
  AND U12774 ( .A(n914), .B(n13081), .Z(n13080) );
  XOR U12775 ( .A(n13082), .B(n13083), .Z(n13074) );
  AND U12776 ( .A(n918), .B(n13073), .Z(n13083) );
  XNOR U12777 ( .A(n13084), .B(n13071), .Z(n13073) );
  XOR U12778 ( .A(n13085), .B(n13086), .Z(n13071) );
  AND U12779 ( .A(n941), .B(n13087), .Z(n13086) );
  IV U12780 ( .A(n13082), .Z(n13084) );
  XOR U12781 ( .A(n13088), .B(n13089), .Z(n13082) );
  AND U12782 ( .A(n925), .B(n13081), .Z(n13089) );
  XNOR U12783 ( .A(n13079), .B(n13088), .Z(n13081) );
  XNOR U12784 ( .A(n13090), .B(n13091), .Z(n13079) );
  AND U12785 ( .A(n929), .B(n13092), .Z(n13091) );
  XOR U12786 ( .A(p_input[1369]), .B(n13090), .Z(n13092) );
  XNOR U12787 ( .A(n13093), .B(n13094), .Z(n13090) );
  AND U12788 ( .A(n933), .B(n13095), .Z(n13094) );
  XOR U12789 ( .A(n13096), .B(n13097), .Z(n13088) );
  AND U12790 ( .A(n937), .B(n13087), .Z(n13097) );
  XNOR U12791 ( .A(n13098), .B(n13085), .Z(n13087) );
  XOR U12792 ( .A(n13099), .B(n13100), .Z(n13085) );
  AND U12793 ( .A(n960), .B(n13101), .Z(n13100) );
  IV U12794 ( .A(n13096), .Z(n13098) );
  XOR U12795 ( .A(n13102), .B(n13103), .Z(n13096) );
  AND U12796 ( .A(n944), .B(n13095), .Z(n13103) );
  XNOR U12797 ( .A(n13093), .B(n13102), .Z(n13095) );
  XNOR U12798 ( .A(n13104), .B(n13105), .Z(n13093) );
  AND U12799 ( .A(n948), .B(n13106), .Z(n13105) );
  XOR U12800 ( .A(p_input[1401]), .B(n13104), .Z(n13106) );
  XNOR U12801 ( .A(n13107), .B(n13108), .Z(n13104) );
  AND U12802 ( .A(n952), .B(n13109), .Z(n13108) );
  XOR U12803 ( .A(n13110), .B(n13111), .Z(n13102) );
  AND U12804 ( .A(n956), .B(n13101), .Z(n13111) );
  XNOR U12805 ( .A(n13112), .B(n13099), .Z(n13101) );
  XOR U12806 ( .A(n13113), .B(n13114), .Z(n13099) );
  AND U12807 ( .A(n979), .B(n13115), .Z(n13114) );
  IV U12808 ( .A(n13110), .Z(n13112) );
  XOR U12809 ( .A(n13116), .B(n13117), .Z(n13110) );
  AND U12810 ( .A(n963), .B(n13109), .Z(n13117) );
  XNOR U12811 ( .A(n13107), .B(n13116), .Z(n13109) );
  XNOR U12812 ( .A(n13118), .B(n13119), .Z(n13107) );
  AND U12813 ( .A(n967), .B(n13120), .Z(n13119) );
  XOR U12814 ( .A(p_input[1433]), .B(n13118), .Z(n13120) );
  XNOR U12815 ( .A(n13121), .B(n13122), .Z(n13118) );
  AND U12816 ( .A(n971), .B(n13123), .Z(n13122) );
  XOR U12817 ( .A(n13124), .B(n13125), .Z(n13116) );
  AND U12818 ( .A(n975), .B(n13115), .Z(n13125) );
  XNOR U12819 ( .A(n13126), .B(n13113), .Z(n13115) );
  XOR U12820 ( .A(n13127), .B(n13128), .Z(n13113) );
  AND U12821 ( .A(n998), .B(n13129), .Z(n13128) );
  IV U12822 ( .A(n13124), .Z(n13126) );
  XOR U12823 ( .A(n13130), .B(n13131), .Z(n13124) );
  AND U12824 ( .A(n982), .B(n13123), .Z(n13131) );
  XNOR U12825 ( .A(n13121), .B(n13130), .Z(n13123) );
  XNOR U12826 ( .A(n13132), .B(n13133), .Z(n13121) );
  AND U12827 ( .A(n986), .B(n13134), .Z(n13133) );
  XOR U12828 ( .A(p_input[1465]), .B(n13132), .Z(n13134) );
  XNOR U12829 ( .A(n13135), .B(n13136), .Z(n13132) );
  AND U12830 ( .A(n990), .B(n13137), .Z(n13136) );
  XOR U12831 ( .A(n13138), .B(n13139), .Z(n13130) );
  AND U12832 ( .A(n994), .B(n13129), .Z(n13139) );
  XNOR U12833 ( .A(n13140), .B(n13127), .Z(n13129) );
  XOR U12834 ( .A(n13141), .B(n13142), .Z(n13127) );
  AND U12835 ( .A(n1017), .B(n13143), .Z(n13142) );
  IV U12836 ( .A(n13138), .Z(n13140) );
  XOR U12837 ( .A(n13144), .B(n13145), .Z(n13138) );
  AND U12838 ( .A(n1001), .B(n13137), .Z(n13145) );
  XNOR U12839 ( .A(n13135), .B(n13144), .Z(n13137) );
  XNOR U12840 ( .A(n13146), .B(n13147), .Z(n13135) );
  AND U12841 ( .A(n1005), .B(n13148), .Z(n13147) );
  XOR U12842 ( .A(p_input[1497]), .B(n13146), .Z(n13148) );
  XNOR U12843 ( .A(n13149), .B(n13150), .Z(n13146) );
  AND U12844 ( .A(n1009), .B(n13151), .Z(n13150) );
  XOR U12845 ( .A(n13152), .B(n13153), .Z(n13144) );
  AND U12846 ( .A(n1013), .B(n13143), .Z(n13153) );
  XNOR U12847 ( .A(n13154), .B(n13141), .Z(n13143) );
  XOR U12848 ( .A(n13155), .B(n13156), .Z(n13141) );
  AND U12849 ( .A(n1036), .B(n13157), .Z(n13156) );
  IV U12850 ( .A(n13152), .Z(n13154) );
  XOR U12851 ( .A(n13158), .B(n13159), .Z(n13152) );
  AND U12852 ( .A(n1020), .B(n13151), .Z(n13159) );
  XNOR U12853 ( .A(n13149), .B(n13158), .Z(n13151) );
  XNOR U12854 ( .A(n13160), .B(n13161), .Z(n13149) );
  AND U12855 ( .A(n1024), .B(n13162), .Z(n13161) );
  XOR U12856 ( .A(p_input[1529]), .B(n13160), .Z(n13162) );
  XNOR U12857 ( .A(n13163), .B(n13164), .Z(n13160) );
  AND U12858 ( .A(n1028), .B(n13165), .Z(n13164) );
  XOR U12859 ( .A(n13166), .B(n13167), .Z(n13158) );
  AND U12860 ( .A(n1032), .B(n13157), .Z(n13167) );
  XNOR U12861 ( .A(n13168), .B(n13155), .Z(n13157) );
  XOR U12862 ( .A(n13169), .B(n13170), .Z(n13155) );
  AND U12863 ( .A(n1055), .B(n13171), .Z(n13170) );
  IV U12864 ( .A(n13166), .Z(n13168) );
  XOR U12865 ( .A(n13172), .B(n13173), .Z(n13166) );
  AND U12866 ( .A(n1039), .B(n13165), .Z(n13173) );
  XNOR U12867 ( .A(n13163), .B(n13172), .Z(n13165) );
  XNOR U12868 ( .A(n13174), .B(n13175), .Z(n13163) );
  AND U12869 ( .A(n1043), .B(n13176), .Z(n13175) );
  XOR U12870 ( .A(p_input[1561]), .B(n13174), .Z(n13176) );
  XNOR U12871 ( .A(n13177), .B(n13178), .Z(n13174) );
  AND U12872 ( .A(n1047), .B(n13179), .Z(n13178) );
  XOR U12873 ( .A(n13180), .B(n13181), .Z(n13172) );
  AND U12874 ( .A(n1051), .B(n13171), .Z(n13181) );
  XNOR U12875 ( .A(n13182), .B(n13169), .Z(n13171) );
  XOR U12876 ( .A(n13183), .B(n13184), .Z(n13169) );
  AND U12877 ( .A(n1074), .B(n13185), .Z(n13184) );
  IV U12878 ( .A(n13180), .Z(n13182) );
  XOR U12879 ( .A(n13186), .B(n13187), .Z(n13180) );
  AND U12880 ( .A(n1058), .B(n13179), .Z(n13187) );
  XNOR U12881 ( .A(n13177), .B(n13186), .Z(n13179) );
  XNOR U12882 ( .A(n13188), .B(n13189), .Z(n13177) );
  AND U12883 ( .A(n1062), .B(n13190), .Z(n13189) );
  XOR U12884 ( .A(p_input[1593]), .B(n13188), .Z(n13190) );
  XNOR U12885 ( .A(n13191), .B(n13192), .Z(n13188) );
  AND U12886 ( .A(n1066), .B(n13193), .Z(n13192) );
  XOR U12887 ( .A(n13194), .B(n13195), .Z(n13186) );
  AND U12888 ( .A(n1070), .B(n13185), .Z(n13195) );
  XNOR U12889 ( .A(n13196), .B(n13183), .Z(n13185) );
  XOR U12890 ( .A(n13197), .B(n13198), .Z(n13183) );
  AND U12891 ( .A(n1093), .B(n13199), .Z(n13198) );
  IV U12892 ( .A(n13194), .Z(n13196) );
  XOR U12893 ( .A(n13200), .B(n13201), .Z(n13194) );
  AND U12894 ( .A(n1077), .B(n13193), .Z(n13201) );
  XNOR U12895 ( .A(n13191), .B(n13200), .Z(n13193) );
  XNOR U12896 ( .A(n13202), .B(n13203), .Z(n13191) );
  AND U12897 ( .A(n1081), .B(n13204), .Z(n13203) );
  XOR U12898 ( .A(p_input[1625]), .B(n13202), .Z(n13204) );
  XNOR U12899 ( .A(n13205), .B(n13206), .Z(n13202) );
  AND U12900 ( .A(n1085), .B(n13207), .Z(n13206) );
  XOR U12901 ( .A(n13208), .B(n13209), .Z(n13200) );
  AND U12902 ( .A(n1089), .B(n13199), .Z(n13209) );
  XNOR U12903 ( .A(n13210), .B(n13197), .Z(n13199) );
  XOR U12904 ( .A(n13211), .B(n13212), .Z(n13197) );
  AND U12905 ( .A(n1112), .B(n13213), .Z(n13212) );
  IV U12906 ( .A(n13208), .Z(n13210) );
  XOR U12907 ( .A(n13214), .B(n13215), .Z(n13208) );
  AND U12908 ( .A(n1096), .B(n13207), .Z(n13215) );
  XNOR U12909 ( .A(n13205), .B(n13214), .Z(n13207) );
  XNOR U12910 ( .A(n13216), .B(n13217), .Z(n13205) );
  AND U12911 ( .A(n1100), .B(n13218), .Z(n13217) );
  XOR U12912 ( .A(p_input[1657]), .B(n13216), .Z(n13218) );
  XNOR U12913 ( .A(n13219), .B(n13220), .Z(n13216) );
  AND U12914 ( .A(n1104), .B(n13221), .Z(n13220) );
  XOR U12915 ( .A(n13222), .B(n13223), .Z(n13214) );
  AND U12916 ( .A(n1108), .B(n13213), .Z(n13223) );
  XNOR U12917 ( .A(n13224), .B(n13211), .Z(n13213) );
  XOR U12918 ( .A(n13225), .B(n13226), .Z(n13211) );
  AND U12919 ( .A(n1131), .B(n13227), .Z(n13226) );
  IV U12920 ( .A(n13222), .Z(n13224) );
  XOR U12921 ( .A(n13228), .B(n13229), .Z(n13222) );
  AND U12922 ( .A(n1115), .B(n13221), .Z(n13229) );
  XNOR U12923 ( .A(n13219), .B(n13228), .Z(n13221) );
  XNOR U12924 ( .A(n13230), .B(n13231), .Z(n13219) );
  AND U12925 ( .A(n1119), .B(n13232), .Z(n13231) );
  XOR U12926 ( .A(p_input[1689]), .B(n13230), .Z(n13232) );
  XNOR U12927 ( .A(n13233), .B(n13234), .Z(n13230) );
  AND U12928 ( .A(n1123), .B(n13235), .Z(n13234) );
  XOR U12929 ( .A(n13236), .B(n13237), .Z(n13228) );
  AND U12930 ( .A(n1127), .B(n13227), .Z(n13237) );
  XNOR U12931 ( .A(n13238), .B(n13225), .Z(n13227) );
  XOR U12932 ( .A(n13239), .B(n13240), .Z(n13225) );
  AND U12933 ( .A(n1150), .B(n13241), .Z(n13240) );
  IV U12934 ( .A(n13236), .Z(n13238) );
  XOR U12935 ( .A(n13242), .B(n13243), .Z(n13236) );
  AND U12936 ( .A(n1134), .B(n13235), .Z(n13243) );
  XNOR U12937 ( .A(n13233), .B(n13242), .Z(n13235) );
  XNOR U12938 ( .A(n13244), .B(n13245), .Z(n13233) );
  AND U12939 ( .A(n1138), .B(n13246), .Z(n13245) );
  XOR U12940 ( .A(p_input[1721]), .B(n13244), .Z(n13246) );
  XNOR U12941 ( .A(n13247), .B(n13248), .Z(n13244) );
  AND U12942 ( .A(n1142), .B(n13249), .Z(n13248) );
  XOR U12943 ( .A(n13250), .B(n13251), .Z(n13242) );
  AND U12944 ( .A(n1146), .B(n13241), .Z(n13251) );
  XNOR U12945 ( .A(n13252), .B(n13239), .Z(n13241) );
  XOR U12946 ( .A(n13253), .B(n13254), .Z(n13239) );
  AND U12947 ( .A(n1169), .B(n13255), .Z(n13254) );
  IV U12948 ( .A(n13250), .Z(n13252) );
  XOR U12949 ( .A(n13256), .B(n13257), .Z(n13250) );
  AND U12950 ( .A(n1153), .B(n13249), .Z(n13257) );
  XNOR U12951 ( .A(n13247), .B(n13256), .Z(n13249) );
  XNOR U12952 ( .A(n13258), .B(n13259), .Z(n13247) );
  AND U12953 ( .A(n1157), .B(n13260), .Z(n13259) );
  XOR U12954 ( .A(p_input[1753]), .B(n13258), .Z(n13260) );
  XNOR U12955 ( .A(n13261), .B(n13262), .Z(n13258) );
  AND U12956 ( .A(n1161), .B(n13263), .Z(n13262) );
  XOR U12957 ( .A(n13264), .B(n13265), .Z(n13256) );
  AND U12958 ( .A(n1165), .B(n13255), .Z(n13265) );
  XNOR U12959 ( .A(n13266), .B(n13253), .Z(n13255) );
  XOR U12960 ( .A(n13267), .B(n13268), .Z(n13253) );
  AND U12961 ( .A(n1188), .B(n13269), .Z(n13268) );
  IV U12962 ( .A(n13264), .Z(n13266) );
  XOR U12963 ( .A(n13270), .B(n13271), .Z(n13264) );
  AND U12964 ( .A(n1172), .B(n13263), .Z(n13271) );
  XNOR U12965 ( .A(n13261), .B(n13270), .Z(n13263) );
  XNOR U12966 ( .A(n13272), .B(n13273), .Z(n13261) );
  AND U12967 ( .A(n1176), .B(n13274), .Z(n13273) );
  XOR U12968 ( .A(p_input[1785]), .B(n13272), .Z(n13274) );
  XNOR U12969 ( .A(n13275), .B(n13276), .Z(n13272) );
  AND U12970 ( .A(n1180), .B(n13277), .Z(n13276) );
  XOR U12971 ( .A(n13278), .B(n13279), .Z(n13270) );
  AND U12972 ( .A(n1184), .B(n13269), .Z(n13279) );
  XNOR U12973 ( .A(n13280), .B(n13267), .Z(n13269) );
  XOR U12974 ( .A(n13281), .B(n13282), .Z(n13267) );
  AND U12975 ( .A(n1207), .B(n13283), .Z(n13282) );
  IV U12976 ( .A(n13278), .Z(n13280) );
  XOR U12977 ( .A(n13284), .B(n13285), .Z(n13278) );
  AND U12978 ( .A(n1191), .B(n13277), .Z(n13285) );
  XNOR U12979 ( .A(n13275), .B(n13284), .Z(n13277) );
  XNOR U12980 ( .A(n13286), .B(n13287), .Z(n13275) );
  AND U12981 ( .A(n1195), .B(n13288), .Z(n13287) );
  XOR U12982 ( .A(p_input[1817]), .B(n13286), .Z(n13288) );
  XNOR U12983 ( .A(n13289), .B(n13290), .Z(n13286) );
  AND U12984 ( .A(n1199), .B(n13291), .Z(n13290) );
  XOR U12985 ( .A(n13292), .B(n13293), .Z(n13284) );
  AND U12986 ( .A(n1203), .B(n13283), .Z(n13293) );
  XNOR U12987 ( .A(n13294), .B(n13281), .Z(n13283) );
  XOR U12988 ( .A(n13295), .B(n13296), .Z(n13281) );
  AND U12989 ( .A(n1226), .B(n13297), .Z(n13296) );
  IV U12990 ( .A(n13292), .Z(n13294) );
  XOR U12991 ( .A(n13298), .B(n13299), .Z(n13292) );
  AND U12992 ( .A(n1210), .B(n13291), .Z(n13299) );
  XNOR U12993 ( .A(n13289), .B(n13298), .Z(n13291) );
  XNOR U12994 ( .A(n13300), .B(n13301), .Z(n13289) );
  AND U12995 ( .A(n1214), .B(n13302), .Z(n13301) );
  XOR U12996 ( .A(p_input[1849]), .B(n13300), .Z(n13302) );
  XNOR U12997 ( .A(n13303), .B(n13304), .Z(n13300) );
  AND U12998 ( .A(n1218), .B(n13305), .Z(n13304) );
  XOR U12999 ( .A(n13306), .B(n13307), .Z(n13298) );
  AND U13000 ( .A(n1222), .B(n13297), .Z(n13307) );
  XNOR U13001 ( .A(n13308), .B(n13295), .Z(n13297) );
  XOR U13002 ( .A(n13309), .B(n13310), .Z(n13295) );
  AND U13003 ( .A(n1245), .B(n13311), .Z(n13310) );
  IV U13004 ( .A(n13306), .Z(n13308) );
  XOR U13005 ( .A(n13312), .B(n13313), .Z(n13306) );
  AND U13006 ( .A(n1229), .B(n13305), .Z(n13313) );
  XNOR U13007 ( .A(n13303), .B(n13312), .Z(n13305) );
  XNOR U13008 ( .A(n13314), .B(n13315), .Z(n13303) );
  AND U13009 ( .A(n1233), .B(n13316), .Z(n13315) );
  XOR U13010 ( .A(p_input[1881]), .B(n13314), .Z(n13316) );
  XNOR U13011 ( .A(n13317), .B(n13318), .Z(n13314) );
  AND U13012 ( .A(n1237), .B(n13319), .Z(n13318) );
  XOR U13013 ( .A(n13320), .B(n13321), .Z(n13312) );
  AND U13014 ( .A(n1241), .B(n13311), .Z(n13321) );
  XNOR U13015 ( .A(n13322), .B(n13309), .Z(n13311) );
  XOR U13016 ( .A(n13323), .B(n13324), .Z(n13309) );
  AND U13017 ( .A(n1264), .B(n13325), .Z(n13324) );
  IV U13018 ( .A(n13320), .Z(n13322) );
  XOR U13019 ( .A(n13326), .B(n13327), .Z(n13320) );
  AND U13020 ( .A(n1248), .B(n13319), .Z(n13327) );
  XNOR U13021 ( .A(n13317), .B(n13326), .Z(n13319) );
  XNOR U13022 ( .A(n13328), .B(n13329), .Z(n13317) );
  AND U13023 ( .A(n1252), .B(n13330), .Z(n13329) );
  XOR U13024 ( .A(p_input[1913]), .B(n13328), .Z(n13330) );
  XNOR U13025 ( .A(n13331), .B(n13332), .Z(n13328) );
  AND U13026 ( .A(n1256), .B(n13333), .Z(n13332) );
  XOR U13027 ( .A(n13334), .B(n13335), .Z(n13326) );
  AND U13028 ( .A(n1260), .B(n13325), .Z(n13335) );
  XNOR U13029 ( .A(n13336), .B(n13323), .Z(n13325) );
  XOR U13030 ( .A(n13337), .B(n13338), .Z(n13323) );
  AND U13031 ( .A(n1282), .B(n13339), .Z(n13338) );
  IV U13032 ( .A(n13334), .Z(n13336) );
  XOR U13033 ( .A(n13340), .B(n13341), .Z(n13334) );
  AND U13034 ( .A(n1267), .B(n13333), .Z(n13341) );
  XNOR U13035 ( .A(n13331), .B(n13340), .Z(n13333) );
  XNOR U13036 ( .A(n13342), .B(n13343), .Z(n13331) );
  AND U13037 ( .A(n1271), .B(n13344), .Z(n13343) );
  XOR U13038 ( .A(p_input[1945]), .B(n13342), .Z(n13344) );
  XOR U13039 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][25] ), .B(n13345), 
        .Z(n13342) );
  AND U13040 ( .A(n1274), .B(n13346), .Z(n13345) );
  XOR U13041 ( .A(n13347), .B(n13348), .Z(n13340) );
  AND U13042 ( .A(n1278), .B(n13339), .Z(n13348) );
  XNOR U13043 ( .A(n13349), .B(n13337), .Z(n13339) );
  XOR U13044 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n13350), .Z(n13337) );
  AND U13045 ( .A(n1290), .B(n13351), .Z(n13350) );
  IV U13046 ( .A(n13347), .Z(n13349) );
  XOR U13047 ( .A(n13352), .B(n13353), .Z(n13347) );
  AND U13048 ( .A(n1285), .B(n13346), .Z(n13353) );
  XOR U13049 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][25] ), .B(n13352), 
        .Z(n13346) );
  XOR U13050 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .B(n13354), 
        .Z(n13352) );
  AND U13051 ( .A(n1287), .B(n13351), .Z(n13354) );
  XOR U13052 ( .A(\knn_comb_/min_val_out[0][25] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .Z(n13351) );
  XOR U13053 ( .A(n89), .B(n13355), .Z(o[24]) );
  AND U13054 ( .A(n122), .B(n13356), .Z(n89) );
  XOR U13055 ( .A(n90), .B(n13355), .Z(n13356) );
  XOR U13056 ( .A(n13357), .B(n13358), .Z(n13355) );
  AND U13057 ( .A(n142), .B(n13359), .Z(n13358) );
  XOR U13058 ( .A(n13360), .B(n19), .Z(n90) );
  AND U13059 ( .A(n125), .B(n13361), .Z(n19) );
  XOR U13060 ( .A(n20), .B(n13360), .Z(n13361) );
  XOR U13061 ( .A(n13362), .B(n13363), .Z(n20) );
  AND U13062 ( .A(n130), .B(n13364), .Z(n13363) );
  XOR U13063 ( .A(p_input[24]), .B(n13362), .Z(n13364) );
  XNOR U13064 ( .A(n13365), .B(n13366), .Z(n13362) );
  AND U13065 ( .A(n134), .B(n13367), .Z(n13366) );
  XOR U13066 ( .A(n13368), .B(n13369), .Z(n13360) );
  AND U13067 ( .A(n138), .B(n13359), .Z(n13369) );
  XNOR U13068 ( .A(n13370), .B(n13357), .Z(n13359) );
  XOR U13069 ( .A(n13371), .B(n13372), .Z(n13357) );
  AND U13070 ( .A(n162), .B(n13373), .Z(n13372) );
  IV U13071 ( .A(n13368), .Z(n13370) );
  XOR U13072 ( .A(n13374), .B(n13375), .Z(n13368) );
  AND U13073 ( .A(n146), .B(n13367), .Z(n13375) );
  XNOR U13074 ( .A(n13365), .B(n13374), .Z(n13367) );
  XNOR U13075 ( .A(n13376), .B(n13377), .Z(n13365) );
  AND U13076 ( .A(n150), .B(n13378), .Z(n13377) );
  XOR U13077 ( .A(p_input[56]), .B(n13376), .Z(n13378) );
  XNOR U13078 ( .A(n13379), .B(n13380), .Z(n13376) );
  AND U13079 ( .A(n154), .B(n13381), .Z(n13380) );
  XOR U13080 ( .A(n13382), .B(n13383), .Z(n13374) );
  AND U13081 ( .A(n158), .B(n13373), .Z(n13383) );
  XNOR U13082 ( .A(n13384), .B(n13371), .Z(n13373) );
  XOR U13083 ( .A(n13385), .B(n13386), .Z(n13371) );
  AND U13084 ( .A(n181), .B(n13387), .Z(n13386) );
  IV U13085 ( .A(n13382), .Z(n13384) );
  XOR U13086 ( .A(n13388), .B(n13389), .Z(n13382) );
  AND U13087 ( .A(n165), .B(n13381), .Z(n13389) );
  XNOR U13088 ( .A(n13379), .B(n13388), .Z(n13381) );
  XNOR U13089 ( .A(n13390), .B(n13391), .Z(n13379) );
  AND U13090 ( .A(n169), .B(n13392), .Z(n13391) );
  XOR U13091 ( .A(p_input[88]), .B(n13390), .Z(n13392) );
  XNOR U13092 ( .A(n13393), .B(n13394), .Z(n13390) );
  AND U13093 ( .A(n173), .B(n13395), .Z(n13394) );
  XOR U13094 ( .A(n13396), .B(n13397), .Z(n13388) );
  AND U13095 ( .A(n177), .B(n13387), .Z(n13397) );
  XNOR U13096 ( .A(n13398), .B(n13385), .Z(n13387) );
  XOR U13097 ( .A(n13399), .B(n13400), .Z(n13385) );
  AND U13098 ( .A(n200), .B(n13401), .Z(n13400) );
  IV U13099 ( .A(n13396), .Z(n13398) );
  XOR U13100 ( .A(n13402), .B(n13403), .Z(n13396) );
  AND U13101 ( .A(n184), .B(n13395), .Z(n13403) );
  XNOR U13102 ( .A(n13393), .B(n13402), .Z(n13395) );
  XNOR U13103 ( .A(n13404), .B(n13405), .Z(n13393) );
  AND U13104 ( .A(n188), .B(n13406), .Z(n13405) );
  XOR U13105 ( .A(p_input[120]), .B(n13404), .Z(n13406) );
  XNOR U13106 ( .A(n13407), .B(n13408), .Z(n13404) );
  AND U13107 ( .A(n192), .B(n13409), .Z(n13408) );
  XOR U13108 ( .A(n13410), .B(n13411), .Z(n13402) );
  AND U13109 ( .A(n196), .B(n13401), .Z(n13411) );
  XNOR U13110 ( .A(n13412), .B(n13399), .Z(n13401) );
  XOR U13111 ( .A(n13413), .B(n13414), .Z(n13399) );
  AND U13112 ( .A(n219), .B(n13415), .Z(n13414) );
  IV U13113 ( .A(n13410), .Z(n13412) );
  XOR U13114 ( .A(n13416), .B(n13417), .Z(n13410) );
  AND U13115 ( .A(n203), .B(n13409), .Z(n13417) );
  XNOR U13116 ( .A(n13407), .B(n13416), .Z(n13409) );
  XNOR U13117 ( .A(n13418), .B(n13419), .Z(n13407) );
  AND U13118 ( .A(n207), .B(n13420), .Z(n13419) );
  XOR U13119 ( .A(p_input[152]), .B(n13418), .Z(n13420) );
  XNOR U13120 ( .A(n13421), .B(n13422), .Z(n13418) );
  AND U13121 ( .A(n211), .B(n13423), .Z(n13422) );
  XOR U13122 ( .A(n13424), .B(n13425), .Z(n13416) );
  AND U13123 ( .A(n215), .B(n13415), .Z(n13425) );
  XNOR U13124 ( .A(n13426), .B(n13413), .Z(n13415) );
  XOR U13125 ( .A(n13427), .B(n13428), .Z(n13413) );
  AND U13126 ( .A(n238), .B(n13429), .Z(n13428) );
  IV U13127 ( .A(n13424), .Z(n13426) );
  XOR U13128 ( .A(n13430), .B(n13431), .Z(n13424) );
  AND U13129 ( .A(n222), .B(n13423), .Z(n13431) );
  XNOR U13130 ( .A(n13421), .B(n13430), .Z(n13423) );
  XNOR U13131 ( .A(n13432), .B(n13433), .Z(n13421) );
  AND U13132 ( .A(n226), .B(n13434), .Z(n13433) );
  XOR U13133 ( .A(p_input[184]), .B(n13432), .Z(n13434) );
  XNOR U13134 ( .A(n13435), .B(n13436), .Z(n13432) );
  AND U13135 ( .A(n230), .B(n13437), .Z(n13436) );
  XOR U13136 ( .A(n13438), .B(n13439), .Z(n13430) );
  AND U13137 ( .A(n234), .B(n13429), .Z(n13439) );
  XNOR U13138 ( .A(n13440), .B(n13427), .Z(n13429) );
  XOR U13139 ( .A(n13441), .B(n13442), .Z(n13427) );
  AND U13140 ( .A(n257), .B(n13443), .Z(n13442) );
  IV U13141 ( .A(n13438), .Z(n13440) );
  XOR U13142 ( .A(n13444), .B(n13445), .Z(n13438) );
  AND U13143 ( .A(n241), .B(n13437), .Z(n13445) );
  XNOR U13144 ( .A(n13435), .B(n13444), .Z(n13437) );
  XNOR U13145 ( .A(n13446), .B(n13447), .Z(n13435) );
  AND U13146 ( .A(n245), .B(n13448), .Z(n13447) );
  XOR U13147 ( .A(p_input[216]), .B(n13446), .Z(n13448) );
  XNOR U13148 ( .A(n13449), .B(n13450), .Z(n13446) );
  AND U13149 ( .A(n249), .B(n13451), .Z(n13450) );
  XOR U13150 ( .A(n13452), .B(n13453), .Z(n13444) );
  AND U13151 ( .A(n253), .B(n13443), .Z(n13453) );
  XNOR U13152 ( .A(n13454), .B(n13441), .Z(n13443) );
  XOR U13153 ( .A(n13455), .B(n13456), .Z(n13441) );
  AND U13154 ( .A(n276), .B(n13457), .Z(n13456) );
  IV U13155 ( .A(n13452), .Z(n13454) );
  XOR U13156 ( .A(n13458), .B(n13459), .Z(n13452) );
  AND U13157 ( .A(n260), .B(n13451), .Z(n13459) );
  XNOR U13158 ( .A(n13449), .B(n13458), .Z(n13451) );
  XNOR U13159 ( .A(n13460), .B(n13461), .Z(n13449) );
  AND U13160 ( .A(n264), .B(n13462), .Z(n13461) );
  XOR U13161 ( .A(p_input[248]), .B(n13460), .Z(n13462) );
  XNOR U13162 ( .A(n13463), .B(n13464), .Z(n13460) );
  AND U13163 ( .A(n268), .B(n13465), .Z(n13464) );
  XOR U13164 ( .A(n13466), .B(n13467), .Z(n13458) );
  AND U13165 ( .A(n272), .B(n13457), .Z(n13467) );
  XNOR U13166 ( .A(n13468), .B(n13455), .Z(n13457) );
  XOR U13167 ( .A(n13469), .B(n13470), .Z(n13455) );
  AND U13168 ( .A(n295), .B(n13471), .Z(n13470) );
  IV U13169 ( .A(n13466), .Z(n13468) );
  XOR U13170 ( .A(n13472), .B(n13473), .Z(n13466) );
  AND U13171 ( .A(n279), .B(n13465), .Z(n13473) );
  XNOR U13172 ( .A(n13463), .B(n13472), .Z(n13465) );
  XNOR U13173 ( .A(n13474), .B(n13475), .Z(n13463) );
  AND U13174 ( .A(n283), .B(n13476), .Z(n13475) );
  XOR U13175 ( .A(p_input[280]), .B(n13474), .Z(n13476) );
  XNOR U13176 ( .A(n13477), .B(n13478), .Z(n13474) );
  AND U13177 ( .A(n287), .B(n13479), .Z(n13478) );
  XOR U13178 ( .A(n13480), .B(n13481), .Z(n13472) );
  AND U13179 ( .A(n291), .B(n13471), .Z(n13481) );
  XNOR U13180 ( .A(n13482), .B(n13469), .Z(n13471) );
  XOR U13181 ( .A(n13483), .B(n13484), .Z(n13469) );
  AND U13182 ( .A(n314), .B(n13485), .Z(n13484) );
  IV U13183 ( .A(n13480), .Z(n13482) );
  XOR U13184 ( .A(n13486), .B(n13487), .Z(n13480) );
  AND U13185 ( .A(n298), .B(n13479), .Z(n13487) );
  XNOR U13186 ( .A(n13477), .B(n13486), .Z(n13479) );
  XNOR U13187 ( .A(n13488), .B(n13489), .Z(n13477) );
  AND U13188 ( .A(n302), .B(n13490), .Z(n13489) );
  XOR U13189 ( .A(p_input[312]), .B(n13488), .Z(n13490) );
  XNOR U13190 ( .A(n13491), .B(n13492), .Z(n13488) );
  AND U13191 ( .A(n306), .B(n13493), .Z(n13492) );
  XOR U13192 ( .A(n13494), .B(n13495), .Z(n13486) );
  AND U13193 ( .A(n310), .B(n13485), .Z(n13495) );
  XNOR U13194 ( .A(n13496), .B(n13483), .Z(n13485) );
  XOR U13195 ( .A(n13497), .B(n13498), .Z(n13483) );
  AND U13196 ( .A(n333), .B(n13499), .Z(n13498) );
  IV U13197 ( .A(n13494), .Z(n13496) );
  XOR U13198 ( .A(n13500), .B(n13501), .Z(n13494) );
  AND U13199 ( .A(n317), .B(n13493), .Z(n13501) );
  XNOR U13200 ( .A(n13491), .B(n13500), .Z(n13493) );
  XNOR U13201 ( .A(n13502), .B(n13503), .Z(n13491) );
  AND U13202 ( .A(n321), .B(n13504), .Z(n13503) );
  XOR U13203 ( .A(p_input[344]), .B(n13502), .Z(n13504) );
  XNOR U13204 ( .A(n13505), .B(n13506), .Z(n13502) );
  AND U13205 ( .A(n325), .B(n13507), .Z(n13506) );
  XOR U13206 ( .A(n13508), .B(n13509), .Z(n13500) );
  AND U13207 ( .A(n329), .B(n13499), .Z(n13509) );
  XNOR U13208 ( .A(n13510), .B(n13497), .Z(n13499) );
  XOR U13209 ( .A(n13511), .B(n13512), .Z(n13497) );
  AND U13210 ( .A(n352), .B(n13513), .Z(n13512) );
  IV U13211 ( .A(n13508), .Z(n13510) );
  XOR U13212 ( .A(n13514), .B(n13515), .Z(n13508) );
  AND U13213 ( .A(n336), .B(n13507), .Z(n13515) );
  XNOR U13214 ( .A(n13505), .B(n13514), .Z(n13507) );
  XNOR U13215 ( .A(n13516), .B(n13517), .Z(n13505) );
  AND U13216 ( .A(n340), .B(n13518), .Z(n13517) );
  XOR U13217 ( .A(p_input[376]), .B(n13516), .Z(n13518) );
  XNOR U13218 ( .A(n13519), .B(n13520), .Z(n13516) );
  AND U13219 ( .A(n344), .B(n13521), .Z(n13520) );
  XOR U13220 ( .A(n13522), .B(n13523), .Z(n13514) );
  AND U13221 ( .A(n348), .B(n13513), .Z(n13523) );
  XNOR U13222 ( .A(n13524), .B(n13511), .Z(n13513) );
  XOR U13223 ( .A(n13525), .B(n13526), .Z(n13511) );
  AND U13224 ( .A(n371), .B(n13527), .Z(n13526) );
  IV U13225 ( .A(n13522), .Z(n13524) );
  XOR U13226 ( .A(n13528), .B(n13529), .Z(n13522) );
  AND U13227 ( .A(n355), .B(n13521), .Z(n13529) );
  XNOR U13228 ( .A(n13519), .B(n13528), .Z(n13521) );
  XNOR U13229 ( .A(n13530), .B(n13531), .Z(n13519) );
  AND U13230 ( .A(n359), .B(n13532), .Z(n13531) );
  XOR U13231 ( .A(p_input[408]), .B(n13530), .Z(n13532) );
  XNOR U13232 ( .A(n13533), .B(n13534), .Z(n13530) );
  AND U13233 ( .A(n363), .B(n13535), .Z(n13534) );
  XOR U13234 ( .A(n13536), .B(n13537), .Z(n13528) );
  AND U13235 ( .A(n367), .B(n13527), .Z(n13537) );
  XNOR U13236 ( .A(n13538), .B(n13525), .Z(n13527) );
  XOR U13237 ( .A(n13539), .B(n13540), .Z(n13525) );
  AND U13238 ( .A(n390), .B(n13541), .Z(n13540) );
  IV U13239 ( .A(n13536), .Z(n13538) );
  XOR U13240 ( .A(n13542), .B(n13543), .Z(n13536) );
  AND U13241 ( .A(n374), .B(n13535), .Z(n13543) );
  XNOR U13242 ( .A(n13533), .B(n13542), .Z(n13535) );
  XNOR U13243 ( .A(n13544), .B(n13545), .Z(n13533) );
  AND U13244 ( .A(n378), .B(n13546), .Z(n13545) );
  XOR U13245 ( .A(p_input[440]), .B(n13544), .Z(n13546) );
  XNOR U13246 ( .A(n13547), .B(n13548), .Z(n13544) );
  AND U13247 ( .A(n382), .B(n13549), .Z(n13548) );
  XOR U13248 ( .A(n13550), .B(n13551), .Z(n13542) );
  AND U13249 ( .A(n386), .B(n13541), .Z(n13551) );
  XNOR U13250 ( .A(n13552), .B(n13539), .Z(n13541) );
  XOR U13251 ( .A(n13553), .B(n13554), .Z(n13539) );
  AND U13252 ( .A(n409), .B(n13555), .Z(n13554) );
  IV U13253 ( .A(n13550), .Z(n13552) );
  XOR U13254 ( .A(n13556), .B(n13557), .Z(n13550) );
  AND U13255 ( .A(n393), .B(n13549), .Z(n13557) );
  XNOR U13256 ( .A(n13547), .B(n13556), .Z(n13549) );
  XNOR U13257 ( .A(n13558), .B(n13559), .Z(n13547) );
  AND U13258 ( .A(n397), .B(n13560), .Z(n13559) );
  XOR U13259 ( .A(p_input[472]), .B(n13558), .Z(n13560) );
  XNOR U13260 ( .A(n13561), .B(n13562), .Z(n13558) );
  AND U13261 ( .A(n401), .B(n13563), .Z(n13562) );
  XOR U13262 ( .A(n13564), .B(n13565), .Z(n13556) );
  AND U13263 ( .A(n405), .B(n13555), .Z(n13565) );
  XNOR U13264 ( .A(n13566), .B(n13553), .Z(n13555) );
  XOR U13265 ( .A(n13567), .B(n13568), .Z(n13553) );
  AND U13266 ( .A(n428), .B(n13569), .Z(n13568) );
  IV U13267 ( .A(n13564), .Z(n13566) );
  XOR U13268 ( .A(n13570), .B(n13571), .Z(n13564) );
  AND U13269 ( .A(n412), .B(n13563), .Z(n13571) );
  XNOR U13270 ( .A(n13561), .B(n13570), .Z(n13563) );
  XNOR U13271 ( .A(n13572), .B(n13573), .Z(n13561) );
  AND U13272 ( .A(n416), .B(n13574), .Z(n13573) );
  XOR U13273 ( .A(p_input[504]), .B(n13572), .Z(n13574) );
  XNOR U13274 ( .A(n13575), .B(n13576), .Z(n13572) );
  AND U13275 ( .A(n420), .B(n13577), .Z(n13576) );
  XOR U13276 ( .A(n13578), .B(n13579), .Z(n13570) );
  AND U13277 ( .A(n424), .B(n13569), .Z(n13579) );
  XNOR U13278 ( .A(n13580), .B(n13567), .Z(n13569) );
  XOR U13279 ( .A(n13581), .B(n13582), .Z(n13567) );
  AND U13280 ( .A(n447), .B(n13583), .Z(n13582) );
  IV U13281 ( .A(n13578), .Z(n13580) );
  XOR U13282 ( .A(n13584), .B(n13585), .Z(n13578) );
  AND U13283 ( .A(n431), .B(n13577), .Z(n13585) );
  XNOR U13284 ( .A(n13575), .B(n13584), .Z(n13577) );
  XNOR U13285 ( .A(n13586), .B(n13587), .Z(n13575) );
  AND U13286 ( .A(n435), .B(n13588), .Z(n13587) );
  XOR U13287 ( .A(p_input[536]), .B(n13586), .Z(n13588) );
  XNOR U13288 ( .A(n13589), .B(n13590), .Z(n13586) );
  AND U13289 ( .A(n439), .B(n13591), .Z(n13590) );
  XOR U13290 ( .A(n13592), .B(n13593), .Z(n13584) );
  AND U13291 ( .A(n443), .B(n13583), .Z(n13593) );
  XNOR U13292 ( .A(n13594), .B(n13581), .Z(n13583) );
  XOR U13293 ( .A(n13595), .B(n13596), .Z(n13581) );
  AND U13294 ( .A(n466), .B(n13597), .Z(n13596) );
  IV U13295 ( .A(n13592), .Z(n13594) );
  XOR U13296 ( .A(n13598), .B(n13599), .Z(n13592) );
  AND U13297 ( .A(n450), .B(n13591), .Z(n13599) );
  XNOR U13298 ( .A(n13589), .B(n13598), .Z(n13591) );
  XNOR U13299 ( .A(n13600), .B(n13601), .Z(n13589) );
  AND U13300 ( .A(n454), .B(n13602), .Z(n13601) );
  XOR U13301 ( .A(p_input[568]), .B(n13600), .Z(n13602) );
  XNOR U13302 ( .A(n13603), .B(n13604), .Z(n13600) );
  AND U13303 ( .A(n458), .B(n13605), .Z(n13604) );
  XOR U13304 ( .A(n13606), .B(n13607), .Z(n13598) );
  AND U13305 ( .A(n462), .B(n13597), .Z(n13607) );
  XNOR U13306 ( .A(n13608), .B(n13595), .Z(n13597) );
  XOR U13307 ( .A(n13609), .B(n13610), .Z(n13595) );
  AND U13308 ( .A(n485), .B(n13611), .Z(n13610) );
  IV U13309 ( .A(n13606), .Z(n13608) );
  XOR U13310 ( .A(n13612), .B(n13613), .Z(n13606) );
  AND U13311 ( .A(n469), .B(n13605), .Z(n13613) );
  XNOR U13312 ( .A(n13603), .B(n13612), .Z(n13605) );
  XNOR U13313 ( .A(n13614), .B(n13615), .Z(n13603) );
  AND U13314 ( .A(n473), .B(n13616), .Z(n13615) );
  XOR U13315 ( .A(p_input[600]), .B(n13614), .Z(n13616) );
  XNOR U13316 ( .A(n13617), .B(n13618), .Z(n13614) );
  AND U13317 ( .A(n477), .B(n13619), .Z(n13618) );
  XOR U13318 ( .A(n13620), .B(n13621), .Z(n13612) );
  AND U13319 ( .A(n481), .B(n13611), .Z(n13621) );
  XNOR U13320 ( .A(n13622), .B(n13609), .Z(n13611) );
  XOR U13321 ( .A(n13623), .B(n13624), .Z(n13609) );
  AND U13322 ( .A(n504), .B(n13625), .Z(n13624) );
  IV U13323 ( .A(n13620), .Z(n13622) );
  XOR U13324 ( .A(n13626), .B(n13627), .Z(n13620) );
  AND U13325 ( .A(n488), .B(n13619), .Z(n13627) );
  XNOR U13326 ( .A(n13617), .B(n13626), .Z(n13619) );
  XNOR U13327 ( .A(n13628), .B(n13629), .Z(n13617) );
  AND U13328 ( .A(n492), .B(n13630), .Z(n13629) );
  XOR U13329 ( .A(p_input[632]), .B(n13628), .Z(n13630) );
  XNOR U13330 ( .A(n13631), .B(n13632), .Z(n13628) );
  AND U13331 ( .A(n496), .B(n13633), .Z(n13632) );
  XOR U13332 ( .A(n13634), .B(n13635), .Z(n13626) );
  AND U13333 ( .A(n500), .B(n13625), .Z(n13635) );
  XNOR U13334 ( .A(n13636), .B(n13623), .Z(n13625) );
  XOR U13335 ( .A(n13637), .B(n13638), .Z(n13623) );
  AND U13336 ( .A(n523), .B(n13639), .Z(n13638) );
  IV U13337 ( .A(n13634), .Z(n13636) );
  XOR U13338 ( .A(n13640), .B(n13641), .Z(n13634) );
  AND U13339 ( .A(n507), .B(n13633), .Z(n13641) );
  XNOR U13340 ( .A(n13631), .B(n13640), .Z(n13633) );
  XNOR U13341 ( .A(n13642), .B(n13643), .Z(n13631) );
  AND U13342 ( .A(n511), .B(n13644), .Z(n13643) );
  XOR U13343 ( .A(p_input[664]), .B(n13642), .Z(n13644) );
  XNOR U13344 ( .A(n13645), .B(n13646), .Z(n13642) );
  AND U13345 ( .A(n515), .B(n13647), .Z(n13646) );
  XOR U13346 ( .A(n13648), .B(n13649), .Z(n13640) );
  AND U13347 ( .A(n519), .B(n13639), .Z(n13649) );
  XNOR U13348 ( .A(n13650), .B(n13637), .Z(n13639) );
  XOR U13349 ( .A(n13651), .B(n13652), .Z(n13637) );
  AND U13350 ( .A(n542), .B(n13653), .Z(n13652) );
  IV U13351 ( .A(n13648), .Z(n13650) );
  XOR U13352 ( .A(n13654), .B(n13655), .Z(n13648) );
  AND U13353 ( .A(n526), .B(n13647), .Z(n13655) );
  XNOR U13354 ( .A(n13645), .B(n13654), .Z(n13647) );
  XNOR U13355 ( .A(n13656), .B(n13657), .Z(n13645) );
  AND U13356 ( .A(n530), .B(n13658), .Z(n13657) );
  XOR U13357 ( .A(p_input[696]), .B(n13656), .Z(n13658) );
  XNOR U13358 ( .A(n13659), .B(n13660), .Z(n13656) );
  AND U13359 ( .A(n534), .B(n13661), .Z(n13660) );
  XOR U13360 ( .A(n13662), .B(n13663), .Z(n13654) );
  AND U13361 ( .A(n538), .B(n13653), .Z(n13663) );
  XNOR U13362 ( .A(n13664), .B(n13651), .Z(n13653) );
  XOR U13363 ( .A(n13665), .B(n13666), .Z(n13651) );
  AND U13364 ( .A(n561), .B(n13667), .Z(n13666) );
  IV U13365 ( .A(n13662), .Z(n13664) );
  XOR U13366 ( .A(n13668), .B(n13669), .Z(n13662) );
  AND U13367 ( .A(n545), .B(n13661), .Z(n13669) );
  XNOR U13368 ( .A(n13659), .B(n13668), .Z(n13661) );
  XNOR U13369 ( .A(n13670), .B(n13671), .Z(n13659) );
  AND U13370 ( .A(n549), .B(n13672), .Z(n13671) );
  XOR U13371 ( .A(p_input[728]), .B(n13670), .Z(n13672) );
  XNOR U13372 ( .A(n13673), .B(n13674), .Z(n13670) );
  AND U13373 ( .A(n553), .B(n13675), .Z(n13674) );
  XOR U13374 ( .A(n13676), .B(n13677), .Z(n13668) );
  AND U13375 ( .A(n557), .B(n13667), .Z(n13677) );
  XNOR U13376 ( .A(n13678), .B(n13665), .Z(n13667) );
  XOR U13377 ( .A(n13679), .B(n13680), .Z(n13665) );
  AND U13378 ( .A(n580), .B(n13681), .Z(n13680) );
  IV U13379 ( .A(n13676), .Z(n13678) );
  XOR U13380 ( .A(n13682), .B(n13683), .Z(n13676) );
  AND U13381 ( .A(n564), .B(n13675), .Z(n13683) );
  XNOR U13382 ( .A(n13673), .B(n13682), .Z(n13675) );
  XNOR U13383 ( .A(n13684), .B(n13685), .Z(n13673) );
  AND U13384 ( .A(n568), .B(n13686), .Z(n13685) );
  XOR U13385 ( .A(p_input[760]), .B(n13684), .Z(n13686) );
  XNOR U13386 ( .A(n13687), .B(n13688), .Z(n13684) );
  AND U13387 ( .A(n572), .B(n13689), .Z(n13688) );
  XOR U13388 ( .A(n13690), .B(n13691), .Z(n13682) );
  AND U13389 ( .A(n576), .B(n13681), .Z(n13691) );
  XNOR U13390 ( .A(n13692), .B(n13679), .Z(n13681) );
  XOR U13391 ( .A(n13693), .B(n13694), .Z(n13679) );
  AND U13392 ( .A(n599), .B(n13695), .Z(n13694) );
  IV U13393 ( .A(n13690), .Z(n13692) );
  XOR U13394 ( .A(n13696), .B(n13697), .Z(n13690) );
  AND U13395 ( .A(n583), .B(n13689), .Z(n13697) );
  XNOR U13396 ( .A(n13687), .B(n13696), .Z(n13689) );
  XNOR U13397 ( .A(n13698), .B(n13699), .Z(n13687) );
  AND U13398 ( .A(n587), .B(n13700), .Z(n13699) );
  XOR U13399 ( .A(p_input[792]), .B(n13698), .Z(n13700) );
  XNOR U13400 ( .A(n13701), .B(n13702), .Z(n13698) );
  AND U13401 ( .A(n591), .B(n13703), .Z(n13702) );
  XOR U13402 ( .A(n13704), .B(n13705), .Z(n13696) );
  AND U13403 ( .A(n595), .B(n13695), .Z(n13705) );
  XNOR U13404 ( .A(n13706), .B(n13693), .Z(n13695) );
  XOR U13405 ( .A(n13707), .B(n13708), .Z(n13693) );
  AND U13406 ( .A(n618), .B(n13709), .Z(n13708) );
  IV U13407 ( .A(n13704), .Z(n13706) );
  XOR U13408 ( .A(n13710), .B(n13711), .Z(n13704) );
  AND U13409 ( .A(n602), .B(n13703), .Z(n13711) );
  XNOR U13410 ( .A(n13701), .B(n13710), .Z(n13703) );
  XNOR U13411 ( .A(n13712), .B(n13713), .Z(n13701) );
  AND U13412 ( .A(n606), .B(n13714), .Z(n13713) );
  XOR U13413 ( .A(p_input[824]), .B(n13712), .Z(n13714) );
  XNOR U13414 ( .A(n13715), .B(n13716), .Z(n13712) );
  AND U13415 ( .A(n610), .B(n13717), .Z(n13716) );
  XOR U13416 ( .A(n13718), .B(n13719), .Z(n13710) );
  AND U13417 ( .A(n614), .B(n13709), .Z(n13719) );
  XNOR U13418 ( .A(n13720), .B(n13707), .Z(n13709) );
  XOR U13419 ( .A(n13721), .B(n13722), .Z(n13707) );
  AND U13420 ( .A(n637), .B(n13723), .Z(n13722) );
  IV U13421 ( .A(n13718), .Z(n13720) );
  XOR U13422 ( .A(n13724), .B(n13725), .Z(n13718) );
  AND U13423 ( .A(n621), .B(n13717), .Z(n13725) );
  XNOR U13424 ( .A(n13715), .B(n13724), .Z(n13717) );
  XNOR U13425 ( .A(n13726), .B(n13727), .Z(n13715) );
  AND U13426 ( .A(n625), .B(n13728), .Z(n13727) );
  XOR U13427 ( .A(p_input[856]), .B(n13726), .Z(n13728) );
  XNOR U13428 ( .A(n13729), .B(n13730), .Z(n13726) );
  AND U13429 ( .A(n629), .B(n13731), .Z(n13730) );
  XOR U13430 ( .A(n13732), .B(n13733), .Z(n13724) );
  AND U13431 ( .A(n633), .B(n13723), .Z(n13733) );
  XNOR U13432 ( .A(n13734), .B(n13721), .Z(n13723) );
  XOR U13433 ( .A(n13735), .B(n13736), .Z(n13721) );
  AND U13434 ( .A(n656), .B(n13737), .Z(n13736) );
  IV U13435 ( .A(n13732), .Z(n13734) );
  XOR U13436 ( .A(n13738), .B(n13739), .Z(n13732) );
  AND U13437 ( .A(n640), .B(n13731), .Z(n13739) );
  XNOR U13438 ( .A(n13729), .B(n13738), .Z(n13731) );
  XNOR U13439 ( .A(n13740), .B(n13741), .Z(n13729) );
  AND U13440 ( .A(n644), .B(n13742), .Z(n13741) );
  XOR U13441 ( .A(p_input[888]), .B(n13740), .Z(n13742) );
  XNOR U13442 ( .A(n13743), .B(n13744), .Z(n13740) );
  AND U13443 ( .A(n648), .B(n13745), .Z(n13744) );
  XOR U13444 ( .A(n13746), .B(n13747), .Z(n13738) );
  AND U13445 ( .A(n652), .B(n13737), .Z(n13747) );
  XNOR U13446 ( .A(n13748), .B(n13735), .Z(n13737) );
  XOR U13447 ( .A(n13749), .B(n13750), .Z(n13735) );
  AND U13448 ( .A(n675), .B(n13751), .Z(n13750) );
  IV U13449 ( .A(n13746), .Z(n13748) );
  XOR U13450 ( .A(n13752), .B(n13753), .Z(n13746) );
  AND U13451 ( .A(n659), .B(n13745), .Z(n13753) );
  XNOR U13452 ( .A(n13743), .B(n13752), .Z(n13745) );
  XNOR U13453 ( .A(n13754), .B(n13755), .Z(n13743) );
  AND U13454 ( .A(n663), .B(n13756), .Z(n13755) );
  XOR U13455 ( .A(p_input[920]), .B(n13754), .Z(n13756) );
  XNOR U13456 ( .A(n13757), .B(n13758), .Z(n13754) );
  AND U13457 ( .A(n667), .B(n13759), .Z(n13758) );
  XOR U13458 ( .A(n13760), .B(n13761), .Z(n13752) );
  AND U13459 ( .A(n671), .B(n13751), .Z(n13761) );
  XNOR U13460 ( .A(n13762), .B(n13749), .Z(n13751) );
  XOR U13461 ( .A(n13763), .B(n13764), .Z(n13749) );
  AND U13462 ( .A(n694), .B(n13765), .Z(n13764) );
  IV U13463 ( .A(n13760), .Z(n13762) );
  XOR U13464 ( .A(n13766), .B(n13767), .Z(n13760) );
  AND U13465 ( .A(n678), .B(n13759), .Z(n13767) );
  XNOR U13466 ( .A(n13757), .B(n13766), .Z(n13759) );
  XNOR U13467 ( .A(n13768), .B(n13769), .Z(n13757) );
  AND U13468 ( .A(n682), .B(n13770), .Z(n13769) );
  XOR U13469 ( .A(p_input[952]), .B(n13768), .Z(n13770) );
  XNOR U13470 ( .A(n13771), .B(n13772), .Z(n13768) );
  AND U13471 ( .A(n686), .B(n13773), .Z(n13772) );
  XOR U13472 ( .A(n13774), .B(n13775), .Z(n13766) );
  AND U13473 ( .A(n690), .B(n13765), .Z(n13775) );
  XNOR U13474 ( .A(n13776), .B(n13763), .Z(n13765) );
  XOR U13475 ( .A(n13777), .B(n13778), .Z(n13763) );
  AND U13476 ( .A(n713), .B(n13779), .Z(n13778) );
  IV U13477 ( .A(n13774), .Z(n13776) );
  XOR U13478 ( .A(n13780), .B(n13781), .Z(n13774) );
  AND U13479 ( .A(n697), .B(n13773), .Z(n13781) );
  XNOR U13480 ( .A(n13771), .B(n13780), .Z(n13773) );
  XNOR U13481 ( .A(n13782), .B(n13783), .Z(n13771) );
  AND U13482 ( .A(n701), .B(n13784), .Z(n13783) );
  XOR U13483 ( .A(p_input[984]), .B(n13782), .Z(n13784) );
  XNOR U13484 ( .A(n13785), .B(n13786), .Z(n13782) );
  AND U13485 ( .A(n705), .B(n13787), .Z(n13786) );
  XOR U13486 ( .A(n13788), .B(n13789), .Z(n13780) );
  AND U13487 ( .A(n709), .B(n13779), .Z(n13789) );
  XNOR U13488 ( .A(n13790), .B(n13777), .Z(n13779) );
  XOR U13489 ( .A(n13791), .B(n13792), .Z(n13777) );
  AND U13490 ( .A(n732), .B(n13793), .Z(n13792) );
  IV U13491 ( .A(n13788), .Z(n13790) );
  XOR U13492 ( .A(n13794), .B(n13795), .Z(n13788) );
  AND U13493 ( .A(n716), .B(n13787), .Z(n13795) );
  XNOR U13494 ( .A(n13785), .B(n13794), .Z(n13787) );
  XNOR U13495 ( .A(n13796), .B(n13797), .Z(n13785) );
  AND U13496 ( .A(n720), .B(n13798), .Z(n13797) );
  XOR U13497 ( .A(p_input[1016]), .B(n13796), .Z(n13798) );
  XNOR U13498 ( .A(n13799), .B(n13800), .Z(n13796) );
  AND U13499 ( .A(n724), .B(n13801), .Z(n13800) );
  XOR U13500 ( .A(n13802), .B(n13803), .Z(n13794) );
  AND U13501 ( .A(n728), .B(n13793), .Z(n13803) );
  XNOR U13502 ( .A(n13804), .B(n13791), .Z(n13793) );
  XOR U13503 ( .A(n13805), .B(n13806), .Z(n13791) );
  AND U13504 ( .A(n751), .B(n13807), .Z(n13806) );
  IV U13505 ( .A(n13802), .Z(n13804) );
  XOR U13506 ( .A(n13808), .B(n13809), .Z(n13802) );
  AND U13507 ( .A(n735), .B(n13801), .Z(n13809) );
  XNOR U13508 ( .A(n13799), .B(n13808), .Z(n13801) );
  XNOR U13509 ( .A(n13810), .B(n13811), .Z(n13799) );
  AND U13510 ( .A(n739), .B(n13812), .Z(n13811) );
  XOR U13511 ( .A(p_input[1048]), .B(n13810), .Z(n13812) );
  XNOR U13512 ( .A(n13813), .B(n13814), .Z(n13810) );
  AND U13513 ( .A(n743), .B(n13815), .Z(n13814) );
  XOR U13514 ( .A(n13816), .B(n13817), .Z(n13808) );
  AND U13515 ( .A(n747), .B(n13807), .Z(n13817) );
  XNOR U13516 ( .A(n13818), .B(n13805), .Z(n13807) );
  XOR U13517 ( .A(n13819), .B(n13820), .Z(n13805) );
  AND U13518 ( .A(n770), .B(n13821), .Z(n13820) );
  IV U13519 ( .A(n13816), .Z(n13818) );
  XOR U13520 ( .A(n13822), .B(n13823), .Z(n13816) );
  AND U13521 ( .A(n754), .B(n13815), .Z(n13823) );
  XNOR U13522 ( .A(n13813), .B(n13822), .Z(n13815) );
  XNOR U13523 ( .A(n13824), .B(n13825), .Z(n13813) );
  AND U13524 ( .A(n758), .B(n13826), .Z(n13825) );
  XOR U13525 ( .A(p_input[1080]), .B(n13824), .Z(n13826) );
  XNOR U13526 ( .A(n13827), .B(n13828), .Z(n13824) );
  AND U13527 ( .A(n762), .B(n13829), .Z(n13828) );
  XOR U13528 ( .A(n13830), .B(n13831), .Z(n13822) );
  AND U13529 ( .A(n766), .B(n13821), .Z(n13831) );
  XNOR U13530 ( .A(n13832), .B(n13819), .Z(n13821) );
  XOR U13531 ( .A(n13833), .B(n13834), .Z(n13819) );
  AND U13532 ( .A(n789), .B(n13835), .Z(n13834) );
  IV U13533 ( .A(n13830), .Z(n13832) );
  XOR U13534 ( .A(n13836), .B(n13837), .Z(n13830) );
  AND U13535 ( .A(n773), .B(n13829), .Z(n13837) );
  XNOR U13536 ( .A(n13827), .B(n13836), .Z(n13829) );
  XNOR U13537 ( .A(n13838), .B(n13839), .Z(n13827) );
  AND U13538 ( .A(n777), .B(n13840), .Z(n13839) );
  XOR U13539 ( .A(p_input[1112]), .B(n13838), .Z(n13840) );
  XNOR U13540 ( .A(n13841), .B(n13842), .Z(n13838) );
  AND U13541 ( .A(n781), .B(n13843), .Z(n13842) );
  XOR U13542 ( .A(n13844), .B(n13845), .Z(n13836) );
  AND U13543 ( .A(n785), .B(n13835), .Z(n13845) );
  XNOR U13544 ( .A(n13846), .B(n13833), .Z(n13835) );
  XOR U13545 ( .A(n13847), .B(n13848), .Z(n13833) );
  AND U13546 ( .A(n808), .B(n13849), .Z(n13848) );
  IV U13547 ( .A(n13844), .Z(n13846) );
  XOR U13548 ( .A(n13850), .B(n13851), .Z(n13844) );
  AND U13549 ( .A(n792), .B(n13843), .Z(n13851) );
  XNOR U13550 ( .A(n13841), .B(n13850), .Z(n13843) );
  XNOR U13551 ( .A(n13852), .B(n13853), .Z(n13841) );
  AND U13552 ( .A(n796), .B(n13854), .Z(n13853) );
  XOR U13553 ( .A(p_input[1144]), .B(n13852), .Z(n13854) );
  XNOR U13554 ( .A(n13855), .B(n13856), .Z(n13852) );
  AND U13555 ( .A(n800), .B(n13857), .Z(n13856) );
  XOR U13556 ( .A(n13858), .B(n13859), .Z(n13850) );
  AND U13557 ( .A(n804), .B(n13849), .Z(n13859) );
  XNOR U13558 ( .A(n13860), .B(n13847), .Z(n13849) );
  XOR U13559 ( .A(n13861), .B(n13862), .Z(n13847) );
  AND U13560 ( .A(n827), .B(n13863), .Z(n13862) );
  IV U13561 ( .A(n13858), .Z(n13860) );
  XOR U13562 ( .A(n13864), .B(n13865), .Z(n13858) );
  AND U13563 ( .A(n811), .B(n13857), .Z(n13865) );
  XNOR U13564 ( .A(n13855), .B(n13864), .Z(n13857) );
  XNOR U13565 ( .A(n13866), .B(n13867), .Z(n13855) );
  AND U13566 ( .A(n815), .B(n13868), .Z(n13867) );
  XOR U13567 ( .A(p_input[1176]), .B(n13866), .Z(n13868) );
  XNOR U13568 ( .A(n13869), .B(n13870), .Z(n13866) );
  AND U13569 ( .A(n819), .B(n13871), .Z(n13870) );
  XOR U13570 ( .A(n13872), .B(n13873), .Z(n13864) );
  AND U13571 ( .A(n823), .B(n13863), .Z(n13873) );
  XNOR U13572 ( .A(n13874), .B(n13861), .Z(n13863) );
  XOR U13573 ( .A(n13875), .B(n13876), .Z(n13861) );
  AND U13574 ( .A(n846), .B(n13877), .Z(n13876) );
  IV U13575 ( .A(n13872), .Z(n13874) );
  XOR U13576 ( .A(n13878), .B(n13879), .Z(n13872) );
  AND U13577 ( .A(n830), .B(n13871), .Z(n13879) );
  XNOR U13578 ( .A(n13869), .B(n13878), .Z(n13871) );
  XNOR U13579 ( .A(n13880), .B(n13881), .Z(n13869) );
  AND U13580 ( .A(n834), .B(n13882), .Z(n13881) );
  XOR U13581 ( .A(p_input[1208]), .B(n13880), .Z(n13882) );
  XNOR U13582 ( .A(n13883), .B(n13884), .Z(n13880) );
  AND U13583 ( .A(n838), .B(n13885), .Z(n13884) );
  XOR U13584 ( .A(n13886), .B(n13887), .Z(n13878) );
  AND U13585 ( .A(n842), .B(n13877), .Z(n13887) );
  XNOR U13586 ( .A(n13888), .B(n13875), .Z(n13877) );
  XOR U13587 ( .A(n13889), .B(n13890), .Z(n13875) );
  AND U13588 ( .A(n865), .B(n13891), .Z(n13890) );
  IV U13589 ( .A(n13886), .Z(n13888) );
  XOR U13590 ( .A(n13892), .B(n13893), .Z(n13886) );
  AND U13591 ( .A(n849), .B(n13885), .Z(n13893) );
  XNOR U13592 ( .A(n13883), .B(n13892), .Z(n13885) );
  XNOR U13593 ( .A(n13894), .B(n13895), .Z(n13883) );
  AND U13594 ( .A(n853), .B(n13896), .Z(n13895) );
  XOR U13595 ( .A(p_input[1240]), .B(n13894), .Z(n13896) );
  XNOR U13596 ( .A(n13897), .B(n13898), .Z(n13894) );
  AND U13597 ( .A(n857), .B(n13899), .Z(n13898) );
  XOR U13598 ( .A(n13900), .B(n13901), .Z(n13892) );
  AND U13599 ( .A(n861), .B(n13891), .Z(n13901) );
  XNOR U13600 ( .A(n13902), .B(n13889), .Z(n13891) );
  XOR U13601 ( .A(n13903), .B(n13904), .Z(n13889) );
  AND U13602 ( .A(n884), .B(n13905), .Z(n13904) );
  IV U13603 ( .A(n13900), .Z(n13902) );
  XOR U13604 ( .A(n13906), .B(n13907), .Z(n13900) );
  AND U13605 ( .A(n868), .B(n13899), .Z(n13907) );
  XNOR U13606 ( .A(n13897), .B(n13906), .Z(n13899) );
  XNOR U13607 ( .A(n13908), .B(n13909), .Z(n13897) );
  AND U13608 ( .A(n872), .B(n13910), .Z(n13909) );
  XOR U13609 ( .A(p_input[1272]), .B(n13908), .Z(n13910) );
  XNOR U13610 ( .A(n13911), .B(n13912), .Z(n13908) );
  AND U13611 ( .A(n876), .B(n13913), .Z(n13912) );
  XOR U13612 ( .A(n13914), .B(n13915), .Z(n13906) );
  AND U13613 ( .A(n880), .B(n13905), .Z(n13915) );
  XNOR U13614 ( .A(n13916), .B(n13903), .Z(n13905) );
  XOR U13615 ( .A(n13917), .B(n13918), .Z(n13903) );
  AND U13616 ( .A(n903), .B(n13919), .Z(n13918) );
  IV U13617 ( .A(n13914), .Z(n13916) );
  XOR U13618 ( .A(n13920), .B(n13921), .Z(n13914) );
  AND U13619 ( .A(n887), .B(n13913), .Z(n13921) );
  XNOR U13620 ( .A(n13911), .B(n13920), .Z(n13913) );
  XNOR U13621 ( .A(n13922), .B(n13923), .Z(n13911) );
  AND U13622 ( .A(n891), .B(n13924), .Z(n13923) );
  XOR U13623 ( .A(p_input[1304]), .B(n13922), .Z(n13924) );
  XNOR U13624 ( .A(n13925), .B(n13926), .Z(n13922) );
  AND U13625 ( .A(n895), .B(n13927), .Z(n13926) );
  XOR U13626 ( .A(n13928), .B(n13929), .Z(n13920) );
  AND U13627 ( .A(n899), .B(n13919), .Z(n13929) );
  XNOR U13628 ( .A(n13930), .B(n13917), .Z(n13919) );
  XOR U13629 ( .A(n13931), .B(n13932), .Z(n13917) );
  AND U13630 ( .A(n922), .B(n13933), .Z(n13932) );
  IV U13631 ( .A(n13928), .Z(n13930) );
  XOR U13632 ( .A(n13934), .B(n13935), .Z(n13928) );
  AND U13633 ( .A(n906), .B(n13927), .Z(n13935) );
  XNOR U13634 ( .A(n13925), .B(n13934), .Z(n13927) );
  XNOR U13635 ( .A(n13936), .B(n13937), .Z(n13925) );
  AND U13636 ( .A(n910), .B(n13938), .Z(n13937) );
  XOR U13637 ( .A(p_input[1336]), .B(n13936), .Z(n13938) );
  XNOR U13638 ( .A(n13939), .B(n13940), .Z(n13936) );
  AND U13639 ( .A(n914), .B(n13941), .Z(n13940) );
  XOR U13640 ( .A(n13942), .B(n13943), .Z(n13934) );
  AND U13641 ( .A(n918), .B(n13933), .Z(n13943) );
  XNOR U13642 ( .A(n13944), .B(n13931), .Z(n13933) );
  XOR U13643 ( .A(n13945), .B(n13946), .Z(n13931) );
  AND U13644 ( .A(n941), .B(n13947), .Z(n13946) );
  IV U13645 ( .A(n13942), .Z(n13944) );
  XOR U13646 ( .A(n13948), .B(n13949), .Z(n13942) );
  AND U13647 ( .A(n925), .B(n13941), .Z(n13949) );
  XNOR U13648 ( .A(n13939), .B(n13948), .Z(n13941) );
  XNOR U13649 ( .A(n13950), .B(n13951), .Z(n13939) );
  AND U13650 ( .A(n929), .B(n13952), .Z(n13951) );
  XOR U13651 ( .A(p_input[1368]), .B(n13950), .Z(n13952) );
  XNOR U13652 ( .A(n13953), .B(n13954), .Z(n13950) );
  AND U13653 ( .A(n933), .B(n13955), .Z(n13954) );
  XOR U13654 ( .A(n13956), .B(n13957), .Z(n13948) );
  AND U13655 ( .A(n937), .B(n13947), .Z(n13957) );
  XNOR U13656 ( .A(n13958), .B(n13945), .Z(n13947) );
  XOR U13657 ( .A(n13959), .B(n13960), .Z(n13945) );
  AND U13658 ( .A(n960), .B(n13961), .Z(n13960) );
  IV U13659 ( .A(n13956), .Z(n13958) );
  XOR U13660 ( .A(n13962), .B(n13963), .Z(n13956) );
  AND U13661 ( .A(n944), .B(n13955), .Z(n13963) );
  XNOR U13662 ( .A(n13953), .B(n13962), .Z(n13955) );
  XNOR U13663 ( .A(n13964), .B(n13965), .Z(n13953) );
  AND U13664 ( .A(n948), .B(n13966), .Z(n13965) );
  XOR U13665 ( .A(p_input[1400]), .B(n13964), .Z(n13966) );
  XNOR U13666 ( .A(n13967), .B(n13968), .Z(n13964) );
  AND U13667 ( .A(n952), .B(n13969), .Z(n13968) );
  XOR U13668 ( .A(n13970), .B(n13971), .Z(n13962) );
  AND U13669 ( .A(n956), .B(n13961), .Z(n13971) );
  XNOR U13670 ( .A(n13972), .B(n13959), .Z(n13961) );
  XOR U13671 ( .A(n13973), .B(n13974), .Z(n13959) );
  AND U13672 ( .A(n979), .B(n13975), .Z(n13974) );
  IV U13673 ( .A(n13970), .Z(n13972) );
  XOR U13674 ( .A(n13976), .B(n13977), .Z(n13970) );
  AND U13675 ( .A(n963), .B(n13969), .Z(n13977) );
  XNOR U13676 ( .A(n13967), .B(n13976), .Z(n13969) );
  XNOR U13677 ( .A(n13978), .B(n13979), .Z(n13967) );
  AND U13678 ( .A(n967), .B(n13980), .Z(n13979) );
  XOR U13679 ( .A(p_input[1432]), .B(n13978), .Z(n13980) );
  XNOR U13680 ( .A(n13981), .B(n13982), .Z(n13978) );
  AND U13681 ( .A(n971), .B(n13983), .Z(n13982) );
  XOR U13682 ( .A(n13984), .B(n13985), .Z(n13976) );
  AND U13683 ( .A(n975), .B(n13975), .Z(n13985) );
  XNOR U13684 ( .A(n13986), .B(n13973), .Z(n13975) );
  XOR U13685 ( .A(n13987), .B(n13988), .Z(n13973) );
  AND U13686 ( .A(n998), .B(n13989), .Z(n13988) );
  IV U13687 ( .A(n13984), .Z(n13986) );
  XOR U13688 ( .A(n13990), .B(n13991), .Z(n13984) );
  AND U13689 ( .A(n982), .B(n13983), .Z(n13991) );
  XNOR U13690 ( .A(n13981), .B(n13990), .Z(n13983) );
  XNOR U13691 ( .A(n13992), .B(n13993), .Z(n13981) );
  AND U13692 ( .A(n986), .B(n13994), .Z(n13993) );
  XOR U13693 ( .A(p_input[1464]), .B(n13992), .Z(n13994) );
  XNOR U13694 ( .A(n13995), .B(n13996), .Z(n13992) );
  AND U13695 ( .A(n990), .B(n13997), .Z(n13996) );
  XOR U13696 ( .A(n13998), .B(n13999), .Z(n13990) );
  AND U13697 ( .A(n994), .B(n13989), .Z(n13999) );
  XNOR U13698 ( .A(n14000), .B(n13987), .Z(n13989) );
  XOR U13699 ( .A(n14001), .B(n14002), .Z(n13987) );
  AND U13700 ( .A(n1017), .B(n14003), .Z(n14002) );
  IV U13701 ( .A(n13998), .Z(n14000) );
  XOR U13702 ( .A(n14004), .B(n14005), .Z(n13998) );
  AND U13703 ( .A(n1001), .B(n13997), .Z(n14005) );
  XNOR U13704 ( .A(n13995), .B(n14004), .Z(n13997) );
  XNOR U13705 ( .A(n14006), .B(n14007), .Z(n13995) );
  AND U13706 ( .A(n1005), .B(n14008), .Z(n14007) );
  XOR U13707 ( .A(p_input[1496]), .B(n14006), .Z(n14008) );
  XNOR U13708 ( .A(n14009), .B(n14010), .Z(n14006) );
  AND U13709 ( .A(n1009), .B(n14011), .Z(n14010) );
  XOR U13710 ( .A(n14012), .B(n14013), .Z(n14004) );
  AND U13711 ( .A(n1013), .B(n14003), .Z(n14013) );
  XNOR U13712 ( .A(n14014), .B(n14001), .Z(n14003) );
  XOR U13713 ( .A(n14015), .B(n14016), .Z(n14001) );
  AND U13714 ( .A(n1036), .B(n14017), .Z(n14016) );
  IV U13715 ( .A(n14012), .Z(n14014) );
  XOR U13716 ( .A(n14018), .B(n14019), .Z(n14012) );
  AND U13717 ( .A(n1020), .B(n14011), .Z(n14019) );
  XNOR U13718 ( .A(n14009), .B(n14018), .Z(n14011) );
  XNOR U13719 ( .A(n14020), .B(n14021), .Z(n14009) );
  AND U13720 ( .A(n1024), .B(n14022), .Z(n14021) );
  XOR U13721 ( .A(p_input[1528]), .B(n14020), .Z(n14022) );
  XNOR U13722 ( .A(n14023), .B(n14024), .Z(n14020) );
  AND U13723 ( .A(n1028), .B(n14025), .Z(n14024) );
  XOR U13724 ( .A(n14026), .B(n14027), .Z(n14018) );
  AND U13725 ( .A(n1032), .B(n14017), .Z(n14027) );
  XNOR U13726 ( .A(n14028), .B(n14015), .Z(n14017) );
  XOR U13727 ( .A(n14029), .B(n14030), .Z(n14015) );
  AND U13728 ( .A(n1055), .B(n14031), .Z(n14030) );
  IV U13729 ( .A(n14026), .Z(n14028) );
  XOR U13730 ( .A(n14032), .B(n14033), .Z(n14026) );
  AND U13731 ( .A(n1039), .B(n14025), .Z(n14033) );
  XNOR U13732 ( .A(n14023), .B(n14032), .Z(n14025) );
  XNOR U13733 ( .A(n14034), .B(n14035), .Z(n14023) );
  AND U13734 ( .A(n1043), .B(n14036), .Z(n14035) );
  XOR U13735 ( .A(p_input[1560]), .B(n14034), .Z(n14036) );
  XNOR U13736 ( .A(n14037), .B(n14038), .Z(n14034) );
  AND U13737 ( .A(n1047), .B(n14039), .Z(n14038) );
  XOR U13738 ( .A(n14040), .B(n14041), .Z(n14032) );
  AND U13739 ( .A(n1051), .B(n14031), .Z(n14041) );
  XNOR U13740 ( .A(n14042), .B(n14029), .Z(n14031) );
  XOR U13741 ( .A(n14043), .B(n14044), .Z(n14029) );
  AND U13742 ( .A(n1074), .B(n14045), .Z(n14044) );
  IV U13743 ( .A(n14040), .Z(n14042) );
  XOR U13744 ( .A(n14046), .B(n14047), .Z(n14040) );
  AND U13745 ( .A(n1058), .B(n14039), .Z(n14047) );
  XNOR U13746 ( .A(n14037), .B(n14046), .Z(n14039) );
  XNOR U13747 ( .A(n14048), .B(n14049), .Z(n14037) );
  AND U13748 ( .A(n1062), .B(n14050), .Z(n14049) );
  XOR U13749 ( .A(p_input[1592]), .B(n14048), .Z(n14050) );
  XNOR U13750 ( .A(n14051), .B(n14052), .Z(n14048) );
  AND U13751 ( .A(n1066), .B(n14053), .Z(n14052) );
  XOR U13752 ( .A(n14054), .B(n14055), .Z(n14046) );
  AND U13753 ( .A(n1070), .B(n14045), .Z(n14055) );
  XNOR U13754 ( .A(n14056), .B(n14043), .Z(n14045) );
  XOR U13755 ( .A(n14057), .B(n14058), .Z(n14043) );
  AND U13756 ( .A(n1093), .B(n14059), .Z(n14058) );
  IV U13757 ( .A(n14054), .Z(n14056) );
  XOR U13758 ( .A(n14060), .B(n14061), .Z(n14054) );
  AND U13759 ( .A(n1077), .B(n14053), .Z(n14061) );
  XNOR U13760 ( .A(n14051), .B(n14060), .Z(n14053) );
  XNOR U13761 ( .A(n14062), .B(n14063), .Z(n14051) );
  AND U13762 ( .A(n1081), .B(n14064), .Z(n14063) );
  XOR U13763 ( .A(p_input[1624]), .B(n14062), .Z(n14064) );
  XNOR U13764 ( .A(n14065), .B(n14066), .Z(n14062) );
  AND U13765 ( .A(n1085), .B(n14067), .Z(n14066) );
  XOR U13766 ( .A(n14068), .B(n14069), .Z(n14060) );
  AND U13767 ( .A(n1089), .B(n14059), .Z(n14069) );
  XNOR U13768 ( .A(n14070), .B(n14057), .Z(n14059) );
  XOR U13769 ( .A(n14071), .B(n14072), .Z(n14057) );
  AND U13770 ( .A(n1112), .B(n14073), .Z(n14072) );
  IV U13771 ( .A(n14068), .Z(n14070) );
  XOR U13772 ( .A(n14074), .B(n14075), .Z(n14068) );
  AND U13773 ( .A(n1096), .B(n14067), .Z(n14075) );
  XNOR U13774 ( .A(n14065), .B(n14074), .Z(n14067) );
  XNOR U13775 ( .A(n14076), .B(n14077), .Z(n14065) );
  AND U13776 ( .A(n1100), .B(n14078), .Z(n14077) );
  XOR U13777 ( .A(p_input[1656]), .B(n14076), .Z(n14078) );
  XNOR U13778 ( .A(n14079), .B(n14080), .Z(n14076) );
  AND U13779 ( .A(n1104), .B(n14081), .Z(n14080) );
  XOR U13780 ( .A(n14082), .B(n14083), .Z(n14074) );
  AND U13781 ( .A(n1108), .B(n14073), .Z(n14083) );
  XNOR U13782 ( .A(n14084), .B(n14071), .Z(n14073) );
  XOR U13783 ( .A(n14085), .B(n14086), .Z(n14071) );
  AND U13784 ( .A(n1131), .B(n14087), .Z(n14086) );
  IV U13785 ( .A(n14082), .Z(n14084) );
  XOR U13786 ( .A(n14088), .B(n14089), .Z(n14082) );
  AND U13787 ( .A(n1115), .B(n14081), .Z(n14089) );
  XNOR U13788 ( .A(n14079), .B(n14088), .Z(n14081) );
  XNOR U13789 ( .A(n14090), .B(n14091), .Z(n14079) );
  AND U13790 ( .A(n1119), .B(n14092), .Z(n14091) );
  XOR U13791 ( .A(p_input[1688]), .B(n14090), .Z(n14092) );
  XNOR U13792 ( .A(n14093), .B(n14094), .Z(n14090) );
  AND U13793 ( .A(n1123), .B(n14095), .Z(n14094) );
  XOR U13794 ( .A(n14096), .B(n14097), .Z(n14088) );
  AND U13795 ( .A(n1127), .B(n14087), .Z(n14097) );
  XNOR U13796 ( .A(n14098), .B(n14085), .Z(n14087) );
  XOR U13797 ( .A(n14099), .B(n14100), .Z(n14085) );
  AND U13798 ( .A(n1150), .B(n14101), .Z(n14100) );
  IV U13799 ( .A(n14096), .Z(n14098) );
  XOR U13800 ( .A(n14102), .B(n14103), .Z(n14096) );
  AND U13801 ( .A(n1134), .B(n14095), .Z(n14103) );
  XNOR U13802 ( .A(n14093), .B(n14102), .Z(n14095) );
  XNOR U13803 ( .A(n14104), .B(n14105), .Z(n14093) );
  AND U13804 ( .A(n1138), .B(n14106), .Z(n14105) );
  XOR U13805 ( .A(p_input[1720]), .B(n14104), .Z(n14106) );
  XNOR U13806 ( .A(n14107), .B(n14108), .Z(n14104) );
  AND U13807 ( .A(n1142), .B(n14109), .Z(n14108) );
  XOR U13808 ( .A(n14110), .B(n14111), .Z(n14102) );
  AND U13809 ( .A(n1146), .B(n14101), .Z(n14111) );
  XNOR U13810 ( .A(n14112), .B(n14099), .Z(n14101) );
  XOR U13811 ( .A(n14113), .B(n14114), .Z(n14099) );
  AND U13812 ( .A(n1169), .B(n14115), .Z(n14114) );
  IV U13813 ( .A(n14110), .Z(n14112) );
  XOR U13814 ( .A(n14116), .B(n14117), .Z(n14110) );
  AND U13815 ( .A(n1153), .B(n14109), .Z(n14117) );
  XNOR U13816 ( .A(n14107), .B(n14116), .Z(n14109) );
  XNOR U13817 ( .A(n14118), .B(n14119), .Z(n14107) );
  AND U13818 ( .A(n1157), .B(n14120), .Z(n14119) );
  XOR U13819 ( .A(p_input[1752]), .B(n14118), .Z(n14120) );
  XNOR U13820 ( .A(n14121), .B(n14122), .Z(n14118) );
  AND U13821 ( .A(n1161), .B(n14123), .Z(n14122) );
  XOR U13822 ( .A(n14124), .B(n14125), .Z(n14116) );
  AND U13823 ( .A(n1165), .B(n14115), .Z(n14125) );
  XNOR U13824 ( .A(n14126), .B(n14113), .Z(n14115) );
  XOR U13825 ( .A(n14127), .B(n14128), .Z(n14113) );
  AND U13826 ( .A(n1188), .B(n14129), .Z(n14128) );
  IV U13827 ( .A(n14124), .Z(n14126) );
  XOR U13828 ( .A(n14130), .B(n14131), .Z(n14124) );
  AND U13829 ( .A(n1172), .B(n14123), .Z(n14131) );
  XNOR U13830 ( .A(n14121), .B(n14130), .Z(n14123) );
  XNOR U13831 ( .A(n14132), .B(n14133), .Z(n14121) );
  AND U13832 ( .A(n1176), .B(n14134), .Z(n14133) );
  XOR U13833 ( .A(p_input[1784]), .B(n14132), .Z(n14134) );
  XNOR U13834 ( .A(n14135), .B(n14136), .Z(n14132) );
  AND U13835 ( .A(n1180), .B(n14137), .Z(n14136) );
  XOR U13836 ( .A(n14138), .B(n14139), .Z(n14130) );
  AND U13837 ( .A(n1184), .B(n14129), .Z(n14139) );
  XNOR U13838 ( .A(n14140), .B(n14127), .Z(n14129) );
  XOR U13839 ( .A(n14141), .B(n14142), .Z(n14127) );
  AND U13840 ( .A(n1207), .B(n14143), .Z(n14142) );
  IV U13841 ( .A(n14138), .Z(n14140) );
  XOR U13842 ( .A(n14144), .B(n14145), .Z(n14138) );
  AND U13843 ( .A(n1191), .B(n14137), .Z(n14145) );
  XNOR U13844 ( .A(n14135), .B(n14144), .Z(n14137) );
  XNOR U13845 ( .A(n14146), .B(n14147), .Z(n14135) );
  AND U13846 ( .A(n1195), .B(n14148), .Z(n14147) );
  XOR U13847 ( .A(p_input[1816]), .B(n14146), .Z(n14148) );
  XNOR U13848 ( .A(n14149), .B(n14150), .Z(n14146) );
  AND U13849 ( .A(n1199), .B(n14151), .Z(n14150) );
  XOR U13850 ( .A(n14152), .B(n14153), .Z(n14144) );
  AND U13851 ( .A(n1203), .B(n14143), .Z(n14153) );
  XNOR U13852 ( .A(n14154), .B(n14141), .Z(n14143) );
  XOR U13853 ( .A(n14155), .B(n14156), .Z(n14141) );
  AND U13854 ( .A(n1226), .B(n14157), .Z(n14156) );
  IV U13855 ( .A(n14152), .Z(n14154) );
  XOR U13856 ( .A(n14158), .B(n14159), .Z(n14152) );
  AND U13857 ( .A(n1210), .B(n14151), .Z(n14159) );
  XNOR U13858 ( .A(n14149), .B(n14158), .Z(n14151) );
  XNOR U13859 ( .A(n14160), .B(n14161), .Z(n14149) );
  AND U13860 ( .A(n1214), .B(n14162), .Z(n14161) );
  XOR U13861 ( .A(p_input[1848]), .B(n14160), .Z(n14162) );
  XNOR U13862 ( .A(n14163), .B(n14164), .Z(n14160) );
  AND U13863 ( .A(n1218), .B(n14165), .Z(n14164) );
  XOR U13864 ( .A(n14166), .B(n14167), .Z(n14158) );
  AND U13865 ( .A(n1222), .B(n14157), .Z(n14167) );
  XNOR U13866 ( .A(n14168), .B(n14155), .Z(n14157) );
  XOR U13867 ( .A(n14169), .B(n14170), .Z(n14155) );
  AND U13868 ( .A(n1245), .B(n14171), .Z(n14170) );
  IV U13869 ( .A(n14166), .Z(n14168) );
  XOR U13870 ( .A(n14172), .B(n14173), .Z(n14166) );
  AND U13871 ( .A(n1229), .B(n14165), .Z(n14173) );
  XNOR U13872 ( .A(n14163), .B(n14172), .Z(n14165) );
  XNOR U13873 ( .A(n14174), .B(n14175), .Z(n14163) );
  AND U13874 ( .A(n1233), .B(n14176), .Z(n14175) );
  XOR U13875 ( .A(p_input[1880]), .B(n14174), .Z(n14176) );
  XNOR U13876 ( .A(n14177), .B(n14178), .Z(n14174) );
  AND U13877 ( .A(n1237), .B(n14179), .Z(n14178) );
  XOR U13878 ( .A(n14180), .B(n14181), .Z(n14172) );
  AND U13879 ( .A(n1241), .B(n14171), .Z(n14181) );
  XNOR U13880 ( .A(n14182), .B(n14169), .Z(n14171) );
  XOR U13881 ( .A(n14183), .B(n14184), .Z(n14169) );
  AND U13882 ( .A(n1264), .B(n14185), .Z(n14184) );
  IV U13883 ( .A(n14180), .Z(n14182) );
  XOR U13884 ( .A(n14186), .B(n14187), .Z(n14180) );
  AND U13885 ( .A(n1248), .B(n14179), .Z(n14187) );
  XNOR U13886 ( .A(n14177), .B(n14186), .Z(n14179) );
  XNOR U13887 ( .A(n14188), .B(n14189), .Z(n14177) );
  AND U13888 ( .A(n1252), .B(n14190), .Z(n14189) );
  XOR U13889 ( .A(p_input[1912]), .B(n14188), .Z(n14190) );
  XNOR U13890 ( .A(n14191), .B(n14192), .Z(n14188) );
  AND U13891 ( .A(n1256), .B(n14193), .Z(n14192) );
  XOR U13892 ( .A(n14194), .B(n14195), .Z(n14186) );
  AND U13893 ( .A(n1260), .B(n14185), .Z(n14195) );
  XNOR U13894 ( .A(n14196), .B(n14183), .Z(n14185) );
  XOR U13895 ( .A(n14197), .B(n14198), .Z(n14183) );
  AND U13896 ( .A(n1282), .B(n14199), .Z(n14198) );
  IV U13897 ( .A(n14194), .Z(n14196) );
  XOR U13898 ( .A(n14200), .B(n14201), .Z(n14194) );
  AND U13899 ( .A(n1267), .B(n14193), .Z(n14201) );
  XNOR U13900 ( .A(n14191), .B(n14200), .Z(n14193) );
  XNOR U13901 ( .A(n14202), .B(n14203), .Z(n14191) );
  AND U13902 ( .A(n1271), .B(n14204), .Z(n14203) );
  XOR U13903 ( .A(p_input[1944]), .B(n14202), .Z(n14204) );
  XOR U13904 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][24] ), .B(n14205), 
        .Z(n14202) );
  AND U13905 ( .A(n1274), .B(n14206), .Z(n14205) );
  XOR U13906 ( .A(n14207), .B(n14208), .Z(n14200) );
  AND U13907 ( .A(n1278), .B(n14199), .Z(n14208) );
  XNOR U13908 ( .A(n14209), .B(n14197), .Z(n14199) );
  XOR U13909 ( .A(\knn_comb_/min_val_out[0][24] ), .B(n14210), .Z(n14197) );
  AND U13910 ( .A(n1290), .B(n14211), .Z(n14210) );
  IV U13911 ( .A(n14207), .Z(n14209) );
  XOR U13912 ( .A(n14212), .B(n14213), .Z(n14207) );
  AND U13913 ( .A(n1285), .B(n14206), .Z(n14213) );
  XOR U13914 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][24] ), .B(n14212), 
        .Z(n14206) );
  XOR U13915 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .B(n14214), 
        .Z(n14212) );
  AND U13916 ( .A(n1287), .B(n14211), .Z(n14214) );
  XOR U13917 ( .A(\knn_comb_/min_val_out[0][24] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .Z(n14211) );
  XOR U13918 ( .A(n91), .B(n14215), .Z(o[23]) );
  AND U13919 ( .A(n122), .B(n14216), .Z(n91) );
  XOR U13920 ( .A(n92), .B(n14215), .Z(n14216) );
  XOR U13921 ( .A(n14217), .B(n14218), .Z(n14215) );
  AND U13922 ( .A(n142), .B(n14219), .Z(n14218) );
  XOR U13923 ( .A(n14220), .B(n21), .Z(n92) );
  AND U13924 ( .A(n125), .B(n14221), .Z(n21) );
  XOR U13925 ( .A(n22), .B(n14220), .Z(n14221) );
  XOR U13926 ( .A(n14222), .B(n14223), .Z(n22) );
  AND U13927 ( .A(n130), .B(n14224), .Z(n14223) );
  XOR U13928 ( .A(p_input[23]), .B(n14222), .Z(n14224) );
  XNOR U13929 ( .A(n14225), .B(n14226), .Z(n14222) );
  AND U13930 ( .A(n134), .B(n14227), .Z(n14226) );
  XOR U13931 ( .A(n14228), .B(n14229), .Z(n14220) );
  AND U13932 ( .A(n138), .B(n14219), .Z(n14229) );
  XNOR U13933 ( .A(n14230), .B(n14217), .Z(n14219) );
  XOR U13934 ( .A(n14231), .B(n14232), .Z(n14217) );
  AND U13935 ( .A(n162), .B(n14233), .Z(n14232) );
  IV U13936 ( .A(n14228), .Z(n14230) );
  XOR U13937 ( .A(n14234), .B(n14235), .Z(n14228) );
  AND U13938 ( .A(n146), .B(n14227), .Z(n14235) );
  XNOR U13939 ( .A(n14225), .B(n14234), .Z(n14227) );
  XNOR U13940 ( .A(n14236), .B(n14237), .Z(n14225) );
  AND U13941 ( .A(n150), .B(n14238), .Z(n14237) );
  XOR U13942 ( .A(p_input[55]), .B(n14236), .Z(n14238) );
  XNOR U13943 ( .A(n14239), .B(n14240), .Z(n14236) );
  AND U13944 ( .A(n154), .B(n14241), .Z(n14240) );
  XOR U13945 ( .A(n14242), .B(n14243), .Z(n14234) );
  AND U13946 ( .A(n158), .B(n14233), .Z(n14243) );
  XNOR U13947 ( .A(n14244), .B(n14231), .Z(n14233) );
  XOR U13948 ( .A(n14245), .B(n14246), .Z(n14231) );
  AND U13949 ( .A(n181), .B(n14247), .Z(n14246) );
  IV U13950 ( .A(n14242), .Z(n14244) );
  XOR U13951 ( .A(n14248), .B(n14249), .Z(n14242) );
  AND U13952 ( .A(n165), .B(n14241), .Z(n14249) );
  XNOR U13953 ( .A(n14239), .B(n14248), .Z(n14241) );
  XNOR U13954 ( .A(n14250), .B(n14251), .Z(n14239) );
  AND U13955 ( .A(n169), .B(n14252), .Z(n14251) );
  XOR U13956 ( .A(p_input[87]), .B(n14250), .Z(n14252) );
  XNOR U13957 ( .A(n14253), .B(n14254), .Z(n14250) );
  AND U13958 ( .A(n173), .B(n14255), .Z(n14254) );
  XOR U13959 ( .A(n14256), .B(n14257), .Z(n14248) );
  AND U13960 ( .A(n177), .B(n14247), .Z(n14257) );
  XNOR U13961 ( .A(n14258), .B(n14245), .Z(n14247) );
  XOR U13962 ( .A(n14259), .B(n14260), .Z(n14245) );
  AND U13963 ( .A(n200), .B(n14261), .Z(n14260) );
  IV U13964 ( .A(n14256), .Z(n14258) );
  XOR U13965 ( .A(n14262), .B(n14263), .Z(n14256) );
  AND U13966 ( .A(n184), .B(n14255), .Z(n14263) );
  XNOR U13967 ( .A(n14253), .B(n14262), .Z(n14255) );
  XNOR U13968 ( .A(n14264), .B(n14265), .Z(n14253) );
  AND U13969 ( .A(n188), .B(n14266), .Z(n14265) );
  XOR U13970 ( .A(p_input[119]), .B(n14264), .Z(n14266) );
  XNOR U13971 ( .A(n14267), .B(n14268), .Z(n14264) );
  AND U13972 ( .A(n192), .B(n14269), .Z(n14268) );
  XOR U13973 ( .A(n14270), .B(n14271), .Z(n14262) );
  AND U13974 ( .A(n196), .B(n14261), .Z(n14271) );
  XNOR U13975 ( .A(n14272), .B(n14259), .Z(n14261) );
  XOR U13976 ( .A(n14273), .B(n14274), .Z(n14259) );
  AND U13977 ( .A(n219), .B(n14275), .Z(n14274) );
  IV U13978 ( .A(n14270), .Z(n14272) );
  XOR U13979 ( .A(n14276), .B(n14277), .Z(n14270) );
  AND U13980 ( .A(n203), .B(n14269), .Z(n14277) );
  XNOR U13981 ( .A(n14267), .B(n14276), .Z(n14269) );
  XNOR U13982 ( .A(n14278), .B(n14279), .Z(n14267) );
  AND U13983 ( .A(n207), .B(n14280), .Z(n14279) );
  XOR U13984 ( .A(p_input[151]), .B(n14278), .Z(n14280) );
  XNOR U13985 ( .A(n14281), .B(n14282), .Z(n14278) );
  AND U13986 ( .A(n211), .B(n14283), .Z(n14282) );
  XOR U13987 ( .A(n14284), .B(n14285), .Z(n14276) );
  AND U13988 ( .A(n215), .B(n14275), .Z(n14285) );
  XNOR U13989 ( .A(n14286), .B(n14273), .Z(n14275) );
  XOR U13990 ( .A(n14287), .B(n14288), .Z(n14273) );
  AND U13991 ( .A(n238), .B(n14289), .Z(n14288) );
  IV U13992 ( .A(n14284), .Z(n14286) );
  XOR U13993 ( .A(n14290), .B(n14291), .Z(n14284) );
  AND U13994 ( .A(n222), .B(n14283), .Z(n14291) );
  XNOR U13995 ( .A(n14281), .B(n14290), .Z(n14283) );
  XNOR U13996 ( .A(n14292), .B(n14293), .Z(n14281) );
  AND U13997 ( .A(n226), .B(n14294), .Z(n14293) );
  XOR U13998 ( .A(p_input[183]), .B(n14292), .Z(n14294) );
  XNOR U13999 ( .A(n14295), .B(n14296), .Z(n14292) );
  AND U14000 ( .A(n230), .B(n14297), .Z(n14296) );
  XOR U14001 ( .A(n14298), .B(n14299), .Z(n14290) );
  AND U14002 ( .A(n234), .B(n14289), .Z(n14299) );
  XNOR U14003 ( .A(n14300), .B(n14287), .Z(n14289) );
  XOR U14004 ( .A(n14301), .B(n14302), .Z(n14287) );
  AND U14005 ( .A(n257), .B(n14303), .Z(n14302) );
  IV U14006 ( .A(n14298), .Z(n14300) );
  XOR U14007 ( .A(n14304), .B(n14305), .Z(n14298) );
  AND U14008 ( .A(n241), .B(n14297), .Z(n14305) );
  XNOR U14009 ( .A(n14295), .B(n14304), .Z(n14297) );
  XNOR U14010 ( .A(n14306), .B(n14307), .Z(n14295) );
  AND U14011 ( .A(n245), .B(n14308), .Z(n14307) );
  XOR U14012 ( .A(p_input[215]), .B(n14306), .Z(n14308) );
  XNOR U14013 ( .A(n14309), .B(n14310), .Z(n14306) );
  AND U14014 ( .A(n249), .B(n14311), .Z(n14310) );
  XOR U14015 ( .A(n14312), .B(n14313), .Z(n14304) );
  AND U14016 ( .A(n253), .B(n14303), .Z(n14313) );
  XNOR U14017 ( .A(n14314), .B(n14301), .Z(n14303) );
  XOR U14018 ( .A(n14315), .B(n14316), .Z(n14301) );
  AND U14019 ( .A(n276), .B(n14317), .Z(n14316) );
  IV U14020 ( .A(n14312), .Z(n14314) );
  XOR U14021 ( .A(n14318), .B(n14319), .Z(n14312) );
  AND U14022 ( .A(n260), .B(n14311), .Z(n14319) );
  XNOR U14023 ( .A(n14309), .B(n14318), .Z(n14311) );
  XNOR U14024 ( .A(n14320), .B(n14321), .Z(n14309) );
  AND U14025 ( .A(n264), .B(n14322), .Z(n14321) );
  XOR U14026 ( .A(p_input[247]), .B(n14320), .Z(n14322) );
  XNOR U14027 ( .A(n14323), .B(n14324), .Z(n14320) );
  AND U14028 ( .A(n268), .B(n14325), .Z(n14324) );
  XOR U14029 ( .A(n14326), .B(n14327), .Z(n14318) );
  AND U14030 ( .A(n272), .B(n14317), .Z(n14327) );
  XNOR U14031 ( .A(n14328), .B(n14315), .Z(n14317) );
  XOR U14032 ( .A(n14329), .B(n14330), .Z(n14315) );
  AND U14033 ( .A(n295), .B(n14331), .Z(n14330) );
  IV U14034 ( .A(n14326), .Z(n14328) );
  XOR U14035 ( .A(n14332), .B(n14333), .Z(n14326) );
  AND U14036 ( .A(n279), .B(n14325), .Z(n14333) );
  XNOR U14037 ( .A(n14323), .B(n14332), .Z(n14325) );
  XNOR U14038 ( .A(n14334), .B(n14335), .Z(n14323) );
  AND U14039 ( .A(n283), .B(n14336), .Z(n14335) );
  XOR U14040 ( .A(p_input[279]), .B(n14334), .Z(n14336) );
  XNOR U14041 ( .A(n14337), .B(n14338), .Z(n14334) );
  AND U14042 ( .A(n287), .B(n14339), .Z(n14338) );
  XOR U14043 ( .A(n14340), .B(n14341), .Z(n14332) );
  AND U14044 ( .A(n291), .B(n14331), .Z(n14341) );
  XNOR U14045 ( .A(n14342), .B(n14329), .Z(n14331) );
  XOR U14046 ( .A(n14343), .B(n14344), .Z(n14329) );
  AND U14047 ( .A(n314), .B(n14345), .Z(n14344) );
  IV U14048 ( .A(n14340), .Z(n14342) );
  XOR U14049 ( .A(n14346), .B(n14347), .Z(n14340) );
  AND U14050 ( .A(n298), .B(n14339), .Z(n14347) );
  XNOR U14051 ( .A(n14337), .B(n14346), .Z(n14339) );
  XNOR U14052 ( .A(n14348), .B(n14349), .Z(n14337) );
  AND U14053 ( .A(n302), .B(n14350), .Z(n14349) );
  XOR U14054 ( .A(p_input[311]), .B(n14348), .Z(n14350) );
  XNOR U14055 ( .A(n14351), .B(n14352), .Z(n14348) );
  AND U14056 ( .A(n306), .B(n14353), .Z(n14352) );
  XOR U14057 ( .A(n14354), .B(n14355), .Z(n14346) );
  AND U14058 ( .A(n310), .B(n14345), .Z(n14355) );
  XNOR U14059 ( .A(n14356), .B(n14343), .Z(n14345) );
  XOR U14060 ( .A(n14357), .B(n14358), .Z(n14343) );
  AND U14061 ( .A(n333), .B(n14359), .Z(n14358) );
  IV U14062 ( .A(n14354), .Z(n14356) );
  XOR U14063 ( .A(n14360), .B(n14361), .Z(n14354) );
  AND U14064 ( .A(n317), .B(n14353), .Z(n14361) );
  XNOR U14065 ( .A(n14351), .B(n14360), .Z(n14353) );
  XNOR U14066 ( .A(n14362), .B(n14363), .Z(n14351) );
  AND U14067 ( .A(n321), .B(n14364), .Z(n14363) );
  XOR U14068 ( .A(p_input[343]), .B(n14362), .Z(n14364) );
  XNOR U14069 ( .A(n14365), .B(n14366), .Z(n14362) );
  AND U14070 ( .A(n325), .B(n14367), .Z(n14366) );
  XOR U14071 ( .A(n14368), .B(n14369), .Z(n14360) );
  AND U14072 ( .A(n329), .B(n14359), .Z(n14369) );
  XNOR U14073 ( .A(n14370), .B(n14357), .Z(n14359) );
  XOR U14074 ( .A(n14371), .B(n14372), .Z(n14357) );
  AND U14075 ( .A(n352), .B(n14373), .Z(n14372) );
  IV U14076 ( .A(n14368), .Z(n14370) );
  XOR U14077 ( .A(n14374), .B(n14375), .Z(n14368) );
  AND U14078 ( .A(n336), .B(n14367), .Z(n14375) );
  XNOR U14079 ( .A(n14365), .B(n14374), .Z(n14367) );
  XNOR U14080 ( .A(n14376), .B(n14377), .Z(n14365) );
  AND U14081 ( .A(n340), .B(n14378), .Z(n14377) );
  XOR U14082 ( .A(p_input[375]), .B(n14376), .Z(n14378) );
  XNOR U14083 ( .A(n14379), .B(n14380), .Z(n14376) );
  AND U14084 ( .A(n344), .B(n14381), .Z(n14380) );
  XOR U14085 ( .A(n14382), .B(n14383), .Z(n14374) );
  AND U14086 ( .A(n348), .B(n14373), .Z(n14383) );
  XNOR U14087 ( .A(n14384), .B(n14371), .Z(n14373) );
  XOR U14088 ( .A(n14385), .B(n14386), .Z(n14371) );
  AND U14089 ( .A(n371), .B(n14387), .Z(n14386) );
  IV U14090 ( .A(n14382), .Z(n14384) );
  XOR U14091 ( .A(n14388), .B(n14389), .Z(n14382) );
  AND U14092 ( .A(n355), .B(n14381), .Z(n14389) );
  XNOR U14093 ( .A(n14379), .B(n14388), .Z(n14381) );
  XNOR U14094 ( .A(n14390), .B(n14391), .Z(n14379) );
  AND U14095 ( .A(n359), .B(n14392), .Z(n14391) );
  XOR U14096 ( .A(p_input[407]), .B(n14390), .Z(n14392) );
  XNOR U14097 ( .A(n14393), .B(n14394), .Z(n14390) );
  AND U14098 ( .A(n363), .B(n14395), .Z(n14394) );
  XOR U14099 ( .A(n14396), .B(n14397), .Z(n14388) );
  AND U14100 ( .A(n367), .B(n14387), .Z(n14397) );
  XNOR U14101 ( .A(n14398), .B(n14385), .Z(n14387) );
  XOR U14102 ( .A(n14399), .B(n14400), .Z(n14385) );
  AND U14103 ( .A(n390), .B(n14401), .Z(n14400) );
  IV U14104 ( .A(n14396), .Z(n14398) );
  XOR U14105 ( .A(n14402), .B(n14403), .Z(n14396) );
  AND U14106 ( .A(n374), .B(n14395), .Z(n14403) );
  XNOR U14107 ( .A(n14393), .B(n14402), .Z(n14395) );
  XNOR U14108 ( .A(n14404), .B(n14405), .Z(n14393) );
  AND U14109 ( .A(n378), .B(n14406), .Z(n14405) );
  XOR U14110 ( .A(p_input[439]), .B(n14404), .Z(n14406) );
  XNOR U14111 ( .A(n14407), .B(n14408), .Z(n14404) );
  AND U14112 ( .A(n382), .B(n14409), .Z(n14408) );
  XOR U14113 ( .A(n14410), .B(n14411), .Z(n14402) );
  AND U14114 ( .A(n386), .B(n14401), .Z(n14411) );
  XNOR U14115 ( .A(n14412), .B(n14399), .Z(n14401) );
  XOR U14116 ( .A(n14413), .B(n14414), .Z(n14399) );
  AND U14117 ( .A(n409), .B(n14415), .Z(n14414) );
  IV U14118 ( .A(n14410), .Z(n14412) );
  XOR U14119 ( .A(n14416), .B(n14417), .Z(n14410) );
  AND U14120 ( .A(n393), .B(n14409), .Z(n14417) );
  XNOR U14121 ( .A(n14407), .B(n14416), .Z(n14409) );
  XNOR U14122 ( .A(n14418), .B(n14419), .Z(n14407) );
  AND U14123 ( .A(n397), .B(n14420), .Z(n14419) );
  XOR U14124 ( .A(p_input[471]), .B(n14418), .Z(n14420) );
  XNOR U14125 ( .A(n14421), .B(n14422), .Z(n14418) );
  AND U14126 ( .A(n401), .B(n14423), .Z(n14422) );
  XOR U14127 ( .A(n14424), .B(n14425), .Z(n14416) );
  AND U14128 ( .A(n405), .B(n14415), .Z(n14425) );
  XNOR U14129 ( .A(n14426), .B(n14413), .Z(n14415) );
  XOR U14130 ( .A(n14427), .B(n14428), .Z(n14413) );
  AND U14131 ( .A(n428), .B(n14429), .Z(n14428) );
  IV U14132 ( .A(n14424), .Z(n14426) );
  XOR U14133 ( .A(n14430), .B(n14431), .Z(n14424) );
  AND U14134 ( .A(n412), .B(n14423), .Z(n14431) );
  XNOR U14135 ( .A(n14421), .B(n14430), .Z(n14423) );
  XNOR U14136 ( .A(n14432), .B(n14433), .Z(n14421) );
  AND U14137 ( .A(n416), .B(n14434), .Z(n14433) );
  XOR U14138 ( .A(p_input[503]), .B(n14432), .Z(n14434) );
  XNOR U14139 ( .A(n14435), .B(n14436), .Z(n14432) );
  AND U14140 ( .A(n420), .B(n14437), .Z(n14436) );
  XOR U14141 ( .A(n14438), .B(n14439), .Z(n14430) );
  AND U14142 ( .A(n424), .B(n14429), .Z(n14439) );
  XNOR U14143 ( .A(n14440), .B(n14427), .Z(n14429) );
  XOR U14144 ( .A(n14441), .B(n14442), .Z(n14427) );
  AND U14145 ( .A(n447), .B(n14443), .Z(n14442) );
  IV U14146 ( .A(n14438), .Z(n14440) );
  XOR U14147 ( .A(n14444), .B(n14445), .Z(n14438) );
  AND U14148 ( .A(n431), .B(n14437), .Z(n14445) );
  XNOR U14149 ( .A(n14435), .B(n14444), .Z(n14437) );
  XNOR U14150 ( .A(n14446), .B(n14447), .Z(n14435) );
  AND U14151 ( .A(n435), .B(n14448), .Z(n14447) );
  XOR U14152 ( .A(p_input[535]), .B(n14446), .Z(n14448) );
  XNOR U14153 ( .A(n14449), .B(n14450), .Z(n14446) );
  AND U14154 ( .A(n439), .B(n14451), .Z(n14450) );
  XOR U14155 ( .A(n14452), .B(n14453), .Z(n14444) );
  AND U14156 ( .A(n443), .B(n14443), .Z(n14453) );
  XNOR U14157 ( .A(n14454), .B(n14441), .Z(n14443) );
  XOR U14158 ( .A(n14455), .B(n14456), .Z(n14441) );
  AND U14159 ( .A(n466), .B(n14457), .Z(n14456) );
  IV U14160 ( .A(n14452), .Z(n14454) );
  XOR U14161 ( .A(n14458), .B(n14459), .Z(n14452) );
  AND U14162 ( .A(n450), .B(n14451), .Z(n14459) );
  XNOR U14163 ( .A(n14449), .B(n14458), .Z(n14451) );
  XNOR U14164 ( .A(n14460), .B(n14461), .Z(n14449) );
  AND U14165 ( .A(n454), .B(n14462), .Z(n14461) );
  XOR U14166 ( .A(p_input[567]), .B(n14460), .Z(n14462) );
  XNOR U14167 ( .A(n14463), .B(n14464), .Z(n14460) );
  AND U14168 ( .A(n458), .B(n14465), .Z(n14464) );
  XOR U14169 ( .A(n14466), .B(n14467), .Z(n14458) );
  AND U14170 ( .A(n462), .B(n14457), .Z(n14467) );
  XNOR U14171 ( .A(n14468), .B(n14455), .Z(n14457) );
  XOR U14172 ( .A(n14469), .B(n14470), .Z(n14455) );
  AND U14173 ( .A(n485), .B(n14471), .Z(n14470) );
  IV U14174 ( .A(n14466), .Z(n14468) );
  XOR U14175 ( .A(n14472), .B(n14473), .Z(n14466) );
  AND U14176 ( .A(n469), .B(n14465), .Z(n14473) );
  XNOR U14177 ( .A(n14463), .B(n14472), .Z(n14465) );
  XNOR U14178 ( .A(n14474), .B(n14475), .Z(n14463) );
  AND U14179 ( .A(n473), .B(n14476), .Z(n14475) );
  XOR U14180 ( .A(p_input[599]), .B(n14474), .Z(n14476) );
  XNOR U14181 ( .A(n14477), .B(n14478), .Z(n14474) );
  AND U14182 ( .A(n477), .B(n14479), .Z(n14478) );
  XOR U14183 ( .A(n14480), .B(n14481), .Z(n14472) );
  AND U14184 ( .A(n481), .B(n14471), .Z(n14481) );
  XNOR U14185 ( .A(n14482), .B(n14469), .Z(n14471) );
  XOR U14186 ( .A(n14483), .B(n14484), .Z(n14469) );
  AND U14187 ( .A(n504), .B(n14485), .Z(n14484) );
  IV U14188 ( .A(n14480), .Z(n14482) );
  XOR U14189 ( .A(n14486), .B(n14487), .Z(n14480) );
  AND U14190 ( .A(n488), .B(n14479), .Z(n14487) );
  XNOR U14191 ( .A(n14477), .B(n14486), .Z(n14479) );
  XNOR U14192 ( .A(n14488), .B(n14489), .Z(n14477) );
  AND U14193 ( .A(n492), .B(n14490), .Z(n14489) );
  XOR U14194 ( .A(p_input[631]), .B(n14488), .Z(n14490) );
  XNOR U14195 ( .A(n14491), .B(n14492), .Z(n14488) );
  AND U14196 ( .A(n496), .B(n14493), .Z(n14492) );
  XOR U14197 ( .A(n14494), .B(n14495), .Z(n14486) );
  AND U14198 ( .A(n500), .B(n14485), .Z(n14495) );
  XNOR U14199 ( .A(n14496), .B(n14483), .Z(n14485) );
  XOR U14200 ( .A(n14497), .B(n14498), .Z(n14483) );
  AND U14201 ( .A(n523), .B(n14499), .Z(n14498) );
  IV U14202 ( .A(n14494), .Z(n14496) );
  XOR U14203 ( .A(n14500), .B(n14501), .Z(n14494) );
  AND U14204 ( .A(n507), .B(n14493), .Z(n14501) );
  XNOR U14205 ( .A(n14491), .B(n14500), .Z(n14493) );
  XNOR U14206 ( .A(n14502), .B(n14503), .Z(n14491) );
  AND U14207 ( .A(n511), .B(n14504), .Z(n14503) );
  XOR U14208 ( .A(p_input[663]), .B(n14502), .Z(n14504) );
  XNOR U14209 ( .A(n14505), .B(n14506), .Z(n14502) );
  AND U14210 ( .A(n515), .B(n14507), .Z(n14506) );
  XOR U14211 ( .A(n14508), .B(n14509), .Z(n14500) );
  AND U14212 ( .A(n519), .B(n14499), .Z(n14509) );
  XNOR U14213 ( .A(n14510), .B(n14497), .Z(n14499) );
  XOR U14214 ( .A(n14511), .B(n14512), .Z(n14497) );
  AND U14215 ( .A(n542), .B(n14513), .Z(n14512) );
  IV U14216 ( .A(n14508), .Z(n14510) );
  XOR U14217 ( .A(n14514), .B(n14515), .Z(n14508) );
  AND U14218 ( .A(n526), .B(n14507), .Z(n14515) );
  XNOR U14219 ( .A(n14505), .B(n14514), .Z(n14507) );
  XNOR U14220 ( .A(n14516), .B(n14517), .Z(n14505) );
  AND U14221 ( .A(n530), .B(n14518), .Z(n14517) );
  XOR U14222 ( .A(p_input[695]), .B(n14516), .Z(n14518) );
  XNOR U14223 ( .A(n14519), .B(n14520), .Z(n14516) );
  AND U14224 ( .A(n534), .B(n14521), .Z(n14520) );
  XOR U14225 ( .A(n14522), .B(n14523), .Z(n14514) );
  AND U14226 ( .A(n538), .B(n14513), .Z(n14523) );
  XNOR U14227 ( .A(n14524), .B(n14511), .Z(n14513) );
  XOR U14228 ( .A(n14525), .B(n14526), .Z(n14511) );
  AND U14229 ( .A(n561), .B(n14527), .Z(n14526) );
  IV U14230 ( .A(n14522), .Z(n14524) );
  XOR U14231 ( .A(n14528), .B(n14529), .Z(n14522) );
  AND U14232 ( .A(n545), .B(n14521), .Z(n14529) );
  XNOR U14233 ( .A(n14519), .B(n14528), .Z(n14521) );
  XNOR U14234 ( .A(n14530), .B(n14531), .Z(n14519) );
  AND U14235 ( .A(n549), .B(n14532), .Z(n14531) );
  XOR U14236 ( .A(p_input[727]), .B(n14530), .Z(n14532) );
  XNOR U14237 ( .A(n14533), .B(n14534), .Z(n14530) );
  AND U14238 ( .A(n553), .B(n14535), .Z(n14534) );
  XOR U14239 ( .A(n14536), .B(n14537), .Z(n14528) );
  AND U14240 ( .A(n557), .B(n14527), .Z(n14537) );
  XNOR U14241 ( .A(n14538), .B(n14525), .Z(n14527) );
  XOR U14242 ( .A(n14539), .B(n14540), .Z(n14525) );
  AND U14243 ( .A(n580), .B(n14541), .Z(n14540) );
  IV U14244 ( .A(n14536), .Z(n14538) );
  XOR U14245 ( .A(n14542), .B(n14543), .Z(n14536) );
  AND U14246 ( .A(n564), .B(n14535), .Z(n14543) );
  XNOR U14247 ( .A(n14533), .B(n14542), .Z(n14535) );
  XNOR U14248 ( .A(n14544), .B(n14545), .Z(n14533) );
  AND U14249 ( .A(n568), .B(n14546), .Z(n14545) );
  XOR U14250 ( .A(p_input[759]), .B(n14544), .Z(n14546) );
  XNOR U14251 ( .A(n14547), .B(n14548), .Z(n14544) );
  AND U14252 ( .A(n572), .B(n14549), .Z(n14548) );
  XOR U14253 ( .A(n14550), .B(n14551), .Z(n14542) );
  AND U14254 ( .A(n576), .B(n14541), .Z(n14551) );
  XNOR U14255 ( .A(n14552), .B(n14539), .Z(n14541) );
  XOR U14256 ( .A(n14553), .B(n14554), .Z(n14539) );
  AND U14257 ( .A(n599), .B(n14555), .Z(n14554) );
  IV U14258 ( .A(n14550), .Z(n14552) );
  XOR U14259 ( .A(n14556), .B(n14557), .Z(n14550) );
  AND U14260 ( .A(n583), .B(n14549), .Z(n14557) );
  XNOR U14261 ( .A(n14547), .B(n14556), .Z(n14549) );
  XNOR U14262 ( .A(n14558), .B(n14559), .Z(n14547) );
  AND U14263 ( .A(n587), .B(n14560), .Z(n14559) );
  XOR U14264 ( .A(p_input[791]), .B(n14558), .Z(n14560) );
  XNOR U14265 ( .A(n14561), .B(n14562), .Z(n14558) );
  AND U14266 ( .A(n591), .B(n14563), .Z(n14562) );
  XOR U14267 ( .A(n14564), .B(n14565), .Z(n14556) );
  AND U14268 ( .A(n595), .B(n14555), .Z(n14565) );
  XNOR U14269 ( .A(n14566), .B(n14553), .Z(n14555) );
  XOR U14270 ( .A(n14567), .B(n14568), .Z(n14553) );
  AND U14271 ( .A(n618), .B(n14569), .Z(n14568) );
  IV U14272 ( .A(n14564), .Z(n14566) );
  XOR U14273 ( .A(n14570), .B(n14571), .Z(n14564) );
  AND U14274 ( .A(n602), .B(n14563), .Z(n14571) );
  XNOR U14275 ( .A(n14561), .B(n14570), .Z(n14563) );
  XNOR U14276 ( .A(n14572), .B(n14573), .Z(n14561) );
  AND U14277 ( .A(n606), .B(n14574), .Z(n14573) );
  XOR U14278 ( .A(p_input[823]), .B(n14572), .Z(n14574) );
  XNOR U14279 ( .A(n14575), .B(n14576), .Z(n14572) );
  AND U14280 ( .A(n610), .B(n14577), .Z(n14576) );
  XOR U14281 ( .A(n14578), .B(n14579), .Z(n14570) );
  AND U14282 ( .A(n614), .B(n14569), .Z(n14579) );
  XNOR U14283 ( .A(n14580), .B(n14567), .Z(n14569) );
  XOR U14284 ( .A(n14581), .B(n14582), .Z(n14567) );
  AND U14285 ( .A(n637), .B(n14583), .Z(n14582) );
  IV U14286 ( .A(n14578), .Z(n14580) );
  XOR U14287 ( .A(n14584), .B(n14585), .Z(n14578) );
  AND U14288 ( .A(n621), .B(n14577), .Z(n14585) );
  XNOR U14289 ( .A(n14575), .B(n14584), .Z(n14577) );
  XNOR U14290 ( .A(n14586), .B(n14587), .Z(n14575) );
  AND U14291 ( .A(n625), .B(n14588), .Z(n14587) );
  XOR U14292 ( .A(p_input[855]), .B(n14586), .Z(n14588) );
  XNOR U14293 ( .A(n14589), .B(n14590), .Z(n14586) );
  AND U14294 ( .A(n629), .B(n14591), .Z(n14590) );
  XOR U14295 ( .A(n14592), .B(n14593), .Z(n14584) );
  AND U14296 ( .A(n633), .B(n14583), .Z(n14593) );
  XNOR U14297 ( .A(n14594), .B(n14581), .Z(n14583) );
  XOR U14298 ( .A(n14595), .B(n14596), .Z(n14581) );
  AND U14299 ( .A(n656), .B(n14597), .Z(n14596) );
  IV U14300 ( .A(n14592), .Z(n14594) );
  XOR U14301 ( .A(n14598), .B(n14599), .Z(n14592) );
  AND U14302 ( .A(n640), .B(n14591), .Z(n14599) );
  XNOR U14303 ( .A(n14589), .B(n14598), .Z(n14591) );
  XNOR U14304 ( .A(n14600), .B(n14601), .Z(n14589) );
  AND U14305 ( .A(n644), .B(n14602), .Z(n14601) );
  XOR U14306 ( .A(p_input[887]), .B(n14600), .Z(n14602) );
  XNOR U14307 ( .A(n14603), .B(n14604), .Z(n14600) );
  AND U14308 ( .A(n648), .B(n14605), .Z(n14604) );
  XOR U14309 ( .A(n14606), .B(n14607), .Z(n14598) );
  AND U14310 ( .A(n652), .B(n14597), .Z(n14607) );
  XNOR U14311 ( .A(n14608), .B(n14595), .Z(n14597) );
  XOR U14312 ( .A(n14609), .B(n14610), .Z(n14595) );
  AND U14313 ( .A(n675), .B(n14611), .Z(n14610) );
  IV U14314 ( .A(n14606), .Z(n14608) );
  XOR U14315 ( .A(n14612), .B(n14613), .Z(n14606) );
  AND U14316 ( .A(n659), .B(n14605), .Z(n14613) );
  XNOR U14317 ( .A(n14603), .B(n14612), .Z(n14605) );
  XNOR U14318 ( .A(n14614), .B(n14615), .Z(n14603) );
  AND U14319 ( .A(n663), .B(n14616), .Z(n14615) );
  XOR U14320 ( .A(p_input[919]), .B(n14614), .Z(n14616) );
  XNOR U14321 ( .A(n14617), .B(n14618), .Z(n14614) );
  AND U14322 ( .A(n667), .B(n14619), .Z(n14618) );
  XOR U14323 ( .A(n14620), .B(n14621), .Z(n14612) );
  AND U14324 ( .A(n671), .B(n14611), .Z(n14621) );
  XNOR U14325 ( .A(n14622), .B(n14609), .Z(n14611) );
  XOR U14326 ( .A(n14623), .B(n14624), .Z(n14609) );
  AND U14327 ( .A(n694), .B(n14625), .Z(n14624) );
  IV U14328 ( .A(n14620), .Z(n14622) );
  XOR U14329 ( .A(n14626), .B(n14627), .Z(n14620) );
  AND U14330 ( .A(n678), .B(n14619), .Z(n14627) );
  XNOR U14331 ( .A(n14617), .B(n14626), .Z(n14619) );
  XNOR U14332 ( .A(n14628), .B(n14629), .Z(n14617) );
  AND U14333 ( .A(n682), .B(n14630), .Z(n14629) );
  XOR U14334 ( .A(p_input[951]), .B(n14628), .Z(n14630) );
  XNOR U14335 ( .A(n14631), .B(n14632), .Z(n14628) );
  AND U14336 ( .A(n686), .B(n14633), .Z(n14632) );
  XOR U14337 ( .A(n14634), .B(n14635), .Z(n14626) );
  AND U14338 ( .A(n690), .B(n14625), .Z(n14635) );
  XNOR U14339 ( .A(n14636), .B(n14623), .Z(n14625) );
  XOR U14340 ( .A(n14637), .B(n14638), .Z(n14623) );
  AND U14341 ( .A(n713), .B(n14639), .Z(n14638) );
  IV U14342 ( .A(n14634), .Z(n14636) );
  XOR U14343 ( .A(n14640), .B(n14641), .Z(n14634) );
  AND U14344 ( .A(n697), .B(n14633), .Z(n14641) );
  XNOR U14345 ( .A(n14631), .B(n14640), .Z(n14633) );
  XNOR U14346 ( .A(n14642), .B(n14643), .Z(n14631) );
  AND U14347 ( .A(n701), .B(n14644), .Z(n14643) );
  XOR U14348 ( .A(p_input[983]), .B(n14642), .Z(n14644) );
  XNOR U14349 ( .A(n14645), .B(n14646), .Z(n14642) );
  AND U14350 ( .A(n705), .B(n14647), .Z(n14646) );
  XOR U14351 ( .A(n14648), .B(n14649), .Z(n14640) );
  AND U14352 ( .A(n709), .B(n14639), .Z(n14649) );
  XNOR U14353 ( .A(n14650), .B(n14637), .Z(n14639) );
  XOR U14354 ( .A(n14651), .B(n14652), .Z(n14637) );
  AND U14355 ( .A(n732), .B(n14653), .Z(n14652) );
  IV U14356 ( .A(n14648), .Z(n14650) );
  XOR U14357 ( .A(n14654), .B(n14655), .Z(n14648) );
  AND U14358 ( .A(n716), .B(n14647), .Z(n14655) );
  XNOR U14359 ( .A(n14645), .B(n14654), .Z(n14647) );
  XNOR U14360 ( .A(n14656), .B(n14657), .Z(n14645) );
  AND U14361 ( .A(n720), .B(n14658), .Z(n14657) );
  XOR U14362 ( .A(p_input[1015]), .B(n14656), .Z(n14658) );
  XNOR U14363 ( .A(n14659), .B(n14660), .Z(n14656) );
  AND U14364 ( .A(n724), .B(n14661), .Z(n14660) );
  XOR U14365 ( .A(n14662), .B(n14663), .Z(n14654) );
  AND U14366 ( .A(n728), .B(n14653), .Z(n14663) );
  XNOR U14367 ( .A(n14664), .B(n14651), .Z(n14653) );
  XOR U14368 ( .A(n14665), .B(n14666), .Z(n14651) );
  AND U14369 ( .A(n751), .B(n14667), .Z(n14666) );
  IV U14370 ( .A(n14662), .Z(n14664) );
  XOR U14371 ( .A(n14668), .B(n14669), .Z(n14662) );
  AND U14372 ( .A(n735), .B(n14661), .Z(n14669) );
  XNOR U14373 ( .A(n14659), .B(n14668), .Z(n14661) );
  XNOR U14374 ( .A(n14670), .B(n14671), .Z(n14659) );
  AND U14375 ( .A(n739), .B(n14672), .Z(n14671) );
  XOR U14376 ( .A(p_input[1047]), .B(n14670), .Z(n14672) );
  XNOR U14377 ( .A(n14673), .B(n14674), .Z(n14670) );
  AND U14378 ( .A(n743), .B(n14675), .Z(n14674) );
  XOR U14379 ( .A(n14676), .B(n14677), .Z(n14668) );
  AND U14380 ( .A(n747), .B(n14667), .Z(n14677) );
  XNOR U14381 ( .A(n14678), .B(n14665), .Z(n14667) );
  XOR U14382 ( .A(n14679), .B(n14680), .Z(n14665) );
  AND U14383 ( .A(n770), .B(n14681), .Z(n14680) );
  IV U14384 ( .A(n14676), .Z(n14678) );
  XOR U14385 ( .A(n14682), .B(n14683), .Z(n14676) );
  AND U14386 ( .A(n754), .B(n14675), .Z(n14683) );
  XNOR U14387 ( .A(n14673), .B(n14682), .Z(n14675) );
  XNOR U14388 ( .A(n14684), .B(n14685), .Z(n14673) );
  AND U14389 ( .A(n758), .B(n14686), .Z(n14685) );
  XOR U14390 ( .A(p_input[1079]), .B(n14684), .Z(n14686) );
  XNOR U14391 ( .A(n14687), .B(n14688), .Z(n14684) );
  AND U14392 ( .A(n762), .B(n14689), .Z(n14688) );
  XOR U14393 ( .A(n14690), .B(n14691), .Z(n14682) );
  AND U14394 ( .A(n766), .B(n14681), .Z(n14691) );
  XNOR U14395 ( .A(n14692), .B(n14679), .Z(n14681) );
  XOR U14396 ( .A(n14693), .B(n14694), .Z(n14679) );
  AND U14397 ( .A(n789), .B(n14695), .Z(n14694) );
  IV U14398 ( .A(n14690), .Z(n14692) );
  XOR U14399 ( .A(n14696), .B(n14697), .Z(n14690) );
  AND U14400 ( .A(n773), .B(n14689), .Z(n14697) );
  XNOR U14401 ( .A(n14687), .B(n14696), .Z(n14689) );
  XNOR U14402 ( .A(n14698), .B(n14699), .Z(n14687) );
  AND U14403 ( .A(n777), .B(n14700), .Z(n14699) );
  XOR U14404 ( .A(p_input[1111]), .B(n14698), .Z(n14700) );
  XNOR U14405 ( .A(n14701), .B(n14702), .Z(n14698) );
  AND U14406 ( .A(n781), .B(n14703), .Z(n14702) );
  XOR U14407 ( .A(n14704), .B(n14705), .Z(n14696) );
  AND U14408 ( .A(n785), .B(n14695), .Z(n14705) );
  XNOR U14409 ( .A(n14706), .B(n14693), .Z(n14695) );
  XOR U14410 ( .A(n14707), .B(n14708), .Z(n14693) );
  AND U14411 ( .A(n808), .B(n14709), .Z(n14708) );
  IV U14412 ( .A(n14704), .Z(n14706) );
  XOR U14413 ( .A(n14710), .B(n14711), .Z(n14704) );
  AND U14414 ( .A(n792), .B(n14703), .Z(n14711) );
  XNOR U14415 ( .A(n14701), .B(n14710), .Z(n14703) );
  XNOR U14416 ( .A(n14712), .B(n14713), .Z(n14701) );
  AND U14417 ( .A(n796), .B(n14714), .Z(n14713) );
  XOR U14418 ( .A(p_input[1143]), .B(n14712), .Z(n14714) );
  XNOR U14419 ( .A(n14715), .B(n14716), .Z(n14712) );
  AND U14420 ( .A(n800), .B(n14717), .Z(n14716) );
  XOR U14421 ( .A(n14718), .B(n14719), .Z(n14710) );
  AND U14422 ( .A(n804), .B(n14709), .Z(n14719) );
  XNOR U14423 ( .A(n14720), .B(n14707), .Z(n14709) );
  XOR U14424 ( .A(n14721), .B(n14722), .Z(n14707) );
  AND U14425 ( .A(n827), .B(n14723), .Z(n14722) );
  IV U14426 ( .A(n14718), .Z(n14720) );
  XOR U14427 ( .A(n14724), .B(n14725), .Z(n14718) );
  AND U14428 ( .A(n811), .B(n14717), .Z(n14725) );
  XNOR U14429 ( .A(n14715), .B(n14724), .Z(n14717) );
  XNOR U14430 ( .A(n14726), .B(n14727), .Z(n14715) );
  AND U14431 ( .A(n815), .B(n14728), .Z(n14727) );
  XOR U14432 ( .A(p_input[1175]), .B(n14726), .Z(n14728) );
  XNOR U14433 ( .A(n14729), .B(n14730), .Z(n14726) );
  AND U14434 ( .A(n819), .B(n14731), .Z(n14730) );
  XOR U14435 ( .A(n14732), .B(n14733), .Z(n14724) );
  AND U14436 ( .A(n823), .B(n14723), .Z(n14733) );
  XNOR U14437 ( .A(n14734), .B(n14721), .Z(n14723) );
  XOR U14438 ( .A(n14735), .B(n14736), .Z(n14721) );
  AND U14439 ( .A(n846), .B(n14737), .Z(n14736) );
  IV U14440 ( .A(n14732), .Z(n14734) );
  XOR U14441 ( .A(n14738), .B(n14739), .Z(n14732) );
  AND U14442 ( .A(n830), .B(n14731), .Z(n14739) );
  XNOR U14443 ( .A(n14729), .B(n14738), .Z(n14731) );
  XNOR U14444 ( .A(n14740), .B(n14741), .Z(n14729) );
  AND U14445 ( .A(n834), .B(n14742), .Z(n14741) );
  XOR U14446 ( .A(p_input[1207]), .B(n14740), .Z(n14742) );
  XNOR U14447 ( .A(n14743), .B(n14744), .Z(n14740) );
  AND U14448 ( .A(n838), .B(n14745), .Z(n14744) );
  XOR U14449 ( .A(n14746), .B(n14747), .Z(n14738) );
  AND U14450 ( .A(n842), .B(n14737), .Z(n14747) );
  XNOR U14451 ( .A(n14748), .B(n14735), .Z(n14737) );
  XOR U14452 ( .A(n14749), .B(n14750), .Z(n14735) );
  AND U14453 ( .A(n865), .B(n14751), .Z(n14750) );
  IV U14454 ( .A(n14746), .Z(n14748) );
  XOR U14455 ( .A(n14752), .B(n14753), .Z(n14746) );
  AND U14456 ( .A(n849), .B(n14745), .Z(n14753) );
  XNOR U14457 ( .A(n14743), .B(n14752), .Z(n14745) );
  XNOR U14458 ( .A(n14754), .B(n14755), .Z(n14743) );
  AND U14459 ( .A(n853), .B(n14756), .Z(n14755) );
  XOR U14460 ( .A(p_input[1239]), .B(n14754), .Z(n14756) );
  XNOR U14461 ( .A(n14757), .B(n14758), .Z(n14754) );
  AND U14462 ( .A(n857), .B(n14759), .Z(n14758) );
  XOR U14463 ( .A(n14760), .B(n14761), .Z(n14752) );
  AND U14464 ( .A(n861), .B(n14751), .Z(n14761) );
  XNOR U14465 ( .A(n14762), .B(n14749), .Z(n14751) );
  XOR U14466 ( .A(n14763), .B(n14764), .Z(n14749) );
  AND U14467 ( .A(n884), .B(n14765), .Z(n14764) );
  IV U14468 ( .A(n14760), .Z(n14762) );
  XOR U14469 ( .A(n14766), .B(n14767), .Z(n14760) );
  AND U14470 ( .A(n868), .B(n14759), .Z(n14767) );
  XNOR U14471 ( .A(n14757), .B(n14766), .Z(n14759) );
  XNOR U14472 ( .A(n14768), .B(n14769), .Z(n14757) );
  AND U14473 ( .A(n872), .B(n14770), .Z(n14769) );
  XOR U14474 ( .A(p_input[1271]), .B(n14768), .Z(n14770) );
  XNOR U14475 ( .A(n14771), .B(n14772), .Z(n14768) );
  AND U14476 ( .A(n876), .B(n14773), .Z(n14772) );
  XOR U14477 ( .A(n14774), .B(n14775), .Z(n14766) );
  AND U14478 ( .A(n880), .B(n14765), .Z(n14775) );
  XNOR U14479 ( .A(n14776), .B(n14763), .Z(n14765) );
  XOR U14480 ( .A(n14777), .B(n14778), .Z(n14763) );
  AND U14481 ( .A(n903), .B(n14779), .Z(n14778) );
  IV U14482 ( .A(n14774), .Z(n14776) );
  XOR U14483 ( .A(n14780), .B(n14781), .Z(n14774) );
  AND U14484 ( .A(n887), .B(n14773), .Z(n14781) );
  XNOR U14485 ( .A(n14771), .B(n14780), .Z(n14773) );
  XNOR U14486 ( .A(n14782), .B(n14783), .Z(n14771) );
  AND U14487 ( .A(n891), .B(n14784), .Z(n14783) );
  XOR U14488 ( .A(p_input[1303]), .B(n14782), .Z(n14784) );
  XNOR U14489 ( .A(n14785), .B(n14786), .Z(n14782) );
  AND U14490 ( .A(n895), .B(n14787), .Z(n14786) );
  XOR U14491 ( .A(n14788), .B(n14789), .Z(n14780) );
  AND U14492 ( .A(n899), .B(n14779), .Z(n14789) );
  XNOR U14493 ( .A(n14790), .B(n14777), .Z(n14779) );
  XOR U14494 ( .A(n14791), .B(n14792), .Z(n14777) );
  AND U14495 ( .A(n922), .B(n14793), .Z(n14792) );
  IV U14496 ( .A(n14788), .Z(n14790) );
  XOR U14497 ( .A(n14794), .B(n14795), .Z(n14788) );
  AND U14498 ( .A(n906), .B(n14787), .Z(n14795) );
  XNOR U14499 ( .A(n14785), .B(n14794), .Z(n14787) );
  XNOR U14500 ( .A(n14796), .B(n14797), .Z(n14785) );
  AND U14501 ( .A(n910), .B(n14798), .Z(n14797) );
  XOR U14502 ( .A(p_input[1335]), .B(n14796), .Z(n14798) );
  XNOR U14503 ( .A(n14799), .B(n14800), .Z(n14796) );
  AND U14504 ( .A(n914), .B(n14801), .Z(n14800) );
  XOR U14505 ( .A(n14802), .B(n14803), .Z(n14794) );
  AND U14506 ( .A(n918), .B(n14793), .Z(n14803) );
  XNOR U14507 ( .A(n14804), .B(n14791), .Z(n14793) );
  XOR U14508 ( .A(n14805), .B(n14806), .Z(n14791) );
  AND U14509 ( .A(n941), .B(n14807), .Z(n14806) );
  IV U14510 ( .A(n14802), .Z(n14804) );
  XOR U14511 ( .A(n14808), .B(n14809), .Z(n14802) );
  AND U14512 ( .A(n925), .B(n14801), .Z(n14809) );
  XNOR U14513 ( .A(n14799), .B(n14808), .Z(n14801) );
  XNOR U14514 ( .A(n14810), .B(n14811), .Z(n14799) );
  AND U14515 ( .A(n929), .B(n14812), .Z(n14811) );
  XOR U14516 ( .A(p_input[1367]), .B(n14810), .Z(n14812) );
  XNOR U14517 ( .A(n14813), .B(n14814), .Z(n14810) );
  AND U14518 ( .A(n933), .B(n14815), .Z(n14814) );
  XOR U14519 ( .A(n14816), .B(n14817), .Z(n14808) );
  AND U14520 ( .A(n937), .B(n14807), .Z(n14817) );
  XNOR U14521 ( .A(n14818), .B(n14805), .Z(n14807) );
  XOR U14522 ( .A(n14819), .B(n14820), .Z(n14805) );
  AND U14523 ( .A(n960), .B(n14821), .Z(n14820) );
  IV U14524 ( .A(n14816), .Z(n14818) );
  XOR U14525 ( .A(n14822), .B(n14823), .Z(n14816) );
  AND U14526 ( .A(n944), .B(n14815), .Z(n14823) );
  XNOR U14527 ( .A(n14813), .B(n14822), .Z(n14815) );
  XNOR U14528 ( .A(n14824), .B(n14825), .Z(n14813) );
  AND U14529 ( .A(n948), .B(n14826), .Z(n14825) );
  XOR U14530 ( .A(p_input[1399]), .B(n14824), .Z(n14826) );
  XNOR U14531 ( .A(n14827), .B(n14828), .Z(n14824) );
  AND U14532 ( .A(n952), .B(n14829), .Z(n14828) );
  XOR U14533 ( .A(n14830), .B(n14831), .Z(n14822) );
  AND U14534 ( .A(n956), .B(n14821), .Z(n14831) );
  XNOR U14535 ( .A(n14832), .B(n14819), .Z(n14821) );
  XOR U14536 ( .A(n14833), .B(n14834), .Z(n14819) );
  AND U14537 ( .A(n979), .B(n14835), .Z(n14834) );
  IV U14538 ( .A(n14830), .Z(n14832) );
  XOR U14539 ( .A(n14836), .B(n14837), .Z(n14830) );
  AND U14540 ( .A(n963), .B(n14829), .Z(n14837) );
  XNOR U14541 ( .A(n14827), .B(n14836), .Z(n14829) );
  XNOR U14542 ( .A(n14838), .B(n14839), .Z(n14827) );
  AND U14543 ( .A(n967), .B(n14840), .Z(n14839) );
  XOR U14544 ( .A(p_input[1431]), .B(n14838), .Z(n14840) );
  XNOR U14545 ( .A(n14841), .B(n14842), .Z(n14838) );
  AND U14546 ( .A(n971), .B(n14843), .Z(n14842) );
  XOR U14547 ( .A(n14844), .B(n14845), .Z(n14836) );
  AND U14548 ( .A(n975), .B(n14835), .Z(n14845) );
  XNOR U14549 ( .A(n14846), .B(n14833), .Z(n14835) );
  XOR U14550 ( .A(n14847), .B(n14848), .Z(n14833) );
  AND U14551 ( .A(n998), .B(n14849), .Z(n14848) );
  IV U14552 ( .A(n14844), .Z(n14846) );
  XOR U14553 ( .A(n14850), .B(n14851), .Z(n14844) );
  AND U14554 ( .A(n982), .B(n14843), .Z(n14851) );
  XNOR U14555 ( .A(n14841), .B(n14850), .Z(n14843) );
  XNOR U14556 ( .A(n14852), .B(n14853), .Z(n14841) );
  AND U14557 ( .A(n986), .B(n14854), .Z(n14853) );
  XOR U14558 ( .A(p_input[1463]), .B(n14852), .Z(n14854) );
  XNOR U14559 ( .A(n14855), .B(n14856), .Z(n14852) );
  AND U14560 ( .A(n990), .B(n14857), .Z(n14856) );
  XOR U14561 ( .A(n14858), .B(n14859), .Z(n14850) );
  AND U14562 ( .A(n994), .B(n14849), .Z(n14859) );
  XNOR U14563 ( .A(n14860), .B(n14847), .Z(n14849) );
  XOR U14564 ( .A(n14861), .B(n14862), .Z(n14847) );
  AND U14565 ( .A(n1017), .B(n14863), .Z(n14862) );
  IV U14566 ( .A(n14858), .Z(n14860) );
  XOR U14567 ( .A(n14864), .B(n14865), .Z(n14858) );
  AND U14568 ( .A(n1001), .B(n14857), .Z(n14865) );
  XNOR U14569 ( .A(n14855), .B(n14864), .Z(n14857) );
  XNOR U14570 ( .A(n14866), .B(n14867), .Z(n14855) );
  AND U14571 ( .A(n1005), .B(n14868), .Z(n14867) );
  XOR U14572 ( .A(p_input[1495]), .B(n14866), .Z(n14868) );
  XNOR U14573 ( .A(n14869), .B(n14870), .Z(n14866) );
  AND U14574 ( .A(n1009), .B(n14871), .Z(n14870) );
  XOR U14575 ( .A(n14872), .B(n14873), .Z(n14864) );
  AND U14576 ( .A(n1013), .B(n14863), .Z(n14873) );
  XNOR U14577 ( .A(n14874), .B(n14861), .Z(n14863) );
  XOR U14578 ( .A(n14875), .B(n14876), .Z(n14861) );
  AND U14579 ( .A(n1036), .B(n14877), .Z(n14876) );
  IV U14580 ( .A(n14872), .Z(n14874) );
  XOR U14581 ( .A(n14878), .B(n14879), .Z(n14872) );
  AND U14582 ( .A(n1020), .B(n14871), .Z(n14879) );
  XNOR U14583 ( .A(n14869), .B(n14878), .Z(n14871) );
  XNOR U14584 ( .A(n14880), .B(n14881), .Z(n14869) );
  AND U14585 ( .A(n1024), .B(n14882), .Z(n14881) );
  XOR U14586 ( .A(p_input[1527]), .B(n14880), .Z(n14882) );
  XNOR U14587 ( .A(n14883), .B(n14884), .Z(n14880) );
  AND U14588 ( .A(n1028), .B(n14885), .Z(n14884) );
  XOR U14589 ( .A(n14886), .B(n14887), .Z(n14878) );
  AND U14590 ( .A(n1032), .B(n14877), .Z(n14887) );
  XNOR U14591 ( .A(n14888), .B(n14875), .Z(n14877) );
  XOR U14592 ( .A(n14889), .B(n14890), .Z(n14875) );
  AND U14593 ( .A(n1055), .B(n14891), .Z(n14890) );
  IV U14594 ( .A(n14886), .Z(n14888) );
  XOR U14595 ( .A(n14892), .B(n14893), .Z(n14886) );
  AND U14596 ( .A(n1039), .B(n14885), .Z(n14893) );
  XNOR U14597 ( .A(n14883), .B(n14892), .Z(n14885) );
  XNOR U14598 ( .A(n14894), .B(n14895), .Z(n14883) );
  AND U14599 ( .A(n1043), .B(n14896), .Z(n14895) );
  XOR U14600 ( .A(p_input[1559]), .B(n14894), .Z(n14896) );
  XNOR U14601 ( .A(n14897), .B(n14898), .Z(n14894) );
  AND U14602 ( .A(n1047), .B(n14899), .Z(n14898) );
  XOR U14603 ( .A(n14900), .B(n14901), .Z(n14892) );
  AND U14604 ( .A(n1051), .B(n14891), .Z(n14901) );
  XNOR U14605 ( .A(n14902), .B(n14889), .Z(n14891) );
  XOR U14606 ( .A(n14903), .B(n14904), .Z(n14889) );
  AND U14607 ( .A(n1074), .B(n14905), .Z(n14904) );
  IV U14608 ( .A(n14900), .Z(n14902) );
  XOR U14609 ( .A(n14906), .B(n14907), .Z(n14900) );
  AND U14610 ( .A(n1058), .B(n14899), .Z(n14907) );
  XNOR U14611 ( .A(n14897), .B(n14906), .Z(n14899) );
  XNOR U14612 ( .A(n14908), .B(n14909), .Z(n14897) );
  AND U14613 ( .A(n1062), .B(n14910), .Z(n14909) );
  XOR U14614 ( .A(p_input[1591]), .B(n14908), .Z(n14910) );
  XNOR U14615 ( .A(n14911), .B(n14912), .Z(n14908) );
  AND U14616 ( .A(n1066), .B(n14913), .Z(n14912) );
  XOR U14617 ( .A(n14914), .B(n14915), .Z(n14906) );
  AND U14618 ( .A(n1070), .B(n14905), .Z(n14915) );
  XNOR U14619 ( .A(n14916), .B(n14903), .Z(n14905) );
  XOR U14620 ( .A(n14917), .B(n14918), .Z(n14903) );
  AND U14621 ( .A(n1093), .B(n14919), .Z(n14918) );
  IV U14622 ( .A(n14914), .Z(n14916) );
  XOR U14623 ( .A(n14920), .B(n14921), .Z(n14914) );
  AND U14624 ( .A(n1077), .B(n14913), .Z(n14921) );
  XNOR U14625 ( .A(n14911), .B(n14920), .Z(n14913) );
  XNOR U14626 ( .A(n14922), .B(n14923), .Z(n14911) );
  AND U14627 ( .A(n1081), .B(n14924), .Z(n14923) );
  XOR U14628 ( .A(p_input[1623]), .B(n14922), .Z(n14924) );
  XNOR U14629 ( .A(n14925), .B(n14926), .Z(n14922) );
  AND U14630 ( .A(n1085), .B(n14927), .Z(n14926) );
  XOR U14631 ( .A(n14928), .B(n14929), .Z(n14920) );
  AND U14632 ( .A(n1089), .B(n14919), .Z(n14929) );
  XNOR U14633 ( .A(n14930), .B(n14917), .Z(n14919) );
  XOR U14634 ( .A(n14931), .B(n14932), .Z(n14917) );
  AND U14635 ( .A(n1112), .B(n14933), .Z(n14932) );
  IV U14636 ( .A(n14928), .Z(n14930) );
  XOR U14637 ( .A(n14934), .B(n14935), .Z(n14928) );
  AND U14638 ( .A(n1096), .B(n14927), .Z(n14935) );
  XNOR U14639 ( .A(n14925), .B(n14934), .Z(n14927) );
  XNOR U14640 ( .A(n14936), .B(n14937), .Z(n14925) );
  AND U14641 ( .A(n1100), .B(n14938), .Z(n14937) );
  XOR U14642 ( .A(p_input[1655]), .B(n14936), .Z(n14938) );
  XNOR U14643 ( .A(n14939), .B(n14940), .Z(n14936) );
  AND U14644 ( .A(n1104), .B(n14941), .Z(n14940) );
  XOR U14645 ( .A(n14942), .B(n14943), .Z(n14934) );
  AND U14646 ( .A(n1108), .B(n14933), .Z(n14943) );
  XNOR U14647 ( .A(n14944), .B(n14931), .Z(n14933) );
  XOR U14648 ( .A(n14945), .B(n14946), .Z(n14931) );
  AND U14649 ( .A(n1131), .B(n14947), .Z(n14946) );
  IV U14650 ( .A(n14942), .Z(n14944) );
  XOR U14651 ( .A(n14948), .B(n14949), .Z(n14942) );
  AND U14652 ( .A(n1115), .B(n14941), .Z(n14949) );
  XNOR U14653 ( .A(n14939), .B(n14948), .Z(n14941) );
  XNOR U14654 ( .A(n14950), .B(n14951), .Z(n14939) );
  AND U14655 ( .A(n1119), .B(n14952), .Z(n14951) );
  XOR U14656 ( .A(p_input[1687]), .B(n14950), .Z(n14952) );
  XNOR U14657 ( .A(n14953), .B(n14954), .Z(n14950) );
  AND U14658 ( .A(n1123), .B(n14955), .Z(n14954) );
  XOR U14659 ( .A(n14956), .B(n14957), .Z(n14948) );
  AND U14660 ( .A(n1127), .B(n14947), .Z(n14957) );
  XNOR U14661 ( .A(n14958), .B(n14945), .Z(n14947) );
  XOR U14662 ( .A(n14959), .B(n14960), .Z(n14945) );
  AND U14663 ( .A(n1150), .B(n14961), .Z(n14960) );
  IV U14664 ( .A(n14956), .Z(n14958) );
  XOR U14665 ( .A(n14962), .B(n14963), .Z(n14956) );
  AND U14666 ( .A(n1134), .B(n14955), .Z(n14963) );
  XNOR U14667 ( .A(n14953), .B(n14962), .Z(n14955) );
  XNOR U14668 ( .A(n14964), .B(n14965), .Z(n14953) );
  AND U14669 ( .A(n1138), .B(n14966), .Z(n14965) );
  XOR U14670 ( .A(p_input[1719]), .B(n14964), .Z(n14966) );
  XNOR U14671 ( .A(n14967), .B(n14968), .Z(n14964) );
  AND U14672 ( .A(n1142), .B(n14969), .Z(n14968) );
  XOR U14673 ( .A(n14970), .B(n14971), .Z(n14962) );
  AND U14674 ( .A(n1146), .B(n14961), .Z(n14971) );
  XNOR U14675 ( .A(n14972), .B(n14959), .Z(n14961) );
  XOR U14676 ( .A(n14973), .B(n14974), .Z(n14959) );
  AND U14677 ( .A(n1169), .B(n14975), .Z(n14974) );
  IV U14678 ( .A(n14970), .Z(n14972) );
  XOR U14679 ( .A(n14976), .B(n14977), .Z(n14970) );
  AND U14680 ( .A(n1153), .B(n14969), .Z(n14977) );
  XNOR U14681 ( .A(n14967), .B(n14976), .Z(n14969) );
  XNOR U14682 ( .A(n14978), .B(n14979), .Z(n14967) );
  AND U14683 ( .A(n1157), .B(n14980), .Z(n14979) );
  XOR U14684 ( .A(p_input[1751]), .B(n14978), .Z(n14980) );
  XNOR U14685 ( .A(n14981), .B(n14982), .Z(n14978) );
  AND U14686 ( .A(n1161), .B(n14983), .Z(n14982) );
  XOR U14687 ( .A(n14984), .B(n14985), .Z(n14976) );
  AND U14688 ( .A(n1165), .B(n14975), .Z(n14985) );
  XNOR U14689 ( .A(n14986), .B(n14973), .Z(n14975) );
  XOR U14690 ( .A(n14987), .B(n14988), .Z(n14973) );
  AND U14691 ( .A(n1188), .B(n14989), .Z(n14988) );
  IV U14692 ( .A(n14984), .Z(n14986) );
  XOR U14693 ( .A(n14990), .B(n14991), .Z(n14984) );
  AND U14694 ( .A(n1172), .B(n14983), .Z(n14991) );
  XNOR U14695 ( .A(n14981), .B(n14990), .Z(n14983) );
  XNOR U14696 ( .A(n14992), .B(n14993), .Z(n14981) );
  AND U14697 ( .A(n1176), .B(n14994), .Z(n14993) );
  XOR U14698 ( .A(p_input[1783]), .B(n14992), .Z(n14994) );
  XNOR U14699 ( .A(n14995), .B(n14996), .Z(n14992) );
  AND U14700 ( .A(n1180), .B(n14997), .Z(n14996) );
  XOR U14701 ( .A(n14998), .B(n14999), .Z(n14990) );
  AND U14702 ( .A(n1184), .B(n14989), .Z(n14999) );
  XNOR U14703 ( .A(n15000), .B(n14987), .Z(n14989) );
  XOR U14704 ( .A(n15001), .B(n15002), .Z(n14987) );
  AND U14705 ( .A(n1207), .B(n15003), .Z(n15002) );
  IV U14706 ( .A(n14998), .Z(n15000) );
  XOR U14707 ( .A(n15004), .B(n15005), .Z(n14998) );
  AND U14708 ( .A(n1191), .B(n14997), .Z(n15005) );
  XNOR U14709 ( .A(n14995), .B(n15004), .Z(n14997) );
  XNOR U14710 ( .A(n15006), .B(n15007), .Z(n14995) );
  AND U14711 ( .A(n1195), .B(n15008), .Z(n15007) );
  XOR U14712 ( .A(p_input[1815]), .B(n15006), .Z(n15008) );
  XNOR U14713 ( .A(n15009), .B(n15010), .Z(n15006) );
  AND U14714 ( .A(n1199), .B(n15011), .Z(n15010) );
  XOR U14715 ( .A(n15012), .B(n15013), .Z(n15004) );
  AND U14716 ( .A(n1203), .B(n15003), .Z(n15013) );
  XNOR U14717 ( .A(n15014), .B(n15001), .Z(n15003) );
  XOR U14718 ( .A(n15015), .B(n15016), .Z(n15001) );
  AND U14719 ( .A(n1226), .B(n15017), .Z(n15016) );
  IV U14720 ( .A(n15012), .Z(n15014) );
  XOR U14721 ( .A(n15018), .B(n15019), .Z(n15012) );
  AND U14722 ( .A(n1210), .B(n15011), .Z(n15019) );
  XNOR U14723 ( .A(n15009), .B(n15018), .Z(n15011) );
  XNOR U14724 ( .A(n15020), .B(n15021), .Z(n15009) );
  AND U14725 ( .A(n1214), .B(n15022), .Z(n15021) );
  XOR U14726 ( .A(p_input[1847]), .B(n15020), .Z(n15022) );
  XNOR U14727 ( .A(n15023), .B(n15024), .Z(n15020) );
  AND U14728 ( .A(n1218), .B(n15025), .Z(n15024) );
  XOR U14729 ( .A(n15026), .B(n15027), .Z(n15018) );
  AND U14730 ( .A(n1222), .B(n15017), .Z(n15027) );
  XNOR U14731 ( .A(n15028), .B(n15015), .Z(n15017) );
  XOR U14732 ( .A(n15029), .B(n15030), .Z(n15015) );
  AND U14733 ( .A(n1245), .B(n15031), .Z(n15030) );
  IV U14734 ( .A(n15026), .Z(n15028) );
  XOR U14735 ( .A(n15032), .B(n15033), .Z(n15026) );
  AND U14736 ( .A(n1229), .B(n15025), .Z(n15033) );
  XNOR U14737 ( .A(n15023), .B(n15032), .Z(n15025) );
  XNOR U14738 ( .A(n15034), .B(n15035), .Z(n15023) );
  AND U14739 ( .A(n1233), .B(n15036), .Z(n15035) );
  XOR U14740 ( .A(p_input[1879]), .B(n15034), .Z(n15036) );
  XNOR U14741 ( .A(n15037), .B(n15038), .Z(n15034) );
  AND U14742 ( .A(n1237), .B(n15039), .Z(n15038) );
  XOR U14743 ( .A(n15040), .B(n15041), .Z(n15032) );
  AND U14744 ( .A(n1241), .B(n15031), .Z(n15041) );
  XNOR U14745 ( .A(n15042), .B(n15029), .Z(n15031) );
  XOR U14746 ( .A(n15043), .B(n15044), .Z(n15029) );
  AND U14747 ( .A(n1264), .B(n15045), .Z(n15044) );
  IV U14748 ( .A(n15040), .Z(n15042) );
  XOR U14749 ( .A(n15046), .B(n15047), .Z(n15040) );
  AND U14750 ( .A(n1248), .B(n15039), .Z(n15047) );
  XNOR U14751 ( .A(n15037), .B(n15046), .Z(n15039) );
  XNOR U14752 ( .A(n15048), .B(n15049), .Z(n15037) );
  AND U14753 ( .A(n1252), .B(n15050), .Z(n15049) );
  XOR U14754 ( .A(p_input[1911]), .B(n15048), .Z(n15050) );
  XNOR U14755 ( .A(n15051), .B(n15052), .Z(n15048) );
  AND U14756 ( .A(n1256), .B(n15053), .Z(n15052) );
  XOR U14757 ( .A(n15054), .B(n15055), .Z(n15046) );
  AND U14758 ( .A(n1260), .B(n15045), .Z(n15055) );
  XNOR U14759 ( .A(n15056), .B(n15043), .Z(n15045) );
  XOR U14760 ( .A(n15057), .B(n15058), .Z(n15043) );
  AND U14761 ( .A(n1282), .B(n15059), .Z(n15058) );
  IV U14762 ( .A(n15054), .Z(n15056) );
  XOR U14763 ( .A(n15060), .B(n15061), .Z(n15054) );
  AND U14764 ( .A(n1267), .B(n15053), .Z(n15061) );
  XNOR U14765 ( .A(n15051), .B(n15060), .Z(n15053) );
  XNOR U14766 ( .A(n15062), .B(n15063), .Z(n15051) );
  AND U14767 ( .A(n1271), .B(n15064), .Z(n15063) );
  XOR U14768 ( .A(p_input[1943]), .B(n15062), .Z(n15064) );
  XOR U14769 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][23] ), .B(n15065), 
        .Z(n15062) );
  AND U14770 ( .A(n1274), .B(n15066), .Z(n15065) );
  XOR U14771 ( .A(n15067), .B(n15068), .Z(n15060) );
  AND U14772 ( .A(n1278), .B(n15059), .Z(n15068) );
  XNOR U14773 ( .A(n15069), .B(n15057), .Z(n15059) );
  XOR U14774 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n15070), .Z(n15057) );
  AND U14775 ( .A(n1290), .B(n15071), .Z(n15070) );
  IV U14776 ( .A(n15067), .Z(n15069) );
  XOR U14777 ( .A(n15072), .B(n15073), .Z(n15067) );
  AND U14778 ( .A(n1285), .B(n15066), .Z(n15073) );
  XOR U14779 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][23] ), .B(n15072), 
        .Z(n15066) );
  XOR U14780 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .B(n15074), 
        .Z(n15072) );
  AND U14781 ( .A(n1287), .B(n15071), .Z(n15074) );
  XOR U14782 ( .A(n15075), .B(n15076), .Z(n15071) );
  IV U14783 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .Z(n15076)
         );
  IV U14784 ( .A(\knn_comb_/min_val_out[0][23] ), .Z(n15075) );
  XOR U14785 ( .A(n93), .B(n15077), .Z(o[22]) );
  AND U14786 ( .A(n122), .B(n15078), .Z(n93) );
  XOR U14787 ( .A(n94), .B(n15077), .Z(n15078) );
  XOR U14788 ( .A(n15079), .B(n15080), .Z(n15077) );
  AND U14789 ( .A(n142), .B(n15081), .Z(n15080) );
  XOR U14790 ( .A(n15082), .B(n23), .Z(n94) );
  AND U14791 ( .A(n125), .B(n15083), .Z(n23) );
  XOR U14792 ( .A(n24), .B(n15082), .Z(n15083) );
  XOR U14793 ( .A(n15084), .B(n15085), .Z(n24) );
  AND U14794 ( .A(n130), .B(n15086), .Z(n15085) );
  XOR U14795 ( .A(p_input[22]), .B(n15084), .Z(n15086) );
  XNOR U14796 ( .A(n15087), .B(n15088), .Z(n15084) );
  AND U14797 ( .A(n134), .B(n15089), .Z(n15088) );
  XOR U14798 ( .A(n15090), .B(n15091), .Z(n15082) );
  AND U14799 ( .A(n138), .B(n15081), .Z(n15091) );
  XNOR U14800 ( .A(n15092), .B(n15079), .Z(n15081) );
  XOR U14801 ( .A(n15093), .B(n15094), .Z(n15079) );
  AND U14802 ( .A(n162), .B(n15095), .Z(n15094) );
  IV U14803 ( .A(n15090), .Z(n15092) );
  XOR U14804 ( .A(n15096), .B(n15097), .Z(n15090) );
  AND U14805 ( .A(n146), .B(n15089), .Z(n15097) );
  XNOR U14806 ( .A(n15087), .B(n15096), .Z(n15089) );
  XNOR U14807 ( .A(n15098), .B(n15099), .Z(n15087) );
  AND U14808 ( .A(n150), .B(n15100), .Z(n15099) );
  XOR U14809 ( .A(p_input[54]), .B(n15098), .Z(n15100) );
  XNOR U14810 ( .A(n15101), .B(n15102), .Z(n15098) );
  AND U14811 ( .A(n154), .B(n15103), .Z(n15102) );
  XOR U14812 ( .A(n15104), .B(n15105), .Z(n15096) );
  AND U14813 ( .A(n158), .B(n15095), .Z(n15105) );
  XNOR U14814 ( .A(n15106), .B(n15093), .Z(n15095) );
  XOR U14815 ( .A(n15107), .B(n15108), .Z(n15093) );
  AND U14816 ( .A(n181), .B(n15109), .Z(n15108) );
  IV U14817 ( .A(n15104), .Z(n15106) );
  XOR U14818 ( .A(n15110), .B(n15111), .Z(n15104) );
  AND U14819 ( .A(n165), .B(n15103), .Z(n15111) );
  XNOR U14820 ( .A(n15101), .B(n15110), .Z(n15103) );
  XNOR U14821 ( .A(n15112), .B(n15113), .Z(n15101) );
  AND U14822 ( .A(n169), .B(n15114), .Z(n15113) );
  XOR U14823 ( .A(p_input[86]), .B(n15112), .Z(n15114) );
  XNOR U14824 ( .A(n15115), .B(n15116), .Z(n15112) );
  AND U14825 ( .A(n173), .B(n15117), .Z(n15116) );
  XOR U14826 ( .A(n15118), .B(n15119), .Z(n15110) );
  AND U14827 ( .A(n177), .B(n15109), .Z(n15119) );
  XNOR U14828 ( .A(n15120), .B(n15107), .Z(n15109) );
  XOR U14829 ( .A(n15121), .B(n15122), .Z(n15107) );
  AND U14830 ( .A(n200), .B(n15123), .Z(n15122) );
  IV U14831 ( .A(n15118), .Z(n15120) );
  XOR U14832 ( .A(n15124), .B(n15125), .Z(n15118) );
  AND U14833 ( .A(n184), .B(n15117), .Z(n15125) );
  XNOR U14834 ( .A(n15115), .B(n15124), .Z(n15117) );
  XNOR U14835 ( .A(n15126), .B(n15127), .Z(n15115) );
  AND U14836 ( .A(n188), .B(n15128), .Z(n15127) );
  XOR U14837 ( .A(p_input[118]), .B(n15126), .Z(n15128) );
  XNOR U14838 ( .A(n15129), .B(n15130), .Z(n15126) );
  AND U14839 ( .A(n192), .B(n15131), .Z(n15130) );
  XOR U14840 ( .A(n15132), .B(n15133), .Z(n15124) );
  AND U14841 ( .A(n196), .B(n15123), .Z(n15133) );
  XNOR U14842 ( .A(n15134), .B(n15121), .Z(n15123) );
  XOR U14843 ( .A(n15135), .B(n15136), .Z(n15121) );
  AND U14844 ( .A(n219), .B(n15137), .Z(n15136) );
  IV U14845 ( .A(n15132), .Z(n15134) );
  XOR U14846 ( .A(n15138), .B(n15139), .Z(n15132) );
  AND U14847 ( .A(n203), .B(n15131), .Z(n15139) );
  XNOR U14848 ( .A(n15129), .B(n15138), .Z(n15131) );
  XNOR U14849 ( .A(n15140), .B(n15141), .Z(n15129) );
  AND U14850 ( .A(n207), .B(n15142), .Z(n15141) );
  XOR U14851 ( .A(p_input[150]), .B(n15140), .Z(n15142) );
  XNOR U14852 ( .A(n15143), .B(n15144), .Z(n15140) );
  AND U14853 ( .A(n211), .B(n15145), .Z(n15144) );
  XOR U14854 ( .A(n15146), .B(n15147), .Z(n15138) );
  AND U14855 ( .A(n215), .B(n15137), .Z(n15147) );
  XNOR U14856 ( .A(n15148), .B(n15135), .Z(n15137) );
  XOR U14857 ( .A(n15149), .B(n15150), .Z(n15135) );
  AND U14858 ( .A(n238), .B(n15151), .Z(n15150) );
  IV U14859 ( .A(n15146), .Z(n15148) );
  XOR U14860 ( .A(n15152), .B(n15153), .Z(n15146) );
  AND U14861 ( .A(n222), .B(n15145), .Z(n15153) );
  XNOR U14862 ( .A(n15143), .B(n15152), .Z(n15145) );
  XNOR U14863 ( .A(n15154), .B(n15155), .Z(n15143) );
  AND U14864 ( .A(n226), .B(n15156), .Z(n15155) );
  XOR U14865 ( .A(p_input[182]), .B(n15154), .Z(n15156) );
  XNOR U14866 ( .A(n15157), .B(n15158), .Z(n15154) );
  AND U14867 ( .A(n230), .B(n15159), .Z(n15158) );
  XOR U14868 ( .A(n15160), .B(n15161), .Z(n15152) );
  AND U14869 ( .A(n234), .B(n15151), .Z(n15161) );
  XNOR U14870 ( .A(n15162), .B(n15149), .Z(n15151) );
  XOR U14871 ( .A(n15163), .B(n15164), .Z(n15149) );
  AND U14872 ( .A(n257), .B(n15165), .Z(n15164) );
  IV U14873 ( .A(n15160), .Z(n15162) );
  XOR U14874 ( .A(n15166), .B(n15167), .Z(n15160) );
  AND U14875 ( .A(n241), .B(n15159), .Z(n15167) );
  XNOR U14876 ( .A(n15157), .B(n15166), .Z(n15159) );
  XNOR U14877 ( .A(n15168), .B(n15169), .Z(n15157) );
  AND U14878 ( .A(n245), .B(n15170), .Z(n15169) );
  XOR U14879 ( .A(p_input[214]), .B(n15168), .Z(n15170) );
  XNOR U14880 ( .A(n15171), .B(n15172), .Z(n15168) );
  AND U14881 ( .A(n249), .B(n15173), .Z(n15172) );
  XOR U14882 ( .A(n15174), .B(n15175), .Z(n15166) );
  AND U14883 ( .A(n253), .B(n15165), .Z(n15175) );
  XNOR U14884 ( .A(n15176), .B(n15163), .Z(n15165) );
  XOR U14885 ( .A(n15177), .B(n15178), .Z(n15163) );
  AND U14886 ( .A(n276), .B(n15179), .Z(n15178) );
  IV U14887 ( .A(n15174), .Z(n15176) );
  XOR U14888 ( .A(n15180), .B(n15181), .Z(n15174) );
  AND U14889 ( .A(n260), .B(n15173), .Z(n15181) );
  XNOR U14890 ( .A(n15171), .B(n15180), .Z(n15173) );
  XNOR U14891 ( .A(n15182), .B(n15183), .Z(n15171) );
  AND U14892 ( .A(n264), .B(n15184), .Z(n15183) );
  XOR U14893 ( .A(p_input[246]), .B(n15182), .Z(n15184) );
  XNOR U14894 ( .A(n15185), .B(n15186), .Z(n15182) );
  AND U14895 ( .A(n268), .B(n15187), .Z(n15186) );
  XOR U14896 ( .A(n15188), .B(n15189), .Z(n15180) );
  AND U14897 ( .A(n272), .B(n15179), .Z(n15189) );
  XNOR U14898 ( .A(n15190), .B(n15177), .Z(n15179) );
  XOR U14899 ( .A(n15191), .B(n15192), .Z(n15177) );
  AND U14900 ( .A(n295), .B(n15193), .Z(n15192) );
  IV U14901 ( .A(n15188), .Z(n15190) );
  XOR U14902 ( .A(n15194), .B(n15195), .Z(n15188) );
  AND U14903 ( .A(n279), .B(n15187), .Z(n15195) );
  XNOR U14904 ( .A(n15185), .B(n15194), .Z(n15187) );
  XNOR U14905 ( .A(n15196), .B(n15197), .Z(n15185) );
  AND U14906 ( .A(n283), .B(n15198), .Z(n15197) );
  XOR U14907 ( .A(p_input[278]), .B(n15196), .Z(n15198) );
  XNOR U14908 ( .A(n15199), .B(n15200), .Z(n15196) );
  AND U14909 ( .A(n287), .B(n15201), .Z(n15200) );
  XOR U14910 ( .A(n15202), .B(n15203), .Z(n15194) );
  AND U14911 ( .A(n291), .B(n15193), .Z(n15203) );
  XNOR U14912 ( .A(n15204), .B(n15191), .Z(n15193) );
  XOR U14913 ( .A(n15205), .B(n15206), .Z(n15191) );
  AND U14914 ( .A(n314), .B(n15207), .Z(n15206) );
  IV U14915 ( .A(n15202), .Z(n15204) );
  XOR U14916 ( .A(n15208), .B(n15209), .Z(n15202) );
  AND U14917 ( .A(n298), .B(n15201), .Z(n15209) );
  XNOR U14918 ( .A(n15199), .B(n15208), .Z(n15201) );
  XNOR U14919 ( .A(n15210), .B(n15211), .Z(n15199) );
  AND U14920 ( .A(n302), .B(n15212), .Z(n15211) );
  XOR U14921 ( .A(p_input[310]), .B(n15210), .Z(n15212) );
  XNOR U14922 ( .A(n15213), .B(n15214), .Z(n15210) );
  AND U14923 ( .A(n306), .B(n15215), .Z(n15214) );
  XOR U14924 ( .A(n15216), .B(n15217), .Z(n15208) );
  AND U14925 ( .A(n310), .B(n15207), .Z(n15217) );
  XNOR U14926 ( .A(n15218), .B(n15205), .Z(n15207) );
  XOR U14927 ( .A(n15219), .B(n15220), .Z(n15205) );
  AND U14928 ( .A(n333), .B(n15221), .Z(n15220) );
  IV U14929 ( .A(n15216), .Z(n15218) );
  XOR U14930 ( .A(n15222), .B(n15223), .Z(n15216) );
  AND U14931 ( .A(n317), .B(n15215), .Z(n15223) );
  XNOR U14932 ( .A(n15213), .B(n15222), .Z(n15215) );
  XNOR U14933 ( .A(n15224), .B(n15225), .Z(n15213) );
  AND U14934 ( .A(n321), .B(n15226), .Z(n15225) );
  XOR U14935 ( .A(p_input[342]), .B(n15224), .Z(n15226) );
  XNOR U14936 ( .A(n15227), .B(n15228), .Z(n15224) );
  AND U14937 ( .A(n325), .B(n15229), .Z(n15228) );
  XOR U14938 ( .A(n15230), .B(n15231), .Z(n15222) );
  AND U14939 ( .A(n329), .B(n15221), .Z(n15231) );
  XNOR U14940 ( .A(n15232), .B(n15219), .Z(n15221) );
  XOR U14941 ( .A(n15233), .B(n15234), .Z(n15219) );
  AND U14942 ( .A(n352), .B(n15235), .Z(n15234) );
  IV U14943 ( .A(n15230), .Z(n15232) );
  XOR U14944 ( .A(n15236), .B(n15237), .Z(n15230) );
  AND U14945 ( .A(n336), .B(n15229), .Z(n15237) );
  XNOR U14946 ( .A(n15227), .B(n15236), .Z(n15229) );
  XNOR U14947 ( .A(n15238), .B(n15239), .Z(n15227) );
  AND U14948 ( .A(n340), .B(n15240), .Z(n15239) );
  XOR U14949 ( .A(p_input[374]), .B(n15238), .Z(n15240) );
  XNOR U14950 ( .A(n15241), .B(n15242), .Z(n15238) );
  AND U14951 ( .A(n344), .B(n15243), .Z(n15242) );
  XOR U14952 ( .A(n15244), .B(n15245), .Z(n15236) );
  AND U14953 ( .A(n348), .B(n15235), .Z(n15245) );
  XNOR U14954 ( .A(n15246), .B(n15233), .Z(n15235) );
  XOR U14955 ( .A(n15247), .B(n15248), .Z(n15233) );
  AND U14956 ( .A(n371), .B(n15249), .Z(n15248) );
  IV U14957 ( .A(n15244), .Z(n15246) );
  XOR U14958 ( .A(n15250), .B(n15251), .Z(n15244) );
  AND U14959 ( .A(n355), .B(n15243), .Z(n15251) );
  XNOR U14960 ( .A(n15241), .B(n15250), .Z(n15243) );
  XNOR U14961 ( .A(n15252), .B(n15253), .Z(n15241) );
  AND U14962 ( .A(n359), .B(n15254), .Z(n15253) );
  XOR U14963 ( .A(p_input[406]), .B(n15252), .Z(n15254) );
  XNOR U14964 ( .A(n15255), .B(n15256), .Z(n15252) );
  AND U14965 ( .A(n363), .B(n15257), .Z(n15256) );
  XOR U14966 ( .A(n15258), .B(n15259), .Z(n15250) );
  AND U14967 ( .A(n367), .B(n15249), .Z(n15259) );
  XNOR U14968 ( .A(n15260), .B(n15247), .Z(n15249) );
  XOR U14969 ( .A(n15261), .B(n15262), .Z(n15247) );
  AND U14970 ( .A(n390), .B(n15263), .Z(n15262) );
  IV U14971 ( .A(n15258), .Z(n15260) );
  XOR U14972 ( .A(n15264), .B(n15265), .Z(n15258) );
  AND U14973 ( .A(n374), .B(n15257), .Z(n15265) );
  XNOR U14974 ( .A(n15255), .B(n15264), .Z(n15257) );
  XNOR U14975 ( .A(n15266), .B(n15267), .Z(n15255) );
  AND U14976 ( .A(n378), .B(n15268), .Z(n15267) );
  XOR U14977 ( .A(p_input[438]), .B(n15266), .Z(n15268) );
  XNOR U14978 ( .A(n15269), .B(n15270), .Z(n15266) );
  AND U14979 ( .A(n382), .B(n15271), .Z(n15270) );
  XOR U14980 ( .A(n15272), .B(n15273), .Z(n15264) );
  AND U14981 ( .A(n386), .B(n15263), .Z(n15273) );
  XNOR U14982 ( .A(n15274), .B(n15261), .Z(n15263) );
  XOR U14983 ( .A(n15275), .B(n15276), .Z(n15261) );
  AND U14984 ( .A(n409), .B(n15277), .Z(n15276) );
  IV U14985 ( .A(n15272), .Z(n15274) );
  XOR U14986 ( .A(n15278), .B(n15279), .Z(n15272) );
  AND U14987 ( .A(n393), .B(n15271), .Z(n15279) );
  XNOR U14988 ( .A(n15269), .B(n15278), .Z(n15271) );
  XNOR U14989 ( .A(n15280), .B(n15281), .Z(n15269) );
  AND U14990 ( .A(n397), .B(n15282), .Z(n15281) );
  XOR U14991 ( .A(p_input[470]), .B(n15280), .Z(n15282) );
  XNOR U14992 ( .A(n15283), .B(n15284), .Z(n15280) );
  AND U14993 ( .A(n401), .B(n15285), .Z(n15284) );
  XOR U14994 ( .A(n15286), .B(n15287), .Z(n15278) );
  AND U14995 ( .A(n405), .B(n15277), .Z(n15287) );
  XNOR U14996 ( .A(n15288), .B(n15275), .Z(n15277) );
  XOR U14997 ( .A(n15289), .B(n15290), .Z(n15275) );
  AND U14998 ( .A(n428), .B(n15291), .Z(n15290) );
  IV U14999 ( .A(n15286), .Z(n15288) );
  XOR U15000 ( .A(n15292), .B(n15293), .Z(n15286) );
  AND U15001 ( .A(n412), .B(n15285), .Z(n15293) );
  XNOR U15002 ( .A(n15283), .B(n15292), .Z(n15285) );
  XNOR U15003 ( .A(n15294), .B(n15295), .Z(n15283) );
  AND U15004 ( .A(n416), .B(n15296), .Z(n15295) );
  XOR U15005 ( .A(p_input[502]), .B(n15294), .Z(n15296) );
  XNOR U15006 ( .A(n15297), .B(n15298), .Z(n15294) );
  AND U15007 ( .A(n420), .B(n15299), .Z(n15298) );
  XOR U15008 ( .A(n15300), .B(n15301), .Z(n15292) );
  AND U15009 ( .A(n424), .B(n15291), .Z(n15301) );
  XNOR U15010 ( .A(n15302), .B(n15289), .Z(n15291) );
  XOR U15011 ( .A(n15303), .B(n15304), .Z(n15289) );
  AND U15012 ( .A(n447), .B(n15305), .Z(n15304) );
  IV U15013 ( .A(n15300), .Z(n15302) );
  XOR U15014 ( .A(n15306), .B(n15307), .Z(n15300) );
  AND U15015 ( .A(n431), .B(n15299), .Z(n15307) );
  XNOR U15016 ( .A(n15297), .B(n15306), .Z(n15299) );
  XNOR U15017 ( .A(n15308), .B(n15309), .Z(n15297) );
  AND U15018 ( .A(n435), .B(n15310), .Z(n15309) );
  XOR U15019 ( .A(p_input[534]), .B(n15308), .Z(n15310) );
  XNOR U15020 ( .A(n15311), .B(n15312), .Z(n15308) );
  AND U15021 ( .A(n439), .B(n15313), .Z(n15312) );
  XOR U15022 ( .A(n15314), .B(n15315), .Z(n15306) );
  AND U15023 ( .A(n443), .B(n15305), .Z(n15315) );
  XNOR U15024 ( .A(n15316), .B(n15303), .Z(n15305) );
  XOR U15025 ( .A(n15317), .B(n15318), .Z(n15303) );
  AND U15026 ( .A(n466), .B(n15319), .Z(n15318) );
  IV U15027 ( .A(n15314), .Z(n15316) );
  XOR U15028 ( .A(n15320), .B(n15321), .Z(n15314) );
  AND U15029 ( .A(n450), .B(n15313), .Z(n15321) );
  XNOR U15030 ( .A(n15311), .B(n15320), .Z(n15313) );
  XNOR U15031 ( .A(n15322), .B(n15323), .Z(n15311) );
  AND U15032 ( .A(n454), .B(n15324), .Z(n15323) );
  XOR U15033 ( .A(p_input[566]), .B(n15322), .Z(n15324) );
  XNOR U15034 ( .A(n15325), .B(n15326), .Z(n15322) );
  AND U15035 ( .A(n458), .B(n15327), .Z(n15326) );
  XOR U15036 ( .A(n15328), .B(n15329), .Z(n15320) );
  AND U15037 ( .A(n462), .B(n15319), .Z(n15329) );
  XNOR U15038 ( .A(n15330), .B(n15317), .Z(n15319) );
  XOR U15039 ( .A(n15331), .B(n15332), .Z(n15317) );
  AND U15040 ( .A(n485), .B(n15333), .Z(n15332) );
  IV U15041 ( .A(n15328), .Z(n15330) );
  XOR U15042 ( .A(n15334), .B(n15335), .Z(n15328) );
  AND U15043 ( .A(n469), .B(n15327), .Z(n15335) );
  XNOR U15044 ( .A(n15325), .B(n15334), .Z(n15327) );
  XNOR U15045 ( .A(n15336), .B(n15337), .Z(n15325) );
  AND U15046 ( .A(n473), .B(n15338), .Z(n15337) );
  XOR U15047 ( .A(p_input[598]), .B(n15336), .Z(n15338) );
  XNOR U15048 ( .A(n15339), .B(n15340), .Z(n15336) );
  AND U15049 ( .A(n477), .B(n15341), .Z(n15340) );
  XOR U15050 ( .A(n15342), .B(n15343), .Z(n15334) );
  AND U15051 ( .A(n481), .B(n15333), .Z(n15343) );
  XNOR U15052 ( .A(n15344), .B(n15331), .Z(n15333) );
  XOR U15053 ( .A(n15345), .B(n15346), .Z(n15331) );
  AND U15054 ( .A(n504), .B(n15347), .Z(n15346) );
  IV U15055 ( .A(n15342), .Z(n15344) );
  XOR U15056 ( .A(n15348), .B(n15349), .Z(n15342) );
  AND U15057 ( .A(n488), .B(n15341), .Z(n15349) );
  XNOR U15058 ( .A(n15339), .B(n15348), .Z(n15341) );
  XNOR U15059 ( .A(n15350), .B(n15351), .Z(n15339) );
  AND U15060 ( .A(n492), .B(n15352), .Z(n15351) );
  XOR U15061 ( .A(p_input[630]), .B(n15350), .Z(n15352) );
  XNOR U15062 ( .A(n15353), .B(n15354), .Z(n15350) );
  AND U15063 ( .A(n496), .B(n15355), .Z(n15354) );
  XOR U15064 ( .A(n15356), .B(n15357), .Z(n15348) );
  AND U15065 ( .A(n500), .B(n15347), .Z(n15357) );
  XNOR U15066 ( .A(n15358), .B(n15345), .Z(n15347) );
  XOR U15067 ( .A(n15359), .B(n15360), .Z(n15345) );
  AND U15068 ( .A(n523), .B(n15361), .Z(n15360) );
  IV U15069 ( .A(n15356), .Z(n15358) );
  XOR U15070 ( .A(n15362), .B(n15363), .Z(n15356) );
  AND U15071 ( .A(n507), .B(n15355), .Z(n15363) );
  XNOR U15072 ( .A(n15353), .B(n15362), .Z(n15355) );
  XNOR U15073 ( .A(n15364), .B(n15365), .Z(n15353) );
  AND U15074 ( .A(n511), .B(n15366), .Z(n15365) );
  XOR U15075 ( .A(p_input[662]), .B(n15364), .Z(n15366) );
  XNOR U15076 ( .A(n15367), .B(n15368), .Z(n15364) );
  AND U15077 ( .A(n515), .B(n15369), .Z(n15368) );
  XOR U15078 ( .A(n15370), .B(n15371), .Z(n15362) );
  AND U15079 ( .A(n519), .B(n15361), .Z(n15371) );
  XNOR U15080 ( .A(n15372), .B(n15359), .Z(n15361) );
  XOR U15081 ( .A(n15373), .B(n15374), .Z(n15359) );
  AND U15082 ( .A(n542), .B(n15375), .Z(n15374) );
  IV U15083 ( .A(n15370), .Z(n15372) );
  XOR U15084 ( .A(n15376), .B(n15377), .Z(n15370) );
  AND U15085 ( .A(n526), .B(n15369), .Z(n15377) );
  XNOR U15086 ( .A(n15367), .B(n15376), .Z(n15369) );
  XNOR U15087 ( .A(n15378), .B(n15379), .Z(n15367) );
  AND U15088 ( .A(n530), .B(n15380), .Z(n15379) );
  XOR U15089 ( .A(p_input[694]), .B(n15378), .Z(n15380) );
  XNOR U15090 ( .A(n15381), .B(n15382), .Z(n15378) );
  AND U15091 ( .A(n534), .B(n15383), .Z(n15382) );
  XOR U15092 ( .A(n15384), .B(n15385), .Z(n15376) );
  AND U15093 ( .A(n538), .B(n15375), .Z(n15385) );
  XNOR U15094 ( .A(n15386), .B(n15373), .Z(n15375) );
  XOR U15095 ( .A(n15387), .B(n15388), .Z(n15373) );
  AND U15096 ( .A(n561), .B(n15389), .Z(n15388) );
  IV U15097 ( .A(n15384), .Z(n15386) );
  XOR U15098 ( .A(n15390), .B(n15391), .Z(n15384) );
  AND U15099 ( .A(n545), .B(n15383), .Z(n15391) );
  XNOR U15100 ( .A(n15381), .B(n15390), .Z(n15383) );
  XNOR U15101 ( .A(n15392), .B(n15393), .Z(n15381) );
  AND U15102 ( .A(n549), .B(n15394), .Z(n15393) );
  XOR U15103 ( .A(p_input[726]), .B(n15392), .Z(n15394) );
  XNOR U15104 ( .A(n15395), .B(n15396), .Z(n15392) );
  AND U15105 ( .A(n553), .B(n15397), .Z(n15396) );
  XOR U15106 ( .A(n15398), .B(n15399), .Z(n15390) );
  AND U15107 ( .A(n557), .B(n15389), .Z(n15399) );
  XNOR U15108 ( .A(n15400), .B(n15387), .Z(n15389) );
  XOR U15109 ( .A(n15401), .B(n15402), .Z(n15387) );
  AND U15110 ( .A(n580), .B(n15403), .Z(n15402) );
  IV U15111 ( .A(n15398), .Z(n15400) );
  XOR U15112 ( .A(n15404), .B(n15405), .Z(n15398) );
  AND U15113 ( .A(n564), .B(n15397), .Z(n15405) );
  XNOR U15114 ( .A(n15395), .B(n15404), .Z(n15397) );
  XNOR U15115 ( .A(n15406), .B(n15407), .Z(n15395) );
  AND U15116 ( .A(n568), .B(n15408), .Z(n15407) );
  XOR U15117 ( .A(p_input[758]), .B(n15406), .Z(n15408) );
  XNOR U15118 ( .A(n15409), .B(n15410), .Z(n15406) );
  AND U15119 ( .A(n572), .B(n15411), .Z(n15410) );
  XOR U15120 ( .A(n15412), .B(n15413), .Z(n15404) );
  AND U15121 ( .A(n576), .B(n15403), .Z(n15413) );
  XNOR U15122 ( .A(n15414), .B(n15401), .Z(n15403) );
  XOR U15123 ( .A(n15415), .B(n15416), .Z(n15401) );
  AND U15124 ( .A(n599), .B(n15417), .Z(n15416) );
  IV U15125 ( .A(n15412), .Z(n15414) );
  XOR U15126 ( .A(n15418), .B(n15419), .Z(n15412) );
  AND U15127 ( .A(n583), .B(n15411), .Z(n15419) );
  XNOR U15128 ( .A(n15409), .B(n15418), .Z(n15411) );
  XNOR U15129 ( .A(n15420), .B(n15421), .Z(n15409) );
  AND U15130 ( .A(n587), .B(n15422), .Z(n15421) );
  XOR U15131 ( .A(p_input[790]), .B(n15420), .Z(n15422) );
  XNOR U15132 ( .A(n15423), .B(n15424), .Z(n15420) );
  AND U15133 ( .A(n591), .B(n15425), .Z(n15424) );
  XOR U15134 ( .A(n15426), .B(n15427), .Z(n15418) );
  AND U15135 ( .A(n595), .B(n15417), .Z(n15427) );
  XNOR U15136 ( .A(n15428), .B(n15415), .Z(n15417) );
  XOR U15137 ( .A(n15429), .B(n15430), .Z(n15415) );
  AND U15138 ( .A(n618), .B(n15431), .Z(n15430) );
  IV U15139 ( .A(n15426), .Z(n15428) );
  XOR U15140 ( .A(n15432), .B(n15433), .Z(n15426) );
  AND U15141 ( .A(n602), .B(n15425), .Z(n15433) );
  XNOR U15142 ( .A(n15423), .B(n15432), .Z(n15425) );
  XNOR U15143 ( .A(n15434), .B(n15435), .Z(n15423) );
  AND U15144 ( .A(n606), .B(n15436), .Z(n15435) );
  XOR U15145 ( .A(p_input[822]), .B(n15434), .Z(n15436) );
  XNOR U15146 ( .A(n15437), .B(n15438), .Z(n15434) );
  AND U15147 ( .A(n610), .B(n15439), .Z(n15438) );
  XOR U15148 ( .A(n15440), .B(n15441), .Z(n15432) );
  AND U15149 ( .A(n614), .B(n15431), .Z(n15441) );
  XNOR U15150 ( .A(n15442), .B(n15429), .Z(n15431) );
  XOR U15151 ( .A(n15443), .B(n15444), .Z(n15429) );
  AND U15152 ( .A(n637), .B(n15445), .Z(n15444) );
  IV U15153 ( .A(n15440), .Z(n15442) );
  XOR U15154 ( .A(n15446), .B(n15447), .Z(n15440) );
  AND U15155 ( .A(n621), .B(n15439), .Z(n15447) );
  XNOR U15156 ( .A(n15437), .B(n15446), .Z(n15439) );
  XNOR U15157 ( .A(n15448), .B(n15449), .Z(n15437) );
  AND U15158 ( .A(n625), .B(n15450), .Z(n15449) );
  XOR U15159 ( .A(p_input[854]), .B(n15448), .Z(n15450) );
  XNOR U15160 ( .A(n15451), .B(n15452), .Z(n15448) );
  AND U15161 ( .A(n629), .B(n15453), .Z(n15452) );
  XOR U15162 ( .A(n15454), .B(n15455), .Z(n15446) );
  AND U15163 ( .A(n633), .B(n15445), .Z(n15455) );
  XNOR U15164 ( .A(n15456), .B(n15443), .Z(n15445) );
  XOR U15165 ( .A(n15457), .B(n15458), .Z(n15443) );
  AND U15166 ( .A(n656), .B(n15459), .Z(n15458) );
  IV U15167 ( .A(n15454), .Z(n15456) );
  XOR U15168 ( .A(n15460), .B(n15461), .Z(n15454) );
  AND U15169 ( .A(n640), .B(n15453), .Z(n15461) );
  XNOR U15170 ( .A(n15451), .B(n15460), .Z(n15453) );
  XNOR U15171 ( .A(n15462), .B(n15463), .Z(n15451) );
  AND U15172 ( .A(n644), .B(n15464), .Z(n15463) );
  XOR U15173 ( .A(p_input[886]), .B(n15462), .Z(n15464) );
  XNOR U15174 ( .A(n15465), .B(n15466), .Z(n15462) );
  AND U15175 ( .A(n648), .B(n15467), .Z(n15466) );
  XOR U15176 ( .A(n15468), .B(n15469), .Z(n15460) );
  AND U15177 ( .A(n652), .B(n15459), .Z(n15469) );
  XNOR U15178 ( .A(n15470), .B(n15457), .Z(n15459) );
  XOR U15179 ( .A(n15471), .B(n15472), .Z(n15457) );
  AND U15180 ( .A(n675), .B(n15473), .Z(n15472) );
  IV U15181 ( .A(n15468), .Z(n15470) );
  XOR U15182 ( .A(n15474), .B(n15475), .Z(n15468) );
  AND U15183 ( .A(n659), .B(n15467), .Z(n15475) );
  XNOR U15184 ( .A(n15465), .B(n15474), .Z(n15467) );
  XNOR U15185 ( .A(n15476), .B(n15477), .Z(n15465) );
  AND U15186 ( .A(n663), .B(n15478), .Z(n15477) );
  XOR U15187 ( .A(p_input[918]), .B(n15476), .Z(n15478) );
  XNOR U15188 ( .A(n15479), .B(n15480), .Z(n15476) );
  AND U15189 ( .A(n667), .B(n15481), .Z(n15480) );
  XOR U15190 ( .A(n15482), .B(n15483), .Z(n15474) );
  AND U15191 ( .A(n671), .B(n15473), .Z(n15483) );
  XNOR U15192 ( .A(n15484), .B(n15471), .Z(n15473) );
  XOR U15193 ( .A(n15485), .B(n15486), .Z(n15471) );
  AND U15194 ( .A(n694), .B(n15487), .Z(n15486) );
  IV U15195 ( .A(n15482), .Z(n15484) );
  XOR U15196 ( .A(n15488), .B(n15489), .Z(n15482) );
  AND U15197 ( .A(n678), .B(n15481), .Z(n15489) );
  XNOR U15198 ( .A(n15479), .B(n15488), .Z(n15481) );
  XNOR U15199 ( .A(n15490), .B(n15491), .Z(n15479) );
  AND U15200 ( .A(n682), .B(n15492), .Z(n15491) );
  XOR U15201 ( .A(p_input[950]), .B(n15490), .Z(n15492) );
  XNOR U15202 ( .A(n15493), .B(n15494), .Z(n15490) );
  AND U15203 ( .A(n686), .B(n15495), .Z(n15494) );
  XOR U15204 ( .A(n15496), .B(n15497), .Z(n15488) );
  AND U15205 ( .A(n690), .B(n15487), .Z(n15497) );
  XNOR U15206 ( .A(n15498), .B(n15485), .Z(n15487) );
  XOR U15207 ( .A(n15499), .B(n15500), .Z(n15485) );
  AND U15208 ( .A(n713), .B(n15501), .Z(n15500) );
  IV U15209 ( .A(n15496), .Z(n15498) );
  XOR U15210 ( .A(n15502), .B(n15503), .Z(n15496) );
  AND U15211 ( .A(n697), .B(n15495), .Z(n15503) );
  XNOR U15212 ( .A(n15493), .B(n15502), .Z(n15495) );
  XNOR U15213 ( .A(n15504), .B(n15505), .Z(n15493) );
  AND U15214 ( .A(n701), .B(n15506), .Z(n15505) );
  XOR U15215 ( .A(p_input[982]), .B(n15504), .Z(n15506) );
  XNOR U15216 ( .A(n15507), .B(n15508), .Z(n15504) );
  AND U15217 ( .A(n705), .B(n15509), .Z(n15508) );
  XOR U15218 ( .A(n15510), .B(n15511), .Z(n15502) );
  AND U15219 ( .A(n709), .B(n15501), .Z(n15511) );
  XNOR U15220 ( .A(n15512), .B(n15499), .Z(n15501) );
  XOR U15221 ( .A(n15513), .B(n15514), .Z(n15499) );
  AND U15222 ( .A(n732), .B(n15515), .Z(n15514) );
  IV U15223 ( .A(n15510), .Z(n15512) );
  XOR U15224 ( .A(n15516), .B(n15517), .Z(n15510) );
  AND U15225 ( .A(n716), .B(n15509), .Z(n15517) );
  XNOR U15226 ( .A(n15507), .B(n15516), .Z(n15509) );
  XNOR U15227 ( .A(n15518), .B(n15519), .Z(n15507) );
  AND U15228 ( .A(n720), .B(n15520), .Z(n15519) );
  XOR U15229 ( .A(p_input[1014]), .B(n15518), .Z(n15520) );
  XNOR U15230 ( .A(n15521), .B(n15522), .Z(n15518) );
  AND U15231 ( .A(n724), .B(n15523), .Z(n15522) );
  XOR U15232 ( .A(n15524), .B(n15525), .Z(n15516) );
  AND U15233 ( .A(n728), .B(n15515), .Z(n15525) );
  XNOR U15234 ( .A(n15526), .B(n15513), .Z(n15515) );
  XOR U15235 ( .A(n15527), .B(n15528), .Z(n15513) );
  AND U15236 ( .A(n751), .B(n15529), .Z(n15528) );
  IV U15237 ( .A(n15524), .Z(n15526) );
  XOR U15238 ( .A(n15530), .B(n15531), .Z(n15524) );
  AND U15239 ( .A(n735), .B(n15523), .Z(n15531) );
  XNOR U15240 ( .A(n15521), .B(n15530), .Z(n15523) );
  XNOR U15241 ( .A(n15532), .B(n15533), .Z(n15521) );
  AND U15242 ( .A(n739), .B(n15534), .Z(n15533) );
  XOR U15243 ( .A(p_input[1046]), .B(n15532), .Z(n15534) );
  XNOR U15244 ( .A(n15535), .B(n15536), .Z(n15532) );
  AND U15245 ( .A(n743), .B(n15537), .Z(n15536) );
  XOR U15246 ( .A(n15538), .B(n15539), .Z(n15530) );
  AND U15247 ( .A(n747), .B(n15529), .Z(n15539) );
  XNOR U15248 ( .A(n15540), .B(n15527), .Z(n15529) );
  XOR U15249 ( .A(n15541), .B(n15542), .Z(n15527) );
  AND U15250 ( .A(n770), .B(n15543), .Z(n15542) );
  IV U15251 ( .A(n15538), .Z(n15540) );
  XOR U15252 ( .A(n15544), .B(n15545), .Z(n15538) );
  AND U15253 ( .A(n754), .B(n15537), .Z(n15545) );
  XNOR U15254 ( .A(n15535), .B(n15544), .Z(n15537) );
  XNOR U15255 ( .A(n15546), .B(n15547), .Z(n15535) );
  AND U15256 ( .A(n758), .B(n15548), .Z(n15547) );
  XOR U15257 ( .A(p_input[1078]), .B(n15546), .Z(n15548) );
  XNOR U15258 ( .A(n15549), .B(n15550), .Z(n15546) );
  AND U15259 ( .A(n762), .B(n15551), .Z(n15550) );
  XOR U15260 ( .A(n15552), .B(n15553), .Z(n15544) );
  AND U15261 ( .A(n766), .B(n15543), .Z(n15553) );
  XNOR U15262 ( .A(n15554), .B(n15541), .Z(n15543) );
  XOR U15263 ( .A(n15555), .B(n15556), .Z(n15541) );
  AND U15264 ( .A(n789), .B(n15557), .Z(n15556) );
  IV U15265 ( .A(n15552), .Z(n15554) );
  XOR U15266 ( .A(n15558), .B(n15559), .Z(n15552) );
  AND U15267 ( .A(n773), .B(n15551), .Z(n15559) );
  XNOR U15268 ( .A(n15549), .B(n15558), .Z(n15551) );
  XNOR U15269 ( .A(n15560), .B(n15561), .Z(n15549) );
  AND U15270 ( .A(n777), .B(n15562), .Z(n15561) );
  XOR U15271 ( .A(p_input[1110]), .B(n15560), .Z(n15562) );
  XNOR U15272 ( .A(n15563), .B(n15564), .Z(n15560) );
  AND U15273 ( .A(n781), .B(n15565), .Z(n15564) );
  XOR U15274 ( .A(n15566), .B(n15567), .Z(n15558) );
  AND U15275 ( .A(n785), .B(n15557), .Z(n15567) );
  XNOR U15276 ( .A(n15568), .B(n15555), .Z(n15557) );
  XOR U15277 ( .A(n15569), .B(n15570), .Z(n15555) );
  AND U15278 ( .A(n808), .B(n15571), .Z(n15570) );
  IV U15279 ( .A(n15566), .Z(n15568) );
  XOR U15280 ( .A(n15572), .B(n15573), .Z(n15566) );
  AND U15281 ( .A(n792), .B(n15565), .Z(n15573) );
  XNOR U15282 ( .A(n15563), .B(n15572), .Z(n15565) );
  XNOR U15283 ( .A(n15574), .B(n15575), .Z(n15563) );
  AND U15284 ( .A(n796), .B(n15576), .Z(n15575) );
  XOR U15285 ( .A(p_input[1142]), .B(n15574), .Z(n15576) );
  XNOR U15286 ( .A(n15577), .B(n15578), .Z(n15574) );
  AND U15287 ( .A(n800), .B(n15579), .Z(n15578) );
  XOR U15288 ( .A(n15580), .B(n15581), .Z(n15572) );
  AND U15289 ( .A(n804), .B(n15571), .Z(n15581) );
  XNOR U15290 ( .A(n15582), .B(n15569), .Z(n15571) );
  XOR U15291 ( .A(n15583), .B(n15584), .Z(n15569) );
  AND U15292 ( .A(n827), .B(n15585), .Z(n15584) );
  IV U15293 ( .A(n15580), .Z(n15582) );
  XOR U15294 ( .A(n15586), .B(n15587), .Z(n15580) );
  AND U15295 ( .A(n811), .B(n15579), .Z(n15587) );
  XNOR U15296 ( .A(n15577), .B(n15586), .Z(n15579) );
  XNOR U15297 ( .A(n15588), .B(n15589), .Z(n15577) );
  AND U15298 ( .A(n815), .B(n15590), .Z(n15589) );
  XOR U15299 ( .A(p_input[1174]), .B(n15588), .Z(n15590) );
  XNOR U15300 ( .A(n15591), .B(n15592), .Z(n15588) );
  AND U15301 ( .A(n819), .B(n15593), .Z(n15592) );
  XOR U15302 ( .A(n15594), .B(n15595), .Z(n15586) );
  AND U15303 ( .A(n823), .B(n15585), .Z(n15595) );
  XNOR U15304 ( .A(n15596), .B(n15583), .Z(n15585) );
  XOR U15305 ( .A(n15597), .B(n15598), .Z(n15583) );
  AND U15306 ( .A(n846), .B(n15599), .Z(n15598) );
  IV U15307 ( .A(n15594), .Z(n15596) );
  XOR U15308 ( .A(n15600), .B(n15601), .Z(n15594) );
  AND U15309 ( .A(n830), .B(n15593), .Z(n15601) );
  XNOR U15310 ( .A(n15591), .B(n15600), .Z(n15593) );
  XNOR U15311 ( .A(n15602), .B(n15603), .Z(n15591) );
  AND U15312 ( .A(n834), .B(n15604), .Z(n15603) );
  XOR U15313 ( .A(p_input[1206]), .B(n15602), .Z(n15604) );
  XNOR U15314 ( .A(n15605), .B(n15606), .Z(n15602) );
  AND U15315 ( .A(n838), .B(n15607), .Z(n15606) );
  XOR U15316 ( .A(n15608), .B(n15609), .Z(n15600) );
  AND U15317 ( .A(n842), .B(n15599), .Z(n15609) );
  XNOR U15318 ( .A(n15610), .B(n15597), .Z(n15599) );
  XOR U15319 ( .A(n15611), .B(n15612), .Z(n15597) );
  AND U15320 ( .A(n865), .B(n15613), .Z(n15612) );
  IV U15321 ( .A(n15608), .Z(n15610) );
  XOR U15322 ( .A(n15614), .B(n15615), .Z(n15608) );
  AND U15323 ( .A(n849), .B(n15607), .Z(n15615) );
  XNOR U15324 ( .A(n15605), .B(n15614), .Z(n15607) );
  XNOR U15325 ( .A(n15616), .B(n15617), .Z(n15605) );
  AND U15326 ( .A(n853), .B(n15618), .Z(n15617) );
  XOR U15327 ( .A(p_input[1238]), .B(n15616), .Z(n15618) );
  XNOR U15328 ( .A(n15619), .B(n15620), .Z(n15616) );
  AND U15329 ( .A(n857), .B(n15621), .Z(n15620) );
  XOR U15330 ( .A(n15622), .B(n15623), .Z(n15614) );
  AND U15331 ( .A(n861), .B(n15613), .Z(n15623) );
  XNOR U15332 ( .A(n15624), .B(n15611), .Z(n15613) );
  XOR U15333 ( .A(n15625), .B(n15626), .Z(n15611) );
  AND U15334 ( .A(n884), .B(n15627), .Z(n15626) );
  IV U15335 ( .A(n15622), .Z(n15624) );
  XOR U15336 ( .A(n15628), .B(n15629), .Z(n15622) );
  AND U15337 ( .A(n868), .B(n15621), .Z(n15629) );
  XNOR U15338 ( .A(n15619), .B(n15628), .Z(n15621) );
  XNOR U15339 ( .A(n15630), .B(n15631), .Z(n15619) );
  AND U15340 ( .A(n872), .B(n15632), .Z(n15631) );
  XOR U15341 ( .A(p_input[1270]), .B(n15630), .Z(n15632) );
  XNOR U15342 ( .A(n15633), .B(n15634), .Z(n15630) );
  AND U15343 ( .A(n876), .B(n15635), .Z(n15634) );
  XOR U15344 ( .A(n15636), .B(n15637), .Z(n15628) );
  AND U15345 ( .A(n880), .B(n15627), .Z(n15637) );
  XNOR U15346 ( .A(n15638), .B(n15625), .Z(n15627) );
  XOR U15347 ( .A(n15639), .B(n15640), .Z(n15625) );
  AND U15348 ( .A(n903), .B(n15641), .Z(n15640) );
  IV U15349 ( .A(n15636), .Z(n15638) );
  XOR U15350 ( .A(n15642), .B(n15643), .Z(n15636) );
  AND U15351 ( .A(n887), .B(n15635), .Z(n15643) );
  XNOR U15352 ( .A(n15633), .B(n15642), .Z(n15635) );
  XNOR U15353 ( .A(n15644), .B(n15645), .Z(n15633) );
  AND U15354 ( .A(n891), .B(n15646), .Z(n15645) );
  XOR U15355 ( .A(p_input[1302]), .B(n15644), .Z(n15646) );
  XNOR U15356 ( .A(n15647), .B(n15648), .Z(n15644) );
  AND U15357 ( .A(n895), .B(n15649), .Z(n15648) );
  XOR U15358 ( .A(n15650), .B(n15651), .Z(n15642) );
  AND U15359 ( .A(n899), .B(n15641), .Z(n15651) );
  XNOR U15360 ( .A(n15652), .B(n15639), .Z(n15641) );
  XOR U15361 ( .A(n15653), .B(n15654), .Z(n15639) );
  AND U15362 ( .A(n922), .B(n15655), .Z(n15654) );
  IV U15363 ( .A(n15650), .Z(n15652) );
  XOR U15364 ( .A(n15656), .B(n15657), .Z(n15650) );
  AND U15365 ( .A(n906), .B(n15649), .Z(n15657) );
  XNOR U15366 ( .A(n15647), .B(n15656), .Z(n15649) );
  XNOR U15367 ( .A(n15658), .B(n15659), .Z(n15647) );
  AND U15368 ( .A(n910), .B(n15660), .Z(n15659) );
  XOR U15369 ( .A(p_input[1334]), .B(n15658), .Z(n15660) );
  XNOR U15370 ( .A(n15661), .B(n15662), .Z(n15658) );
  AND U15371 ( .A(n914), .B(n15663), .Z(n15662) );
  XOR U15372 ( .A(n15664), .B(n15665), .Z(n15656) );
  AND U15373 ( .A(n918), .B(n15655), .Z(n15665) );
  XNOR U15374 ( .A(n15666), .B(n15653), .Z(n15655) );
  XOR U15375 ( .A(n15667), .B(n15668), .Z(n15653) );
  AND U15376 ( .A(n941), .B(n15669), .Z(n15668) );
  IV U15377 ( .A(n15664), .Z(n15666) );
  XOR U15378 ( .A(n15670), .B(n15671), .Z(n15664) );
  AND U15379 ( .A(n925), .B(n15663), .Z(n15671) );
  XNOR U15380 ( .A(n15661), .B(n15670), .Z(n15663) );
  XNOR U15381 ( .A(n15672), .B(n15673), .Z(n15661) );
  AND U15382 ( .A(n929), .B(n15674), .Z(n15673) );
  XOR U15383 ( .A(p_input[1366]), .B(n15672), .Z(n15674) );
  XNOR U15384 ( .A(n15675), .B(n15676), .Z(n15672) );
  AND U15385 ( .A(n933), .B(n15677), .Z(n15676) );
  XOR U15386 ( .A(n15678), .B(n15679), .Z(n15670) );
  AND U15387 ( .A(n937), .B(n15669), .Z(n15679) );
  XNOR U15388 ( .A(n15680), .B(n15667), .Z(n15669) );
  XOR U15389 ( .A(n15681), .B(n15682), .Z(n15667) );
  AND U15390 ( .A(n960), .B(n15683), .Z(n15682) );
  IV U15391 ( .A(n15678), .Z(n15680) );
  XOR U15392 ( .A(n15684), .B(n15685), .Z(n15678) );
  AND U15393 ( .A(n944), .B(n15677), .Z(n15685) );
  XNOR U15394 ( .A(n15675), .B(n15684), .Z(n15677) );
  XNOR U15395 ( .A(n15686), .B(n15687), .Z(n15675) );
  AND U15396 ( .A(n948), .B(n15688), .Z(n15687) );
  XOR U15397 ( .A(p_input[1398]), .B(n15686), .Z(n15688) );
  XNOR U15398 ( .A(n15689), .B(n15690), .Z(n15686) );
  AND U15399 ( .A(n952), .B(n15691), .Z(n15690) );
  XOR U15400 ( .A(n15692), .B(n15693), .Z(n15684) );
  AND U15401 ( .A(n956), .B(n15683), .Z(n15693) );
  XNOR U15402 ( .A(n15694), .B(n15681), .Z(n15683) );
  XOR U15403 ( .A(n15695), .B(n15696), .Z(n15681) );
  AND U15404 ( .A(n979), .B(n15697), .Z(n15696) );
  IV U15405 ( .A(n15692), .Z(n15694) );
  XOR U15406 ( .A(n15698), .B(n15699), .Z(n15692) );
  AND U15407 ( .A(n963), .B(n15691), .Z(n15699) );
  XNOR U15408 ( .A(n15689), .B(n15698), .Z(n15691) );
  XNOR U15409 ( .A(n15700), .B(n15701), .Z(n15689) );
  AND U15410 ( .A(n967), .B(n15702), .Z(n15701) );
  XOR U15411 ( .A(p_input[1430]), .B(n15700), .Z(n15702) );
  XNOR U15412 ( .A(n15703), .B(n15704), .Z(n15700) );
  AND U15413 ( .A(n971), .B(n15705), .Z(n15704) );
  XOR U15414 ( .A(n15706), .B(n15707), .Z(n15698) );
  AND U15415 ( .A(n975), .B(n15697), .Z(n15707) );
  XNOR U15416 ( .A(n15708), .B(n15695), .Z(n15697) );
  XOR U15417 ( .A(n15709), .B(n15710), .Z(n15695) );
  AND U15418 ( .A(n998), .B(n15711), .Z(n15710) );
  IV U15419 ( .A(n15706), .Z(n15708) );
  XOR U15420 ( .A(n15712), .B(n15713), .Z(n15706) );
  AND U15421 ( .A(n982), .B(n15705), .Z(n15713) );
  XNOR U15422 ( .A(n15703), .B(n15712), .Z(n15705) );
  XNOR U15423 ( .A(n15714), .B(n15715), .Z(n15703) );
  AND U15424 ( .A(n986), .B(n15716), .Z(n15715) );
  XOR U15425 ( .A(p_input[1462]), .B(n15714), .Z(n15716) );
  XNOR U15426 ( .A(n15717), .B(n15718), .Z(n15714) );
  AND U15427 ( .A(n990), .B(n15719), .Z(n15718) );
  XOR U15428 ( .A(n15720), .B(n15721), .Z(n15712) );
  AND U15429 ( .A(n994), .B(n15711), .Z(n15721) );
  XNOR U15430 ( .A(n15722), .B(n15709), .Z(n15711) );
  XOR U15431 ( .A(n15723), .B(n15724), .Z(n15709) );
  AND U15432 ( .A(n1017), .B(n15725), .Z(n15724) );
  IV U15433 ( .A(n15720), .Z(n15722) );
  XOR U15434 ( .A(n15726), .B(n15727), .Z(n15720) );
  AND U15435 ( .A(n1001), .B(n15719), .Z(n15727) );
  XNOR U15436 ( .A(n15717), .B(n15726), .Z(n15719) );
  XNOR U15437 ( .A(n15728), .B(n15729), .Z(n15717) );
  AND U15438 ( .A(n1005), .B(n15730), .Z(n15729) );
  XOR U15439 ( .A(p_input[1494]), .B(n15728), .Z(n15730) );
  XNOR U15440 ( .A(n15731), .B(n15732), .Z(n15728) );
  AND U15441 ( .A(n1009), .B(n15733), .Z(n15732) );
  XOR U15442 ( .A(n15734), .B(n15735), .Z(n15726) );
  AND U15443 ( .A(n1013), .B(n15725), .Z(n15735) );
  XNOR U15444 ( .A(n15736), .B(n15723), .Z(n15725) );
  XOR U15445 ( .A(n15737), .B(n15738), .Z(n15723) );
  AND U15446 ( .A(n1036), .B(n15739), .Z(n15738) );
  IV U15447 ( .A(n15734), .Z(n15736) );
  XOR U15448 ( .A(n15740), .B(n15741), .Z(n15734) );
  AND U15449 ( .A(n1020), .B(n15733), .Z(n15741) );
  XNOR U15450 ( .A(n15731), .B(n15740), .Z(n15733) );
  XNOR U15451 ( .A(n15742), .B(n15743), .Z(n15731) );
  AND U15452 ( .A(n1024), .B(n15744), .Z(n15743) );
  XOR U15453 ( .A(p_input[1526]), .B(n15742), .Z(n15744) );
  XNOR U15454 ( .A(n15745), .B(n15746), .Z(n15742) );
  AND U15455 ( .A(n1028), .B(n15747), .Z(n15746) );
  XOR U15456 ( .A(n15748), .B(n15749), .Z(n15740) );
  AND U15457 ( .A(n1032), .B(n15739), .Z(n15749) );
  XNOR U15458 ( .A(n15750), .B(n15737), .Z(n15739) );
  XOR U15459 ( .A(n15751), .B(n15752), .Z(n15737) );
  AND U15460 ( .A(n1055), .B(n15753), .Z(n15752) );
  IV U15461 ( .A(n15748), .Z(n15750) );
  XOR U15462 ( .A(n15754), .B(n15755), .Z(n15748) );
  AND U15463 ( .A(n1039), .B(n15747), .Z(n15755) );
  XNOR U15464 ( .A(n15745), .B(n15754), .Z(n15747) );
  XNOR U15465 ( .A(n15756), .B(n15757), .Z(n15745) );
  AND U15466 ( .A(n1043), .B(n15758), .Z(n15757) );
  XOR U15467 ( .A(p_input[1558]), .B(n15756), .Z(n15758) );
  XNOR U15468 ( .A(n15759), .B(n15760), .Z(n15756) );
  AND U15469 ( .A(n1047), .B(n15761), .Z(n15760) );
  XOR U15470 ( .A(n15762), .B(n15763), .Z(n15754) );
  AND U15471 ( .A(n1051), .B(n15753), .Z(n15763) );
  XNOR U15472 ( .A(n15764), .B(n15751), .Z(n15753) );
  XOR U15473 ( .A(n15765), .B(n15766), .Z(n15751) );
  AND U15474 ( .A(n1074), .B(n15767), .Z(n15766) );
  IV U15475 ( .A(n15762), .Z(n15764) );
  XOR U15476 ( .A(n15768), .B(n15769), .Z(n15762) );
  AND U15477 ( .A(n1058), .B(n15761), .Z(n15769) );
  XNOR U15478 ( .A(n15759), .B(n15768), .Z(n15761) );
  XNOR U15479 ( .A(n15770), .B(n15771), .Z(n15759) );
  AND U15480 ( .A(n1062), .B(n15772), .Z(n15771) );
  XOR U15481 ( .A(p_input[1590]), .B(n15770), .Z(n15772) );
  XNOR U15482 ( .A(n15773), .B(n15774), .Z(n15770) );
  AND U15483 ( .A(n1066), .B(n15775), .Z(n15774) );
  XOR U15484 ( .A(n15776), .B(n15777), .Z(n15768) );
  AND U15485 ( .A(n1070), .B(n15767), .Z(n15777) );
  XNOR U15486 ( .A(n15778), .B(n15765), .Z(n15767) );
  XOR U15487 ( .A(n15779), .B(n15780), .Z(n15765) );
  AND U15488 ( .A(n1093), .B(n15781), .Z(n15780) );
  IV U15489 ( .A(n15776), .Z(n15778) );
  XOR U15490 ( .A(n15782), .B(n15783), .Z(n15776) );
  AND U15491 ( .A(n1077), .B(n15775), .Z(n15783) );
  XNOR U15492 ( .A(n15773), .B(n15782), .Z(n15775) );
  XNOR U15493 ( .A(n15784), .B(n15785), .Z(n15773) );
  AND U15494 ( .A(n1081), .B(n15786), .Z(n15785) );
  XOR U15495 ( .A(p_input[1622]), .B(n15784), .Z(n15786) );
  XNOR U15496 ( .A(n15787), .B(n15788), .Z(n15784) );
  AND U15497 ( .A(n1085), .B(n15789), .Z(n15788) );
  XOR U15498 ( .A(n15790), .B(n15791), .Z(n15782) );
  AND U15499 ( .A(n1089), .B(n15781), .Z(n15791) );
  XNOR U15500 ( .A(n15792), .B(n15779), .Z(n15781) );
  XOR U15501 ( .A(n15793), .B(n15794), .Z(n15779) );
  AND U15502 ( .A(n1112), .B(n15795), .Z(n15794) );
  IV U15503 ( .A(n15790), .Z(n15792) );
  XOR U15504 ( .A(n15796), .B(n15797), .Z(n15790) );
  AND U15505 ( .A(n1096), .B(n15789), .Z(n15797) );
  XNOR U15506 ( .A(n15787), .B(n15796), .Z(n15789) );
  XNOR U15507 ( .A(n15798), .B(n15799), .Z(n15787) );
  AND U15508 ( .A(n1100), .B(n15800), .Z(n15799) );
  XOR U15509 ( .A(p_input[1654]), .B(n15798), .Z(n15800) );
  XNOR U15510 ( .A(n15801), .B(n15802), .Z(n15798) );
  AND U15511 ( .A(n1104), .B(n15803), .Z(n15802) );
  XOR U15512 ( .A(n15804), .B(n15805), .Z(n15796) );
  AND U15513 ( .A(n1108), .B(n15795), .Z(n15805) );
  XNOR U15514 ( .A(n15806), .B(n15793), .Z(n15795) );
  XOR U15515 ( .A(n15807), .B(n15808), .Z(n15793) );
  AND U15516 ( .A(n1131), .B(n15809), .Z(n15808) );
  IV U15517 ( .A(n15804), .Z(n15806) );
  XOR U15518 ( .A(n15810), .B(n15811), .Z(n15804) );
  AND U15519 ( .A(n1115), .B(n15803), .Z(n15811) );
  XNOR U15520 ( .A(n15801), .B(n15810), .Z(n15803) );
  XNOR U15521 ( .A(n15812), .B(n15813), .Z(n15801) );
  AND U15522 ( .A(n1119), .B(n15814), .Z(n15813) );
  XOR U15523 ( .A(p_input[1686]), .B(n15812), .Z(n15814) );
  XNOR U15524 ( .A(n15815), .B(n15816), .Z(n15812) );
  AND U15525 ( .A(n1123), .B(n15817), .Z(n15816) );
  XOR U15526 ( .A(n15818), .B(n15819), .Z(n15810) );
  AND U15527 ( .A(n1127), .B(n15809), .Z(n15819) );
  XNOR U15528 ( .A(n15820), .B(n15807), .Z(n15809) );
  XOR U15529 ( .A(n15821), .B(n15822), .Z(n15807) );
  AND U15530 ( .A(n1150), .B(n15823), .Z(n15822) );
  IV U15531 ( .A(n15818), .Z(n15820) );
  XOR U15532 ( .A(n15824), .B(n15825), .Z(n15818) );
  AND U15533 ( .A(n1134), .B(n15817), .Z(n15825) );
  XNOR U15534 ( .A(n15815), .B(n15824), .Z(n15817) );
  XNOR U15535 ( .A(n15826), .B(n15827), .Z(n15815) );
  AND U15536 ( .A(n1138), .B(n15828), .Z(n15827) );
  XOR U15537 ( .A(p_input[1718]), .B(n15826), .Z(n15828) );
  XNOR U15538 ( .A(n15829), .B(n15830), .Z(n15826) );
  AND U15539 ( .A(n1142), .B(n15831), .Z(n15830) );
  XOR U15540 ( .A(n15832), .B(n15833), .Z(n15824) );
  AND U15541 ( .A(n1146), .B(n15823), .Z(n15833) );
  XNOR U15542 ( .A(n15834), .B(n15821), .Z(n15823) );
  XOR U15543 ( .A(n15835), .B(n15836), .Z(n15821) );
  AND U15544 ( .A(n1169), .B(n15837), .Z(n15836) );
  IV U15545 ( .A(n15832), .Z(n15834) );
  XOR U15546 ( .A(n15838), .B(n15839), .Z(n15832) );
  AND U15547 ( .A(n1153), .B(n15831), .Z(n15839) );
  XNOR U15548 ( .A(n15829), .B(n15838), .Z(n15831) );
  XNOR U15549 ( .A(n15840), .B(n15841), .Z(n15829) );
  AND U15550 ( .A(n1157), .B(n15842), .Z(n15841) );
  XOR U15551 ( .A(p_input[1750]), .B(n15840), .Z(n15842) );
  XNOR U15552 ( .A(n15843), .B(n15844), .Z(n15840) );
  AND U15553 ( .A(n1161), .B(n15845), .Z(n15844) );
  XOR U15554 ( .A(n15846), .B(n15847), .Z(n15838) );
  AND U15555 ( .A(n1165), .B(n15837), .Z(n15847) );
  XNOR U15556 ( .A(n15848), .B(n15835), .Z(n15837) );
  XOR U15557 ( .A(n15849), .B(n15850), .Z(n15835) );
  AND U15558 ( .A(n1188), .B(n15851), .Z(n15850) );
  IV U15559 ( .A(n15846), .Z(n15848) );
  XOR U15560 ( .A(n15852), .B(n15853), .Z(n15846) );
  AND U15561 ( .A(n1172), .B(n15845), .Z(n15853) );
  XNOR U15562 ( .A(n15843), .B(n15852), .Z(n15845) );
  XNOR U15563 ( .A(n15854), .B(n15855), .Z(n15843) );
  AND U15564 ( .A(n1176), .B(n15856), .Z(n15855) );
  XOR U15565 ( .A(p_input[1782]), .B(n15854), .Z(n15856) );
  XNOR U15566 ( .A(n15857), .B(n15858), .Z(n15854) );
  AND U15567 ( .A(n1180), .B(n15859), .Z(n15858) );
  XOR U15568 ( .A(n15860), .B(n15861), .Z(n15852) );
  AND U15569 ( .A(n1184), .B(n15851), .Z(n15861) );
  XNOR U15570 ( .A(n15862), .B(n15849), .Z(n15851) );
  XOR U15571 ( .A(n15863), .B(n15864), .Z(n15849) );
  AND U15572 ( .A(n1207), .B(n15865), .Z(n15864) );
  IV U15573 ( .A(n15860), .Z(n15862) );
  XOR U15574 ( .A(n15866), .B(n15867), .Z(n15860) );
  AND U15575 ( .A(n1191), .B(n15859), .Z(n15867) );
  XNOR U15576 ( .A(n15857), .B(n15866), .Z(n15859) );
  XNOR U15577 ( .A(n15868), .B(n15869), .Z(n15857) );
  AND U15578 ( .A(n1195), .B(n15870), .Z(n15869) );
  XOR U15579 ( .A(p_input[1814]), .B(n15868), .Z(n15870) );
  XNOR U15580 ( .A(n15871), .B(n15872), .Z(n15868) );
  AND U15581 ( .A(n1199), .B(n15873), .Z(n15872) );
  XOR U15582 ( .A(n15874), .B(n15875), .Z(n15866) );
  AND U15583 ( .A(n1203), .B(n15865), .Z(n15875) );
  XNOR U15584 ( .A(n15876), .B(n15863), .Z(n15865) );
  XOR U15585 ( .A(n15877), .B(n15878), .Z(n15863) );
  AND U15586 ( .A(n1226), .B(n15879), .Z(n15878) );
  IV U15587 ( .A(n15874), .Z(n15876) );
  XOR U15588 ( .A(n15880), .B(n15881), .Z(n15874) );
  AND U15589 ( .A(n1210), .B(n15873), .Z(n15881) );
  XNOR U15590 ( .A(n15871), .B(n15880), .Z(n15873) );
  XNOR U15591 ( .A(n15882), .B(n15883), .Z(n15871) );
  AND U15592 ( .A(n1214), .B(n15884), .Z(n15883) );
  XOR U15593 ( .A(p_input[1846]), .B(n15882), .Z(n15884) );
  XNOR U15594 ( .A(n15885), .B(n15886), .Z(n15882) );
  AND U15595 ( .A(n1218), .B(n15887), .Z(n15886) );
  XOR U15596 ( .A(n15888), .B(n15889), .Z(n15880) );
  AND U15597 ( .A(n1222), .B(n15879), .Z(n15889) );
  XNOR U15598 ( .A(n15890), .B(n15877), .Z(n15879) );
  XOR U15599 ( .A(n15891), .B(n15892), .Z(n15877) );
  AND U15600 ( .A(n1245), .B(n15893), .Z(n15892) );
  IV U15601 ( .A(n15888), .Z(n15890) );
  XOR U15602 ( .A(n15894), .B(n15895), .Z(n15888) );
  AND U15603 ( .A(n1229), .B(n15887), .Z(n15895) );
  XNOR U15604 ( .A(n15885), .B(n15894), .Z(n15887) );
  XNOR U15605 ( .A(n15896), .B(n15897), .Z(n15885) );
  AND U15606 ( .A(n1233), .B(n15898), .Z(n15897) );
  XOR U15607 ( .A(p_input[1878]), .B(n15896), .Z(n15898) );
  XNOR U15608 ( .A(n15899), .B(n15900), .Z(n15896) );
  AND U15609 ( .A(n1237), .B(n15901), .Z(n15900) );
  XOR U15610 ( .A(n15902), .B(n15903), .Z(n15894) );
  AND U15611 ( .A(n1241), .B(n15893), .Z(n15903) );
  XNOR U15612 ( .A(n15904), .B(n15891), .Z(n15893) );
  XOR U15613 ( .A(n15905), .B(n15906), .Z(n15891) );
  AND U15614 ( .A(n1264), .B(n15907), .Z(n15906) );
  IV U15615 ( .A(n15902), .Z(n15904) );
  XOR U15616 ( .A(n15908), .B(n15909), .Z(n15902) );
  AND U15617 ( .A(n1248), .B(n15901), .Z(n15909) );
  XNOR U15618 ( .A(n15899), .B(n15908), .Z(n15901) );
  XNOR U15619 ( .A(n15910), .B(n15911), .Z(n15899) );
  AND U15620 ( .A(n1252), .B(n15912), .Z(n15911) );
  XOR U15621 ( .A(p_input[1910]), .B(n15910), .Z(n15912) );
  XNOR U15622 ( .A(n15913), .B(n15914), .Z(n15910) );
  AND U15623 ( .A(n1256), .B(n15915), .Z(n15914) );
  XOR U15624 ( .A(n15916), .B(n15917), .Z(n15908) );
  AND U15625 ( .A(n1260), .B(n15907), .Z(n15917) );
  XNOR U15626 ( .A(n15918), .B(n15905), .Z(n15907) );
  XOR U15627 ( .A(n15919), .B(n15920), .Z(n15905) );
  AND U15628 ( .A(n1282), .B(n15921), .Z(n15920) );
  IV U15629 ( .A(n15916), .Z(n15918) );
  XOR U15630 ( .A(n15922), .B(n15923), .Z(n15916) );
  AND U15631 ( .A(n1267), .B(n15915), .Z(n15923) );
  XNOR U15632 ( .A(n15913), .B(n15922), .Z(n15915) );
  XNOR U15633 ( .A(n15924), .B(n15925), .Z(n15913) );
  AND U15634 ( .A(n1271), .B(n15926), .Z(n15925) );
  XOR U15635 ( .A(p_input[1942]), .B(n15924), .Z(n15926) );
  XOR U15636 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][22] ), .B(n15927), 
        .Z(n15924) );
  AND U15637 ( .A(n1274), .B(n15928), .Z(n15927) );
  XOR U15638 ( .A(n15929), .B(n15930), .Z(n15922) );
  AND U15639 ( .A(n1278), .B(n15921), .Z(n15930) );
  XNOR U15640 ( .A(n15931), .B(n15919), .Z(n15921) );
  XOR U15641 ( .A(\knn_comb_/min_val_out[0][22] ), .B(n15932), .Z(n15919) );
  AND U15642 ( .A(n1290), .B(n15933), .Z(n15932) );
  IV U15643 ( .A(n15929), .Z(n15931) );
  XOR U15644 ( .A(n15934), .B(n15935), .Z(n15929) );
  AND U15645 ( .A(n1285), .B(n15928), .Z(n15935) );
  XOR U15646 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][22] ), .B(n15934), 
        .Z(n15928) );
  XOR U15647 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .B(n15936), 
        .Z(n15934) );
  AND U15648 ( .A(n1287), .B(n15933), .Z(n15936) );
  XOR U15649 ( .A(\knn_comb_/min_val_out[0][22] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .Z(n15933) );
  XOR U15650 ( .A(n95), .B(n15937), .Z(o[21]) );
  AND U15651 ( .A(n122), .B(n15938), .Z(n95) );
  XOR U15652 ( .A(n96), .B(n15937), .Z(n15938) );
  XOR U15653 ( .A(n15939), .B(n15940), .Z(n15937) );
  AND U15654 ( .A(n142), .B(n15941), .Z(n15940) );
  XOR U15655 ( .A(n15942), .B(n25), .Z(n96) );
  AND U15656 ( .A(n125), .B(n15943), .Z(n25) );
  XOR U15657 ( .A(n26), .B(n15942), .Z(n15943) );
  XOR U15658 ( .A(n15944), .B(n15945), .Z(n26) );
  AND U15659 ( .A(n130), .B(n15946), .Z(n15945) );
  XOR U15660 ( .A(p_input[21]), .B(n15944), .Z(n15946) );
  XNOR U15661 ( .A(n15947), .B(n15948), .Z(n15944) );
  AND U15662 ( .A(n134), .B(n15949), .Z(n15948) );
  XOR U15663 ( .A(n15950), .B(n15951), .Z(n15942) );
  AND U15664 ( .A(n138), .B(n15941), .Z(n15951) );
  XNOR U15665 ( .A(n15952), .B(n15939), .Z(n15941) );
  XOR U15666 ( .A(n15953), .B(n15954), .Z(n15939) );
  AND U15667 ( .A(n162), .B(n15955), .Z(n15954) );
  IV U15668 ( .A(n15950), .Z(n15952) );
  XOR U15669 ( .A(n15956), .B(n15957), .Z(n15950) );
  AND U15670 ( .A(n146), .B(n15949), .Z(n15957) );
  XNOR U15671 ( .A(n15947), .B(n15956), .Z(n15949) );
  XNOR U15672 ( .A(n15958), .B(n15959), .Z(n15947) );
  AND U15673 ( .A(n150), .B(n15960), .Z(n15959) );
  XOR U15674 ( .A(p_input[53]), .B(n15958), .Z(n15960) );
  XNOR U15675 ( .A(n15961), .B(n15962), .Z(n15958) );
  AND U15676 ( .A(n154), .B(n15963), .Z(n15962) );
  XOR U15677 ( .A(n15964), .B(n15965), .Z(n15956) );
  AND U15678 ( .A(n158), .B(n15955), .Z(n15965) );
  XNOR U15679 ( .A(n15966), .B(n15953), .Z(n15955) );
  XOR U15680 ( .A(n15967), .B(n15968), .Z(n15953) );
  AND U15681 ( .A(n181), .B(n15969), .Z(n15968) );
  IV U15682 ( .A(n15964), .Z(n15966) );
  XOR U15683 ( .A(n15970), .B(n15971), .Z(n15964) );
  AND U15684 ( .A(n165), .B(n15963), .Z(n15971) );
  XNOR U15685 ( .A(n15961), .B(n15970), .Z(n15963) );
  XNOR U15686 ( .A(n15972), .B(n15973), .Z(n15961) );
  AND U15687 ( .A(n169), .B(n15974), .Z(n15973) );
  XOR U15688 ( .A(p_input[85]), .B(n15972), .Z(n15974) );
  XNOR U15689 ( .A(n15975), .B(n15976), .Z(n15972) );
  AND U15690 ( .A(n173), .B(n15977), .Z(n15976) );
  XOR U15691 ( .A(n15978), .B(n15979), .Z(n15970) );
  AND U15692 ( .A(n177), .B(n15969), .Z(n15979) );
  XNOR U15693 ( .A(n15980), .B(n15967), .Z(n15969) );
  XOR U15694 ( .A(n15981), .B(n15982), .Z(n15967) );
  AND U15695 ( .A(n200), .B(n15983), .Z(n15982) );
  IV U15696 ( .A(n15978), .Z(n15980) );
  XOR U15697 ( .A(n15984), .B(n15985), .Z(n15978) );
  AND U15698 ( .A(n184), .B(n15977), .Z(n15985) );
  XNOR U15699 ( .A(n15975), .B(n15984), .Z(n15977) );
  XNOR U15700 ( .A(n15986), .B(n15987), .Z(n15975) );
  AND U15701 ( .A(n188), .B(n15988), .Z(n15987) );
  XOR U15702 ( .A(p_input[117]), .B(n15986), .Z(n15988) );
  XNOR U15703 ( .A(n15989), .B(n15990), .Z(n15986) );
  AND U15704 ( .A(n192), .B(n15991), .Z(n15990) );
  XOR U15705 ( .A(n15992), .B(n15993), .Z(n15984) );
  AND U15706 ( .A(n196), .B(n15983), .Z(n15993) );
  XNOR U15707 ( .A(n15994), .B(n15981), .Z(n15983) );
  XOR U15708 ( .A(n15995), .B(n15996), .Z(n15981) );
  AND U15709 ( .A(n219), .B(n15997), .Z(n15996) );
  IV U15710 ( .A(n15992), .Z(n15994) );
  XOR U15711 ( .A(n15998), .B(n15999), .Z(n15992) );
  AND U15712 ( .A(n203), .B(n15991), .Z(n15999) );
  XNOR U15713 ( .A(n15989), .B(n15998), .Z(n15991) );
  XNOR U15714 ( .A(n16000), .B(n16001), .Z(n15989) );
  AND U15715 ( .A(n207), .B(n16002), .Z(n16001) );
  XOR U15716 ( .A(p_input[149]), .B(n16000), .Z(n16002) );
  XNOR U15717 ( .A(n16003), .B(n16004), .Z(n16000) );
  AND U15718 ( .A(n211), .B(n16005), .Z(n16004) );
  XOR U15719 ( .A(n16006), .B(n16007), .Z(n15998) );
  AND U15720 ( .A(n215), .B(n15997), .Z(n16007) );
  XNOR U15721 ( .A(n16008), .B(n15995), .Z(n15997) );
  XOR U15722 ( .A(n16009), .B(n16010), .Z(n15995) );
  AND U15723 ( .A(n238), .B(n16011), .Z(n16010) );
  IV U15724 ( .A(n16006), .Z(n16008) );
  XOR U15725 ( .A(n16012), .B(n16013), .Z(n16006) );
  AND U15726 ( .A(n222), .B(n16005), .Z(n16013) );
  XNOR U15727 ( .A(n16003), .B(n16012), .Z(n16005) );
  XNOR U15728 ( .A(n16014), .B(n16015), .Z(n16003) );
  AND U15729 ( .A(n226), .B(n16016), .Z(n16015) );
  XOR U15730 ( .A(p_input[181]), .B(n16014), .Z(n16016) );
  XNOR U15731 ( .A(n16017), .B(n16018), .Z(n16014) );
  AND U15732 ( .A(n230), .B(n16019), .Z(n16018) );
  XOR U15733 ( .A(n16020), .B(n16021), .Z(n16012) );
  AND U15734 ( .A(n234), .B(n16011), .Z(n16021) );
  XNOR U15735 ( .A(n16022), .B(n16009), .Z(n16011) );
  XOR U15736 ( .A(n16023), .B(n16024), .Z(n16009) );
  AND U15737 ( .A(n257), .B(n16025), .Z(n16024) );
  IV U15738 ( .A(n16020), .Z(n16022) );
  XOR U15739 ( .A(n16026), .B(n16027), .Z(n16020) );
  AND U15740 ( .A(n241), .B(n16019), .Z(n16027) );
  XNOR U15741 ( .A(n16017), .B(n16026), .Z(n16019) );
  XNOR U15742 ( .A(n16028), .B(n16029), .Z(n16017) );
  AND U15743 ( .A(n245), .B(n16030), .Z(n16029) );
  XOR U15744 ( .A(p_input[213]), .B(n16028), .Z(n16030) );
  XNOR U15745 ( .A(n16031), .B(n16032), .Z(n16028) );
  AND U15746 ( .A(n249), .B(n16033), .Z(n16032) );
  XOR U15747 ( .A(n16034), .B(n16035), .Z(n16026) );
  AND U15748 ( .A(n253), .B(n16025), .Z(n16035) );
  XNOR U15749 ( .A(n16036), .B(n16023), .Z(n16025) );
  XOR U15750 ( .A(n16037), .B(n16038), .Z(n16023) );
  AND U15751 ( .A(n276), .B(n16039), .Z(n16038) );
  IV U15752 ( .A(n16034), .Z(n16036) );
  XOR U15753 ( .A(n16040), .B(n16041), .Z(n16034) );
  AND U15754 ( .A(n260), .B(n16033), .Z(n16041) );
  XNOR U15755 ( .A(n16031), .B(n16040), .Z(n16033) );
  XNOR U15756 ( .A(n16042), .B(n16043), .Z(n16031) );
  AND U15757 ( .A(n264), .B(n16044), .Z(n16043) );
  XOR U15758 ( .A(p_input[245]), .B(n16042), .Z(n16044) );
  XNOR U15759 ( .A(n16045), .B(n16046), .Z(n16042) );
  AND U15760 ( .A(n268), .B(n16047), .Z(n16046) );
  XOR U15761 ( .A(n16048), .B(n16049), .Z(n16040) );
  AND U15762 ( .A(n272), .B(n16039), .Z(n16049) );
  XNOR U15763 ( .A(n16050), .B(n16037), .Z(n16039) );
  XOR U15764 ( .A(n16051), .B(n16052), .Z(n16037) );
  AND U15765 ( .A(n295), .B(n16053), .Z(n16052) );
  IV U15766 ( .A(n16048), .Z(n16050) );
  XOR U15767 ( .A(n16054), .B(n16055), .Z(n16048) );
  AND U15768 ( .A(n279), .B(n16047), .Z(n16055) );
  XNOR U15769 ( .A(n16045), .B(n16054), .Z(n16047) );
  XNOR U15770 ( .A(n16056), .B(n16057), .Z(n16045) );
  AND U15771 ( .A(n283), .B(n16058), .Z(n16057) );
  XOR U15772 ( .A(p_input[277]), .B(n16056), .Z(n16058) );
  XNOR U15773 ( .A(n16059), .B(n16060), .Z(n16056) );
  AND U15774 ( .A(n287), .B(n16061), .Z(n16060) );
  XOR U15775 ( .A(n16062), .B(n16063), .Z(n16054) );
  AND U15776 ( .A(n291), .B(n16053), .Z(n16063) );
  XNOR U15777 ( .A(n16064), .B(n16051), .Z(n16053) );
  XOR U15778 ( .A(n16065), .B(n16066), .Z(n16051) );
  AND U15779 ( .A(n314), .B(n16067), .Z(n16066) );
  IV U15780 ( .A(n16062), .Z(n16064) );
  XOR U15781 ( .A(n16068), .B(n16069), .Z(n16062) );
  AND U15782 ( .A(n298), .B(n16061), .Z(n16069) );
  XNOR U15783 ( .A(n16059), .B(n16068), .Z(n16061) );
  XNOR U15784 ( .A(n16070), .B(n16071), .Z(n16059) );
  AND U15785 ( .A(n302), .B(n16072), .Z(n16071) );
  XOR U15786 ( .A(p_input[309]), .B(n16070), .Z(n16072) );
  XNOR U15787 ( .A(n16073), .B(n16074), .Z(n16070) );
  AND U15788 ( .A(n306), .B(n16075), .Z(n16074) );
  XOR U15789 ( .A(n16076), .B(n16077), .Z(n16068) );
  AND U15790 ( .A(n310), .B(n16067), .Z(n16077) );
  XNOR U15791 ( .A(n16078), .B(n16065), .Z(n16067) );
  XOR U15792 ( .A(n16079), .B(n16080), .Z(n16065) );
  AND U15793 ( .A(n333), .B(n16081), .Z(n16080) );
  IV U15794 ( .A(n16076), .Z(n16078) );
  XOR U15795 ( .A(n16082), .B(n16083), .Z(n16076) );
  AND U15796 ( .A(n317), .B(n16075), .Z(n16083) );
  XNOR U15797 ( .A(n16073), .B(n16082), .Z(n16075) );
  XNOR U15798 ( .A(n16084), .B(n16085), .Z(n16073) );
  AND U15799 ( .A(n321), .B(n16086), .Z(n16085) );
  XOR U15800 ( .A(p_input[341]), .B(n16084), .Z(n16086) );
  XNOR U15801 ( .A(n16087), .B(n16088), .Z(n16084) );
  AND U15802 ( .A(n325), .B(n16089), .Z(n16088) );
  XOR U15803 ( .A(n16090), .B(n16091), .Z(n16082) );
  AND U15804 ( .A(n329), .B(n16081), .Z(n16091) );
  XNOR U15805 ( .A(n16092), .B(n16079), .Z(n16081) );
  XOR U15806 ( .A(n16093), .B(n16094), .Z(n16079) );
  AND U15807 ( .A(n352), .B(n16095), .Z(n16094) );
  IV U15808 ( .A(n16090), .Z(n16092) );
  XOR U15809 ( .A(n16096), .B(n16097), .Z(n16090) );
  AND U15810 ( .A(n336), .B(n16089), .Z(n16097) );
  XNOR U15811 ( .A(n16087), .B(n16096), .Z(n16089) );
  XNOR U15812 ( .A(n16098), .B(n16099), .Z(n16087) );
  AND U15813 ( .A(n340), .B(n16100), .Z(n16099) );
  XOR U15814 ( .A(p_input[373]), .B(n16098), .Z(n16100) );
  XNOR U15815 ( .A(n16101), .B(n16102), .Z(n16098) );
  AND U15816 ( .A(n344), .B(n16103), .Z(n16102) );
  XOR U15817 ( .A(n16104), .B(n16105), .Z(n16096) );
  AND U15818 ( .A(n348), .B(n16095), .Z(n16105) );
  XNOR U15819 ( .A(n16106), .B(n16093), .Z(n16095) );
  XOR U15820 ( .A(n16107), .B(n16108), .Z(n16093) );
  AND U15821 ( .A(n371), .B(n16109), .Z(n16108) );
  IV U15822 ( .A(n16104), .Z(n16106) );
  XOR U15823 ( .A(n16110), .B(n16111), .Z(n16104) );
  AND U15824 ( .A(n355), .B(n16103), .Z(n16111) );
  XNOR U15825 ( .A(n16101), .B(n16110), .Z(n16103) );
  XNOR U15826 ( .A(n16112), .B(n16113), .Z(n16101) );
  AND U15827 ( .A(n359), .B(n16114), .Z(n16113) );
  XOR U15828 ( .A(p_input[405]), .B(n16112), .Z(n16114) );
  XNOR U15829 ( .A(n16115), .B(n16116), .Z(n16112) );
  AND U15830 ( .A(n363), .B(n16117), .Z(n16116) );
  XOR U15831 ( .A(n16118), .B(n16119), .Z(n16110) );
  AND U15832 ( .A(n367), .B(n16109), .Z(n16119) );
  XNOR U15833 ( .A(n16120), .B(n16107), .Z(n16109) );
  XOR U15834 ( .A(n16121), .B(n16122), .Z(n16107) );
  AND U15835 ( .A(n390), .B(n16123), .Z(n16122) );
  IV U15836 ( .A(n16118), .Z(n16120) );
  XOR U15837 ( .A(n16124), .B(n16125), .Z(n16118) );
  AND U15838 ( .A(n374), .B(n16117), .Z(n16125) );
  XNOR U15839 ( .A(n16115), .B(n16124), .Z(n16117) );
  XNOR U15840 ( .A(n16126), .B(n16127), .Z(n16115) );
  AND U15841 ( .A(n378), .B(n16128), .Z(n16127) );
  XOR U15842 ( .A(p_input[437]), .B(n16126), .Z(n16128) );
  XNOR U15843 ( .A(n16129), .B(n16130), .Z(n16126) );
  AND U15844 ( .A(n382), .B(n16131), .Z(n16130) );
  XOR U15845 ( .A(n16132), .B(n16133), .Z(n16124) );
  AND U15846 ( .A(n386), .B(n16123), .Z(n16133) );
  XNOR U15847 ( .A(n16134), .B(n16121), .Z(n16123) );
  XOR U15848 ( .A(n16135), .B(n16136), .Z(n16121) );
  AND U15849 ( .A(n409), .B(n16137), .Z(n16136) );
  IV U15850 ( .A(n16132), .Z(n16134) );
  XOR U15851 ( .A(n16138), .B(n16139), .Z(n16132) );
  AND U15852 ( .A(n393), .B(n16131), .Z(n16139) );
  XNOR U15853 ( .A(n16129), .B(n16138), .Z(n16131) );
  XNOR U15854 ( .A(n16140), .B(n16141), .Z(n16129) );
  AND U15855 ( .A(n397), .B(n16142), .Z(n16141) );
  XOR U15856 ( .A(p_input[469]), .B(n16140), .Z(n16142) );
  XNOR U15857 ( .A(n16143), .B(n16144), .Z(n16140) );
  AND U15858 ( .A(n401), .B(n16145), .Z(n16144) );
  XOR U15859 ( .A(n16146), .B(n16147), .Z(n16138) );
  AND U15860 ( .A(n405), .B(n16137), .Z(n16147) );
  XNOR U15861 ( .A(n16148), .B(n16135), .Z(n16137) );
  XOR U15862 ( .A(n16149), .B(n16150), .Z(n16135) );
  AND U15863 ( .A(n428), .B(n16151), .Z(n16150) );
  IV U15864 ( .A(n16146), .Z(n16148) );
  XOR U15865 ( .A(n16152), .B(n16153), .Z(n16146) );
  AND U15866 ( .A(n412), .B(n16145), .Z(n16153) );
  XNOR U15867 ( .A(n16143), .B(n16152), .Z(n16145) );
  XNOR U15868 ( .A(n16154), .B(n16155), .Z(n16143) );
  AND U15869 ( .A(n416), .B(n16156), .Z(n16155) );
  XOR U15870 ( .A(p_input[501]), .B(n16154), .Z(n16156) );
  XNOR U15871 ( .A(n16157), .B(n16158), .Z(n16154) );
  AND U15872 ( .A(n420), .B(n16159), .Z(n16158) );
  XOR U15873 ( .A(n16160), .B(n16161), .Z(n16152) );
  AND U15874 ( .A(n424), .B(n16151), .Z(n16161) );
  XNOR U15875 ( .A(n16162), .B(n16149), .Z(n16151) );
  XOR U15876 ( .A(n16163), .B(n16164), .Z(n16149) );
  AND U15877 ( .A(n447), .B(n16165), .Z(n16164) );
  IV U15878 ( .A(n16160), .Z(n16162) );
  XOR U15879 ( .A(n16166), .B(n16167), .Z(n16160) );
  AND U15880 ( .A(n431), .B(n16159), .Z(n16167) );
  XNOR U15881 ( .A(n16157), .B(n16166), .Z(n16159) );
  XNOR U15882 ( .A(n16168), .B(n16169), .Z(n16157) );
  AND U15883 ( .A(n435), .B(n16170), .Z(n16169) );
  XOR U15884 ( .A(p_input[533]), .B(n16168), .Z(n16170) );
  XNOR U15885 ( .A(n16171), .B(n16172), .Z(n16168) );
  AND U15886 ( .A(n439), .B(n16173), .Z(n16172) );
  XOR U15887 ( .A(n16174), .B(n16175), .Z(n16166) );
  AND U15888 ( .A(n443), .B(n16165), .Z(n16175) );
  XNOR U15889 ( .A(n16176), .B(n16163), .Z(n16165) );
  XOR U15890 ( .A(n16177), .B(n16178), .Z(n16163) );
  AND U15891 ( .A(n466), .B(n16179), .Z(n16178) );
  IV U15892 ( .A(n16174), .Z(n16176) );
  XOR U15893 ( .A(n16180), .B(n16181), .Z(n16174) );
  AND U15894 ( .A(n450), .B(n16173), .Z(n16181) );
  XNOR U15895 ( .A(n16171), .B(n16180), .Z(n16173) );
  XNOR U15896 ( .A(n16182), .B(n16183), .Z(n16171) );
  AND U15897 ( .A(n454), .B(n16184), .Z(n16183) );
  XOR U15898 ( .A(p_input[565]), .B(n16182), .Z(n16184) );
  XNOR U15899 ( .A(n16185), .B(n16186), .Z(n16182) );
  AND U15900 ( .A(n458), .B(n16187), .Z(n16186) );
  XOR U15901 ( .A(n16188), .B(n16189), .Z(n16180) );
  AND U15902 ( .A(n462), .B(n16179), .Z(n16189) );
  XNOR U15903 ( .A(n16190), .B(n16177), .Z(n16179) );
  XOR U15904 ( .A(n16191), .B(n16192), .Z(n16177) );
  AND U15905 ( .A(n485), .B(n16193), .Z(n16192) );
  IV U15906 ( .A(n16188), .Z(n16190) );
  XOR U15907 ( .A(n16194), .B(n16195), .Z(n16188) );
  AND U15908 ( .A(n469), .B(n16187), .Z(n16195) );
  XNOR U15909 ( .A(n16185), .B(n16194), .Z(n16187) );
  XNOR U15910 ( .A(n16196), .B(n16197), .Z(n16185) );
  AND U15911 ( .A(n473), .B(n16198), .Z(n16197) );
  XOR U15912 ( .A(p_input[597]), .B(n16196), .Z(n16198) );
  XNOR U15913 ( .A(n16199), .B(n16200), .Z(n16196) );
  AND U15914 ( .A(n477), .B(n16201), .Z(n16200) );
  XOR U15915 ( .A(n16202), .B(n16203), .Z(n16194) );
  AND U15916 ( .A(n481), .B(n16193), .Z(n16203) );
  XNOR U15917 ( .A(n16204), .B(n16191), .Z(n16193) );
  XOR U15918 ( .A(n16205), .B(n16206), .Z(n16191) );
  AND U15919 ( .A(n504), .B(n16207), .Z(n16206) );
  IV U15920 ( .A(n16202), .Z(n16204) );
  XOR U15921 ( .A(n16208), .B(n16209), .Z(n16202) );
  AND U15922 ( .A(n488), .B(n16201), .Z(n16209) );
  XNOR U15923 ( .A(n16199), .B(n16208), .Z(n16201) );
  XNOR U15924 ( .A(n16210), .B(n16211), .Z(n16199) );
  AND U15925 ( .A(n492), .B(n16212), .Z(n16211) );
  XOR U15926 ( .A(p_input[629]), .B(n16210), .Z(n16212) );
  XNOR U15927 ( .A(n16213), .B(n16214), .Z(n16210) );
  AND U15928 ( .A(n496), .B(n16215), .Z(n16214) );
  XOR U15929 ( .A(n16216), .B(n16217), .Z(n16208) );
  AND U15930 ( .A(n500), .B(n16207), .Z(n16217) );
  XNOR U15931 ( .A(n16218), .B(n16205), .Z(n16207) );
  XOR U15932 ( .A(n16219), .B(n16220), .Z(n16205) );
  AND U15933 ( .A(n523), .B(n16221), .Z(n16220) );
  IV U15934 ( .A(n16216), .Z(n16218) );
  XOR U15935 ( .A(n16222), .B(n16223), .Z(n16216) );
  AND U15936 ( .A(n507), .B(n16215), .Z(n16223) );
  XNOR U15937 ( .A(n16213), .B(n16222), .Z(n16215) );
  XNOR U15938 ( .A(n16224), .B(n16225), .Z(n16213) );
  AND U15939 ( .A(n511), .B(n16226), .Z(n16225) );
  XOR U15940 ( .A(p_input[661]), .B(n16224), .Z(n16226) );
  XNOR U15941 ( .A(n16227), .B(n16228), .Z(n16224) );
  AND U15942 ( .A(n515), .B(n16229), .Z(n16228) );
  XOR U15943 ( .A(n16230), .B(n16231), .Z(n16222) );
  AND U15944 ( .A(n519), .B(n16221), .Z(n16231) );
  XNOR U15945 ( .A(n16232), .B(n16219), .Z(n16221) );
  XOR U15946 ( .A(n16233), .B(n16234), .Z(n16219) );
  AND U15947 ( .A(n542), .B(n16235), .Z(n16234) );
  IV U15948 ( .A(n16230), .Z(n16232) );
  XOR U15949 ( .A(n16236), .B(n16237), .Z(n16230) );
  AND U15950 ( .A(n526), .B(n16229), .Z(n16237) );
  XNOR U15951 ( .A(n16227), .B(n16236), .Z(n16229) );
  XNOR U15952 ( .A(n16238), .B(n16239), .Z(n16227) );
  AND U15953 ( .A(n530), .B(n16240), .Z(n16239) );
  XOR U15954 ( .A(p_input[693]), .B(n16238), .Z(n16240) );
  XNOR U15955 ( .A(n16241), .B(n16242), .Z(n16238) );
  AND U15956 ( .A(n534), .B(n16243), .Z(n16242) );
  XOR U15957 ( .A(n16244), .B(n16245), .Z(n16236) );
  AND U15958 ( .A(n538), .B(n16235), .Z(n16245) );
  XNOR U15959 ( .A(n16246), .B(n16233), .Z(n16235) );
  XOR U15960 ( .A(n16247), .B(n16248), .Z(n16233) );
  AND U15961 ( .A(n561), .B(n16249), .Z(n16248) );
  IV U15962 ( .A(n16244), .Z(n16246) );
  XOR U15963 ( .A(n16250), .B(n16251), .Z(n16244) );
  AND U15964 ( .A(n545), .B(n16243), .Z(n16251) );
  XNOR U15965 ( .A(n16241), .B(n16250), .Z(n16243) );
  XNOR U15966 ( .A(n16252), .B(n16253), .Z(n16241) );
  AND U15967 ( .A(n549), .B(n16254), .Z(n16253) );
  XOR U15968 ( .A(p_input[725]), .B(n16252), .Z(n16254) );
  XNOR U15969 ( .A(n16255), .B(n16256), .Z(n16252) );
  AND U15970 ( .A(n553), .B(n16257), .Z(n16256) );
  XOR U15971 ( .A(n16258), .B(n16259), .Z(n16250) );
  AND U15972 ( .A(n557), .B(n16249), .Z(n16259) );
  XNOR U15973 ( .A(n16260), .B(n16247), .Z(n16249) );
  XOR U15974 ( .A(n16261), .B(n16262), .Z(n16247) );
  AND U15975 ( .A(n580), .B(n16263), .Z(n16262) );
  IV U15976 ( .A(n16258), .Z(n16260) );
  XOR U15977 ( .A(n16264), .B(n16265), .Z(n16258) );
  AND U15978 ( .A(n564), .B(n16257), .Z(n16265) );
  XNOR U15979 ( .A(n16255), .B(n16264), .Z(n16257) );
  XNOR U15980 ( .A(n16266), .B(n16267), .Z(n16255) );
  AND U15981 ( .A(n568), .B(n16268), .Z(n16267) );
  XOR U15982 ( .A(p_input[757]), .B(n16266), .Z(n16268) );
  XNOR U15983 ( .A(n16269), .B(n16270), .Z(n16266) );
  AND U15984 ( .A(n572), .B(n16271), .Z(n16270) );
  XOR U15985 ( .A(n16272), .B(n16273), .Z(n16264) );
  AND U15986 ( .A(n576), .B(n16263), .Z(n16273) );
  XNOR U15987 ( .A(n16274), .B(n16261), .Z(n16263) );
  XOR U15988 ( .A(n16275), .B(n16276), .Z(n16261) );
  AND U15989 ( .A(n599), .B(n16277), .Z(n16276) );
  IV U15990 ( .A(n16272), .Z(n16274) );
  XOR U15991 ( .A(n16278), .B(n16279), .Z(n16272) );
  AND U15992 ( .A(n583), .B(n16271), .Z(n16279) );
  XNOR U15993 ( .A(n16269), .B(n16278), .Z(n16271) );
  XNOR U15994 ( .A(n16280), .B(n16281), .Z(n16269) );
  AND U15995 ( .A(n587), .B(n16282), .Z(n16281) );
  XOR U15996 ( .A(p_input[789]), .B(n16280), .Z(n16282) );
  XNOR U15997 ( .A(n16283), .B(n16284), .Z(n16280) );
  AND U15998 ( .A(n591), .B(n16285), .Z(n16284) );
  XOR U15999 ( .A(n16286), .B(n16287), .Z(n16278) );
  AND U16000 ( .A(n595), .B(n16277), .Z(n16287) );
  XNOR U16001 ( .A(n16288), .B(n16275), .Z(n16277) );
  XOR U16002 ( .A(n16289), .B(n16290), .Z(n16275) );
  AND U16003 ( .A(n618), .B(n16291), .Z(n16290) );
  IV U16004 ( .A(n16286), .Z(n16288) );
  XOR U16005 ( .A(n16292), .B(n16293), .Z(n16286) );
  AND U16006 ( .A(n602), .B(n16285), .Z(n16293) );
  XNOR U16007 ( .A(n16283), .B(n16292), .Z(n16285) );
  XNOR U16008 ( .A(n16294), .B(n16295), .Z(n16283) );
  AND U16009 ( .A(n606), .B(n16296), .Z(n16295) );
  XOR U16010 ( .A(p_input[821]), .B(n16294), .Z(n16296) );
  XNOR U16011 ( .A(n16297), .B(n16298), .Z(n16294) );
  AND U16012 ( .A(n610), .B(n16299), .Z(n16298) );
  XOR U16013 ( .A(n16300), .B(n16301), .Z(n16292) );
  AND U16014 ( .A(n614), .B(n16291), .Z(n16301) );
  XNOR U16015 ( .A(n16302), .B(n16289), .Z(n16291) );
  XOR U16016 ( .A(n16303), .B(n16304), .Z(n16289) );
  AND U16017 ( .A(n637), .B(n16305), .Z(n16304) );
  IV U16018 ( .A(n16300), .Z(n16302) );
  XOR U16019 ( .A(n16306), .B(n16307), .Z(n16300) );
  AND U16020 ( .A(n621), .B(n16299), .Z(n16307) );
  XNOR U16021 ( .A(n16297), .B(n16306), .Z(n16299) );
  XNOR U16022 ( .A(n16308), .B(n16309), .Z(n16297) );
  AND U16023 ( .A(n625), .B(n16310), .Z(n16309) );
  XOR U16024 ( .A(p_input[853]), .B(n16308), .Z(n16310) );
  XNOR U16025 ( .A(n16311), .B(n16312), .Z(n16308) );
  AND U16026 ( .A(n629), .B(n16313), .Z(n16312) );
  XOR U16027 ( .A(n16314), .B(n16315), .Z(n16306) );
  AND U16028 ( .A(n633), .B(n16305), .Z(n16315) );
  XNOR U16029 ( .A(n16316), .B(n16303), .Z(n16305) );
  XOR U16030 ( .A(n16317), .B(n16318), .Z(n16303) );
  AND U16031 ( .A(n656), .B(n16319), .Z(n16318) );
  IV U16032 ( .A(n16314), .Z(n16316) );
  XOR U16033 ( .A(n16320), .B(n16321), .Z(n16314) );
  AND U16034 ( .A(n640), .B(n16313), .Z(n16321) );
  XNOR U16035 ( .A(n16311), .B(n16320), .Z(n16313) );
  XNOR U16036 ( .A(n16322), .B(n16323), .Z(n16311) );
  AND U16037 ( .A(n644), .B(n16324), .Z(n16323) );
  XOR U16038 ( .A(p_input[885]), .B(n16322), .Z(n16324) );
  XNOR U16039 ( .A(n16325), .B(n16326), .Z(n16322) );
  AND U16040 ( .A(n648), .B(n16327), .Z(n16326) );
  XOR U16041 ( .A(n16328), .B(n16329), .Z(n16320) );
  AND U16042 ( .A(n652), .B(n16319), .Z(n16329) );
  XNOR U16043 ( .A(n16330), .B(n16317), .Z(n16319) );
  XOR U16044 ( .A(n16331), .B(n16332), .Z(n16317) );
  AND U16045 ( .A(n675), .B(n16333), .Z(n16332) );
  IV U16046 ( .A(n16328), .Z(n16330) );
  XOR U16047 ( .A(n16334), .B(n16335), .Z(n16328) );
  AND U16048 ( .A(n659), .B(n16327), .Z(n16335) );
  XNOR U16049 ( .A(n16325), .B(n16334), .Z(n16327) );
  XNOR U16050 ( .A(n16336), .B(n16337), .Z(n16325) );
  AND U16051 ( .A(n663), .B(n16338), .Z(n16337) );
  XOR U16052 ( .A(p_input[917]), .B(n16336), .Z(n16338) );
  XNOR U16053 ( .A(n16339), .B(n16340), .Z(n16336) );
  AND U16054 ( .A(n667), .B(n16341), .Z(n16340) );
  XOR U16055 ( .A(n16342), .B(n16343), .Z(n16334) );
  AND U16056 ( .A(n671), .B(n16333), .Z(n16343) );
  XNOR U16057 ( .A(n16344), .B(n16331), .Z(n16333) );
  XOR U16058 ( .A(n16345), .B(n16346), .Z(n16331) );
  AND U16059 ( .A(n694), .B(n16347), .Z(n16346) );
  IV U16060 ( .A(n16342), .Z(n16344) );
  XOR U16061 ( .A(n16348), .B(n16349), .Z(n16342) );
  AND U16062 ( .A(n678), .B(n16341), .Z(n16349) );
  XNOR U16063 ( .A(n16339), .B(n16348), .Z(n16341) );
  XNOR U16064 ( .A(n16350), .B(n16351), .Z(n16339) );
  AND U16065 ( .A(n682), .B(n16352), .Z(n16351) );
  XOR U16066 ( .A(p_input[949]), .B(n16350), .Z(n16352) );
  XNOR U16067 ( .A(n16353), .B(n16354), .Z(n16350) );
  AND U16068 ( .A(n686), .B(n16355), .Z(n16354) );
  XOR U16069 ( .A(n16356), .B(n16357), .Z(n16348) );
  AND U16070 ( .A(n690), .B(n16347), .Z(n16357) );
  XNOR U16071 ( .A(n16358), .B(n16345), .Z(n16347) );
  XOR U16072 ( .A(n16359), .B(n16360), .Z(n16345) );
  AND U16073 ( .A(n713), .B(n16361), .Z(n16360) );
  IV U16074 ( .A(n16356), .Z(n16358) );
  XOR U16075 ( .A(n16362), .B(n16363), .Z(n16356) );
  AND U16076 ( .A(n697), .B(n16355), .Z(n16363) );
  XNOR U16077 ( .A(n16353), .B(n16362), .Z(n16355) );
  XNOR U16078 ( .A(n16364), .B(n16365), .Z(n16353) );
  AND U16079 ( .A(n701), .B(n16366), .Z(n16365) );
  XOR U16080 ( .A(p_input[981]), .B(n16364), .Z(n16366) );
  XNOR U16081 ( .A(n16367), .B(n16368), .Z(n16364) );
  AND U16082 ( .A(n705), .B(n16369), .Z(n16368) );
  XOR U16083 ( .A(n16370), .B(n16371), .Z(n16362) );
  AND U16084 ( .A(n709), .B(n16361), .Z(n16371) );
  XNOR U16085 ( .A(n16372), .B(n16359), .Z(n16361) );
  XOR U16086 ( .A(n16373), .B(n16374), .Z(n16359) );
  AND U16087 ( .A(n732), .B(n16375), .Z(n16374) );
  IV U16088 ( .A(n16370), .Z(n16372) );
  XOR U16089 ( .A(n16376), .B(n16377), .Z(n16370) );
  AND U16090 ( .A(n716), .B(n16369), .Z(n16377) );
  XNOR U16091 ( .A(n16367), .B(n16376), .Z(n16369) );
  XNOR U16092 ( .A(n16378), .B(n16379), .Z(n16367) );
  AND U16093 ( .A(n720), .B(n16380), .Z(n16379) );
  XOR U16094 ( .A(p_input[1013]), .B(n16378), .Z(n16380) );
  XNOR U16095 ( .A(n16381), .B(n16382), .Z(n16378) );
  AND U16096 ( .A(n724), .B(n16383), .Z(n16382) );
  XOR U16097 ( .A(n16384), .B(n16385), .Z(n16376) );
  AND U16098 ( .A(n728), .B(n16375), .Z(n16385) );
  XNOR U16099 ( .A(n16386), .B(n16373), .Z(n16375) );
  XOR U16100 ( .A(n16387), .B(n16388), .Z(n16373) );
  AND U16101 ( .A(n751), .B(n16389), .Z(n16388) );
  IV U16102 ( .A(n16384), .Z(n16386) );
  XOR U16103 ( .A(n16390), .B(n16391), .Z(n16384) );
  AND U16104 ( .A(n735), .B(n16383), .Z(n16391) );
  XNOR U16105 ( .A(n16381), .B(n16390), .Z(n16383) );
  XNOR U16106 ( .A(n16392), .B(n16393), .Z(n16381) );
  AND U16107 ( .A(n739), .B(n16394), .Z(n16393) );
  XOR U16108 ( .A(p_input[1045]), .B(n16392), .Z(n16394) );
  XNOR U16109 ( .A(n16395), .B(n16396), .Z(n16392) );
  AND U16110 ( .A(n743), .B(n16397), .Z(n16396) );
  XOR U16111 ( .A(n16398), .B(n16399), .Z(n16390) );
  AND U16112 ( .A(n747), .B(n16389), .Z(n16399) );
  XNOR U16113 ( .A(n16400), .B(n16387), .Z(n16389) );
  XOR U16114 ( .A(n16401), .B(n16402), .Z(n16387) );
  AND U16115 ( .A(n770), .B(n16403), .Z(n16402) );
  IV U16116 ( .A(n16398), .Z(n16400) );
  XOR U16117 ( .A(n16404), .B(n16405), .Z(n16398) );
  AND U16118 ( .A(n754), .B(n16397), .Z(n16405) );
  XNOR U16119 ( .A(n16395), .B(n16404), .Z(n16397) );
  XNOR U16120 ( .A(n16406), .B(n16407), .Z(n16395) );
  AND U16121 ( .A(n758), .B(n16408), .Z(n16407) );
  XOR U16122 ( .A(p_input[1077]), .B(n16406), .Z(n16408) );
  XNOR U16123 ( .A(n16409), .B(n16410), .Z(n16406) );
  AND U16124 ( .A(n762), .B(n16411), .Z(n16410) );
  XOR U16125 ( .A(n16412), .B(n16413), .Z(n16404) );
  AND U16126 ( .A(n766), .B(n16403), .Z(n16413) );
  XNOR U16127 ( .A(n16414), .B(n16401), .Z(n16403) );
  XOR U16128 ( .A(n16415), .B(n16416), .Z(n16401) );
  AND U16129 ( .A(n789), .B(n16417), .Z(n16416) );
  IV U16130 ( .A(n16412), .Z(n16414) );
  XOR U16131 ( .A(n16418), .B(n16419), .Z(n16412) );
  AND U16132 ( .A(n773), .B(n16411), .Z(n16419) );
  XNOR U16133 ( .A(n16409), .B(n16418), .Z(n16411) );
  XNOR U16134 ( .A(n16420), .B(n16421), .Z(n16409) );
  AND U16135 ( .A(n777), .B(n16422), .Z(n16421) );
  XOR U16136 ( .A(p_input[1109]), .B(n16420), .Z(n16422) );
  XNOR U16137 ( .A(n16423), .B(n16424), .Z(n16420) );
  AND U16138 ( .A(n781), .B(n16425), .Z(n16424) );
  XOR U16139 ( .A(n16426), .B(n16427), .Z(n16418) );
  AND U16140 ( .A(n785), .B(n16417), .Z(n16427) );
  XNOR U16141 ( .A(n16428), .B(n16415), .Z(n16417) );
  XOR U16142 ( .A(n16429), .B(n16430), .Z(n16415) );
  AND U16143 ( .A(n808), .B(n16431), .Z(n16430) );
  IV U16144 ( .A(n16426), .Z(n16428) );
  XOR U16145 ( .A(n16432), .B(n16433), .Z(n16426) );
  AND U16146 ( .A(n792), .B(n16425), .Z(n16433) );
  XNOR U16147 ( .A(n16423), .B(n16432), .Z(n16425) );
  XNOR U16148 ( .A(n16434), .B(n16435), .Z(n16423) );
  AND U16149 ( .A(n796), .B(n16436), .Z(n16435) );
  XOR U16150 ( .A(p_input[1141]), .B(n16434), .Z(n16436) );
  XNOR U16151 ( .A(n16437), .B(n16438), .Z(n16434) );
  AND U16152 ( .A(n800), .B(n16439), .Z(n16438) );
  XOR U16153 ( .A(n16440), .B(n16441), .Z(n16432) );
  AND U16154 ( .A(n804), .B(n16431), .Z(n16441) );
  XNOR U16155 ( .A(n16442), .B(n16429), .Z(n16431) );
  XOR U16156 ( .A(n16443), .B(n16444), .Z(n16429) );
  AND U16157 ( .A(n827), .B(n16445), .Z(n16444) );
  IV U16158 ( .A(n16440), .Z(n16442) );
  XOR U16159 ( .A(n16446), .B(n16447), .Z(n16440) );
  AND U16160 ( .A(n811), .B(n16439), .Z(n16447) );
  XNOR U16161 ( .A(n16437), .B(n16446), .Z(n16439) );
  XNOR U16162 ( .A(n16448), .B(n16449), .Z(n16437) );
  AND U16163 ( .A(n815), .B(n16450), .Z(n16449) );
  XOR U16164 ( .A(p_input[1173]), .B(n16448), .Z(n16450) );
  XNOR U16165 ( .A(n16451), .B(n16452), .Z(n16448) );
  AND U16166 ( .A(n819), .B(n16453), .Z(n16452) );
  XOR U16167 ( .A(n16454), .B(n16455), .Z(n16446) );
  AND U16168 ( .A(n823), .B(n16445), .Z(n16455) );
  XNOR U16169 ( .A(n16456), .B(n16443), .Z(n16445) );
  XOR U16170 ( .A(n16457), .B(n16458), .Z(n16443) );
  AND U16171 ( .A(n846), .B(n16459), .Z(n16458) );
  IV U16172 ( .A(n16454), .Z(n16456) );
  XOR U16173 ( .A(n16460), .B(n16461), .Z(n16454) );
  AND U16174 ( .A(n830), .B(n16453), .Z(n16461) );
  XNOR U16175 ( .A(n16451), .B(n16460), .Z(n16453) );
  XNOR U16176 ( .A(n16462), .B(n16463), .Z(n16451) );
  AND U16177 ( .A(n834), .B(n16464), .Z(n16463) );
  XOR U16178 ( .A(p_input[1205]), .B(n16462), .Z(n16464) );
  XNOR U16179 ( .A(n16465), .B(n16466), .Z(n16462) );
  AND U16180 ( .A(n838), .B(n16467), .Z(n16466) );
  XOR U16181 ( .A(n16468), .B(n16469), .Z(n16460) );
  AND U16182 ( .A(n842), .B(n16459), .Z(n16469) );
  XNOR U16183 ( .A(n16470), .B(n16457), .Z(n16459) );
  XOR U16184 ( .A(n16471), .B(n16472), .Z(n16457) );
  AND U16185 ( .A(n865), .B(n16473), .Z(n16472) );
  IV U16186 ( .A(n16468), .Z(n16470) );
  XOR U16187 ( .A(n16474), .B(n16475), .Z(n16468) );
  AND U16188 ( .A(n849), .B(n16467), .Z(n16475) );
  XNOR U16189 ( .A(n16465), .B(n16474), .Z(n16467) );
  XNOR U16190 ( .A(n16476), .B(n16477), .Z(n16465) );
  AND U16191 ( .A(n853), .B(n16478), .Z(n16477) );
  XOR U16192 ( .A(p_input[1237]), .B(n16476), .Z(n16478) );
  XNOR U16193 ( .A(n16479), .B(n16480), .Z(n16476) );
  AND U16194 ( .A(n857), .B(n16481), .Z(n16480) );
  XOR U16195 ( .A(n16482), .B(n16483), .Z(n16474) );
  AND U16196 ( .A(n861), .B(n16473), .Z(n16483) );
  XNOR U16197 ( .A(n16484), .B(n16471), .Z(n16473) );
  XOR U16198 ( .A(n16485), .B(n16486), .Z(n16471) );
  AND U16199 ( .A(n884), .B(n16487), .Z(n16486) );
  IV U16200 ( .A(n16482), .Z(n16484) );
  XOR U16201 ( .A(n16488), .B(n16489), .Z(n16482) );
  AND U16202 ( .A(n868), .B(n16481), .Z(n16489) );
  XNOR U16203 ( .A(n16479), .B(n16488), .Z(n16481) );
  XNOR U16204 ( .A(n16490), .B(n16491), .Z(n16479) );
  AND U16205 ( .A(n872), .B(n16492), .Z(n16491) );
  XOR U16206 ( .A(p_input[1269]), .B(n16490), .Z(n16492) );
  XNOR U16207 ( .A(n16493), .B(n16494), .Z(n16490) );
  AND U16208 ( .A(n876), .B(n16495), .Z(n16494) );
  XOR U16209 ( .A(n16496), .B(n16497), .Z(n16488) );
  AND U16210 ( .A(n880), .B(n16487), .Z(n16497) );
  XNOR U16211 ( .A(n16498), .B(n16485), .Z(n16487) );
  XOR U16212 ( .A(n16499), .B(n16500), .Z(n16485) );
  AND U16213 ( .A(n903), .B(n16501), .Z(n16500) );
  IV U16214 ( .A(n16496), .Z(n16498) );
  XOR U16215 ( .A(n16502), .B(n16503), .Z(n16496) );
  AND U16216 ( .A(n887), .B(n16495), .Z(n16503) );
  XNOR U16217 ( .A(n16493), .B(n16502), .Z(n16495) );
  XNOR U16218 ( .A(n16504), .B(n16505), .Z(n16493) );
  AND U16219 ( .A(n891), .B(n16506), .Z(n16505) );
  XOR U16220 ( .A(p_input[1301]), .B(n16504), .Z(n16506) );
  XNOR U16221 ( .A(n16507), .B(n16508), .Z(n16504) );
  AND U16222 ( .A(n895), .B(n16509), .Z(n16508) );
  XOR U16223 ( .A(n16510), .B(n16511), .Z(n16502) );
  AND U16224 ( .A(n899), .B(n16501), .Z(n16511) );
  XNOR U16225 ( .A(n16512), .B(n16499), .Z(n16501) );
  XOR U16226 ( .A(n16513), .B(n16514), .Z(n16499) );
  AND U16227 ( .A(n922), .B(n16515), .Z(n16514) );
  IV U16228 ( .A(n16510), .Z(n16512) );
  XOR U16229 ( .A(n16516), .B(n16517), .Z(n16510) );
  AND U16230 ( .A(n906), .B(n16509), .Z(n16517) );
  XNOR U16231 ( .A(n16507), .B(n16516), .Z(n16509) );
  XNOR U16232 ( .A(n16518), .B(n16519), .Z(n16507) );
  AND U16233 ( .A(n910), .B(n16520), .Z(n16519) );
  XOR U16234 ( .A(p_input[1333]), .B(n16518), .Z(n16520) );
  XNOR U16235 ( .A(n16521), .B(n16522), .Z(n16518) );
  AND U16236 ( .A(n914), .B(n16523), .Z(n16522) );
  XOR U16237 ( .A(n16524), .B(n16525), .Z(n16516) );
  AND U16238 ( .A(n918), .B(n16515), .Z(n16525) );
  XNOR U16239 ( .A(n16526), .B(n16513), .Z(n16515) );
  XOR U16240 ( .A(n16527), .B(n16528), .Z(n16513) );
  AND U16241 ( .A(n941), .B(n16529), .Z(n16528) );
  IV U16242 ( .A(n16524), .Z(n16526) );
  XOR U16243 ( .A(n16530), .B(n16531), .Z(n16524) );
  AND U16244 ( .A(n925), .B(n16523), .Z(n16531) );
  XNOR U16245 ( .A(n16521), .B(n16530), .Z(n16523) );
  XNOR U16246 ( .A(n16532), .B(n16533), .Z(n16521) );
  AND U16247 ( .A(n929), .B(n16534), .Z(n16533) );
  XOR U16248 ( .A(p_input[1365]), .B(n16532), .Z(n16534) );
  XNOR U16249 ( .A(n16535), .B(n16536), .Z(n16532) );
  AND U16250 ( .A(n933), .B(n16537), .Z(n16536) );
  XOR U16251 ( .A(n16538), .B(n16539), .Z(n16530) );
  AND U16252 ( .A(n937), .B(n16529), .Z(n16539) );
  XNOR U16253 ( .A(n16540), .B(n16527), .Z(n16529) );
  XOR U16254 ( .A(n16541), .B(n16542), .Z(n16527) );
  AND U16255 ( .A(n960), .B(n16543), .Z(n16542) );
  IV U16256 ( .A(n16538), .Z(n16540) );
  XOR U16257 ( .A(n16544), .B(n16545), .Z(n16538) );
  AND U16258 ( .A(n944), .B(n16537), .Z(n16545) );
  XNOR U16259 ( .A(n16535), .B(n16544), .Z(n16537) );
  XNOR U16260 ( .A(n16546), .B(n16547), .Z(n16535) );
  AND U16261 ( .A(n948), .B(n16548), .Z(n16547) );
  XOR U16262 ( .A(p_input[1397]), .B(n16546), .Z(n16548) );
  XNOR U16263 ( .A(n16549), .B(n16550), .Z(n16546) );
  AND U16264 ( .A(n952), .B(n16551), .Z(n16550) );
  XOR U16265 ( .A(n16552), .B(n16553), .Z(n16544) );
  AND U16266 ( .A(n956), .B(n16543), .Z(n16553) );
  XNOR U16267 ( .A(n16554), .B(n16541), .Z(n16543) );
  XOR U16268 ( .A(n16555), .B(n16556), .Z(n16541) );
  AND U16269 ( .A(n979), .B(n16557), .Z(n16556) );
  IV U16270 ( .A(n16552), .Z(n16554) );
  XOR U16271 ( .A(n16558), .B(n16559), .Z(n16552) );
  AND U16272 ( .A(n963), .B(n16551), .Z(n16559) );
  XNOR U16273 ( .A(n16549), .B(n16558), .Z(n16551) );
  XNOR U16274 ( .A(n16560), .B(n16561), .Z(n16549) );
  AND U16275 ( .A(n967), .B(n16562), .Z(n16561) );
  XOR U16276 ( .A(p_input[1429]), .B(n16560), .Z(n16562) );
  XNOR U16277 ( .A(n16563), .B(n16564), .Z(n16560) );
  AND U16278 ( .A(n971), .B(n16565), .Z(n16564) );
  XOR U16279 ( .A(n16566), .B(n16567), .Z(n16558) );
  AND U16280 ( .A(n975), .B(n16557), .Z(n16567) );
  XNOR U16281 ( .A(n16568), .B(n16555), .Z(n16557) );
  XOR U16282 ( .A(n16569), .B(n16570), .Z(n16555) );
  AND U16283 ( .A(n998), .B(n16571), .Z(n16570) );
  IV U16284 ( .A(n16566), .Z(n16568) );
  XOR U16285 ( .A(n16572), .B(n16573), .Z(n16566) );
  AND U16286 ( .A(n982), .B(n16565), .Z(n16573) );
  XNOR U16287 ( .A(n16563), .B(n16572), .Z(n16565) );
  XNOR U16288 ( .A(n16574), .B(n16575), .Z(n16563) );
  AND U16289 ( .A(n986), .B(n16576), .Z(n16575) );
  XOR U16290 ( .A(p_input[1461]), .B(n16574), .Z(n16576) );
  XNOR U16291 ( .A(n16577), .B(n16578), .Z(n16574) );
  AND U16292 ( .A(n990), .B(n16579), .Z(n16578) );
  XOR U16293 ( .A(n16580), .B(n16581), .Z(n16572) );
  AND U16294 ( .A(n994), .B(n16571), .Z(n16581) );
  XNOR U16295 ( .A(n16582), .B(n16569), .Z(n16571) );
  XOR U16296 ( .A(n16583), .B(n16584), .Z(n16569) );
  AND U16297 ( .A(n1017), .B(n16585), .Z(n16584) );
  IV U16298 ( .A(n16580), .Z(n16582) );
  XOR U16299 ( .A(n16586), .B(n16587), .Z(n16580) );
  AND U16300 ( .A(n1001), .B(n16579), .Z(n16587) );
  XNOR U16301 ( .A(n16577), .B(n16586), .Z(n16579) );
  XNOR U16302 ( .A(n16588), .B(n16589), .Z(n16577) );
  AND U16303 ( .A(n1005), .B(n16590), .Z(n16589) );
  XOR U16304 ( .A(p_input[1493]), .B(n16588), .Z(n16590) );
  XNOR U16305 ( .A(n16591), .B(n16592), .Z(n16588) );
  AND U16306 ( .A(n1009), .B(n16593), .Z(n16592) );
  XOR U16307 ( .A(n16594), .B(n16595), .Z(n16586) );
  AND U16308 ( .A(n1013), .B(n16585), .Z(n16595) );
  XNOR U16309 ( .A(n16596), .B(n16583), .Z(n16585) );
  XOR U16310 ( .A(n16597), .B(n16598), .Z(n16583) );
  AND U16311 ( .A(n1036), .B(n16599), .Z(n16598) );
  IV U16312 ( .A(n16594), .Z(n16596) );
  XOR U16313 ( .A(n16600), .B(n16601), .Z(n16594) );
  AND U16314 ( .A(n1020), .B(n16593), .Z(n16601) );
  XNOR U16315 ( .A(n16591), .B(n16600), .Z(n16593) );
  XNOR U16316 ( .A(n16602), .B(n16603), .Z(n16591) );
  AND U16317 ( .A(n1024), .B(n16604), .Z(n16603) );
  XOR U16318 ( .A(p_input[1525]), .B(n16602), .Z(n16604) );
  XNOR U16319 ( .A(n16605), .B(n16606), .Z(n16602) );
  AND U16320 ( .A(n1028), .B(n16607), .Z(n16606) );
  XOR U16321 ( .A(n16608), .B(n16609), .Z(n16600) );
  AND U16322 ( .A(n1032), .B(n16599), .Z(n16609) );
  XNOR U16323 ( .A(n16610), .B(n16597), .Z(n16599) );
  XOR U16324 ( .A(n16611), .B(n16612), .Z(n16597) );
  AND U16325 ( .A(n1055), .B(n16613), .Z(n16612) );
  IV U16326 ( .A(n16608), .Z(n16610) );
  XOR U16327 ( .A(n16614), .B(n16615), .Z(n16608) );
  AND U16328 ( .A(n1039), .B(n16607), .Z(n16615) );
  XNOR U16329 ( .A(n16605), .B(n16614), .Z(n16607) );
  XNOR U16330 ( .A(n16616), .B(n16617), .Z(n16605) );
  AND U16331 ( .A(n1043), .B(n16618), .Z(n16617) );
  XOR U16332 ( .A(p_input[1557]), .B(n16616), .Z(n16618) );
  XNOR U16333 ( .A(n16619), .B(n16620), .Z(n16616) );
  AND U16334 ( .A(n1047), .B(n16621), .Z(n16620) );
  XOR U16335 ( .A(n16622), .B(n16623), .Z(n16614) );
  AND U16336 ( .A(n1051), .B(n16613), .Z(n16623) );
  XNOR U16337 ( .A(n16624), .B(n16611), .Z(n16613) );
  XOR U16338 ( .A(n16625), .B(n16626), .Z(n16611) );
  AND U16339 ( .A(n1074), .B(n16627), .Z(n16626) );
  IV U16340 ( .A(n16622), .Z(n16624) );
  XOR U16341 ( .A(n16628), .B(n16629), .Z(n16622) );
  AND U16342 ( .A(n1058), .B(n16621), .Z(n16629) );
  XNOR U16343 ( .A(n16619), .B(n16628), .Z(n16621) );
  XNOR U16344 ( .A(n16630), .B(n16631), .Z(n16619) );
  AND U16345 ( .A(n1062), .B(n16632), .Z(n16631) );
  XOR U16346 ( .A(p_input[1589]), .B(n16630), .Z(n16632) );
  XNOR U16347 ( .A(n16633), .B(n16634), .Z(n16630) );
  AND U16348 ( .A(n1066), .B(n16635), .Z(n16634) );
  XOR U16349 ( .A(n16636), .B(n16637), .Z(n16628) );
  AND U16350 ( .A(n1070), .B(n16627), .Z(n16637) );
  XNOR U16351 ( .A(n16638), .B(n16625), .Z(n16627) );
  XOR U16352 ( .A(n16639), .B(n16640), .Z(n16625) );
  AND U16353 ( .A(n1093), .B(n16641), .Z(n16640) );
  IV U16354 ( .A(n16636), .Z(n16638) );
  XOR U16355 ( .A(n16642), .B(n16643), .Z(n16636) );
  AND U16356 ( .A(n1077), .B(n16635), .Z(n16643) );
  XNOR U16357 ( .A(n16633), .B(n16642), .Z(n16635) );
  XNOR U16358 ( .A(n16644), .B(n16645), .Z(n16633) );
  AND U16359 ( .A(n1081), .B(n16646), .Z(n16645) );
  XOR U16360 ( .A(p_input[1621]), .B(n16644), .Z(n16646) );
  XNOR U16361 ( .A(n16647), .B(n16648), .Z(n16644) );
  AND U16362 ( .A(n1085), .B(n16649), .Z(n16648) );
  XOR U16363 ( .A(n16650), .B(n16651), .Z(n16642) );
  AND U16364 ( .A(n1089), .B(n16641), .Z(n16651) );
  XNOR U16365 ( .A(n16652), .B(n16639), .Z(n16641) );
  XOR U16366 ( .A(n16653), .B(n16654), .Z(n16639) );
  AND U16367 ( .A(n1112), .B(n16655), .Z(n16654) );
  IV U16368 ( .A(n16650), .Z(n16652) );
  XOR U16369 ( .A(n16656), .B(n16657), .Z(n16650) );
  AND U16370 ( .A(n1096), .B(n16649), .Z(n16657) );
  XNOR U16371 ( .A(n16647), .B(n16656), .Z(n16649) );
  XNOR U16372 ( .A(n16658), .B(n16659), .Z(n16647) );
  AND U16373 ( .A(n1100), .B(n16660), .Z(n16659) );
  XOR U16374 ( .A(p_input[1653]), .B(n16658), .Z(n16660) );
  XNOR U16375 ( .A(n16661), .B(n16662), .Z(n16658) );
  AND U16376 ( .A(n1104), .B(n16663), .Z(n16662) );
  XOR U16377 ( .A(n16664), .B(n16665), .Z(n16656) );
  AND U16378 ( .A(n1108), .B(n16655), .Z(n16665) );
  XNOR U16379 ( .A(n16666), .B(n16653), .Z(n16655) );
  XOR U16380 ( .A(n16667), .B(n16668), .Z(n16653) );
  AND U16381 ( .A(n1131), .B(n16669), .Z(n16668) );
  IV U16382 ( .A(n16664), .Z(n16666) );
  XOR U16383 ( .A(n16670), .B(n16671), .Z(n16664) );
  AND U16384 ( .A(n1115), .B(n16663), .Z(n16671) );
  XNOR U16385 ( .A(n16661), .B(n16670), .Z(n16663) );
  XNOR U16386 ( .A(n16672), .B(n16673), .Z(n16661) );
  AND U16387 ( .A(n1119), .B(n16674), .Z(n16673) );
  XOR U16388 ( .A(p_input[1685]), .B(n16672), .Z(n16674) );
  XNOR U16389 ( .A(n16675), .B(n16676), .Z(n16672) );
  AND U16390 ( .A(n1123), .B(n16677), .Z(n16676) );
  XOR U16391 ( .A(n16678), .B(n16679), .Z(n16670) );
  AND U16392 ( .A(n1127), .B(n16669), .Z(n16679) );
  XNOR U16393 ( .A(n16680), .B(n16667), .Z(n16669) );
  XOR U16394 ( .A(n16681), .B(n16682), .Z(n16667) );
  AND U16395 ( .A(n1150), .B(n16683), .Z(n16682) );
  IV U16396 ( .A(n16678), .Z(n16680) );
  XOR U16397 ( .A(n16684), .B(n16685), .Z(n16678) );
  AND U16398 ( .A(n1134), .B(n16677), .Z(n16685) );
  XNOR U16399 ( .A(n16675), .B(n16684), .Z(n16677) );
  XNOR U16400 ( .A(n16686), .B(n16687), .Z(n16675) );
  AND U16401 ( .A(n1138), .B(n16688), .Z(n16687) );
  XOR U16402 ( .A(p_input[1717]), .B(n16686), .Z(n16688) );
  XNOR U16403 ( .A(n16689), .B(n16690), .Z(n16686) );
  AND U16404 ( .A(n1142), .B(n16691), .Z(n16690) );
  XOR U16405 ( .A(n16692), .B(n16693), .Z(n16684) );
  AND U16406 ( .A(n1146), .B(n16683), .Z(n16693) );
  XNOR U16407 ( .A(n16694), .B(n16681), .Z(n16683) );
  XOR U16408 ( .A(n16695), .B(n16696), .Z(n16681) );
  AND U16409 ( .A(n1169), .B(n16697), .Z(n16696) );
  IV U16410 ( .A(n16692), .Z(n16694) );
  XOR U16411 ( .A(n16698), .B(n16699), .Z(n16692) );
  AND U16412 ( .A(n1153), .B(n16691), .Z(n16699) );
  XNOR U16413 ( .A(n16689), .B(n16698), .Z(n16691) );
  XNOR U16414 ( .A(n16700), .B(n16701), .Z(n16689) );
  AND U16415 ( .A(n1157), .B(n16702), .Z(n16701) );
  XOR U16416 ( .A(p_input[1749]), .B(n16700), .Z(n16702) );
  XNOR U16417 ( .A(n16703), .B(n16704), .Z(n16700) );
  AND U16418 ( .A(n1161), .B(n16705), .Z(n16704) );
  XOR U16419 ( .A(n16706), .B(n16707), .Z(n16698) );
  AND U16420 ( .A(n1165), .B(n16697), .Z(n16707) );
  XNOR U16421 ( .A(n16708), .B(n16695), .Z(n16697) );
  XOR U16422 ( .A(n16709), .B(n16710), .Z(n16695) );
  AND U16423 ( .A(n1188), .B(n16711), .Z(n16710) );
  IV U16424 ( .A(n16706), .Z(n16708) );
  XOR U16425 ( .A(n16712), .B(n16713), .Z(n16706) );
  AND U16426 ( .A(n1172), .B(n16705), .Z(n16713) );
  XNOR U16427 ( .A(n16703), .B(n16712), .Z(n16705) );
  XNOR U16428 ( .A(n16714), .B(n16715), .Z(n16703) );
  AND U16429 ( .A(n1176), .B(n16716), .Z(n16715) );
  XOR U16430 ( .A(p_input[1781]), .B(n16714), .Z(n16716) );
  XNOR U16431 ( .A(n16717), .B(n16718), .Z(n16714) );
  AND U16432 ( .A(n1180), .B(n16719), .Z(n16718) );
  XOR U16433 ( .A(n16720), .B(n16721), .Z(n16712) );
  AND U16434 ( .A(n1184), .B(n16711), .Z(n16721) );
  XNOR U16435 ( .A(n16722), .B(n16709), .Z(n16711) );
  XOR U16436 ( .A(n16723), .B(n16724), .Z(n16709) );
  AND U16437 ( .A(n1207), .B(n16725), .Z(n16724) );
  IV U16438 ( .A(n16720), .Z(n16722) );
  XOR U16439 ( .A(n16726), .B(n16727), .Z(n16720) );
  AND U16440 ( .A(n1191), .B(n16719), .Z(n16727) );
  XNOR U16441 ( .A(n16717), .B(n16726), .Z(n16719) );
  XNOR U16442 ( .A(n16728), .B(n16729), .Z(n16717) );
  AND U16443 ( .A(n1195), .B(n16730), .Z(n16729) );
  XOR U16444 ( .A(p_input[1813]), .B(n16728), .Z(n16730) );
  XNOR U16445 ( .A(n16731), .B(n16732), .Z(n16728) );
  AND U16446 ( .A(n1199), .B(n16733), .Z(n16732) );
  XOR U16447 ( .A(n16734), .B(n16735), .Z(n16726) );
  AND U16448 ( .A(n1203), .B(n16725), .Z(n16735) );
  XNOR U16449 ( .A(n16736), .B(n16723), .Z(n16725) );
  XOR U16450 ( .A(n16737), .B(n16738), .Z(n16723) );
  AND U16451 ( .A(n1226), .B(n16739), .Z(n16738) );
  IV U16452 ( .A(n16734), .Z(n16736) );
  XOR U16453 ( .A(n16740), .B(n16741), .Z(n16734) );
  AND U16454 ( .A(n1210), .B(n16733), .Z(n16741) );
  XNOR U16455 ( .A(n16731), .B(n16740), .Z(n16733) );
  XNOR U16456 ( .A(n16742), .B(n16743), .Z(n16731) );
  AND U16457 ( .A(n1214), .B(n16744), .Z(n16743) );
  XOR U16458 ( .A(p_input[1845]), .B(n16742), .Z(n16744) );
  XNOR U16459 ( .A(n16745), .B(n16746), .Z(n16742) );
  AND U16460 ( .A(n1218), .B(n16747), .Z(n16746) );
  XOR U16461 ( .A(n16748), .B(n16749), .Z(n16740) );
  AND U16462 ( .A(n1222), .B(n16739), .Z(n16749) );
  XNOR U16463 ( .A(n16750), .B(n16737), .Z(n16739) );
  XOR U16464 ( .A(n16751), .B(n16752), .Z(n16737) );
  AND U16465 ( .A(n1245), .B(n16753), .Z(n16752) );
  IV U16466 ( .A(n16748), .Z(n16750) );
  XOR U16467 ( .A(n16754), .B(n16755), .Z(n16748) );
  AND U16468 ( .A(n1229), .B(n16747), .Z(n16755) );
  XNOR U16469 ( .A(n16745), .B(n16754), .Z(n16747) );
  XNOR U16470 ( .A(n16756), .B(n16757), .Z(n16745) );
  AND U16471 ( .A(n1233), .B(n16758), .Z(n16757) );
  XOR U16472 ( .A(p_input[1877]), .B(n16756), .Z(n16758) );
  XNOR U16473 ( .A(n16759), .B(n16760), .Z(n16756) );
  AND U16474 ( .A(n1237), .B(n16761), .Z(n16760) );
  XOR U16475 ( .A(n16762), .B(n16763), .Z(n16754) );
  AND U16476 ( .A(n1241), .B(n16753), .Z(n16763) );
  XNOR U16477 ( .A(n16764), .B(n16751), .Z(n16753) );
  XOR U16478 ( .A(n16765), .B(n16766), .Z(n16751) );
  AND U16479 ( .A(n1264), .B(n16767), .Z(n16766) );
  IV U16480 ( .A(n16762), .Z(n16764) );
  XOR U16481 ( .A(n16768), .B(n16769), .Z(n16762) );
  AND U16482 ( .A(n1248), .B(n16761), .Z(n16769) );
  XNOR U16483 ( .A(n16759), .B(n16768), .Z(n16761) );
  XNOR U16484 ( .A(n16770), .B(n16771), .Z(n16759) );
  AND U16485 ( .A(n1252), .B(n16772), .Z(n16771) );
  XOR U16486 ( .A(p_input[1909]), .B(n16770), .Z(n16772) );
  XNOR U16487 ( .A(n16773), .B(n16774), .Z(n16770) );
  AND U16488 ( .A(n1256), .B(n16775), .Z(n16774) );
  XOR U16489 ( .A(n16776), .B(n16777), .Z(n16768) );
  AND U16490 ( .A(n1260), .B(n16767), .Z(n16777) );
  XNOR U16491 ( .A(n16778), .B(n16765), .Z(n16767) );
  XOR U16492 ( .A(n16779), .B(n16780), .Z(n16765) );
  AND U16493 ( .A(n1282), .B(n16781), .Z(n16780) );
  IV U16494 ( .A(n16776), .Z(n16778) );
  XOR U16495 ( .A(n16782), .B(n16783), .Z(n16776) );
  AND U16496 ( .A(n1267), .B(n16775), .Z(n16783) );
  XNOR U16497 ( .A(n16773), .B(n16782), .Z(n16775) );
  XNOR U16498 ( .A(n16784), .B(n16785), .Z(n16773) );
  AND U16499 ( .A(n1271), .B(n16786), .Z(n16785) );
  XOR U16500 ( .A(p_input[1941]), .B(n16784), .Z(n16786) );
  XOR U16501 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][21] ), .B(n16787), 
        .Z(n16784) );
  AND U16502 ( .A(n1274), .B(n16788), .Z(n16787) );
  XOR U16503 ( .A(n16789), .B(n16790), .Z(n16782) );
  AND U16504 ( .A(n1278), .B(n16781), .Z(n16790) );
  XNOR U16505 ( .A(n16791), .B(n16779), .Z(n16781) );
  XOR U16506 ( .A(\knn_comb_/min_val_out[0][21] ), .B(n16792), .Z(n16779) );
  AND U16507 ( .A(n1290), .B(n16793), .Z(n16792) );
  IV U16508 ( .A(n16789), .Z(n16791) );
  XOR U16509 ( .A(n16794), .B(n16795), .Z(n16789) );
  AND U16510 ( .A(n1285), .B(n16788), .Z(n16795) );
  XOR U16511 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][21] ), .B(n16794), 
        .Z(n16788) );
  XOR U16512 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .B(n16796), 
        .Z(n16794) );
  AND U16513 ( .A(n1287), .B(n16793), .Z(n16796) );
  XOR U16514 ( .A(\knn_comb_/min_val_out[0][21] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .Z(n16793) );
  XOR U16515 ( .A(n97), .B(n16797), .Z(o[20]) );
  AND U16516 ( .A(n122), .B(n16798), .Z(n97) );
  XOR U16517 ( .A(n98), .B(n16797), .Z(n16798) );
  XOR U16518 ( .A(n16799), .B(n16800), .Z(n16797) );
  AND U16519 ( .A(n142), .B(n16801), .Z(n16800) );
  XOR U16520 ( .A(n16802), .B(n27), .Z(n98) );
  AND U16521 ( .A(n125), .B(n16803), .Z(n27) );
  XOR U16522 ( .A(n28), .B(n16802), .Z(n16803) );
  XOR U16523 ( .A(n16804), .B(n16805), .Z(n28) );
  AND U16524 ( .A(n130), .B(n16806), .Z(n16805) );
  XOR U16525 ( .A(p_input[20]), .B(n16804), .Z(n16806) );
  XNOR U16526 ( .A(n16807), .B(n16808), .Z(n16804) );
  AND U16527 ( .A(n134), .B(n16809), .Z(n16808) );
  XOR U16528 ( .A(n16810), .B(n16811), .Z(n16802) );
  AND U16529 ( .A(n138), .B(n16801), .Z(n16811) );
  XNOR U16530 ( .A(n16812), .B(n16799), .Z(n16801) );
  XOR U16531 ( .A(n16813), .B(n16814), .Z(n16799) );
  AND U16532 ( .A(n162), .B(n16815), .Z(n16814) );
  IV U16533 ( .A(n16810), .Z(n16812) );
  XOR U16534 ( .A(n16816), .B(n16817), .Z(n16810) );
  AND U16535 ( .A(n146), .B(n16809), .Z(n16817) );
  XNOR U16536 ( .A(n16807), .B(n16816), .Z(n16809) );
  XNOR U16537 ( .A(n16818), .B(n16819), .Z(n16807) );
  AND U16538 ( .A(n150), .B(n16820), .Z(n16819) );
  XOR U16539 ( .A(p_input[52]), .B(n16818), .Z(n16820) );
  XNOR U16540 ( .A(n16821), .B(n16822), .Z(n16818) );
  AND U16541 ( .A(n154), .B(n16823), .Z(n16822) );
  XOR U16542 ( .A(n16824), .B(n16825), .Z(n16816) );
  AND U16543 ( .A(n158), .B(n16815), .Z(n16825) );
  XNOR U16544 ( .A(n16826), .B(n16813), .Z(n16815) );
  XOR U16545 ( .A(n16827), .B(n16828), .Z(n16813) );
  AND U16546 ( .A(n181), .B(n16829), .Z(n16828) );
  IV U16547 ( .A(n16824), .Z(n16826) );
  XOR U16548 ( .A(n16830), .B(n16831), .Z(n16824) );
  AND U16549 ( .A(n165), .B(n16823), .Z(n16831) );
  XNOR U16550 ( .A(n16821), .B(n16830), .Z(n16823) );
  XNOR U16551 ( .A(n16832), .B(n16833), .Z(n16821) );
  AND U16552 ( .A(n169), .B(n16834), .Z(n16833) );
  XOR U16553 ( .A(p_input[84]), .B(n16832), .Z(n16834) );
  XNOR U16554 ( .A(n16835), .B(n16836), .Z(n16832) );
  AND U16555 ( .A(n173), .B(n16837), .Z(n16836) );
  XOR U16556 ( .A(n16838), .B(n16839), .Z(n16830) );
  AND U16557 ( .A(n177), .B(n16829), .Z(n16839) );
  XNOR U16558 ( .A(n16840), .B(n16827), .Z(n16829) );
  XOR U16559 ( .A(n16841), .B(n16842), .Z(n16827) );
  AND U16560 ( .A(n200), .B(n16843), .Z(n16842) );
  IV U16561 ( .A(n16838), .Z(n16840) );
  XOR U16562 ( .A(n16844), .B(n16845), .Z(n16838) );
  AND U16563 ( .A(n184), .B(n16837), .Z(n16845) );
  XNOR U16564 ( .A(n16835), .B(n16844), .Z(n16837) );
  XNOR U16565 ( .A(n16846), .B(n16847), .Z(n16835) );
  AND U16566 ( .A(n188), .B(n16848), .Z(n16847) );
  XOR U16567 ( .A(p_input[116]), .B(n16846), .Z(n16848) );
  XNOR U16568 ( .A(n16849), .B(n16850), .Z(n16846) );
  AND U16569 ( .A(n192), .B(n16851), .Z(n16850) );
  XOR U16570 ( .A(n16852), .B(n16853), .Z(n16844) );
  AND U16571 ( .A(n196), .B(n16843), .Z(n16853) );
  XNOR U16572 ( .A(n16854), .B(n16841), .Z(n16843) );
  XOR U16573 ( .A(n16855), .B(n16856), .Z(n16841) );
  AND U16574 ( .A(n219), .B(n16857), .Z(n16856) );
  IV U16575 ( .A(n16852), .Z(n16854) );
  XOR U16576 ( .A(n16858), .B(n16859), .Z(n16852) );
  AND U16577 ( .A(n203), .B(n16851), .Z(n16859) );
  XNOR U16578 ( .A(n16849), .B(n16858), .Z(n16851) );
  XNOR U16579 ( .A(n16860), .B(n16861), .Z(n16849) );
  AND U16580 ( .A(n207), .B(n16862), .Z(n16861) );
  XOR U16581 ( .A(p_input[148]), .B(n16860), .Z(n16862) );
  XNOR U16582 ( .A(n16863), .B(n16864), .Z(n16860) );
  AND U16583 ( .A(n211), .B(n16865), .Z(n16864) );
  XOR U16584 ( .A(n16866), .B(n16867), .Z(n16858) );
  AND U16585 ( .A(n215), .B(n16857), .Z(n16867) );
  XNOR U16586 ( .A(n16868), .B(n16855), .Z(n16857) );
  XOR U16587 ( .A(n16869), .B(n16870), .Z(n16855) );
  AND U16588 ( .A(n238), .B(n16871), .Z(n16870) );
  IV U16589 ( .A(n16866), .Z(n16868) );
  XOR U16590 ( .A(n16872), .B(n16873), .Z(n16866) );
  AND U16591 ( .A(n222), .B(n16865), .Z(n16873) );
  XNOR U16592 ( .A(n16863), .B(n16872), .Z(n16865) );
  XNOR U16593 ( .A(n16874), .B(n16875), .Z(n16863) );
  AND U16594 ( .A(n226), .B(n16876), .Z(n16875) );
  XOR U16595 ( .A(p_input[180]), .B(n16874), .Z(n16876) );
  XNOR U16596 ( .A(n16877), .B(n16878), .Z(n16874) );
  AND U16597 ( .A(n230), .B(n16879), .Z(n16878) );
  XOR U16598 ( .A(n16880), .B(n16881), .Z(n16872) );
  AND U16599 ( .A(n234), .B(n16871), .Z(n16881) );
  XNOR U16600 ( .A(n16882), .B(n16869), .Z(n16871) );
  XOR U16601 ( .A(n16883), .B(n16884), .Z(n16869) );
  AND U16602 ( .A(n257), .B(n16885), .Z(n16884) );
  IV U16603 ( .A(n16880), .Z(n16882) );
  XOR U16604 ( .A(n16886), .B(n16887), .Z(n16880) );
  AND U16605 ( .A(n241), .B(n16879), .Z(n16887) );
  XNOR U16606 ( .A(n16877), .B(n16886), .Z(n16879) );
  XNOR U16607 ( .A(n16888), .B(n16889), .Z(n16877) );
  AND U16608 ( .A(n245), .B(n16890), .Z(n16889) );
  XOR U16609 ( .A(p_input[212]), .B(n16888), .Z(n16890) );
  XNOR U16610 ( .A(n16891), .B(n16892), .Z(n16888) );
  AND U16611 ( .A(n249), .B(n16893), .Z(n16892) );
  XOR U16612 ( .A(n16894), .B(n16895), .Z(n16886) );
  AND U16613 ( .A(n253), .B(n16885), .Z(n16895) );
  XNOR U16614 ( .A(n16896), .B(n16883), .Z(n16885) );
  XOR U16615 ( .A(n16897), .B(n16898), .Z(n16883) );
  AND U16616 ( .A(n276), .B(n16899), .Z(n16898) );
  IV U16617 ( .A(n16894), .Z(n16896) );
  XOR U16618 ( .A(n16900), .B(n16901), .Z(n16894) );
  AND U16619 ( .A(n260), .B(n16893), .Z(n16901) );
  XNOR U16620 ( .A(n16891), .B(n16900), .Z(n16893) );
  XNOR U16621 ( .A(n16902), .B(n16903), .Z(n16891) );
  AND U16622 ( .A(n264), .B(n16904), .Z(n16903) );
  XOR U16623 ( .A(p_input[244]), .B(n16902), .Z(n16904) );
  XNOR U16624 ( .A(n16905), .B(n16906), .Z(n16902) );
  AND U16625 ( .A(n268), .B(n16907), .Z(n16906) );
  XOR U16626 ( .A(n16908), .B(n16909), .Z(n16900) );
  AND U16627 ( .A(n272), .B(n16899), .Z(n16909) );
  XNOR U16628 ( .A(n16910), .B(n16897), .Z(n16899) );
  XOR U16629 ( .A(n16911), .B(n16912), .Z(n16897) );
  AND U16630 ( .A(n295), .B(n16913), .Z(n16912) );
  IV U16631 ( .A(n16908), .Z(n16910) );
  XOR U16632 ( .A(n16914), .B(n16915), .Z(n16908) );
  AND U16633 ( .A(n279), .B(n16907), .Z(n16915) );
  XNOR U16634 ( .A(n16905), .B(n16914), .Z(n16907) );
  XNOR U16635 ( .A(n16916), .B(n16917), .Z(n16905) );
  AND U16636 ( .A(n283), .B(n16918), .Z(n16917) );
  XOR U16637 ( .A(p_input[276]), .B(n16916), .Z(n16918) );
  XNOR U16638 ( .A(n16919), .B(n16920), .Z(n16916) );
  AND U16639 ( .A(n287), .B(n16921), .Z(n16920) );
  XOR U16640 ( .A(n16922), .B(n16923), .Z(n16914) );
  AND U16641 ( .A(n291), .B(n16913), .Z(n16923) );
  XNOR U16642 ( .A(n16924), .B(n16911), .Z(n16913) );
  XOR U16643 ( .A(n16925), .B(n16926), .Z(n16911) );
  AND U16644 ( .A(n314), .B(n16927), .Z(n16926) );
  IV U16645 ( .A(n16922), .Z(n16924) );
  XOR U16646 ( .A(n16928), .B(n16929), .Z(n16922) );
  AND U16647 ( .A(n298), .B(n16921), .Z(n16929) );
  XNOR U16648 ( .A(n16919), .B(n16928), .Z(n16921) );
  XNOR U16649 ( .A(n16930), .B(n16931), .Z(n16919) );
  AND U16650 ( .A(n302), .B(n16932), .Z(n16931) );
  XOR U16651 ( .A(p_input[308]), .B(n16930), .Z(n16932) );
  XNOR U16652 ( .A(n16933), .B(n16934), .Z(n16930) );
  AND U16653 ( .A(n306), .B(n16935), .Z(n16934) );
  XOR U16654 ( .A(n16936), .B(n16937), .Z(n16928) );
  AND U16655 ( .A(n310), .B(n16927), .Z(n16937) );
  XNOR U16656 ( .A(n16938), .B(n16925), .Z(n16927) );
  XOR U16657 ( .A(n16939), .B(n16940), .Z(n16925) );
  AND U16658 ( .A(n333), .B(n16941), .Z(n16940) );
  IV U16659 ( .A(n16936), .Z(n16938) );
  XOR U16660 ( .A(n16942), .B(n16943), .Z(n16936) );
  AND U16661 ( .A(n317), .B(n16935), .Z(n16943) );
  XNOR U16662 ( .A(n16933), .B(n16942), .Z(n16935) );
  XNOR U16663 ( .A(n16944), .B(n16945), .Z(n16933) );
  AND U16664 ( .A(n321), .B(n16946), .Z(n16945) );
  XOR U16665 ( .A(p_input[340]), .B(n16944), .Z(n16946) );
  XNOR U16666 ( .A(n16947), .B(n16948), .Z(n16944) );
  AND U16667 ( .A(n325), .B(n16949), .Z(n16948) );
  XOR U16668 ( .A(n16950), .B(n16951), .Z(n16942) );
  AND U16669 ( .A(n329), .B(n16941), .Z(n16951) );
  XNOR U16670 ( .A(n16952), .B(n16939), .Z(n16941) );
  XOR U16671 ( .A(n16953), .B(n16954), .Z(n16939) );
  AND U16672 ( .A(n352), .B(n16955), .Z(n16954) );
  IV U16673 ( .A(n16950), .Z(n16952) );
  XOR U16674 ( .A(n16956), .B(n16957), .Z(n16950) );
  AND U16675 ( .A(n336), .B(n16949), .Z(n16957) );
  XNOR U16676 ( .A(n16947), .B(n16956), .Z(n16949) );
  XNOR U16677 ( .A(n16958), .B(n16959), .Z(n16947) );
  AND U16678 ( .A(n340), .B(n16960), .Z(n16959) );
  XOR U16679 ( .A(p_input[372]), .B(n16958), .Z(n16960) );
  XNOR U16680 ( .A(n16961), .B(n16962), .Z(n16958) );
  AND U16681 ( .A(n344), .B(n16963), .Z(n16962) );
  XOR U16682 ( .A(n16964), .B(n16965), .Z(n16956) );
  AND U16683 ( .A(n348), .B(n16955), .Z(n16965) );
  XNOR U16684 ( .A(n16966), .B(n16953), .Z(n16955) );
  XOR U16685 ( .A(n16967), .B(n16968), .Z(n16953) );
  AND U16686 ( .A(n371), .B(n16969), .Z(n16968) );
  IV U16687 ( .A(n16964), .Z(n16966) );
  XOR U16688 ( .A(n16970), .B(n16971), .Z(n16964) );
  AND U16689 ( .A(n355), .B(n16963), .Z(n16971) );
  XNOR U16690 ( .A(n16961), .B(n16970), .Z(n16963) );
  XNOR U16691 ( .A(n16972), .B(n16973), .Z(n16961) );
  AND U16692 ( .A(n359), .B(n16974), .Z(n16973) );
  XOR U16693 ( .A(p_input[404]), .B(n16972), .Z(n16974) );
  XNOR U16694 ( .A(n16975), .B(n16976), .Z(n16972) );
  AND U16695 ( .A(n363), .B(n16977), .Z(n16976) );
  XOR U16696 ( .A(n16978), .B(n16979), .Z(n16970) );
  AND U16697 ( .A(n367), .B(n16969), .Z(n16979) );
  XNOR U16698 ( .A(n16980), .B(n16967), .Z(n16969) );
  XOR U16699 ( .A(n16981), .B(n16982), .Z(n16967) );
  AND U16700 ( .A(n390), .B(n16983), .Z(n16982) );
  IV U16701 ( .A(n16978), .Z(n16980) );
  XOR U16702 ( .A(n16984), .B(n16985), .Z(n16978) );
  AND U16703 ( .A(n374), .B(n16977), .Z(n16985) );
  XNOR U16704 ( .A(n16975), .B(n16984), .Z(n16977) );
  XNOR U16705 ( .A(n16986), .B(n16987), .Z(n16975) );
  AND U16706 ( .A(n378), .B(n16988), .Z(n16987) );
  XOR U16707 ( .A(p_input[436]), .B(n16986), .Z(n16988) );
  XNOR U16708 ( .A(n16989), .B(n16990), .Z(n16986) );
  AND U16709 ( .A(n382), .B(n16991), .Z(n16990) );
  XOR U16710 ( .A(n16992), .B(n16993), .Z(n16984) );
  AND U16711 ( .A(n386), .B(n16983), .Z(n16993) );
  XNOR U16712 ( .A(n16994), .B(n16981), .Z(n16983) );
  XOR U16713 ( .A(n16995), .B(n16996), .Z(n16981) );
  AND U16714 ( .A(n409), .B(n16997), .Z(n16996) );
  IV U16715 ( .A(n16992), .Z(n16994) );
  XOR U16716 ( .A(n16998), .B(n16999), .Z(n16992) );
  AND U16717 ( .A(n393), .B(n16991), .Z(n16999) );
  XNOR U16718 ( .A(n16989), .B(n16998), .Z(n16991) );
  XNOR U16719 ( .A(n17000), .B(n17001), .Z(n16989) );
  AND U16720 ( .A(n397), .B(n17002), .Z(n17001) );
  XOR U16721 ( .A(p_input[468]), .B(n17000), .Z(n17002) );
  XNOR U16722 ( .A(n17003), .B(n17004), .Z(n17000) );
  AND U16723 ( .A(n401), .B(n17005), .Z(n17004) );
  XOR U16724 ( .A(n17006), .B(n17007), .Z(n16998) );
  AND U16725 ( .A(n405), .B(n16997), .Z(n17007) );
  XNOR U16726 ( .A(n17008), .B(n16995), .Z(n16997) );
  XOR U16727 ( .A(n17009), .B(n17010), .Z(n16995) );
  AND U16728 ( .A(n428), .B(n17011), .Z(n17010) );
  IV U16729 ( .A(n17006), .Z(n17008) );
  XOR U16730 ( .A(n17012), .B(n17013), .Z(n17006) );
  AND U16731 ( .A(n412), .B(n17005), .Z(n17013) );
  XNOR U16732 ( .A(n17003), .B(n17012), .Z(n17005) );
  XNOR U16733 ( .A(n17014), .B(n17015), .Z(n17003) );
  AND U16734 ( .A(n416), .B(n17016), .Z(n17015) );
  XOR U16735 ( .A(p_input[500]), .B(n17014), .Z(n17016) );
  XNOR U16736 ( .A(n17017), .B(n17018), .Z(n17014) );
  AND U16737 ( .A(n420), .B(n17019), .Z(n17018) );
  XOR U16738 ( .A(n17020), .B(n17021), .Z(n17012) );
  AND U16739 ( .A(n424), .B(n17011), .Z(n17021) );
  XNOR U16740 ( .A(n17022), .B(n17009), .Z(n17011) );
  XOR U16741 ( .A(n17023), .B(n17024), .Z(n17009) );
  AND U16742 ( .A(n447), .B(n17025), .Z(n17024) );
  IV U16743 ( .A(n17020), .Z(n17022) );
  XOR U16744 ( .A(n17026), .B(n17027), .Z(n17020) );
  AND U16745 ( .A(n431), .B(n17019), .Z(n17027) );
  XNOR U16746 ( .A(n17017), .B(n17026), .Z(n17019) );
  XNOR U16747 ( .A(n17028), .B(n17029), .Z(n17017) );
  AND U16748 ( .A(n435), .B(n17030), .Z(n17029) );
  XOR U16749 ( .A(p_input[532]), .B(n17028), .Z(n17030) );
  XNOR U16750 ( .A(n17031), .B(n17032), .Z(n17028) );
  AND U16751 ( .A(n439), .B(n17033), .Z(n17032) );
  XOR U16752 ( .A(n17034), .B(n17035), .Z(n17026) );
  AND U16753 ( .A(n443), .B(n17025), .Z(n17035) );
  XNOR U16754 ( .A(n17036), .B(n17023), .Z(n17025) );
  XOR U16755 ( .A(n17037), .B(n17038), .Z(n17023) );
  AND U16756 ( .A(n466), .B(n17039), .Z(n17038) );
  IV U16757 ( .A(n17034), .Z(n17036) );
  XOR U16758 ( .A(n17040), .B(n17041), .Z(n17034) );
  AND U16759 ( .A(n450), .B(n17033), .Z(n17041) );
  XNOR U16760 ( .A(n17031), .B(n17040), .Z(n17033) );
  XNOR U16761 ( .A(n17042), .B(n17043), .Z(n17031) );
  AND U16762 ( .A(n454), .B(n17044), .Z(n17043) );
  XOR U16763 ( .A(p_input[564]), .B(n17042), .Z(n17044) );
  XNOR U16764 ( .A(n17045), .B(n17046), .Z(n17042) );
  AND U16765 ( .A(n458), .B(n17047), .Z(n17046) );
  XOR U16766 ( .A(n17048), .B(n17049), .Z(n17040) );
  AND U16767 ( .A(n462), .B(n17039), .Z(n17049) );
  XNOR U16768 ( .A(n17050), .B(n17037), .Z(n17039) );
  XOR U16769 ( .A(n17051), .B(n17052), .Z(n17037) );
  AND U16770 ( .A(n485), .B(n17053), .Z(n17052) );
  IV U16771 ( .A(n17048), .Z(n17050) );
  XOR U16772 ( .A(n17054), .B(n17055), .Z(n17048) );
  AND U16773 ( .A(n469), .B(n17047), .Z(n17055) );
  XNOR U16774 ( .A(n17045), .B(n17054), .Z(n17047) );
  XNOR U16775 ( .A(n17056), .B(n17057), .Z(n17045) );
  AND U16776 ( .A(n473), .B(n17058), .Z(n17057) );
  XOR U16777 ( .A(p_input[596]), .B(n17056), .Z(n17058) );
  XNOR U16778 ( .A(n17059), .B(n17060), .Z(n17056) );
  AND U16779 ( .A(n477), .B(n17061), .Z(n17060) );
  XOR U16780 ( .A(n17062), .B(n17063), .Z(n17054) );
  AND U16781 ( .A(n481), .B(n17053), .Z(n17063) );
  XNOR U16782 ( .A(n17064), .B(n17051), .Z(n17053) );
  XOR U16783 ( .A(n17065), .B(n17066), .Z(n17051) );
  AND U16784 ( .A(n504), .B(n17067), .Z(n17066) );
  IV U16785 ( .A(n17062), .Z(n17064) );
  XOR U16786 ( .A(n17068), .B(n17069), .Z(n17062) );
  AND U16787 ( .A(n488), .B(n17061), .Z(n17069) );
  XNOR U16788 ( .A(n17059), .B(n17068), .Z(n17061) );
  XNOR U16789 ( .A(n17070), .B(n17071), .Z(n17059) );
  AND U16790 ( .A(n492), .B(n17072), .Z(n17071) );
  XOR U16791 ( .A(p_input[628]), .B(n17070), .Z(n17072) );
  XNOR U16792 ( .A(n17073), .B(n17074), .Z(n17070) );
  AND U16793 ( .A(n496), .B(n17075), .Z(n17074) );
  XOR U16794 ( .A(n17076), .B(n17077), .Z(n17068) );
  AND U16795 ( .A(n500), .B(n17067), .Z(n17077) );
  XNOR U16796 ( .A(n17078), .B(n17065), .Z(n17067) );
  XOR U16797 ( .A(n17079), .B(n17080), .Z(n17065) );
  AND U16798 ( .A(n523), .B(n17081), .Z(n17080) );
  IV U16799 ( .A(n17076), .Z(n17078) );
  XOR U16800 ( .A(n17082), .B(n17083), .Z(n17076) );
  AND U16801 ( .A(n507), .B(n17075), .Z(n17083) );
  XNOR U16802 ( .A(n17073), .B(n17082), .Z(n17075) );
  XNOR U16803 ( .A(n17084), .B(n17085), .Z(n17073) );
  AND U16804 ( .A(n511), .B(n17086), .Z(n17085) );
  XOR U16805 ( .A(p_input[660]), .B(n17084), .Z(n17086) );
  XNOR U16806 ( .A(n17087), .B(n17088), .Z(n17084) );
  AND U16807 ( .A(n515), .B(n17089), .Z(n17088) );
  XOR U16808 ( .A(n17090), .B(n17091), .Z(n17082) );
  AND U16809 ( .A(n519), .B(n17081), .Z(n17091) );
  XNOR U16810 ( .A(n17092), .B(n17079), .Z(n17081) );
  XOR U16811 ( .A(n17093), .B(n17094), .Z(n17079) );
  AND U16812 ( .A(n542), .B(n17095), .Z(n17094) );
  IV U16813 ( .A(n17090), .Z(n17092) );
  XOR U16814 ( .A(n17096), .B(n17097), .Z(n17090) );
  AND U16815 ( .A(n526), .B(n17089), .Z(n17097) );
  XNOR U16816 ( .A(n17087), .B(n17096), .Z(n17089) );
  XNOR U16817 ( .A(n17098), .B(n17099), .Z(n17087) );
  AND U16818 ( .A(n530), .B(n17100), .Z(n17099) );
  XOR U16819 ( .A(p_input[692]), .B(n17098), .Z(n17100) );
  XNOR U16820 ( .A(n17101), .B(n17102), .Z(n17098) );
  AND U16821 ( .A(n534), .B(n17103), .Z(n17102) );
  XOR U16822 ( .A(n17104), .B(n17105), .Z(n17096) );
  AND U16823 ( .A(n538), .B(n17095), .Z(n17105) );
  XNOR U16824 ( .A(n17106), .B(n17093), .Z(n17095) );
  XOR U16825 ( .A(n17107), .B(n17108), .Z(n17093) );
  AND U16826 ( .A(n561), .B(n17109), .Z(n17108) );
  IV U16827 ( .A(n17104), .Z(n17106) );
  XOR U16828 ( .A(n17110), .B(n17111), .Z(n17104) );
  AND U16829 ( .A(n545), .B(n17103), .Z(n17111) );
  XNOR U16830 ( .A(n17101), .B(n17110), .Z(n17103) );
  XNOR U16831 ( .A(n17112), .B(n17113), .Z(n17101) );
  AND U16832 ( .A(n549), .B(n17114), .Z(n17113) );
  XOR U16833 ( .A(p_input[724]), .B(n17112), .Z(n17114) );
  XNOR U16834 ( .A(n17115), .B(n17116), .Z(n17112) );
  AND U16835 ( .A(n553), .B(n17117), .Z(n17116) );
  XOR U16836 ( .A(n17118), .B(n17119), .Z(n17110) );
  AND U16837 ( .A(n557), .B(n17109), .Z(n17119) );
  XNOR U16838 ( .A(n17120), .B(n17107), .Z(n17109) );
  XOR U16839 ( .A(n17121), .B(n17122), .Z(n17107) );
  AND U16840 ( .A(n580), .B(n17123), .Z(n17122) );
  IV U16841 ( .A(n17118), .Z(n17120) );
  XOR U16842 ( .A(n17124), .B(n17125), .Z(n17118) );
  AND U16843 ( .A(n564), .B(n17117), .Z(n17125) );
  XNOR U16844 ( .A(n17115), .B(n17124), .Z(n17117) );
  XNOR U16845 ( .A(n17126), .B(n17127), .Z(n17115) );
  AND U16846 ( .A(n568), .B(n17128), .Z(n17127) );
  XOR U16847 ( .A(p_input[756]), .B(n17126), .Z(n17128) );
  XNOR U16848 ( .A(n17129), .B(n17130), .Z(n17126) );
  AND U16849 ( .A(n572), .B(n17131), .Z(n17130) );
  XOR U16850 ( .A(n17132), .B(n17133), .Z(n17124) );
  AND U16851 ( .A(n576), .B(n17123), .Z(n17133) );
  XNOR U16852 ( .A(n17134), .B(n17121), .Z(n17123) );
  XOR U16853 ( .A(n17135), .B(n17136), .Z(n17121) );
  AND U16854 ( .A(n599), .B(n17137), .Z(n17136) );
  IV U16855 ( .A(n17132), .Z(n17134) );
  XOR U16856 ( .A(n17138), .B(n17139), .Z(n17132) );
  AND U16857 ( .A(n583), .B(n17131), .Z(n17139) );
  XNOR U16858 ( .A(n17129), .B(n17138), .Z(n17131) );
  XNOR U16859 ( .A(n17140), .B(n17141), .Z(n17129) );
  AND U16860 ( .A(n587), .B(n17142), .Z(n17141) );
  XOR U16861 ( .A(p_input[788]), .B(n17140), .Z(n17142) );
  XNOR U16862 ( .A(n17143), .B(n17144), .Z(n17140) );
  AND U16863 ( .A(n591), .B(n17145), .Z(n17144) );
  XOR U16864 ( .A(n17146), .B(n17147), .Z(n17138) );
  AND U16865 ( .A(n595), .B(n17137), .Z(n17147) );
  XNOR U16866 ( .A(n17148), .B(n17135), .Z(n17137) );
  XOR U16867 ( .A(n17149), .B(n17150), .Z(n17135) );
  AND U16868 ( .A(n618), .B(n17151), .Z(n17150) );
  IV U16869 ( .A(n17146), .Z(n17148) );
  XOR U16870 ( .A(n17152), .B(n17153), .Z(n17146) );
  AND U16871 ( .A(n602), .B(n17145), .Z(n17153) );
  XNOR U16872 ( .A(n17143), .B(n17152), .Z(n17145) );
  XNOR U16873 ( .A(n17154), .B(n17155), .Z(n17143) );
  AND U16874 ( .A(n606), .B(n17156), .Z(n17155) );
  XOR U16875 ( .A(p_input[820]), .B(n17154), .Z(n17156) );
  XNOR U16876 ( .A(n17157), .B(n17158), .Z(n17154) );
  AND U16877 ( .A(n610), .B(n17159), .Z(n17158) );
  XOR U16878 ( .A(n17160), .B(n17161), .Z(n17152) );
  AND U16879 ( .A(n614), .B(n17151), .Z(n17161) );
  XNOR U16880 ( .A(n17162), .B(n17149), .Z(n17151) );
  XOR U16881 ( .A(n17163), .B(n17164), .Z(n17149) );
  AND U16882 ( .A(n637), .B(n17165), .Z(n17164) );
  IV U16883 ( .A(n17160), .Z(n17162) );
  XOR U16884 ( .A(n17166), .B(n17167), .Z(n17160) );
  AND U16885 ( .A(n621), .B(n17159), .Z(n17167) );
  XNOR U16886 ( .A(n17157), .B(n17166), .Z(n17159) );
  XNOR U16887 ( .A(n17168), .B(n17169), .Z(n17157) );
  AND U16888 ( .A(n625), .B(n17170), .Z(n17169) );
  XOR U16889 ( .A(p_input[852]), .B(n17168), .Z(n17170) );
  XNOR U16890 ( .A(n17171), .B(n17172), .Z(n17168) );
  AND U16891 ( .A(n629), .B(n17173), .Z(n17172) );
  XOR U16892 ( .A(n17174), .B(n17175), .Z(n17166) );
  AND U16893 ( .A(n633), .B(n17165), .Z(n17175) );
  XNOR U16894 ( .A(n17176), .B(n17163), .Z(n17165) );
  XOR U16895 ( .A(n17177), .B(n17178), .Z(n17163) );
  AND U16896 ( .A(n656), .B(n17179), .Z(n17178) );
  IV U16897 ( .A(n17174), .Z(n17176) );
  XOR U16898 ( .A(n17180), .B(n17181), .Z(n17174) );
  AND U16899 ( .A(n640), .B(n17173), .Z(n17181) );
  XNOR U16900 ( .A(n17171), .B(n17180), .Z(n17173) );
  XNOR U16901 ( .A(n17182), .B(n17183), .Z(n17171) );
  AND U16902 ( .A(n644), .B(n17184), .Z(n17183) );
  XOR U16903 ( .A(p_input[884]), .B(n17182), .Z(n17184) );
  XNOR U16904 ( .A(n17185), .B(n17186), .Z(n17182) );
  AND U16905 ( .A(n648), .B(n17187), .Z(n17186) );
  XOR U16906 ( .A(n17188), .B(n17189), .Z(n17180) );
  AND U16907 ( .A(n652), .B(n17179), .Z(n17189) );
  XNOR U16908 ( .A(n17190), .B(n17177), .Z(n17179) );
  XOR U16909 ( .A(n17191), .B(n17192), .Z(n17177) );
  AND U16910 ( .A(n675), .B(n17193), .Z(n17192) );
  IV U16911 ( .A(n17188), .Z(n17190) );
  XOR U16912 ( .A(n17194), .B(n17195), .Z(n17188) );
  AND U16913 ( .A(n659), .B(n17187), .Z(n17195) );
  XNOR U16914 ( .A(n17185), .B(n17194), .Z(n17187) );
  XNOR U16915 ( .A(n17196), .B(n17197), .Z(n17185) );
  AND U16916 ( .A(n663), .B(n17198), .Z(n17197) );
  XOR U16917 ( .A(p_input[916]), .B(n17196), .Z(n17198) );
  XNOR U16918 ( .A(n17199), .B(n17200), .Z(n17196) );
  AND U16919 ( .A(n667), .B(n17201), .Z(n17200) );
  XOR U16920 ( .A(n17202), .B(n17203), .Z(n17194) );
  AND U16921 ( .A(n671), .B(n17193), .Z(n17203) );
  XNOR U16922 ( .A(n17204), .B(n17191), .Z(n17193) );
  XOR U16923 ( .A(n17205), .B(n17206), .Z(n17191) );
  AND U16924 ( .A(n694), .B(n17207), .Z(n17206) );
  IV U16925 ( .A(n17202), .Z(n17204) );
  XOR U16926 ( .A(n17208), .B(n17209), .Z(n17202) );
  AND U16927 ( .A(n678), .B(n17201), .Z(n17209) );
  XNOR U16928 ( .A(n17199), .B(n17208), .Z(n17201) );
  XNOR U16929 ( .A(n17210), .B(n17211), .Z(n17199) );
  AND U16930 ( .A(n682), .B(n17212), .Z(n17211) );
  XOR U16931 ( .A(p_input[948]), .B(n17210), .Z(n17212) );
  XNOR U16932 ( .A(n17213), .B(n17214), .Z(n17210) );
  AND U16933 ( .A(n686), .B(n17215), .Z(n17214) );
  XOR U16934 ( .A(n17216), .B(n17217), .Z(n17208) );
  AND U16935 ( .A(n690), .B(n17207), .Z(n17217) );
  XNOR U16936 ( .A(n17218), .B(n17205), .Z(n17207) );
  XOR U16937 ( .A(n17219), .B(n17220), .Z(n17205) );
  AND U16938 ( .A(n713), .B(n17221), .Z(n17220) );
  IV U16939 ( .A(n17216), .Z(n17218) );
  XOR U16940 ( .A(n17222), .B(n17223), .Z(n17216) );
  AND U16941 ( .A(n697), .B(n17215), .Z(n17223) );
  XNOR U16942 ( .A(n17213), .B(n17222), .Z(n17215) );
  XNOR U16943 ( .A(n17224), .B(n17225), .Z(n17213) );
  AND U16944 ( .A(n701), .B(n17226), .Z(n17225) );
  XOR U16945 ( .A(p_input[980]), .B(n17224), .Z(n17226) );
  XNOR U16946 ( .A(n17227), .B(n17228), .Z(n17224) );
  AND U16947 ( .A(n705), .B(n17229), .Z(n17228) );
  XOR U16948 ( .A(n17230), .B(n17231), .Z(n17222) );
  AND U16949 ( .A(n709), .B(n17221), .Z(n17231) );
  XNOR U16950 ( .A(n17232), .B(n17219), .Z(n17221) );
  XOR U16951 ( .A(n17233), .B(n17234), .Z(n17219) );
  AND U16952 ( .A(n732), .B(n17235), .Z(n17234) );
  IV U16953 ( .A(n17230), .Z(n17232) );
  XOR U16954 ( .A(n17236), .B(n17237), .Z(n17230) );
  AND U16955 ( .A(n716), .B(n17229), .Z(n17237) );
  XNOR U16956 ( .A(n17227), .B(n17236), .Z(n17229) );
  XNOR U16957 ( .A(n17238), .B(n17239), .Z(n17227) );
  AND U16958 ( .A(n720), .B(n17240), .Z(n17239) );
  XOR U16959 ( .A(p_input[1012]), .B(n17238), .Z(n17240) );
  XNOR U16960 ( .A(n17241), .B(n17242), .Z(n17238) );
  AND U16961 ( .A(n724), .B(n17243), .Z(n17242) );
  XOR U16962 ( .A(n17244), .B(n17245), .Z(n17236) );
  AND U16963 ( .A(n728), .B(n17235), .Z(n17245) );
  XNOR U16964 ( .A(n17246), .B(n17233), .Z(n17235) );
  XOR U16965 ( .A(n17247), .B(n17248), .Z(n17233) );
  AND U16966 ( .A(n751), .B(n17249), .Z(n17248) );
  IV U16967 ( .A(n17244), .Z(n17246) );
  XOR U16968 ( .A(n17250), .B(n17251), .Z(n17244) );
  AND U16969 ( .A(n735), .B(n17243), .Z(n17251) );
  XNOR U16970 ( .A(n17241), .B(n17250), .Z(n17243) );
  XNOR U16971 ( .A(n17252), .B(n17253), .Z(n17241) );
  AND U16972 ( .A(n739), .B(n17254), .Z(n17253) );
  XOR U16973 ( .A(p_input[1044]), .B(n17252), .Z(n17254) );
  XNOR U16974 ( .A(n17255), .B(n17256), .Z(n17252) );
  AND U16975 ( .A(n743), .B(n17257), .Z(n17256) );
  XOR U16976 ( .A(n17258), .B(n17259), .Z(n17250) );
  AND U16977 ( .A(n747), .B(n17249), .Z(n17259) );
  XNOR U16978 ( .A(n17260), .B(n17247), .Z(n17249) );
  XOR U16979 ( .A(n17261), .B(n17262), .Z(n17247) );
  AND U16980 ( .A(n770), .B(n17263), .Z(n17262) );
  IV U16981 ( .A(n17258), .Z(n17260) );
  XOR U16982 ( .A(n17264), .B(n17265), .Z(n17258) );
  AND U16983 ( .A(n754), .B(n17257), .Z(n17265) );
  XNOR U16984 ( .A(n17255), .B(n17264), .Z(n17257) );
  XNOR U16985 ( .A(n17266), .B(n17267), .Z(n17255) );
  AND U16986 ( .A(n758), .B(n17268), .Z(n17267) );
  XOR U16987 ( .A(p_input[1076]), .B(n17266), .Z(n17268) );
  XNOR U16988 ( .A(n17269), .B(n17270), .Z(n17266) );
  AND U16989 ( .A(n762), .B(n17271), .Z(n17270) );
  XOR U16990 ( .A(n17272), .B(n17273), .Z(n17264) );
  AND U16991 ( .A(n766), .B(n17263), .Z(n17273) );
  XNOR U16992 ( .A(n17274), .B(n17261), .Z(n17263) );
  XOR U16993 ( .A(n17275), .B(n17276), .Z(n17261) );
  AND U16994 ( .A(n789), .B(n17277), .Z(n17276) );
  IV U16995 ( .A(n17272), .Z(n17274) );
  XOR U16996 ( .A(n17278), .B(n17279), .Z(n17272) );
  AND U16997 ( .A(n773), .B(n17271), .Z(n17279) );
  XNOR U16998 ( .A(n17269), .B(n17278), .Z(n17271) );
  XNOR U16999 ( .A(n17280), .B(n17281), .Z(n17269) );
  AND U17000 ( .A(n777), .B(n17282), .Z(n17281) );
  XOR U17001 ( .A(p_input[1108]), .B(n17280), .Z(n17282) );
  XNOR U17002 ( .A(n17283), .B(n17284), .Z(n17280) );
  AND U17003 ( .A(n781), .B(n17285), .Z(n17284) );
  XOR U17004 ( .A(n17286), .B(n17287), .Z(n17278) );
  AND U17005 ( .A(n785), .B(n17277), .Z(n17287) );
  XNOR U17006 ( .A(n17288), .B(n17275), .Z(n17277) );
  XOR U17007 ( .A(n17289), .B(n17290), .Z(n17275) );
  AND U17008 ( .A(n808), .B(n17291), .Z(n17290) );
  IV U17009 ( .A(n17286), .Z(n17288) );
  XOR U17010 ( .A(n17292), .B(n17293), .Z(n17286) );
  AND U17011 ( .A(n792), .B(n17285), .Z(n17293) );
  XNOR U17012 ( .A(n17283), .B(n17292), .Z(n17285) );
  XNOR U17013 ( .A(n17294), .B(n17295), .Z(n17283) );
  AND U17014 ( .A(n796), .B(n17296), .Z(n17295) );
  XOR U17015 ( .A(p_input[1140]), .B(n17294), .Z(n17296) );
  XNOR U17016 ( .A(n17297), .B(n17298), .Z(n17294) );
  AND U17017 ( .A(n800), .B(n17299), .Z(n17298) );
  XOR U17018 ( .A(n17300), .B(n17301), .Z(n17292) );
  AND U17019 ( .A(n804), .B(n17291), .Z(n17301) );
  XNOR U17020 ( .A(n17302), .B(n17289), .Z(n17291) );
  XOR U17021 ( .A(n17303), .B(n17304), .Z(n17289) );
  AND U17022 ( .A(n827), .B(n17305), .Z(n17304) );
  IV U17023 ( .A(n17300), .Z(n17302) );
  XOR U17024 ( .A(n17306), .B(n17307), .Z(n17300) );
  AND U17025 ( .A(n811), .B(n17299), .Z(n17307) );
  XNOR U17026 ( .A(n17297), .B(n17306), .Z(n17299) );
  XNOR U17027 ( .A(n17308), .B(n17309), .Z(n17297) );
  AND U17028 ( .A(n815), .B(n17310), .Z(n17309) );
  XOR U17029 ( .A(p_input[1172]), .B(n17308), .Z(n17310) );
  XNOR U17030 ( .A(n17311), .B(n17312), .Z(n17308) );
  AND U17031 ( .A(n819), .B(n17313), .Z(n17312) );
  XOR U17032 ( .A(n17314), .B(n17315), .Z(n17306) );
  AND U17033 ( .A(n823), .B(n17305), .Z(n17315) );
  XNOR U17034 ( .A(n17316), .B(n17303), .Z(n17305) );
  XOR U17035 ( .A(n17317), .B(n17318), .Z(n17303) );
  AND U17036 ( .A(n846), .B(n17319), .Z(n17318) );
  IV U17037 ( .A(n17314), .Z(n17316) );
  XOR U17038 ( .A(n17320), .B(n17321), .Z(n17314) );
  AND U17039 ( .A(n830), .B(n17313), .Z(n17321) );
  XNOR U17040 ( .A(n17311), .B(n17320), .Z(n17313) );
  XNOR U17041 ( .A(n17322), .B(n17323), .Z(n17311) );
  AND U17042 ( .A(n834), .B(n17324), .Z(n17323) );
  XOR U17043 ( .A(p_input[1204]), .B(n17322), .Z(n17324) );
  XNOR U17044 ( .A(n17325), .B(n17326), .Z(n17322) );
  AND U17045 ( .A(n838), .B(n17327), .Z(n17326) );
  XOR U17046 ( .A(n17328), .B(n17329), .Z(n17320) );
  AND U17047 ( .A(n842), .B(n17319), .Z(n17329) );
  XNOR U17048 ( .A(n17330), .B(n17317), .Z(n17319) );
  XOR U17049 ( .A(n17331), .B(n17332), .Z(n17317) );
  AND U17050 ( .A(n865), .B(n17333), .Z(n17332) );
  IV U17051 ( .A(n17328), .Z(n17330) );
  XOR U17052 ( .A(n17334), .B(n17335), .Z(n17328) );
  AND U17053 ( .A(n849), .B(n17327), .Z(n17335) );
  XNOR U17054 ( .A(n17325), .B(n17334), .Z(n17327) );
  XNOR U17055 ( .A(n17336), .B(n17337), .Z(n17325) );
  AND U17056 ( .A(n853), .B(n17338), .Z(n17337) );
  XOR U17057 ( .A(p_input[1236]), .B(n17336), .Z(n17338) );
  XNOR U17058 ( .A(n17339), .B(n17340), .Z(n17336) );
  AND U17059 ( .A(n857), .B(n17341), .Z(n17340) );
  XOR U17060 ( .A(n17342), .B(n17343), .Z(n17334) );
  AND U17061 ( .A(n861), .B(n17333), .Z(n17343) );
  XNOR U17062 ( .A(n17344), .B(n17331), .Z(n17333) );
  XOR U17063 ( .A(n17345), .B(n17346), .Z(n17331) );
  AND U17064 ( .A(n884), .B(n17347), .Z(n17346) );
  IV U17065 ( .A(n17342), .Z(n17344) );
  XOR U17066 ( .A(n17348), .B(n17349), .Z(n17342) );
  AND U17067 ( .A(n868), .B(n17341), .Z(n17349) );
  XNOR U17068 ( .A(n17339), .B(n17348), .Z(n17341) );
  XNOR U17069 ( .A(n17350), .B(n17351), .Z(n17339) );
  AND U17070 ( .A(n872), .B(n17352), .Z(n17351) );
  XOR U17071 ( .A(p_input[1268]), .B(n17350), .Z(n17352) );
  XNOR U17072 ( .A(n17353), .B(n17354), .Z(n17350) );
  AND U17073 ( .A(n876), .B(n17355), .Z(n17354) );
  XOR U17074 ( .A(n17356), .B(n17357), .Z(n17348) );
  AND U17075 ( .A(n880), .B(n17347), .Z(n17357) );
  XNOR U17076 ( .A(n17358), .B(n17345), .Z(n17347) );
  XOR U17077 ( .A(n17359), .B(n17360), .Z(n17345) );
  AND U17078 ( .A(n903), .B(n17361), .Z(n17360) );
  IV U17079 ( .A(n17356), .Z(n17358) );
  XOR U17080 ( .A(n17362), .B(n17363), .Z(n17356) );
  AND U17081 ( .A(n887), .B(n17355), .Z(n17363) );
  XNOR U17082 ( .A(n17353), .B(n17362), .Z(n17355) );
  XNOR U17083 ( .A(n17364), .B(n17365), .Z(n17353) );
  AND U17084 ( .A(n891), .B(n17366), .Z(n17365) );
  XOR U17085 ( .A(p_input[1300]), .B(n17364), .Z(n17366) );
  XNOR U17086 ( .A(n17367), .B(n17368), .Z(n17364) );
  AND U17087 ( .A(n895), .B(n17369), .Z(n17368) );
  XOR U17088 ( .A(n17370), .B(n17371), .Z(n17362) );
  AND U17089 ( .A(n899), .B(n17361), .Z(n17371) );
  XNOR U17090 ( .A(n17372), .B(n17359), .Z(n17361) );
  XOR U17091 ( .A(n17373), .B(n17374), .Z(n17359) );
  AND U17092 ( .A(n922), .B(n17375), .Z(n17374) );
  IV U17093 ( .A(n17370), .Z(n17372) );
  XOR U17094 ( .A(n17376), .B(n17377), .Z(n17370) );
  AND U17095 ( .A(n906), .B(n17369), .Z(n17377) );
  XNOR U17096 ( .A(n17367), .B(n17376), .Z(n17369) );
  XNOR U17097 ( .A(n17378), .B(n17379), .Z(n17367) );
  AND U17098 ( .A(n910), .B(n17380), .Z(n17379) );
  XOR U17099 ( .A(p_input[1332]), .B(n17378), .Z(n17380) );
  XNOR U17100 ( .A(n17381), .B(n17382), .Z(n17378) );
  AND U17101 ( .A(n914), .B(n17383), .Z(n17382) );
  XOR U17102 ( .A(n17384), .B(n17385), .Z(n17376) );
  AND U17103 ( .A(n918), .B(n17375), .Z(n17385) );
  XNOR U17104 ( .A(n17386), .B(n17373), .Z(n17375) );
  XOR U17105 ( .A(n17387), .B(n17388), .Z(n17373) );
  AND U17106 ( .A(n941), .B(n17389), .Z(n17388) );
  IV U17107 ( .A(n17384), .Z(n17386) );
  XOR U17108 ( .A(n17390), .B(n17391), .Z(n17384) );
  AND U17109 ( .A(n925), .B(n17383), .Z(n17391) );
  XNOR U17110 ( .A(n17381), .B(n17390), .Z(n17383) );
  XNOR U17111 ( .A(n17392), .B(n17393), .Z(n17381) );
  AND U17112 ( .A(n929), .B(n17394), .Z(n17393) );
  XOR U17113 ( .A(p_input[1364]), .B(n17392), .Z(n17394) );
  XNOR U17114 ( .A(n17395), .B(n17396), .Z(n17392) );
  AND U17115 ( .A(n933), .B(n17397), .Z(n17396) );
  XOR U17116 ( .A(n17398), .B(n17399), .Z(n17390) );
  AND U17117 ( .A(n937), .B(n17389), .Z(n17399) );
  XNOR U17118 ( .A(n17400), .B(n17387), .Z(n17389) );
  XOR U17119 ( .A(n17401), .B(n17402), .Z(n17387) );
  AND U17120 ( .A(n960), .B(n17403), .Z(n17402) );
  IV U17121 ( .A(n17398), .Z(n17400) );
  XOR U17122 ( .A(n17404), .B(n17405), .Z(n17398) );
  AND U17123 ( .A(n944), .B(n17397), .Z(n17405) );
  XNOR U17124 ( .A(n17395), .B(n17404), .Z(n17397) );
  XNOR U17125 ( .A(n17406), .B(n17407), .Z(n17395) );
  AND U17126 ( .A(n948), .B(n17408), .Z(n17407) );
  XOR U17127 ( .A(p_input[1396]), .B(n17406), .Z(n17408) );
  XNOR U17128 ( .A(n17409), .B(n17410), .Z(n17406) );
  AND U17129 ( .A(n952), .B(n17411), .Z(n17410) );
  XOR U17130 ( .A(n17412), .B(n17413), .Z(n17404) );
  AND U17131 ( .A(n956), .B(n17403), .Z(n17413) );
  XNOR U17132 ( .A(n17414), .B(n17401), .Z(n17403) );
  XOR U17133 ( .A(n17415), .B(n17416), .Z(n17401) );
  AND U17134 ( .A(n979), .B(n17417), .Z(n17416) );
  IV U17135 ( .A(n17412), .Z(n17414) );
  XOR U17136 ( .A(n17418), .B(n17419), .Z(n17412) );
  AND U17137 ( .A(n963), .B(n17411), .Z(n17419) );
  XNOR U17138 ( .A(n17409), .B(n17418), .Z(n17411) );
  XNOR U17139 ( .A(n17420), .B(n17421), .Z(n17409) );
  AND U17140 ( .A(n967), .B(n17422), .Z(n17421) );
  XOR U17141 ( .A(p_input[1428]), .B(n17420), .Z(n17422) );
  XNOR U17142 ( .A(n17423), .B(n17424), .Z(n17420) );
  AND U17143 ( .A(n971), .B(n17425), .Z(n17424) );
  XOR U17144 ( .A(n17426), .B(n17427), .Z(n17418) );
  AND U17145 ( .A(n975), .B(n17417), .Z(n17427) );
  XNOR U17146 ( .A(n17428), .B(n17415), .Z(n17417) );
  XOR U17147 ( .A(n17429), .B(n17430), .Z(n17415) );
  AND U17148 ( .A(n998), .B(n17431), .Z(n17430) );
  IV U17149 ( .A(n17426), .Z(n17428) );
  XOR U17150 ( .A(n17432), .B(n17433), .Z(n17426) );
  AND U17151 ( .A(n982), .B(n17425), .Z(n17433) );
  XNOR U17152 ( .A(n17423), .B(n17432), .Z(n17425) );
  XNOR U17153 ( .A(n17434), .B(n17435), .Z(n17423) );
  AND U17154 ( .A(n986), .B(n17436), .Z(n17435) );
  XOR U17155 ( .A(p_input[1460]), .B(n17434), .Z(n17436) );
  XNOR U17156 ( .A(n17437), .B(n17438), .Z(n17434) );
  AND U17157 ( .A(n990), .B(n17439), .Z(n17438) );
  XOR U17158 ( .A(n17440), .B(n17441), .Z(n17432) );
  AND U17159 ( .A(n994), .B(n17431), .Z(n17441) );
  XNOR U17160 ( .A(n17442), .B(n17429), .Z(n17431) );
  XOR U17161 ( .A(n17443), .B(n17444), .Z(n17429) );
  AND U17162 ( .A(n1017), .B(n17445), .Z(n17444) );
  IV U17163 ( .A(n17440), .Z(n17442) );
  XOR U17164 ( .A(n17446), .B(n17447), .Z(n17440) );
  AND U17165 ( .A(n1001), .B(n17439), .Z(n17447) );
  XNOR U17166 ( .A(n17437), .B(n17446), .Z(n17439) );
  XNOR U17167 ( .A(n17448), .B(n17449), .Z(n17437) );
  AND U17168 ( .A(n1005), .B(n17450), .Z(n17449) );
  XOR U17169 ( .A(p_input[1492]), .B(n17448), .Z(n17450) );
  XNOR U17170 ( .A(n17451), .B(n17452), .Z(n17448) );
  AND U17171 ( .A(n1009), .B(n17453), .Z(n17452) );
  XOR U17172 ( .A(n17454), .B(n17455), .Z(n17446) );
  AND U17173 ( .A(n1013), .B(n17445), .Z(n17455) );
  XNOR U17174 ( .A(n17456), .B(n17443), .Z(n17445) );
  XOR U17175 ( .A(n17457), .B(n17458), .Z(n17443) );
  AND U17176 ( .A(n1036), .B(n17459), .Z(n17458) );
  IV U17177 ( .A(n17454), .Z(n17456) );
  XOR U17178 ( .A(n17460), .B(n17461), .Z(n17454) );
  AND U17179 ( .A(n1020), .B(n17453), .Z(n17461) );
  XNOR U17180 ( .A(n17451), .B(n17460), .Z(n17453) );
  XNOR U17181 ( .A(n17462), .B(n17463), .Z(n17451) );
  AND U17182 ( .A(n1024), .B(n17464), .Z(n17463) );
  XOR U17183 ( .A(p_input[1524]), .B(n17462), .Z(n17464) );
  XNOR U17184 ( .A(n17465), .B(n17466), .Z(n17462) );
  AND U17185 ( .A(n1028), .B(n17467), .Z(n17466) );
  XOR U17186 ( .A(n17468), .B(n17469), .Z(n17460) );
  AND U17187 ( .A(n1032), .B(n17459), .Z(n17469) );
  XNOR U17188 ( .A(n17470), .B(n17457), .Z(n17459) );
  XOR U17189 ( .A(n17471), .B(n17472), .Z(n17457) );
  AND U17190 ( .A(n1055), .B(n17473), .Z(n17472) );
  IV U17191 ( .A(n17468), .Z(n17470) );
  XOR U17192 ( .A(n17474), .B(n17475), .Z(n17468) );
  AND U17193 ( .A(n1039), .B(n17467), .Z(n17475) );
  XNOR U17194 ( .A(n17465), .B(n17474), .Z(n17467) );
  XNOR U17195 ( .A(n17476), .B(n17477), .Z(n17465) );
  AND U17196 ( .A(n1043), .B(n17478), .Z(n17477) );
  XOR U17197 ( .A(p_input[1556]), .B(n17476), .Z(n17478) );
  XNOR U17198 ( .A(n17479), .B(n17480), .Z(n17476) );
  AND U17199 ( .A(n1047), .B(n17481), .Z(n17480) );
  XOR U17200 ( .A(n17482), .B(n17483), .Z(n17474) );
  AND U17201 ( .A(n1051), .B(n17473), .Z(n17483) );
  XNOR U17202 ( .A(n17484), .B(n17471), .Z(n17473) );
  XOR U17203 ( .A(n17485), .B(n17486), .Z(n17471) );
  AND U17204 ( .A(n1074), .B(n17487), .Z(n17486) );
  IV U17205 ( .A(n17482), .Z(n17484) );
  XOR U17206 ( .A(n17488), .B(n17489), .Z(n17482) );
  AND U17207 ( .A(n1058), .B(n17481), .Z(n17489) );
  XNOR U17208 ( .A(n17479), .B(n17488), .Z(n17481) );
  XNOR U17209 ( .A(n17490), .B(n17491), .Z(n17479) );
  AND U17210 ( .A(n1062), .B(n17492), .Z(n17491) );
  XOR U17211 ( .A(p_input[1588]), .B(n17490), .Z(n17492) );
  XNOR U17212 ( .A(n17493), .B(n17494), .Z(n17490) );
  AND U17213 ( .A(n1066), .B(n17495), .Z(n17494) );
  XOR U17214 ( .A(n17496), .B(n17497), .Z(n17488) );
  AND U17215 ( .A(n1070), .B(n17487), .Z(n17497) );
  XNOR U17216 ( .A(n17498), .B(n17485), .Z(n17487) );
  XOR U17217 ( .A(n17499), .B(n17500), .Z(n17485) );
  AND U17218 ( .A(n1093), .B(n17501), .Z(n17500) );
  IV U17219 ( .A(n17496), .Z(n17498) );
  XOR U17220 ( .A(n17502), .B(n17503), .Z(n17496) );
  AND U17221 ( .A(n1077), .B(n17495), .Z(n17503) );
  XNOR U17222 ( .A(n17493), .B(n17502), .Z(n17495) );
  XNOR U17223 ( .A(n17504), .B(n17505), .Z(n17493) );
  AND U17224 ( .A(n1081), .B(n17506), .Z(n17505) );
  XOR U17225 ( .A(p_input[1620]), .B(n17504), .Z(n17506) );
  XNOR U17226 ( .A(n17507), .B(n17508), .Z(n17504) );
  AND U17227 ( .A(n1085), .B(n17509), .Z(n17508) );
  XOR U17228 ( .A(n17510), .B(n17511), .Z(n17502) );
  AND U17229 ( .A(n1089), .B(n17501), .Z(n17511) );
  XNOR U17230 ( .A(n17512), .B(n17499), .Z(n17501) );
  XOR U17231 ( .A(n17513), .B(n17514), .Z(n17499) );
  AND U17232 ( .A(n1112), .B(n17515), .Z(n17514) );
  IV U17233 ( .A(n17510), .Z(n17512) );
  XOR U17234 ( .A(n17516), .B(n17517), .Z(n17510) );
  AND U17235 ( .A(n1096), .B(n17509), .Z(n17517) );
  XNOR U17236 ( .A(n17507), .B(n17516), .Z(n17509) );
  XNOR U17237 ( .A(n17518), .B(n17519), .Z(n17507) );
  AND U17238 ( .A(n1100), .B(n17520), .Z(n17519) );
  XOR U17239 ( .A(p_input[1652]), .B(n17518), .Z(n17520) );
  XNOR U17240 ( .A(n17521), .B(n17522), .Z(n17518) );
  AND U17241 ( .A(n1104), .B(n17523), .Z(n17522) );
  XOR U17242 ( .A(n17524), .B(n17525), .Z(n17516) );
  AND U17243 ( .A(n1108), .B(n17515), .Z(n17525) );
  XNOR U17244 ( .A(n17526), .B(n17513), .Z(n17515) );
  XOR U17245 ( .A(n17527), .B(n17528), .Z(n17513) );
  AND U17246 ( .A(n1131), .B(n17529), .Z(n17528) );
  IV U17247 ( .A(n17524), .Z(n17526) );
  XOR U17248 ( .A(n17530), .B(n17531), .Z(n17524) );
  AND U17249 ( .A(n1115), .B(n17523), .Z(n17531) );
  XNOR U17250 ( .A(n17521), .B(n17530), .Z(n17523) );
  XNOR U17251 ( .A(n17532), .B(n17533), .Z(n17521) );
  AND U17252 ( .A(n1119), .B(n17534), .Z(n17533) );
  XOR U17253 ( .A(p_input[1684]), .B(n17532), .Z(n17534) );
  XNOR U17254 ( .A(n17535), .B(n17536), .Z(n17532) );
  AND U17255 ( .A(n1123), .B(n17537), .Z(n17536) );
  XOR U17256 ( .A(n17538), .B(n17539), .Z(n17530) );
  AND U17257 ( .A(n1127), .B(n17529), .Z(n17539) );
  XNOR U17258 ( .A(n17540), .B(n17527), .Z(n17529) );
  XOR U17259 ( .A(n17541), .B(n17542), .Z(n17527) );
  AND U17260 ( .A(n1150), .B(n17543), .Z(n17542) );
  IV U17261 ( .A(n17538), .Z(n17540) );
  XOR U17262 ( .A(n17544), .B(n17545), .Z(n17538) );
  AND U17263 ( .A(n1134), .B(n17537), .Z(n17545) );
  XNOR U17264 ( .A(n17535), .B(n17544), .Z(n17537) );
  XNOR U17265 ( .A(n17546), .B(n17547), .Z(n17535) );
  AND U17266 ( .A(n1138), .B(n17548), .Z(n17547) );
  XOR U17267 ( .A(p_input[1716]), .B(n17546), .Z(n17548) );
  XNOR U17268 ( .A(n17549), .B(n17550), .Z(n17546) );
  AND U17269 ( .A(n1142), .B(n17551), .Z(n17550) );
  XOR U17270 ( .A(n17552), .B(n17553), .Z(n17544) );
  AND U17271 ( .A(n1146), .B(n17543), .Z(n17553) );
  XNOR U17272 ( .A(n17554), .B(n17541), .Z(n17543) );
  XOR U17273 ( .A(n17555), .B(n17556), .Z(n17541) );
  AND U17274 ( .A(n1169), .B(n17557), .Z(n17556) );
  IV U17275 ( .A(n17552), .Z(n17554) );
  XOR U17276 ( .A(n17558), .B(n17559), .Z(n17552) );
  AND U17277 ( .A(n1153), .B(n17551), .Z(n17559) );
  XNOR U17278 ( .A(n17549), .B(n17558), .Z(n17551) );
  XNOR U17279 ( .A(n17560), .B(n17561), .Z(n17549) );
  AND U17280 ( .A(n1157), .B(n17562), .Z(n17561) );
  XOR U17281 ( .A(p_input[1748]), .B(n17560), .Z(n17562) );
  XNOR U17282 ( .A(n17563), .B(n17564), .Z(n17560) );
  AND U17283 ( .A(n1161), .B(n17565), .Z(n17564) );
  XOR U17284 ( .A(n17566), .B(n17567), .Z(n17558) );
  AND U17285 ( .A(n1165), .B(n17557), .Z(n17567) );
  XNOR U17286 ( .A(n17568), .B(n17555), .Z(n17557) );
  XOR U17287 ( .A(n17569), .B(n17570), .Z(n17555) );
  AND U17288 ( .A(n1188), .B(n17571), .Z(n17570) );
  IV U17289 ( .A(n17566), .Z(n17568) );
  XOR U17290 ( .A(n17572), .B(n17573), .Z(n17566) );
  AND U17291 ( .A(n1172), .B(n17565), .Z(n17573) );
  XNOR U17292 ( .A(n17563), .B(n17572), .Z(n17565) );
  XNOR U17293 ( .A(n17574), .B(n17575), .Z(n17563) );
  AND U17294 ( .A(n1176), .B(n17576), .Z(n17575) );
  XOR U17295 ( .A(p_input[1780]), .B(n17574), .Z(n17576) );
  XNOR U17296 ( .A(n17577), .B(n17578), .Z(n17574) );
  AND U17297 ( .A(n1180), .B(n17579), .Z(n17578) );
  XOR U17298 ( .A(n17580), .B(n17581), .Z(n17572) );
  AND U17299 ( .A(n1184), .B(n17571), .Z(n17581) );
  XNOR U17300 ( .A(n17582), .B(n17569), .Z(n17571) );
  XOR U17301 ( .A(n17583), .B(n17584), .Z(n17569) );
  AND U17302 ( .A(n1207), .B(n17585), .Z(n17584) );
  IV U17303 ( .A(n17580), .Z(n17582) );
  XOR U17304 ( .A(n17586), .B(n17587), .Z(n17580) );
  AND U17305 ( .A(n1191), .B(n17579), .Z(n17587) );
  XNOR U17306 ( .A(n17577), .B(n17586), .Z(n17579) );
  XNOR U17307 ( .A(n17588), .B(n17589), .Z(n17577) );
  AND U17308 ( .A(n1195), .B(n17590), .Z(n17589) );
  XOR U17309 ( .A(p_input[1812]), .B(n17588), .Z(n17590) );
  XNOR U17310 ( .A(n17591), .B(n17592), .Z(n17588) );
  AND U17311 ( .A(n1199), .B(n17593), .Z(n17592) );
  XOR U17312 ( .A(n17594), .B(n17595), .Z(n17586) );
  AND U17313 ( .A(n1203), .B(n17585), .Z(n17595) );
  XNOR U17314 ( .A(n17596), .B(n17583), .Z(n17585) );
  XOR U17315 ( .A(n17597), .B(n17598), .Z(n17583) );
  AND U17316 ( .A(n1226), .B(n17599), .Z(n17598) );
  IV U17317 ( .A(n17594), .Z(n17596) );
  XOR U17318 ( .A(n17600), .B(n17601), .Z(n17594) );
  AND U17319 ( .A(n1210), .B(n17593), .Z(n17601) );
  XNOR U17320 ( .A(n17591), .B(n17600), .Z(n17593) );
  XNOR U17321 ( .A(n17602), .B(n17603), .Z(n17591) );
  AND U17322 ( .A(n1214), .B(n17604), .Z(n17603) );
  XOR U17323 ( .A(p_input[1844]), .B(n17602), .Z(n17604) );
  XNOR U17324 ( .A(n17605), .B(n17606), .Z(n17602) );
  AND U17325 ( .A(n1218), .B(n17607), .Z(n17606) );
  XOR U17326 ( .A(n17608), .B(n17609), .Z(n17600) );
  AND U17327 ( .A(n1222), .B(n17599), .Z(n17609) );
  XNOR U17328 ( .A(n17610), .B(n17597), .Z(n17599) );
  XOR U17329 ( .A(n17611), .B(n17612), .Z(n17597) );
  AND U17330 ( .A(n1245), .B(n17613), .Z(n17612) );
  IV U17331 ( .A(n17608), .Z(n17610) );
  XOR U17332 ( .A(n17614), .B(n17615), .Z(n17608) );
  AND U17333 ( .A(n1229), .B(n17607), .Z(n17615) );
  XNOR U17334 ( .A(n17605), .B(n17614), .Z(n17607) );
  XNOR U17335 ( .A(n17616), .B(n17617), .Z(n17605) );
  AND U17336 ( .A(n1233), .B(n17618), .Z(n17617) );
  XOR U17337 ( .A(p_input[1876]), .B(n17616), .Z(n17618) );
  XNOR U17338 ( .A(n17619), .B(n17620), .Z(n17616) );
  AND U17339 ( .A(n1237), .B(n17621), .Z(n17620) );
  XOR U17340 ( .A(n17622), .B(n17623), .Z(n17614) );
  AND U17341 ( .A(n1241), .B(n17613), .Z(n17623) );
  XNOR U17342 ( .A(n17624), .B(n17611), .Z(n17613) );
  XOR U17343 ( .A(n17625), .B(n17626), .Z(n17611) );
  AND U17344 ( .A(n1264), .B(n17627), .Z(n17626) );
  IV U17345 ( .A(n17622), .Z(n17624) );
  XOR U17346 ( .A(n17628), .B(n17629), .Z(n17622) );
  AND U17347 ( .A(n1248), .B(n17621), .Z(n17629) );
  XNOR U17348 ( .A(n17619), .B(n17628), .Z(n17621) );
  XNOR U17349 ( .A(n17630), .B(n17631), .Z(n17619) );
  AND U17350 ( .A(n1252), .B(n17632), .Z(n17631) );
  XOR U17351 ( .A(p_input[1908]), .B(n17630), .Z(n17632) );
  XNOR U17352 ( .A(n17633), .B(n17634), .Z(n17630) );
  AND U17353 ( .A(n1256), .B(n17635), .Z(n17634) );
  XOR U17354 ( .A(n17636), .B(n17637), .Z(n17628) );
  AND U17355 ( .A(n1260), .B(n17627), .Z(n17637) );
  XNOR U17356 ( .A(n17638), .B(n17625), .Z(n17627) );
  XOR U17357 ( .A(n17639), .B(n17640), .Z(n17625) );
  AND U17358 ( .A(n1282), .B(n17641), .Z(n17640) );
  IV U17359 ( .A(n17636), .Z(n17638) );
  XOR U17360 ( .A(n17642), .B(n17643), .Z(n17636) );
  AND U17361 ( .A(n1267), .B(n17635), .Z(n17643) );
  XNOR U17362 ( .A(n17633), .B(n17642), .Z(n17635) );
  XNOR U17363 ( .A(n17644), .B(n17645), .Z(n17633) );
  AND U17364 ( .A(n1271), .B(n17646), .Z(n17645) );
  XOR U17365 ( .A(p_input[1940]), .B(n17644), .Z(n17646) );
  XOR U17366 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][20] ), .B(n17647), 
        .Z(n17644) );
  AND U17367 ( .A(n1274), .B(n17648), .Z(n17647) );
  XOR U17368 ( .A(n17649), .B(n17650), .Z(n17642) );
  AND U17369 ( .A(n1278), .B(n17641), .Z(n17650) );
  XNOR U17370 ( .A(n17651), .B(n17639), .Z(n17641) );
  XOR U17371 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n17652), .Z(n17639) );
  AND U17372 ( .A(n1290), .B(n17653), .Z(n17652) );
  IV U17373 ( .A(n17649), .Z(n17651) );
  XOR U17374 ( .A(n17654), .B(n17655), .Z(n17649) );
  AND U17375 ( .A(n1285), .B(n17648), .Z(n17655) );
  XOR U17376 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][20] ), .B(n17654), 
        .Z(n17648) );
  XOR U17377 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .B(n17656), 
        .Z(n17654) );
  AND U17378 ( .A(n1287), .B(n17653), .Z(n17656) );
  XOR U17379 ( .A(n17657), .B(n17658), .Z(n17653) );
  IV U17380 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .Z(n17658)
         );
  IV U17381 ( .A(\knn_comb_/min_val_out[0][20] ), .Z(n17657) );
  XOR U17382 ( .A(n6465), .B(n17659), .Z(o[1]) );
  AND U17383 ( .A(n122), .B(n17660), .Z(n6465) );
  XOR U17384 ( .A(n6466), .B(n17659), .Z(n17660) );
  XOR U17385 ( .A(n17661), .B(n17662), .Z(n17659) );
  AND U17386 ( .A(n142), .B(n17663), .Z(n17662) );
  XOR U17387 ( .A(n17664), .B(n69), .Z(n6466) );
  AND U17388 ( .A(n125), .B(n17665), .Z(n69) );
  XOR U17389 ( .A(n70), .B(n17664), .Z(n17665) );
  XOR U17390 ( .A(n17666), .B(n17667), .Z(n70) );
  AND U17391 ( .A(n130), .B(n17668), .Z(n17667) );
  XOR U17392 ( .A(p_input[1]), .B(n17666), .Z(n17668) );
  XNOR U17393 ( .A(n17669), .B(n17670), .Z(n17666) );
  AND U17394 ( .A(n134), .B(n17671), .Z(n17670) );
  XOR U17395 ( .A(n17672), .B(n17673), .Z(n17664) );
  AND U17396 ( .A(n138), .B(n17663), .Z(n17673) );
  XNOR U17397 ( .A(n17674), .B(n17661), .Z(n17663) );
  XOR U17398 ( .A(n17675), .B(n17676), .Z(n17661) );
  AND U17399 ( .A(n162), .B(n17677), .Z(n17676) );
  IV U17400 ( .A(n17672), .Z(n17674) );
  XOR U17401 ( .A(n17678), .B(n17679), .Z(n17672) );
  AND U17402 ( .A(n146), .B(n17671), .Z(n17679) );
  XNOR U17403 ( .A(n17669), .B(n17678), .Z(n17671) );
  XNOR U17404 ( .A(n17680), .B(n17681), .Z(n17669) );
  AND U17405 ( .A(n150), .B(n17682), .Z(n17681) );
  XOR U17406 ( .A(p_input[33]), .B(n17680), .Z(n17682) );
  XNOR U17407 ( .A(n17683), .B(n17684), .Z(n17680) );
  AND U17408 ( .A(n154), .B(n17685), .Z(n17684) );
  XOR U17409 ( .A(n17686), .B(n17687), .Z(n17678) );
  AND U17410 ( .A(n158), .B(n17677), .Z(n17687) );
  XNOR U17411 ( .A(n17688), .B(n17675), .Z(n17677) );
  XOR U17412 ( .A(n17689), .B(n17690), .Z(n17675) );
  AND U17413 ( .A(n181), .B(n17691), .Z(n17690) );
  IV U17414 ( .A(n17686), .Z(n17688) );
  XOR U17415 ( .A(n17692), .B(n17693), .Z(n17686) );
  AND U17416 ( .A(n165), .B(n17685), .Z(n17693) );
  XNOR U17417 ( .A(n17683), .B(n17692), .Z(n17685) );
  XNOR U17418 ( .A(n17694), .B(n17695), .Z(n17683) );
  AND U17419 ( .A(n169), .B(n17696), .Z(n17695) );
  XOR U17420 ( .A(p_input[65]), .B(n17694), .Z(n17696) );
  XNOR U17421 ( .A(n17697), .B(n17698), .Z(n17694) );
  AND U17422 ( .A(n173), .B(n17699), .Z(n17698) );
  XOR U17423 ( .A(n17700), .B(n17701), .Z(n17692) );
  AND U17424 ( .A(n177), .B(n17691), .Z(n17701) );
  XNOR U17425 ( .A(n17702), .B(n17689), .Z(n17691) );
  XOR U17426 ( .A(n17703), .B(n17704), .Z(n17689) );
  AND U17427 ( .A(n200), .B(n17705), .Z(n17704) );
  IV U17428 ( .A(n17700), .Z(n17702) );
  XOR U17429 ( .A(n17706), .B(n17707), .Z(n17700) );
  AND U17430 ( .A(n184), .B(n17699), .Z(n17707) );
  XNOR U17431 ( .A(n17697), .B(n17706), .Z(n17699) );
  XNOR U17432 ( .A(n17708), .B(n17709), .Z(n17697) );
  AND U17433 ( .A(n188), .B(n17710), .Z(n17709) );
  XOR U17434 ( .A(p_input[97]), .B(n17708), .Z(n17710) );
  XNOR U17435 ( .A(n17711), .B(n17712), .Z(n17708) );
  AND U17436 ( .A(n192), .B(n17713), .Z(n17712) );
  XOR U17437 ( .A(n17714), .B(n17715), .Z(n17706) );
  AND U17438 ( .A(n196), .B(n17705), .Z(n17715) );
  XNOR U17439 ( .A(n17716), .B(n17703), .Z(n17705) );
  XOR U17440 ( .A(n17717), .B(n17718), .Z(n17703) );
  AND U17441 ( .A(n219), .B(n17719), .Z(n17718) );
  IV U17442 ( .A(n17714), .Z(n17716) );
  XOR U17443 ( .A(n17720), .B(n17721), .Z(n17714) );
  AND U17444 ( .A(n203), .B(n17713), .Z(n17721) );
  XNOR U17445 ( .A(n17711), .B(n17720), .Z(n17713) );
  XNOR U17446 ( .A(n17722), .B(n17723), .Z(n17711) );
  AND U17447 ( .A(n207), .B(n17724), .Z(n17723) );
  XOR U17448 ( .A(p_input[129]), .B(n17722), .Z(n17724) );
  XNOR U17449 ( .A(n17725), .B(n17726), .Z(n17722) );
  AND U17450 ( .A(n211), .B(n17727), .Z(n17726) );
  XOR U17451 ( .A(n17728), .B(n17729), .Z(n17720) );
  AND U17452 ( .A(n215), .B(n17719), .Z(n17729) );
  XNOR U17453 ( .A(n17730), .B(n17717), .Z(n17719) );
  XOR U17454 ( .A(n17731), .B(n17732), .Z(n17717) );
  AND U17455 ( .A(n238), .B(n17733), .Z(n17732) );
  IV U17456 ( .A(n17728), .Z(n17730) );
  XOR U17457 ( .A(n17734), .B(n17735), .Z(n17728) );
  AND U17458 ( .A(n222), .B(n17727), .Z(n17735) );
  XNOR U17459 ( .A(n17725), .B(n17734), .Z(n17727) );
  XNOR U17460 ( .A(n17736), .B(n17737), .Z(n17725) );
  AND U17461 ( .A(n226), .B(n17738), .Z(n17737) );
  XOR U17462 ( .A(p_input[161]), .B(n17736), .Z(n17738) );
  XNOR U17463 ( .A(n17739), .B(n17740), .Z(n17736) );
  AND U17464 ( .A(n230), .B(n17741), .Z(n17740) );
  XOR U17465 ( .A(n17742), .B(n17743), .Z(n17734) );
  AND U17466 ( .A(n234), .B(n17733), .Z(n17743) );
  XNOR U17467 ( .A(n17744), .B(n17731), .Z(n17733) );
  XOR U17468 ( .A(n17745), .B(n17746), .Z(n17731) );
  AND U17469 ( .A(n257), .B(n17747), .Z(n17746) );
  IV U17470 ( .A(n17742), .Z(n17744) );
  XOR U17471 ( .A(n17748), .B(n17749), .Z(n17742) );
  AND U17472 ( .A(n241), .B(n17741), .Z(n17749) );
  XNOR U17473 ( .A(n17739), .B(n17748), .Z(n17741) );
  XNOR U17474 ( .A(n17750), .B(n17751), .Z(n17739) );
  AND U17475 ( .A(n245), .B(n17752), .Z(n17751) );
  XOR U17476 ( .A(p_input[193]), .B(n17750), .Z(n17752) );
  XNOR U17477 ( .A(n17753), .B(n17754), .Z(n17750) );
  AND U17478 ( .A(n249), .B(n17755), .Z(n17754) );
  XOR U17479 ( .A(n17756), .B(n17757), .Z(n17748) );
  AND U17480 ( .A(n253), .B(n17747), .Z(n17757) );
  XNOR U17481 ( .A(n17758), .B(n17745), .Z(n17747) );
  XOR U17482 ( .A(n17759), .B(n17760), .Z(n17745) );
  AND U17483 ( .A(n276), .B(n17761), .Z(n17760) );
  IV U17484 ( .A(n17756), .Z(n17758) );
  XOR U17485 ( .A(n17762), .B(n17763), .Z(n17756) );
  AND U17486 ( .A(n260), .B(n17755), .Z(n17763) );
  XNOR U17487 ( .A(n17753), .B(n17762), .Z(n17755) );
  XNOR U17488 ( .A(n17764), .B(n17765), .Z(n17753) );
  AND U17489 ( .A(n264), .B(n17766), .Z(n17765) );
  XOR U17490 ( .A(p_input[225]), .B(n17764), .Z(n17766) );
  XNOR U17491 ( .A(n17767), .B(n17768), .Z(n17764) );
  AND U17492 ( .A(n268), .B(n17769), .Z(n17768) );
  XOR U17493 ( .A(n17770), .B(n17771), .Z(n17762) );
  AND U17494 ( .A(n272), .B(n17761), .Z(n17771) );
  XNOR U17495 ( .A(n17772), .B(n17759), .Z(n17761) );
  XOR U17496 ( .A(n17773), .B(n17774), .Z(n17759) );
  AND U17497 ( .A(n295), .B(n17775), .Z(n17774) );
  IV U17498 ( .A(n17770), .Z(n17772) );
  XOR U17499 ( .A(n17776), .B(n17777), .Z(n17770) );
  AND U17500 ( .A(n279), .B(n17769), .Z(n17777) );
  XNOR U17501 ( .A(n17767), .B(n17776), .Z(n17769) );
  XNOR U17502 ( .A(n17778), .B(n17779), .Z(n17767) );
  AND U17503 ( .A(n283), .B(n17780), .Z(n17779) );
  XOR U17504 ( .A(p_input[257]), .B(n17778), .Z(n17780) );
  XNOR U17505 ( .A(n17781), .B(n17782), .Z(n17778) );
  AND U17506 ( .A(n287), .B(n17783), .Z(n17782) );
  XOR U17507 ( .A(n17784), .B(n17785), .Z(n17776) );
  AND U17508 ( .A(n291), .B(n17775), .Z(n17785) );
  XNOR U17509 ( .A(n17786), .B(n17773), .Z(n17775) );
  XOR U17510 ( .A(n17787), .B(n17788), .Z(n17773) );
  AND U17511 ( .A(n314), .B(n17789), .Z(n17788) );
  IV U17512 ( .A(n17784), .Z(n17786) );
  XOR U17513 ( .A(n17790), .B(n17791), .Z(n17784) );
  AND U17514 ( .A(n298), .B(n17783), .Z(n17791) );
  XNOR U17515 ( .A(n17781), .B(n17790), .Z(n17783) );
  XNOR U17516 ( .A(n17792), .B(n17793), .Z(n17781) );
  AND U17517 ( .A(n302), .B(n17794), .Z(n17793) );
  XOR U17518 ( .A(p_input[289]), .B(n17792), .Z(n17794) );
  XNOR U17519 ( .A(n17795), .B(n17796), .Z(n17792) );
  AND U17520 ( .A(n306), .B(n17797), .Z(n17796) );
  XOR U17521 ( .A(n17798), .B(n17799), .Z(n17790) );
  AND U17522 ( .A(n310), .B(n17789), .Z(n17799) );
  XNOR U17523 ( .A(n17800), .B(n17787), .Z(n17789) );
  XOR U17524 ( .A(n17801), .B(n17802), .Z(n17787) );
  AND U17525 ( .A(n333), .B(n17803), .Z(n17802) );
  IV U17526 ( .A(n17798), .Z(n17800) );
  XOR U17527 ( .A(n17804), .B(n17805), .Z(n17798) );
  AND U17528 ( .A(n317), .B(n17797), .Z(n17805) );
  XNOR U17529 ( .A(n17795), .B(n17804), .Z(n17797) );
  XNOR U17530 ( .A(n17806), .B(n17807), .Z(n17795) );
  AND U17531 ( .A(n321), .B(n17808), .Z(n17807) );
  XOR U17532 ( .A(p_input[321]), .B(n17806), .Z(n17808) );
  XNOR U17533 ( .A(n17809), .B(n17810), .Z(n17806) );
  AND U17534 ( .A(n325), .B(n17811), .Z(n17810) );
  XOR U17535 ( .A(n17812), .B(n17813), .Z(n17804) );
  AND U17536 ( .A(n329), .B(n17803), .Z(n17813) );
  XNOR U17537 ( .A(n17814), .B(n17801), .Z(n17803) );
  XOR U17538 ( .A(n17815), .B(n17816), .Z(n17801) );
  AND U17539 ( .A(n352), .B(n17817), .Z(n17816) );
  IV U17540 ( .A(n17812), .Z(n17814) );
  XOR U17541 ( .A(n17818), .B(n17819), .Z(n17812) );
  AND U17542 ( .A(n336), .B(n17811), .Z(n17819) );
  XNOR U17543 ( .A(n17809), .B(n17818), .Z(n17811) );
  XNOR U17544 ( .A(n17820), .B(n17821), .Z(n17809) );
  AND U17545 ( .A(n340), .B(n17822), .Z(n17821) );
  XOR U17546 ( .A(p_input[353]), .B(n17820), .Z(n17822) );
  XNOR U17547 ( .A(n17823), .B(n17824), .Z(n17820) );
  AND U17548 ( .A(n344), .B(n17825), .Z(n17824) );
  XOR U17549 ( .A(n17826), .B(n17827), .Z(n17818) );
  AND U17550 ( .A(n348), .B(n17817), .Z(n17827) );
  XNOR U17551 ( .A(n17828), .B(n17815), .Z(n17817) );
  XOR U17552 ( .A(n17829), .B(n17830), .Z(n17815) );
  AND U17553 ( .A(n371), .B(n17831), .Z(n17830) );
  IV U17554 ( .A(n17826), .Z(n17828) );
  XOR U17555 ( .A(n17832), .B(n17833), .Z(n17826) );
  AND U17556 ( .A(n355), .B(n17825), .Z(n17833) );
  XNOR U17557 ( .A(n17823), .B(n17832), .Z(n17825) );
  XNOR U17558 ( .A(n17834), .B(n17835), .Z(n17823) );
  AND U17559 ( .A(n359), .B(n17836), .Z(n17835) );
  XOR U17560 ( .A(p_input[385]), .B(n17834), .Z(n17836) );
  XNOR U17561 ( .A(n17837), .B(n17838), .Z(n17834) );
  AND U17562 ( .A(n363), .B(n17839), .Z(n17838) );
  XOR U17563 ( .A(n17840), .B(n17841), .Z(n17832) );
  AND U17564 ( .A(n367), .B(n17831), .Z(n17841) );
  XNOR U17565 ( .A(n17842), .B(n17829), .Z(n17831) );
  XOR U17566 ( .A(n17843), .B(n17844), .Z(n17829) );
  AND U17567 ( .A(n390), .B(n17845), .Z(n17844) );
  IV U17568 ( .A(n17840), .Z(n17842) );
  XOR U17569 ( .A(n17846), .B(n17847), .Z(n17840) );
  AND U17570 ( .A(n374), .B(n17839), .Z(n17847) );
  XNOR U17571 ( .A(n17837), .B(n17846), .Z(n17839) );
  XNOR U17572 ( .A(n17848), .B(n17849), .Z(n17837) );
  AND U17573 ( .A(n378), .B(n17850), .Z(n17849) );
  XOR U17574 ( .A(p_input[417]), .B(n17848), .Z(n17850) );
  XNOR U17575 ( .A(n17851), .B(n17852), .Z(n17848) );
  AND U17576 ( .A(n382), .B(n17853), .Z(n17852) );
  XOR U17577 ( .A(n17854), .B(n17855), .Z(n17846) );
  AND U17578 ( .A(n386), .B(n17845), .Z(n17855) );
  XNOR U17579 ( .A(n17856), .B(n17843), .Z(n17845) );
  XOR U17580 ( .A(n17857), .B(n17858), .Z(n17843) );
  AND U17581 ( .A(n409), .B(n17859), .Z(n17858) );
  IV U17582 ( .A(n17854), .Z(n17856) );
  XOR U17583 ( .A(n17860), .B(n17861), .Z(n17854) );
  AND U17584 ( .A(n393), .B(n17853), .Z(n17861) );
  XNOR U17585 ( .A(n17851), .B(n17860), .Z(n17853) );
  XNOR U17586 ( .A(n17862), .B(n17863), .Z(n17851) );
  AND U17587 ( .A(n397), .B(n17864), .Z(n17863) );
  XOR U17588 ( .A(p_input[449]), .B(n17862), .Z(n17864) );
  XNOR U17589 ( .A(n17865), .B(n17866), .Z(n17862) );
  AND U17590 ( .A(n401), .B(n17867), .Z(n17866) );
  XOR U17591 ( .A(n17868), .B(n17869), .Z(n17860) );
  AND U17592 ( .A(n405), .B(n17859), .Z(n17869) );
  XNOR U17593 ( .A(n17870), .B(n17857), .Z(n17859) );
  XOR U17594 ( .A(n17871), .B(n17872), .Z(n17857) );
  AND U17595 ( .A(n428), .B(n17873), .Z(n17872) );
  IV U17596 ( .A(n17868), .Z(n17870) );
  XOR U17597 ( .A(n17874), .B(n17875), .Z(n17868) );
  AND U17598 ( .A(n412), .B(n17867), .Z(n17875) );
  XNOR U17599 ( .A(n17865), .B(n17874), .Z(n17867) );
  XNOR U17600 ( .A(n17876), .B(n17877), .Z(n17865) );
  AND U17601 ( .A(n416), .B(n17878), .Z(n17877) );
  XOR U17602 ( .A(p_input[481]), .B(n17876), .Z(n17878) );
  XNOR U17603 ( .A(n17879), .B(n17880), .Z(n17876) );
  AND U17604 ( .A(n420), .B(n17881), .Z(n17880) );
  XOR U17605 ( .A(n17882), .B(n17883), .Z(n17874) );
  AND U17606 ( .A(n424), .B(n17873), .Z(n17883) );
  XNOR U17607 ( .A(n17884), .B(n17871), .Z(n17873) );
  XOR U17608 ( .A(n17885), .B(n17886), .Z(n17871) );
  AND U17609 ( .A(n447), .B(n17887), .Z(n17886) );
  IV U17610 ( .A(n17882), .Z(n17884) );
  XOR U17611 ( .A(n17888), .B(n17889), .Z(n17882) );
  AND U17612 ( .A(n431), .B(n17881), .Z(n17889) );
  XNOR U17613 ( .A(n17879), .B(n17888), .Z(n17881) );
  XNOR U17614 ( .A(n17890), .B(n17891), .Z(n17879) );
  AND U17615 ( .A(n435), .B(n17892), .Z(n17891) );
  XOR U17616 ( .A(p_input[513]), .B(n17890), .Z(n17892) );
  XNOR U17617 ( .A(n17893), .B(n17894), .Z(n17890) );
  AND U17618 ( .A(n439), .B(n17895), .Z(n17894) );
  XOR U17619 ( .A(n17896), .B(n17897), .Z(n17888) );
  AND U17620 ( .A(n443), .B(n17887), .Z(n17897) );
  XNOR U17621 ( .A(n17898), .B(n17885), .Z(n17887) );
  XOR U17622 ( .A(n17899), .B(n17900), .Z(n17885) );
  AND U17623 ( .A(n466), .B(n17901), .Z(n17900) );
  IV U17624 ( .A(n17896), .Z(n17898) );
  XOR U17625 ( .A(n17902), .B(n17903), .Z(n17896) );
  AND U17626 ( .A(n450), .B(n17895), .Z(n17903) );
  XNOR U17627 ( .A(n17893), .B(n17902), .Z(n17895) );
  XNOR U17628 ( .A(n17904), .B(n17905), .Z(n17893) );
  AND U17629 ( .A(n454), .B(n17906), .Z(n17905) );
  XOR U17630 ( .A(p_input[545]), .B(n17904), .Z(n17906) );
  XNOR U17631 ( .A(n17907), .B(n17908), .Z(n17904) );
  AND U17632 ( .A(n458), .B(n17909), .Z(n17908) );
  XOR U17633 ( .A(n17910), .B(n17911), .Z(n17902) );
  AND U17634 ( .A(n462), .B(n17901), .Z(n17911) );
  XNOR U17635 ( .A(n17912), .B(n17899), .Z(n17901) );
  XOR U17636 ( .A(n17913), .B(n17914), .Z(n17899) );
  AND U17637 ( .A(n485), .B(n17915), .Z(n17914) );
  IV U17638 ( .A(n17910), .Z(n17912) );
  XOR U17639 ( .A(n17916), .B(n17917), .Z(n17910) );
  AND U17640 ( .A(n469), .B(n17909), .Z(n17917) );
  XNOR U17641 ( .A(n17907), .B(n17916), .Z(n17909) );
  XNOR U17642 ( .A(n17918), .B(n17919), .Z(n17907) );
  AND U17643 ( .A(n473), .B(n17920), .Z(n17919) );
  XOR U17644 ( .A(p_input[577]), .B(n17918), .Z(n17920) );
  XNOR U17645 ( .A(n17921), .B(n17922), .Z(n17918) );
  AND U17646 ( .A(n477), .B(n17923), .Z(n17922) );
  XOR U17647 ( .A(n17924), .B(n17925), .Z(n17916) );
  AND U17648 ( .A(n481), .B(n17915), .Z(n17925) );
  XNOR U17649 ( .A(n17926), .B(n17913), .Z(n17915) );
  XOR U17650 ( .A(n17927), .B(n17928), .Z(n17913) );
  AND U17651 ( .A(n504), .B(n17929), .Z(n17928) );
  IV U17652 ( .A(n17924), .Z(n17926) );
  XOR U17653 ( .A(n17930), .B(n17931), .Z(n17924) );
  AND U17654 ( .A(n488), .B(n17923), .Z(n17931) );
  XNOR U17655 ( .A(n17921), .B(n17930), .Z(n17923) );
  XNOR U17656 ( .A(n17932), .B(n17933), .Z(n17921) );
  AND U17657 ( .A(n492), .B(n17934), .Z(n17933) );
  XOR U17658 ( .A(p_input[609]), .B(n17932), .Z(n17934) );
  XNOR U17659 ( .A(n17935), .B(n17936), .Z(n17932) );
  AND U17660 ( .A(n496), .B(n17937), .Z(n17936) );
  XOR U17661 ( .A(n17938), .B(n17939), .Z(n17930) );
  AND U17662 ( .A(n500), .B(n17929), .Z(n17939) );
  XNOR U17663 ( .A(n17940), .B(n17927), .Z(n17929) );
  XOR U17664 ( .A(n17941), .B(n17942), .Z(n17927) );
  AND U17665 ( .A(n523), .B(n17943), .Z(n17942) );
  IV U17666 ( .A(n17938), .Z(n17940) );
  XOR U17667 ( .A(n17944), .B(n17945), .Z(n17938) );
  AND U17668 ( .A(n507), .B(n17937), .Z(n17945) );
  XNOR U17669 ( .A(n17935), .B(n17944), .Z(n17937) );
  XNOR U17670 ( .A(n17946), .B(n17947), .Z(n17935) );
  AND U17671 ( .A(n511), .B(n17948), .Z(n17947) );
  XOR U17672 ( .A(p_input[641]), .B(n17946), .Z(n17948) );
  XNOR U17673 ( .A(n17949), .B(n17950), .Z(n17946) );
  AND U17674 ( .A(n515), .B(n17951), .Z(n17950) );
  XOR U17675 ( .A(n17952), .B(n17953), .Z(n17944) );
  AND U17676 ( .A(n519), .B(n17943), .Z(n17953) );
  XNOR U17677 ( .A(n17954), .B(n17941), .Z(n17943) );
  XOR U17678 ( .A(n17955), .B(n17956), .Z(n17941) );
  AND U17679 ( .A(n542), .B(n17957), .Z(n17956) );
  IV U17680 ( .A(n17952), .Z(n17954) );
  XOR U17681 ( .A(n17958), .B(n17959), .Z(n17952) );
  AND U17682 ( .A(n526), .B(n17951), .Z(n17959) );
  XNOR U17683 ( .A(n17949), .B(n17958), .Z(n17951) );
  XNOR U17684 ( .A(n17960), .B(n17961), .Z(n17949) );
  AND U17685 ( .A(n530), .B(n17962), .Z(n17961) );
  XOR U17686 ( .A(p_input[673]), .B(n17960), .Z(n17962) );
  XNOR U17687 ( .A(n17963), .B(n17964), .Z(n17960) );
  AND U17688 ( .A(n534), .B(n17965), .Z(n17964) );
  XOR U17689 ( .A(n17966), .B(n17967), .Z(n17958) );
  AND U17690 ( .A(n538), .B(n17957), .Z(n17967) );
  XNOR U17691 ( .A(n17968), .B(n17955), .Z(n17957) );
  XOR U17692 ( .A(n17969), .B(n17970), .Z(n17955) );
  AND U17693 ( .A(n561), .B(n17971), .Z(n17970) );
  IV U17694 ( .A(n17966), .Z(n17968) );
  XOR U17695 ( .A(n17972), .B(n17973), .Z(n17966) );
  AND U17696 ( .A(n545), .B(n17965), .Z(n17973) );
  XNOR U17697 ( .A(n17963), .B(n17972), .Z(n17965) );
  XNOR U17698 ( .A(n17974), .B(n17975), .Z(n17963) );
  AND U17699 ( .A(n549), .B(n17976), .Z(n17975) );
  XOR U17700 ( .A(p_input[705]), .B(n17974), .Z(n17976) );
  XNOR U17701 ( .A(n17977), .B(n17978), .Z(n17974) );
  AND U17702 ( .A(n553), .B(n17979), .Z(n17978) );
  XOR U17703 ( .A(n17980), .B(n17981), .Z(n17972) );
  AND U17704 ( .A(n557), .B(n17971), .Z(n17981) );
  XNOR U17705 ( .A(n17982), .B(n17969), .Z(n17971) );
  XOR U17706 ( .A(n17983), .B(n17984), .Z(n17969) );
  AND U17707 ( .A(n580), .B(n17985), .Z(n17984) );
  IV U17708 ( .A(n17980), .Z(n17982) );
  XOR U17709 ( .A(n17986), .B(n17987), .Z(n17980) );
  AND U17710 ( .A(n564), .B(n17979), .Z(n17987) );
  XNOR U17711 ( .A(n17977), .B(n17986), .Z(n17979) );
  XNOR U17712 ( .A(n17988), .B(n17989), .Z(n17977) );
  AND U17713 ( .A(n568), .B(n17990), .Z(n17989) );
  XOR U17714 ( .A(p_input[737]), .B(n17988), .Z(n17990) );
  XNOR U17715 ( .A(n17991), .B(n17992), .Z(n17988) );
  AND U17716 ( .A(n572), .B(n17993), .Z(n17992) );
  XOR U17717 ( .A(n17994), .B(n17995), .Z(n17986) );
  AND U17718 ( .A(n576), .B(n17985), .Z(n17995) );
  XNOR U17719 ( .A(n17996), .B(n17983), .Z(n17985) );
  XOR U17720 ( .A(n17997), .B(n17998), .Z(n17983) );
  AND U17721 ( .A(n599), .B(n17999), .Z(n17998) );
  IV U17722 ( .A(n17994), .Z(n17996) );
  XOR U17723 ( .A(n18000), .B(n18001), .Z(n17994) );
  AND U17724 ( .A(n583), .B(n17993), .Z(n18001) );
  XNOR U17725 ( .A(n17991), .B(n18000), .Z(n17993) );
  XNOR U17726 ( .A(n18002), .B(n18003), .Z(n17991) );
  AND U17727 ( .A(n587), .B(n18004), .Z(n18003) );
  XOR U17728 ( .A(p_input[769]), .B(n18002), .Z(n18004) );
  XNOR U17729 ( .A(n18005), .B(n18006), .Z(n18002) );
  AND U17730 ( .A(n591), .B(n18007), .Z(n18006) );
  XOR U17731 ( .A(n18008), .B(n18009), .Z(n18000) );
  AND U17732 ( .A(n595), .B(n17999), .Z(n18009) );
  XNOR U17733 ( .A(n18010), .B(n17997), .Z(n17999) );
  XOR U17734 ( .A(n18011), .B(n18012), .Z(n17997) );
  AND U17735 ( .A(n618), .B(n18013), .Z(n18012) );
  IV U17736 ( .A(n18008), .Z(n18010) );
  XOR U17737 ( .A(n18014), .B(n18015), .Z(n18008) );
  AND U17738 ( .A(n602), .B(n18007), .Z(n18015) );
  XNOR U17739 ( .A(n18005), .B(n18014), .Z(n18007) );
  XNOR U17740 ( .A(n18016), .B(n18017), .Z(n18005) );
  AND U17741 ( .A(n606), .B(n18018), .Z(n18017) );
  XOR U17742 ( .A(p_input[801]), .B(n18016), .Z(n18018) );
  XNOR U17743 ( .A(n18019), .B(n18020), .Z(n18016) );
  AND U17744 ( .A(n610), .B(n18021), .Z(n18020) );
  XOR U17745 ( .A(n18022), .B(n18023), .Z(n18014) );
  AND U17746 ( .A(n614), .B(n18013), .Z(n18023) );
  XNOR U17747 ( .A(n18024), .B(n18011), .Z(n18013) );
  XOR U17748 ( .A(n18025), .B(n18026), .Z(n18011) );
  AND U17749 ( .A(n637), .B(n18027), .Z(n18026) );
  IV U17750 ( .A(n18022), .Z(n18024) );
  XOR U17751 ( .A(n18028), .B(n18029), .Z(n18022) );
  AND U17752 ( .A(n621), .B(n18021), .Z(n18029) );
  XNOR U17753 ( .A(n18019), .B(n18028), .Z(n18021) );
  XNOR U17754 ( .A(n18030), .B(n18031), .Z(n18019) );
  AND U17755 ( .A(n625), .B(n18032), .Z(n18031) );
  XOR U17756 ( .A(p_input[833]), .B(n18030), .Z(n18032) );
  XNOR U17757 ( .A(n18033), .B(n18034), .Z(n18030) );
  AND U17758 ( .A(n629), .B(n18035), .Z(n18034) );
  XOR U17759 ( .A(n18036), .B(n18037), .Z(n18028) );
  AND U17760 ( .A(n633), .B(n18027), .Z(n18037) );
  XNOR U17761 ( .A(n18038), .B(n18025), .Z(n18027) );
  XOR U17762 ( .A(n18039), .B(n18040), .Z(n18025) );
  AND U17763 ( .A(n656), .B(n18041), .Z(n18040) );
  IV U17764 ( .A(n18036), .Z(n18038) );
  XOR U17765 ( .A(n18042), .B(n18043), .Z(n18036) );
  AND U17766 ( .A(n640), .B(n18035), .Z(n18043) );
  XNOR U17767 ( .A(n18033), .B(n18042), .Z(n18035) );
  XNOR U17768 ( .A(n18044), .B(n18045), .Z(n18033) );
  AND U17769 ( .A(n644), .B(n18046), .Z(n18045) );
  XOR U17770 ( .A(p_input[865]), .B(n18044), .Z(n18046) );
  XNOR U17771 ( .A(n18047), .B(n18048), .Z(n18044) );
  AND U17772 ( .A(n648), .B(n18049), .Z(n18048) );
  XOR U17773 ( .A(n18050), .B(n18051), .Z(n18042) );
  AND U17774 ( .A(n652), .B(n18041), .Z(n18051) );
  XNOR U17775 ( .A(n18052), .B(n18039), .Z(n18041) );
  XOR U17776 ( .A(n18053), .B(n18054), .Z(n18039) );
  AND U17777 ( .A(n675), .B(n18055), .Z(n18054) );
  IV U17778 ( .A(n18050), .Z(n18052) );
  XOR U17779 ( .A(n18056), .B(n18057), .Z(n18050) );
  AND U17780 ( .A(n659), .B(n18049), .Z(n18057) );
  XNOR U17781 ( .A(n18047), .B(n18056), .Z(n18049) );
  XNOR U17782 ( .A(n18058), .B(n18059), .Z(n18047) );
  AND U17783 ( .A(n663), .B(n18060), .Z(n18059) );
  XOR U17784 ( .A(p_input[897]), .B(n18058), .Z(n18060) );
  XNOR U17785 ( .A(n18061), .B(n18062), .Z(n18058) );
  AND U17786 ( .A(n667), .B(n18063), .Z(n18062) );
  XOR U17787 ( .A(n18064), .B(n18065), .Z(n18056) );
  AND U17788 ( .A(n671), .B(n18055), .Z(n18065) );
  XNOR U17789 ( .A(n18066), .B(n18053), .Z(n18055) );
  XOR U17790 ( .A(n18067), .B(n18068), .Z(n18053) );
  AND U17791 ( .A(n694), .B(n18069), .Z(n18068) );
  IV U17792 ( .A(n18064), .Z(n18066) );
  XOR U17793 ( .A(n18070), .B(n18071), .Z(n18064) );
  AND U17794 ( .A(n678), .B(n18063), .Z(n18071) );
  XNOR U17795 ( .A(n18061), .B(n18070), .Z(n18063) );
  XNOR U17796 ( .A(n18072), .B(n18073), .Z(n18061) );
  AND U17797 ( .A(n682), .B(n18074), .Z(n18073) );
  XOR U17798 ( .A(p_input[929]), .B(n18072), .Z(n18074) );
  XNOR U17799 ( .A(n18075), .B(n18076), .Z(n18072) );
  AND U17800 ( .A(n686), .B(n18077), .Z(n18076) );
  XOR U17801 ( .A(n18078), .B(n18079), .Z(n18070) );
  AND U17802 ( .A(n690), .B(n18069), .Z(n18079) );
  XNOR U17803 ( .A(n18080), .B(n18067), .Z(n18069) );
  XOR U17804 ( .A(n18081), .B(n18082), .Z(n18067) );
  AND U17805 ( .A(n713), .B(n18083), .Z(n18082) );
  IV U17806 ( .A(n18078), .Z(n18080) );
  XOR U17807 ( .A(n18084), .B(n18085), .Z(n18078) );
  AND U17808 ( .A(n697), .B(n18077), .Z(n18085) );
  XNOR U17809 ( .A(n18075), .B(n18084), .Z(n18077) );
  XNOR U17810 ( .A(n18086), .B(n18087), .Z(n18075) );
  AND U17811 ( .A(n701), .B(n18088), .Z(n18087) );
  XOR U17812 ( .A(p_input[961]), .B(n18086), .Z(n18088) );
  XNOR U17813 ( .A(n18089), .B(n18090), .Z(n18086) );
  AND U17814 ( .A(n705), .B(n18091), .Z(n18090) );
  XOR U17815 ( .A(n18092), .B(n18093), .Z(n18084) );
  AND U17816 ( .A(n709), .B(n18083), .Z(n18093) );
  XNOR U17817 ( .A(n18094), .B(n18081), .Z(n18083) );
  XOR U17818 ( .A(n18095), .B(n18096), .Z(n18081) );
  AND U17819 ( .A(n732), .B(n18097), .Z(n18096) );
  IV U17820 ( .A(n18092), .Z(n18094) );
  XOR U17821 ( .A(n18098), .B(n18099), .Z(n18092) );
  AND U17822 ( .A(n716), .B(n18091), .Z(n18099) );
  XNOR U17823 ( .A(n18089), .B(n18098), .Z(n18091) );
  XNOR U17824 ( .A(n18100), .B(n18101), .Z(n18089) );
  AND U17825 ( .A(n720), .B(n18102), .Z(n18101) );
  XOR U17826 ( .A(p_input[993]), .B(n18100), .Z(n18102) );
  XNOR U17827 ( .A(n18103), .B(n18104), .Z(n18100) );
  AND U17828 ( .A(n724), .B(n18105), .Z(n18104) );
  XOR U17829 ( .A(n18106), .B(n18107), .Z(n18098) );
  AND U17830 ( .A(n728), .B(n18097), .Z(n18107) );
  XNOR U17831 ( .A(n18108), .B(n18095), .Z(n18097) );
  XOR U17832 ( .A(n18109), .B(n18110), .Z(n18095) );
  AND U17833 ( .A(n751), .B(n18111), .Z(n18110) );
  IV U17834 ( .A(n18106), .Z(n18108) );
  XOR U17835 ( .A(n18112), .B(n18113), .Z(n18106) );
  AND U17836 ( .A(n735), .B(n18105), .Z(n18113) );
  XNOR U17837 ( .A(n18103), .B(n18112), .Z(n18105) );
  XNOR U17838 ( .A(n18114), .B(n18115), .Z(n18103) );
  AND U17839 ( .A(n739), .B(n18116), .Z(n18115) );
  XOR U17840 ( .A(p_input[1025]), .B(n18114), .Z(n18116) );
  XNOR U17841 ( .A(n18117), .B(n18118), .Z(n18114) );
  AND U17842 ( .A(n743), .B(n18119), .Z(n18118) );
  XOR U17843 ( .A(n18120), .B(n18121), .Z(n18112) );
  AND U17844 ( .A(n747), .B(n18111), .Z(n18121) );
  XNOR U17845 ( .A(n18122), .B(n18109), .Z(n18111) );
  XOR U17846 ( .A(n18123), .B(n18124), .Z(n18109) );
  AND U17847 ( .A(n770), .B(n18125), .Z(n18124) );
  IV U17848 ( .A(n18120), .Z(n18122) );
  XOR U17849 ( .A(n18126), .B(n18127), .Z(n18120) );
  AND U17850 ( .A(n754), .B(n18119), .Z(n18127) );
  XNOR U17851 ( .A(n18117), .B(n18126), .Z(n18119) );
  XNOR U17852 ( .A(n18128), .B(n18129), .Z(n18117) );
  AND U17853 ( .A(n758), .B(n18130), .Z(n18129) );
  XOR U17854 ( .A(p_input[1057]), .B(n18128), .Z(n18130) );
  XNOR U17855 ( .A(n18131), .B(n18132), .Z(n18128) );
  AND U17856 ( .A(n762), .B(n18133), .Z(n18132) );
  XOR U17857 ( .A(n18134), .B(n18135), .Z(n18126) );
  AND U17858 ( .A(n766), .B(n18125), .Z(n18135) );
  XNOR U17859 ( .A(n18136), .B(n18123), .Z(n18125) );
  XOR U17860 ( .A(n18137), .B(n18138), .Z(n18123) );
  AND U17861 ( .A(n789), .B(n18139), .Z(n18138) );
  IV U17862 ( .A(n18134), .Z(n18136) );
  XOR U17863 ( .A(n18140), .B(n18141), .Z(n18134) );
  AND U17864 ( .A(n773), .B(n18133), .Z(n18141) );
  XNOR U17865 ( .A(n18131), .B(n18140), .Z(n18133) );
  XNOR U17866 ( .A(n18142), .B(n18143), .Z(n18131) );
  AND U17867 ( .A(n777), .B(n18144), .Z(n18143) );
  XOR U17868 ( .A(p_input[1089]), .B(n18142), .Z(n18144) );
  XNOR U17869 ( .A(n18145), .B(n18146), .Z(n18142) );
  AND U17870 ( .A(n781), .B(n18147), .Z(n18146) );
  XOR U17871 ( .A(n18148), .B(n18149), .Z(n18140) );
  AND U17872 ( .A(n785), .B(n18139), .Z(n18149) );
  XNOR U17873 ( .A(n18150), .B(n18137), .Z(n18139) );
  XOR U17874 ( .A(n18151), .B(n18152), .Z(n18137) );
  AND U17875 ( .A(n808), .B(n18153), .Z(n18152) );
  IV U17876 ( .A(n18148), .Z(n18150) );
  XOR U17877 ( .A(n18154), .B(n18155), .Z(n18148) );
  AND U17878 ( .A(n792), .B(n18147), .Z(n18155) );
  XNOR U17879 ( .A(n18145), .B(n18154), .Z(n18147) );
  XNOR U17880 ( .A(n18156), .B(n18157), .Z(n18145) );
  AND U17881 ( .A(n796), .B(n18158), .Z(n18157) );
  XOR U17882 ( .A(p_input[1121]), .B(n18156), .Z(n18158) );
  XNOR U17883 ( .A(n18159), .B(n18160), .Z(n18156) );
  AND U17884 ( .A(n800), .B(n18161), .Z(n18160) );
  XOR U17885 ( .A(n18162), .B(n18163), .Z(n18154) );
  AND U17886 ( .A(n804), .B(n18153), .Z(n18163) );
  XNOR U17887 ( .A(n18164), .B(n18151), .Z(n18153) );
  XOR U17888 ( .A(n18165), .B(n18166), .Z(n18151) );
  AND U17889 ( .A(n827), .B(n18167), .Z(n18166) );
  IV U17890 ( .A(n18162), .Z(n18164) );
  XOR U17891 ( .A(n18168), .B(n18169), .Z(n18162) );
  AND U17892 ( .A(n811), .B(n18161), .Z(n18169) );
  XNOR U17893 ( .A(n18159), .B(n18168), .Z(n18161) );
  XNOR U17894 ( .A(n18170), .B(n18171), .Z(n18159) );
  AND U17895 ( .A(n815), .B(n18172), .Z(n18171) );
  XOR U17896 ( .A(p_input[1153]), .B(n18170), .Z(n18172) );
  XNOR U17897 ( .A(n18173), .B(n18174), .Z(n18170) );
  AND U17898 ( .A(n819), .B(n18175), .Z(n18174) );
  XOR U17899 ( .A(n18176), .B(n18177), .Z(n18168) );
  AND U17900 ( .A(n823), .B(n18167), .Z(n18177) );
  XNOR U17901 ( .A(n18178), .B(n18165), .Z(n18167) );
  XOR U17902 ( .A(n18179), .B(n18180), .Z(n18165) );
  AND U17903 ( .A(n846), .B(n18181), .Z(n18180) );
  IV U17904 ( .A(n18176), .Z(n18178) );
  XOR U17905 ( .A(n18182), .B(n18183), .Z(n18176) );
  AND U17906 ( .A(n830), .B(n18175), .Z(n18183) );
  XNOR U17907 ( .A(n18173), .B(n18182), .Z(n18175) );
  XNOR U17908 ( .A(n18184), .B(n18185), .Z(n18173) );
  AND U17909 ( .A(n834), .B(n18186), .Z(n18185) );
  XOR U17910 ( .A(p_input[1185]), .B(n18184), .Z(n18186) );
  XNOR U17911 ( .A(n18187), .B(n18188), .Z(n18184) );
  AND U17912 ( .A(n838), .B(n18189), .Z(n18188) );
  XOR U17913 ( .A(n18190), .B(n18191), .Z(n18182) );
  AND U17914 ( .A(n842), .B(n18181), .Z(n18191) );
  XNOR U17915 ( .A(n18192), .B(n18179), .Z(n18181) );
  XOR U17916 ( .A(n18193), .B(n18194), .Z(n18179) );
  AND U17917 ( .A(n865), .B(n18195), .Z(n18194) );
  IV U17918 ( .A(n18190), .Z(n18192) );
  XOR U17919 ( .A(n18196), .B(n18197), .Z(n18190) );
  AND U17920 ( .A(n849), .B(n18189), .Z(n18197) );
  XNOR U17921 ( .A(n18187), .B(n18196), .Z(n18189) );
  XNOR U17922 ( .A(n18198), .B(n18199), .Z(n18187) );
  AND U17923 ( .A(n853), .B(n18200), .Z(n18199) );
  XOR U17924 ( .A(p_input[1217]), .B(n18198), .Z(n18200) );
  XNOR U17925 ( .A(n18201), .B(n18202), .Z(n18198) );
  AND U17926 ( .A(n857), .B(n18203), .Z(n18202) );
  XOR U17927 ( .A(n18204), .B(n18205), .Z(n18196) );
  AND U17928 ( .A(n861), .B(n18195), .Z(n18205) );
  XNOR U17929 ( .A(n18206), .B(n18193), .Z(n18195) );
  XOR U17930 ( .A(n18207), .B(n18208), .Z(n18193) );
  AND U17931 ( .A(n884), .B(n18209), .Z(n18208) );
  IV U17932 ( .A(n18204), .Z(n18206) );
  XOR U17933 ( .A(n18210), .B(n18211), .Z(n18204) );
  AND U17934 ( .A(n868), .B(n18203), .Z(n18211) );
  XNOR U17935 ( .A(n18201), .B(n18210), .Z(n18203) );
  XNOR U17936 ( .A(n18212), .B(n18213), .Z(n18201) );
  AND U17937 ( .A(n872), .B(n18214), .Z(n18213) );
  XOR U17938 ( .A(p_input[1249]), .B(n18212), .Z(n18214) );
  XNOR U17939 ( .A(n18215), .B(n18216), .Z(n18212) );
  AND U17940 ( .A(n876), .B(n18217), .Z(n18216) );
  XOR U17941 ( .A(n18218), .B(n18219), .Z(n18210) );
  AND U17942 ( .A(n880), .B(n18209), .Z(n18219) );
  XNOR U17943 ( .A(n18220), .B(n18207), .Z(n18209) );
  XOR U17944 ( .A(n18221), .B(n18222), .Z(n18207) );
  AND U17945 ( .A(n903), .B(n18223), .Z(n18222) );
  IV U17946 ( .A(n18218), .Z(n18220) );
  XOR U17947 ( .A(n18224), .B(n18225), .Z(n18218) );
  AND U17948 ( .A(n887), .B(n18217), .Z(n18225) );
  XNOR U17949 ( .A(n18215), .B(n18224), .Z(n18217) );
  XNOR U17950 ( .A(n18226), .B(n18227), .Z(n18215) );
  AND U17951 ( .A(n891), .B(n18228), .Z(n18227) );
  XOR U17952 ( .A(p_input[1281]), .B(n18226), .Z(n18228) );
  XNOR U17953 ( .A(n18229), .B(n18230), .Z(n18226) );
  AND U17954 ( .A(n895), .B(n18231), .Z(n18230) );
  XOR U17955 ( .A(n18232), .B(n18233), .Z(n18224) );
  AND U17956 ( .A(n899), .B(n18223), .Z(n18233) );
  XNOR U17957 ( .A(n18234), .B(n18221), .Z(n18223) );
  XOR U17958 ( .A(n18235), .B(n18236), .Z(n18221) );
  AND U17959 ( .A(n922), .B(n18237), .Z(n18236) );
  IV U17960 ( .A(n18232), .Z(n18234) );
  XOR U17961 ( .A(n18238), .B(n18239), .Z(n18232) );
  AND U17962 ( .A(n906), .B(n18231), .Z(n18239) );
  XNOR U17963 ( .A(n18229), .B(n18238), .Z(n18231) );
  XNOR U17964 ( .A(n18240), .B(n18241), .Z(n18229) );
  AND U17965 ( .A(n910), .B(n18242), .Z(n18241) );
  XOR U17966 ( .A(p_input[1313]), .B(n18240), .Z(n18242) );
  XNOR U17967 ( .A(n18243), .B(n18244), .Z(n18240) );
  AND U17968 ( .A(n914), .B(n18245), .Z(n18244) );
  XOR U17969 ( .A(n18246), .B(n18247), .Z(n18238) );
  AND U17970 ( .A(n918), .B(n18237), .Z(n18247) );
  XNOR U17971 ( .A(n18248), .B(n18235), .Z(n18237) );
  XOR U17972 ( .A(n18249), .B(n18250), .Z(n18235) );
  AND U17973 ( .A(n941), .B(n18251), .Z(n18250) );
  IV U17974 ( .A(n18246), .Z(n18248) );
  XOR U17975 ( .A(n18252), .B(n18253), .Z(n18246) );
  AND U17976 ( .A(n925), .B(n18245), .Z(n18253) );
  XNOR U17977 ( .A(n18243), .B(n18252), .Z(n18245) );
  XNOR U17978 ( .A(n18254), .B(n18255), .Z(n18243) );
  AND U17979 ( .A(n929), .B(n18256), .Z(n18255) );
  XOR U17980 ( .A(p_input[1345]), .B(n18254), .Z(n18256) );
  XNOR U17981 ( .A(n18257), .B(n18258), .Z(n18254) );
  AND U17982 ( .A(n933), .B(n18259), .Z(n18258) );
  XOR U17983 ( .A(n18260), .B(n18261), .Z(n18252) );
  AND U17984 ( .A(n937), .B(n18251), .Z(n18261) );
  XNOR U17985 ( .A(n18262), .B(n18249), .Z(n18251) );
  XOR U17986 ( .A(n18263), .B(n18264), .Z(n18249) );
  AND U17987 ( .A(n960), .B(n18265), .Z(n18264) );
  IV U17988 ( .A(n18260), .Z(n18262) );
  XOR U17989 ( .A(n18266), .B(n18267), .Z(n18260) );
  AND U17990 ( .A(n944), .B(n18259), .Z(n18267) );
  XNOR U17991 ( .A(n18257), .B(n18266), .Z(n18259) );
  XNOR U17992 ( .A(n18268), .B(n18269), .Z(n18257) );
  AND U17993 ( .A(n948), .B(n18270), .Z(n18269) );
  XOR U17994 ( .A(p_input[1377]), .B(n18268), .Z(n18270) );
  XNOR U17995 ( .A(n18271), .B(n18272), .Z(n18268) );
  AND U17996 ( .A(n952), .B(n18273), .Z(n18272) );
  XOR U17997 ( .A(n18274), .B(n18275), .Z(n18266) );
  AND U17998 ( .A(n956), .B(n18265), .Z(n18275) );
  XNOR U17999 ( .A(n18276), .B(n18263), .Z(n18265) );
  XOR U18000 ( .A(n18277), .B(n18278), .Z(n18263) );
  AND U18001 ( .A(n979), .B(n18279), .Z(n18278) );
  IV U18002 ( .A(n18274), .Z(n18276) );
  XOR U18003 ( .A(n18280), .B(n18281), .Z(n18274) );
  AND U18004 ( .A(n963), .B(n18273), .Z(n18281) );
  XNOR U18005 ( .A(n18271), .B(n18280), .Z(n18273) );
  XNOR U18006 ( .A(n18282), .B(n18283), .Z(n18271) );
  AND U18007 ( .A(n967), .B(n18284), .Z(n18283) );
  XOR U18008 ( .A(p_input[1409]), .B(n18282), .Z(n18284) );
  XNOR U18009 ( .A(n18285), .B(n18286), .Z(n18282) );
  AND U18010 ( .A(n971), .B(n18287), .Z(n18286) );
  XOR U18011 ( .A(n18288), .B(n18289), .Z(n18280) );
  AND U18012 ( .A(n975), .B(n18279), .Z(n18289) );
  XNOR U18013 ( .A(n18290), .B(n18277), .Z(n18279) );
  XOR U18014 ( .A(n18291), .B(n18292), .Z(n18277) );
  AND U18015 ( .A(n998), .B(n18293), .Z(n18292) );
  IV U18016 ( .A(n18288), .Z(n18290) );
  XOR U18017 ( .A(n18294), .B(n18295), .Z(n18288) );
  AND U18018 ( .A(n982), .B(n18287), .Z(n18295) );
  XNOR U18019 ( .A(n18285), .B(n18294), .Z(n18287) );
  XNOR U18020 ( .A(n18296), .B(n18297), .Z(n18285) );
  AND U18021 ( .A(n986), .B(n18298), .Z(n18297) );
  XOR U18022 ( .A(p_input[1441]), .B(n18296), .Z(n18298) );
  XNOR U18023 ( .A(n18299), .B(n18300), .Z(n18296) );
  AND U18024 ( .A(n990), .B(n18301), .Z(n18300) );
  XOR U18025 ( .A(n18302), .B(n18303), .Z(n18294) );
  AND U18026 ( .A(n994), .B(n18293), .Z(n18303) );
  XNOR U18027 ( .A(n18304), .B(n18291), .Z(n18293) );
  XOR U18028 ( .A(n18305), .B(n18306), .Z(n18291) );
  AND U18029 ( .A(n1017), .B(n18307), .Z(n18306) );
  IV U18030 ( .A(n18302), .Z(n18304) );
  XOR U18031 ( .A(n18308), .B(n18309), .Z(n18302) );
  AND U18032 ( .A(n1001), .B(n18301), .Z(n18309) );
  XNOR U18033 ( .A(n18299), .B(n18308), .Z(n18301) );
  XNOR U18034 ( .A(n18310), .B(n18311), .Z(n18299) );
  AND U18035 ( .A(n1005), .B(n18312), .Z(n18311) );
  XOR U18036 ( .A(p_input[1473]), .B(n18310), .Z(n18312) );
  XNOR U18037 ( .A(n18313), .B(n18314), .Z(n18310) );
  AND U18038 ( .A(n1009), .B(n18315), .Z(n18314) );
  XOR U18039 ( .A(n18316), .B(n18317), .Z(n18308) );
  AND U18040 ( .A(n1013), .B(n18307), .Z(n18317) );
  XNOR U18041 ( .A(n18318), .B(n18305), .Z(n18307) );
  XOR U18042 ( .A(n18319), .B(n18320), .Z(n18305) );
  AND U18043 ( .A(n1036), .B(n18321), .Z(n18320) );
  IV U18044 ( .A(n18316), .Z(n18318) );
  XOR U18045 ( .A(n18322), .B(n18323), .Z(n18316) );
  AND U18046 ( .A(n1020), .B(n18315), .Z(n18323) );
  XNOR U18047 ( .A(n18313), .B(n18322), .Z(n18315) );
  XNOR U18048 ( .A(n18324), .B(n18325), .Z(n18313) );
  AND U18049 ( .A(n1024), .B(n18326), .Z(n18325) );
  XOR U18050 ( .A(p_input[1505]), .B(n18324), .Z(n18326) );
  XNOR U18051 ( .A(n18327), .B(n18328), .Z(n18324) );
  AND U18052 ( .A(n1028), .B(n18329), .Z(n18328) );
  XOR U18053 ( .A(n18330), .B(n18331), .Z(n18322) );
  AND U18054 ( .A(n1032), .B(n18321), .Z(n18331) );
  XNOR U18055 ( .A(n18332), .B(n18319), .Z(n18321) );
  XOR U18056 ( .A(n18333), .B(n18334), .Z(n18319) );
  AND U18057 ( .A(n1055), .B(n18335), .Z(n18334) );
  IV U18058 ( .A(n18330), .Z(n18332) );
  XOR U18059 ( .A(n18336), .B(n18337), .Z(n18330) );
  AND U18060 ( .A(n1039), .B(n18329), .Z(n18337) );
  XNOR U18061 ( .A(n18327), .B(n18336), .Z(n18329) );
  XNOR U18062 ( .A(n18338), .B(n18339), .Z(n18327) );
  AND U18063 ( .A(n1043), .B(n18340), .Z(n18339) );
  XOR U18064 ( .A(p_input[1537]), .B(n18338), .Z(n18340) );
  XNOR U18065 ( .A(n18341), .B(n18342), .Z(n18338) );
  AND U18066 ( .A(n1047), .B(n18343), .Z(n18342) );
  XOR U18067 ( .A(n18344), .B(n18345), .Z(n18336) );
  AND U18068 ( .A(n1051), .B(n18335), .Z(n18345) );
  XNOR U18069 ( .A(n18346), .B(n18333), .Z(n18335) );
  XOR U18070 ( .A(n18347), .B(n18348), .Z(n18333) );
  AND U18071 ( .A(n1074), .B(n18349), .Z(n18348) );
  IV U18072 ( .A(n18344), .Z(n18346) );
  XOR U18073 ( .A(n18350), .B(n18351), .Z(n18344) );
  AND U18074 ( .A(n1058), .B(n18343), .Z(n18351) );
  XNOR U18075 ( .A(n18341), .B(n18350), .Z(n18343) );
  XNOR U18076 ( .A(n18352), .B(n18353), .Z(n18341) );
  AND U18077 ( .A(n1062), .B(n18354), .Z(n18353) );
  XOR U18078 ( .A(p_input[1569]), .B(n18352), .Z(n18354) );
  XNOR U18079 ( .A(n18355), .B(n18356), .Z(n18352) );
  AND U18080 ( .A(n1066), .B(n18357), .Z(n18356) );
  XOR U18081 ( .A(n18358), .B(n18359), .Z(n18350) );
  AND U18082 ( .A(n1070), .B(n18349), .Z(n18359) );
  XNOR U18083 ( .A(n18360), .B(n18347), .Z(n18349) );
  XOR U18084 ( .A(n18361), .B(n18362), .Z(n18347) );
  AND U18085 ( .A(n1093), .B(n18363), .Z(n18362) );
  IV U18086 ( .A(n18358), .Z(n18360) );
  XOR U18087 ( .A(n18364), .B(n18365), .Z(n18358) );
  AND U18088 ( .A(n1077), .B(n18357), .Z(n18365) );
  XNOR U18089 ( .A(n18355), .B(n18364), .Z(n18357) );
  XNOR U18090 ( .A(n18366), .B(n18367), .Z(n18355) );
  AND U18091 ( .A(n1081), .B(n18368), .Z(n18367) );
  XOR U18092 ( .A(p_input[1601]), .B(n18366), .Z(n18368) );
  XNOR U18093 ( .A(n18369), .B(n18370), .Z(n18366) );
  AND U18094 ( .A(n1085), .B(n18371), .Z(n18370) );
  XOR U18095 ( .A(n18372), .B(n18373), .Z(n18364) );
  AND U18096 ( .A(n1089), .B(n18363), .Z(n18373) );
  XNOR U18097 ( .A(n18374), .B(n18361), .Z(n18363) );
  XOR U18098 ( .A(n18375), .B(n18376), .Z(n18361) );
  AND U18099 ( .A(n1112), .B(n18377), .Z(n18376) );
  IV U18100 ( .A(n18372), .Z(n18374) );
  XOR U18101 ( .A(n18378), .B(n18379), .Z(n18372) );
  AND U18102 ( .A(n1096), .B(n18371), .Z(n18379) );
  XNOR U18103 ( .A(n18369), .B(n18378), .Z(n18371) );
  XNOR U18104 ( .A(n18380), .B(n18381), .Z(n18369) );
  AND U18105 ( .A(n1100), .B(n18382), .Z(n18381) );
  XOR U18106 ( .A(p_input[1633]), .B(n18380), .Z(n18382) );
  XNOR U18107 ( .A(n18383), .B(n18384), .Z(n18380) );
  AND U18108 ( .A(n1104), .B(n18385), .Z(n18384) );
  XOR U18109 ( .A(n18386), .B(n18387), .Z(n18378) );
  AND U18110 ( .A(n1108), .B(n18377), .Z(n18387) );
  XNOR U18111 ( .A(n18388), .B(n18375), .Z(n18377) );
  XOR U18112 ( .A(n18389), .B(n18390), .Z(n18375) );
  AND U18113 ( .A(n1131), .B(n18391), .Z(n18390) );
  IV U18114 ( .A(n18386), .Z(n18388) );
  XOR U18115 ( .A(n18392), .B(n18393), .Z(n18386) );
  AND U18116 ( .A(n1115), .B(n18385), .Z(n18393) );
  XNOR U18117 ( .A(n18383), .B(n18392), .Z(n18385) );
  XNOR U18118 ( .A(n18394), .B(n18395), .Z(n18383) );
  AND U18119 ( .A(n1119), .B(n18396), .Z(n18395) );
  XOR U18120 ( .A(p_input[1665]), .B(n18394), .Z(n18396) );
  XNOR U18121 ( .A(n18397), .B(n18398), .Z(n18394) );
  AND U18122 ( .A(n1123), .B(n18399), .Z(n18398) );
  XOR U18123 ( .A(n18400), .B(n18401), .Z(n18392) );
  AND U18124 ( .A(n1127), .B(n18391), .Z(n18401) );
  XNOR U18125 ( .A(n18402), .B(n18389), .Z(n18391) );
  XOR U18126 ( .A(n18403), .B(n18404), .Z(n18389) );
  AND U18127 ( .A(n1150), .B(n18405), .Z(n18404) );
  IV U18128 ( .A(n18400), .Z(n18402) );
  XOR U18129 ( .A(n18406), .B(n18407), .Z(n18400) );
  AND U18130 ( .A(n1134), .B(n18399), .Z(n18407) );
  XNOR U18131 ( .A(n18397), .B(n18406), .Z(n18399) );
  XNOR U18132 ( .A(n18408), .B(n18409), .Z(n18397) );
  AND U18133 ( .A(n1138), .B(n18410), .Z(n18409) );
  XOR U18134 ( .A(p_input[1697]), .B(n18408), .Z(n18410) );
  XNOR U18135 ( .A(n18411), .B(n18412), .Z(n18408) );
  AND U18136 ( .A(n1142), .B(n18413), .Z(n18412) );
  XOR U18137 ( .A(n18414), .B(n18415), .Z(n18406) );
  AND U18138 ( .A(n1146), .B(n18405), .Z(n18415) );
  XNOR U18139 ( .A(n18416), .B(n18403), .Z(n18405) );
  XOR U18140 ( .A(n18417), .B(n18418), .Z(n18403) );
  AND U18141 ( .A(n1169), .B(n18419), .Z(n18418) );
  IV U18142 ( .A(n18414), .Z(n18416) );
  XOR U18143 ( .A(n18420), .B(n18421), .Z(n18414) );
  AND U18144 ( .A(n1153), .B(n18413), .Z(n18421) );
  XNOR U18145 ( .A(n18411), .B(n18420), .Z(n18413) );
  XNOR U18146 ( .A(n18422), .B(n18423), .Z(n18411) );
  AND U18147 ( .A(n1157), .B(n18424), .Z(n18423) );
  XOR U18148 ( .A(p_input[1729]), .B(n18422), .Z(n18424) );
  XNOR U18149 ( .A(n18425), .B(n18426), .Z(n18422) );
  AND U18150 ( .A(n1161), .B(n18427), .Z(n18426) );
  XOR U18151 ( .A(n18428), .B(n18429), .Z(n18420) );
  AND U18152 ( .A(n1165), .B(n18419), .Z(n18429) );
  XNOR U18153 ( .A(n18430), .B(n18417), .Z(n18419) );
  XOR U18154 ( .A(n18431), .B(n18432), .Z(n18417) );
  AND U18155 ( .A(n1188), .B(n18433), .Z(n18432) );
  IV U18156 ( .A(n18428), .Z(n18430) );
  XOR U18157 ( .A(n18434), .B(n18435), .Z(n18428) );
  AND U18158 ( .A(n1172), .B(n18427), .Z(n18435) );
  XNOR U18159 ( .A(n18425), .B(n18434), .Z(n18427) );
  XNOR U18160 ( .A(n18436), .B(n18437), .Z(n18425) );
  AND U18161 ( .A(n1176), .B(n18438), .Z(n18437) );
  XOR U18162 ( .A(p_input[1761]), .B(n18436), .Z(n18438) );
  XNOR U18163 ( .A(n18439), .B(n18440), .Z(n18436) );
  AND U18164 ( .A(n1180), .B(n18441), .Z(n18440) );
  XOR U18165 ( .A(n18442), .B(n18443), .Z(n18434) );
  AND U18166 ( .A(n1184), .B(n18433), .Z(n18443) );
  XNOR U18167 ( .A(n18444), .B(n18431), .Z(n18433) );
  XOR U18168 ( .A(n18445), .B(n18446), .Z(n18431) );
  AND U18169 ( .A(n1207), .B(n18447), .Z(n18446) );
  IV U18170 ( .A(n18442), .Z(n18444) );
  XOR U18171 ( .A(n18448), .B(n18449), .Z(n18442) );
  AND U18172 ( .A(n1191), .B(n18441), .Z(n18449) );
  XNOR U18173 ( .A(n18439), .B(n18448), .Z(n18441) );
  XNOR U18174 ( .A(n18450), .B(n18451), .Z(n18439) );
  AND U18175 ( .A(n1195), .B(n18452), .Z(n18451) );
  XOR U18176 ( .A(p_input[1793]), .B(n18450), .Z(n18452) );
  XNOR U18177 ( .A(n18453), .B(n18454), .Z(n18450) );
  AND U18178 ( .A(n1199), .B(n18455), .Z(n18454) );
  XOR U18179 ( .A(n18456), .B(n18457), .Z(n18448) );
  AND U18180 ( .A(n1203), .B(n18447), .Z(n18457) );
  XNOR U18181 ( .A(n18458), .B(n18445), .Z(n18447) );
  XOR U18182 ( .A(n18459), .B(n18460), .Z(n18445) );
  AND U18183 ( .A(n1226), .B(n18461), .Z(n18460) );
  IV U18184 ( .A(n18456), .Z(n18458) );
  XOR U18185 ( .A(n18462), .B(n18463), .Z(n18456) );
  AND U18186 ( .A(n1210), .B(n18455), .Z(n18463) );
  XNOR U18187 ( .A(n18453), .B(n18462), .Z(n18455) );
  XNOR U18188 ( .A(n18464), .B(n18465), .Z(n18453) );
  AND U18189 ( .A(n1214), .B(n18466), .Z(n18465) );
  XOR U18190 ( .A(p_input[1825]), .B(n18464), .Z(n18466) );
  XNOR U18191 ( .A(n18467), .B(n18468), .Z(n18464) );
  AND U18192 ( .A(n1218), .B(n18469), .Z(n18468) );
  XOR U18193 ( .A(n18470), .B(n18471), .Z(n18462) );
  AND U18194 ( .A(n1222), .B(n18461), .Z(n18471) );
  XNOR U18195 ( .A(n18472), .B(n18459), .Z(n18461) );
  XOR U18196 ( .A(n18473), .B(n18474), .Z(n18459) );
  AND U18197 ( .A(n1245), .B(n18475), .Z(n18474) );
  IV U18198 ( .A(n18470), .Z(n18472) );
  XOR U18199 ( .A(n18476), .B(n18477), .Z(n18470) );
  AND U18200 ( .A(n1229), .B(n18469), .Z(n18477) );
  XNOR U18201 ( .A(n18467), .B(n18476), .Z(n18469) );
  XNOR U18202 ( .A(n18478), .B(n18479), .Z(n18467) );
  AND U18203 ( .A(n1233), .B(n18480), .Z(n18479) );
  XOR U18204 ( .A(p_input[1857]), .B(n18478), .Z(n18480) );
  XNOR U18205 ( .A(n18481), .B(n18482), .Z(n18478) );
  AND U18206 ( .A(n1237), .B(n18483), .Z(n18482) );
  XOR U18207 ( .A(n18484), .B(n18485), .Z(n18476) );
  AND U18208 ( .A(n1241), .B(n18475), .Z(n18485) );
  XNOR U18209 ( .A(n18486), .B(n18473), .Z(n18475) );
  XOR U18210 ( .A(n18487), .B(n18488), .Z(n18473) );
  AND U18211 ( .A(n1264), .B(n18489), .Z(n18488) );
  IV U18212 ( .A(n18484), .Z(n18486) );
  XOR U18213 ( .A(n18490), .B(n18491), .Z(n18484) );
  AND U18214 ( .A(n1248), .B(n18483), .Z(n18491) );
  XNOR U18215 ( .A(n18481), .B(n18490), .Z(n18483) );
  XNOR U18216 ( .A(n18492), .B(n18493), .Z(n18481) );
  AND U18217 ( .A(n1252), .B(n18494), .Z(n18493) );
  XOR U18218 ( .A(p_input[1889]), .B(n18492), .Z(n18494) );
  XNOR U18219 ( .A(n18495), .B(n18496), .Z(n18492) );
  AND U18220 ( .A(n1256), .B(n18497), .Z(n18496) );
  XOR U18221 ( .A(n18498), .B(n18499), .Z(n18490) );
  AND U18222 ( .A(n1260), .B(n18489), .Z(n18499) );
  XNOR U18223 ( .A(n18500), .B(n18487), .Z(n18489) );
  XOR U18224 ( .A(n18501), .B(n18502), .Z(n18487) );
  AND U18225 ( .A(n1282), .B(n18503), .Z(n18502) );
  IV U18226 ( .A(n18498), .Z(n18500) );
  XOR U18227 ( .A(n18504), .B(n18505), .Z(n18498) );
  AND U18228 ( .A(n1267), .B(n18497), .Z(n18505) );
  XNOR U18229 ( .A(n18495), .B(n18504), .Z(n18497) );
  XNOR U18230 ( .A(n18506), .B(n18507), .Z(n18495) );
  AND U18231 ( .A(n1271), .B(n18508), .Z(n18507) );
  XOR U18232 ( .A(p_input[1921]), .B(n18506), .Z(n18508) );
  XOR U18233 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n18509), 
        .Z(n18506) );
  AND U18234 ( .A(n1274), .B(n18510), .Z(n18509) );
  XOR U18235 ( .A(n18511), .B(n18512), .Z(n18504) );
  AND U18236 ( .A(n1278), .B(n18503), .Z(n18512) );
  XNOR U18237 ( .A(n18513), .B(n18501), .Z(n18503) );
  XOR U18238 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n18514), .Z(n18501) );
  AND U18239 ( .A(n1290), .B(n18515), .Z(n18514) );
  IV U18240 ( .A(n18511), .Z(n18513) );
  XOR U18241 ( .A(n18516), .B(n18517), .Z(n18511) );
  AND U18242 ( .A(n1285), .B(n18510), .Z(n18517) );
  XOR U18243 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n18516), 
        .Z(n18510) );
  XOR U18244 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(n18518), 
        .Z(n18516) );
  AND U18245 ( .A(n1287), .B(n18515), .Z(n18518) );
  XOR U18246 ( .A(\knn_comb_/min_val_out[0][1] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n18515) );
  XOR U18247 ( .A(n99), .B(n18519), .Z(o[19]) );
  AND U18248 ( .A(n122), .B(n18520), .Z(n99) );
  XOR U18249 ( .A(n100), .B(n18519), .Z(n18520) );
  XOR U18250 ( .A(n18521), .B(n18522), .Z(n18519) );
  AND U18251 ( .A(n142), .B(n18523), .Z(n18522) );
  XOR U18252 ( .A(n18524), .B(n29), .Z(n100) );
  AND U18253 ( .A(n125), .B(n18525), .Z(n29) );
  XOR U18254 ( .A(n30), .B(n18524), .Z(n18525) );
  XOR U18255 ( .A(n18526), .B(n18527), .Z(n30) );
  AND U18256 ( .A(n130), .B(n18528), .Z(n18527) );
  XOR U18257 ( .A(p_input[19]), .B(n18526), .Z(n18528) );
  XNOR U18258 ( .A(n18529), .B(n18530), .Z(n18526) );
  AND U18259 ( .A(n134), .B(n18531), .Z(n18530) );
  XOR U18260 ( .A(n18532), .B(n18533), .Z(n18524) );
  AND U18261 ( .A(n138), .B(n18523), .Z(n18533) );
  XNOR U18262 ( .A(n18534), .B(n18521), .Z(n18523) );
  XOR U18263 ( .A(n18535), .B(n18536), .Z(n18521) );
  AND U18264 ( .A(n162), .B(n18537), .Z(n18536) );
  IV U18265 ( .A(n18532), .Z(n18534) );
  XOR U18266 ( .A(n18538), .B(n18539), .Z(n18532) );
  AND U18267 ( .A(n146), .B(n18531), .Z(n18539) );
  XNOR U18268 ( .A(n18529), .B(n18538), .Z(n18531) );
  XNOR U18269 ( .A(n18540), .B(n18541), .Z(n18529) );
  AND U18270 ( .A(n150), .B(n18542), .Z(n18541) );
  XOR U18271 ( .A(p_input[51]), .B(n18540), .Z(n18542) );
  XNOR U18272 ( .A(n18543), .B(n18544), .Z(n18540) );
  AND U18273 ( .A(n154), .B(n18545), .Z(n18544) );
  XOR U18274 ( .A(n18546), .B(n18547), .Z(n18538) );
  AND U18275 ( .A(n158), .B(n18537), .Z(n18547) );
  XNOR U18276 ( .A(n18548), .B(n18535), .Z(n18537) );
  XOR U18277 ( .A(n18549), .B(n18550), .Z(n18535) );
  AND U18278 ( .A(n181), .B(n18551), .Z(n18550) );
  IV U18279 ( .A(n18546), .Z(n18548) );
  XOR U18280 ( .A(n18552), .B(n18553), .Z(n18546) );
  AND U18281 ( .A(n165), .B(n18545), .Z(n18553) );
  XNOR U18282 ( .A(n18543), .B(n18552), .Z(n18545) );
  XNOR U18283 ( .A(n18554), .B(n18555), .Z(n18543) );
  AND U18284 ( .A(n169), .B(n18556), .Z(n18555) );
  XOR U18285 ( .A(p_input[83]), .B(n18554), .Z(n18556) );
  XNOR U18286 ( .A(n18557), .B(n18558), .Z(n18554) );
  AND U18287 ( .A(n173), .B(n18559), .Z(n18558) );
  XOR U18288 ( .A(n18560), .B(n18561), .Z(n18552) );
  AND U18289 ( .A(n177), .B(n18551), .Z(n18561) );
  XNOR U18290 ( .A(n18562), .B(n18549), .Z(n18551) );
  XOR U18291 ( .A(n18563), .B(n18564), .Z(n18549) );
  AND U18292 ( .A(n200), .B(n18565), .Z(n18564) );
  IV U18293 ( .A(n18560), .Z(n18562) );
  XOR U18294 ( .A(n18566), .B(n18567), .Z(n18560) );
  AND U18295 ( .A(n184), .B(n18559), .Z(n18567) );
  XNOR U18296 ( .A(n18557), .B(n18566), .Z(n18559) );
  XNOR U18297 ( .A(n18568), .B(n18569), .Z(n18557) );
  AND U18298 ( .A(n188), .B(n18570), .Z(n18569) );
  XOR U18299 ( .A(p_input[115]), .B(n18568), .Z(n18570) );
  XNOR U18300 ( .A(n18571), .B(n18572), .Z(n18568) );
  AND U18301 ( .A(n192), .B(n18573), .Z(n18572) );
  XOR U18302 ( .A(n18574), .B(n18575), .Z(n18566) );
  AND U18303 ( .A(n196), .B(n18565), .Z(n18575) );
  XNOR U18304 ( .A(n18576), .B(n18563), .Z(n18565) );
  XOR U18305 ( .A(n18577), .B(n18578), .Z(n18563) );
  AND U18306 ( .A(n219), .B(n18579), .Z(n18578) );
  IV U18307 ( .A(n18574), .Z(n18576) );
  XOR U18308 ( .A(n18580), .B(n18581), .Z(n18574) );
  AND U18309 ( .A(n203), .B(n18573), .Z(n18581) );
  XNOR U18310 ( .A(n18571), .B(n18580), .Z(n18573) );
  XNOR U18311 ( .A(n18582), .B(n18583), .Z(n18571) );
  AND U18312 ( .A(n207), .B(n18584), .Z(n18583) );
  XOR U18313 ( .A(p_input[147]), .B(n18582), .Z(n18584) );
  XNOR U18314 ( .A(n18585), .B(n18586), .Z(n18582) );
  AND U18315 ( .A(n211), .B(n18587), .Z(n18586) );
  XOR U18316 ( .A(n18588), .B(n18589), .Z(n18580) );
  AND U18317 ( .A(n215), .B(n18579), .Z(n18589) );
  XNOR U18318 ( .A(n18590), .B(n18577), .Z(n18579) );
  XOR U18319 ( .A(n18591), .B(n18592), .Z(n18577) );
  AND U18320 ( .A(n238), .B(n18593), .Z(n18592) );
  IV U18321 ( .A(n18588), .Z(n18590) );
  XOR U18322 ( .A(n18594), .B(n18595), .Z(n18588) );
  AND U18323 ( .A(n222), .B(n18587), .Z(n18595) );
  XNOR U18324 ( .A(n18585), .B(n18594), .Z(n18587) );
  XNOR U18325 ( .A(n18596), .B(n18597), .Z(n18585) );
  AND U18326 ( .A(n226), .B(n18598), .Z(n18597) );
  XOR U18327 ( .A(p_input[179]), .B(n18596), .Z(n18598) );
  XNOR U18328 ( .A(n18599), .B(n18600), .Z(n18596) );
  AND U18329 ( .A(n230), .B(n18601), .Z(n18600) );
  XOR U18330 ( .A(n18602), .B(n18603), .Z(n18594) );
  AND U18331 ( .A(n234), .B(n18593), .Z(n18603) );
  XNOR U18332 ( .A(n18604), .B(n18591), .Z(n18593) );
  XOR U18333 ( .A(n18605), .B(n18606), .Z(n18591) );
  AND U18334 ( .A(n257), .B(n18607), .Z(n18606) );
  IV U18335 ( .A(n18602), .Z(n18604) );
  XOR U18336 ( .A(n18608), .B(n18609), .Z(n18602) );
  AND U18337 ( .A(n241), .B(n18601), .Z(n18609) );
  XNOR U18338 ( .A(n18599), .B(n18608), .Z(n18601) );
  XNOR U18339 ( .A(n18610), .B(n18611), .Z(n18599) );
  AND U18340 ( .A(n245), .B(n18612), .Z(n18611) );
  XOR U18341 ( .A(p_input[211]), .B(n18610), .Z(n18612) );
  XNOR U18342 ( .A(n18613), .B(n18614), .Z(n18610) );
  AND U18343 ( .A(n249), .B(n18615), .Z(n18614) );
  XOR U18344 ( .A(n18616), .B(n18617), .Z(n18608) );
  AND U18345 ( .A(n253), .B(n18607), .Z(n18617) );
  XNOR U18346 ( .A(n18618), .B(n18605), .Z(n18607) );
  XOR U18347 ( .A(n18619), .B(n18620), .Z(n18605) );
  AND U18348 ( .A(n276), .B(n18621), .Z(n18620) );
  IV U18349 ( .A(n18616), .Z(n18618) );
  XOR U18350 ( .A(n18622), .B(n18623), .Z(n18616) );
  AND U18351 ( .A(n260), .B(n18615), .Z(n18623) );
  XNOR U18352 ( .A(n18613), .B(n18622), .Z(n18615) );
  XNOR U18353 ( .A(n18624), .B(n18625), .Z(n18613) );
  AND U18354 ( .A(n264), .B(n18626), .Z(n18625) );
  XOR U18355 ( .A(p_input[243]), .B(n18624), .Z(n18626) );
  XNOR U18356 ( .A(n18627), .B(n18628), .Z(n18624) );
  AND U18357 ( .A(n268), .B(n18629), .Z(n18628) );
  XOR U18358 ( .A(n18630), .B(n18631), .Z(n18622) );
  AND U18359 ( .A(n272), .B(n18621), .Z(n18631) );
  XNOR U18360 ( .A(n18632), .B(n18619), .Z(n18621) );
  XOR U18361 ( .A(n18633), .B(n18634), .Z(n18619) );
  AND U18362 ( .A(n295), .B(n18635), .Z(n18634) );
  IV U18363 ( .A(n18630), .Z(n18632) );
  XOR U18364 ( .A(n18636), .B(n18637), .Z(n18630) );
  AND U18365 ( .A(n279), .B(n18629), .Z(n18637) );
  XNOR U18366 ( .A(n18627), .B(n18636), .Z(n18629) );
  XNOR U18367 ( .A(n18638), .B(n18639), .Z(n18627) );
  AND U18368 ( .A(n283), .B(n18640), .Z(n18639) );
  XOR U18369 ( .A(p_input[275]), .B(n18638), .Z(n18640) );
  XNOR U18370 ( .A(n18641), .B(n18642), .Z(n18638) );
  AND U18371 ( .A(n287), .B(n18643), .Z(n18642) );
  XOR U18372 ( .A(n18644), .B(n18645), .Z(n18636) );
  AND U18373 ( .A(n291), .B(n18635), .Z(n18645) );
  XNOR U18374 ( .A(n18646), .B(n18633), .Z(n18635) );
  XOR U18375 ( .A(n18647), .B(n18648), .Z(n18633) );
  AND U18376 ( .A(n314), .B(n18649), .Z(n18648) );
  IV U18377 ( .A(n18644), .Z(n18646) );
  XOR U18378 ( .A(n18650), .B(n18651), .Z(n18644) );
  AND U18379 ( .A(n298), .B(n18643), .Z(n18651) );
  XNOR U18380 ( .A(n18641), .B(n18650), .Z(n18643) );
  XNOR U18381 ( .A(n18652), .B(n18653), .Z(n18641) );
  AND U18382 ( .A(n302), .B(n18654), .Z(n18653) );
  XOR U18383 ( .A(p_input[307]), .B(n18652), .Z(n18654) );
  XNOR U18384 ( .A(n18655), .B(n18656), .Z(n18652) );
  AND U18385 ( .A(n306), .B(n18657), .Z(n18656) );
  XOR U18386 ( .A(n18658), .B(n18659), .Z(n18650) );
  AND U18387 ( .A(n310), .B(n18649), .Z(n18659) );
  XNOR U18388 ( .A(n18660), .B(n18647), .Z(n18649) );
  XOR U18389 ( .A(n18661), .B(n18662), .Z(n18647) );
  AND U18390 ( .A(n333), .B(n18663), .Z(n18662) );
  IV U18391 ( .A(n18658), .Z(n18660) );
  XOR U18392 ( .A(n18664), .B(n18665), .Z(n18658) );
  AND U18393 ( .A(n317), .B(n18657), .Z(n18665) );
  XNOR U18394 ( .A(n18655), .B(n18664), .Z(n18657) );
  XNOR U18395 ( .A(n18666), .B(n18667), .Z(n18655) );
  AND U18396 ( .A(n321), .B(n18668), .Z(n18667) );
  XOR U18397 ( .A(p_input[339]), .B(n18666), .Z(n18668) );
  XNOR U18398 ( .A(n18669), .B(n18670), .Z(n18666) );
  AND U18399 ( .A(n325), .B(n18671), .Z(n18670) );
  XOR U18400 ( .A(n18672), .B(n18673), .Z(n18664) );
  AND U18401 ( .A(n329), .B(n18663), .Z(n18673) );
  XNOR U18402 ( .A(n18674), .B(n18661), .Z(n18663) );
  XOR U18403 ( .A(n18675), .B(n18676), .Z(n18661) );
  AND U18404 ( .A(n352), .B(n18677), .Z(n18676) );
  IV U18405 ( .A(n18672), .Z(n18674) );
  XOR U18406 ( .A(n18678), .B(n18679), .Z(n18672) );
  AND U18407 ( .A(n336), .B(n18671), .Z(n18679) );
  XNOR U18408 ( .A(n18669), .B(n18678), .Z(n18671) );
  XNOR U18409 ( .A(n18680), .B(n18681), .Z(n18669) );
  AND U18410 ( .A(n340), .B(n18682), .Z(n18681) );
  XOR U18411 ( .A(p_input[371]), .B(n18680), .Z(n18682) );
  XNOR U18412 ( .A(n18683), .B(n18684), .Z(n18680) );
  AND U18413 ( .A(n344), .B(n18685), .Z(n18684) );
  XOR U18414 ( .A(n18686), .B(n18687), .Z(n18678) );
  AND U18415 ( .A(n348), .B(n18677), .Z(n18687) );
  XNOR U18416 ( .A(n18688), .B(n18675), .Z(n18677) );
  XOR U18417 ( .A(n18689), .B(n18690), .Z(n18675) );
  AND U18418 ( .A(n371), .B(n18691), .Z(n18690) );
  IV U18419 ( .A(n18686), .Z(n18688) );
  XOR U18420 ( .A(n18692), .B(n18693), .Z(n18686) );
  AND U18421 ( .A(n355), .B(n18685), .Z(n18693) );
  XNOR U18422 ( .A(n18683), .B(n18692), .Z(n18685) );
  XNOR U18423 ( .A(n18694), .B(n18695), .Z(n18683) );
  AND U18424 ( .A(n359), .B(n18696), .Z(n18695) );
  XOR U18425 ( .A(p_input[403]), .B(n18694), .Z(n18696) );
  XNOR U18426 ( .A(n18697), .B(n18698), .Z(n18694) );
  AND U18427 ( .A(n363), .B(n18699), .Z(n18698) );
  XOR U18428 ( .A(n18700), .B(n18701), .Z(n18692) );
  AND U18429 ( .A(n367), .B(n18691), .Z(n18701) );
  XNOR U18430 ( .A(n18702), .B(n18689), .Z(n18691) );
  XOR U18431 ( .A(n18703), .B(n18704), .Z(n18689) );
  AND U18432 ( .A(n390), .B(n18705), .Z(n18704) );
  IV U18433 ( .A(n18700), .Z(n18702) );
  XOR U18434 ( .A(n18706), .B(n18707), .Z(n18700) );
  AND U18435 ( .A(n374), .B(n18699), .Z(n18707) );
  XNOR U18436 ( .A(n18697), .B(n18706), .Z(n18699) );
  XNOR U18437 ( .A(n18708), .B(n18709), .Z(n18697) );
  AND U18438 ( .A(n378), .B(n18710), .Z(n18709) );
  XOR U18439 ( .A(p_input[435]), .B(n18708), .Z(n18710) );
  XNOR U18440 ( .A(n18711), .B(n18712), .Z(n18708) );
  AND U18441 ( .A(n382), .B(n18713), .Z(n18712) );
  XOR U18442 ( .A(n18714), .B(n18715), .Z(n18706) );
  AND U18443 ( .A(n386), .B(n18705), .Z(n18715) );
  XNOR U18444 ( .A(n18716), .B(n18703), .Z(n18705) );
  XOR U18445 ( .A(n18717), .B(n18718), .Z(n18703) );
  AND U18446 ( .A(n409), .B(n18719), .Z(n18718) );
  IV U18447 ( .A(n18714), .Z(n18716) );
  XOR U18448 ( .A(n18720), .B(n18721), .Z(n18714) );
  AND U18449 ( .A(n393), .B(n18713), .Z(n18721) );
  XNOR U18450 ( .A(n18711), .B(n18720), .Z(n18713) );
  XNOR U18451 ( .A(n18722), .B(n18723), .Z(n18711) );
  AND U18452 ( .A(n397), .B(n18724), .Z(n18723) );
  XOR U18453 ( .A(p_input[467]), .B(n18722), .Z(n18724) );
  XNOR U18454 ( .A(n18725), .B(n18726), .Z(n18722) );
  AND U18455 ( .A(n401), .B(n18727), .Z(n18726) );
  XOR U18456 ( .A(n18728), .B(n18729), .Z(n18720) );
  AND U18457 ( .A(n405), .B(n18719), .Z(n18729) );
  XNOR U18458 ( .A(n18730), .B(n18717), .Z(n18719) );
  XOR U18459 ( .A(n18731), .B(n18732), .Z(n18717) );
  AND U18460 ( .A(n428), .B(n18733), .Z(n18732) );
  IV U18461 ( .A(n18728), .Z(n18730) );
  XOR U18462 ( .A(n18734), .B(n18735), .Z(n18728) );
  AND U18463 ( .A(n412), .B(n18727), .Z(n18735) );
  XNOR U18464 ( .A(n18725), .B(n18734), .Z(n18727) );
  XNOR U18465 ( .A(n18736), .B(n18737), .Z(n18725) );
  AND U18466 ( .A(n416), .B(n18738), .Z(n18737) );
  XOR U18467 ( .A(p_input[499]), .B(n18736), .Z(n18738) );
  XNOR U18468 ( .A(n18739), .B(n18740), .Z(n18736) );
  AND U18469 ( .A(n420), .B(n18741), .Z(n18740) );
  XOR U18470 ( .A(n18742), .B(n18743), .Z(n18734) );
  AND U18471 ( .A(n424), .B(n18733), .Z(n18743) );
  XNOR U18472 ( .A(n18744), .B(n18731), .Z(n18733) );
  XOR U18473 ( .A(n18745), .B(n18746), .Z(n18731) );
  AND U18474 ( .A(n447), .B(n18747), .Z(n18746) );
  IV U18475 ( .A(n18742), .Z(n18744) );
  XOR U18476 ( .A(n18748), .B(n18749), .Z(n18742) );
  AND U18477 ( .A(n431), .B(n18741), .Z(n18749) );
  XNOR U18478 ( .A(n18739), .B(n18748), .Z(n18741) );
  XNOR U18479 ( .A(n18750), .B(n18751), .Z(n18739) );
  AND U18480 ( .A(n435), .B(n18752), .Z(n18751) );
  XOR U18481 ( .A(p_input[531]), .B(n18750), .Z(n18752) );
  XNOR U18482 ( .A(n18753), .B(n18754), .Z(n18750) );
  AND U18483 ( .A(n439), .B(n18755), .Z(n18754) );
  XOR U18484 ( .A(n18756), .B(n18757), .Z(n18748) );
  AND U18485 ( .A(n443), .B(n18747), .Z(n18757) );
  XNOR U18486 ( .A(n18758), .B(n18745), .Z(n18747) );
  XOR U18487 ( .A(n18759), .B(n18760), .Z(n18745) );
  AND U18488 ( .A(n466), .B(n18761), .Z(n18760) );
  IV U18489 ( .A(n18756), .Z(n18758) );
  XOR U18490 ( .A(n18762), .B(n18763), .Z(n18756) );
  AND U18491 ( .A(n450), .B(n18755), .Z(n18763) );
  XNOR U18492 ( .A(n18753), .B(n18762), .Z(n18755) );
  XNOR U18493 ( .A(n18764), .B(n18765), .Z(n18753) );
  AND U18494 ( .A(n454), .B(n18766), .Z(n18765) );
  XOR U18495 ( .A(p_input[563]), .B(n18764), .Z(n18766) );
  XNOR U18496 ( .A(n18767), .B(n18768), .Z(n18764) );
  AND U18497 ( .A(n458), .B(n18769), .Z(n18768) );
  XOR U18498 ( .A(n18770), .B(n18771), .Z(n18762) );
  AND U18499 ( .A(n462), .B(n18761), .Z(n18771) );
  XNOR U18500 ( .A(n18772), .B(n18759), .Z(n18761) );
  XOR U18501 ( .A(n18773), .B(n18774), .Z(n18759) );
  AND U18502 ( .A(n485), .B(n18775), .Z(n18774) );
  IV U18503 ( .A(n18770), .Z(n18772) );
  XOR U18504 ( .A(n18776), .B(n18777), .Z(n18770) );
  AND U18505 ( .A(n469), .B(n18769), .Z(n18777) );
  XNOR U18506 ( .A(n18767), .B(n18776), .Z(n18769) );
  XNOR U18507 ( .A(n18778), .B(n18779), .Z(n18767) );
  AND U18508 ( .A(n473), .B(n18780), .Z(n18779) );
  XOR U18509 ( .A(p_input[595]), .B(n18778), .Z(n18780) );
  XNOR U18510 ( .A(n18781), .B(n18782), .Z(n18778) );
  AND U18511 ( .A(n477), .B(n18783), .Z(n18782) );
  XOR U18512 ( .A(n18784), .B(n18785), .Z(n18776) );
  AND U18513 ( .A(n481), .B(n18775), .Z(n18785) );
  XNOR U18514 ( .A(n18786), .B(n18773), .Z(n18775) );
  XOR U18515 ( .A(n18787), .B(n18788), .Z(n18773) );
  AND U18516 ( .A(n504), .B(n18789), .Z(n18788) );
  IV U18517 ( .A(n18784), .Z(n18786) );
  XOR U18518 ( .A(n18790), .B(n18791), .Z(n18784) );
  AND U18519 ( .A(n488), .B(n18783), .Z(n18791) );
  XNOR U18520 ( .A(n18781), .B(n18790), .Z(n18783) );
  XNOR U18521 ( .A(n18792), .B(n18793), .Z(n18781) );
  AND U18522 ( .A(n492), .B(n18794), .Z(n18793) );
  XOR U18523 ( .A(p_input[627]), .B(n18792), .Z(n18794) );
  XNOR U18524 ( .A(n18795), .B(n18796), .Z(n18792) );
  AND U18525 ( .A(n496), .B(n18797), .Z(n18796) );
  XOR U18526 ( .A(n18798), .B(n18799), .Z(n18790) );
  AND U18527 ( .A(n500), .B(n18789), .Z(n18799) );
  XNOR U18528 ( .A(n18800), .B(n18787), .Z(n18789) );
  XOR U18529 ( .A(n18801), .B(n18802), .Z(n18787) );
  AND U18530 ( .A(n523), .B(n18803), .Z(n18802) );
  IV U18531 ( .A(n18798), .Z(n18800) );
  XOR U18532 ( .A(n18804), .B(n18805), .Z(n18798) );
  AND U18533 ( .A(n507), .B(n18797), .Z(n18805) );
  XNOR U18534 ( .A(n18795), .B(n18804), .Z(n18797) );
  XNOR U18535 ( .A(n18806), .B(n18807), .Z(n18795) );
  AND U18536 ( .A(n511), .B(n18808), .Z(n18807) );
  XOR U18537 ( .A(p_input[659]), .B(n18806), .Z(n18808) );
  XNOR U18538 ( .A(n18809), .B(n18810), .Z(n18806) );
  AND U18539 ( .A(n515), .B(n18811), .Z(n18810) );
  XOR U18540 ( .A(n18812), .B(n18813), .Z(n18804) );
  AND U18541 ( .A(n519), .B(n18803), .Z(n18813) );
  XNOR U18542 ( .A(n18814), .B(n18801), .Z(n18803) );
  XOR U18543 ( .A(n18815), .B(n18816), .Z(n18801) );
  AND U18544 ( .A(n542), .B(n18817), .Z(n18816) );
  IV U18545 ( .A(n18812), .Z(n18814) );
  XOR U18546 ( .A(n18818), .B(n18819), .Z(n18812) );
  AND U18547 ( .A(n526), .B(n18811), .Z(n18819) );
  XNOR U18548 ( .A(n18809), .B(n18818), .Z(n18811) );
  XNOR U18549 ( .A(n18820), .B(n18821), .Z(n18809) );
  AND U18550 ( .A(n530), .B(n18822), .Z(n18821) );
  XOR U18551 ( .A(p_input[691]), .B(n18820), .Z(n18822) );
  XNOR U18552 ( .A(n18823), .B(n18824), .Z(n18820) );
  AND U18553 ( .A(n534), .B(n18825), .Z(n18824) );
  XOR U18554 ( .A(n18826), .B(n18827), .Z(n18818) );
  AND U18555 ( .A(n538), .B(n18817), .Z(n18827) );
  XNOR U18556 ( .A(n18828), .B(n18815), .Z(n18817) );
  XOR U18557 ( .A(n18829), .B(n18830), .Z(n18815) );
  AND U18558 ( .A(n561), .B(n18831), .Z(n18830) );
  IV U18559 ( .A(n18826), .Z(n18828) );
  XOR U18560 ( .A(n18832), .B(n18833), .Z(n18826) );
  AND U18561 ( .A(n545), .B(n18825), .Z(n18833) );
  XNOR U18562 ( .A(n18823), .B(n18832), .Z(n18825) );
  XNOR U18563 ( .A(n18834), .B(n18835), .Z(n18823) );
  AND U18564 ( .A(n549), .B(n18836), .Z(n18835) );
  XOR U18565 ( .A(p_input[723]), .B(n18834), .Z(n18836) );
  XNOR U18566 ( .A(n18837), .B(n18838), .Z(n18834) );
  AND U18567 ( .A(n553), .B(n18839), .Z(n18838) );
  XOR U18568 ( .A(n18840), .B(n18841), .Z(n18832) );
  AND U18569 ( .A(n557), .B(n18831), .Z(n18841) );
  XNOR U18570 ( .A(n18842), .B(n18829), .Z(n18831) );
  XOR U18571 ( .A(n18843), .B(n18844), .Z(n18829) );
  AND U18572 ( .A(n580), .B(n18845), .Z(n18844) );
  IV U18573 ( .A(n18840), .Z(n18842) );
  XOR U18574 ( .A(n18846), .B(n18847), .Z(n18840) );
  AND U18575 ( .A(n564), .B(n18839), .Z(n18847) );
  XNOR U18576 ( .A(n18837), .B(n18846), .Z(n18839) );
  XNOR U18577 ( .A(n18848), .B(n18849), .Z(n18837) );
  AND U18578 ( .A(n568), .B(n18850), .Z(n18849) );
  XOR U18579 ( .A(p_input[755]), .B(n18848), .Z(n18850) );
  XNOR U18580 ( .A(n18851), .B(n18852), .Z(n18848) );
  AND U18581 ( .A(n572), .B(n18853), .Z(n18852) );
  XOR U18582 ( .A(n18854), .B(n18855), .Z(n18846) );
  AND U18583 ( .A(n576), .B(n18845), .Z(n18855) );
  XNOR U18584 ( .A(n18856), .B(n18843), .Z(n18845) );
  XOR U18585 ( .A(n18857), .B(n18858), .Z(n18843) );
  AND U18586 ( .A(n599), .B(n18859), .Z(n18858) );
  IV U18587 ( .A(n18854), .Z(n18856) );
  XOR U18588 ( .A(n18860), .B(n18861), .Z(n18854) );
  AND U18589 ( .A(n583), .B(n18853), .Z(n18861) );
  XNOR U18590 ( .A(n18851), .B(n18860), .Z(n18853) );
  XNOR U18591 ( .A(n18862), .B(n18863), .Z(n18851) );
  AND U18592 ( .A(n587), .B(n18864), .Z(n18863) );
  XOR U18593 ( .A(p_input[787]), .B(n18862), .Z(n18864) );
  XNOR U18594 ( .A(n18865), .B(n18866), .Z(n18862) );
  AND U18595 ( .A(n591), .B(n18867), .Z(n18866) );
  XOR U18596 ( .A(n18868), .B(n18869), .Z(n18860) );
  AND U18597 ( .A(n595), .B(n18859), .Z(n18869) );
  XNOR U18598 ( .A(n18870), .B(n18857), .Z(n18859) );
  XOR U18599 ( .A(n18871), .B(n18872), .Z(n18857) );
  AND U18600 ( .A(n618), .B(n18873), .Z(n18872) );
  IV U18601 ( .A(n18868), .Z(n18870) );
  XOR U18602 ( .A(n18874), .B(n18875), .Z(n18868) );
  AND U18603 ( .A(n602), .B(n18867), .Z(n18875) );
  XNOR U18604 ( .A(n18865), .B(n18874), .Z(n18867) );
  XNOR U18605 ( .A(n18876), .B(n18877), .Z(n18865) );
  AND U18606 ( .A(n606), .B(n18878), .Z(n18877) );
  XOR U18607 ( .A(p_input[819]), .B(n18876), .Z(n18878) );
  XNOR U18608 ( .A(n18879), .B(n18880), .Z(n18876) );
  AND U18609 ( .A(n610), .B(n18881), .Z(n18880) );
  XOR U18610 ( .A(n18882), .B(n18883), .Z(n18874) );
  AND U18611 ( .A(n614), .B(n18873), .Z(n18883) );
  XNOR U18612 ( .A(n18884), .B(n18871), .Z(n18873) );
  XOR U18613 ( .A(n18885), .B(n18886), .Z(n18871) );
  AND U18614 ( .A(n637), .B(n18887), .Z(n18886) );
  IV U18615 ( .A(n18882), .Z(n18884) );
  XOR U18616 ( .A(n18888), .B(n18889), .Z(n18882) );
  AND U18617 ( .A(n621), .B(n18881), .Z(n18889) );
  XNOR U18618 ( .A(n18879), .B(n18888), .Z(n18881) );
  XNOR U18619 ( .A(n18890), .B(n18891), .Z(n18879) );
  AND U18620 ( .A(n625), .B(n18892), .Z(n18891) );
  XOR U18621 ( .A(p_input[851]), .B(n18890), .Z(n18892) );
  XNOR U18622 ( .A(n18893), .B(n18894), .Z(n18890) );
  AND U18623 ( .A(n629), .B(n18895), .Z(n18894) );
  XOR U18624 ( .A(n18896), .B(n18897), .Z(n18888) );
  AND U18625 ( .A(n633), .B(n18887), .Z(n18897) );
  XNOR U18626 ( .A(n18898), .B(n18885), .Z(n18887) );
  XOR U18627 ( .A(n18899), .B(n18900), .Z(n18885) );
  AND U18628 ( .A(n656), .B(n18901), .Z(n18900) );
  IV U18629 ( .A(n18896), .Z(n18898) );
  XOR U18630 ( .A(n18902), .B(n18903), .Z(n18896) );
  AND U18631 ( .A(n640), .B(n18895), .Z(n18903) );
  XNOR U18632 ( .A(n18893), .B(n18902), .Z(n18895) );
  XNOR U18633 ( .A(n18904), .B(n18905), .Z(n18893) );
  AND U18634 ( .A(n644), .B(n18906), .Z(n18905) );
  XOR U18635 ( .A(p_input[883]), .B(n18904), .Z(n18906) );
  XNOR U18636 ( .A(n18907), .B(n18908), .Z(n18904) );
  AND U18637 ( .A(n648), .B(n18909), .Z(n18908) );
  XOR U18638 ( .A(n18910), .B(n18911), .Z(n18902) );
  AND U18639 ( .A(n652), .B(n18901), .Z(n18911) );
  XNOR U18640 ( .A(n18912), .B(n18899), .Z(n18901) );
  XOR U18641 ( .A(n18913), .B(n18914), .Z(n18899) );
  AND U18642 ( .A(n675), .B(n18915), .Z(n18914) );
  IV U18643 ( .A(n18910), .Z(n18912) );
  XOR U18644 ( .A(n18916), .B(n18917), .Z(n18910) );
  AND U18645 ( .A(n659), .B(n18909), .Z(n18917) );
  XNOR U18646 ( .A(n18907), .B(n18916), .Z(n18909) );
  XNOR U18647 ( .A(n18918), .B(n18919), .Z(n18907) );
  AND U18648 ( .A(n663), .B(n18920), .Z(n18919) );
  XOR U18649 ( .A(p_input[915]), .B(n18918), .Z(n18920) );
  XNOR U18650 ( .A(n18921), .B(n18922), .Z(n18918) );
  AND U18651 ( .A(n667), .B(n18923), .Z(n18922) );
  XOR U18652 ( .A(n18924), .B(n18925), .Z(n18916) );
  AND U18653 ( .A(n671), .B(n18915), .Z(n18925) );
  XNOR U18654 ( .A(n18926), .B(n18913), .Z(n18915) );
  XOR U18655 ( .A(n18927), .B(n18928), .Z(n18913) );
  AND U18656 ( .A(n694), .B(n18929), .Z(n18928) );
  IV U18657 ( .A(n18924), .Z(n18926) );
  XOR U18658 ( .A(n18930), .B(n18931), .Z(n18924) );
  AND U18659 ( .A(n678), .B(n18923), .Z(n18931) );
  XNOR U18660 ( .A(n18921), .B(n18930), .Z(n18923) );
  XNOR U18661 ( .A(n18932), .B(n18933), .Z(n18921) );
  AND U18662 ( .A(n682), .B(n18934), .Z(n18933) );
  XOR U18663 ( .A(p_input[947]), .B(n18932), .Z(n18934) );
  XNOR U18664 ( .A(n18935), .B(n18936), .Z(n18932) );
  AND U18665 ( .A(n686), .B(n18937), .Z(n18936) );
  XOR U18666 ( .A(n18938), .B(n18939), .Z(n18930) );
  AND U18667 ( .A(n690), .B(n18929), .Z(n18939) );
  XNOR U18668 ( .A(n18940), .B(n18927), .Z(n18929) );
  XOR U18669 ( .A(n18941), .B(n18942), .Z(n18927) );
  AND U18670 ( .A(n713), .B(n18943), .Z(n18942) );
  IV U18671 ( .A(n18938), .Z(n18940) );
  XOR U18672 ( .A(n18944), .B(n18945), .Z(n18938) );
  AND U18673 ( .A(n697), .B(n18937), .Z(n18945) );
  XNOR U18674 ( .A(n18935), .B(n18944), .Z(n18937) );
  XNOR U18675 ( .A(n18946), .B(n18947), .Z(n18935) );
  AND U18676 ( .A(n701), .B(n18948), .Z(n18947) );
  XOR U18677 ( .A(p_input[979]), .B(n18946), .Z(n18948) );
  XNOR U18678 ( .A(n18949), .B(n18950), .Z(n18946) );
  AND U18679 ( .A(n705), .B(n18951), .Z(n18950) );
  XOR U18680 ( .A(n18952), .B(n18953), .Z(n18944) );
  AND U18681 ( .A(n709), .B(n18943), .Z(n18953) );
  XNOR U18682 ( .A(n18954), .B(n18941), .Z(n18943) );
  XOR U18683 ( .A(n18955), .B(n18956), .Z(n18941) );
  AND U18684 ( .A(n732), .B(n18957), .Z(n18956) );
  IV U18685 ( .A(n18952), .Z(n18954) );
  XOR U18686 ( .A(n18958), .B(n18959), .Z(n18952) );
  AND U18687 ( .A(n716), .B(n18951), .Z(n18959) );
  XNOR U18688 ( .A(n18949), .B(n18958), .Z(n18951) );
  XNOR U18689 ( .A(n18960), .B(n18961), .Z(n18949) );
  AND U18690 ( .A(n720), .B(n18962), .Z(n18961) );
  XOR U18691 ( .A(p_input[1011]), .B(n18960), .Z(n18962) );
  XNOR U18692 ( .A(n18963), .B(n18964), .Z(n18960) );
  AND U18693 ( .A(n724), .B(n18965), .Z(n18964) );
  XOR U18694 ( .A(n18966), .B(n18967), .Z(n18958) );
  AND U18695 ( .A(n728), .B(n18957), .Z(n18967) );
  XNOR U18696 ( .A(n18968), .B(n18955), .Z(n18957) );
  XOR U18697 ( .A(n18969), .B(n18970), .Z(n18955) );
  AND U18698 ( .A(n751), .B(n18971), .Z(n18970) );
  IV U18699 ( .A(n18966), .Z(n18968) );
  XOR U18700 ( .A(n18972), .B(n18973), .Z(n18966) );
  AND U18701 ( .A(n735), .B(n18965), .Z(n18973) );
  XNOR U18702 ( .A(n18963), .B(n18972), .Z(n18965) );
  XNOR U18703 ( .A(n18974), .B(n18975), .Z(n18963) );
  AND U18704 ( .A(n739), .B(n18976), .Z(n18975) );
  XOR U18705 ( .A(p_input[1043]), .B(n18974), .Z(n18976) );
  XNOR U18706 ( .A(n18977), .B(n18978), .Z(n18974) );
  AND U18707 ( .A(n743), .B(n18979), .Z(n18978) );
  XOR U18708 ( .A(n18980), .B(n18981), .Z(n18972) );
  AND U18709 ( .A(n747), .B(n18971), .Z(n18981) );
  XNOR U18710 ( .A(n18982), .B(n18969), .Z(n18971) );
  XOR U18711 ( .A(n18983), .B(n18984), .Z(n18969) );
  AND U18712 ( .A(n770), .B(n18985), .Z(n18984) );
  IV U18713 ( .A(n18980), .Z(n18982) );
  XOR U18714 ( .A(n18986), .B(n18987), .Z(n18980) );
  AND U18715 ( .A(n754), .B(n18979), .Z(n18987) );
  XNOR U18716 ( .A(n18977), .B(n18986), .Z(n18979) );
  XNOR U18717 ( .A(n18988), .B(n18989), .Z(n18977) );
  AND U18718 ( .A(n758), .B(n18990), .Z(n18989) );
  XOR U18719 ( .A(p_input[1075]), .B(n18988), .Z(n18990) );
  XNOR U18720 ( .A(n18991), .B(n18992), .Z(n18988) );
  AND U18721 ( .A(n762), .B(n18993), .Z(n18992) );
  XOR U18722 ( .A(n18994), .B(n18995), .Z(n18986) );
  AND U18723 ( .A(n766), .B(n18985), .Z(n18995) );
  XNOR U18724 ( .A(n18996), .B(n18983), .Z(n18985) );
  XOR U18725 ( .A(n18997), .B(n18998), .Z(n18983) );
  AND U18726 ( .A(n789), .B(n18999), .Z(n18998) );
  IV U18727 ( .A(n18994), .Z(n18996) );
  XOR U18728 ( .A(n19000), .B(n19001), .Z(n18994) );
  AND U18729 ( .A(n773), .B(n18993), .Z(n19001) );
  XNOR U18730 ( .A(n18991), .B(n19000), .Z(n18993) );
  XNOR U18731 ( .A(n19002), .B(n19003), .Z(n18991) );
  AND U18732 ( .A(n777), .B(n19004), .Z(n19003) );
  XOR U18733 ( .A(p_input[1107]), .B(n19002), .Z(n19004) );
  XNOR U18734 ( .A(n19005), .B(n19006), .Z(n19002) );
  AND U18735 ( .A(n781), .B(n19007), .Z(n19006) );
  XOR U18736 ( .A(n19008), .B(n19009), .Z(n19000) );
  AND U18737 ( .A(n785), .B(n18999), .Z(n19009) );
  XNOR U18738 ( .A(n19010), .B(n18997), .Z(n18999) );
  XOR U18739 ( .A(n19011), .B(n19012), .Z(n18997) );
  AND U18740 ( .A(n808), .B(n19013), .Z(n19012) );
  IV U18741 ( .A(n19008), .Z(n19010) );
  XOR U18742 ( .A(n19014), .B(n19015), .Z(n19008) );
  AND U18743 ( .A(n792), .B(n19007), .Z(n19015) );
  XNOR U18744 ( .A(n19005), .B(n19014), .Z(n19007) );
  XNOR U18745 ( .A(n19016), .B(n19017), .Z(n19005) );
  AND U18746 ( .A(n796), .B(n19018), .Z(n19017) );
  XOR U18747 ( .A(p_input[1139]), .B(n19016), .Z(n19018) );
  XNOR U18748 ( .A(n19019), .B(n19020), .Z(n19016) );
  AND U18749 ( .A(n800), .B(n19021), .Z(n19020) );
  XOR U18750 ( .A(n19022), .B(n19023), .Z(n19014) );
  AND U18751 ( .A(n804), .B(n19013), .Z(n19023) );
  XNOR U18752 ( .A(n19024), .B(n19011), .Z(n19013) );
  XOR U18753 ( .A(n19025), .B(n19026), .Z(n19011) );
  AND U18754 ( .A(n827), .B(n19027), .Z(n19026) );
  IV U18755 ( .A(n19022), .Z(n19024) );
  XOR U18756 ( .A(n19028), .B(n19029), .Z(n19022) );
  AND U18757 ( .A(n811), .B(n19021), .Z(n19029) );
  XNOR U18758 ( .A(n19019), .B(n19028), .Z(n19021) );
  XNOR U18759 ( .A(n19030), .B(n19031), .Z(n19019) );
  AND U18760 ( .A(n815), .B(n19032), .Z(n19031) );
  XOR U18761 ( .A(p_input[1171]), .B(n19030), .Z(n19032) );
  XNOR U18762 ( .A(n19033), .B(n19034), .Z(n19030) );
  AND U18763 ( .A(n819), .B(n19035), .Z(n19034) );
  XOR U18764 ( .A(n19036), .B(n19037), .Z(n19028) );
  AND U18765 ( .A(n823), .B(n19027), .Z(n19037) );
  XNOR U18766 ( .A(n19038), .B(n19025), .Z(n19027) );
  XOR U18767 ( .A(n19039), .B(n19040), .Z(n19025) );
  AND U18768 ( .A(n846), .B(n19041), .Z(n19040) );
  IV U18769 ( .A(n19036), .Z(n19038) );
  XOR U18770 ( .A(n19042), .B(n19043), .Z(n19036) );
  AND U18771 ( .A(n830), .B(n19035), .Z(n19043) );
  XNOR U18772 ( .A(n19033), .B(n19042), .Z(n19035) );
  XNOR U18773 ( .A(n19044), .B(n19045), .Z(n19033) );
  AND U18774 ( .A(n834), .B(n19046), .Z(n19045) );
  XOR U18775 ( .A(p_input[1203]), .B(n19044), .Z(n19046) );
  XNOR U18776 ( .A(n19047), .B(n19048), .Z(n19044) );
  AND U18777 ( .A(n838), .B(n19049), .Z(n19048) );
  XOR U18778 ( .A(n19050), .B(n19051), .Z(n19042) );
  AND U18779 ( .A(n842), .B(n19041), .Z(n19051) );
  XNOR U18780 ( .A(n19052), .B(n19039), .Z(n19041) );
  XOR U18781 ( .A(n19053), .B(n19054), .Z(n19039) );
  AND U18782 ( .A(n865), .B(n19055), .Z(n19054) );
  IV U18783 ( .A(n19050), .Z(n19052) );
  XOR U18784 ( .A(n19056), .B(n19057), .Z(n19050) );
  AND U18785 ( .A(n849), .B(n19049), .Z(n19057) );
  XNOR U18786 ( .A(n19047), .B(n19056), .Z(n19049) );
  XNOR U18787 ( .A(n19058), .B(n19059), .Z(n19047) );
  AND U18788 ( .A(n853), .B(n19060), .Z(n19059) );
  XOR U18789 ( .A(p_input[1235]), .B(n19058), .Z(n19060) );
  XNOR U18790 ( .A(n19061), .B(n19062), .Z(n19058) );
  AND U18791 ( .A(n857), .B(n19063), .Z(n19062) );
  XOR U18792 ( .A(n19064), .B(n19065), .Z(n19056) );
  AND U18793 ( .A(n861), .B(n19055), .Z(n19065) );
  XNOR U18794 ( .A(n19066), .B(n19053), .Z(n19055) );
  XOR U18795 ( .A(n19067), .B(n19068), .Z(n19053) );
  AND U18796 ( .A(n884), .B(n19069), .Z(n19068) );
  IV U18797 ( .A(n19064), .Z(n19066) );
  XOR U18798 ( .A(n19070), .B(n19071), .Z(n19064) );
  AND U18799 ( .A(n868), .B(n19063), .Z(n19071) );
  XNOR U18800 ( .A(n19061), .B(n19070), .Z(n19063) );
  XNOR U18801 ( .A(n19072), .B(n19073), .Z(n19061) );
  AND U18802 ( .A(n872), .B(n19074), .Z(n19073) );
  XOR U18803 ( .A(p_input[1267]), .B(n19072), .Z(n19074) );
  XNOR U18804 ( .A(n19075), .B(n19076), .Z(n19072) );
  AND U18805 ( .A(n876), .B(n19077), .Z(n19076) );
  XOR U18806 ( .A(n19078), .B(n19079), .Z(n19070) );
  AND U18807 ( .A(n880), .B(n19069), .Z(n19079) );
  XNOR U18808 ( .A(n19080), .B(n19067), .Z(n19069) );
  XOR U18809 ( .A(n19081), .B(n19082), .Z(n19067) );
  AND U18810 ( .A(n903), .B(n19083), .Z(n19082) );
  IV U18811 ( .A(n19078), .Z(n19080) );
  XOR U18812 ( .A(n19084), .B(n19085), .Z(n19078) );
  AND U18813 ( .A(n887), .B(n19077), .Z(n19085) );
  XNOR U18814 ( .A(n19075), .B(n19084), .Z(n19077) );
  XNOR U18815 ( .A(n19086), .B(n19087), .Z(n19075) );
  AND U18816 ( .A(n891), .B(n19088), .Z(n19087) );
  XOR U18817 ( .A(p_input[1299]), .B(n19086), .Z(n19088) );
  XNOR U18818 ( .A(n19089), .B(n19090), .Z(n19086) );
  AND U18819 ( .A(n895), .B(n19091), .Z(n19090) );
  XOR U18820 ( .A(n19092), .B(n19093), .Z(n19084) );
  AND U18821 ( .A(n899), .B(n19083), .Z(n19093) );
  XNOR U18822 ( .A(n19094), .B(n19081), .Z(n19083) );
  XOR U18823 ( .A(n19095), .B(n19096), .Z(n19081) );
  AND U18824 ( .A(n922), .B(n19097), .Z(n19096) );
  IV U18825 ( .A(n19092), .Z(n19094) );
  XOR U18826 ( .A(n19098), .B(n19099), .Z(n19092) );
  AND U18827 ( .A(n906), .B(n19091), .Z(n19099) );
  XNOR U18828 ( .A(n19089), .B(n19098), .Z(n19091) );
  XNOR U18829 ( .A(n19100), .B(n19101), .Z(n19089) );
  AND U18830 ( .A(n910), .B(n19102), .Z(n19101) );
  XOR U18831 ( .A(p_input[1331]), .B(n19100), .Z(n19102) );
  XNOR U18832 ( .A(n19103), .B(n19104), .Z(n19100) );
  AND U18833 ( .A(n914), .B(n19105), .Z(n19104) );
  XOR U18834 ( .A(n19106), .B(n19107), .Z(n19098) );
  AND U18835 ( .A(n918), .B(n19097), .Z(n19107) );
  XNOR U18836 ( .A(n19108), .B(n19095), .Z(n19097) );
  XOR U18837 ( .A(n19109), .B(n19110), .Z(n19095) );
  AND U18838 ( .A(n941), .B(n19111), .Z(n19110) );
  IV U18839 ( .A(n19106), .Z(n19108) );
  XOR U18840 ( .A(n19112), .B(n19113), .Z(n19106) );
  AND U18841 ( .A(n925), .B(n19105), .Z(n19113) );
  XNOR U18842 ( .A(n19103), .B(n19112), .Z(n19105) );
  XNOR U18843 ( .A(n19114), .B(n19115), .Z(n19103) );
  AND U18844 ( .A(n929), .B(n19116), .Z(n19115) );
  XOR U18845 ( .A(p_input[1363]), .B(n19114), .Z(n19116) );
  XNOR U18846 ( .A(n19117), .B(n19118), .Z(n19114) );
  AND U18847 ( .A(n933), .B(n19119), .Z(n19118) );
  XOR U18848 ( .A(n19120), .B(n19121), .Z(n19112) );
  AND U18849 ( .A(n937), .B(n19111), .Z(n19121) );
  XNOR U18850 ( .A(n19122), .B(n19109), .Z(n19111) );
  XOR U18851 ( .A(n19123), .B(n19124), .Z(n19109) );
  AND U18852 ( .A(n960), .B(n19125), .Z(n19124) );
  IV U18853 ( .A(n19120), .Z(n19122) );
  XOR U18854 ( .A(n19126), .B(n19127), .Z(n19120) );
  AND U18855 ( .A(n944), .B(n19119), .Z(n19127) );
  XNOR U18856 ( .A(n19117), .B(n19126), .Z(n19119) );
  XNOR U18857 ( .A(n19128), .B(n19129), .Z(n19117) );
  AND U18858 ( .A(n948), .B(n19130), .Z(n19129) );
  XOR U18859 ( .A(p_input[1395]), .B(n19128), .Z(n19130) );
  XNOR U18860 ( .A(n19131), .B(n19132), .Z(n19128) );
  AND U18861 ( .A(n952), .B(n19133), .Z(n19132) );
  XOR U18862 ( .A(n19134), .B(n19135), .Z(n19126) );
  AND U18863 ( .A(n956), .B(n19125), .Z(n19135) );
  XNOR U18864 ( .A(n19136), .B(n19123), .Z(n19125) );
  XOR U18865 ( .A(n19137), .B(n19138), .Z(n19123) );
  AND U18866 ( .A(n979), .B(n19139), .Z(n19138) );
  IV U18867 ( .A(n19134), .Z(n19136) );
  XOR U18868 ( .A(n19140), .B(n19141), .Z(n19134) );
  AND U18869 ( .A(n963), .B(n19133), .Z(n19141) );
  XNOR U18870 ( .A(n19131), .B(n19140), .Z(n19133) );
  XNOR U18871 ( .A(n19142), .B(n19143), .Z(n19131) );
  AND U18872 ( .A(n967), .B(n19144), .Z(n19143) );
  XOR U18873 ( .A(p_input[1427]), .B(n19142), .Z(n19144) );
  XNOR U18874 ( .A(n19145), .B(n19146), .Z(n19142) );
  AND U18875 ( .A(n971), .B(n19147), .Z(n19146) );
  XOR U18876 ( .A(n19148), .B(n19149), .Z(n19140) );
  AND U18877 ( .A(n975), .B(n19139), .Z(n19149) );
  XNOR U18878 ( .A(n19150), .B(n19137), .Z(n19139) );
  XOR U18879 ( .A(n19151), .B(n19152), .Z(n19137) );
  AND U18880 ( .A(n998), .B(n19153), .Z(n19152) );
  IV U18881 ( .A(n19148), .Z(n19150) );
  XOR U18882 ( .A(n19154), .B(n19155), .Z(n19148) );
  AND U18883 ( .A(n982), .B(n19147), .Z(n19155) );
  XNOR U18884 ( .A(n19145), .B(n19154), .Z(n19147) );
  XNOR U18885 ( .A(n19156), .B(n19157), .Z(n19145) );
  AND U18886 ( .A(n986), .B(n19158), .Z(n19157) );
  XOR U18887 ( .A(p_input[1459]), .B(n19156), .Z(n19158) );
  XNOR U18888 ( .A(n19159), .B(n19160), .Z(n19156) );
  AND U18889 ( .A(n990), .B(n19161), .Z(n19160) );
  XOR U18890 ( .A(n19162), .B(n19163), .Z(n19154) );
  AND U18891 ( .A(n994), .B(n19153), .Z(n19163) );
  XNOR U18892 ( .A(n19164), .B(n19151), .Z(n19153) );
  XOR U18893 ( .A(n19165), .B(n19166), .Z(n19151) );
  AND U18894 ( .A(n1017), .B(n19167), .Z(n19166) );
  IV U18895 ( .A(n19162), .Z(n19164) );
  XOR U18896 ( .A(n19168), .B(n19169), .Z(n19162) );
  AND U18897 ( .A(n1001), .B(n19161), .Z(n19169) );
  XNOR U18898 ( .A(n19159), .B(n19168), .Z(n19161) );
  XNOR U18899 ( .A(n19170), .B(n19171), .Z(n19159) );
  AND U18900 ( .A(n1005), .B(n19172), .Z(n19171) );
  XOR U18901 ( .A(p_input[1491]), .B(n19170), .Z(n19172) );
  XNOR U18902 ( .A(n19173), .B(n19174), .Z(n19170) );
  AND U18903 ( .A(n1009), .B(n19175), .Z(n19174) );
  XOR U18904 ( .A(n19176), .B(n19177), .Z(n19168) );
  AND U18905 ( .A(n1013), .B(n19167), .Z(n19177) );
  XNOR U18906 ( .A(n19178), .B(n19165), .Z(n19167) );
  XOR U18907 ( .A(n19179), .B(n19180), .Z(n19165) );
  AND U18908 ( .A(n1036), .B(n19181), .Z(n19180) );
  IV U18909 ( .A(n19176), .Z(n19178) );
  XOR U18910 ( .A(n19182), .B(n19183), .Z(n19176) );
  AND U18911 ( .A(n1020), .B(n19175), .Z(n19183) );
  XNOR U18912 ( .A(n19173), .B(n19182), .Z(n19175) );
  XNOR U18913 ( .A(n19184), .B(n19185), .Z(n19173) );
  AND U18914 ( .A(n1024), .B(n19186), .Z(n19185) );
  XOR U18915 ( .A(p_input[1523]), .B(n19184), .Z(n19186) );
  XNOR U18916 ( .A(n19187), .B(n19188), .Z(n19184) );
  AND U18917 ( .A(n1028), .B(n19189), .Z(n19188) );
  XOR U18918 ( .A(n19190), .B(n19191), .Z(n19182) );
  AND U18919 ( .A(n1032), .B(n19181), .Z(n19191) );
  XNOR U18920 ( .A(n19192), .B(n19179), .Z(n19181) );
  XOR U18921 ( .A(n19193), .B(n19194), .Z(n19179) );
  AND U18922 ( .A(n1055), .B(n19195), .Z(n19194) );
  IV U18923 ( .A(n19190), .Z(n19192) );
  XOR U18924 ( .A(n19196), .B(n19197), .Z(n19190) );
  AND U18925 ( .A(n1039), .B(n19189), .Z(n19197) );
  XNOR U18926 ( .A(n19187), .B(n19196), .Z(n19189) );
  XNOR U18927 ( .A(n19198), .B(n19199), .Z(n19187) );
  AND U18928 ( .A(n1043), .B(n19200), .Z(n19199) );
  XOR U18929 ( .A(p_input[1555]), .B(n19198), .Z(n19200) );
  XNOR U18930 ( .A(n19201), .B(n19202), .Z(n19198) );
  AND U18931 ( .A(n1047), .B(n19203), .Z(n19202) );
  XOR U18932 ( .A(n19204), .B(n19205), .Z(n19196) );
  AND U18933 ( .A(n1051), .B(n19195), .Z(n19205) );
  XNOR U18934 ( .A(n19206), .B(n19193), .Z(n19195) );
  XOR U18935 ( .A(n19207), .B(n19208), .Z(n19193) );
  AND U18936 ( .A(n1074), .B(n19209), .Z(n19208) );
  IV U18937 ( .A(n19204), .Z(n19206) );
  XOR U18938 ( .A(n19210), .B(n19211), .Z(n19204) );
  AND U18939 ( .A(n1058), .B(n19203), .Z(n19211) );
  XNOR U18940 ( .A(n19201), .B(n19210), .Z(n19203) );
  XNOR U18941 ( .A(n19212), .B(n19213), .Z(n19201) );
  AND U18942 ( .A(n1062), .B(n19214), .Z(n19213) );
  XOR U18943 ( .A(p_input[1587]), .B(n19212), .Z(n19214) );
  XNOR U18944 ( .A(n19215), .B(n19216), .Z(n19212) );
  AND U18945 ( .A(n1066), .B(n19217), .Z(n19216) );
  XOR U18946 ( .A(n19218), .B(n19219), .Z(n19210) );
  AND U18947 ( .A(n1070), .B(n19209), .Z(n19219) );
  XNOR U18948 ( .A(n19220), .B(n19207), .Z(n19209) );
  XOR U18949 ( .A(n19221), .B(n19222), .Z(n19207) );
  AND U18950 ( .A(n1093), .B(n19223), .Z(n19222) );
  IV U18951 ( .A(n19218), .Z(n19220) );
  XOR U18952 ( .A(n19224), .B(n19225), .Z(n19218) );
  AND U18953 ( .A(n1077), .B(n19217), .Z(n19225) );
  XNOR U18954 ( .A(n19215), .B(n19224), .Z(n19217) );
  XNOR U18955 ( .A(n19226), .B(n19227), .Z(n19215) );
  AND U18956 ( .A(n1081), .B(n19228), .Z(n19227) );
  XOR U18957 ( .A(p_input[1619]), .B(n19226), .Z(n19228) );
  XNOR U18958 ( .A(n19229), .B(n19230), .Z(n19226) );
  AND U18959 ( .A(n1085), .B(n19231), .Z(n19230) );
  XOR U18960 ( .A(n19232), .B(n19233), .Z(n19224) );
  AND U18961 ( .A(n1089), .B(n19223), .Z(n19233) );
  XNOR U18962 ( .A(n19234), .B(n19221), .Z(n19223) );
  XOR U18963 ( .A(n19235), .B(n19236), .Z(n19221) );
  AND U18964 ( .A(n1112), .B(n19237), .Z(n19236) );
  IV U18965 ( .A(n19232), .Z(n19234) );
  XOR U18966 ( .A(n19238), .B(n19239), .Z(n19232) );
  AND U18967 ( .A(n1096), .B(n19231), .Z(n19239) );
  XNOR U18968 ( .A(n19229), .B(n19238), .Z(n19231) );
  XNOR U18969 ( .A(n19240), .B(n19241), .Z(n19229) );
  AND U18970 ( .A(n1100), .B(n19242), .Z(n19241) );
  XOR U18971 ( .A(p_input[1651]), .B(n19240), .Z(n19242) );
  XNOR U18972 ( .A(n19243), .B(n19244), .Z(n19240) );
  AND U18973 ( .A(n1104), .B(n19245), .Z(n19244) );
  XOR U18974 ( .A(n19246), .B(n19247), .Z(n19238) );
  AND U18975 ( .A(n1108), .B(n19237), .Z(n19247) );
  XNOR U18976 ( .A(n19248), .B(n19235), .Z(n19237) );
  XOR U18977 ( .A(n19249), .B(n19250), .Z(n19235) );
  AND U18978 ( .A(n1131), .B(n19251), .Z(n19250) );
  IV U18979 ( .A(n19246), .Z(n19248) );
  XOR U18980 ( .A(n19252), .B(n19253), .Z(n19246) );
  AND U18981 ( .A(n1115), .B(n19245), .Z(n19253) );
  XNOR U18982 ( .A(n19243), .B(n19252), .Z(n19245) );
  XNOR U18983 ( .A(n19254), .B(n19255), .Z(n19243) );
  AND U18984 ( .A(n1119), .B(n19256), .Z(n19255) );
  XOR U18985 ( .A(p_input[1683]), .B(n19254), .Z(n19256) );
  XNOR U18986 ( .A(n19257), .B(n19258), .Z(n19254) );
  AND U18987 ( .A(n1123), .B(n19259), .Z(n19258) );
  XOR U18988 ( .A(n19260), .B(n19261), .Z(n19252) );
  AND U18989 ( .A(n1127), .B(n19251), .Z(n19261) );
  XNOR U18990 ( .A(n19262), .B(n19249), .Z(n19251) );
  XOR U18991 ( .A(n19263), .B(n19264), .Z(n19249) );
  AND U18992 ( .A(n1150), .B(n19265), .Z(n19264) );
  IV U18993 ( .A(n19260), .Z(n19262) );
  XOR U18994 ( .A(n19266), .B(n19267), .Z(n19260) );
  AND U18995 ( .A(n1134), .B(n19259), .Z(n19267) );
  XNOR U18996 ( .A(n19257), .B(n19266), .Z(n19259) );
  XNOR U18997 ( .A(n19268), .B(n19269), .Z(n19257) );
  AND U18998 ( .A(n1138), .B(n19270), .Z(n19269) );
  XOR U18999 ( .A(p_input[1715]), .B(n19268), .Z(n19270) );
  XNOR U19000 ( .A(n19271), .B(n19272), .Z(n19268) );
  AND U19001 ( .A(n1142), .B(n19273), .Z(n19272) );
  XOR U19002 ( .A(n19274), .B(n19275), .Z(n19266) );
  AND U19003 ( .A(n1146), .B(n19265), .Z(n19275) );
  XNOR U19004 ( .A(n19276), .B(n19263), .Z(n19265) );
  XOR U19005 ( .A(n19277), .B(n19278), .Z(n19263) );
  AND U19006 ( .A(n1169), .B(n19279), .Z(n19278) );
  IV U19007 ( .A(n19274), .Z(n19276) );
  XOR U19008 ( .A(n19280), .B(n19281), .Z(n19274) );
  AND U19009 ( .A(n1153), .B(n19273), .Z(n19281) );
  XNOR U19010 ( .A(n19271), .B(n19280), .Z(n19273) );
  XNOR U19011 ( .A(n19282), .B(n19283), .Z(n19271) );
  AND U19012 ( .A(n1157), .B(n19284), .Z(n19283) );
  XOR U19013 ( .A(p_input[1747]), .B(n19282), .Z(n19284) );
  XNOR U19014 ( .A(n19285), .B(n19286), .Z(n19282) );
  AND U19015 ( .A(n1161), .B(n19287), .Z(n19286) );
  XOR U19016 ( .A(n19288), .B(n19289), .Z(n19280) );
  AND U19017 ( .A(n1165), .B(n19279), .Z(n19289) );
  XNOR U19018 ( .A(n19290), .B(n19277), .Z(n19279) );
  XOR U19019 ( .A(n19291), .B(n19292), .Z(n19277) );
  AND U19020 ( .A(n1188), .B(n19293), .Z(n19292) );
  IV U19021 ( .A(n19288), .Z(n19290) );
  XOR U19022 ( .A(n19294), .B(n19295), .Z(n19288) );
  AND U19023 ( .A(n1172), .B(n19287), .Z(n19295) );
  XNOR U19024 ( .A(n19285), .B(n19294), .Z(n19287) );
  XNOR U19025 ( .A(n19296), .B(n19297), .Z(n19285) );
  AND U19026 ( .A(n1176), .B(n19298), .Z(n19297) );
  XOR U19027 ( .A(p_input[1779]), .B(n19296), .Z(n19298) );
  XNOR U19028 ( .A(n19299), .B(n19300), .Z(n19296) );
  AND U19029 ( .A(n1180), .B(n19301), .Z(n19300) );
  XOR U19030 ( .A(n19302), .B(n19303), .Z(n19294) );
  AND U19031 ( .A(n1184), .B(n19293), .Z(n19303) );
  XNOR U19032 ( .A(n19304), .B(n19291), .Z(n19293) );
  XOR U19033 ( .A(n19305), .B(n19306), .Z(n19291) );
  AND U19034 ( .A(n1207), .B(n19307), .Z(n19306) );
  IV U19035 ( .A(n19302), .Z(n19304) );
  XOR U19036 ( .A(n19308), .B(n19309), .Z(n19302) );
  AND U19037 ( .A(n1191), .B(n19301), .Z(n19309) );
  XNOR U19038 ( .A(n19299), .B(n19308), .Z(n19301) );
  XNOR U19039 ( .A(n19310), .B(n19311), .Z(n19299) );
  AND U19040 ( .A(n1195), .B(n19312), .Z(n19311) );
  XOR U19041 ( .A(p_input[1811]), .B(n19310), .Z(n19312) );
  XNOR U19042 ( .A(n19313), .B(n19314), .Z(n19310) );
  AND U19043 ( .A(n1199), .B(n19315), .Z(n19314) );
  XOR U19044 ( .A(n19316), .B(n19317), .Z(n19308) );
  AND U19045 ( .A(n1203), .B(n19307), .Z(n19317) );
  XNOR U19046 ( .A(n19318), .B(n19305), .Z(n19307) );
  XOR U19047 ( .A(n19319), .B(n19320), .Z(n19305) );
  AND U19048 ( .A(n1226), .B(n19321), .Z(n19320) );
  IV U19049 ( .A(n19316), .Z(n19318) );
  XOR U19050 ( .A(n19322), .B(n19323), .Z(n19316) );
  AND U19051 ( .A(n1210), .B(n19315), .Z(n19323) );
  XNOR U19052 ( .A(n19313), .B(n19322), .Z(n19315) );
  XNOR U19053 ( .A(n19324), .B(n19325), .Z(n19313) );
  AND U19054 ( .A(n1214), .B(n19326), .Z(n19325) );
  XOR U19055 ( .A(p_input[1843]), .B(n19324), .Z(n19326) );
  XNOR U19056 ( .A(n19327), .B(n19328), .Z(n19324) );
  AND U19057 ( .A(n1218), .B(n19329), .Z(n19328) );
  XOR U19058 ( .A(n19330), .B(n19331), .Z(n19322) );
  AND U19059 ( .A(n1222), .B(n19321), .Z(n19331) );
  XNOR U19060 ( .A(n19332), .B(n19319), .Z(n19321) );
  XOR U19061 ( .A(n19333), .B(n19334), .Z(n19319) );
  AND U19062 ( .A(n1245), .B(n19335), .Z(n19334) );
  IV U19063 ( .A(n19330), .Z(n19332) );
  XOR U19064 ( .A(n19336), .B(n19337), .Z(n19330) );
  AND U19065 ( .A(n1229), .B(n19329), .Z(n19337) );
  XNOR U19066 ( .A(n19327), .B(n19336), .Z(n19329) );
  XNOR U19067 ( .A(n19338), .B(n19339), .Z(n19327) );
  AND U19068 ( .A(n1233), .B(n19340), .Z(n19339) );
  XOR U19069 ( .A(p_input[1875]), .B(n19338), .Z(n19340) );
  XNOR U19070 ( .A(n19341), .B(n19342), .Z(n19338) );
  AND U19071 ( .A(n1237), .B(n19343), .Z(n19342) );
  XOR U19072 ( .A(n19344), .B(n19345), .Z(n19336) );
  AND U19073 ( .A(n1241), .B(n19335), .Z(n19345) );
  XNOR U19074 ( .A(n19346), .B(n19333), .Z(n19335) );
  XOR U19075 ( .A(n19347), .B(n19348), .Z(n19333) );
  AND U19076 ( .A(n1264), .B(n19349), .Z(n19348) );
  IV U19077 ( .A(n19344), .Z(n19346) );
  XOR U19078 ( .A(n19350), .B(n19351), .Z(n19344) );
  AND U19079 ( .A(n1248), .B(n19343), .Z(n19351) );
  XNOR U19080 ( .A(n19341), .B(n19350), .Z(n19343) );
  XNOR U19081 ( .A(n19352), .B(n19353), .Z(n19341) );
  AND U19082 ( .A(n1252), .B(n19354), .Z(n19353) );
  XOR U19083 ( .A(p_input[1907]), .B(n19352), .Z(n19354) );
  XNOR U19084 ( .A(n19355), .B(n19356), .Z(n19352) );
  AND U19085 ( .A(n1256), .B(n19357), .Z(n19356) );
  XOR U19086 ( .A(n19358), .B(n19359), .Z(n19350) );
  AND U19087 ( .A(n1260), .B(n19349), .Z(n19359) );
  XNOR U19088 ( .A(n19360), .B(n19347), .Z(n19349) );
  XOR U19089 ( .A(n19361), .B(n19362), .Z(n19347) );
  AND U19090 ( .A(n1282), .B(n19363), .Z(n19362) );
  IV U19091 ( .A(n19358), .Z(n19360) );
  XOR U19092 ( .A(n19364), .B(n19365), .Z(n19358) );
  AND U19093 ( .A(n1267), .B(n19357), .Z(n19365) );
  XNOR U19094 ( .A(n19355), .B(n19364), .Z(n19357) );
  XNOR U19095 ( .A(n19366), .B(n19367), .Z(n19355) );
  AND U19096 ( .A(n1271), .B(n19368), .Z(n19367) );
  XOR U19097 ( .A(p_input[1939]), .B(n19366), .Z(n19368) );
  XOR U19098 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][19] ), .B(n19369), 
        .Z(n19366) );
  AND U19099 ( .A(n1274), .B(n19370), .Z(n19369) );
  XOR U19100 ( .A(n19371), .B(n19372), .Z(n19364) );
  AND U19101 ( .A(n1278), .B(n19363), .Z(n19372) );
  XNOR U19102 ( .A(n19373), .B(n19361), .Z(n19363) );
  XOR U19103 ( .A(\knn_comb_/min_val_out[0][19] ), .B(n19374), .Z(n19361) );
  AND U19104 ( .A(n1290), .B(n19375), .Z(n19374) );
  IV U19105 ( .A(n19371), .Z(n19373) );
  XOR U19106 ( .A(n19376), .B(n19377), .Z(n19371) );
  AND U19107 ( .A(n1285), .B(n19370), .Z(n19377) );
  XOR U19108 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][19] ), .B(n19376), 
        .Z(n19370) );
  XOR U19109 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .B(n19378), 
        .Z(n19376) );
  AND U19110 ( .A(n1287), .B(n19375), .Z(n19378) );
  XOR U19111 ( .A(\knn_comb_/min_val_out[0][19] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .Z(n19375) );
  XOR U19112 ( .A(n101), .B(n19379), .Z(o[18]) );
  AND U19113 ( .A(n122), .B(n19380), .Z(n101) );
  XOR U19114 ( .A(n102), .B(n19379), .Z(n19380) );
  XOR U19115 ( .A(n19381), .B(n19382), .Z(n19379) );
  AND U19116 ( .A(n142), .B(n19383), .Z(n19382) );
  XOR U19117 ( .A(n19384), .B(n31), .Z(n102) );
  AND U19118 ( .A(n125), .B(n19385), .Z(n31) );
  XOR U19119 ( .A(n32), .B(n19384), .Z(n19385) );
  XOR U19120 ( .A(n19386), .B(n19387), .Z(n32) );
  AND U19121 ( .A(n130), .B(n19388), .Z(n19387) );
  XOR U19122 ( .A(p_input[18]), .B(n19386), .Z(n19388) );
  XNOR U19123 ( .A(n19389), .B(n19390), .Z(n19386) );
  AND U19124 ( .A(n134), .B(n19391), .Z(n19390) );
  XOR U19125 ( .A(n19392), .B(n19393), .Z(n19384) );
  AND U19126 ( .A(n138), .B(n19383), .Z(n19393) );
  XNOR U19127 ( .A(n19394), .B(n19381), .Z(n19383) );
  XOR U19128 ( .A(n19395), .B(n19396), .Z(n19381) );
  AND U19129 ( .A(n162), .B(n19397), .Z(n19396) );
  IV U19130 ( .A(n19392), .Z(n19394) );
  XOR U19131 ( .A(n19398), .B(n19399), .Z(n19392) );
  AND U19132 ( .A(n146), .B(n19391), .Z(n19399) );
  XNOR U19133 ( .A(n19389), .B(n19398), .Z(n19391) );
  XNOR U19134 ( .A(n19400), .B(n19401), .Z(n19389) );
  AND U19135 ( .A(n150), .B(n19402), .Z(n19401) );
  XOR U19136 ( .A(p_input[50]), .B(n19400), .Z(n19402) );
  XNOR U19137 ( .A(n19403), .B(n19404), .Z(n19400) );
  AND U19138 ( .A(n154), .B(n19405), .Z(n19404) );
  XOR U19139 ( .A(n19406), .B(n19407), .Z(n19398) );
  AND U19140 ( .A(n158), .B(n19397), .Z(n19407) );
  XNOR U19141 ( .A(n19408), .B(n19395), .Z(n19397) );
  XOR U19142 ( .A(n19409), .B(n19410), .Z(n19395) );
  AND U19143 ( .A(n181), .B(n19411), .Z(n19410) );
  IV U19144 ( .A(n19406), .Z(n19408) );
  XOR U19145 ( .A(n19412), .B(n19413), .Z(n19406) );
  AND U19146 ( .A(n165), .B(n19405), .Z(n19413) );
  XNOR U19147 ( .A(n19403), .B(n19412), .Z(n19405) );
  XNOR U19148 ( .A(n19414), .B(n19415), .Z(n19403) );
  AND U19149 ( .A(n169), .B(n19416), .Z(n19415) );
  XOR U19150 ( .A(p_input[82]), .B(n19414), .Z(n19416) );
  XNOR U19151 ( .A(n19417), .B(n19418), .Z(n19414) );
  AND U19152 ( .A(n173), .B(n19419), .Z(n19418) );
  XOR U19153 ( .A(n19420), .B(n19421), .Z(n19412) );
  AND U19154 ( .A(n177), .B(n19411), .Z(n19421) );
  XNOR U19155 ( .A(n19422), .B(n19409), .Z(n19411) );
  XOR U19156 ( .A(n19423), .B(n19424), .Z(n19409) );
  AND U19157 ( .A(n200), .B(n19425), .Z(n19424) );
  IV U19158 ( .A(n19420), .Z(n19422) );
  XOR U19159 ( .A(n19426), .B(n19427), .Z(n19420) );
  AND U19160 ( .A(n184), .B(n19419), .Z(n19427) );
  XNOR U19161 ( .A(n19417), .B(n19426), .Z(n19419) );
  XNOR U19162 ( .A(n19428), .B(n19429), .Z(n19417) );
  AND U19163 ( .A(n188), .B(n19430), .Z(n19429) );
  XOR U19164 ( .A(p_input[114]), .B(n19428), .Z(n19430) );
  XNOR U19165 ( .A(n19431), .B(n19432), .Z(n19428) );
  AND U19166 ( .A(n192), .B(n19433), .Z(n19432) );
  XOR U19167 ( .A(n19434), .B(n19435), .Z(n19426) );
  AND U19168 ( .A(n196), .B(n19425), .Z(n19435) );
  XNOR U19169 ( .A(n19436), .B(n19423), .Z(n19425) );
  XOR U19170 ( .A(n19437), .B(n19438), .Z(n19423) );
  AND U19171 ( .A(n219), .B(n19439), .Z(n19438) );
  IV U19172 ( .A(n19434), .Z(n19436) );
  XOR U19173 ( .A(n19440), .B(n19441), .Z(n19434) );
  AND U19174 ( .A(n203), .B(n19433), .Z(n19441) );
  XNOR U19175 ( .A(n19431), .B(n19440), .Z(n19433) );
  XNOR U19176 ( .A(n19442), .B(n19443), .Z(n19431) );
  AND U19177 ( .A(n207), .B(n19444), .Z(n19443) );
  XOR U19178 ( .A(p_input[146]), .B(n19442), .Z(n19444) );
  XNOR U19179 ( .A(n19445), .B(n19446), .Z(n19442) );
  AND U19180 ( .A(n211), .B(n19447), .Z(n19446) );
  XOR U19181 ( .A(n19448), .B(n19449), .Z(n19440) );
  AND U19182 ( .A(n215), .B(n19439), .Z(n19449) );
  XNOR U19183 ( .A(n19450), .B(n19437), .Z(n19439) );
  XOR U19184 ( .A(n19451), .B(n19452), .Z(n19437) );
  AND U19185 ( .A(n238), .B(n19453), .Z(n19452) );
  IV U19186 ( .A(n19448), .Z(n19450) );
  XOR U19187 ( .A(n19454), .B(n19455), .Z(n19448) );
  AND U19188 ( .A(n222), .B(n19447), .Z(n19455) );
  XNOR U19189 ( .A(n19445), .B(n19454), .Z(n19447) );
  XNOR U19190 ( .A(n19456), .B(n19457), .Z(n19445) );
  AND U19191 ( .A(n226), .B(n19458), .Z(n19457) );
  XOR U19192 ( .A(p_input[178]), .B(n19456), .Z(n19458) );
  XNOR U19193 ( .A(n19459), .B(n19460), .Z(n19456) );
  AND U19194 ( .A(n230), .B(n19461), .Z(n19460) );
  XOR U19195 ( .A(n19462), .B(n19463), .Z(n19454) );
  AND U19196 ( .A(n234), .B(n19453), .Z(n19463) );
  XNOR U19197 ( .A(n19464), .B(n19451), .Z(n19453) );
  XOR U19198 ( .A(n19465), .B(n19466), .Z(n19451) );
  AND U19199 ( .A(n257), .B(n19467), .Z(n19466) );
  IV U19200 ( .A(n19462), .Z(n19464) );
  XOR U19201 ( .A(n19468), .B(n19469), .Z(n19462) );
  AND U19202 ( .A(n241), .B(n19461), .Z(n19469) );
  XNOR U19203 ( .A(n19459), .B(n19468), .Z(n19461) );
  XNOR U19204 ( .A(n19470), .B(n19471), .Z(n19459) );
  AND U19205 ( .A(n245), .B(n19472), .Z(n19471) );
  XOR U19206 ( .A(p_input[210]), .B(n19470), .Z(n19472) );
  XNOR U19207 ( .A(n19473), .B(n19474), .Z(n19470) );
  AND U19208 ( .A(n249), .B(n19475), .Z(n19474) );
  XOR U19209 ( .A(n19476), .B(n19477), .Z(n19468) );
  AND U19210 ( .A(n253), .B(n19467), .Z(n19477) );
  XNOR U19211 ( .A(n19478), .B(n19465), .Z(n19467) );
  XOR U19212 ( .A(n19479), .B(n19480), .Z(n19465) );
  AND U19213 ( .A(n276), .B(n19481), .Z(n19480) );
  IV U19214 ( .A(n19476), .Z(n19478) );
  XOR U19215 ( .A(n19482), .B(n19483), .Z(n19476) );
  AND U19216 ( .A(n260), .B(n19475), .Z(n19483) );
  XNOR U19217 ( .A(n19473), .B(n19482), .Z(n19475) );
  XNOR U19218 ( .A(n19484), .B(n19485), .Z(n19473) );
  AND U19219 ( .A(n264), .B(n19486), .Z(n19485) );
  XOR U19220 ( .A(p_input[242]), .B(n19484), .Z(n19486) );
  XNOR U19221 ( .A(n19487), .B(n19488), .Z(n19484) );
  AND U19222 ( .A(n268), .B(n19489), .Z(n19488) );
  XOR U19223 ( .A(n19490), .B(n19491), .Z(n19482) );
  AND U19224 ( .A(n272), .B(n19481), .Z(n19491) );
  XNOR U19225 ( .A(n19492), .B(n19479), .Z(n19481) );
  XOR U19226 ( .A(n19493), .B(n19494), .Z(n19479) );
  AND U19227 ( .A(n295), .B(n19495), .Z(n19494) );
  IV U19228 ( .A(n19490), .Z(n19492) );
  XOR U19229 ( .A(n19496), .B(n19497), .Z(n19490) );
  AND U19230 ( .A(n279), .B(n19489), .Z(n19497) );
  XNOR U19231 ( .A(n19487), .B(n19496), .Z(n19489) );
  XNOR U19232 ( .A(n19498), .B(n19499), .Z(n19487) );
  AND U19233 ( .A(n283), .B(n19500), .Z(n19499) );
  XOR U19234 ( .A(p_input[274]), .B(n19498), .Z(n19500) );
  XNOR U19235 ( .A(n19501), .B(n19502), .Z(n19498) );
  AND U19236 ( .A(n287), .B(n19503), .Z(n19502) );
  XOR U19237 ( .A(n19504), .B(n19505), .Z(n19496) );
  AND U19238 ( .A(n291), .B(n19495), .Z(n19505) );
  XNOR U19239 ( .A(n19506), .B(n19493), .Z(n19495) );
  XOR U19240 ( .A(n19507), .B(n19508), .Z(n19493) );
  AND U19241 ( .A(n314), .B(n19509), .Z(n19508) );
  IV U19242 ( .A(n19504), .Z(n19506) );
  XOR U19243 ( .A(n19510), .B(n19511), .Z(n19504) );
  AND U19244 ( .A(n298), .B(n19503), .Z(n19511) );
  XNOR U19245 ( .A(n19501), .B(n19510), .Z(n19503) );
  XNOR U19246 ( .A(n19512), .B(n19513), .Z(n19501) );
  AND U19247 ( .A(n302), .B(n19514), .Z(n19513) );
  XOR U19248 ( .A(p_input[306]), .B(n19512), .Z(n19514) );
  XNOR U19249 ( .A(n19515), .B(n19516), .Z(n19512) );
  AND U19250 ( .A(n306), .B(n19517), .Z(n19516) );
  XOR U19251 ( .A(n19518), .B(n19519), .Z(n19510) );
  AND U19252 ( .A(n310), .B(n19509), .Z(n19519) );
  XNOR U19253 ( .A(n19520), .B(n19507), .Z(n19509) );
  XOR U19254 ( .A(n19521), .B(n19522), .Z(n19507) );
  AND U19255 ( .A(n333), .B(n19523), .Z(n19522) );
  IV U19256 ( .A(n19518), .Z(n19520) );
  XOR U19257 ( .A(n19524), .B(n19525), .Z(n19518) );
  AND U19258 ( .A(n317), .B(n19517), .Z(n19525) );
  XNOR U19259 ( .A(n19515), .B(n19524), .Z(n19517) );
  XNOR U19260 ( .A(n19526), .B(n19527), .Z(n19515) );
  AND U19261 ( .A(n321), .B(n19528), .Z(n19527) );
  XOR U19262 ( .A(p_input[338]), .B(n19526), .Z(n19528) );
  XNOR U19263 ( .A(n19529), .B(n19530), .Z(n19526) );
  AND U19264 ( .A(n325), .B(n19531), .Z(n19530) );
  XOR U19265 ( .A(n19532), .B(n19533), .Z(n19524) );
  AND U19266 ( .A(n329), .B(n19523), .Z(n19533) );
  XNOR U19267 ( .A(n19534), .B(n19521), .Z(n19523) );
  XOR U19268 ( .A(n19535), .B(n19536), .Z(n19521) );
  AND U19269 ( .A(n352), .B(n19537), .Z(n19536) );
  IV U19270 ( .A(n19532), .Z(n19534) );
  XOR U19271 ( .A(n19538), .B(n19539), .Z(n19532) );
  AND U19272 ( .A(n336), .B(n19531), .Z(n19539) );
  XNOR U19273 ( .A(n19529), .B(n19538), .Z(n19531) );
  XNOR U19274 ( .A(n19540), .B(n19541), .Z(n19529) );
  AND U19275 ( .A(n340), .B(n19542), .Z(n19541) );
  XOR U19276 ( .A(p_input[370]), .B(n19540), .Z(n19542) );
  XNOR U19277 ( .A(n19543), .B(n19544), .Z(n19540) );
  AND U19278 ( .A(n344), .B(n19545), .Z(n19544) );
  XOR U19279 ( .A(n19546), .B(n19547), .Z(n19538) );
  AND U19280 ( .A(n348), .B(n19537), .Z(n19547) );
  XNOR U19281 ( .A(n19548), .B(n19535), .Z(n19537) );
  XOR U19282 ( .A(n19549), .B(n19550), .Z(n19535) );
  AND U19283 ( .A(n371), .B(n19551), .Z(n19550) );
  IV U19284 ( .A(n19546), .Z(n19548) );
  XOR U19285 ( .A(n19552), .B(n19553), .Z(n19546) );
  AND U19286 ( .A(n355), .B(n19545), .Z(n19553) );
  XNOR U19287 ( .A(n19543), .B(n19552), .Z(n19545) );
  XNOR U19288 ( .A(n19554), .B(n19555), .Z(n19543) );
  AND U19289 ( .A(n359), .B(n19556), .Z(n19555) );
  XOR U19290 ( .A(p_input[402]), .B(n19554), .Z(n19556) );
  XNOR U19291 ( .A(n19557), .B(n19558), .Z(n19554) );
  AND U19292 ( .A(n363), .B(n19559), .Z(n19558) );
  XOR U19293 ( .A(n19560), .B(n19561), .Z(n19552) );
  AND U19294 ( .A(n367), .B(n19551), .Z(n19561) );
  XNOR U19295 ( .A(n19562), .B(n19549), .Z(n19551) );
  XOR U19296 ( .A(n19563), .B(n19564), .Z(n19549) );
  AND U19297 ( .A(n390), .B(n19565), .Z(n19564) );
  IV U19298 ( .A(n19560), .Z(n19562) );
  XOR U19299 ( .A(n19566), .B(n19567), .Z(n19560) );
  AND U19300 ( .A(n374), .B(n19559), .Z(n19567) );
  XNOR U19301 ( .A(n19557), .B(n19566), .Z(n19559) );
  XNOR U19302 ( .A(n19568), .B(n19569), .Z(n19557) );
  AND U19303 ( .A(n378), .B(n19570), .Z(n19569) );
  XOR U19304 ( .A(p_input[434]), .B(n19568), .Z(n19570) );
  XNOR U19305 ( .A(n19571), .B(n19572), .Z(n19568) );
  AND U19306 ( .A(n382), .B(n19573), .Z(n19572) );
  XOR U19307 ( .A(n19574), .B(n19575), .Z(n19566) );
  AND U19308 ( .A(n386), .B(n19565), .Z(n19575) );
  XNOR U19309 ( .A(n19576), .B(n19563), .Z(n19565) );
  XOR U19310 ( .A(n19577), .B(n19578), .Z(n19563) );
  AND U19311 ( .A(n409), .B(n19579), .Z(n19578) );
  IV U19312 ( .A(n19574), .Z(n19576) );
  XOR U19313 ( .A(n19580), .B(n19581), .Z(n19574) );
  AND U19314 ( .A(n393), .B(n19573), .Z(n19581) );
  XNOR U19315 ( .A(n19571), .B(n19580), .Z(n19573) );
  XNOR U19316 ( .A(n19582), .B(n19583), .Z(n19571) );
  AND U19317 ( .A(n397), .B(n19584), .Z(n19583) );
  XOR U19318 ( .A(p_input[466]), .B(n19582), .Z(n19584) );
  XNOR U19319 ( .A(n19585), .B(n19586), .Z(n19582) );
  AND U19320 ( .A(n401), .B(n19587), .Z(n19586) );
  XOR U19321 ( .A(n19588), .B(n19589), .Z(n19580) );
  AND U19322 ( .A(n405), .B(n19579), .Z(n19589) );
  XNOR U19323 ( .A(n19590), .B(n19577), .Z(n19579) );
  XOR U19324 ( .A(n19591), .B(n19592), .Z(n19577) );
  AND U19325 ( .A(n428), .B(n19593), .Z(n19592) );
  IV U19326 ( .A(n19588), .Z(n19590) );
  XOR U19327 ( .A(n19594), .B(n19595), .Z(n19588) );
  AND U19328 ( .A(n412), .B(n19587), .Z(n19595) );
  XNOR U19329 ( .A(n19585), .B(n19594), .Z(n19587) );
  XNOR U19330 ( .A(n19596), .B(n19597), .Z(n19585) );
  AND U19331 ( .A(n416), .B(n19598), .Z(n19597) );
  XOR U19332 ( .A(p_input[498]), .B(n19596), .Z(n19598) );
  XNOR U19333 ( .A(n19599), .B(n19600), .Z(n19596) );
  AND U19334 ( .A(n420), .B(n19601), .Z(n19600) );
  XOR U19335 ( .A(n19602), .B(n19603), .Z(n19594) );
  AND U19336 ( .A(n424), .B(n19593), .Z(n19603) );
  XNOR U19337 ( .A(n19604), .B(n19591), .Z(n19593) );
  XOR U19338 ( .A(n19605), .B(n19606), .Z(n19591) );
  AND U19339 ( .A(n447), .B(n19607), .Z(n19606) );
  IV U19340 ( .A(n19602), .Z(n19604) );
  XOR U19341 ( .A(n19608), .B(n19609), .Z(n19602) );
  AND U19342 ( .A(n431), .B(n19601), .Z(n19609) );
  XNOR U19343 ( .A(n19599), .B(n19608), .Z(n19601) );
  XNOR U19344 ( .A(n19610), .B(n19611), .Z(n19599) );
  AND U19345 ( .A(n435), .B(n19612), .Z(n19611) );
  XOR U19346 ( .A(p_input[530]), .B(n19610), .Z(n19612) );
  XNOR U19347 ( .A(n19613), .B(n19614), .Z(n19610) );
  AND U19348 ( .A(n439), .B(n19615), .Z(n19614) );
  XOR U19349 ( .A(n19616), .B(n19617), .Z(n19608) );
  AND U19350 ( .A(n443), .B(n19607), .Z(n19617) );
  XNOR U19351 ( .A(n19618), .B(n19605), .Z(n19607) );
  XOR U19352 ( .A(n19619), .B(n19620), .Z(n19605) );
  AND U19353 ( .A(n466), .B(n19621), .Z(n19620) );
  IV U19354 ( .A(n19616), .Z(n19618) );
  XOR U19355 ( .A(n19622), .B(n19623), .Z(n19616) );
  AND U19356 ( .A(n450), .B(n19615), .Z(n19623) );
  XNOR U19357 ( .A(n19613), .B(n19622), .Z(n19615) );
  XNOR U19358 ( .A(n19624), .B(n19625), .Z(n19613) );
  AND U19359 ( .A(n454), .B(n19626), .Z(n19625) );
  XOR U19360 ( .A(p_input[562]), .B(n19624), .Z(n19626) );
  XNOR U19361 ( .A(n19627), .B(n19628), .Z(n19624) );
  AND U19362 ( .A(n458), .B(n19629), .Z(n19628) );
  XOR U19363 ( .A(n19630), .B(n19631), .Z(n19622) );
  AND U19364 ( .A(n462), .B(n19621), .Z(n19631) );
  XNOR U19365 ( .A(n19632), .B(n19619), .Z(n19621) );
  XOR U19366 ( .A(n19633), .B(n19634), .Z(n19619) );
  AND U19367 ( .A(n485), .B(n19635), .Z(n19634) );
  IV U19368 ( .A(n19630), .Z(n19632) );
  XOR U19369 ( .A(n19636), .B(n19637), .Z(n19630) );
  AND U19370 ( .A(n469), .B(n19629), .Z(n19637) );
  XNOR U19371 ( .A(n19627), .B(n19636), .Z(n19629) );
  XNOR U19372 ( .A(n19638), .B(n19639), .Z(n19627) );
  AND U19373 ( .A(n473), .B(n19640), .Z(n19639) );
  XOR U19374 ( .A(p_input[594]), .B(n19638), .Z(n19640) );
  XNOR U19375 ( .A(n19641), .B(n19642), .Z(n19638) );
  AND U19376 ( .A(n477), .B(n19643), .Z(n19642) );
  XOR U19377 ( .A(n19644), .B(n19645), .Z(n19636) );
  AND U19378 ( .A(n481), .B(n19635), .Z(n19645) );
  XNOR U19379 ( .A(n19646), .B(n19633), .Z(n19635) );
  XOR U19380 ( .A(n19647), .B(n19648), .Z(n19633) );
  AND U19381 ( .A(n504), .B(n19649), .Z(n19648) );
  IV U19382 ( .A(n19644), .Z(n19646) );
  XOR U19383 ( .A(n19650), .B(n19651), .Z(n19644) );
  AND U19384 ( .A(n488), .B(n19643), .Z(n19651) );
  XNOR U19385 ( .A(n19641), .B(n19650), .Z(n19643) );
  XNOR U19386 ( .A(n19652), .B(n19653), .Z(n19641) );
  AND U19387 ( .A(n492), .B(n19654), .Z(n19653) );
  XOR U19388 ( .A(p_input[626]), .B(n19652), .Z(n19654) );
  XNOR U19389 ( .A(n19655), .B(n19656), .Z(n19652) );
  AND U19390 ( .A(n496), .B(n19657), .Z(n19656) );
  XOR U19391 ( .A(n19658), .B(n19659), .Z(n19650) );
  AND U19392 ( .A(n500), .B(n19649), .Z(n19659) );
  XNOR U19393 ( .A(n19660), .B(n19647), .Z(n19649) );
  XOR U19394 ( .A(n19661), .B(n19662), .Z(n19647) );
  AND U19395 ( .A(n523), .B(n19663), .Z(n19662) );
  IV U19396 ( .A(n19658), .Z(n19660) );
  XOR U19397 ( .A(n19664), .B(n19665), .Z(n19658) );
  AND U19398 ( .A(n507), .B(n19657), .Z(n19665) );
  XNOR U19399 ( .A(n19655), .B(n19664), .Z(n19657) );
  XNOR U19400 ( .A(n19666), .B(n19667), .Z(n19655) );
  AND U19401 ( .A(n511), .B(n19668), .Z(n19667) );
  XOR U19402 ( .A(p_input[658]), .B(n19666), .Z(n19668) );
  XNOR U19403 ( .A(n19669), .B(n19670), .Z(n19666) );
  AND U19404 ( .A(n515), .B(n19671), .Z(n19670) );
  XOR U19405 ( .A(n19672), .B(n19673), .Z(n19664) );
  AND U19406 ( .A(n519), .B(n19663), .Z(n19673) );
  XNOR U19407 ( .A(n19674), .B(n19661), .Z(n19663) );
  XOR U19408 ( .A(n19675), .B(n19676), .Z(n19661) );
  AND U19409 ( .A(n542), .B(n19677), .Z(n19676) );
  IV U19410 ( .A(n19672), .Z(n19674) );
  XOR U19411 ( .A(n19678), .B(n19679), .Z(n19672) );
  AND U19412 ( .A(n526), .B(n19671), .Z(n19679) );
  XNOR U19413 ( .A(n19669), .B(n19678), .Z(n19671) );
  XNOR U19414 ( .A(n19680), .B(n19681), .Z(n19669) );
  AND U19415 ( .A(n530), .B(n19682), .Z(n19681) );
  XOR U19416 ( .A(p_input[690]), .B(n19680), .Z(n19682) );
  XNOR U19417 ( .A(n19683), .B(n19684), .Z(n19680) );
  AND U19418 ( .A(n534), .B(n19685), .Z(n19684) );
  XOR U19419 ( .A(n19686), .B(n19687), .Z(n19678) );
  AND U19420 ( .A(n538), .B(n19677), .Z(n19687) );
  XNOR U19421 ( .A(n19688), .B(n19675), .Z(n19677) );
  XOR U19422 ( .A(n19689), .B(n19690), .Z(n19675) );
  AND U19423 ( .A(n561), .B(n19691), .Z(n19690) );
  IV U19424 ( .A(n19686), .Z(n19688) );
  XOR U19425 ( .A(n19692), .B(n19693), .Z(n19686) );
  AND U19426 ( .A(n545), .B(n19685), .Z(n19693) );
  XNOR U19427 ( .A(n19683), .B(n19692), .Z(n19685) );
  XNOR U19428 ( .A(n19694), .B(n19695), .Z(n19683) );
  AND U19429 ( .A(n549), .B(n19696), .Z(n19695) );
  XOR U19430 ( .A(p_input[722]), .B(n19694), .Z(n19696) );
  XNOR U19431 ( .A(n19697), .B(n19698), .Z(n19694) );
  AND U19432 ( .A(n553), .B(n19699), .Z(n19698) );
  XOR U19433 ( .A(n19700), .B(n19701), .Z(n19692) );
  AND U19434 ( .A(n557), .B(n19691), .Z(n19701) );
  XNOR U19435 ( .A(n19702), .B(n19689), .Z(n19691) );
  XOR U19436 ( .A(n19703), .B(n19704), .Z(n19689) );
  AND U19437 ( .A(n580), .B(n19705), .Z(n19704) );
  IV U19438 ( .A(n19700), .Z(n19702) );
  XOR U19439 ( .A(n19706), .B(n19707), .Z(n19700) );
  AND U19440 ( .A(n564), .B(n19699), .Z(n19707) );
  XNOR U19441 ( .A(n19697), .B(n19706), .Z(n19699) );
  XNOR U19442 ( .A(n19708), .B(n19709), .Z(n19697) );
  AND U19443 ( .A(n568), .B(n19710), .Z(n19709) );
  XOR U19444 ( .A(p_input[754]), .B(n19708), .Z(n19710) );
  XNOR U19445 ( .A(n19711), .B(n19712), .Z(n19708) );
  AND U19446 ( .A(n572), .B(n19713), .Z(n19712) );
  XOR U19447 ( .A(n19714), .B(n19715), .Z(n19706) );
  AND U19448 ( .A(n576), .B(n19705), .Z(n19715) );
  XNOR U19449 ( .A(n19716), .B(n19703), .Z(n19705) );
  XOR U19450 ( .A(n19717), .B(n19718), .Z(n19703) );
  AND U19451 ( .A(n599), .B(n19719), .Z(n19718) );
  IV U19452 ( .A(n19714), .Z(n19716) );
  XOR U19453 ( .A(n19720), .B(n19721), .Z(n19714) );
  AND U19454 ( .A(n583), .B(n19713), .Z(n19721) );
  XNOR U19455 ( .A(n19711), .B(n19720), .Z(n19713) );
  XNOR U19456 ( .A(n19722), .B(n19723), .Z(n19711) );
  AND U19457 ( .A(n587), .B(n19724), .Z(n19723) );
  XOR U19458 ( .A(p_input[786]), .B(n19722), .Z(n19724) );
  XNOR U19459 ( .A(n19725), .B(n19726), .Z(n19722) );
  AND U19460 ( .A(n591), .B(n19727), .Z(n19726) );
  XOR U19461 ( .A(n19728), .B(n19729), .Z(n19720) );
  AND U19462 ( .A(n595), .B(n19719), .Z(n19729) );
  XNOR U19463 ( .A(n19730), .B(n19717), .Z(n19719) );
  XOR U19464 ( .A(n19731), .B(n19732), .Z(n19717) );
  AND U19465 ( .A(n618), .B(n19733), .Z(n19732) );
  IV U19466 ( .A(n19728), .Z(n19730) );
  XOR U19467 ( .A(n19734), .B(n19735), .Z(n19728) );
  AND U19468 ( .A(n602), .B(n19727), .Z(n19735) );
  XNOR U19469 ( .A(n19725), .B(n19734), .Z(n19727) );
  XNOR U19470 ( .A(n19736), .B(n19737), .Z(n19725) );
  AND U19471 ( .A(n606), .B(n19738), .Z(n19737) );
  XOR U19472 ( .A(p_input[818]), .B(n19736), .Z(n19738) );
  XNOR U19473 ( .A(n19739), .B(n19740), .Z(n19736) );
  AND U19474 ( .A(n610), .B(n19741), .Z(n19740) );
  XOR U19475 ( .A(n19742), .B(n19743), .Z(n19734) );
  AND U19476 ( .A(n614), .B(n19733), .Z(n19743) );
  XNOR U19477 ( .A(n19744), .B(n19731), .Z(n19733) );
  XOR U19478 ( .A(n19745), .B(n19746), .Z(n19731) );
  AND U19479 ( .A(n637), .B(n19747), .Z(n19746) );
  IV U19480 ( .A(n19742), .Z(n19744) );
  XOR U19481 ( .A(n19748), .B(n19749), .Z(n19742) );
  AND U19482 ( .A(n621), .B(n19741), .Z(n19749) );
  XNOR U19483 ( .A(n19739), .B(n19748), .Z(n19741) );
  XNOR U19484 ( .A(n19750), .B(n19751), .Z(n19739) );
  AND U19485 ( .A(n625), .B(n19752), .Z(n19751) );
  XOR U19486 ( .A(p_input[850]), .B(n19750), .Z(n19752) );
  XNOR U19487 ( .A(n19753), .B(n19754), .Z(n19750) );
  AND U19488 ( .A(n629), .B(n19755), .Z(n19754) );
  XOR U19489 ( .A(n19756), .B(n19757), .Z(n19748) );
  AND U19490 ( .A(n633), .B(n19747), .Z(n19757) );
  XNOR U19491 ( .A(n19758), .B(n19745), .Z(n19747) );
  XOR U19492 ( .A(n19759), .B(n19760), .Z(n19745) );
  AND U19493 ( .A(n656), .B(n19761), .Z(n19760) );
  IV U19494 ( .A(n19756), .Z(n19758) );
  XOR U19495 ( .A(n19762), .B(n19763), .Z(n19756) );
  AND U19496 ( .A(n640), .B(n19755), .Z(n19763) );
  XNOR U19497 ( .A(n19753), .B(n19762), .Z(n19755) );
  XNOR U19498 ( .A(n19764), .B(n19765), .Z(n19753) );
  AND U19499 ( .A(n644), .B(n19766), .Z(n19765) );
  XOR U19500 ( .A(p_input[882]), .B(n19764), .Z(n19766) );
  XNOR U19501 ( .A(n19767), .B(n19768), .Z(n19764) );
  AND U19502 ( .A(n648), .B(n19769), .Z(n19768) );
  XOR U19503 ( .A(n19770), .B(n19771), .Z(n19762) );
  AND U19504 ( .A(n652), .B(n19761), .Z(n19771) );
  XNOR U19505 ( .A(n19772), .B(n19759), .Z(n19761) );
  XOR U19506 ( .A(n19773), .B(n19774), .Z(n19759) );
  AND U19507 ( .A(n675), .B(n19775), .Z(n19774) );
  IV U19508 ( .A(n19770), .Z(n19772) );
  XOR U19509 ( .A(n19776), .B(n19777), .Z(n19770) );
  AND U19510 ( .A(n659), .B(n19769), .Z(n19777) );
  XNOR U19511 ( .A(n19767), .B(n19776), .Z(n19769) );
  XNOR U19512 ( .A(n19778), .B(n19779), .Z(n19767) );
  AND U19513 ( .A(n663), .B(n19780), .Z(n19779) );
  XOR U19514 ( .A(p_input[914]), .B(n19778), .Z(n19780) );
  XNOR U19515 ( .A(n19781), .B(n19782), .Z(n19778) );
  AND U19516 ( .A(n667), .B(n19783), .Z(n19782) );
  XOR U19517 ( .A(n19784), .B(n19785), .Z(n19776) );
  AND U19518 ( .A(n671), .B(n19775), .Z(n19785) );
  XNOR U19519 ( .A(n19786), .B(n19773), .Z(n19775) );
  XOR U19520 ( .A(n19787), .B(n19788), .Z(n19773) );
  AND U19521 ( .A(n694), .B(n19789), .Z(n19788) );
  IV U19522 ( .A(n19784), .Z(n19786) );
  XOR U19523 ( .A(n19790), .B(n19791), .Z(n19784) );
  AND U19524 ( .A(n678), .B(n19783), .Z(n19791) );
  XNOR U19525 ( .A(n19781), .B(n19790), .Z(n19783) );
  XNOR U19526 ( .A(n19792), .B(n19793), .Z(n19781) );
  AND U19527 ( .A(n682), .B(n19794), .Z(n19793) );
  XOR U19528 ( .A(p_input[946]), .B(n19792), .Z(n19794) );
  XNOR U19529 ( .A(n19795), .B(n19796), .Z(n19792) );
  AND U19530 ( .A(n686), .B(n19797), .Z(n19796) );
  XOR U19531 ( .A(n19798), .B(n19799), .Z(n19790) );
  AND U19532 ( .A(n690), .B(n19789), .Z(n19799) );
  XNOR U19533 ( .A(n19800), .B(n19787), .Z(n19789) );
  XOR U19534 ( .A(n19801), .B(n19802), .Z(n19787) );
  AND U19535 ( .A(n713), .B(n19803), .Z(n19802) );
  IV U19536 ( .A(n19798), .Z(n19800) );
  XOR U19537 ( .A(n19804), .B(n19805), .Z(n19798) );
  AND U19538 ( .A(n697), .B(n19797), .Z(n19805) );
  XNOR U19539 ( .A(n19795), .B(n19804), .Z(n19797) );
  XNOR U19540 ( .A(n19806), .B(n19807), .Z(n19795) );
  AND U19541 ( .A(n701), .B(n19808), .Z(n19807) );
  XOR U19542 ( .A(p_input[978]), .B(n19806), .Z(n19808) );
  XNOR U19543 ( .A(n19809), .B(n19810), .Z(n19806) );
  AND U19544 ( .A(n705), .B(n19811), .Z(n19810) );
  XOR U19545 ( .A(n19812), .B(n19813), .Z(n19804) );
  AND U19546 ( .A(n709), .B(n19803), .Z(n19813) );
  XNOR U19547 ( .A(n19814), .B(n19801), .Z(n19803) );
  XOR U19548 ( .A(n19815), .B(n19816), .Z(n19801) );
  AND U19549 ( .A(n732), .B(n19817), .Z(n19816) );
  IV U19550 ( .A(n19812), .Z(n19814) );
  XOR U19551 ( .A(n19818), .B(n19819), .Z(n19812) );
  AND U19552 ( .A(n716), .B(n19811), .Z(n19819) );
  XNOR U19553 ( .A(n19809), .B(n19818), .Z(n19811) );
  XNOR U19554 ( .A(n19820), .B(n19821), .Z(n19809) );
  AND U19555 ( .A(n720), .B(n19822), .Z(n19821) );
  XOR U19556 ( .A(p_input[1010]), .B(n19820), .Z(n19822) );
  XNOR U19557 ( .A(n19823), .B(n19824), .Z(n19820) );
  AND U19558 ( .A(n724), .B(n19825), .Z(n19824) );
  XOR U19559 ( .A(n19826), .B(n19827), .Z(n19818) );
  AND U19560 ( .A(n728), .B(n19817), .Z(n19827) );
  XNOR U19561 ( .A(n19828), .B(n19815), .Z(n19817) );
  XOR U19562 ( .A(n19829), .B(n19830), .Z(n19815) );
  AND U19563 ( .A(n751), .B(n19831), .Z(n19830) );
  IV U19564 ( .A(n19826), .Z(n19828) );
  XOR U19565 ( .A(n19832), .B(n19833), .Z(n19826) );
  AND U19566 ( .A(n735), .B(n19825), .Z(n19833) );
  XNOR U19567 ( .A(n19823), .B(n19832), .Z(n19825) );
  XNOR U19568 ( .A(n19834), .B(n19835), .Z(n19823) );
  AND U19569 ( .A(n739), .B(n19836), .Z(n19835) );
  XOR U19570 ( .A(p_input[1042]), .B(n19834), .Z(n19836) );
  XNOR U19571 ( .A(n19837), .B(n19838), .Z(n19834) );
  AND U19572 ( .A(n743), .B(n19839), .Z(n19838) );
  XOR U19573 ( .A(n19840), .B(n19841), .Z(n19832) );
  AND U19574 ( .A(n747), .B(n19831), .Z(n19841) );
  XNOR U19575 ( .A(n19842), .B(n19829), .Z(n19831) );
  XOR U19576 ( .A(n19843), .B(n19844), .Z(n19829) );
  AND U19577 ( .A(n770), .B(n19845), .Z(n19844) );
  IV U19578 ( .A(n19840), .Z(n19842) );
  XOR U19579 ( .A(n19846), .B(n19847), .Z(n19840) );
  AND U19580 ( .A(n754), .B(n19839), .Z(n19847) );
  XNOR U19581 ( .A(n19837), .B(n19846), .Z(n19839) );
  XNOR U19582 ( .A(n19848), .B(n19849), .Z(n19837) );
  AND U19583 ( .A(n758), .B(n19850), .Z(n19849) );
  XOR U19584 ( .A(p_input[1074]), .B(n19848), .Z(n19850) );
  XNOR U19585 ( .A(n19851), .B(n19852), .Z(n19848) );
  AND U19586 ( .A(n762), .B(n19853), .Z(n19852) );
  XOR U19587 ( .A(n19854), .B(n19855), .Z(n19846) );
  AND U19588 ( .A(n766), .B(n19845), .Z(n19855) );
  XNOR U19589 ( .A(n19856), .B(n19843), .Z(n19845) );
  XOR U19590 ( .A(n19857), .B(n19858), .Z(n19843) );
  AND U19591 ( .A(n789), .B(n19859), .Z(n19858) );
  IV U19592 ( .A(n19854), .Z(n19856) );
  XOR U19593 ( .A(n19860), .B(n19861), .Z(n19854) );
  AND U19594 ( .A(n773), .B(n19853), .Z(n19861) );
  XNOR U19595 ( .A(n19851), .B(n19860), .Z(n19853) );
  XNOR U19596 ( .A(n19862), .B(n19863), .Z(n19851) );
  AND U19597 ( .A(n777), .B(n19864), .Z(n19863) );
  XOR U19598 ( .A(p_input[1106]), .B(n19862), .Z(n19864) );
  XNOR U19599 ( .A(n19865), .B(n19866), .Z(n19862) );
  AND U19600 ( .A(n781), .B(n19867), .Z(n19866) );
  XOR U19601 ( .A(n19868), .B(n19869), .Z(n19860) );
  AND U19602 ( .A(n785), .B(n19859), .Z(n19869) );
  XNOR U19603 ( .A(n19870), .B(n19857), .Z(n19859) );
  XOR U19604 ( .A(n19871), .B(n19872), .Z(n19857) );
  AND U19605 ( .A(n808), .B(n19873), .Z(n19872) );
  IV U19606 ( .A(n19868), .Z(n19870) );
  XOR U19607 ( .A(n19874), .B(n19875), .Z(n19868) );
  AND U19608 ( .A(n792), .B(n19867), .Z(n19875) );
  XNOR U19609 ( .A(n19865), .B(n19874), .Z(n19867) );
  XNOR U19610 ( .A(n19876), .B(n19877), .Z(n19865) );
  AND U19611 ( .A(n796), .B(n19878), .Z(n19877) );
  XOR U19612 ( .A(p_input[1138]), .B(n19876), .Z(n19878) );
  XNOR U19613 ( .A(n19879), .B(n19880), .Z(n19876) );
  AND U19614 ( .A(n800), .B(n19881), .Z(n19880) );
  XOR U19615 ( .A(n19882), .B(n19883), .Z(n19874) );
  AND U19616 ( .A(n804), .B(n19873), .Z(n19883) );
  XNOR U19617 ( .A(n19884), .B(n19871), .Z(n19873) );
  XOR U19618 ( .A(n19885), .B(n19886), .Z(n19871) );
  AND U19619 ( .A(n827), .B(n19887), .Z(n19886) );
  IV U19620 ( .A(n19882), .Z(n19884) );
  XOR U19621 ( .A(n19888), .B(n19889), .Z(n19882) );
  AND U19622 ( .A(n811), .B(n19881), .Z(n19889) );
  XNOR U19623 ( .A(n19879), .B(n19888), .Z(n19881) );
  XNOR U19624 ( .A(n19890), .B(n19891), .Z(n19879) );
  AND U19625 ( .A(n815), .B(n19892), .Z(n19891) );
  XOR U19626 ( .A(p_input[1170]), .B(n19890), .Z(n19892) );
  XNOR U19627 ( .A(n19893), .B(n19894), .Z(n19890) );
  AND U19628 ( .A(n819), .B(n19895), .Z(n19894) );
  XOR U19629 ( .A(n19896), .B(n19897), .Z(n19888) );
  AND U19630 ( .A(n823), .B(n19887), .Z(n19897) );
  XNOR U19631 ( .A(n19898), .B(n19885), .Z(n19887) );
  XOR U19632 ( .A(n19899), .B(n19900), .Z(n19885) );
  AND U19633 ( .A(n846), .B(n19901), .Z(n19900) );
  IV U19634 ( .A(n19896), .Z(n19898) );
  XOR U19635 ( .A(n19902), .B(n19903), .Z(n19896) );
  AND U19636 ( .A(n830), .B(n19895), .Z(n19903) );
  XNOR U19637 ( .A(n19893), .B(n19902), .Z(n19895) );
  XNOR U19638 ( .A(n19904), .B(n19905), .Z(n19893) );
  AND U19639 ( .A(n834), .B(n19906), .Z(n19905) );
  XOR U19640 ( .A(p_input[1202]), .B(n19904), .Z(n19906) );
  XNOR U19641 ( .A(n19907), .B(n19908), .Z(n19904) );
  AND U19642 ( .A(n838), .B(n19909), .Z(n19908) );
  XOR U19643 ( .A(n19910), .B(n19911), .Z(n19902) );
  AND U19644 ( .A(n842), .B(n19901), .Z(n19911) );
  XNOR U19645 ( .A(n19912), .B(n19899), .Z(n19901) );
  XOR U19646 ( .A(n19913), .B(n19914), .Z(n19899) );
  AND U19647 ( .A(n865), .B(n19915), .Z(n19914) );
  IV U19648 ( .A(n19910), .Z(n19912) );
  XOR U19649 ( .A(n19916), .B(n19917), .Z(n19910) );
  AND U19650 ( .A(n849), .B(n19909), .Z(n19917) );
  XNOR U19651 ( .A(n19907), .B(n19916), .Z(n19909) );
  XNOR U19652 ( .A(n19918), .B(n19919), .Z(n19907) );
  AND U19653 ( .A(n853), .B(n19920), .Z(n19919) );
  XOR U19654 ( .A(p_input[1234]), .B(n19918), .Z(n19920) );
  XNOR U19655 ( .A(n19921), .B(n19922), .Z(n19918) );
  AND U19656 ( .A(n857), .B(n19923), .Z(n19922) );
  XOR U19657 ( .A(n19924), .B(n19925), .Z(n19916) );
  AND U19658 ( .A(n861), .B(n19915), .Z(n19925) );
  XNOR U19659 ( .A(n19926), .B(n19913), .Z(n19915) );
  XOR U19660 ( .A(n19927), .B(n19928), .Z(n19913) );
  AND U19661 ( .A(n884), .B(n19929), .Z(n19928) );
  IV U19662 ( .A(n19924), .Z(n19926) );
  XOR U19663 ( .A(n19930), .B(n19931), .Z(n19924) );
  AND U19664 ( .A(n868), .B(n19923), .Z(n19931) );
  XNOR U19665 ( .A(n19921), .B(n19930), .Z(n19923) );
  XNOR U19666 ( .A(n19932), .B(n19933), .Z(n19921) );
  AND U19667 ( .A(n872), .B(n19934), .Z(n19933) );
  XOR U19668 ( .A(p_input[1266]), .B(n19932), .Z(n19934) );
  XNOR U19669 ( .A(n19935), .B(n19936), .Z(n19932) );
  AND U19670 ( .A(n876), .B(n19937), .Z(n19936) );
  XOR U19671 ( .A(n19938), .B(n19939), .Z(n19930) );
  AND U19672 ( .A(n880), .B(n19929), .Z(n19939) );
  XNOR U19673 ( .A(n19940), .B(n19927), .Z(n19929) );
  XOR U19674 ( .A(n19941), .B(n19942), .Z(n19927) );
  AND U19675 ( .A(n903), .B(n19943), .Z(n19942) );
  IV U19676 ( .A(n19938), .Z(n19940) );
  XOR U19677 ( .A(n19944), .B(n19945), .Z(n19938) );
  AND U19678 ( .A(n887), .B(n19937), .Z(n19945) );
  XNOR U19679 ( .A(n19935), .B(n19944), .Z(n19937) );
  XNOR U19680 ( .A(n19946), .B(n19947), .Z(n19935) );
  AND U19681 ( .A(n891), .B(n19948), .Z(n19947) );
  XOR U19682 ( .A(p_input[1298]), .B(n19946), .Z(n19948) );
  XNOR U19683 ( .A(n19949), .B(n19950), .Z(n19946) );
  AND U19684 ( .A(n895), .B(n19951), .Z(n19950) );
  XOR U19685 ( .A(n19952), .B(n19953), .Z(n19944) );
  AND U19686 ( .A(n899), .B(n19943), .Z(n19953) );
  XNOR U19687 ( .A(n19954), .B(n19941), .Z(n19943) );
  XOR U19688 ( .A(n19955), .B(n19956), .Z(n19941) );
  AND U19689 ( .A(n922), .B(n19957), .Z(n19956) );
  IV U19690 ( .A(n19952), .Z(n19954) );
  XOR U19691 ( .A(n19958), .B(n19959), .Z(n19952) );
  AND U19692 ( .A(n906), .B(n19951), .Z(n19959) );
  XNOR U19693 ( .A(n19949), .B(n19958), .Z(n19951) );
  XNOR U19694 ( .A(n19960), .B(n19961), .Z(n19949) );
  AND U19695 ( .A(n910), .B(n19962), .Z(n19961) );
  XOR U19696 ( .A(p_input[1330]), .B(n19960), .Z(n19962) );
  XNOR U19697 ( .A(n19963), .B(n19964), .Z(n19960) );
  AND U19698 ( .A(n914), .B(n19965), .Z(n19964) );
  XOR U19699 ( .A(n19966), .B(n19967), .Z(n19958) );
  AND U19700 ( .A(n918), .B(n19957), .Z(n19967) );
  XNOR U19701 ( .A(n19968), .B(n19955), .Z(n19957) );
  XOR U19702 ( .A(n19969), .B(n19970), .Z(n19955) );
  AND U19703 ( .A(n941), .B(n19971), .Z(n19970) );
  IV U19704 ( .A(n19966), .Z(n19968) );
  XOR U19705 ( .A(n19972), .B(n19973), .Z(n19966) );
  AND U19706 ( .A(n925), .B(n19965), .Z(n19973) );
  XNOR U19707 ( .A(n19963), .B(n19972), .Z(n19965) );
  XNOR U19708 ( .A(n19974), .B(n19975), .Z(n19963) );
  AND U19709 ( .A(n929), .B(n19976), .Z(n19975) );
  XOR U19710 ( .A(p_input[1362]), .B(n19974), .Z(n19976) );
  XNOR U19711 ( .A(n19977), .B(n19978), .Z(n19974) );
  AND U19712 ( .A(n933), .B(n19979), .Z(n19978) );
  XOR U19713 ( .A(n19980), .B(n19981), .Z(n19972) );
  AND U19714 ( .A(n937), .B(n19971), .Z(n19981) );
  XNOR U19715 ( .A(n19982), .B(n19969), .Z(n19971) );
  XOR U19716 ( .A(n19983), .B(n19984), .Z(n19969) );
  AND U19717 ( .A(n960), .B(n19985), .Z(n19984) );
  IV U19718 ( .A(n19980), .Z(n19982) );
  XOR U19719 ( .A(n19986), .B(n19987), .Z(n19980) );
  AND U19720 ( .A(n944), .B(n19979), .Z(n19987) );
  XNOR U19721 ( .A(n19977), .B(n19986), .Z(n19979) );
  XNOR U19722 ( .A(n19988), .B(n19989), .Z(n19977) );
  AND U19723 ( .A(n948), .B(n19990), .Z(n19989) );
  XOR U19724 ( .A(p_input[1394]), .B(n19988), .Z(n19990) );
  XNOR U19725 ( .A(n19991), .B(n19992), .Z(n19988) );
  AND U19726 ( .A(n952), .B(n19993), .Z(n19992) );
  XOR U19727 ( .A(n19994), .B(n19995), .Z(n19986) );
  AND U19728 ( .A(n956), .B(n19985), .Z(n19995) );
  XNOR U19729 ( .A(n19996), .B(n19983), .Z(n19985) );
  XOR U19730 ( .A(n19997), .B(n19998), .Z(n19983) );
  AND U19731 ( .A(n979), .B(n19999), .Z(n19998) );
  IV U19732 ( .A(n19994), .Z(n19996) );
  XOR U19733 ( .A(n20000), .B(n20001), .Z(n19994) );
  AND U19734 ( .A(n963), .B(n19993), .Z(n20001) );
  XNOR U19735 ( .A(n19991), .B(n20000), .Z(n19993) );
  XNOR U19736 ( .A(n20002), .B(n20003), .Z(n19991) );
  AND U19737 ( .A(n967), .B(n20004), .Z(n20003) );
  XOR U19738 ( .A(p_input[1426]), .B(n20002), .Z(n20004) );
  XNOR U19739 ( .A(n20005), .B(n20006), .Z(n20002) );
  AND U19740 ( .A(n971), .B(n20007), .Z(n20006) );
  XOR U19741 ( .A(n20008), .B(n20009), .Z(n20000) );
  AND U19742 ( .A(n975), .B(n19999), .Z(n20009) );
  XNOR U19743 ( .A(n20010), .B(n19997), .Z(n19999) );
  XOR U19744 ( .A(n20011), .B(n20012), .Z(n19997) );
  AND U19745 ( .A(n998), .B(n20013), .Z(n20012) );
  IV U19746 ( .A(n20008), .Z(n20010) );
  XOR U19747 ( .A(n20014), .B(n20015), .Z(n20008) );
  AND U19748 ( .A(n982), .B(n20007), .Z(n20015) );
  XNOR U19749 ( .A(n20005), .B(n20014), .Z(n20007) );
  XNOR U19750 ( .A(n20016), .B(n20017), .Z(n20005) );
  AND U19751 ( .A(n986), .B(n20018), .Z(n20017) );
  XOR U19752 ( .A(p_input[1458]), .B(n20016), .Z(n20018) );
  XNOR U19753 ( .A(n20019), .B(n20020), .Z(n20016) );
  AND U19754 ( .A(n990), .B(n20021), .Z(n20020) );
  XOR U19755 ( .A(n20022), .B(n20023), .Z(n20014) );
  AND U19756 ( .A(n994), .B(n20013), .Z(n20023) );
  XNOR U19757 ( .A(n20024), .B(n20011), .Z(n20013) );
  XOR U19758 ( .A(n20025), .B(n20026), .Z(n20011) );
  AND U19759 ( .A(n1017), .B(n20027), .Z(n20026) );
  IV U19760 ( .A(n20022), .Z(n20024) );
  XOR U19761 ( .A(n20028), .B(n20029), .Z(n20022) );
  AND U19762 ( .A(n1001), .B(n20021), .Z(n20029) );
  XNOR U19763 ( .A(n20019), .B(n20028), .Z(n20021) );
  XNOR U19764 ( .A(n20030), .B(n20031), .Z(n20019) );
  AND U19765 ( .A(n1005), .B(n20032), .Z(n20031) );
  XOR U19766 ( .A(p_input[1490]), .B(n20030), .Z(n20032) );
  XNOR U19767 ( .A(n20033), .B(n20034), .Z(n20030) );
  AND U19768 ( .A(n1009), .B(n20035), .Z(n20034) );
  XOR U19769 ( .A(n20036), .B(n20037), .Z(n20028) );
  AND U19770 ( .A(n1013), .B(n20027), .Z(n20037) );
  XNOR U19771 ( .A(n20038), .B(n20025), .Z(n20027) );
  XOR U19772 ( .A(n20039), .B(n20040), .Z(n20025) );
  AND U19773 ( .A(n1036), .B(n20041), .Z(n20040) );
  IV U19774 ( .A(n20036), .Z(n20038) );
  XOR U19775 ( .A(n20042), .B(n20043), .Z(n20036) );
  AND U19776 ( .A(n1020), .B(n20035), .Z(n20043) );
  XNOR U19777 ( .A(n20033), .B(n20042), .Z(n20035) );
  XNOR U19778 ( .A(n20044), .B(n20045), .Z(n20033) );
  AND U19779 ( .A(n1024), .B(n20046), .Z(n20045) );
  XOR U19780 ( .A(p_input[1522]), .B(n20044), .Z(n20046) );
  XNOR U19781 ( .A(n20047), .B(n20048), .Z(n20044) );
  AND U19782 ( .A(n1028), .B(n20049), .Z(n20048) );
  XOR U19783 ( .A(n20050), .B(n20051), .Z(n20042) );
  AND U19784 ( .A(n1032), .B(n20041), .Z(n20051) );
  XNOR U19785 ( .A(n20052), .B(n20039), .Z(n20041) );
  XOR U19786 ( .A(n20053), .B(n20054), .Z(n20039) );
  AND U19787 ( .A(n1055), .B(n20055), .Z(n20054) );
  IV U19788 ( .A(n20050), .Z(n20052) );
  XOR U19789 ( .A(n20056), .B(n20057), .Z(n20050) );
  AND U19790 ( .A(n1039), .B(n20049), .Z(n20057) );
  XNOR U19791 ( .A(n20047), .B(n20056), .Z(n20049) );
  XNOR U19792 ( .A(n20058), .B(n20059), .Z(n20047) );
  AND U19793 ( .A(n1043), .B(n20060), .Z(n20059) );
  XOR U19794 ( .A(p_input[1554]), .B(n20058), .Z(n20060) );
  XNOR U19795 ( .A(n20061), .B(n20062), .Z(n20058) );
  AND U19796 ( .A(n1047), .B(n20063), .Z(n20062) );
  XOR U19797 ( .A(n20064), .B(n20065), .Z(n20056) );
  AND U19798 ( .A(n1051), .B(n20055), .Z(n20065) );
  XNOR U19799 ( .A(n20066), .B(n20053), .Z(n20055) );
  XOR U19800 ( .A(n20067), .B(n20068), .Z(n20053) );
  AND U19801 ( .A(n1074), .B(n20069), .Z(n20068) );
  IV U19802 ( .A(n20064), .Z(n20066) );
  XOR U19803 ( .A(n20070), .B(n20071), .Z(n20064) );
  AND U19804 ( .A(n1058), .B(n20063), .Z(n20071) );
  XNOR U19805 ( .A(n20061), .B(n20070), .Z(n20063) );
  XNOR U19806 ( .A(n20072), .B(n20073), .Z(n20061) );
  AND U19807 ( .A(n1062), .B(n20074), .Z(n20073) );
  XOR U19808 ( .A(p_input[1586]), .B(n20072), .Z(n20074) );
  XNOR U19809 ( .A(n20075), .B(n20076), .Z(n20072) );
  AND U19810 ( .A(n1066), .B(n20077), .Z(n20076) );
  XOR U19811 ( .A(n20078), .B(n20079), .Z(n20070) );
  AND U19812 ( .A(n1070), .B(n20069), .Z(n20079) );
  XNOR U19813 ( .A(n20080), .B(n20067), .Z(n20069) );
  XOR U19814 ( .A(n20081), .B(n20082), .Z(n20067) );
  AND U19815 ( .A(n1093), .B(n20083), .Z(n20082) );
  IV U19816 ( .A(n20078), .Z(n20080) );
  XOR U19817 ( .A(n20084), .B(n20085), .Z(n20078) );
  AND U19818 ( .A(n1077), .B(n20077), .Z(n20085) );
  XNOR U19819 ( .A(n20075), .B(n20084), .Z(n20077) );
  XNOR U19820 ( .A(n20086), .B(n20087), .Z(n20075) );
  AND U19821 ( .A(n1081), .B(n20088), .Z(n20087) );
  XOR U19822 ( .A(p_input[1618]), .B(n20086), .Z(n20088) );
  XNOR U19823 ( .A(n20089), .B(n20090), .Z(n20086) );
  AND U19824 ( .A(n1085), .B(n20091), .Z(n20090) );
  XOR U19825 ( .A(n20092), .B(n20093), .Z(n20084) );
  AND U19826 ( .A(n1089), .B(n20083), .Z(n20093) );
  XNOR U19827 ( .A(n20094), .B(n20081), .Z(n20083) );
  XOR U19828 ( .A(n20095), .B(n20096), .Z(n20081) );
  AND U19829 ( .A(n1112), .B(n20097), .Z(n20096) );
  IV U19830 ( .A(n20092), .Z(n20094) );
  XOR U19831 ( .A(n20098), .B(n20099), .Z(n20092) );
  AND U19832 ( .A(n1096), .B(n20091), .Z(n20099) );
  XNOR U19833 ( .A(n20089), .B(n20098), .Z(n20091) );
  XNOR U19834 ( .A(n20100), .B(n20101), .Z(n20089) );
  AND U19835 ( .A(n1100), .B(n20102), .Z(n20101) );
  XOR U19836 ( .A(p_input[1650]), .B(n20100), .Z(n20102) );
  XNOR U19837 ( .A(n20103), .B(n20104), .Z(n20100) );
  AND U19838 ( .A(n1104), .B(n20105), .Z(n20104) );
  XOR U19839 ( .A(n20106), .B(n20107), .Z(n20098) );
  AND U19840 ( .A(n1108), .B(n20097), .Z(n20107) );
  XNOR U19841 ( .A(n20108), .B(n20095), .Z(n20097) );
  XOR U19842 ( .A(n20109), .B(n20110), .Z(n20095) );
  AND U19843 ( .A(n1131), .B(n20111), .Z(n20110) );
  IV U19844 ( .A(n20106), .Z(n20108) );
  XOR U19845 ( .A(n20112), .B(n20113), .Z(n20106) );
  AND U19846 ( .A(n1115), .B(n20105), .Z(n20113) );
  XNOR U19847 ( .A(n20103), .B(n20112), .Z(n20105) );
  XNOR U19848 ( .A(n20114), .B(n20115), .Z(n20103) );
  AND U19849 ( .A(n1119), .B(n20116), .Z(n20115) );
  XOR U19850 ( .A(p_input[1682]), .B(n20114), .Z(n20116) );
  XNOR U19851 ( .A(n20117), .B(n20118), .Z(n20114) );
  AND U19852 ( .A(n1123), .B(n20119), .Z(n20118) );
  XOR U19853 ( .A(n20120), .B(n20121), .Z(n20112) );
  AND U19854 ( .A(n1127), .B(n20111), .Z(n20121) );
  XNOR U19855 ( .A(n20122), .B(n20109), .Z(n20111) );
  XOR U19856 ( .A(n20123), .B(n20124), .Z(n20109) );
  AND U19857 ( .A(n1150), .B(n20125), .Z(n20124) );
  IV U19858 ( .A(n20120), .Z(n20122) );
  XOR U19859 ( .A(n20126), .B(n20127), .Z(n20120) );
  AND U19860 ( .A(n1134), .B(n20119), .Z(n20127) );
  XNOR U19861 ( .A(n20117), .B(n20126), .Z(n20119) );
  XNOR U19862 ( .A(n20128), .B(n20129), .Z(n20117) );
  AND U19863 ( .A(n1138), .B(n20130), .Z(n20129) );
  XOR U19864 ( .A(p_input[1714]), .B(n20128), .Z(n20130) );
  XNOR U19865 ( .A(n20131), .B(n20132), .Z(n20128) );
  AND U19866 ( .A(n1142), .B(n20133), .Z(n20132) );
  XOR U19867 ( .A(n20134), .B(n20135), .Z(n20126) );
  AND U19868 ( .A(n1146), .B(n20125), .Z(n20135) );
  XNOR U19869 ( .A(n20136), .B(n20123), .Z(n20125) );
  XOR U19870 ( .A(n20137), .B(n20138), .Z(n20123) );
  AND U19871 ( .A(n1169), .B(n20139), .Z(n20138) );
  IV U19872 ( .A(n20134), .Z(n20136) );
  XOR U19873 ( .A(n20140), .B(n20141), .Z(n20134) );
  AND U19874 ( .A(n1153), .B(n20133), .Z(n20141) );
  XNOR U19875 ( .A(n20131), .B(n20140), .Z(n20133) );
  XNOR U19876 ( .A(n20142), .B(n20143), .Z(n20131) );
  AND U19877 ( .A(n1157), .B(n20144), .Z(n20143) );
  XOR U19878 ( .A(p_input[1746]), .B(n20142), .Z(n20144) );
  XNOR U19879 ( .A(n20145), .B(n20146), .Z(n20142) );
  AND U19880 ( .A(n1161), .B(n20147), .Z(n20146) );
  XOR U19881 ( .A(n20148), .B(n20149), .Z(n20140) );
  AND U19882 ( .A(n1165), .B(n20139), .Z(n20149) );
  XNOR U19883 ( .A(n20150), .B(n20137), .Z(n20139) );
  XOR U19884 ( .A(n20151), .B(n20152), .Z(n20137) );
  AND U19885 ( .A(n1188), .B(n20153), .Z(n20152) );
  IV U19886 ( .A(n20148), .Z(n20150) );
  XOR U19887 ( .A(n20154), .B(n20155), .Z(n20148) );
  AND U19888 ( .A(n1172), .B(n20147), .Z(n20155) );
  XNOR U19889 ( .A(n20145), .B(n20154), .Z(n20147) );
  XNOR U19890 ( .A(n20156), .B(n20157), .Z(n20145) );
  AND U19891 ( .A(n1176), .B(n20158), .Z(n20157) );
  XOR U19892 ( .A(p_input[1778]), .B(n20156), .Z(n20158) );
  XNOR U19893 ( .A(n20159), .B(n20160), .Z(n20156) );
  AND U19894 ( .A(n1180), .B(n20161), .Z(n20160) );
  XOR U19895 ( .A(n20162), .B(n20163), .Z(n20154) );
  AND U19896 ( .A(n1184), .B(n20153), .Z(n20163) );
  XNOR U19897 ( .A(n20164), .B(n20151), .Z(n20153) );
  XOR U19898 ( .A(n20165), .B(n20166), .Z(n20151) );
  AND U19899 ( .A(n1207), .B(n20167), .Z(n20166) );
  IV U19900 ( .A(n20162), .Z(n20164) );
  XOR U19901 ( .A(n20168), .B(n20169), .Z(n20162) );
  AND U19902 ( .A(n1191), .B(n20161), .Z(n20169) );
  XNOR U19903 ( .A(n20159), .B(n20168), .Z(n20161) );
  XNOR U19904 ( .A(n20170), .B(n20171), .Z(n20159) );
  AND U19905 ( .A(n1195), .B(n20172), .Z(n20171) );
  XOR U19906 ( .A(p_input[1810]), .B(n20170), .Z(n20172) );
  XNOR U19907 ( .A(n20173), .B(n20174), .Z(n20170) );
  AND U19908 ( .A(n1199), .B(n20175), .Z(n20174) );
  XOR U19909 ( .A(n20176), .B(n20177), .Z(n20168) );
  AND U19910 ( .A(n1203), .B(n20167), .Z(n20177) );
  XNOR U19911 ( .A(n20178), .B(n20165), .Z(n20167) );
  XOR U19912 ( .A(n20179), .B(n20180), .Z(n20165) );
  AND U19913 ( .A(n1226), .B(n20181), .Z(n20180) );
  IV U19914 ( .A(n20176), .Z(n20178) );
  XOR U19915 ( .A(n20182), .B(n20183), .Z(n20176) );
  AND U19916 ( .A(n1210), .B(n20175), .Z(n20183) );
  XNOR U19917 ( .A(n20173), .B(n20182), .Z(n20175) );
  XNOR U19918 ( .A(n20184), .B(n20185), .Z(n20173) );
  AND U19919 ( .A(n1214), .B(n20186), .Z(n20185) );
  XOR U19920 ( .A(p_input[1842]), .B(n20184), .Z(n20186) );
  XNOR U19921 ( .A(n20187), .B(n20188), .Z(n20184) );
  AND U19922 ( .A(n1218), .B(n20189), .Z(n20188) );
  XOR U19923 ( .A(n20190), .B(n20191), .Z(n20182) );
  AND U19924 ( .A(n1222), .B(n20181), .Z(n20191) );
  XNOR U19925 ( .A(n20192), .B(n20179), .Z(n20181) );
  XOR U19926 ( .A(n20193), .B(n20194), .Z(n20179) );
  AND U19927 ( .A(n1245), .B(n20195), .Z(n20194) );
  IV U19928 ( .A(n20190), .Z(n20192) );
  XOR U19929 ( .A(n20196), .B(n20197), .Z(n20190) );
  AND U19930 ( .A(n1229), .B(n20189), .Z(n20197) );
  XNOR U19931 ( .A(n20187), .B(n20196), .Z(n20189) );
  XNOR U19932 ( .A(n20198), .B(n20199), .Z(n20187) );
  AND U19933 ( .A(n1233), .B(n20200), .Z(n20199) );
  XOR U19934 ( .A(p_input[1874]), .B(n20198), .Z(n20200) );
  XNOR U19935 ( .A(n20201), .B(n20202), .Z(n20198) );
  AND U19936 ( .A(n1237), .B(n20203), .Z(n20202) );
  XOR U19937 ( .A(n20204), .B(n20205), .Z(n20196) );
  AND U19938 ( .A(n1241), .B(n20195), .Z(n20205) );
  XNOR U19939 ( .A(n20206), .B(n20193), .Z(n20195) );
  XOR U19940 ( .A(n20207), .B(n20208), .Z(n20193) );
  AND U19941 ( .A(n1264), .B(n20209), .Z(n20208) );
  IV U19942 ( .A(n20204), .Z(n20206) );
  XOR U19943 ( .A(n20210), .B(n20211), .Z(n20204) );
  AND U19944 ( .A(n1248), .B(n20203), .Z(n20211) );
  XNOR U19945 ( .A(n20201), .B(n20210), .Z(n20203) );
  XNOR U19946 ( .A(n20212), .B(n20213), .Z(n20201) );
  AND U19947 ( .A(n1252), .B(n20214), .Z(n20213) );
  XOR U19948 ( .A(p_input[1906]), .B(n20212), .Z(n20214) );
  XNOR U19949 ( .A(n20215), .B(n20216), .Z(n20212) );
  AND U19950 ( .A(n1256), .B(n20217), .Z(n20216) );
  XOR U19951 ( .A(n20218), .B(n20219), .Z(n20210) );
  AND U19952 ( .A(n1260), .B(n20209), .Z(n20219) );
  XNOR U19953 ( .A(n20220), .B(n20207), .Z(n20209) );
  XOR U19954 ( .A(n20221), .B(n20222), .Z(n20207) );
  AND U19955 ( .A(n1282), .B(n20223), .Z(n20222) );
  IV U19956 ( .A(n20218), .Z(n20220) );
  XOR U19957 ( .A(n20224), .B(n20225), .Z(n20218) );
  AND U19958 ( .A(n1267), .B(n20217), .Z(n20225) );
  XNOR U19959 ( .A(n20215), .B(n20224), .Z(n20217) );
  XNOR U19960 ( .A(n20226), .B(n20227), .Z(n20215) );
  AND U19961 ( .A(n1271), .B(n20228), .Z(n20227) );
  XOR U19962 ( .A(p_input[1938]), .B(n20226), .Z(n20228) );
  XOR U19963 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][18] ), .B(n20229), 
        .Z(n20226) );
  AND U19964 ( .A(n1274), .B(n20230), .Z(n20229) );
  XOR U19965 ( .A(n20231), .B(n20232), .Z(n20224) );
  AND U19966 ( .A(n1278), .B(n20223), .Z(n20232) );
  XNOR U19967 ( .A(n20233), .B(n20221), .Z(n20223) );
  XOR U19968 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n20234), .Z(n20221) );
  AND U19969 ( .A(n1290), .B(n20235), .Z(n20234) );
  IV U19970 ( .A(n20231), .Z(n20233) );
  XOR U19971 ( .A(n20236), .B(n20237), .Z(n20231) );
  AND U19972 ( .A(n1285), .B(n20230), .Z(n20237) );
  XOR U19973 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][18] ), .B(n20236), 
        .Z(n20230) );
  XOR U19974 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .B(n20238), 
        .Z(n20236) );
  AND U19975 ( .A(n1287), .B(n20235), .Z(n20238) );
  XOR U19976 ( .A(\knn_comb_/min_val_out[0][18] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .Z(n20235) );
  XOR U19977 ( .A(n105), .B(n20239), .Z(o[17]) );
  AND U19978 ( .A(n122), .B(n20240), .Z(n105) );
  XOR U19979 ( .A(n106), .B(n20239), .Z(n20240) );
  XOR U19980 ( .A(n20241), .B(n20242), .Z(n20239) );
  AND U19981 ( .A(n142), .B(n20243), .Z(n20242) );
  XOR U19982 ( .A(n20244), .B(n33), .Z(n106) );
  AND U19983 ( .A(n125), .B(n20245), .Z(n33) );
  XOR U19984 ( .A(n34), .B(n20244), .Z(n20245) );
  XOR U19985 ( .A(n20246), .B(n20247), .Z(n34) );
  AND U19986 ( .A(n130), .B(n20248), .Z(n20247) );
  XOR U19987 ( .A(p_input[17]), .B(n20246), .Z(n20248) );
  XNOR U19988 ( .A(n20249), .B(n20250), .Z(n20246) );
  AND U19989 ( .A(n134), .B(n20251), .Z(n20250) );
  XOR U19990 ( .A(n20252), .B(n20253), .Z(n20244) );
  AND U19991 ( .A(n138), .B(n20243), .Z(n20253) );
  XNOR U19992 ( .A(n20254), .B(n20241), .Z(n20243) );
  XOR U19993 ( .A(n20255), .B(n20256), .Z(n20241) );
  AND U19994 ( .A(n162), .B(n20257), .Z(n20256) );
  IV U19995 ( .A(n20252), .Z(n20254) );
  XOR U19996 ( .A(n20258), .B(n20259), .Z(n20252) );
  AND U19997 ( .A(n146), .B(n20251), .Z(n20259) );
  XNOR U19998 ( .A(n20249), .B(n20258), .Z(n20251) );
  XNOR U19999 ( .A(n20260), .B(n20261), .Z(n20249) );
  AND U20000 ( .A(n150), .B(n20262), .Z(n20261) );
  XOR U20001 ( .A(p_input[49]), .B(n20260), .Z(n20262) );
  XNOR U20002 ( .A(n20263), .B(n20264), .Z(n20260) );
  AND U20003 ( .A(n154), .B(n20265), .Z(n20264) );
  XOR U20004 ( .A(n20266), .B(n20267), .Z(n20258) );
  AND U20005 ( .A(n158), .B(n20257), .Z(n20267) );
  XNOR U20006 ( .A(n20268), .B(n20255), .Z(n20257) );
  XOR U20007 ( .A(n20269), .B(n20270), .Z(n20255) );
  AND U20008 ( .A(n181), .B(n20271), .Z(n20270) );
  IV U20009 ( .A(n20266), .Z(n20268) );
  XOR U20010 ( .A(n20272), .B(n20273), .Z(n20266) );
  AND U20011 ( .A(n165), .B(n20265), .Z(n20273) );
  XNOR U20012 ( .A(n20263), .B(n20272), .Z(n20265) );
  XNOR U20013 ( .A(n20274), .B(n20275), .Z(n20263) );
  AND U20014 ( .A(n169), .B(n20276), .Z(n20275) );
  XOR U20015 ( .A(p_input[81]), .B(n20274), .Z(n20276) );
  XNOR U20016 ( .A(n20277), .B(n20278), .Z(n20274) );
  AND U20017 ( .A(n173), .B(n20279), .Z(n20278) );
  XOR U20018 ( .A(n20280), .B(n20281), .Z(n20272) );
  AND U20019 ( .A(n177), .B(n20271), .Z(n20281) );
  XNOR U20020 ( .A(n20282), .B(n20269), .Z(n20271) );
  XOR U20021 ( .A(n20283), .B(n20284), .Z(n20269) );
  AND U20022 ( .A(n200), .B(n20285), .Z(n20284) );
  IV U20023 ( .A(n20280), .Z(n20282) );
  XOR U20024 ( .A(n20286), .B(n20287), .Z(n20280) );
  AND U20025 ( .A(n184), .B(n20279), .Z(n20287) );
  XNOR U20026 ( .A(n20277), .B(n20286), .Z(n20279) );
  XNOR U20027 ( .A(n20288), .B(n20289), .Z(n20277) );
  AND U20028 ( .A(n188), .B(n20290), .Z(n20289) );
  XOR U20029 ( .A(p_input[113]), .B(n20288), .Z(n20290) );
  XNOR U20030 ( .A(n20291), .B(n20292), .Z(n20288) );
  AND U20031 ( .A(n192), .B(n20293), .Z(n20292) );
  XOR U20032 ( .A(n20294), .B(n20295), .Z(n20286) );
  AND U20033 ( .A(n196), .B(n20285), .Z(n20295) );
  XNOR U20034 ( .A(n20296), .B(n20283), .Z(n20285) );
  XOR U20035 ( .A(n20297), .B(n20298), .Z(n20283) );
  AND U20036 ( .A(n219), .B(n20299), .Z(n20298) );
  IV U20037 ( .A(n20294), .Z(n20296) );
  XOR U20038 ( .A(n20300), .B(n20301), .Z(n20294) );
  AND U20039 ( .A(n203), .B(n20293), .Z(n20301) );
  XNOR U20040 ( .A(n20291), .B(n20300), .Z(n20293) );
  XNOR U20041 ( .A(n20302), .B(n20303), .Z(n20291) );
  AND U20042 ( .A(n207), .B(n20304), .Z(n20303) );
  XOR U20043 ( .A(p_input[145]), .B(n20302), .Z(n20304) );
  XNOR U20044 ( .A(n20305), .B(n20306), .Z(n20302) );
  AND U20045 ( .A(n211), .B(n20307), .Z(n20306) );
  XOR U20046 ( .A(n20308), .B(n20309), .Z(n20300) );
  AND U20047 ( .A(n215), .B(n20299), .Z(n20309) );
  XNOR U20048 ( .A(n20310), .B(n20297), .Z(n20299) );
  XOR U20049 ( .A(n20311), .B(n20312), .Z(n20297) );
  AND U20050 ( .A(n238), .B(n20313), .Z(n20312) );
  IV U20051 ( .A(n20308), .Z(n20310) );
  XOR U20052 ( .A(n20314), .B(n20315), .Z(n20308) );
  AND U20053 ( .A(n222), .B(n20307), .Z(n20315) );
  XNOR U20054 ( .A(n20305), .B(n20314), .Z(n20307) );
  XNOR U20055 ( .A(n20316), .B(n20317), .Z(n20305) );
  AND U20056 ( .A(n226), .B(n20318), .Z(n20317) );
  XOR U20057 ( .A(p_input[177]), .B(n20316), .Z(n20318) );
  XNOR U20058 ( .A(n20319), .B(n20320), .Z(n20316) );
  AND U20059 ( .A(n230), .B(n20321), .Z(n20320) );
  XOR U20060 ( .A(n20322), .B(n20323), .Z(n20314) );
  AND U20061 ( .A(n234), .B(n20313), .Z(n20323) );
  XNOR U20062 ( .A(n20324), .B(n20311), .Z(n20313) );
  XOR U20063 ( .A(n20325), .B(n20326), .Z(n20311) );
  AND U20064 ( .A(n257), .B(n20327), .Z(n20326) );
  IV U20065 ( .A(n20322), .Z(n20324) );
  XOR U20066 ( .A(n20328), .B(n20329), .Z(n20322) );
  AND U20067 ( .A(n241), .B(n20321), .Z(n20329) );
  XNOR U20068 ( .A(n20319), .B(n20328), .Z(n20321) );
  XNOR U20069 ( .A(n20330), .B(n20331), .Z(n20319) );
  AND U20070 ( .A(n245), .B(n20332), .Z(n20331) );
  XOR U20071 ( .A(p_input[209]), .B(n20330), .Z(n20332) );
  XNOR U20072 ( .A(n20333), .B(n20334), .Z(n20330) );
  AND U20073 ( .A(n249), .B(n20335), .Z(n20334) );
  XOR U20074 ( .A(n20336), .B(n20337), .Z(n20328) );
  AND U20075 ( .A(n253), .B(n20327), .Z(n20337) );
  XNOR U20076 ( .A(n20338), .B(n20325), .Z(n20327) );
  XOR U20077 ( .A(n20339), .B(n20340), .Z(n20325) );
  AND U20078 ( .A(n276), .B(n20341), .Z(n20340) );
  IV U20079 ( .A(n20336), .Z(n20338) );
  XOR U20080 ( .A(n20342), .B(n20343), .Z(n20336) );
  AND U20081 ( .A(n260), .B(n20335), .Z(n20343) );
  XNOR U20082 ( .A(n20333), .B(n20342), .Z(n20335) );
  XNOR U20083 ( .A(n20344), .B(n20345), .Z(n20333) );
  AND U20084 ( .A(n264), .B(n20346), .Z(n20345) );
  XOR U20085 ( .A(p_input[241]), .B(n20344), .Z(n20346) );
  XNOR U20086 ( .A(n20347), .B(n20348), .Z(n20344) );
  AND U20087 ( .A(n268), .B(n20349), .Z(n20348) );
  XOR U20088 ( .A(n20350), .B(n20351), .Z(n20342) );
  AND U20089 ( .A(n272), .B(n20341), .Z(n20351) );
  XNOR U20090 ( .A(n20352), .B(n20339), .Z(n20341) );
  XOR U20091 ( .A(n20353), .B(n20354), .Z(n20339) );
  AND U20092 ( .A(n295), .B(n20355), .Z(n20354) );
  IV U20093 ( .A(n20350), .Z(n20352) );
  XOR U20094 ( .A(n20356), .B(n20357), .Z(n20350) );
  AND U20095 ( .A(n279), .B(n20349), .Z(n20357) );
  XNOR U20096 ( .A(n20347), .B(n20356), .Z(n20349) );
  XNOR U20097 ( .A(n20358), .B(n20359), .Z(n20347) );
  AND U20098 ( .A(n283), .B(n20360), .Z(n20359) );
  XOR U20099 ( .A(p_input[273]), .B(n20358), .Z(n20360) );
  XNOR U20100 ( .A(n20361), .B(n20362), .Z(n20358) );
  AND U20101 ( .A(n287), .B(n20363), .Z(n20362) );
  XOR U20102 ( .A(n20364), .B(n20365), .Z(n20356) );
  AND U20103 ( .A(n291), .B(n20355), .Z(n20365) );
  XNOR U20104 ( .A(n20366), .B(n20353), .Z(n20355) );
  XOR U20105 ( .A(n20367), .B(n20368), .Z(n20353) );
  AND U20106 ( .A(n314), .B(n20369), .Z(n20368) );
  IV U20107 ( .A(n20364), .Z(n20366) );
  XOR U20108 ( .A(n20370), .B(n20371), .Z(n20364) );
  AND U20109 ( .A(n298), .B(n20363), .Z(n20371) );
  XNOR U20110 ( .A(n20361), .B(n20370), .Z(n20363) );
  XNOR U20111 ( .A(n20372), .B(n20373), .Z(n20361) );
  AND U20112 ( .A(n302), .B(n20374), .Z(n20373) );
  XOR U20113 ( .A(p_input[305]), .B(n20372), .Z(n20374) );
  XNOR U20114 ( .A(n20375), .B(n20376), .Z(n20372) );
  AND U20115 ( .A(n306), .B(n20377), .Z(n20376) );
  XOR U20116 ( .A(n20378), .B(n20379), .Z(n20370) );
  AND U20117 ( .A(n310), .B(n20369), .Z(n20379) );
  XNOR U20118 ( .A(n20380), .B(n20367), .Z(n20369) );
  XOR U20119 ( .A(n20381), .B(n20382), .Z(n20367) );
  AND U20120 ( .A(n333), .B(n20383), .Z(n20382) );
  IV U20121 ( .A(n20378), .Z(n20380) );
  XOR U20122 ( .A(n20384), .B(n20385), .Z(n20378) );
  AND U20123 ( .A(n317), .B(n20377), .Z(n20385) );
  XNOR U20124 ( .A(n20375), .B(n20384), .Z(n20377) );
  XNOR U20125 ( .A(n20386), .B(n20387), .Z(n20375) );
  AND U20126 ( .A(n321), .B(n20388), .Z(n20387) );
  XOR U20127 ( .A(p_input[337]), .B(n20386), .Z(n20388) );
  XNOR U20128 ( .A(n20389), .B(n20390), .Z(n20386) );
  AND U20129 ( .A(n325), .B(n20391), .Z(n20390) );
  XOR U20130 ( .A(n20392), .B(n20393), .Z(n20384) );
  AND U20131 ( .A(n329), .B(n20383), .Z(n20393) );
  XNOR U20132 ( .A(n20394), .B(n20381), .Z(n20383) );
  XOR U20133 ( .A(n20395), .B(n20396), .Z(n20381) );
  AND U20134 ( .A(n352), .B(n20397), .Z(n20396) );
  IV U20135 ( .A(n20392), .Z(n20394) );
  XOR U20136 ( .A(n20398), .B(n20399), .Z(n20392) );
  AND U20137 ( .A(n336), .B(n20391), .Z(n20399) );
  XNOR U20138 ( .A(n20389), .B(n20398), .Z(n20391) );
  XNOR U20139 ( .A(n20400), .B(n20401), .Z(n20389) );
  AND U20140 ( .A(n340), .B(n20402), .Z(n20401) );
  XOR U20141 ( .A(p_input[369]), .B(n20400), .Z(n20402) );
  XNOR U20142 ( .A(n20403), .B(n20404), .Z(n20400) );
  AND U20143 ( .A(n344), .B(n20405), .Z(n20404) );
  XOR U20144 ( .A(n20406), .B(n20407), .Z(n20398) );
  AND U20145 ( .A(n348), .B(n20397), .Z(n20407) );
  XNOR U20146 ( .A(n20408), .B(n20395), .Z(n20397) );
  XOR U20147 ( .A(n20409), .B(n20410), .Z(n20395) );
  AND U20148 ( .A(n371), .B(n20411), .Z(n20410) );
  IV U20149 ( .A(n20406), .Z(n20408) );
  XOR U20150 ( .A(n20412), .B(n20413), .Z(n20406) );
  AND U20151 ( .A(n355), .B(n20405), .Z(n20413) );
  XNOR U20152 ( .A(n20403), .B(n20412), .Z(n20405) );
  XNOR U20153 ( .A(n20414), .B(n20415), .Z(n20403) );
  AND U20154 ( .A(n359), .B(n20416), .Z(n20415) );
  XOR U20155 ( .A(p_input[401]), .B(n20414), .Z(n20416) );
  XNOR U20156 ( .A(n20417), .B(n20418), .Z(n20414) );
  AND U20157 ( .A(n363), .B(n20419), .Z(n20418) );
  XOR U20158 ( .A(n20420), .B(n20421), .Z(n20412) );
  AND U20159 ( .A(n367), .B(n20411), .Z(n20421) );
  XNOR U20160 ( .A(n20422), .B(n20409), .Z(n20411) );
  XOR U20161 ( .A(n20423), .B(n20424), .Z(n20409) );
  AND U20162 ( .A(n390), .B(n20425), .Z(n20424) );
  IV U20163 ( .A(n20420), .Z(n20422) );
  XOR U20164 ( .A(n20426), .B(n20427), .Z(n20420) );
  AND U20165 ( .A(n374), .B(n20419), .Z(n20427) );
  XNOR U20166 ( .A(n20417), .B(n20426), .Z(n20419) );
  XNOR U20167 ( .A(n20428), .B(n20429), .Z(n20417) );
  AND U20168 ( .A(n378), .B(n20430), .Z(n20429) );
  XOR U20169 ( .A(p_input[433]), .B(n20428), .Z(n20430) );
  XNOR U20170 ( .A(n20431), .B(n20432), .Z(n20428) );
  AND U20171 ( .A(n382), .B(n20433), .Z(n20432) );
  XOR U20172 ( .A(n20434), .B(n20435), .Z(n20426) );
  AND U20173 ( .A(n386), .B(n20425), .Z(n20435) );
  XNOR U20174 ( .A(n20436), .B(n20423), .Z(n20425) );
  XOR U20175 ( .A(n20437), .B(n20438), .Z(n20423) );
  AND U20176 ( .A(n409), .B(n20439), .Z(n20438) );
  IV U20177 ( .A(n20434), .Z(n20436) );
  XOR U20178 ( .A(n20440), .B(n20441), .Z(n20434) );
  AND U20179 ( .A(n393), .B(n20433), .Z(n20441) );
  XNOR U20180 ( .A(n20431), .B(n20440), .Z(n20433) );
  XNOR U20181 ( .A(n20442), .B(n20443), .Z(n20431) );
  AND U20182 ( .A(n397), .B(n20444), .Z(n20443) );
  XOR U20183 ( .A(p_input[465]), .B(n20442), .Z(n20444) );
  XNOR U20184 ( .A(n20445), .B(n20446), .Z(n20442) );
  AND U20185 ( .A(n401), .B(n20447), .Z(n20446) );
  XOR U20186 ( .A(n20448), .B(n20449), .Z(n20440) );
  AND U20187 ( .A(n405), .B(n20439), .Z(n20449) );
  XNOR U20188 ( .A(n20450), .B(n20437), .Z(n20439) );
  XOR U20189 ( .A(n20451), .B(n20452), .Z(n20437) );
  AND U20190 ( .A(n428), .B(n20453), .Z(n20452) );
  IV U20191 ( .A(n20448), .Z(n20450) );
  XOR U20192 ( .A(n20454), .B(n20455), .Z(n20448) );
  AND U20193 ( .A(n412), .B(n20447), .Z(n20455) );
  XNOR U20194 ( .A(n20445), .B(n20454), .Z(n20447) );
  XNOR U20195 ( .A(n20456), .B(n20457), .Z(n20445) );
  AND U20196 ( .A(n416), .B(n20458), .Z(n20457) );
  XOR U20197 ( .A(p_input[497]), .B(n20456), .Z(n20458) );
  XNOR U20198 ( .A(n20459), .B(n20460), .Z(n20456) );
  AND U20199 ( .A(n420), .B(n20461), .Z(n20460) );
  XOR U20200 ( .A(n20462), .B(n20463), .Z(n20454) );
  AND U20201 ( .A(n424), .B(n20453), .Z(n20463) );
  XNOR U20202 ( .A(n20464), .B(n20451), .Z(n20453) );
  XOR U20203 ( .A(n20465), .B(n20466), .Z(n20451) );
  AND U20204 ( .A(n447), .B(n20467), .Z(n20466) );
  IV U20205 ( .A(n20462), .Z(n20464) );
  XOR U20206 ( .A(n20468), .B(n20469), .Z(n20462) );
  AND U20207 ( .A(n431), .B(n20461), .Z(n20469) );
  XNOR U20208 ( .A(n20459), .B(n20468), .Z(n20461) );
  XNOR U20209 ( .A(n20470), .B(n20471), .Z(n20459) );
  AND U20210 ( .A(n435), .B(n20472), .Z(n20471) );
  XOR U20211 ( .A(p_input[529]), .B(n20470), .Z(n20472) );
  XNOR U20212 ( .A(n20473), .B(n20474), .Z(n20470) );
  AND U20213 ( .A(n439), .B(n20475), .Z(n20474) );
  XOR U20214 ( .A(n20476), .B(n20477), .Z(n20468) );
  AND U20215 ( .A(n443), .B(n20467), .Z(n20477) );
  XNOR U20216 ( .A(n20478), .B(n20465), .Z(n20467) );
  XOR U20217 ( .A(n20479), .B(n20480), .Z(n20465) );
  AND U20218 ( .A(n466), .B(n20481), .Z(n20480) );
  IV U20219 ( .A(n20476), .Z(n20478) );
  XOR U20220 ( .A(n20482), .B(n20483), .Z(n20476) );
  AND U20221 ( .A(n450), .B(n20475), .Z(n20483) );
  XNOR U20222 ( .A(n20473), .B(n20482), .Z(n20475) );
  XNOR U20223 ( .A(n20484), .B(n20485), .Z(n20473) );
  AND U20224 ( .A(n454), .B(n20486), .Z(n20485) );
  XOR U20225 ( .A(p_input[561]), .B(n20484), .Z(n20486) );
  XNOR U20226 ( .A(n20487), .B(n20488), .Z(n20484) );
  AND U20227 ( .A(n458), .B(n20489), .Z(n20488) );
  XOR U20228 ( .A(n20490), .B(n20491), .Z(n20482) );
  AND U20229 ( .A(n462), .B(n20481), .Z(n20491) );
  XNOR U20230 ( .A(n20492), .B(n20479), .Z(n20481) );
  XOR U20231 ( .A(n20493), .B(n20494), .Z(n20479) );
  AND U20232 ( .A(n485), .B(n20495), .Z(n20494) );
  IV U20233 ( .A(n20490), .Z(n20492) );
  XOR U20234 ( .A(n20496), .B(n20497), .Z(n20490) );
  AND U20235 ( .A(n469), .B(n20489), .Z(n20497) );
  XNOR U20236 ( .A(n20487), .B(n20496), .Z(n20489) );
  XNOR U20237 ( .A(n20498), .B(n20499), .Z(n20487) );
  AND U20238 ( .A(n473), .B(n20500), .Z(n20499) );
  XOR U20239 ( .A(p_input[593]), .B(n20498), .Z(n20500) );
  XNOR U20240 ( .A(n20501), .B(n20502), .Z(n20498) );
  AND U20241 ( .A(n477), .B(n20503), .Z(n20502) );
  XOR U20242 ( .A(n20504), .B(n20505), .Z(n20496) );
  AND U20243 ( .A(n481), .B(n20495), .Z(n20505) );
  XNOR U20244 ( .A(n20506), .B(n20493), .Z(n20495) );
  XOR U20245 ( .A(n20507), .B(n20508), .Z(n20493) );
  AND U20246 ( .A(n504), .B(n20509), .Z(n20508) );
  IV U20247 ( .A(n20504), .Z(n20506) );
  XOR U20248 ( .A(n20510), .B(n20511), .Z(n20504) );
  AND U20249 ( .A(n488), .B(n20503), .Z(n20511) );
  XNOR U20250 ( .A(n20501), .B(n20510), .Z(n20503) );
  XNOR U20251 ( .A(n20512), .B(n20513), .Z(n20501) );
  AND U20252 ( .A(n492), .B(n20514), .Z(n20513) );
  XOR U20253 ( .A(p_input[625]), .B(n20512), .Z(n20514) );
  XNOR U20254 ( .A(n20515), .B(n20516), .Z(n20512) );
  AND U20255 ( .A(n496), .B(n20517), .Z(n20516) );
  XOR U20256 ( .A(n20518), .B(n20519), .Z(n20510) );
  AND U20257 ( .A(n500), .B(n20509), .Z(n20519) );
  XNOR U20258 ( .A(n20520), .B(n20507), .Z(n20509) );
  XOR U20259 ( .A(n20521), .B(n20522), .Z(n20507) );
  AND U20260 ( .A(n523), .B(n20523), .Z(n20522) );
  IV U20261 ( .A(n20518), .Z(n20520) );
  XOR U20262 ( .A(n20524), .B(n20525), .Z(n20518) );
  AND U20263 ( .A(n507), .B(n20517), .Z(n20525) );
  XNOR U20264 ( .A(n20515), .B(n20524), .Z(n20517) );
  XNOR U20265 ( .A(n20526), .B(n20527), .Z(n20515) );
  AND U20266 ( .A(n511), .B(n20528), .Z(n20527) );
  XOR U20267 ( .A(p_input[657]), .B(n20526), .Z(n20528) );
  XNOR U20268 ( .A(n20529), .B(n20530), .Z(n20526) );
  AND U20269 ( .A(n515), .B(n20531), .Z(n20530) );
  XOR U20270 ( .A(n20532), .B(n20533), .Z(n20524) );
  AND U20271 ( .A(n519), .B(n20523), .Z(n20533) );
  XNOR U20272 ( .A(n20534), .B(n20521), .Z(n20523) );
  XOR U20273 ( .A(n20535), .B(n20536), .Z(n20521) );
  AND U20274 ( .A(n542), .B(n20537), .Z(n20536) );
  IV U20275 ( .A(n20532), .Z(n20534) );
  XOR U20276 ( .A(n20538), .B(n20539), .Z(n20532) );
  AND U20277 ( .A(n526), .B(n20531), .Z(n20539) );
  XNOR U20278 ( .A(n20529), .B(n20538), .Z(n20531) );
  XNOR U20279 ( .A(n20540), .B(n20541), .Z(n20529) );
  AND U20280 ( .A(n530), .B(n20542), .Z(n20541) );
  XOR U20281 ( .A(p_input[689]), .B(n20540), .Z(n20542) );
  XNOR U20282 ( .A(n20543), .B(n20544), .Z(n20540) );
  AND U20283 ( .A(n534), .B(n20545), .Z(n20544) );
  XOR U20284 ( .A(n20546), .B(n20547), .Z(n20538) );
  AND U20285 ( .A(n538), .B(n20537), .Z(n20547) );
  XNOR U20286 ( .A(n20548), .B(n20535), .Z(n20537) );
  XOR U20287 ( .A(n20549), .B(n20550), .Z(n20535) );
  AND U20288 ( .A(n561), .B(n20551), .Z(n20550) );
  IV U20289 ( .A(n20546), .Z(n20548) );
  XOR U20290 ( .A(n20552), .B(n20553), .Z(n20546) );
  AND U20291 ( .A(n545), .B(n20545), .Z(n20553) );
  XNOR U20292 ( .A(n20543), .B(n20552), .Z(n20545) );
  XNOR U20293 ( .A(n20554), .B(n20555), .Z(n20543) );
  AND U20294 ( .A(n549), .B(n20556), .Z(n20555) );
  XOR U20295 ( .A(p_input[721]), .B(n20554), .Z(n20556) );
  XNOR U20296 ( .A(n20557), .B(n20558), .Z(n20554) );
  AND U20297 ( .A(n553), .B(n20559), .Z(n20558) );
  XOR U20298 ( .A(n20560), .B(n20561), .Z(n20552) );
  AND U20299 ( .A(n557), .B(n20551), .Z(n20561) );
  XNOR U20300 ( .A(n20562), .B(n20549), .Z(n20551) );
  XOR U20301 ( .A(n20563), .B(n20564), .Z(n20549) );
  AND U20302 ( .A(n580), .B(n20565), .Z(n20564) );
  IV U20303 ( .A(n20560), .Z(n20562) );
  XOR U20304 ( .A(n20566), .B(n20567), .Z(n20560) );
  AND U20305 ( .A(n564), .B(n20559), .Z(n20567) );
  XNOR U20306 ( .A(n20557), .B(n20566), .Z(n20559) );
  XNOR U20307 ( .A(n20568), .B(n20569), .Z(n20557) );
  AND U20308 ( .A(n568), .B(n20570), .Z(n20569) );
  XOR U20309 ( .A(p_input[753]), .B(n20568), .Z(n20570) );
  XNOR U20310 ( .A(n20571), .B(n20572), .Z(n20568) );
  AND U20311 ( .A(n572), .B(n20573), .Z(n20572) );
  XOR U20312 ( .A(n20574), .B(n20575), .Z(n20566) );
  AND U20313 ( .A(n576), .B(n20565), .Z(n20575) );
  XNOR U20314 ( .A(n20576), .B(n20563), .Z(n20565) );
  XOR U20315 ( .A(n20577), .B(n20578), .Z(n20563) );
  AND U20316 ( .A(n599), .B(n20579), .Z(n20578) );
  IV U20317 ( .A(n20574), .Z(n20576) );
  XOR U20318 ( .A(n20580), .B(n20581), .Z(n20574) );
  AND U20319 ( .A(n583), .B(n20573), .Z(n20581) );
  XNOR U20320 ( .A(n20571), .B(n20580), .Z(n20573) );
  XNOR U20321 ( .A(n20582), .B(n20583), .Z(n20571) );
  AND U20322 ( .A(n587), .B(n20584), .Z(n20583) );
  XOR U20323 ( .A(p_input[785]), .B(n20582), .Z(n20584) );
  XNOR U20324 ( .A(n20585), .B(n20586), .Z(n20582) );
  AND U20325 ( .A(n591), .B(n20587), .Z(n20586) );
  XOR U20326 ( .A(n20588), .B(n20589), .Z(n20580) );
  AND U20327 ( .A(n595), .B(n20579), .Z(n20589) );
  XNOR U20328 ( .A(n20590), .B(n20577), .Z(n20579) );
  XOR U20329 ( .A(n20591), .B(n20592), .Z(n20577) );
  AND U20330 ( .A(n618), .B(n20593), .Z(n20592) );
  IV U20331 ( .A(n20588), .Z(n20590) );
  XOR U20332 ( .A(n20594), .B(n20595), .Z(n20588) );
  AND U20333 ( .A(n602), .B(n20587), .Z(n20595) );
  XNOR U20334 ( .A(n20585), .B(n20594), .Z(n20587) );
  XNOR U20335 ( .A(n20596), .B(n20597), .Z(n20585) );
  AND U20336 ( .A(n606), .B(n20598), .Z(n20597) );
  XOR U20337 ( .A(p_input[817]), .B(n20596), .Z(n20598) );
  XNOR U20338 ( .A(n20599), .B(n20600), .Z(n20596) );
  AND U20339 ( .A(n610), .B(n20601), .Z(n20600) );
  XOR U20340 ( .A(n20602), .B(n20603), .Z(n20594) );
  AND U20341 ( .A(n614), .B(n20593), .Z(n20603) );
  XNOR U20342 ( .A(n20604), .B(n20591), .Z(n20593) );
  XOR U20343 ( .A(n20605), .B(n20606), .Z(n20591) );
  AND U20344 ( .A(n637), .B(n20607), .Z(n20606) );
  IV U20345 ( .A(n20602), .Z(n20604) );
  XOR U20346 ( .A(n20608), .B(n20609), .Z(n20602) );
  AND U20347 ( .A(n621), .B(n20601), .Z(n20609) );
  XNOR U20348 ( .A(n20599), .B(n20608), .Z(n20601) );
  XNOR U20349 ( .A(n20610), .B(n20611), .Z(n20599) );
  AND U20350 ( .A(n625), .B(n20612), .Z(n20611) );
  XOR U20351 ( .A(p_input[849]), .B(n20610), .Z(n20612) );
  XNOR U20352 ( .A(n20613), .B(n20614), .Z(n20610) );
  AND U20353 ( .A(n629), .B(n20615), .Z(n20614) );
  XOR U20354 ( .A(n20616), .B(n20617), .Z(n20608) );
  AND U20355 ( .A(n633), .B(n20607), .Z(n20617) );
  XNOR U20356 ( .A(n20618), .B(n20605), .Z(n20607) );
  XOR U20357 ( .A(n20619), .B(n20620), .Z(n20605) );
  AND U20358 ( .A(n656), .B(n20621), .Z(n20620) );
  IV U20359 ( .A(n20616), .Z(n20618) );
  XOR U20360 ( .A(n20622), .B(n20623), .Z(n20616) );
  AND U20361 ( .A(n640), .B(n20615), .Z(n20623) );
  XNOR U20362 ( .A(n20613), .B(n20622), .Z(n20615) );
  XNOR U20363 ( .A(n20624), .B(n20625), .Z(n20613) );
  AND U20364 ( .A(n644), .B(n20626), .Z(n20625) );
  XOR U20365 ( .A(p_input[881]), .B(n20624), .Z(n20626) );
  XNOR U20366 ( .A(n20627), .B(n20628), .Z(n20624) );
  AND U20367 ( .A(n648), .B(n20629), .Z(n20628) );
  XOR U20368 ( .A(n20630), .B(n20631), .Z(n20622) );
  AND U20369 ( .A(n652), .B(n20621), .Z(n20631) );
  XNOR U20370 ( .A(n20632), .B(n20619), .Z(n20621) );
  XOR U20371 ( .A(n20633), .B(n20634), .Z(n20619) );
  AND U20372 ( .A(n675), .B(n20635), .Z(n20634) );
  IV U20373 ( .A(n20630), .Z(n20632) );
  XOR U20374 ( .A(n20636), .B(n20637), .Z(n20630) );
  AND U20375 ( .A(n659), .B(n20629), .Z(n20637) );
  XNOR U20376 ( .A(n20627), .B(n20636), .Z(n20629) );
  XNOR U20377 ( .A(n20638), .B(n20639), .Z(n20627) );
  AND U20378 ( .A(n663), .B(n20640), .Z(n20639) );
  XOR U20379 ( .A(p_input[913]), .B(n20638), .Z(n20640) );
  XNOR U20380 ( .A(n20641), .B(n20642), .Z(n20638) );
  AND U20381 ( .A(n667), .B(n20643), .Z(n20642) );
  XOR U20382 ( .A(n20644), .B(n20645), .Z(n20636) );
  AND U20383 ( .A(n671), .B(n20635), .Z(n20645) );
  XNOR U20384 ( .A(n20646), .B(n20633), .Z(n20635) );
  XOR U20385 ( .A(n20647), .B(n20648), .Z(n20633) );
  AND U20386 ( .A(n694), .B(n20649), .Z(n20648) );
  IV U20387 ( .A(n20644), .Z(n20646) );
  XOR U20388 ( .A(n20650), .B(n20651), .Z(n20644) );
  AND U20389 ( .A(n678), .B(n20643), .Z(n20651) );
  XNOR U20390 ( .A(n20641), .B(n20650), .Z(n20643) );
  XNOR U20391 ( .A(n20652), .B(n20653), .Z(n20641) );
  AND U20392 ( .A(n682), .B(n20654), .Z(n20653) );
  XOR U20393 ( .A(p_input[945]), .B(n20652), .Z(n20654) );
  XNOR U20394 ( .A(n20655), .B(n20656), .Z(n20652) );
  AND U20395 ( .A(n686), .B(n20657), .Z(n20656) );
  XOR U20396 ( .A(n20658), .B(n20659), .Z(n20650) );
  AND U20397 ( .A(n690), .B(n20649), .Z(n20659) );
  XNOR U20398 ( .A(n20660), .B(n20647), .Z(n20649) );
  XOR U20399 ( .A(n20661), .B(n20662), .Z(n20647) );
  AND U20400 ( .A(n713), .B(n20663), .Z(n20662) );
  IV U20401 ( .A(n20658), .Z(n20660) );
  XOR U20402 ( .A(n20664), .B(n20665), .Z(n20658) );
  AND U20403 ( .A(n697), .B(n20657), .Z(n20665) );
  XNOR U20404 ( .A(n20655), .B(n20664), .Z(n20657) );
  XNOR U20405 ( .A(n20666), .B(n20667), .Z(n20655) );
  AND U20406 ( .A(n701), .B(n20668), .Z(n20667) );
  XOR U20407 ( .A(p_input[977]), .B(n20666), .Z(n20668) );
  XNOR U20408 ( .A(n20669), .B(n20670), .Z(n20666) );
  AND U20409 ( .A(n705), .B(n20671), .Z(n20670) );
  XOR U20410 ( .A(n20672), .B(n20673), .Z(n20664) );
  AND U20411 ( .A(n709), .B(n20663), .Z(n20673) );
  XNOR U20412 ( .A(n20674), .B(n20661), .Z(n20663) );
  XOR U20413 ( .A(n20675), .B(n20676), .Z(n20661) );
  AND U20414 ( .A(n732), .B(n20677), .Z(n20676) );
  IV U20415 ( .A(n20672), .Z(n20674) );
  XOR U20416 ( .A(n20678), .B(n20679), .Z(n20672) );
  AND U20417 ( .A(n716), .B(n20671), .Z(n20679) );
  XNOR U20418 ( .A(n20669), .B(n20678), .Z(n20671) );
  XNOR U20419 ( .A(n20680), .B(n20681), .Z(n20669) );
  AND U20420 ( .A(n720), .B(n20682), .Z(n20681) );
  XOR U20421 ( .A(p_input[1009]), .B(n20680), .Z(n20682) );
  XNOR U20422 ( .A(n20683), .B(n20684), .Z(n20680) );
  AND U20423 ( .A(n724), .B(n20685), .Z(n20684) );
  XOR U20424 ( .A(n20686), .B(n20687), .Z(n20678) );
  AND U20425 ( .A(n728), .B(n20677), .Z(n20687) );
  XNOR U20426 ( .A(n20688), .B(n20675), .Z(n20677) );
  XOR U20427 ( .A(n20689), .B(n20690), .Z(n20675) );
  AND U20428 ( .A(n751), .B(n20691), .Z(n20690) );
  IV U20429 ( .A(n20686), .Z(n20688) );
  XOR U20430 ( .A(n20692), .B(n20693), .Z(n20686) );
  AND U20431 ( .A(n735), .B(n20685), .Z(n20693) );
  XNOR U20432 ( .A(n20683), .B(n20692), .Z(n20685) );
  XNOR U20433 ( .A(n20694), .B(n20695), .Z(n20683) );
  AND U20434 ( .A(n739), .B(n20696), .Z(n20695) );
  XOR U20435 ( .A(p_input[1041]), .B(n20694), .Z(n20696) );
  XNOR U20436 ( .A(n20697), .B(n20698), .Z(n20694) );
  AND U20437 ( .A(n743), .B(n20699), .Z(n20698) );
  XOR U20438 ( .A(n20700), .B(n20701), .Z(n20692) );
  AND U20439 ( .A(n747), .B(n20691), .Z(n20701) );
  XNOR U20440 ( .A(n20702), .B(n20689), .Z(n20691) );
  XOR U20441 ( .A(n20703), .B(n20704), .Z(n20689) );
  AND U20442 ( .A(n770), .B(n20705), .Z(n20704) );
  IV U20443 ( .A(n20700), .Z(n20702) );
  XOR U20444 ( .A(n20706), .B(n20707), .Z(n20700) );
  AND U20445 ( .A(n754), .B(n20699), .Z(n20707) );
  XNOR U20446 ( .A(n20697), .B(n20706), .Z(n20699) );
  XNOR U20447 ( .A(n20708), .B(n20709), .Z(n20697) );
  AND U20448 ( .A(n758), .B(n20710), .Z(n20709) );
  XOR U20449 ( .A(p_input[1073]), .B(n20708), .Z(n20710) );
  XNOR U20450 ( .A(n20711), .B(n20712), .Z(n20708) );
  AND U20451 ( .A(n762), .B(n20713), .Z(n20712) );
  XOR U20452 ( .A(n20714), .B(n20715), .Z(n20706) );
  AND U20453 ( .A(n766), .B(n20705), .Z(n20715) );
  XNOR U20454 ( .A(n20716), .B(n20703), .Z(n20705) );
  XOR U20455 ( .A(n20717), .B(n20718), .Z(n20703) );
  AND U20456 ( .A(n789), .B(n20719), .Z(n20718) );
  IV U20457 ( .A(n20714), .Z(n20716) );
  XOR U20458 ( .A(n20720), .B(n20721), .Z(n20714) );
  AND U20459 ( .A(n773), .B(n20713), .Z(n20721) );
  XNOR U20460 ( .A(n20711), .B(n20720), .Z(n20713) );
  XNOR U20461 ( .A(n20722), .B(n20723), .Z(n20711) );
  AND U20462 ( .A(n777), .B(n20724), .Z(n20723) );
  XOR U20463 ( .A(p_input[1105]), .B(n20722), .Z(n20724) );
  XNOR U20464 ( .A(n20725), .B(n20726), .Z(n20722) );
  AND U20465 ( .A(n781), .B(n20727), .Z(n20726) );
  XOR U20466 ( .A(n20728), .B(n20729), .Z(n20720) );
  AND U20467 ( .A(n785), .B(n20719), .Z(n20729) );
  XNOR U20468 ( .A(n20730), .B(n20717), .Z(n20719) );
  XOR U20469 ( .A(n20731), .B(n20732), .Z(n20717) );
  AND U20470 ( .A(n808), .B(n20733), .Z(n20732) );
  IV U20471 ( .A(n20728), .Z(n20730) );
  XOR U20472 ( .A(n20734), .B(n20735), .Z(n20728) );
  AND U20473 ( .A(n792), .B(n20727), .Z(n20735) );
  XNOR U20474 ( .A(n20725), .B(n20734), .Z(n20727) );
  XNOR U20475 ( .A(n20736), .B(n20737), .Z(n20725) );
  AND U20476 ( .A(n796), .B(n20738), .Z(n20737) );
  XOR U20477 ( .A(p_input[1137]), .B(n20736), .Z(n20738) );
  XNOR U20478 ( .A(n20739), .B(n20740), .Z(n20736) );
  AND U20479 ( .A(n800), .B(n20741), .Z(n20740) );
  XOR U20480 ( .A(n20742), .B(n20743), .Z(n20734) );
  AND U20481 ( .A(n804), .B(n20733), .Z(n20743) );
  XNOR U20482 ( .A(n20744), .B(n20731), .Z(n20733) );
  XOR U20483 ( .A(n20745), .B(n20746), .Z(n20731) );
  AND U20484 ( .A(n827), .B(n20747), .Z(n20746) );
  IV U20485 ( .A(n20742), .Z(n20744) );
  XOR U20486 ( .A(n20748), .B(n20749), .Z(n20742) );
  AND U20487 ( .A(n811), .B(n20741), .Z(n20749) );
  XNOR U20488 ( .A(n20739), .B(n20748), .Z(n20741) );
  XNOR U20489 ( .A(n20750), .B(n20751), .Z(n20739) );
  AND U20490 ( .A(n815), .B(n20752), .Z(n20751) );
  XOR U20491 ( .A(p_input[1169]), .B(n20750), .Z(n20752) );
  XNOR U20492 ( .A(n20753), .B(n20754), .Z(n20750) );
  AND U20493 ( .A(n819), .B(n20755), .Z(n20754) );
  XOR U20494 ( .A(n20756), .B(n20757), .Z(n20748) );
  AND U20495 ( .A(n823), .B(n20747), .Z(n20757) );
  XNOR U20496 ( .A(n20758), .B(n20745), .Z(n20747) );
  XOR U20497 ( .A(n20759), .B(n20760), .Z(n20745) );
  AND U20498 ( .A(n846), .B(n20761), .Z(n20760) );
  IV U20499 ( .A(n20756), .Z(n20758) );
  XOR U20500 ( .A(n20762), .B(n20763), .Z(n20756) );
  AND U20501 ( .A(n830), .B(n20755), .Z(n20763) );
  XNOR U20502 ( .A(n20753), .B(n20762), .Z(n20755) );
  XNOR U20503 ( .A(n20764), .B(n20765), .Z(n20753) );
  AND U20504 ( .A(n834), .B(n20766), .Z(n20765) );
  XOR U20505 ( .A(p_input[1201]), .B(n20764), .Z(n20766) );
  XNOR U20506 ( .A(n20767), .B(n20768), .Z(n20764) );
  AND U20507 ( .A(n838), .B(n20769), .Z(n20768) );
  XOR U20508 ( .A(n20770), .B(n20771), .Z(n20762) );
  AND U20509 ( .A(n842), .B(n20761), .Z(n20771) );
  XNOR U20510 ( .A(n20772), .B(n20759), .Z(n20761) );
  XOR U20511 ( .A(n20773), .B(n20774), .Z(n20759) );
  AND U20512 ( .A(n865), .B(n20775), .Z(n20774) );
  IV U20513 ( .A(n20770), .Z(n20772) );
  XOR U20514 ( .A(n20776), .B(n20777), .Z(n20770) );
  AND U20515 ( .A(n849), .B(n20769), .Z(n20777) );
  XNOR U20516 ( .A(n20767), .B(n20776), .Z(n20769) );
  XNOR U20517 ( .A(n20778), .B(n20779), .Z(n20767) );
  AND U20518 ( .A(n853), .B(n20780), .Z(n20779) );
  XOR U20519 ( .A(p_input[1233]), .B(n20778), .Z(n20780) );
  XNOR U20520 ( .A(n20781), .B(n20782), .Z(n20778) );
  AND U20521 ( .A(n857), .B(n20783), .Z(n20782) );
  XOR U20522 ( .A(n20784), .B(n20785), .Z(n20776) );
  AND U20523 ( .A(n861), .B(n20775), .Z(n20785) );
  XNOR U20524 ( .A(n20786), .B(n20773), .Z(n20775) );
  XOR U20525 ( .A(n20787), .B(n20788), .Z(n20773) );
  AND U20526 ( .A(n884), .B(n20789), .Z(n20788) );
  IV U20527 ( .A(n20784), .Z(n20786) );
  XOR U20528 ( .A(n20790), .B(n20791), .Z(n20784) );
  AND U20529 ( .A(n868), .B(n20783), .Z(n20791) );
  XNOR U20530 ( .A(n20781), .B(n20790), .Z(n20783) );
  XNOR U20531 ( .A(n20792), .B(n20793), .Z(n20781) );
  AND U20532 ( .A(n872), .B(n20794), .Z(n20793) );
  XOR U20533 ( .A(p_input[1265]), .B(n20792), .Z(n20794) );
  XNOR U20534 ( .A(n20795), .B(n20796), .Z(n20792) );
  AND U20535 ( .A(n876), .B(n20797), .Z(n20796) );
  XOR U20536 ( .A(n20798), .B(n20799), .Z(n20790) );
  AND U20537 ( .A(n880), .B(n20789), .Z(n20799) );
  XNOR U20538 ( .A(n20800), .B(n20787), .Z(n20789) );
  XOR U20539 ( .A(n20801), .B(n20802), .Z(n20787) );
  AND U20540 ( .A(n903), .B(n20803), .Z(n20802) );
  IV U20541 ( .A(n20798), .Z(n20800) );
  XOR U20542 ( .A(n20804), .B(n20805), .Z(n20798) );
  AND U20543 ( .A(n887), .B(n20797), .Z(n20805) );
  XNOR U20544 ( .A(n20795), .B(n20804), .Z(n20797) );
  XNOR U20545 ( .A(n20806), .B(n20807), .Z(n20795) );
  AND U20546 ( .A(n891), .B(n20808), .Z(n20807) );
  XOR U20547 ( .A(p_input[1297]), .B(n20806), .Z(n20808) );
  XNOR U20548 ( .A(n20809), .B(n20810), .Z(n20806) );
  AND U20549 ( .A(n895), .B(n20811), .Z(n20810) );
  XOR U20550 ( .A(n20812), .B(n20813), .Z(n20804) );
  AND U20551 ( .A(n899), .B(n20803), .Z(n20813) );
  XNOR U20552 ( .A(n20814), .B(n20801), .Z(n20803) );
  XOR U20553 ( .A(n20815), .B(n20816), .Z(n20801) );
  AND U20554 ( .A(n922), .B(n20817), .Z(n20816) );
  IV U20555 ( .A(n20812), .Z(n20814) );
  XOR U20556 ( .A(n20818), .B(n20819), .Z(n20812) );
  AND U20557 ( .A(n906), .B(n20811), .Z(n20819) );
  XNOR U20558 ( .A(n20809), .B(n20818), .Z(n20811) );
  XNOR U20559 ( .A(n20820), .B(n20821), .Z(n20809) );
  AND U20560 ( .A(n910), .B(n20822), .Z(n20821) );
  XOR U20561 ( .A(p_input[1329]), .B(n20820), .Z(n20822) );
  XNOR U20562 ( .A(n20823), .B(n20824), .Z(n20820) );
  AND U20563 ( .A(n914), .B(n20825), .Z(n20824) );
  XOR U20564 ( .A(n20826), .B(n20827), .Z(n20818) );
  AND U20565 ( .A(n918), .B(n20817), .Z(n20827) );
  XNOR U20566 ( .A(n20828), .B(n20815), .Z(n20817) );
  XOR U20567 ( .A(n20829), .B(n20830), .Z(n20815) );
  AND U20568 ( .A(n941), .B(n20831), .Z(n20830) );
  IV U20569 ( .A(n20826), .Z(n20828) );
  XOR U20570 ( .A(n20832), .B(n20833), .Z(n20826) );
  AND U20571 ( .A(n925), .B(n20825), .Z(n20833) );
  XNOR U20572 ( .A(n20823), .B(n20832), .Z(n20825) );
  XNOR U20573 ( .A(n20834), .B(n20835), .Z(n20823) );
  AND U20574 ( .A(n929), .B(n20836), .Z(n20835) );
  XOR U20575 ( .A(p_input[1361]), .B(n20834), .Z(n20836) );
  XNOR U20576 ( .A(n20837), .B(n20838), .Z(n20834) );
  AND U20577 ( .A(n933), .B(n20839), .Z(n20838) );
  XOR U20578 ( .A(n20840), .B(n20841), .Z(n20832) );
  AND U20579 ( .A(n937), .B(n20831), .Z(n20841) );
  XNOR U20580 ( .A(n20842), .B(n20829), .Z(n20831) );
  XOR U20581 ( .A(n20843), .B(n20844), .Z(n20829) );
  AND U20582 ( .A(n960), .B(n20845), .Z(n20844) );
  IV U20583 ( .A(n20840), .Z(n20842) );
  XOR U20584 ( .A(n20846), .B(n20847), .Z(n20840) );
  AND U20585 ( .A(n944), .B(n20839), .Z(n20847) );
  XNOR U20586 ( .A(n20837), .B(n20846), .Z(n20839) );
  XNOR U20587 ( .A(n20848), .B(n20849), .Z(n20837) );
  AND U20588 ( .A(n948), .B(n20850), .Z(n20849) );
  XOR U20589 ( .A(p_input[1393]), .B(n20848), .Z(n20850) );
  XNOR U20590 ( .A(n20851), .B(n20852), .Z(n20848) );
  AND U20591 ( .A(n952), .B(n20853), .Z(n20852) );
  XOR U20592 ( .A(n20854), .B(n20855), .Z(n20846) );
  AND U20593 ( .A(n956), .B(n20845), .Z(n20855) );
  XNOR U20594 ( .A(n20856), .B(n20843), .Z(n20845) );
  XOR U20595 ( .A(n20857), .B(n20858), .Z(n20843) );
  AND U20596 ( .A(n979), .B(n20859), .Z(n20858) );
  IV U20597 ( .A(n20854), .Z(n20856) );
  XOR U20598 ( .A(n20860), .B(n20861), .Z(n20854) );
  AND U20599 ( .A(n963), .B(n20853), .Z(n20861) );
  XNOR U20600 ( .A(n20851), .B(n20860), .Z(n20853) );
  XNOR U20601 ( .A(n20862), .B(n20863), .Z(n20851) );
  AND U20602 ( .A(n967), .B(n20864), .Z(n20863) );
  XOR U20603 ( .A(p_input[1425]), .B(n20862), .Z(n20864) );
  XNOR U20604 ( .A(n20865), .B(n20866), .Z(n20862) );
  AND U20605 ( .A(n971), .B(n20867), .Z(n20866) );
  XOR U20606 ( .A(n20868), .B(n20869), .Z(n20860) );
  AND U20607 ( .A(n975), .B(n20859), .Z(n20869) );
  XNOR U20608 ( .A(n20870), .B(n20857), .Z(n20859) );
  XOR U20609 ( .A(n20871), .B(n20872), .Z(n20857) );
  AND U20610 ( .A(n998), .B(n20873), .Z(n20872) );
  IV U20611 ( .A(n20868), .Z(n20870) );
  XOR U20612 ( .A(n20874), .B(n20875), .Z(n20868) );
  AND U20613 ( .A(n982), .B(n20867), .Z(n20875) );
  XNOR U20614 ( .A(n20865), .B(n20874), .Z(n20867) );
  XNOR U20615 ( .A(n20876), .B(n20877), .Z(n20865) );
  AND U20616 ( .A(n986), .B(n20878), .Z(n20877) );
  XOR U20617 ( .A(p_input[1457]), .B(n20876), .Z(n20878) );
  XNOR U20618 ( .A(n20879), .B(n20880), .Z(n20876) );
  AND U20619 ( .A(n990), .B(n20881), .Z(n20880) );
  XOR U20620 ( .A(n20882), .B(n20883), .Z(n20874) );
  AND U20621 ( .A(n994), .B(n20873), .Z(n20883) );
  XNOR U20622 ( .A(n20884), .B(n20871), .Z(n20873) );
  XOR U20623 ( .A(n20885), .B(n20886), .Z(n20871) );
  AND U20624 ( .A(n1017), .B(n20887), .Z(n20886) );
  IV U20625 ( .A(n20882), .Z(n20884) );
  XOR U20626 ( .A(n20888), .B(n20889), .Z(n20882) );
  AND U20627 ( .A(n1001), .B(n20881), .Z(n20889) );
  XNOR U20628 ( .A(n20879), .B(n20888), .Z(n20881) );
  XNOR U20629 ( .A(n20890), .B(n20891), .Z(n20879) );
  AND U20630 ( .A(n1005), .B(n20892), .Z(n20891) );
  XOR U20631 ( .A(p_input[1489]), .B(n20890), .Z(n20892) );
  XNOR U20632 ( .A(n20893), .B(n20894), .Z(n20890) );
  AND U20633 ( .A(n1009), .B(n20895), .Z(n20894) );
  XOR U20634 ( .A(n20896), .B(n20897), .Z(n20888) );
  AND U20635 ( .A(n1013), .B(n20887), .Z(n20897) );
  XNOR U20636 ( .A(n20898), .B(n20885), .Z(n20887) );
  XOR U20637 ( .A(n20899), .B(n20900), .Z(n20885) );
  AND U20638 ( .A(n1036), .B(n20901), .Z(n20900) );
  IV U20639 ( .A(n20896), .Z(n20898) );
  XOR U20640 ( .A(n20902), .B(n20903), .Z(n20896) );
  AND U20641 ( .A(n1020), .B(n20895), .Z(n20903) );
  XNOR U20642 ( .A(n20893), .B(n20902), .Z(n20895) );
  XNOR U20643 ( .A(n20904), .B(n20905), .Z(n20893) );
  AND U20644 ( .A(n1024), .B(n20906), .Z(n20905) );
  XOR U20645 ( .A(p_input[1521]), .B(n20904), .Z(n20906) );
  XNOR U20646 ( .A(n20907), .B(n20908), .Z(n20904) );
  AND U20647 ( .A(n1028), .B(n20909), .Z(n20908) );
  XOR U20648 ( .A(n20910), .B(n20911), .Z(n20902) );
  AND U20649 ( .A(n1032), .B(n20901), .Z(n20911) );
  XNOR U20650 ( .A(n20912), .B(n20899), .Z(n20901) );
  XOR U20651 ( .A(n20913), .B(n20914), .Z(n20899) );
  AND U20652 ( .A(n1055), .B(n20915), .Z(n20914) );
  IV U20653 ( .A(n20910), .Z(n20912) );
  XOR U20654 ( .A(n20916), .B(n20917), .Z(n20910) );
  AND U20655 ( .A(n1039), .B(n20909), .Z(n20917) );
  XNOR U20656 ( .A(n20907), .B(n20916), .Z(n20909) );
  XNOR U20657 ( .A(n20918), .B(n20919), .Z(n20907) );
  AND U20658 ( .A(n1043), .B(n20920), .Z(n20919) );
  XOR U20659 ( .A(p_input[1553]), .B(n20918), .Z(n20920) );
  XNOR U20660 ( .A(n20921), .B(n20922), .Z(n20918) );
  AND U20661 ( .A(n1047), .B(n20923), .Z(n20922) );
  XOR U20662 ( .A(n20924), .B(n20925), .Z(n20916) );
  AND U20663 ( .A(n1051), .B(n20915), .Z(n20925) );
  XNOR U20664 ( .A(n20926), .B(n20913), .Z(n20915) );
  XOR U20665 ( .A(n20927), .B(n20928), .Z(n20913) );
  AND U20666 ( .A(n1074), .B(n20929), .Z(n20928) );
  IV U20667 ( .A(n20924), .Z(n20926) );
  XOR U20668 ( .A(n20930), .B(n20931), .Z(n20924) );
  AND U20669 ( .A(n1058), .B(n20923), .Z(n20931) );
  XNOR U20670 ( .A(n20921), .B(n20930), .Z(n20923) );
  XNOR U20671 ( .A(n20932), .B(n20933), .Z(n20921) );
  AND U20672 ( .A(n1062), .B(n20934), .Z(n20933) );
  XOR U20673 ( .A(p_input[1585]), .B(n20932), .Z(n20934) );
  XNOR U20674 ( .A(n20935), .B(n20936), .Z(n20932) );
  AND U20675 ( .A(n1066), .B(n20937), .Z(n20936) );
  XOR U20676 ( .A(n20938), .B(n20939), .Z(n20930) );
  AND U20677 ( .A(n1070), .B(n20929), .Z(n20939) );
  XNOR U20678 ( .A(n20940), .B(n20927), .Z(n20929) );
  XOR U20679 ( .A(n20941), .B(n20942), .Z(n20927) );
  AND U20680 ( .A(n1093), .B(n20943), .Z(n20942) );
  IV U20681 ( .A(n20938), .Z(n20940) );
  XOR U20682 ( .A(n20944), .B(n20945), .Z(n20938) );
  AND U20683 ( .A(n1077), .B(n20937), .Z(n20945) );
  XNOR U20684 ( .A(n20935), .B(n20944), .Z(n20937) );
  XNOR U20685 ( .A(n20946), .B(n20947), .Z(n20935) );
  AND U20686 ( .A(n1081), .B(n20948), .Z(n20947) );
  XOR U20687 ( .A(p_input[1617]), .B(n20946), .Z(n20948) );
  XNOR U20688 ( .A(n20949), .B(n20950), .Z(n20946) );
  AND U20689 ( .A(n1085), .B(n20951), .Z(n20950) );
  XOR U20690 ( .A(n20952), .B(n20953), .Z(n20944) );
  AND U20691 ( .A(n1089), .B(n20943), .Z(n20953) );
  XNOR U20692 ( .A(n20954), .B(n20941), .Z(n20943) );
  XOR U20693 ( .A(n20955), .B(n20956), .Z(n20941) );
  AND U20694 ( .A(n1112), .B(n20957), .Z(n20956) );
  IV U20695 ( .A(n20952), .Z(n20954) );
  XOR U20696 ( .A(n20958), .B(n20959), .Z(n20952) );
  AND U20697 ( .A(n1096), .B(n20951), .Z(n20959) );
  XNOR U20698 ( .A(n20949), .B(n20958), .Z(n20951) );
  XNOR U20699 ( .A(n20960), .B(n20961), .Z(n20949) );
  AND U20700 ( .A(n1100), .B(n20962), .Z(n20961) );
  XOR U20701 ( .A(p_input[1649]), .B(n20960), .Z(n20962) );
  XNOR U20702 ( .A(n20963), .B(n20964), .Z(n20960) );
  AND U20703 ( .A(n1104), .B(n20965), .Z(n20964) );
  XOR U20704 ( .A(n20966), .B(n20967), .Z(n20958) );
  AND U20705 ( .A(n1108), .B(n20957), .Z(n20967) );
  XNOR U20706 ( .A(n20968), .B(n20955), .Z(n20957) );
  XOR U20707 ( .A(n20969), .B(n20970), .Z(n20955) );
  AND U20708 ( .A(n1131), .B(n20971), .Z(n20970) );
  IV U20709 ( .A(n20966), .Z(n20968) );
  XOR U20710 ( .A(n20972), .B(n20973), .Z(n20966) );
  AND U20711 ( .A(n1115), .B(n20965), .Z(n20973) );
  XNOR U20712 ( .A(n20963), .B(n20972), .Z(n20965) );
  XNOR U20713 ( .A(n20974), .B(n20975), .Z(n20963) );
  AND U20714 ( .A(n1119), .B(n20976), .Z(n20975) );
  XOR U20715 ( .A(p_input[1681]), .B(n20974), .Z(n20976) );
  XNOR U20716 ( .A(n20977), .B(n20978), .Z(n20974) );
  AND U20717 ( .A(n1123), .B(n20979), .Z(n20978) );
  XOR U20718 ( .A(n20980), .B(n20981), .Z(n20972) );
  AND U20719 ( .A(n1127), .B(n20971), .Z(n20981) );
  XNOR U20720 ( .A(n20982), .B(n20969), .Z(n20971) );
  XOR U20721 ( .A(n20983), .B(n20984), .Z(n20969) );
  AND U20722 ( .A(n1150), .B(n20985), .Z(n20984) );
  IV U20723 ( .A(n20980), .Z(n20982) );
  XOR U20724 ( .A(n20986), .B(n20987), .Z(n20980) );
  AND U20725 ( .A(n1134), .B(n20979), .Z(n20987) );
  XNOR U20726 ( .A(n20977), .B(n20986), .Z(n20979) );
  XNOR U20727 ( .A(n20988), .B(n20989), .Z(n20977) );
  AND U20728 ( .A(n1138), .B(n20990), .Z(n20989) );
  XOR U20729 ( .A(p_input[1713]), .B(n20988), .Z(n20990) );
  XNOR U20730 ( .A(n20991), .B(n20992), .Z(n20988) );
  AND U20731 ( .A(n1142), .B(n20993), .Z(n20992) );
  XOR U20732 ( .A(n20994), .B(n20995), .Z(n20986) );
  AND U20733 ( .A(n1146), .B(n20985), .Z(n20995) );
  XNOR U20734 ( .A(n20996), .B(n20983), .Z(n20985) );
  XOR U20735 ( .A(n20997), .B(n20998), .Z(n20983) );
  AND U20736 ( .A(n1169), .B(n20999), .Z(n20998) );
  IV U20737 ( .A(n20994), .Z(n20996) );
  XOR U20738 ( .A(n21000), .B(n21001), .Z(n20994) );
  AND U20739 ( .A(n1153), .B(n20993), .Z(n21001) );
  XNOR U20740 ( .A(n20991), .B(n21000), .Z(n20993) );
  XNOR U20741 ( .A(n21002), .B(n21003), .Z(n20991) );
  AND U20742 ( .A(n1157), .B(n21004), .Z(n21003) );
  XOR U20743 ( .A(p_input[1745]), .B(n21002), .Z(n21004) );
  XNOR U20744 ( .A(n21005), .B(n21006), .Z(n21002) );
  AND U20745 ( .A(n1161), .B(n21007), .Z(n21006) );
  XOR U20746 ( .A(n21008), .B(n21009), .Z(n21000) );
  AND U20747 ( .A(n1165), .B(n20999), .Z(n21009) );
  XNOR U20748 ( .A(n21010), .B(n20997), .Z(n20999) );
  XOR U20749 ( .A(n21011), .B(n21012), .Z(n20997) );
  AND U20750 ( .A(n1188), .B(n21013), .Z(n21012) );
  IV U20751 ( .A(n21008), .Z(n21010) );
  XOR U20752 ( .A(n21014), .B(n21015), .Z(n21008) );
  AND U20753 ( .A(n1172), .B(n21007), .Z(n21015) );
  XNOR U20754 ( .A(n21005), .B(n21014), .Z(n21007) );
  XNOR U20755 ( .A(n21016), .B(n21017), .Z(n21005) );
  AND U20756 ( .A(n1176), .B(n21018), .Z(n21017) );
  XOR U20757 ( .A(p_input[1777]), .B(n21016), .Z(n21018) );
  XNOR U20758 ( .A(n21019), .B(n21020), .Z(n21016) );
  AND U20759 ( .A(n1180), .B(n21021), .Z(n21020) );
  XOR U20760 ( .A(n21022), .B(n21023), .Z(n21014) );
  AND U20761 ( .A(n1184), .B(n21013), .Z(n21023) );
  XNOR U20762 ( .A(n21024), .B(n21011), .Z(n21013) );
  XOR U20763 ( .A(n21025), .B(n21026), .Z(n21011) );
  AND U20764 ( .A(n1207), .B(n21027), .Z(n21026) );
  IV U20765 ( .A(n21022), .Z(n21024) );
  XOR U20766 ( .A(n21028), .B(n21029), .Z(n21022) );
  AND U20767 ( .A(n1191), .B(n21021), .Z(n21029) );
  XNOR U20768 ( .A(n21019), .B(n21028), .Z(n21021) );
  XNOR U20769 ( .A(n21030), .B(n21031), .Z(n21019) );
  AND U20770 ( .A(n1195), .B(n21032), .Z(n21031) );
  XOR U20771 ( .A(p_input[1809]), .B(n21030), .Z(n21032) );
  XNOR U20772 ( .A(n21033), .B(n21034), .Z(n21030) );
  AND U20773 ( .A(n1199), .B(n21035), .Z(n21034) );
  XOR U20774 ( .A(n21036), .B(n21037), .Z(n21028) );
  AND U20775 ( .A(n1203), .B(n21027), .Z(n21037) );
  XNOR U20776 ( .A(n21038), .B(n21025), .Z(n21027) );
  XOR U20777 ( .A(n21039), .B(n21040), .Z(n21025) );
  AND U20778 ( .A(n1226), .B(n21041), .Z(n21040) );
  IV U20779 ( .A(n21036), .Z(n21038) );
  XOR U20780 ( .A(n21042), .B(n21043), .Z(n21036) );
  AND U20781 ( .A(n1210), .B(n21035), .Z(n21043) );
  XNOR U20782 ( .A(n21033), .B(n21042), .Z(n21035) );
  XNOR U20783 ( .A(n21044), .B(n21045), .Z(n21033) );
  AND U20784 ( .A(n1214), .B(n21046), .Z(n21045) );
  XOR U20785 ( .A(p_input[1841]), .B(n21044), .Z(n21046) );
  XNOR U20786 ( .A(n21047), .B(n21048), .Z(n21044) );
  AND U20787 ( .A(n1218), .B(n21049), .Z(n21048) );
  XOR U20788 ( .A(n21050), .B(n21051), .Z(n21042) );
  AND U20789 ( .A(n1222), .B(n21041), .Z(n21051) );
  XNOR U20790 ( .A(n21052), .B(n21039), .Z(n21041) );
  XOR U20791 ( .A(n21053), .B(n21054), .Z(n21039) );
  AND U20792 ( .A(n1245), .B(n21055), .Z(n21054) );
  IV U20793 ( .A(n21050), .Z(n21052) );
  XOR U20794 ( .A(n21056), .B(n21057), .Z(n21050) );
  AND U20795 ( .A(n1229), .B(n21049), .Z(n21057) );
  XNOR U20796 ( .A(n21047), .B(n21056), .Z(n21049) );
  XNOR U20797 ( .A(n21058), .B(n21059), .Z(n21047) );
  AND U20798 ( .A(n1233), .B(n21060), .Z(n21059) );
  XOR U20799 ( .A(p_input[1873]), .B(n21058), .Z(n21060) );
  XNOR U20800 ( .A(n21061), .B(n21062), .Z(n21058) );
  AND U20801 ( .A(n1237), .B(n21063), .Z(n21062) );
  XOR U20802 ( .A(n21064), .B(n21065), .Z(n21056) );
  AND U20803 ( .A(n1241), .B(n21055), .Z(n21065) );
  XNOR U20804 ( .A(n21066), .B(n21053), .Z(n21055) );
  XOR U20805 ( .A(n21067), .B(n21068), .Z(n21053) );
  AND U20806 ( .A(n1264), .B(n21069), .Z(n21068) );
  IV U20807 ( .A(n21064), .Z(n21066) );
  XOR U20808 ( .A(n21070), .B(n21071), .Z(n21064) );
  AND U20809 ( .A(n1248), .B(n21063), .Z(n21071) );
  XNOR U20810 ( .A(n21061), .B(n21070), .Z(n21063) );
  XNOR U20811 ( .A(n21072), .B(n21073), .Z(n21061) );
  AND U20812 ( .A(n1252), .B(n21074), .Z(n21073) );
  XOR U20813 ( .A(p_input[1905]), .B(n21072), .Z(n21074) );
  XNOR U20814 ( .A(n21075), .B(n21076), .Z(n21072) );
  AND U20815 ( .A(n1256), .B(n21077), .Z(n21076) );
  XOR U20816 ( .A(n21078), .B(n21079), .Z(n21070) );
  AND U20817 ( .A(n1260), .B(n21069), .Z(n21079) );
  XNOR U20818 ( .A(n21080), .B(n21067), .Z(n21069) );
  XOR U20819 ( .A(n21081), .B(n21082), .Z(n21067) );
  AND U20820 ( .A(n1282), .B(n21083), .Z(n21082) );
  IV U20821 ( .A(n21078), .Z(n21080) );
  XOR U20822 ( .A(n21084), .B(n21085), .Z(n21078) );
  AND U20823 ( .A(n1267), .B(n21077), .Z(n21085) );
  XNOR U20824 ( .A(n21075), .B(n21084), .Z(n21077) );
  XNOR U20825 ( .A(n21086), .B(n21087), .Z(n21075) );
  AND U20826 ( .A(n1271), .B(n21088), .Z(n21087) );
  XOR U20827 ( .A(p_input[1937]), .B(n21086), .Z(n21088) );
  XOR U20828 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][17] ), .B(n21089), 
        .Z(n21086) );
  AND U20829 ( .A(n1274), .B(n21090), .Z(n21089) );
  XOR U20830 ( .A(n21091), .B(n21092), .Z(n21084) );
  AND U20831 ( .A(n1278), .B(n21083), .Z(n21092) );
  XNOR U20832 ( .A(n21093), .B(n21081), .Z(n21083) );
  XOR U20833 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n21094), .Z(n21081) );
  AND U20834 ( .A(n1290), .B(n21095), .Z(n21094) );
  IV U20835 ( .A(n21091), .Z(n21093) );
  XOR U20836 ( .A(n21096), .B(n21097), .Z(n21091) );
  AND U20837 ( .A(n1285), .B(n21090), .Z(n21097) );
  XOR U20838 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][17] ), .B(n21096), 
        .Z(n21090) );
  XOR U20839 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .B(n21098), 
        .Z(n21096) );
  AND U20840 ( .A(n1287), .B(n21095), .Z(n21098) );
  XOR U20841 ( .A(\knn_comb_/min_val_out[0][17] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .Z(n21095) );
  XOR U20842 ( .A(n107), .B(n21099), .Z(o[16]) );
  AND U20843 ( .A(n122), .B(n21100), .Z(n107) );
  XOR U20844 ( .A(n108), .B(n21099), .Z(n21100) );
  XOR U20845 ( .A(n21101), .B(n21102), .Z(n21099) );
  AND U20846 ( .A(n142), .B(n21103), .Z(n21102) );
  XOR U20847 ( .A(n21104), .B(n35), .Z(n108) );
  AND U20848 ( .A(n125), .B(n21105), .Z(n35) );
  XOR U20849 ( .A(n36), .B(n21104), .Z(n21105) );
  XOR U20850 ( .A(n21106), .B(n21107), .Z(n36) );
  AND U20851 ( .A(n130), .B(n21108), .Z(n21107) );
  XOR U20852 ( .A(p_input[16]), .B(n21106), .Z(n21108) );
  XNOR U20853 ( .A(n21109), .B(n21110), .Z(n21106) );
  AND U20854 ( .A(n134), .B(n21111), .Z(n21110) );
  XOR U20855 ( .A(n21112), .B(n21113), .Z(n21104) );
  AND U20856 ( .A(n138), .B(n21103), .Z(n21113) );
  XNOR U20857 ( .A(n21114), .B(n21101), .Z(n21103) );
  XOR U20858 ( .A(n21115), .B(n21116), .Z(n21101) );
  AND U20859 ( .A(n162), .B(n21117), .Z(n21116) );
  IV U20860 ( .A(n21112), .Z(n21114) );
  XOR U20861 ( .A(n21118), .B(n21119), .Z(n21112) );
  AND U20862 ( .A(n146), .B(n21111), .Z(n21119) );
  XNOR U20863 ( .A(n21109), .B(n21118), .Z(n21111) );
  XNOR U20864 ( .A(n21120), .B(n21121), .Z(n21109) );
  AND U20865 ( .A(n150), .B(n21122), .Z(n21121) );
  XOR U20866 ( .A(p_input[48]), .B(n21120), .Z(n21122) );
  XNOR U20867 ( .A(n21123), .B(n21124), .Z(n21120) );
  AND U20868 ( .A(n154), .B(n21125), .Z(n21124) );
  XOR U20869 ( .A(n21126), .B(n21127), .Z(n21118) );
  AND U20870 ( .A(n158), .B(n21117), .Z(n21127) );
  XNOR U20871 ( .A(n21128), .B(n21115), .Z(n21117) );
  XOR U20872 ( .A(n21129), .B(n21130), .Z(n21115) );
  AND U20873 ( .A(n181), .B(n21131), .Z(n21130) );
  IV U20874 ( .A(n21126), .Z(n21128) );
  XOR U20875 ( .A(n21132), .B(n21133), .Z(n21126) );
  AND U20876 ( .A(n165), .B(n21125), .Z(n21133) );
  XNOR U20877 ( .A(n21123), .B(n21132), .Z(n21125) );
  XNOR U20878 ( .A(n21134), .B(n21135), .Z(n21123) );
  AND U20879 ( .A(n169), .B(n21136), .Z(n21135) );
  XOR U20880 ( .A(p_input[80]), .B(n21134), .Z(n21136) );
  XNOR U20881 ( .A(n21137), .B(n21138), .Z(n21134) );
  AND U20882 ( .A(n173), .B(n21139), .Z(n21138) );
  XOR U20883 ( .A(n21140), .B(n21141), .Z(n21132) );
  AND U20884 ( .A(n177), .B(n21131), .Z(n21141) );
  XNOR U20885 ( .A(n21142), .B(n21129), .Z(n21131) );
  XOR U20886 ( .A(n21143), .B(n21144), .Z(n21129) );
  AND U20887 ( .A(n200), .B(n21145), .Z(n21144) );
  IV U20888 ( .A(n21140), .Z(n21142) );
  XOR U20889 ( .A(n21146), .B(n21147), .Z(n21140) );
  AND U20890 ( .A(n184), .B(n21139), .Z(n21147) );
  XNOR U20891 ( .A(n21137), .B(n21146), .Z(n21139) );
  XNOR U20892 ( .A(n21148), .B(n21149), .Z(n21137) );
  AND U20893 ( .A(n188), .B(n21150), .Z(n21149) );
  XOR U20894 ( .A(p_input[112]), .B(n21148), .Z(n21150) );
  XNOR U20895 ( .A(n21151), .B(n21152), .Z(n21148) );
  AND U20896 ( .A(n192), .B(n21153), .Z(n21152) );
  XOR U20897 ( .A(n21154), .B(n21155), .Z(n21146) );
  AND U20898 ( .A(n196), .B(n21145), .Z(n21155) );
  XNOR U20899 ( .A(n21156), .B(n21143), .Z(n21145) );
  XOR U20900 ( .A(n21157), .B(n21158), .Z(n21143) );
  AND U20901 ( .A(n219), .B(n21159), .Z(n21158) );
  IV U20902 ( .A(n21154), .Z(n21156) );
  XOR U20903 ( .A(n21160), .B(n21161), .Z(n21154) );
  AND U20904 ( .A(n203), .B(n21153), .Z(n21161) );
  XNOR U20905 ( .A(n21151), .B(n21160), .Z(n21153) );
  XNOR U20906 ( .A(n21162), .B(n21163), .Z(n21151) );
  AND U20907 ( .A(n207), .B(n21164), .Z(n21163) );
  XOR U20908 ( .A(p_input[144]), .B(n21162), .Z(n21164) );
  XNOR U20909 ( .A(n21165), .B(n21166), .Z(n21162) );
  AND U20910 ( .A(n211), .B(n21167), .Z(n21166) );
  XOR U20911 ( .A(n21168), .B(n21169), .Z(n21160) );
  AND U20912 ( .A(n215), .B(n21159), .Z(n21169) );
  XNOR U20913 ( .A(n21170), .B(n21157), .Z(n21159) );
  XOR U20914 ( .A(n21171), .B(n21172), .Z(n21157) );
  AND U20915 ( .A(n238), .B(n21173), .Z(n21172) );
  IV U20916 ( .A(n21168), .Z(n21170) );
  XOR U20917 ( .A(n21174), .B(n21175), .Z(n21168) );
  AND U20918 ( .A(n222), .B(n21167), .Z(n21175) );
  XNOR U20919 ( .A(n21165), .B(n21174), .Z(n21167) );
  XNOR U20920 ( .A(n21176), .B(n21177), .Z(n21165) );
  AND U20921 ( .A(n226), .B(n21178), .Z(n21177) );
  XOR U20922 ( .A(p_input[176]), .B(n21176), .Z(n21178) );
  XNOR U20923 ( .A(n21179), .B(n21180), .Z(n21176) );
  AND U20924 ( .A(n230), .B(n21181), .Z(n21180) );
  XOR U20925 ( .A(n21182), .B(n21183), .Z(n21174) );
  AND U20926 ( .A(n234), .B(n21173), .Z(n21183) );
  XNOR U20927 ( .A(n21184), .B(n21171), .Z(n21173) );
  XOR U20928 ( .A(n21185), .B(n21186), .Z(n21171) );
  AND U20929 ( .A(n257), .B(n21187), .Z(n21186) );
  IV U20930 ( .A(n21182), .Z(n21184) );
  XOR U20931 ( .A(n21188), .B(n21189), .Z(n21182) );
  AND U20932 ( .A(n241), .B(n21181), .Z(n21189) );
  XNOR U20933 ( .A(n21179), .B(n21188), .Z(n21181) );
  XNOR U20934 ( .A(n21190), .B(n21191), .Z(n21179) );
  AND U20935 ( .A(n245), .B(n21192), .Z(n21191) );
  XOR U20936 ( .A(p_input[208]), .B(n21190), .Z(n21192) );
  XNOR U20937 ( .A(n21193), .B(n21194), .Z(n21190) );
  AND U20938 ( .A(n249), .B(n21195), .Z(n21194) );
  XOR U20939 ( .A(n21196), .B(n21197), .Z(n21188) );
  AND U20940 ( .A(n253), .B(n21187), .Z(n21197) );
  XNOR U20941 ( .A(n21198), .B(n21185), .Z(n21187) );
  XOR U20942 ( .A(n21199), .B(n21200), .Z(n21185) );
  AND U20943 ( .A(n276), .B(n21201), .Z(n21200) );
  IV U20944 ( .A(n21196), .Z(n21198) );
  XOR U20945 ( .A(n21202), .B(n21203), .Z(n21196) );
  AND U20946 ( .A(n260), .B(n21195), .Z(n21203) );
  XNOR U20947 ( .A(n21193), .B(n21202), .Z(n21195) );
  XNOR U20948 ( .A(n21204), .B(n21205), .Z(n21193) );
  AND U20949 ( .A(n264), .B(n21206), .Z(n21205) );
  XOR U20950 ( .A(p_input[240]), .B(n21204), .Z(n21206) );
  XNOR U20951 ( .A(n21207), .B(n21208), .Z(n21204) );
  AND U20952 ( .A(n268), .B(n21209), .Z(n21208) );
  XOR U20953 ( .A(n21210), .B(n21211), .Z(n21202) );
  AND U20954 ( .A(n272), .B(n21201), .Z(n21211) );
  XNOR U20955 ( .A(n21212), .B(n21199), .Z(n21201) );
  XOR U20956 ( .A(n21213), .B(n21214), .Z(n21199) );
  AND U20957 ( .A(n295), .B(n21215), .Z(n21214) );
  IV U20958 ( .A(n21210), .Z(n21212) );
  XOR U20959 ( .A(n21216), .B(n21217), .Z(n21210) );
  AND U20960 ( .A(n279), .B(n21209), .Z(n21217) );
  XNOR U20961 ( .A(n21207), .B(n21216), .Z(n21209) );
  XNOR U20962 ( .A(n21218), .B(n21219), .Z(n21207) );
  AND U20963 ( .A(n283), .B(n21220), .Z(n21219) );
  XOR U20964 ( .A(p_input[272]), .B(n21218), .Z(n21220) );
  XNOR U20965 ( .A(n21221), .B(n21222), .Z(n21218) );
  AND U20966 ( .A(n287), .B(n21223), .Z(n21222) );
  XOR U20967 ( .A(n21224), .B(n21225), .Z(n21216) );
  AND U20968 ( .A(n291), .B(n21215), .Z(n21225) );
  XNOR U20969 ( .A(n21226), .B(n21213), .Z(n21215) );
  XOR U20970 ( .A(n21227), .B(n21228), .Z(n21213) );
  AND U20971 ( .A(n314), .B(n21229), .Z(n21228) );
  IV U20972 ( .A(n21224), .Z(n21226) );
  XOR U20973 ( .A(n21230), .B(n21231), .Z(n21224) );
  AND U20974 ( .A(n298), .B(n21223), .Z(n21231) );
  XNOR U20975 ( .A(n21221), .B(n21230), .Z(n21223) );
  XNOR U20976 ( .A(n21232), .B(n21233), .Z(n21221) );
  AND U20977 ( .A(n302), .B(n21234), .Z(n21233) );
  XOR U20978 ( .A(p_input[304]), .B(n21232), .Z(n21234) );
  XNOR U20979 ( .A(n21235), .B(n21236), .Z(n21232) );
  AND U20980 ( .A(n306), .B(n21237), .Z(n21236) );
  XOR U20981 ( .A(n21238), .B(n21239), .Z(n21230) );
  AND U20982 ( .A(n310), .B(n21229), .Z(n21239) );
  XNOR U20983 ( .A(n21240), .B(n21227), .Z(n21229) );
  XOR U20984 ( .A(n21241), .B(n21242), .Z(n21227) );
  AND U20985 ( .A(n333), .B(n21243), .Z(n21242) );
  IV U20986 ( .A(n21238), .Z(n21240) );
  XOR U20987 ( .A(n21244), .B(n21245), .Z(n21238) );
  AND U20988 ( .A(n317), .B(n21237), .Z(n21245) );
  XNOR U20989 ( .A(n21235), .B(n21244), .Z(n21237) );
  XNOR U20990 ( .A(n21246), .B(n21247), .Z(n21235) );
  AND U20991 ( .A(n321), .B(n21248), .Z(n21247) );
  XOR U20992 ( .A(p_input[336]), .B(n21246), .Z(n21248) );
  XNOR U20993 ( .A(n21249), .B(n21250), .Z(n21246) );
  AND U20994 ( .A(n325), .B(n21251), .Z(n21250) );
  XOR U20995 ( .A(n21252), .B(n21253), .Z(n21244) );
  AND U20996 ( .A(n329), .B(n21243), .Z(n21253) );
  XNOR U20997 ( .A(n21254), .B(n21241), .Z(n21243) );
  XOR U20998 ( .A(n21255), .B(n21256), .Z(n21241) );
  AND U20999 ( .A(n352), .B(n21257), .Z(n21256) );
  IV U21000 ( .A(n21252), .Z(n21254) );
  XOR U21001 ( .A(n21258), .B(n21259), .Z(n21252) );
  AND U21002 ( .A(n336), .B(n21251), .Z(n21259) );
  XNOR U21003 ( .A(n21249), .B(n21258), .Z(n21251) );
  XNOR U21004 ( .A(n21260), .B(n21261), .Z(n21249) );
  AND U21005 ( .A(n340), .B(n21262), .Z(n21261) );
  XOR U21006 ( .A(p_input[368]), .B(n21260), .Z(n21262) );
  XNOR U21007 ( .A(n21263), .B(n21264), .Z(n21260) );
  AND U21008 ( .A(n344), .B(n21265), .Z(n21264) );
  XOR U21009 ( .A(n21266), .B(n21267), .Z(n21258) );
  AND U21010 ( .A(n348), .B(n21257), .Z(n21267) );
  XNOR U21011 ( .A(n21268), .B(n21255), .Z(n21257) );
  XOR U21012 ( .A(n21269), .B(n21270), .Z(n21255) );
  AND U21013 ( .A(n371), .B(n21271), .Z(n21270) );
  IV U21014 ( .A(n21266), .Z(n21268) );
  XOR U21015 ( .A(n21272), .B(n21273), .Z(n21266) );
  AND U21016 ( .A(n355), .B(n21265), .Z(n21273) );
  XNOR U21017 ( .A(n21263), .B(n21272), .Z(n21265) );
  XNOR U21018 ( .A(n21274), .B(n21275), .Z(n21263) );
  AND U21019 ( .A(n359), .B(n21276), .Z(n21275) );
  XOR U21020 ( .A(p_input[400]), .B(n21274), .Z(n21276) );
  XNOR U21021 ( .A(n21277), .B(n21278), .Z(n21274) );
  AND U21022 ( .A(n363), .B(n21279), .Z(n21278) );
  XOR U21023 ( .A(n21280), .B(n21281), .Z(n21272) );
  AND U21024 ( .A(n367), .B(n21271), .Z(n21281) );
  XNOR U21025 ( .A(n21282), .B(n21269), .Z(n21271) );
  XOR U21026 ( .A(n21283), .B(n21284), .Z(n21269) );
  AND U21027 ( .A(n390), .B(n21285), .Z(n21284) );
  IV U21028 ( .A(n21280), .Z(n21282) );
  XOR U21029 ( .A(n21286), .B(n21287), .Z(n21280) );
  AND U21030 ( .A(n374), .B(n21279), .Z(n21287) );
  XNOR U21031 ( .A(n21277), .B(n21286), .Z(n21279) );
  XNOR U21032 ( .A(n21288), .B(n21289), .Z(n21277) );
  AND U21033 ( .A(n378), .B(n21290), .Z(n21289) );
  XOR U21034 ( .A(p_input[432]), .B(n21288), .Z(n21290) );
  XNOR U21035 ( .A(n21291), .B(n21292), .Z(n21288) );
  AND U21036 ( .A(n382), .B(n21293), .Z(n21292) );
  XOR U21037 ( .A(n21294), .B(n21295), .Z(n21286) );
  AND U21038 ( .A(n386), .B(n21285), .Z(n21295) );
  XNOR U21039 ( .A(n21296), .B(n21283), .Z(n21285) );
  XOR U21040 ( .A(n21297), .B(n21298), .Z(n21283) );
  AND U21041 ( .A(n409), .B(n21299), .Z(n21298) );
  IV U21042 ( .A(n21294), .Z(n21296) );
  XOR U21043 ( .A(n21300), .B(n21301), .Z(n21294) );
  AND U21044 ( .A(n393), .B(n21293), .Z(n21301) );
  XNOR U21045 ( .A(n21291), .B(n21300), .Z(n21293) );
  XNOR U21046 ( .A(n21302), .B(n21303), .Z(n21291) );
  AND U21047 ( .A(n397), .B(n21304), .Z(n21303) );
  XOR U21048 ( .A(p_input[464]), .B(n21302), .Z(n21304) );
  XNOR U21049 ( .A(n21305), .B(n21306), .Z(n21302) );
  AND U21050 ( .A(n401), .B(n21307), .Z(n21306) );
  XOR U21051 ( .A(n21308), .B(n21309), .Z(n21300) );
  AND U21052 ( .A(n405), .B(n21299), .Z(n21309) );
  XNOR U21053 ( .A(n21310), .B(n21297), .Z(n21299) );
  XOR U21054 ( .A(n21311), .B(n21312), .Z(n21297) );
  AND U21055 ( .A(n428), .B(n21313), .Z(n21312) );
  IV U21056 ( .A(n21308), .Z(n21310) );
  XOR U21057 ( .A(n21314), .B(n21315), .Z(n21308) );
  AND U21058 ( .A(n412), .B(n21307), .Z(n21315) );
  XNOR U21059 ( .A(n21305), .B(n21314), .Z(n21307) );
  XNOR U21060 ( .A(n21316), .B(n21317), .Z(n21305) );
  AND U21061 ( .A(n416), .B(n21318), .Z(n21317) );
  XOR U21062 ( .A(p_input[496]), .B(n21316), .Z(n21318) );
  XNOR U21063 ( .A(n21319), .B(n21320), .Z(n21316) );
  AND U21064 ( .A(n420), .B(n21321), .Z(n21320) );
  XOR U21065 ( .A(n21322), .B(n21323), .Z(n21314) );
  AND U21066 ( .A(n424), .B(n21313), .Z(n21323) );
  XNOR U21067 ( .A(n21324), .B(n21311), .Z(n21313) );
  XOR U21068 ( .A(n21325), .B(n21326), .Z(n21311) );
  AND U21069 ( .A(n447), .B(n21327), .Z(n21326) );
  IV U21070 ( .A(n21322), .Z(n21324) );
  XOR U21071 ( .A(n21328), .B(n21329), .Z(n21322) );
  AND U21072 ( .A(n431), .B(n21321), .Z(n21329) );
  XNOR U21073 ( .A(n21319), .B(n21328), .Z(n21321) );
  XNOR U21074 ( .A(n21330), .B(n21331), .Z(n21319) );
  AND U21075 ( .A(n435), .B(n21332), .Z(n21331) );
  XOR U21076 ( .A(p_input[528]), .B(n21330), .Z(n21332) );
  XNOR U21077 ( .A(n21333), .B(n21334), .Z(n21330) );
  AND U21078 ( .A(n439), .B(n21335), .Z(n21334) );
  XOR U21079 ( .A(n21336), .B(n21337), .Z(n21328) );
  AND U21080 ( .A(n443), .B(n21327), .Z(n21337) );
  XNOR U21081 ( .A(n21338), .B(n21325), .Z(n21327) );
  XOR U21082 ( .A(n21339), .B(n21340), .Z(n21325) );
  AND U21083 ( .A(n466), .B(n21341), .Z(n21340) );
  IV U21084 ( .A(n21336), .Z(n21338) );
  XOR U21085 ( .A(n21342), .B(n21343), .Z(n21336) );
  AND U21086 ( .A(n450), .B(n21335), .Z(n21343) );
  XNOR U21087 ( .A(n21333), .B(n21342), .Z(n21335) );
  XNOR U21088 ( .A(n21344), .B(n21345), .Z(n21333) );
  AND U21089 ( .A(n454), .B(n21346), .Z(n21345) );
  XOR U21090 ( .A(p_input[560]), .B(n21344), .Z(n21346) );
  XNOR U21091 ( .A(n21347), .B(n21348), .Z(n21344) );
  AND U21092 ( .A(n458), .B(n21349), .Z(n21348) );
  XOR U21093 ( .A(n21350), .B(n21351), .Z(n21342) );
  AND U21094 ( .A(n462), .B(n21341), .Z(n21351) );
  XNOR U21095 ( .A(n21352), .B(n21339), .Z(n21341) );
  XOR U21096 ( .A(n21353), .B(n21354), .Z(n21339) );
  AND U21097 ( .A(n485), .B(n21355), .Z(n21354) );
  IV U21098 ( .A(n21350), .Z(n21352) );
  XOR U21099 ( .A(n21356), .B(n21357), .Z(n21350) );
  AND U21100 ( .A(n469), .B(n21349), .Z(n21357) );
  XNOR U21101 ( .A(n21347), .B(n21356), .Z(n21349) );
  XNOR U21102 ( .A(n21358), .B(n21359), .Z(n21347) );
  AND U21103 ( .A(n473), .B(n21360), .Z(n21359) );
  XOR U21104 ( .A(p_input[592]), .B(n21358), .Z(n21360) );
  XNOR U21105 ( .A(n21361), .B(n21362), .Z(n21358) );
  AND U21106 ( .A(n477), .B(n21363), .Z(n21362) );
  XOR U21107 ( .A(n21364), .B(n21365), .Z(n21356) );
  AND U21108 ( .A(n481), .B(n21355), .Z(n21365) );
  XNOR U21109 ( .A(n21366), .B(n21353), .Z(n21355) );
  XOR U21110 ( .A(n21367), .B(n21368), .Z(n21353) );
  AND U21111 ( .A(n504), .B(n21369), .Z(n21368) );
  IV U21112 ( .A(n21364), .Z(n21366) );
  XOR U21113 ( .A(n21370), .B(n21371), .Z(n21364) );
  AND U21114 ( .A(n488), .B(n21363), .Z(n21371) );
  XNOR U21115 ( .A(n21361), .B(n21370), .Z(n21363) );
  XNOR U21116 ( .A(n21372), .B(n21373), .Z(n21361) );
  AND U21117 ( .A(n492), .B(n21374), .Z(n21373) );
  XOR U21118 ( .A(p_input[624]), .B(n21372), .Z(n21374) );
  XNOR U21119 ( .A(n21375), .B(n21376), .Z(n21372) );
  AND U21120 ( .A(n496), .B(n21377), .Z(n21376) );
  XOR U21121 ( .A(n21378), .B(n21379), .Z(n21370) );
  AND U21122 ( .A(n500), .B(n21369), .Z(n21379) );
  XNOR U21123 ( .A(n21380), .B(n21367), .Z(n21369) );
  XOR U21124 ( .A(n21381), .B(n21382), .Z(n21367) );
  AND U21125 ( .A(n523), .B(n21383), .Z(n21382) );
  IV U21126 ( .A(n21378), .Z(n21380) );
  XOR U21127 ( .A(n21384), .B(n21385), .Z(n21378) );
  AND U21128 ( .A(n507), .B(n21377), .Z(n21385) );
  XNOR U21129 ( .A(n21375), .B(n21384), .Z(n21377) );
  XNOR U21130 ( .A(n21386), .B(n21387), .Z(n21375) );
  AND U21131 ( .A(n511), .B(n21388), .Z(n21387) );
  XOR U21132 ( .A(p_input[656]), .B(n21386), .Z(n21388) );
  XNOR U21133 ( .A(n21389), .B(n21390), .Z(n21386) );
  AND U21134 ( .A(n515), .B(n21391), .Z(n21390) );
  XOR U21135 ( .A(n21392), .B(n21393), .Z(n21384) );
  AND U21136 ( .A(n519), .B(n21383), .Z(n21393) );
  XNOR U21137 ( .A(n21394), .B(n21381), .Z(n21383) );
  XOR U21138 ( .A(n21395), .B(n21396), .Z(n21381) );
  AND U21139 ( .A(n542), .B(n21397), .Z(n21396) );
  IV U21140 ( .A(n21392), .Z(n21394) );
  XOR U21141 ( .A(n21398), .B(n21399), .Z(n21392) );
  AND U21142 ( .A(n526), .B(n21391), .Z(n21399) );
  XNOR U21143 ( .A(n21389), .B(n21398), .Z(n21391) );
  XNOR U21144 ( .A(n21400), .B(n21401), .Z(n21389) );
  AND U21145 ( .A(n530), .B(n21402), .Z(n21401) );
  XOR U21146 ( .A(p_input[688]), .B(n21400), .Z(n21402) );
  XNOR U21147 ( .A(n21403), .B(n21404), .Z(n21400) );
  AND U21148 ( .A(n534), .B(n21405), .Z(n21404) );
  XOR U21149 ( .A(n21406), .B(n21407), .Z(n21398) );
  AND U21150 ( .A(n538), .B(n21397), .Z(n21407) );
  XNOR U21151 ( .A(n21408), .B(n21395), .Z(n21397) );
  XOR U21152 ( .A(n21409), .B(n21410), .Z(n21395) );
  AND U21153 ( .A(n561), .B(n21411), .Z(n21410) );
  IV U21154 ( .A(n21406), .Z(n21408) );
  XOR U21155 ( .A(n21412), .B(n21413), .Z(n21406) );
  AND U21156 ( .A(n545), .B(n21405), .Z(n21413) );
  XNOR U21157 ( .A(n21403), .B(n21412), .Z(n21405) );
  XNOR U21158 ( .A(n21414), .B(n21415), .Z(n21403) );
  AND U21159 ( .A(n549), .B(n21416), .Z(n21415) );
  XOR U21160 ( .A(p_input[720]), .B(n21414), .Z(n21416) );
  XNOR U21161 ( .A(n21417), .B(n21418), .Z(n21414) );
  AND U21162 ( .A(n553), .B(n21419), .Z(n21418) );
  XOR U21163 ( .A(n21420), .B(n21421), .Z(n21412) );
  AND U21164 ( .A(n557), .B(n21411), .Z(n21421) );
  XNOR U21165 ( .A(n21422), .B(n21409), .Z(n21411) );
  XOR U21166 ( .A(n21423), .B(n21424), .Z(n21409) );
  AND U21167 ( .A(n580), .B(n21425), .Z(n21424) );
  IV U21168 ( .A(n21420), .Z(n21422) );
  XOR U21169 ( .A(n21426), .B(n21427), .Z(n21420) );
  AND U21170 ( .A(n564), .B(n21419), .Z(n21427) );
  XNOR U21171 ( .A(n21417), .B(n21426), .Z(n21419) );
  XNOR U21172 ( .A(n21428), .B(n21429), .Z(n21417) );
  AND U21173 ( .A(n568), .B(n21430), .Z(n21429) );
  XOR U21174 ( .A(p_input[752]), .B(n21428), .Z(n21430) );
  XNOR U21175 ( .A(n21431), .B(n21432), .Z(n21428) );
  AND U21176 ( .A(n572), .B(n21433), .Z(n21432) );
  XOR U21177 ( .A(n21434), .B(n21435), .Z(n21426) );
  AND U21178 ( .A(n576), .B(n21425), .Z(n21435) );
  XNOR U21179 ( .A(n21436), .B(n21423), .Z(n21425) );
  XOR U21180 ( .A(n21437), .B(n21438), .Z(n21423) );
  AND U21181 ( .A(n599), .B(n21439), .Z(n21438) );
  IV U21182 ( .A(n21434), .Z(n21436) );
  XOR U21183 ( .A(n21440), .B(n21441), .Z(n21434) );
  AND U21184 ( .A(n583), .B(n21433), .Z(n21441) );
  XNOR U21185 ( .A(n21431), .B(n21440), .Z(n21433) );
  XNOR U21186 ( .A(n21442), .B(n21443), .Z(n21431) );
  AND U21187 ( .A(n587), .B(n21444), .Z(n21443) );
  XOR U21188 ( .A(p_input[784]), .B(n21442), .Z(n21444) );
  XNOR U21189 ( .A(n21445), .B(n21446), .Z(n21442) );
  AND U21190 ( .A(n591), .B(n21447), .Z(n21446) );
  XOR U21191 ( .A(n21448), .B(n21449), .Z(n21440) );
  AND U21192 ( .A(n595), .B(n21439), .Z(n21449) );
  XNOR U21193 ( .A(n21450), .B(n21437), .Z(n21439) );
  XOR U21194 ( .A(n21451), .B(n21452), .Z(n21437) );
  AND U21195 ( .A(n618), .B(n21453), .Z(n21452) );
  IV U21196 ( .A(n21448), .Z(n21450) );
  XOR U21197 ( .A(n21454), .B(n21455), .Z(n21448) );
  AND U21198 ( .A(n602), .B(n21447), .Z(n21455) );
  XNOR U21199 ( .A(n21445), .B(n21454), .Z(n21447) );
  XNOR U21200 ( .A(n21456), .B(n21457), .Z(n21445) );
  AND U21201 ( .A(n606), .B(n21458), .Z(n21457) );
  XOR U21202 ( .A(p_input[816]), .B(n21456), .Z(n21458) );
  XNOR U21203 ( .A(n21459), .B(n21460), .Z(n21456) );
  AND U21204 ( .A(n610), .B(n21461), .Z(n21460) );
  XOR U21205 ( .A(n21462), .B(n21463), .Z(n21454) );
  AND U21206 ( .A(n614), .B(n21453), .Z(n21463) );
  XNOR U21207 ( .A(n21464), .B(n21451), .Z(n21453) );
  XOR U21208 ( .A(n21465), .B(n21466), .Z(n21451) );
  AND U21209 ( .A(n637), .B(n21467), .Z(n21466) );
  IV U21210 ( .A(n21462), .Z(n21464) );
  XOR U21211 ( .A(n21468), .B(n21469), .Z(n21462) );
  AND U21212 ( .A(n621), .B(n21461), .Z(n21469) );
  XNOR U21213 ( .A(n21459), .B(n21468), .Z(n21461) );
  XNOR U21214 ( .A(n21470), .B(n21471), .Z(n21459) );
  AND U21215 ( .A(n625), .B(n21472), .Z(n21471) );
  XOR U21216 ( .A(p_input[848]), .B(n21470), .Z(n21472) );
  XNOR U21217 ( .A(n21473), .B(n21474), .Z(n21470) );
  AND U21218 ( .A(n629), .B(n21475), .Z(n21474) );
  XOR U21219 ( .A(n21476), .B(n21477), .Z(n21468) );
  AND U21220 ( .A(n633), .B(n21467), .Z(n21477) );
  XNOR U21221 ( .A(n21478), .B(n21465), .Z(n21467) );
  XOR U21222 ( .A(n21479), .B(n21480), .Z(n21465) );
  AND U21223 ( .A(n656), .B(n21481), .Z(n21480) );
  IV U21224 ( .A(n21476), .Z(n21478) );
  XOR U21225 ( .A(n21482), .B(n21483), .Z(n21476) );
  AND U21226 ( .A(n640), .B(n21475), .Z(n21483) );
  XNOR U21227 ( .A(n21473), .B(n21482), .Z(n21475) );
  XNOR U21228 ( .A(n21484), .B(n21485), .Z(n21473) );
  AND U21229 ( .A(n644), .B(n21486), .Z(n21485) );
  XOR U21230 ( .A(p_input[880]), .B(n21484), .Z(n21486) );
  XNOR U21231 ( .A(n21487), .B(n21488), .Z(n21484) );
  AND U21232 ( .A(n648), .B(n21489), .Z(n21488) );
  XOR U21233 ( .A(n21490), .B(n21491), .Z(n21482) );
  AND U21234 ( .A(n652), .B(n21481), .Z(n21491) );
  XNOR U21235 ( .A(n21492), .B(n21479), .Z(n21481) );
  XOR U21236 ( .A(n21493), .B(n21494), .Z(n21479) );
  AND U21237 ( .A(n675), .B(n21495), .Z(n21494) );
  IV U21238 ( .A(n21490), .Z(n21492) );
  XOR U21239 ( .A(n21496), .B(n21497), .Z(n21490) );
  AND U21240 ( .A(n659), .B(n21489), .Z(n21497) );
  XNOR U21241 ( .A(n21487), .B(n21496), .Z(n21489) );
  XNOR U21242 ( .A(n21498), .B(n21499), .Z(n21487) );
  AND U21243 ( .A(n663), .B(n21500), .Z(n21499) );
  XOR U21244 ( .A(p_input[912]), .B(n21498), .Z(n21500) );
  XNOR U21245 ( .A(n21501), .B(n21502), .Z(n21498) );
  AND U21246 ( .A(n667), .B(n21503), .Z(n21502) );
  XOR U21247 ( .A(n21504), .B(n21505), .Z(n21496) );
  AND U21248 ( .A(n671), .B(n21495), .Z(n21505) );
  XNOR U21249 ( .A(n21506), .B(n21493), .Z(n21495) );
  XOR U21250 ( .A(n21507), .B(n21508), .Z(n21493) );
  AND U21251 ( .A(n694), .B(n21509), .Z(n21508) );
  IV U21252 ( .A(n21504), .Z(n21506) );
  XOR U21253 ( .A(n21510), .B(n21511), .Z(n21504) );
  AND U21254 ( .A(n678), .B(n21503), .Z(n21511) );
  XNOR U21255 ( .A(n21501), .B(n21510), .Z(n21503) );
  XNOR U21256 ( .A(n21512), .B(n21513), .Z(n21501) );
  AND U21257 ( .A(n682), .B(n21514), .Z(n21513) );
  XOR U21258 ( .A(p_input[944]), .B(n21512), .Z(n21514) );
  XNOR U21259 ( .A(n21515), .B(n21516), .Z(n21512) );
  AND U21260 ( .A(n686), .B(n21517), .Z(n21516) );
  XOR U21261 ( .A(n21518), .B(n21519), .Z(n21510) );
  AND U21262 ( .A(n690), .B(n21509), .Z(n21519) );
  XNOR U21263 ( .A(n21520), .B(n21507), .Z(n21509) );
  XOR U21264 ( .A(n21521), .B(n21522), .Z(n21507) );
  AND U21265 ( .A(n713), .B(n21523), .Z(n21522) );
  IV U21266 ( .A(n21518), .Z(n21520) );
  XOR U21267 ( .A(n21524), .B(n21525), .Z(n21518) );
  AND U21268 ( .A(n697), .B(n21517), .Z(n21525) );
  XNOR U21269 ( .A(n21515), .B(n21524), .Z(n21517) );
  XNOR U21270 ( .A(n21526), .B(n21527), .Z(n21515) );
  AND U21271 ( .A(n701), .B(n21528), .Z(n21527) );
  XOR U21272 ( .A(p_input[976]), .B(n21526), .Z(n21528) );
  XNOR U21273 ( .A(n21529), .B(n21530), .Z(n21526) );
  AND U21274 ( .A(n705), .B(n21531), .Z(n21530) );
  XOR U21275 ( .A(n21532), .B(n21533), .Z(n21524) );
  AND U21276 ( .A(n709), .B(n21523), .Z(n21533) );
  XNOR U21277 ( .A(n21534), .B(n21521), .Z(n21523) );
  XOR U21278 ( .A(n21535), .B(n21536), .Z(n21521) );
  AND U21279 ( .A(n732), .B(n21537), .Z(n21536) );
  IV U21280 ( .A(n21532), .Z(n21534) );
  XOR U21281 ( .A(n21538), .B(n21539), .Z(n21532) );
  AND U21282 ( .A(n716), .B(n21531), .Z(n21539) );
  XNOR U21283 ( .A(n21529), .B(n21538), .Z(n21531) );
  XNOR U21284 ( .A(n21540), .B(n21541), .Z(n21529) );
  AND U21285 ( .A(n720), .B(n21542), .Z(n21541) );
  XOR U21286 ( .A(p_input[1008]), .B(n21540), .Z(n21542) );
  XNOR U21287 ( .A(n21543), .B(n21544), .Z(n21540) );
  AND U21288 ( .A(n724), .B(n21545), .Z(n21544) );
  XOR U21289 ( .A(n21546), .B(n21547), .Z(n21538) );
  AND U21290 ( .A(n728), .B(n21537), .Z(n21547) );
  XNOR U21291 ( .A(n21548), .B(n21535), .Z(n21537) );
  XOR U21292 ( .A(n21549), .B(n21550), .Z(n21535) );
  AND U21293 ( .A(n751), .B(n21551), .Z(n21550) );
  IV U21294 ( .A(n21546), .Z(n21548) );
  XOR U21295 ( .A(n21552), .B(n21553), .Z(n21546) );
  AND U21296 ( .A(n735), .B(n21545), .Z(n21553) );
  XNOR U21297 ( .A(n21543), .B(n21552), .Z(n21545) );
  XNOR U21298 ( .A(n21554), .B(n21555), .Z(n21543) );
  AND U21299 ( .A(n739), .B(n21556), .Z(n21555) );
  XOR U21300 ( .A(p_input[1040]), .B(n21554), .Z(n21556) );
  XNOR U21301 ( .A(n21557), .B(n21558), .Z(n21554) );
  AND U21302 ( .A(n743), .B(n21559), .Z(n21558) );
  XOR U21303 ( .A(n21560), .B(n21561), .Z(n21552) );
  AND U21304 ( .A(n747), .B(n21551), .Z(n21561) );
  XNOR U21305 ( .A(n21562), .B(n21549), .Z(n21551) );
  XOR U21306 ( .A(n21563), .B(n21564), .Z(n21549) );
  AND U21307 ( .A(n770), .B(n21565), .Z(n21564) );
  IV U21308 ( .A(n21560), .Z(n21562) );
  XOR U21309 ( .A(n21566), .B(n21567), .Z(n21560) );
  AND U21310 ( .A(n754), .B(n21559), .Z(n21567) );
  XNOR U21311 ( .A(n21557), .B(n21566), .Z(n21559) );
  XNOR U21312 ( .A(n21568), .B(n21569), .Z(n21557) );
  AND U21313 ( .A(n758), .B(n21570), .Z(n21569) );
  XOR U21314 ( .A(p_input[1072]), .B(n21568), .Z(n21570) );
  XNOR U21315 ( .A(n21571), .B(n21572), .Z(n21568) );
  AND U21316 ( .A(n762), .B(n21573), .Z(n21572) );
  XOR U21317 ( .A(n21574), .B(n21575), .Z(n21566) );
  AND U21318 ( .A(n766), .B(n21565), .Z(n21575) );
  XNOR U21319 ( .A(n21576), .B(n21563), .Z(n21565) );
  XOR U21320 ( .A(n21577), .B(n21578), .Z(n21563) );
  AND U21321 ( .A(n789), .B(n21579), .Z(n21578) );
  IV U21322 ( .A(n21574), .Z(n21576) );
  XOR U21323 ( .A(n21580), .B(n21581), .Z(n21574) );
  AND U21324 ( .A(n773), .B(n21573), .Z(n21581) );
  XNOR U21325 ( .A(n21571), .B(n21580), .Z(n21573) );
  XNOR U21326 ( .A(n21582), .B(n21583), .Z(n21571) );
  AND U21327 ( .A(n777), .B(n21584), .Z(n21583) );
  XOR U21328 ( .A(p_input[1104]), .B(n21582), .Z(n21584) );
  XNOR U21329 ( .A(n21585), .B(n21586), .Z(n21582) );
  AND U21330 ( .A(n781), .B(n21587), .Z(n21586) );
  XOR U21331 ( .A(n21588), .B(n21589), .Z(n21580) );
  AND U21332 ( .A(n785), .B(n21579), .Z(n21589) );
  XNOR U21333 ( .A(n21590), .B(n21577), .Z(n21579) );
  XOR U21334 ( .A(n21591), .B(n21592), .Z(n21577) );
  AND U21335 ( .A(n808), .B(n21593), .Z(n21592) );
  IV U21336 ( .A(n21588), .Z(n21590) );
  XOR U21337 ( .A(n21594), .B(n21595), .Z(n21588) );
  AND U21338 ( .A(n792), .B(n21587), .Z(n21595) );
  XNOR U21339 ( .A(n21585), .B(n21594), .Z(n21587) );
  XNOR U21340 ( .A(n21596), .B(n21597), .Z(n21585) );
  AND U21341 ( .A(n796), .B(n21598), .Z(n21597) );
  XOR U21342 ( .A(p_input[1136]), .B(n21596), .Z(n21598) );
  XNOR U21343 ( .A(n21599), .B(n21600), .Z(n21596) );
  AND U21344 ( .A(n800), .B(n21601), .Z(n21600) );
  XOR U21345 ( .A(n21602), .B(n21603), .Z(n21594) );
  AND U21346 ( .A(n804), .B(n21593), .Z(n21603) );
  XNOR U21347 ( .A(n21604), .B(n21591), .Z(n21593) );
  XOR U21348 ( .A(n21605), .B(n21606), .Z(n21591) );
  AND U21349 ( .A(n827), .B(n21607), .Z(n21606) );
  IV U21350 ( .A(n21602), .Z(n21604) );
  XOR U21351 ( .A(n21608), .B(n21609), .Z(n21602) );
  AND U21352 ( .A(n811), .B(n21601), .Z(n21609) );
  XNOR U21353 ( .A(n21599), .B(n21608), .Z(n21601) );
  XNOR U21354 ( .A(n21610), .B(n21611), .Z(n21599) );
  AND U21355 ( .A(n815), .B(n21612), .Z(n21611) );
  XOR U21356 ( .A(p_input[1168]), .B(n21610), .Z(n21612) );
  XNOR U21357 ( .A(n21613), .B(n21614), .Z(n21610) );
  AND U21358 ( .A(n819), .B(n21615), .Z(n21614) );
  XOR U21359 ( .A(n21616), .B(n21617), .Z(n21608) );
  AND U21360 ( .A(n823), .B(n21607), .Z(n21617) );
  XNOR U21361 ( .A(n21618), .B(n21605), .Z(n21607) );
  XOR U21362 ( .A(n21619), .B(n21620), .Z(n21605) );
  AND U21363 ( .A(n846), .B(n21621), .Z(n21620) );
  IV U21364 ( .A(n21616), .Z(n21618) );
  XOR U21365 ( .A(n21622), .B(n21623), .Z(n21616) );
  AND U21366 ( .A(n830), .B(n21615), .Z(n21623) );
  XNOR U21367 ( .A(n21613), .B(n21622), .Z(n21615) );
  XNOR U21368 ( .A(n21624), .B(n21625), .Z(n21613) );
  AND U21369 ( .A(n834), .B(n21626), .Z(n21625) );
  XOR U21370 ( .A(p_input[1200]), .B(n21624), .Z(n21626) );
  XNOR U21371 ( .A(n21627), .B(n21628), .Z(n21624) );
  AND U21372 ( .A(n838), .B(n21629), .Z(n21628) );
  XOR U21373 ( .A(n21630), .B(n21631), .Z(n21622) );
  AND U21374 ( .A(n842), .B(n21621), .Z(n21631) );
  XNOR U21375 ( .A(n21632), .B(n21619), .Z(n21621) );
  XOR U21376 ( .A(n21633), .B(n21634), .Z(n21619) );
  AND U21377 ( .A(n865), .B(n21635), .Z(n21634) );
  IV U21378 ( .A(n21630), .Z(n21632) );
  XOR U21379 ( .A(n21636), .B(n21637), .Z(n21630) );
  AND U21380 ( .A(n849), .B(n21629), .Z(n21637) );
  XNOR U21381 ( .A(n21627), .B(n21636), .Z(n21629) );
  XNOR U21382 ( .A(n21638), .B(n21639), .Z(n21627) );
  AND U21383 ( .A(n853), .B(n21640), .Z(n21639) );
  XOR U21384 ( .A(p_input[1232]), .B(n21638), .Z(n21640) );
  XNOR U21385 ( .A(n21641), .B(n21642), .Z(n21638) );
  AND U21386 ( .A(n857), .B(n21643), .Z(n21642) );
  XOR U21387 ( .A(n21644), .B(n21645), .Z(n21636) );
  AND U21388 ( .A(n861), .B(n21635), .Z(n21645) );
  XNOR U21389 ( .A(n21646), .B(n21633), .Z(n21635) );
  XOR U21390 ( .A(n21647), .B(n21648), .Z(n21633) );
  AND U21391 ( .A(n884), .B(n21649), .Z(n21648) );
  IV U21392 ( .A(n21644), .Z(n21646) );
  XOR U21393 ( .A(n21650), .B(n21651), .Z(n21644) );
  AND U21394 ( .A(n868), .B(n21643), .Z(n21651) );
  XNOR U21395 ( .A(n21641), .B(n21650), .Z(n21643) );
  XNOR U21396 ( .A(n21652), .B(n21653), .Z(n21641) );
  AND U21397 ( .A(n872), .B(n21654), .Z(n21653) );
  XOR U21398 ( .A(p_input[1264]), .B(n21652), .Z(n21654) );
  XNOR U21399 ( .A(n21655), .B(n21656), .Z(n21652) );
  AND U21400 ( .A(n876), .B(n21657), .Z(n21656) );
  XOR U21401 ( .A(n21658), .B(n21659), .Z(n21650) );
  AND U21402 ( .A(n880), .B(n21649), .Z(n21659) );
  XNOR U21403 ( .A(n21660), .B(n21647), .Z(n21649) );
  XOR U21404 ( .A(n21661), .B(n21662), .Z(n21647) );
  AND U21405 ( .A(n903), .B(n21663), .Z(n21662) );
  IV U21406 ( .A(n21658), .Z(n21660) );
  XOR U21407 ( .A(n21664), .B(n21665), .Z(n21658) );
  AND U21408 ( .A(n887), .B(n21657), .Z(n21665) );
  XNOR U21409 ( .A(n21655), .B(n21664), .Z(n21657) );
  XNOR U21410 ( .A(n21666), .B(n21667), .Z(n21655) );
  AND U21411 ( .A(n891), .B(n21668), .Z(n21667) );
  XOR U21412 ( .A(p_input[1296]), .B(n21666), .Z(n21668) );
  XNOR U21413 ( .A(n21669), .B(n21670), .Z(n21666) );
  AND U21414 ( .A(n895), .B(n21671), .Z(n21670) );
  XOR U21415 ( .A(n21672), .B(n21673), .Z(n21664) );
  AND U21416 ( .A(n899), .B(n21663), .Z(n21673) );
  XNOR U21417 ( .A(n21674), .B(n21661), .Z(n21663) );
  XOR U21418 ( .A(n21675), .B(n21676), .Z(n21661) );
  AND U21419 ( .A(n922), .B(n21677), .Z(n21676) );
  IV U21420 ( .A(n21672), .Z(n21674) );
  XOR U21421 ( .A(n21678), .B(n21679), .Z(n21672) );
  AND U21422 ( .A(n906), .B(n21671), .Z(n21679) );
  XNOR U21423 ( .A(n21669), .B(n21678), .Z(n21671) );
  XNOR U21424 ( .A(n21680), .B(n21681), .Z(n21669) );
  AND U21425 ( .A(n910), .B(n21682), .Z(n21681) );
  XOR U21426 ( .A(p_input[1328]), .B(n21680), .Z(n21682) );
  XNOR U21427 ( .A(n21683), .B(n21684), .Z(n21680) );
  AND U21428 ( .A(n914), .B(n21685), .Z(n21684) );
  XOR U21429 ( .A(n21686), .B(n21687), .Z(n21678) );
  AND U21430 ( .A(n918), .B(n21677), .Z(n21687) );
  XNOR U21431 ( .A(n21688), .B(n21675), .Z(n21677) );
  XOR U21432 ( .A(n21689), .B(n21690), .Z(n21675) );
  AND U21433 ( .A(n941), .B(n21691), .Z(n21690) );
  IV U21434 ( .A(n21686), .Z(n21688) );
  XOR U21435 ( .A(n21692), .B(n21693), .Z(n21686) );
  AND U21436 ( .A(n925), .B(n21685), .Z(n21693) );
  XNOR U21437 ( .A(n21683), .B(n21692), .Z(n21685) );
  XNOR U21438 ( .A(n21694), .B(n21695), .Z(n21683) );
  AND U21439 ( .A(n929), .B(n21696), .Z(n21695) );
  XOR U21440 ( .A(p_input[1360]), .B(n21694), .Z(n21696) );
  XNOR U21441 ( .A(n21697), .B(n21698), .Z(n21694) );
  AND U21442 ( .A(n933), .B(n21699), .Z(n21698) );
  XOR U21443 ( .A(n21700), .B(n21701), .Z(n21692) );
  AND U21444 ( .A(n937), .B(n21691), .Z(n21701) );
  XNOR U21445 ( .A(n21702), .B(n21689), .Z(n21691) );
  XOR U21446 ( .A(n21703), .B(n21704), .Z(n21689) );
  AND U21447 ( .A(n960), .B(n21705), .Z(n21704) );
  IV U21448 ( .A(n21700), .Z(n21702) );
  XOR U21449 ( .A(n21706), .B(n21707), .Z(n21700) );
  AND U21450 ( .A(n944), .B(n21699), .Z(n21707) );
  XNOR U21451 ( .A(n21697), .B(n21706), .Z(n21699) );
  XNOR U21452 ( .A(n21708), .B(n21709), .Z(n21697) );
  AND U21453 ( .A(n948), .B(n21710), .Z(n21709) );
  XOR U21454 ( .A(p_input[1392]), .B(n21708), .Z(n21710) );
  XNOR U21455 ( .A(n21711), .B(n21712), .Z(n21708) );
  AND U21456 ( .A(n952), .B(n21713), .Z(n21712) );
  XOR U21457 ( .A(n21714), .B(n21715), .Z(n21706) );
  AND U21458 ( .A(n956), .B(n21705), .Z(n21715) );
  XNOR U21459 ( .A(n21716), .B(n21703), .Z(n21705) );
  XOR U21460 ( .A(n21717), .B(n21718), .Z(n21703) );
  AND U21461 ( .A(n979), .B(n21719), .Z(n21718) );
  IV U21462 ( .A(n21714), .Z(n21716) );
  XOR U21463 ( .A(n21720), .B(n21721), .Z(n21714) );
  AND U21464 ( .A(n963), .B(n21713), .Z(n21721) );
  XNOR U21465 ( .A(n21711), .B(n21720), .Z(n21713) );
  XNOR U21466 ( .A(n21722), .B(n21723), .Z(n21711) );
  AND U21467 ( .A(n967), .B(n21724), .Z(n21723) );
  XOR U21468 ( .A(p_input[1424]), .B(n21722), .Z(n21724) );
  XNOR U21469 ( .A(n21725), .B(n21726), .Z(n21722) );
  AND U21470 ( .A(n971), .B(n21727), .Z(n21726) );
  XOR U21471 ( .A(n21728), .B(n21729), .Z(n21720) );
  AND U21472 ( .A(n975), .B(n21719), .Z(n21729) );
  XNOR U21473 ( .A(n21730), .B(n21717), .Z(n21719) );
  XOR U21474 ( .A(n21731), .B(n21732), .Z(n21717) );
  AND U21475 ( .A(n998), .B(n21733), .Z(n21732) );
  IV U21476 ( .A(n21728), .Z(n21730) );
  XOR U21477 ( .A(n21734), .B(n21735), .Z(n21728) );
  AND U21478 ( .A(n982), .B(n21727), .Z(n21735) );
  XNOR U21479 ( .A(n21725), .B(n21734), .Z(n21727) );
  XNOR U21480 ( .A(n21736), .B(n21737), .Z(n21725) );
  AND U21481 ( .A(n986), .B(n21738), .Z(n21737) );
  XOR U21482 ( .A(p_input[1456]), .B(n21736), .Z(n21738) );
  XNOR U21483 ( .A(n21739), .B(n21740), .Z(n21736) );
  AND U21484 ( .A(n990), .B(n21741), .Z(n21740) );
  XOR U21485 ( .A(n21742), .B(n21743), .Z(n21734) );
  AND U21486 ( .A(n994), .B(n21733), .Z(n21743) );
  XNOR U21487 ( .A(n21744), .B(n21731), .Z(n21733) );
  XOR U21488 ( .A(n21745), .B(n21746), .Z(n21731) );
  AND U21489 ( .A(n1017), .B(n21747), .Z(n21746) );
  IV U21490 ( .A(n21742), .Z(n21744) );
  XOR U21491 ( .A(n21748), .B(n21749), .Z(n21742) );
  AND U21492 ( .A(n1001), .B(n21741), .Z(n21749) );
  XNOR U21493 ( .A(n21739), .B(n21748), .Z(n21741) );
  XNOR U21494 ( .A(n21750), .B(n21751), .Z(n21739) );
  AND U21495 ( .A(n1005), .B(n21752), .Z(n21751) );
  XOR U21496 ( .A(p_input[1488]), .B(n21750), .Z(n21752) );
  XNOR U21497 ( .A(n21753), .B(n21754), .Z(n21750) );
  AND U21498 ( .A(n1009), .B(n21755), .Z(n21754) );
  XOR U21499 ( .A(n21756), .B(n21757), .Z(n21748) );
  AND U21500 ( .A(n1013), .B(n21747), .Z(n21757) );
  XNOR U21501 ( .A(n21758), .B(n21745), .Z(n21747) );
  XOR U21502 ( .A(n21759), .B(n21760), .Z(n21745) );
  AND U21503 ( .A(n1036), .B(n21761), .Z(n21760) );
  IV U21504 ( .A(n21756), .Z(n21758) );
  XOR U21505 ( .A(n21762), .B(n21763), .Z(n21756) );
  AND U21506 ( .A(n1020), .B(n21755), .Z(n21763) );
  XNOR U21507 ( .A(n21753), .B(n21762), .Z(n21755) );
  XNOR U21508 ( .A(n21764), .B(n21765), .Z(n21753) );
  AND U21509 ( .A(n1024), .B(n21766), .Z(n21765) );
  XOR U21510 ( .A(p_input[1520]), .B(n21764), .Z(n21766) );
  XNOR U21511 ( .A(n21767), .B(n21768), .Z(n21764) );
  AND U21512 ( .A(n1028), .B(n21769), .Z(n21768) );
  XOR U21513 ( .A(n21770), .B(n21771), .Z(n21762) );
  AND U21514 ( .A(n1032), .B(n21761), .Z(n21771) );
  XNOR U21515 ( .A(n21772), .B(n21759), .Z(n21761) );
  XOR U21516 ( .A(n21773), .B(n21774), .Z(n21759) );
  AND U21517 ( .A(n1055), .B(n21775), .Z(n21774) );
  IV U21518 ( .A(n21770), .Z(n21772) );
  XOR U21519 ( .A(n21776), .B(n21777), .Z(n21770) );
  AND U21520 ( .A(n1039), .B(n21769), .Z(n21777) );
  XNOR U21521 ( .A(n21767), .B(n21776), .Z(n21769) );
  XNOR U21522 ( .A(n21778), .B(n21779), .Z(n21767) );
  AND U21523 ( .A(n1043), .B(n21780), .Z(n21779) );
  XOR U21524 ( .A(p_input[1552]), .B(n21778), .Z(n21780) );
  XNOR U21525 ( .A(n21781), .B(n21782), .Z(n21778) );
  AND U21526 ( .A(n1047), .B(n21783), .Z(n21782) );
  XOR U21527 ( .A(n21784), .B(n21785), .Z(n21776) );
  AND U21528 ( .A(n1051), .B(n21775), .Z(n21785) );
  XNOR U21529 ( .A(n21786), .B(n21773), .Z(n21775) );
  XOR U21530 ( .A(n21787), .B(n21788), .Z(n21773) );
  AND U21531 ( .A(n1074), .B(n21789), .Z(n21788) );
  IV U21532 ( .A(n21784), .Z(n21786) );
  XOR U21533 ( .A(n21790), .B(n21791), .Z(n21784) );
  AND U21534 ( .A(n1058), .B(n21783), .Z(n21791) );
  XNOR U21535 ( .A(n21781), .B(n21790), .Z(n21783) );
  XNOR U21536 ( .A(n21792), .B(n21793), .Z(n21781) );
  AND U21537 ( .A(n1062), .B(n21794), .Z(n21793) );
  XOR U21538 ( .A(p_input[1584]), .B(n21792), .Z(n21794) );
  XNOR U21539 ( .A(n21795), .B(n21796), .Z(n21792) );
  AND U21540 ( .A(n1066), .B(n21797), .Z(n21796) );
  XOR U21541 ( .A(n21798), .B(n21799), .Z(n21790) );
  AND U21542 ( .A(n1070), .B(n21789), .Z(n21799) );
  XNOR U21543 ( .A(n21800), .B(n21787), .Z(n21789) );
  XOR U21544 ( .A(n21801), .B(n21802), .Z(n21787) );
  AND U21545 ( .A(n1093), .B(n21803), .Z(n21802) );
  IV U21546 ( .A(n21798), .Z(n21800) );
  XOR U21547 ( .A(n21804), .B(n21805), .Z(n21798) );
  AND U21548 ( .A(n1077), .B(n21797), .Z(n21805) );
  XNOR U21549 ( .A(n21795), .B(n21804), .Z(n21797) );
  XNOR U21550 ( .A(n21806), .B(n21807), .Z(n21795) );
  AND U21551 ( .A(n1081), .B(n21808), .Z(n21807) );
  XOR U21552 ( .A(p_input[1616]), .B(n21806), .Z(n21808) );
  XNOR U21553 ( .A(n21809), .B(n21810), .Z(n21806) );
  AND U21554 ( .A(n1085), .B(n21811), .Z(n21810) );
  XOR U21555 ( .A(n21812), .B(n21813), .Z(n21804) );
  AND U21556 ( .A(n1089), .B(n21803), .Z(n21813) );
  XNOR U21557 ( .A(n21814), .B(n21801), .Z(n21803) );
  XOR U21558 ( .A(n21815), .B(n21816), .Z(n21801) );
  AND U21559 ( .A(n1112), .B(n21817), .Z(n21816) );
  IV U21560 ( .A(n21812), .Z(n21814) );
  XOR U21561 ( .A(n21818), .B(n21819), .Z(n21812) );
  AND U21562 ( .A(n1096), .B(n21811), .Z(n21819) );
  XNOR U21563 ( .A(n21809), .B(n21818), .Z(n21811) );
  XNOR U21564 ( .A(n21820), .B(n21821), .Z(n21809) );
  AND U21565 ( .A(n1100), .B(n21822), .Z(n21821) );
  XOR U21566 ( .A(p_input[1648]), .B(n21820), .Z(n21822) );
  XNOR U21567 ( .A(n21823), .B(n21824), .Z(n21820) );
  AND U21568 ( .A(n1104), .B(n21825), .Z(n21824) );
  XOR U21569 ( .A(n21826), .B(n21827), .Z(n21818) );
  AND U21570 ( .A(n1108), .B(n21817), .Z(n21827) );
  XNOR U21571 ( .A(n21828), .B(n21815), .Z(n21817) );
  XOR U21572 ( .A(n21829), .B(n21830), .Z(n21815) );
  AND U21573 ( .A(n1131), .B(n21831), .Z(n21830) );
  IV U21574 ( .A(n21826), .Z(n21828) );
  XOR U21575 ( .A(n21832), .B(n21833), .Z(n21826) );
  AND U21576 ( .A(n1115), .B(n21825), .Z(n21833) );
  XNOR U21577 ( .A(n21823), .B(n21832), .Z(n21825) );
  XNOR U21578 ( .A(n21834), .B(n21835), .Z(n21823) );
  AND U21579 ( .A(n1119), .B(n21836), .Z(n21835) );
  XOR U21580 ( .A(p_input[1680]), .B(n21834), .Z(n21836) );
  XNOR U21581 ( .A(n21837), .B(n21838), .Z(n21834) );
  AND U21582 ( .A(n1123), .B(n21839), .Z(n21838) );
  XOR U21583 ( .A(n21840), .B(n21841), .Z(n21832) );
  AND U21584 ( .A(n1127), .B(n21831), .Z(n21841) );
  XNOR U21585 ( .A(n21842), .B(n21829), .Z(n21831) );
  XOR U21586 ( .A(n21843), .B(n21844), .Z(n21829) );
  AND U21587 ( .A(n1150), .B(n21845), .Z(n21844) );
  IV U21588 ( .A(n21840), .Z(n21842) );
  XOR U21589 ( .A(n21846), .B(n21847), .Z(n21840) );
  AND U21590 ( .A(n1134), .B(n21839), .Z(n21847) );
  XNOR U21591 ( .A(n21837), .B(n21846), .Z(n21839) );
  XNOR U21592 ( .A(n21848), .B(n21849), .Z(n21837) );
  AND U21593 ( .A(n1138), .B(n21850), .Z(n21849) );
  XOR U21594 ( .A(p_input[1712]), .B(n21848), .Z(n21850) );
  XNOR U21595 ( .A(n21851), .B(n21852), .Z(n21848) );
  AND U21596 ( .A(n1142), .B(n21853), .Z(n21852) );
  XOR U21597 ( .A(n21854), .B(n21855), .Z(n21846) );
  AND U21598 ( .A(n1146), .B(n21845), .Z(n21855) );
  XNOR U21599 ( .A(n21856), .B(n21843), .Z(n21845) );
  XOR U21600 ( .A(n21857), .B(n21858), .Z(n21843) );
  AND U21601 ( .A(n1169), .B(n21859), .Z(n21858) );
  IV U21602 ( .A(n21854), .Z(n21856) );
  XOR U21603 ( .A(n21860), .B(n21861), .Z(n21854) );
  AND U21604 ( .A(n1153), .B(n21853), .Z(n21861) );
  XNOR U21605 ( .A(n21851), .B(n21860), .Z(n21853) );
  XNOR U21606 ( .A(n21862), .B(n21863), .Z(n21851) );
  AND U21607 ( .A(n1157), .B(n21864), .Z(n21863) );
  XOR U21608 ( .A(p_input[1744]), .B(n21862), .Z(n21864) );
  XNOR U21609 ( .A(n21865), .B(n21866), .Z(n21862) );
  AND U21610 ( .A(n1161), .B(n21867), .Z(n21866) );
  XOR U21611 ( .A(n21868), .B(n21869), .Z(n21860) );
  AND U21612 ( .A(n1165), .B(n21859), .Z(n21869) );
  XNOR U21613 ( .A(n21870), .B(n21857), .Z(n21859) );
  XOR U21614 ( .A(n21871), .B(n21872), .Z(n21857) );
  AND U21615 ( .A(n1188), .B(n21873), .Z(n21872) );
  IV U21616 ( .A(n21868), .Z(n21870) );
  XOR U21617 ( .A(n21874), .B(n21875), .Z(n21868) );
  AND U21618 ( .A(n1172), .B(n21867), .Z(n21875) );
  XNOR U21619 ( .A(n21865), .B(n21874), .Z(n21867) );
  XNOR U21620 ( .A(n21876), .B(n21877), .Z(n21865) );
  AND U21621 ( .A(n1176), .B(n21878), .Z(n21877) );
  XOR U21622 ( .A(p_input[1776]), .B(n21876), .Z(n21878) );
  XNOR U21623 ( .A(n21879), .B(n21880), .Z(n21876) );
  AND U21624 ( .A(n1180), .B(n21881), .Z(n21880) );
  XOR U21625 ( .A(n21882), .B(n21883), .Z(n21874) );
  AND U21626 ( .A(n1184), .B(n21873), .Z(n21883) );
  XNOR U21627 ( .A(n21884), .B(n21871), .Z(n21873) );
  XOR U21628 ( .A(n21885), .B(n21886), .Z(n21871) );
  AND U21629 ( .A(n1207), .B(n21887), .Z(n21886) );
  IV U21630 ( .A(n21882), .Z(n21884) );
  XOR U21631 ( .A(n21888), .B(n21889), .Z(n21882) );
  AND U21632 ( .A(n1191), .B(n21881), .Z(n21889) );
  XNOR U21633 ( .A(n21879), .B(n21888), .Z(n21881) );
  XNOR U21634 ( .A(n21890), .B(n21891), .Z(n21879) );
  AND U21635 ( .A(n1195), .B(n21892), .Z(n21891) );
  XOR U21636 ( .A(p_input[1808]), .B(n21890), .Z(n21892) );
  XNOR U21637 ( .A(n21893), .B(n21894), .Z(n21890) );
  AND U21638 ( .A(n1199), .B(n21895), .Z(n21894) );
  XOR U21639 ( .A(n21896), .B(n21897), .Z(n21888) );
  AND U21640 ( .A(n1203), .B(n21887), .Z(n21897) );
  XNOR U21641 ( .A(n21898), .B(n21885), .Z(n21887) );
  XOR U21642 ( .A(n21899), .B(n21900), .Z(n21885) );
  AND U21643 ( .A(n1226), .B(n21901), .Z(n21900) );
  IV U21644 ( .A(n21896), .Z(n21898) );
  XOR U21645 ( .A(n21902), .B(n21903), .Z(n21896) );
  AND U21646 ( .A(n1210), .B(n21895), .Z(n21903) );
  XNOR U21647 ( .A(n21893), .B(n21902), .Z(n21895) );
  XNOR U21648 ( .A(n21904), .B(n21905), .Z(n21893) );
  AND U21649 ( .A(n1214), .B(n21906), .Z(n21905) );
  XOR U21650 ( .A(p_input[1840]), .B(n21904), .Z(n21906) );
  XNOR U21651 ( .A(n21907), .B(n21908), .Z(n21904) );
  AND U21652 ( .A(n1218), .B(n21909), .Z(n21908) );
  XOR U21653 ( .A(n21910), .B(n21911), .Z(n21902) );
  AND U21654 ( .A(n1222), .B(n21901), .Z(n21911) );
  XNOR U21655 ( .A(n21912), .B(n21899), .Z(n21901) );
  XOR U21656 ( .A(n21913), .B(n21914), .Z(n21899) );
  AND U21657 ( .A(n1245), .B(n21915), .Z(n21914) );
  IV U21658 ( .A(n21910), .Z(n21912) );
  XOR U21659 ( .A(n21916), .B(n21917), .Z(n21910) );
  AND U21660 ( .A(n1229), .B(n21909), .Z(n21917) );
  XNOR U21661 ( .A(n21907), .B(n21916), .Z(n21909) );
  XNOR U21662 ( .A(n21918), .B(n21919), .Z(n21907) );
  AND U21663 ( .A(n1233), .B(n21920), .Z(n21919) );
  XOR U21664 ( .A(p_input[1872]), .B(n21918), .Z(n21920) );
  XNOR U21665 ( .A(n21921), .B(n21922), .Z(n21918) );
  AND U21666 ( .A(n1237), .B(n21923), .Z(n21922) );
  XOR U21667 ( .A(n21924), .B(n21925), .Z(n21916) );
  AND U21668 ( .A(n1241), .B(n21915), .Z(n21925) );
  XNOR U21669 ( .A(n21926), .B(n21913), .Z(n21915) );
  XOR U21670 ( .A(n21927), .B(n21928), .Z(n21913) );
  AND U21671 ( .A(n1264), .B(n21929), .Z(n21928) );
  IV U21672 ( .A(n21924), .Z(n21926) );
  XOR U21673 ( .A(n21930), .B(n21931), .Z(n21924) );
  AND U21674 ( .A(n1248), .B(n21923), .Z(n21931) );
  XNOR U21675 ( .A(n21921), .B(n21930), .Z(n21923) );
  XNOR U21676 ( .A(n21932), .B(n21933), .Z(n21921) );
  AND U21677 ( .A(n1252), .B(n21934), .Z(n21933) );
  XOR U21678 ( .A(p_input[1904]), .B(n21932), .Z(n21934) );
  XNOR U21679 ( .A(n21935), .B(n21936), .Z(n21932) );
  AND U21680 ( .A(n1256), .B(n21937), .Z(n21936) );
  XOR U21681 ( .A(n21938), .B(n21939), .Z(n21930) );
  AND U21682 ( .A(n1260), .B(n21929), .Z(n21939) );
  XNOR U21683 ( .A(n21940), .B(n21927), .Z(n21929) );
  XOR U21684 ( .A(n21941), .B(n21942), .Z(n21927) );
  AND U21685 ( .A(n1282), .B(n21943), .Z(n21942) );
  IV U21686 ( .A(n21938), .Z(n21940) );
  XOR U21687 ( .A(n21944), .B(n21945), .Z(n21938) );
  AND U21688 ( .A(n1267), .B(n21937), .Z(n21945) );
  XNOR U21689 ( .A(n21935), .B(n21944), .Z(n21937) );
  XNOR U21690 ( .A(n21946), .B(n21947), .Z(n21935) );
  AND U21691 ( .A(n1271), .B(n21948), .Z(n21947) );
  XOR U21692 ( .A(p_input[1936]), .B(n21946), .Z(n21948) );
  XOR U21693 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][16] ), .B(n21949), 
        .Z(n21946) );
  AND U21694 ( .A(n1274), .B(n21950), .Z(n21949) );
  XOR U21695 ( .A(n21951), .B(n21952), .Z(n21944) );
  AND U21696 ( .A(n1278), .B(n21943), .Z(n21952) );
  XNOR U21697 ( .A(n21953), .B(n21941), .Z(n21943) );
  XOR U21698 ( .A(\knn_comb_/min_val_out[0][16] ), .B(n21954), .Z(n21941) );
  AND U21699 ( .A(n1290), .B(n21955), .Z(n21954) );
  IV U21700 ( .A(n21951), .Z(n21953) );
  XOR U21701 ( .A(n21956), .B(n21957), .Z(n21951) );
  AND U21702 ( .A(n1285), .B(n21950), .Z(n21957) );
  XOR U21703 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][16] ), .B(n21956), 
        .Z(n21950) );
  XOR U21704 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .B(n21958), 
        .Z(n21956) );
  AND U21705 ( .A(n1287), .B(n21955), .Z(n21958) );
  XOR U21706 ( .A(n21959), .B(n21960), .Z(n21955) );
  IV U21707 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .Z(n21960)
         );
  IV U21708 ( .A(\knn_comb_/min_val_out[0][16] ), .Z(n21959) );
  XOR U21709 ( .A(n109), .B(n21961), .Z(o[15]) );
  AND U21710 ( .A(n122), .B(n21962), .Z(n109) );
  XOR U21711 ( .A(n110), .B(n21961), .Z(n21962) );
  XOR U21712 ( .A(n21963), .B(n21964), .Z(n21961) );
  AND U21713 ( .A(n142), .B(n21965), .Z(n21964) );
  XOR U21714 ( .A(n21966), .B(n39), .Z(n110) );
  AND U21715 ( .A(n125), .B(n21967), .Z(n39) );
  XOR U21716 ( .A(n40), .B(n21966), .Z(n21967) );
  XOR U21717 ( .A(n21968), .B(n21969), .Z(n40) );
  AND U21718 ( .A(n130), .B(n21970), .Z(n21969) );
  XOR U21719 ( .A(p_input[15]), .B(n21968), .Z(n21970) );
  XNOR U21720 ( .A(n21971), .B(n21972), .Z(n21968) );
  AND U21721 ( .A(n134), .B(n21973), .Z(n21972) );
  XOR U21722 ( .A(n21974), .B(n21975), .Z(n21966) );
  AND U21723 ( .A(n138), .B(n21965), .Z(n21975) );
  XNOR U21724 ( .A(n21976), .B(n21963), .Z(n21965) );
  XOR U21725 ( .A(n21977), .B(n21978), .Z(n21963) );
  AND U21726 ( .A(n162), .B(n21979), .Z(n21978) );
  IV U21727 ( .A(n21974), .Z(n21976) );
  XOR U21728 ( .A(n21980), .B(n21981), .Z(n21974) );
  AND U21729 ( .A(n146), .B(n21973), .Z(n21981) );
  XNOR U21730 ( .A(n21971), .B(n21980), .Z(n21973) );
  XNOR U21731 ( .A(n21982), .B(n21983), .Z(n21971) );
  AND U21732 ( .A(n150), .B(n21984), .Z(n21983) );
  XOR U21733 ( .A(p_input[47]), .B(n21982), .Z(n21984) );
  XNOR U21734 ( .A(n21985), .B(n21986), .Z(n21982) );
  AND U21735 ( .A(n154), .B(n21987), .Z(n21986) );
  XOR U21736 ( .A(n21988), .B(n21989), .Z(n21980) );
  AND U21737 ( .A(n158), .B(n21979), .Z(n21989) );
  XNOR U21738 ( .A(n21990), .B(n21977), .Z(n21979) );
  XOR U21739 ( .A(n21991), .B(n21992), .Z(n21977) );
  AND U21740 ( .A(n181), .B(n21993), .Z(n21992) );
  IV U21741 ( .A(n21988), .Z(n21990) );
  XOR U21742 ( .A(n21994), .B(n21995), .Z(n21988) );
  AND U21743 ( .A(n165), .B(n21987), .Z(n21995) );
  XNOR U21744 ( .A(n21985), .B(n21994), .Z(n21987) );
  XNOR U21745 ( .A(n21996), .B(n21997), .Z(n21985) );
  AND U21746 ( .A(n169), .B(n21998), .Z(n21997) );
  XOR U21747 ( .A(p_input[79]), .B(n21996), .Z(n21998) );
  XNOR U21748 ( .A(n21999), .B(n22000), .Z(n21996) );
  AND U21749 ( .A(n173), .B(n22001), .Z(n22000) );
  XOR U21750 ( .A(n22002), .B(n22003), .Z(n21994) );
  AND U21751 ( .A(n177), .B(n21993), .Z(n22003) );
  XNOR U21752 ( .A(n22004), .B(n21991), .Z(n21993) );
  XOR U21753 ( .A(n22005), .B(n22006), .Z(n21991) );
  AND U21754 ( .A(n200), .B(n22007), .Z(n22006) );
  IV U21755 ( .A(n22002), .Z(n22004) );
  XOR U21756 ( .A(n22008), .B(n22009), .Z(n22002) );
  AND U21757 ( .A(n184), .B(n22001), .Z(n22009) );
  XNOR U21758 ( .A(n21999), .B(n22008), .Z(n22001) );
  XNOR U21759 ( .A(n22010), .B(n22011), .Z(n21999) );
  AND U21760 ( .A(n188), .B(n22012), .Z(n22011) );
  XOR U21761 ( .A(p_input[111]), .B(n22010), .Z(n22012) );
  XNOR U21762 ( .A(n22013), .B(n22014), .Z(n22010) );
  AND U21763 ( .A(n192), .B(n22015), .Z(n22014) );
  XOR U21764 ( .A(n22016), .B(n22017), .Z(n22008) );
  AND U21765 ( .A(n196), .B(n22007), .Z(n22017) );
  XNOR U21766 ( .A(n22018), .B(n22005), .Z(n22007) );
  XOR U21767 ( .A(n22019), .B(n22020), .Z(n22005) );
  AND U21768 ( .A(n219), .B(n22021), .Z(n22020) );
  IV U21769 ( .A(n22016), .Z(n22018) );
  XOR U21770 ( .A(n22022), .B(n22023), .Z(n22016) );
  AND U21771 ( .A(n203), .B(n22015), .Z(n22023) );
  XNOR U21772 ( .A(n22013), .B(n22022), .Z(n22015) );
  XNOR U21773 ( .A(n22024), .B(n22025), .Z(n22013) );
  AND U21774 ( .A(n207), .B(n22026), .Z(n22025) );
  XOR U21775 ( .A(p_input[143]), .B(n22024), .Z(n22026) );
  XNOR U21776 ( .A(n22027), .B(n22028), .Z(n22024) );
  AND U21777 ( .A(n211), .B(n22029), .Z(n22028) );
  XOR U21778 ( .A(n22030), .B(n22031), .Z(n22022) );
  AND U21779 ( .A(n215), .B(n22021), .Z(n22031) );
  XNOR U21780 ( .A(n22032), .B(n22019), .Z(n22021) );
  XOR U21781 ( .A(n22033), .B(n22034), .Z(n22019) );
  AND U21782 ( .A(n238), .B(n22035), .Z(n22034) );
  IV U21783 ( .A(n22030), .Z(n22032) );
  XOR U21784 ( .A(n22036), .B(n22037), .Z(n22030) );
  AND U21785 ( .A(n222), .B(n22029), .Z(n22037) );
  XNOR U21786 ( .A(n22027), .B(n22036), .Z(n22029) );
  XNOR U21787 ( .A(n22038), .B(n22039), .Z(n22027) );
  AND U21788 ( .A(n226), .B(n22040), .Z(n22039) );
  XOR U21789 ( .A(p_input[175]), .B(n22038), .Z(n22040) );
  XNOR U21790 ( .A(n22041), .B(n22042), .Z(n22038) );
  AND U21791 ( .A(n230), .B(n22043), .Z(n22042) );
  XOR U21792 ( .A(n22044), .B(n22045), .Z(n22036) );
  AND U21793 ( .A(n234), .B(n22035), .Z(n22045) );
  XNOR U21794 ( .A(n22046), .B(n22033), .Z(n22035) );
  XOR U21795 ( .A(n22047), .B(n22048), .Z(n22033) );
  AND U21796 ( .A(n257), .B(n22049), .Z(n22048) );
  IV U21797 ( .A(n22044), .Z(n22046) );
  XOR U21798 ( .A(n22050), .B(n22051), .Z(n22044) );
  AND U21799 ( .A(n241), .B(n22043), .Z(n22051) );
  XNOR U21800 ( .A(n22041), .B(n22050), .Z(n22043) );
  XNOR U21801 ( .A(n22052), .B(n22053), .Z(n22041) );
  AND U21802 ( .A(n245), .B(n22054), .Z(n22053) );
  XOR U21803 ( .A(p_input[207]), .B(n22052), .Z(n22054) );
  XNOR U21804 ( .A(n22055), .B(n22056), .Z(n22052) );
  AND U21805 ( .A(n249), .B(n22057), .Z(n22056) );
  XOR U21806 ( .A(n22058), .B(n22059), .Z(n22050) );
  AND U21807 ( .A(n253), .B(n22049), .Z(n22059) );
  XNOR U21808 ( .A(n22060), .B(n22047), .Z(n22049) );
  XOR U21809 ( .A(n22061), .B(n22062), .Z(n22047) );
  AND U21810 ( .A(n276), .B(n22063), .Z(n22062) );
  IV U21811 ( .A(n22058), .Z(n22060) );
  XOR U21812 ( .A(n22064), .B(n22065), .Z(n22058) );
  AND U21813 ( .A(n260), .B(n22057), .Z(n22065) );
  XNOR U21814 ( .A(n22055), .B(n22064), .Z(n22057) );
  XNOR U21815 ( .A(n22066), .B(n22067), .Z(n22055) );
  AND U21816 ( .A(n264), .B(n22068), .Z(n22067) );
  XOR U21817 ( .A(p_input[239]), .B(n22066), .Z(n22068) );
  XNOR U21818 ( .A(n22069), .B(n22070), .Z(n22066) );
  AND U21819 ( .A(n268), .B(n22071), .Z(n22070) );
  XOR U21820 ( .A(n22072), .B(n22073), .Z(n22064) );
  AND U21821 ( .A(n272), .B(n22063), .Z(n22073) );
  XNOR U21822 ( .A(n22074), .B(n22061), .Z(n22063) );
  XOR U21823 ( .A(n22075), .B(n22076), .Z(n22061) );
  AND U21824 ( .A(n295), .B(n22077), .Z(n22076) );
  IV U21825 ( .A(n22072), .Z(n22074) );
  XOR U21826 ( .A(n22078), .B(n22079), .Z(n22072) );
  AND U21827 ( .A(n279), .B(n22071), .Z(n22079) );
  XNOR U21828 ( .A(n22069), .B(n22078), .Z(n22071) );
  XNOR U21829 ( .A(n22080), .B(n22081), .Z(n22069) );
  AND U21830 ( .A(n283), .B(n22082), .Z(n22081) );
  XOR U21831 ( .A(p_input[271]), .B(n22080), .Z(n22082) );
  XNOR U21832 ( .A(n22083), .B(n22084), .Z(n22080) );
  AND U21833 ( .A(n287), .B(n22085), .Z(n22084) );
  XOR U21834 ( .A(n22086), .B(n22087), .Z(n22078) );
  AND U21835 ( .A(n291), .B(n22077), .Z(n22087) );
  XNOR U21836 ( .A(n22088), .B(n22075), .Z(n22077) );
  XOR U21837 ( .A(n22089), .B(n22090), .Z(n22075) );
  AND U21838 ( .A(n314), .B(n22091), .Z(n22090) );
  IV U21839 ( .A(n22086), .Z(n22088) );
  XOR U21840 ( .A(n22092), .B(n22093), .Z(n22086) );
  AND U21841 ( .A(n298), .B(n22085), .Z(n22093) );
  XNOR U21842 ( .A(n22083), .B(n22092), .Z(n22085) );
  XNOR U21843 ( .A(n22094), .B(n22095), .Z(n22083) );
  AND U21844 ( .A(n302), .B(n22096), .Z(n22095) );
  XOR U21845 ( .A(p_input[303]), .B(n22094), .Z(n22096) );
  XNOR U21846 ( .A(n22097), .B(n22098), .Z(n22094) );
  AND U21847 ( .A(n306), .B(n22099), .Z(n22098) );
  XOR U21848 ( .A(n22100), .B(n22101), .Z(n22092) );
  AND U21849 ( .A(n310), .B(n22091), .Z(n22101) );
  XNOR U21850 ( .A(n22102), .B(n22089), .Z(n22091) );
  XOR U21851 ( .A(n22103), .B(n22104), .Z(n22089) );
  AND U21852 ( .A(n333), .B(n22105), .Z(n22104) );
  IV U21853 ( .A(n22100), .Z(n22102) );
  XOR U21854 ( .A(n22106), .B(n22107), .Z(n22100) );
  AND U21855 ( .A(n317), .B(n22099), .Z(n22107) );
  XNOR U21856 ( .A(n22097), .B(n22106), .Z(n22099) );
  XNOR U21857 ( .A(n22108), .B(n22109), .Z(n22097) );
  AND U21858 ( .A(n321), .B(n22110), .Z(n22109) );
  XOR U21859 ( .A(p_input[335]), .B(n22108), .Z(n22110) );
  XNOR U21860 ( .A(n22111), .B(n22112), .Z(n22108) );
  AND U21861 ( .A(n325), .B(n22113), .Z(n22112) );
  XOR U21862 ( .A(n22114), .B(n22115), .Z(n22106) );
  AND U21863 ( .A(n329), .B(n22105), .Z(n22115) );
  XNOR U21864 ( .A(n22116), .B(n22103), .Z(n22105) );
  XOR U21865 ( .A(n22117), .B(n22118), .Z(n22103) );
  AND U21866 ( .A(n352), .B(n22119), .Z(n22118) );
  IV U21867 ( .A(n22114), .Z(n22116) );
  XOR U21868 ( .A(n22120), .B(n22121), .Z(n22114) );
  AND U21869 ( .A(n336), .B(n22113), .Z(n22121) );
  XNOR U21870 ( .A(n22111), .B(n22120), .Z(n22113) );
  XNOR U21871 ( .A(n22122), .B(n22123), .Z(n22111) );
  AND U21872 ( .A(n340), .B(n22124), .Z(n22123) );
  XOR U21873 ( .A(p_input[367]), .B(n22122), .Z(n22124) );
  XNOR U21874 ( .A(n22125), .B(n22126), .Z(n22122) );
  AND U21875 ( .A(n344), .B(n22127), .Z(n22126) );
  XOR U21876 ( .A(n22128), .B(n22129), .Z(n22120) );
  AND U21877 ( .A(n348), .B(n22119), .Z(n22129) );
  XNOR U21878 ( .A(n22130), .B(n22117), .Z(n22119) );
  XOR U21879 ( .A(n22131), .B(n22132), .Z(n22117) );
  AND U21880 ( .A(n371), .B(n22133), .Z(n22132) );
  IV U21881 ( .A(n22128), .Z(n22130) );
  XOR U21882 ( .A(n22134), .B(n22135), .Z(n22128) );
  AND U21883 ( .A(n355), .B(n22127), .Z(n22135) );
  XNOR U21884 ( .A(n22125), .B(n22134), .Z(n22127) );
  XNOR U21885 ( .A(n22136), .B(n22137), .Z(n22125) );
  AND U21886 ( .A(n359), .B(n22138), .Z(n22137) );
  XOR U21887 ( .A(p_input[399]), .B(n22136), .Z(n22138) );
  XNOR U21888 ( .A(n22139), .B(n22140), .Z(n22136) );
  AND U21889 ( .A(n363), .B(n22141), .Z(n22140) );
  XOR U21890 ( .A(n22142), .B(n22143), .Z(n22134) );
  AND U21891 ( .A(n367), .B(n22133), .Z(n22143) );
  XNOR U21892 ( .A(n22144), .B(n22131), .Z(n22133) );
  XOR U21893 ( .A(n22145), .B(n22146), .Z(n22131) );
  AND U21894 ( .A(n390), .B(n22147), .Z(n22146) );
  IV U21895 ( .A(n22142), .Z(n22144) );
  XOR U21896 ( .A(n22148), .B(n22149), .Z(n22142) );
  AND U21897 ( .A(n374), .B(n22141), .Z(n22149) );
  XNOR U21898 ( .A(n22139), .B(n22148), .Z(n22141) );
  XNOR U21899 ( .A(n22150), .B(n22151), .Z(n22139) );
  AND U21900 ( .A(n378), .B(n22152), .Z(n22151) );
  XOR U21901 ( .A(p_input[431]), .B(n22150), .Z(n22152) );
  XNOR U21902 ( .A(n22153), .B(n22154), .Z(n22150) );
  AND U21903 ( .A(n382), .B(n22155), .Z(n22154) );
  XOR U21904 ( .A(n22156), .B(n22157), .Z(n22148) );
  AND U21905 ( .A(n386), .B(n22147), .Z(n22157) );
  XNOR U21906 ( .A(n22158), .B(n22145), .Z(n22147) );
  XOR U21907 ( .A(n22159), .B(n22160), .Z(n22145) );
  AND U21908 ( .A(n409), .B(n22161), .Z(n22160) );
  IV U21909 ( .A(n22156), .Z(n22158) );
  XOR U21910 ( .A(n22162), .B(n22163), .Z(n22156) );
  AND U21911 ( .A(n393), .B(n22155), .Z(n22163) );
  XNOR U21912 ( .A(n22153), .B(n22162), .Z(n22155) );
  XNOR U21913 ( .A(n22164), .B(n22165), .Z(n22153) );
  AND U21914 ( .A(n397), .B(n22166), .Z(n22165) );
  XOR U21915 ( .A(p_input[463]), .B(n22164), .Z(n22166) );
  XNOR U21916 ( .A(n22167), .B(n22168), .Z(n22164) );
  AND U21917 ( .A(n401), .B(n22169), .Z(n22168) );
  XOR U21918 ( .A(n22170), .B(n22171), .Z(n22162) );
  AND U21919 ( .A(n405), .B(n22161), .Z(n22171) );
  XNOR U21920 ( .A(n22172), .B(n22159), .Z(n22161) );
  XOR U21921 ( .A(n22173), .B(n22174), .Z(n22159) );
  AND U21922 ( .A(n428), .B(n22175), .Z(n22174) );
  IV U21923 ( .A(n22170), .Z(n22172) );
  XOR U21924 ( .A(n22176), .B(n22177), .Z(n22170) );
  AND U21925 ( .A(n412), .B(n22169), .Z(n22177) );
  XNOR U21926 ( .A(n22167), .B(n22176), .Z(n22169) );
  XNOR U21927 ( .A(n22178), .B(n22179), .Z(n22167) );
  AND U21928 ( .A(n416), .B(n22180), .Z(n22179) );
  XOR U21929 ( .A(p_input[495]), .B(n22178), .Z(n22180) );
  XNOR U21930 ( .A(n22181), .B(n22182), .Z(n22178) );
  AND U21931 ( .A(n420), .B(n22183), .Z(n22182) );
  XOR U21932 ( .A(n22184), .B(n22185), .Z(n22176) );
  AND U21933 ( .A(n424), .B(n22175), .Z(n22185) );
  XNOR U21934 ( .A(n22186), .B(n22173), .Z(n22175) );
  XOR U21935 ( .A(n22187), .B(n22188), .Z(n22173) );
  AND U21936 ( .A(n447), .B(n22189), .Z(n22188) );
  IV U21937 ( .A(n22184), .Z(n22186) );
  XOR U21938 ( .A(n22190), .B(n22191), .Z(n22184) );
  AND U21939 ( .A(n431), .B(n22183), .Z(n22191) );
  XNOR U21940 ( .A(n22181), .B(n22190), .Z(n22183) );
  XNOR U21941 ( .A(n22192), .B(n22193), .Z(n22181) );
  AND U21942 ( .A(n435), .B(n22194), .Z(n22193) );
  XOR U21943 ( .A(p_input[527]), .B(n22192), .Z(n22194) );
  XNOR U21944 ( .A(n22195), .B(n22196), .Z(n22192) );
  AND U21945 ( .A(n439), .B(n22197), .Z(n22196) );
  XOR U21946 ( .A(n22198), .B(n22199), .Z(n22190) );
  AND U21947 ( .A(n443), .B(n22189), .Z(n22199) );
  XNOR U21948 ( .A(n22200), .B(n22187), .Z(n22189) );
  XOR U21949 ( .A(n22201), .B(n22202), .Z(n22187) );
  AND U21950 ( .A(n466), .B(n22203), .Z(n22202) );
  IV U21951 ( .A(n22198), .Z(n22200) );
  XOR U21952 ( .A(n22204), .B(n22205), .Z(n22198) );
  AND U21953 ( .A(n450), .B(n22197), .Z(n22205) );
  XNOR U21954 ( .A(n22195), .B(n22204), .Z(n22197) );
  XNOR U21955 ( .A(n22206), .B(n22207), .Z(n22195) );
  AND U21956 ( .A(n454), .B(n22208), .Z(n22207) );
  XOR U21957 ( .A(p_input[559]), .B(n22206), .Z(n22208) );
  XNOR U21958 ( .A(n22209), .B(n22210), .Z(n22206) );
  AND U21959 ( .A(n458), .B(n22211), .Z(n22210) );
  XOR U21960 ( .A(n22212), .B(n22213), .Z(n22204) );
  AND U21961 ( .A(n462), .B(n22203), .Z(n22213) );
  XNOR U21962 ( .A(n22214), .B(n22201), .Z(n22203) );
  XOR U21963 ( .A(n22215), .B(n22216), .Z(n22201) );
  AND U21964 ( .A(n485), .B(n22217), .Z(n22216) );
  IV U21965 ( .A(n22212), .Z(n22214) );
  XOR U21966 ( .A(n22218), .B(n22219), .Z(n22212) );
  AND U21967 ( .A(n469), .B(n22211), .Z(n22219) );
  XNOR U21968 ( .A(n22209), .B(n22218), .Z(n22211) );
  XNOR U21969 ( .A(n22220), .B(n22221), .Z(n22209) );
  AND U21970 ( .A(n473), .B(n22222), .Z(n22221) );
  XOR U21971 ( .A(p_input[591]), .B(n22220), .Z(n22222) );
  XNOR U21972 ( .A(n22223), .B(n22224), .Z(n22220) );
  AND U21973 ( .A(n477), .B(n22225), .Z(n22224) );
  XOR U21974 ( .A(n22226), .B(n22227), .Z(n22218) );
  AND U21975 ( .A(n481), .B(n22217), .Z(n22227) );
  XNOR U21976 ( .A(n22228), .B(n22215), .Z(n22217) );
  XOR U21977 ( .A(n22229), .B(n22230), .Z(n22215) );
  AND U21978 ( .A(n504), .B(n22231), .Z(n22230) );
  IV U21979 ( .A(n22226), .Z(n22228) );
  XOR U21980 ( .A(n22232), .B(n22233), .Z(n22226) );
  AND U21981 ( .A(n488), .B(n22225), .Z(n22233) );
  XNOR U21982 ( .A(n22223), .B(n22232), .Z(n22225) );
  XNOR U21983 ( .A(n22234), .B(n22235), .Z(n22223) );
  AND U21984 ( .A(n492), .B(n22236), .Z(n22235) );
  XOR U21985 ( .A(p_input[623]), .B(n22234), .Z(n22236) );
  XNOR U21986 ( .A(n22237), .B(n22238), .Z(n22234) );
  AND U21987 ( .A(n496), .B(n22239), .Z(n22238) );
  XOR U21988 ( .A(n22240), .B(n22241), .Z(n22232) );
  AND U21989 ( .A(n500), .B(n22231), .Z(n22241) );
  XNOR U21990 ( .A(n22242), .B(n22229), .Z(n22231) );
  XOR U21991 ( .A(n22243), .B(n22244), .Z(n22229) );
  AND U21992 ( .A(n523), .B(n22245), .Z(n22244) );
  IV U21993 ( .A(n22240), .Z(n22242) );
  XOR U21994 ( .A(n22246), .B(n22247), .Z(n22240) );
  AND U21995 ( .A(n507), .B(n22239), .Z(n22247) );
  XNOR U21996 ( .A(n22237), .B(n22246), .Z(n22239) );
  XNOR U21997 ( .A(n22248), .B(n22249), .Z(n22237) );
  AND U21998 ( .A(n511), .B(n22250), .Z(n22249) );
  XOR U21999 ( .A(p_input[655]), .B(n22248), .Z(n22250) );
  XNOR U22000 ( .A(n22251), .B(n22252), .Z(n22248) );
  AND U22001 ( .A(n515), .B(n22253), .Z(n22252) );
  XOR U22002 ( .A(n22254), .B(n22255), .Z(n22246) );
  AND U22003 ( .A(n519), .B(n22245), .Z(n22255) );
  XNOR U22004 ( .A(n22256), .B(n22243), .Z(n22245) );
  XOR U22005 ( .A(n22257), .B(n22258), .Z(n22243) );
  AND U22006 ( .A(n542), .B(n22259), .Z(n22258) );
  IV U22007 ( .A(n22254), .Z(n22256) );
  XOR U22008 ( .A(n22260), .B(n22261), .Z(n22254) );
  AND U22009 ( .A(n526), .B(n22253), .Z(n22261) );
  XNOR U22010 ( .A(n22251), .B(n22260), .Z(n22253) );
  XNOR U22011 ( .A(n22262), .B(n22263), .Z(n22251) );
  AND U22012 ( .A(n530), .B(n22264), .Z(n22263) );
  XOR U22013 ( .A(p_input[687]), .B(n22262), .Z(n22264) );
  XNOR U22014 ( .A(n22265), .B(n22266), .Z(n22262) );
  AND U22015 ( .A(n534), .B(n22267), .Z(n22266) );
  XOR U22016 ( .A(n22268), .B(n22269), .Z(n22260) );
  AND U22017 ( .A(n538), .B(n22259), .Z(n22269) );
  XNOR U22018 ( .A(n22270), .B(n22257), .Z(n22259) );
  XOR U22019 ( .A(n22271), .B(n22272), .Z(n22257) );
  AND U22020 ( .A(n561), .B(n22273), .Z(n22272) );
  IV U22021 ( .A(n22268), .Z(n22270) );
  XOR U22022 ( .A(n22274), .B(n22275), .Z(n22268) );
  AND U22023 ( .A(n545), .B(n22267), .Z(n22275) );
  XNOR U22024 ( .A(n22265), .B(n22274), .Z(n22267) );
  XNOR U22025 ( .A(n22276), .B(n22277), .Z(n22265) );
  AND U22026 ( .A(n549), .B(n22278), .Z(n22277) );
  XOR U22027 ( .A(p_input[719]), .B(n22276), .Z(n22278) );
  XNOR U22028 ( .A(n22279), .B(n22280), .Z(n22276) );
  AND U22029 ( .A(n553), .B(n22281), .Z(n22280) );
  XOR U22030 ( .A(n22282), .B(n22283), .Z(n22274) );
  AND U22031 ( .A(n557), .B(n22273), .Z(n22283) );
  XNOR U22032 ( .A(n22284), .B(n22271), .Z(n22273) );
  XOR U22033 ( .A(n22285), .B(n22286), .Z(n22271) );
  AND U22034 ( .A(n580), .B(n22287), .Z(n22286) );
  IV U22035 ( .A(n22282), .Z(n22284) );
  XOR U22036 ( .A(n22288), .B(n22289), .Z(n22282) );
  AND U22037 ( .A(n564), .B(n22281), .Z(n22289) );
  XNOR U22038 ( .A(n22279), .B(n22288), .Z(n22281) );
  XNOR U22039 ( .A(n22290), .B(n22291), .Z(n22279) );
  AND U22040 ( .A(n568), .B(n22292), .Z(n22291) );
  XOR U22041 ( .A(p_input[751]), .B(n22290), .Z(n22292) );
  XNOR U22042 ( .A(n22293), .B(n22294), .Z(n22290) );
  AND U22043 ( .A(n572), .B(n22295), .Z(n22294) );
  XOR U22044 ( .A(n22296), .B(n22297), .Z(n22288) );
  AND U22045 ( .A(n576), .B(n22287), .Z(n22297) );
  XNOR U22046 ( .A(n22298), .B(n22285), .Z(n22287) );
  XOR U22047 ( .A(n22299), .B(n22300), .Z(n22285) );
  AND U22048 ( .A(n599), .B(n22301), .Z(n22300) );
  IV U22049 ( .A(n22296), .Z(n22298) );
  XOR U22050 ( .A(n22302), .B(n22303), .Z(n22296) );
  AND U22051 ( .A(n583), .B(n22295), .Z(n22303) );
  XNOR U22052 ( .A(n22293), .B(n22302), .Z(n22295) );
  XNOR U22053 ( .A(n22304), .B(n22305), .Z(n22293) );
  AND U22054 ( .A(n587), .B(n22306), .Z(n22305) );
  XOR U22055 ( .A(p_input[783]), .B(n22304), .Z(n22306) );
  XNOR U22056 ( .A(n22307), .B(n22308), .Z(n22304) );
  AND U22057 ( .A(n591), .B(n22309), .Z(n22308) );
  XOR U22058 ( .A(n22310), .B(n22311), .Z(n22302) );
  AND U22059 ( .A(n595), .B(n22301), .Z(n22311) );
  XNOR U22060 ( .A(n22312), .B(n22299), .Z(n22301) );
  XOR U22061 ( .A(n22313), .B(n22314), .Z(n22299) );
  AND U22062 ( .A(n618), .B(n22315), .Z(n22314) );
  IV U22063 ( .A(n22310), .Z(n22312) );
  XOR U22064 ( .A(n22316), .B(n22317), .Z(n22310) );
  AND U22065 ( .A(n602), .B(n22309), .Z(n22317) );
  XNOR U22066 ( .A(n22307), .B(n22316), .Z(n22309) );
  XNOR U22067 ( .A(n22318), .B(n22319), .Z(n22307) );
  AND U22068 ( .A(n606), .B(n22320), .Z(n22319) );
  XOR U22069 ( .A(p_input[815]), .B(n22318), .Z(n22320) );
  XNOR U22070 ( .A(n22321), .B(n22322), .Z(n22318) );
  AND U22071 ( .A(n610), .B(n22323), .Z(n22322) );
  XOR U22072 ( .A(n22324), .B(n22325), .Z(n22316) );
  AND U22073 ( .A(n614), .B(n22315), .Z(n22325) );
  XNOR U22074 ( .A(n22326), .B(n22313), .Z(n22315) );
  XOR U22075 ( .A(n22327), .B(n22328), .Z(n22313) );
  AND U22076 ( .A(n637), .B(n22329), .Z(n22328) );
  IV U22077 ( .A(n22324), .Z(n22326) );
  XOR U22078 ( .A(n22330), .B(n22331), .Z(n22324) );
  AND U22079 ( .A(n621), .B(n22323), .Z(n22331) );
  XNOR U22080 ( .A(n22321), .B(n22330), .Z(n22323) );
  XNOR U22081 ( .A(n22332), .B(n22333), .Z(n22321) );
  AND U22082 ( .A(n625), .B(n22334), .Z(n22333) );
  XOR U22083 ( .A(p_input[847]), .B(n22332), .Z(n22334) );
  XNOR U22084 ( .A(n22335), .B(n22336), .Z(n22332) );
  AND U22085 ( .A(n629), .B(n22337), .Z(n22336) );
  XOR U22086 ( .A(n22338), .B(n22339), .Z(n22330) );
  AND U22087 ( .A(n633), .B(n22329), .Z(n22339) );
  XNOR U22088 ( .A(n22340), .B(n22327), .Z(n22329) );
  XOR U22089 ( .A(n22341), .B(n22342), .Z(n22327) );
  AND U22090 ( .A(n656), .B(n22343), .Z(n22342) );
  IV U22091 ( .A(n22338), .Z(n22340) );
  XOR U22092 ( .A(n22344), .B(n22345), .Z(n22338) );
  AND U22093 ( .A(n640), .B(n22337), .Z(n22345) );
  XNOR U22094 ( .A(n22335), .B(n22344), .Z(n22337) );
  XNOR U22095 ( .A(n22346), .B(n22347), .Z(n22335) );
  AND U22096 ( .A(n644), .B(n22348), .Z(n22347) );
  XOR U22097 ( .A(p_input[879]), .B(n22346), .Z(n22348) );
  XNOR U22098 ( .A(n22349), .B(n22350), .Z(n22346) );
  AND U22099 ( .A(n648), .B(n22351), .Z(n22350) );
  XOR U22100 ( .A(n22352), .B(n22353), .Z(n22344) );
  AND U22101 ( .A(n652), .B(n22343), .Z(n22353) );
  XNOR U22102 ( .A(n22354), .B(n22341), .Z(n22343) );
  XOR U22103 ( .A(n22355), .B(n22356), .Z(n22341) );
  AND U22104 ( .A(n675), .B(n22357), .Z(n22356) );
  IV U22105 ( .A(n22352), .Z(n22354) );
  XOR U22106 ( .A(n22358), .B(n22359), .Z(n22352) );
  AND U22107 ( .A(n659), .B(n22351), .Z(n22359) );
  XNOR U22108 ( .A(n22349), .B(n22358), .Z(n22351) );
  XNOR U22109 ( .A(n22360), .B(n22361), .Z(n22349) );
  AND U22110 ( .A(n663), .B(n22362), .Z(n22361) );
  XOR U22111 ( .A(p_input[911]), .B(n22360), .Z(n22362) );
  XNOR U22112 ( .A(n22363), .B(n22364), .Z(n22360) );
  AND U22113 ( .A(n667), .B(n22365), .Z(n22364) );
  XOR U22114 ( .A(n22366), .B(n22367), .Z(n22358) );
  AND U22115 ( .A(n671), .B(n22357), .Z(n22367) );
  XNOR U22116 ( .A(n22368), .B(n22355), .Z(n22357) );
  XOR U22117 ( .A(n22369), .B(n22370), .Z(n22355) );
  AND U22118 ( .A(n694), .B(n22371), .Z(n22370) );
  IV U22119 ( .A(n22366), .Z(n22368) );
  XOR U22120 ( .A(n22372), .B(n22373), .Z(n22366) );
  AND U22121 ( .A(n678), .B(n22365), .Z(n22373) );
  XNOR U22122 ( .A(n22363), .B(n22372), .Z(n22365) );
  XNOR U22123 ( .A(n22374), .B(n22375), .Z(n22363) );
  AND U22124 ( .A(n682), .B(n22376), .Z(n22375) );
  XOR U22125 ( .A(p_input[943]), .B(n22374), .Z(n22376) );
  XNOR U22126 ( .A(n22377), .B(n22378), .Z(n22374) );
  AND U22127 ( .A(n686), .B(n22379), .Z(n22378) );
  XOR U22128 ( .A(n22380), .B(n22381), .Z(n22372) );
  AND U22129 ( .A(n690), .B(n22371), .Z(n22381) );
  XNOR U22130 ( .A(n22382), .B(n22369), .Z(n22371) );
  XOR U22131 ( .A(n22383), .B(n22384), .Z(n22369) );
  AND U22132 ( .A(n713), .B(n22385), .Z(n22384) );
  IV U22133 ( .A(n22380), .Z(n22382) );
  XOR U22134 ( .A(n22386), .B(n22387), .Z(n22380) );
  AND U22135 ( .A(n697), .B(n22379), .Z(n22387) );
  XNOR U22136 ( .A(n22377), .B(n22386), .Z(n22379) );
  XNOR U22137 ( .A(n22388), .B(n22389), .Z(n22377) );
  AND U22138 ( .A(n701), .B(n22390), .Z(n22389) );
  XOR U22139 ( .A(p_input[975]), .B(n22388), .Z(n22390) );
  XNOR U22140 ( .A(n22391), .B(n22392), .Z(n22388) );
  AND U22141 ( .A(n705), .B(n22393), .Z(n22392) );
  XOR U22142 ( .A(n22394), .B(n22395), .Z(n22386) );
  AND U22143 ( .A(n709), .B(n22385), .Z(n22395) );
  XNOR U22144 ( .A(n22396), .B(n22383), .Z(n22385) );
  XOR U22145 ( .A(n22397), .B(n22398), .Z(n22383) );
  AND U22146 ( .A(n732), .B(n22399), .Z(n22398) );
  IV U22147 ( .A(n22394), .Z(n22396) );
  XOR U22148 ( .A(n22400), .B(n22401), .Z(n22394) );
  AND U22149 ( .A(n716), .B(n22393), .Z(n22401) );
  XNOR U22150 ( .A(n22391), .B(n22400), .Z(n22393) );
  XNOR U22151 ( .A(n22402), .B(n22403), .Z(n22391) );
  AND U22152 ( .A(n720), .B(n22404), .Z(n22403) );
  XOR U22153 ( .A(p_input[1007]), .B(n22402), .Z(n22404) );
  XNOR U22154 ( .A(n22405), .B(n22406), .Z(n22402) );
  AND U22155 ( .A(n724), .B(n22407), .Z(n22406) );
  XOR U22156 ( .A(n22408), .B(n22409), .Z(n22400) );
  AND U22157 ( .A(n728), .B(n22399), .Z(n22409) );
  XNOR U22158 ( .A(n22410), .B(n22397), .Z(n22399) );
  XOR U22159 ( .A(n22411), .B(n22412), .Z(n22397) );
  AND U22160 ( .A(n751), .B(n22413), .Z(n22412) );
  IV U22161 ( .A(n22408), .Z(n22410) );
  XOR U22162 ( .A(n22414), .B(n22415), .Z(n22408) );
  AND U22163 ( .A(n735), .B(n22407), .Z(n22415) );
  XNOR U22164 ( .A(n22405), .B(n22414), .Z(n22407) );
  XNOR U22165 ( .A(n22416), .B(n22417), .Z(n22405) );
  AND U22166 ( .A(n739), .B(n22418), .Z(n22417) );
  XOR U22167 ( .A(p_input[1039]), .B(n22416), .Z(n22418) );
  XNOR U22168 ( .A(n22419), .B(n22420), .Z(n22416) );
  AND U22169 ( .A(n743), .B(n22421), .Z(n22420) );
  XOR U22170 ( .A(n22422), .B(n22423), .Z(n22414) );
  AND U22171 ( .A(n747), .B(n22413), .Z(n22423) );
  XNOR U22172 ( .A(n22424), .B(n22411), .Z(n22413) );
  XOR U22173 ( .A(n22425), .B(n22426), .Z(n22411) );
  AND U22174 ( .A(n770), .B(n22427), .Z(n22426) );
  IV U22175 ( .A(n22422), .Z(n22424) );
  XOR U22176 ( .A(n22428), .B(n22429), .Z(n22422) );
  AND U22177 ( .A(n754), .B(n22421), .Z(n22429) );
  XNOR U22178 ( .A(n22419), .B(n22428), .Z(n22421) );
  XNOR U22179 ( .A(n22430), .B(n22431), .Z(n22419) );
  AND U22180 ( .A(n758), .B(n22432), .Z(n22431) );
  XOR U22181 ( .A(p_input[1071]), .B(n22430), .Z(n22432) );
  XNOR U22182 ( .A(n22433), .B(n22434), .Z(n22430) );
  AND U22183 ( .A(n762), .B(n22435), .Z(n22434) );
  XOR U22184 ( .A(n22436), .B(n22437), .Z(n22428) );
  AND U22185 ( .A(n766), .B(n22427), .Z(n22437) );
  XNOR U22186 ( .A(n22438), .B(n22425), .Z(n22427) );
  XOR U22187 ( .A(n22439), .B(n22440), .Z(n22425) );
  AND U22188 ( .A(n789), .B(n22441), .Z(n22440) );
  IV U22189 ( .A(n22436), .Z(n22438) );
  XOR U22190 ( .A(n22442), .B(n22443), .Z(n22436) );
  AND U22191 ( .A(n773), .B(n22435), .Z(n22443) );
  XNOR U22192 ( .A(n22433), .B(n22442), .Z(n22435) );
  XNOR U22193 ( .A(n22444), .B(n22445), .Z(n22433) );
  AND U22194 ( .A(n777), .B(n22446), .Z(n22445) );
  XOR U22195 ( .A(p_input[1103]), .B(n22444), .Z(n22446) );
  XNOR U22196 ( .A(n22447), .B(n22448), .Z(n22444) );
  AND U22197 ( .A(n781), .B(n22449), .Z(n22448) );
  XOR U22198 ( .A(n22450), .B(n22451), .Z(n22442) );
  AND U22199 ( .A(n785), .B(n22441), .Z(n22451) );
  XNOR U22200 ( .A(n22452), .B(n22439), .Z(n22441) );
  XOR U22201 ( .A(n22453), .B(n22454), .Z(n22439) );
  AND U22202 ( .A(n808), .B(n22455), .Z(n22454) );
  IV U22203 ( .A(n22450), .Z(n22452) );
  XOR U22204 ( .A(n22456), .B(n22457), .Z(n22450) );
  AND U22205 ( .A(n792), .B(n22449), .Z(n22457) );
  XNOR U22206 ( .A(n22447), .B(n22456), .Z(n22449) );
  XNOR U22207 ( .A(n22458), .B(n22459), .Z(n22447) );
  AND U22208 ( .A(n796), .B(n22460), .Z(n22459) );
  XOR U22209 ( .A(p_input[1135]), .B(n22458), .Z(n22460) );
  XNOR U22210 ( .A(n22461), .B(n22462), .Z(n22458) );
  AND U22211 ( .A(n800), .B(n22463), .Z(n22462) );
  XOR U22212 ( .A(n22464), .B(n22465), .Z(n22456) );
  AND U22213 ( .A(n804), .B(n22455), .Z(n22465) );
  XNOR U22214 ( .A(n22466), .B(n22453), .Z(n22455) );
  XOR U22215 ( .A(n22467), .B(n22468), .Z(n22453) );
  AND U22216 ( .A(n827), .B(n22469), .Z(n22468) );
  IV U22217 ( .A(n22464), .Z(n22466) );
  XOR U22218 ( .A(n22470), .B(n22471), .Z(n22464) );
  AND U22219 ( .A(n811), .B(n22463), .Z(n22471) );
  XNOR U22220 ( .A(n22461), .B(n22470), .Z(n22463) );
  XNOR U22221 ( .A(n22472), .B(n22473), .Z(n22461) );
  AND U22222 ( .A(n815), .B(n22474), .Z(n22473) );
  XOR U22223 ( .A(p_input[1167]), .B(n22472), .Z(n22474) );
  XNOR U22224 ( .A(n22475), .B(n22476), .Z(n22472) );
  AND U22225 ( .A(n819), .B(n22477), .Z(n22476) );
  XOR U22226 ( .A(n22478), .B(n22479), .Z(n22470) );
  AND U22227 ( .A(n823), .B(n22469), .Z(n22479) );
  XNOR U22228 ( .A(n22480), .B(n22467), .Z(n22469) );
  XOR U22229 ( .A(n22481), .B(n22482), .Z(n22467) );
  AND U22230 ( .A(n846), .B(n22483), .Z(n22482) );
  IV U22231 ( .A(n22478), .Z(n22480) );
  XOR U22232 ( .A(n22484), .B(n22485), .Z(n22478) );
  AND U22233 ( .A(n830), .B(n22477), .Z(n22485) );
  XNOR U22234 ( .A(n22475), .B(n22484), .Z(n22477) );
  XNOR U22235 ( .A(n22486), .B(n22487), .Z(n22475) );
  AND U22236 ( .A(n834), .B(n22488), .Z(n22487) );
  XOR U22237 ( .A(p_input[1199]), .B(n22486), .Z(n22488) );
  XNOR U22238 ( .A(n22489), .B(n22490), .Z(n22486) );
  AND U22239 ( .A(n838), .B(n22491), .Z(n22490) );
  XOR U22240 ( .A(n22492), .B(n22493), .Z(n22484) );
  AND U22241 ( .A(n842), .B(n22483), .Z(n22493) );
  XNOR U22242 ( .A(n22494), .B(n22481), .Z(n22483) );
  XOR U22243 ( .A(n22495), .B(n22496), .Z(n22481) );
  AND U22244 ( .A(n865), .B(n22497), .Z(n22496) );
  IV U22245 ( .A(n22492), .Z(n22494) );
  XOR U22246 ( .A(n22498), .B(n22499), .Z(n22492) );
  AND U22247 ( .A(n849), .B(n22491), .Z(n22499) );
  XNOR U22248 ( .A(n22489), .B(n22498), .Z(n22491) );
  XNOR U22249 ( .A(n22500), .B(n22501), .Z(n22489) );
  AND U22250 ( .A(n853), .B(n22502), .Z(n22501) );
  XOR U22251 ( .A(p_input[1231]), .B(n22500), .Z(n22502) );
  XNOR U22252 ( .A(n22503), .B(n22504), .Z(n22500) );
  AND U22253 ( .A(n857), .B(n22505), .Z(n22504) );
  XOR U22254 ( .A(n22506), .B(n22507), .Z(n22498) );
  AND U22255 ( .A(n861), .B(n22497), .Z(n22507) );
  XNOR U22256 ( .A(n22508), .B(n22495), .Z(n22497) );
  XOR U22257 ( .A(n22509), .B(n22510), .Z(n22495) );
  AND U22258 ( .A(n884), .B(n22511), .Z(n22510) );
  IV U22259 ( .A(n22506), .Z(n22508) );
  XOR U22260 ( .A(n22512), .B(n22513), .Z(n22506) );
  AND U22261 ( .A(n868), .B(n22505), .Z(n22513) );
  XNOR U22262 ( .A(n22503), .B(n22512), .Z(n22505) );
  XNOR U22263 ( .A(n22514), .B(n22515), .Z(n22503) );
  AND U22264 ( .A(n872), .B(n22516), .Z(n22515) );
  XOR U22265 ( .A(p_input[1263]), .B(n22514), .Z(n22516) );
  XNOR U22266 ( .A(n22517), .B(n22518), .Z(n22514) );
  AND U22267 ( .A(n876), .B(n22519), .Z(n22518) );
  XOR U22268 ( .A(n22520), .B(n22521), .Z(n22512) );
  AND U22269 ( .A(n880), .B(n22511), .Z(n22521) );
  XNOR U22270 ( .A(n22522), .B(n22509), .Z(n22511) );
  XOR U22271 ( .A(n22523), .B(n22524), .Z(n22509) );
  AND U22272 ( .A(n903), .B(n22525), .Z(n22524) );
  IV U22273 ( .A(n22520), .Z(n22522) );
  XOR U22274 ( .A(n22526), .B(n22527), .Z(n22520) );
  AND U22275 ( .A(n887), .B(n22519), .Z(n22527) );
  XNOR U22276 ( .A(n22517), .B(n22526), .Z(n22519) );
  XNOR U22277 ( .A(n22528), .B(n22529), .Z(n22517) );
  AND U22278 ( .A(n891), .B(n22530), .Z(n22529) );
  XOR U22279 ( .A(p_input[1295]), .B(n22528), .Z(n22530) );
  XNOR U22280 ( .A(n22531), .B(n22532), .Z(n22528) );
  AND U22281 ( .A(n895), .B(n22533), .Z(n22532) );
  XOR U22282 ( .A(n22534), .B(n22535), .Z(n22526) );
  AND U22283 ( .A(n899), .B(n22525), .Z(n22535) );
  XNOR U22284 ( .A(n22536), .B(n22523), .Z(n22525) );
  XOR U22285 ( .A(n22537), .B(n22538), .Z(n22523) );
  AND U22286 ( .A(n922), .B(n22539), .Z(n22538) );
  IV U22287 ( .A(n22534), .Z(n22536) );
  XOR U22288 ( .A(n22540), .B(n22541), .Z(n22534) );
  AND U22289 ( .A(n906), .B(n22533), .Z(n22541) );
  XNOR U22290 ( .A(n22531), .B(n22540), .Z(n22533) );
  XNOR U22291 ( .A(n22542), .B(n22543), .Z(n22531) );
  AND U22292 ( .A(n910), .B(n22544), .Z(n22543) );
  XOR U22293 ( .A(p_input[1327]), .B(n22542), .Z(n22544) );
  XNOR U22294 ( .A(n22545), .B(n22546), .Z(n22542) );
  AND U22295 ( .A(n914), .B(n22547), .Z(n22546) );
  XOR U22296 ( .A(n22548), .B(n22549), .Z(n22540) );
  AND U22297 ( .A(n918), .B(n22539), .Z(n22549) );
  XNOR U22298 ( .A(n22550), .B(n22537), .Z(n22539) );
  XOR U22299 ( .A(n22551), .B(n22552), .Z(n22537) );
  AND U22300 ( .A(n941), .B(n22553), .Z(n22552) );
  IV U22301 ( .A(n22548), .Z(n22550) );
  XOR U22302 ( .A(n22554), .B(n22555), .Z(n22548) );
  AND U22303 ( .A(n925), .B(n22547), .Z(n22555) );
  XNOR U22304 ( .A(n22545), .B(n22554), .Z(n22547) );
  XNOR U22305 ( .A(n22556), .B(n22557), .Z(n22545) );
  AND U22306 ( .A(n929), .B(n22558), .Z(n22557) );
  XOR U22307 ( .A(p_input[1359]), .B(n22556), .Z(n22558) );
  XNOR U22308 ( .A(n22559), .B(n22560), .Z(n22556) );
  AND U22309 ( .A(n933), .B(n22561), .Z(n22560) );
  XOR U22310 ( .A(n22562), .B(n22563), .Z(n22554) );
  AND U22311 ( .A(n937), .B(n22553), .Z(n22563) );
  XNOR U22312 ( .A(n22564), .B(n22551), .Z(n22553) );
  XOR U22313 ( .A(n22565), .B(n22566), .Z(n22551) );
  AND U22314 ( .A(n960), .B(n22567), .Z(n22566) );
  IV U22315 ( .A(n22562), .Z(n22564) );
  XOR U22316 ( .A(n22568), .B(n22569), .Z(n22562) );
  AND U22317 ( .A(n944), .B(n22561), .Z(n22569) );
  XNOR U22318 ( .A(n22559), .B(n22568), .Z(n22561) );
  XNOR U22319 ( .A(n22570), .B(n22571), .Z(n22559) );
  AND U22320 ( .A(n948), .B(n22572), .Z(n22571) );
  XOR U22321 ( .A(p_input[1391]), .B(n22570), .Z(n22572) );
  XNOR U22322 ( .A(n22573), .B(n22574), .Z(n22570) );
  AND U22323 ( .A(n952), .B(n22575), .Z(n22574) );
  XOR U22324 ( .A(n22576), .B(n22577), .Z(n22568) );
  AND U22325 ( .A(n956), .B(n22567), .Z(n22577) );
  XNOR U22326 ( .A(n22578), .B(n22565), .Z(n22567) );
  XOR U22327 ( .A(n22579), .B(n22580), .Z(n22565) );
  AND U22328 ( .A(n979), .B(n22581), .Z(n22580) );
  IV U22329 ( .A(n22576), .Z(n22578) );
  XOR U22330 ( .A(n22582), .B(n22583), .Z(n22576) );
  AND U22331 ( .A(n963), .B(n22575), .Z(n22583) );
  XNOR U22332 ( .A(n22573), .B(n22582), .Z(n22575) );
  XNOR U22333 ( .A(n22584), .B(n22585), .Z(n22573) );
  AND U22334 ( .A(n967), .B(n22586), .Z(n22585) );
  XOR U22335 ( .A(p_input[1423]), .B(n22584), .Z(n22586) );
  XNOR U22336 ( .A(n22587), .B(n22588), .Z(n22584) );
  AND U22337 ( .A(n971), .B(n22589), .Z(n22588) );
  XOR U22338 ( .A(n22590), .B(n22591), .Z(n22582) );
  AND U22339 ( .A(n975), .B(n22581), .Z(n22591) );
  XNOR U22340 ( .A(n22592), .B(n22579), .Z(n22581) );
  XOR U22341 ( .A(n22593), .B(n22594), .Z(n22579) );
  AND U22342 ( .A(n998), .B(n22595), .Z(n22594) );
  IV U22343 ( .A(n22590), .Z(n22592) );
  XOR U22344 ( .A(n22596), .B(n22597), .Z(n22590) );
  AND U22345 ( .A(n982), .B(n22589), .Z(n22597) );
  XNOR U22346 ( .A(n22587), .B(n22596), .Z(n22589) );
  XNOR U22347 ( .A(n22598), .B(n22599), .Z(n22587) );
  AND U22348 ( .A(n986), .B(n22600), .Z(n22599) );
  XOR U22349 ( .A(p_input[1455]), .B(n22598), .Z(n22600) );
  XNOR U22350 ( .A(n22601), .B(n22602), .Z(n22598) );
  AND U22351 ( .A(n990), .B(n22603), .Z(n22602) );
  XOR U22352 ( .A(n22604), .B(n22605), .Z(n22596) );
  AND U22353 ( .A(n994), .B(n22595), .Z(n22605) );
  XNOR U22354 ( .A(n22606), .B(n22593), .Z(n22595) );
  XOR U22355 ( .A(n22607), .B(n22608), .Z(n22593) );
  AND U22356 ( .A(n1017), .B(n22609), .Z(n22608) );
  IV U22357 ( .A(n22604), .Z(n22606) );
  XOR U22358 ( .A(n22610), .B(n22611), .Z(n22604) );
  AND U22359 ( .A(n1001), .B(n22603), .Z(n22611) );
  XNOR U22360 ( .A(n22601), .B(n22610), .Z(n22603) );
  XNOR U22361 ( .A(n22612), .B(n22613), .Z(n22601) );
  AND U22362 ( .A(n1005), .B(n22614), .Z(n22613) );
  XOR U22363 ( .A(p_input[1487]), .B(n22612), .Z(n22614) );
  XNOR U22364 ( .A(n22615), .B(n22616), .Z(n22612) );
  AND U22365 ( .A(n1009), .B(n22617), .Z(n22616) );
  XOR U22366 ( .A(n22618), .B(n22619), .Z(n22610) );
  AND U22367 ( .A(n1013), .B(n22609), .Z(n22619) );
  XNOR U22368 ( .A(n22620), .B(n22607), .Z(n22609) );
  XOR U22369 ( .A(n22621), .B(n22622), .Z(n22607) );
  AND U22370 ( .A(n1036), .B(n22623), .Z(n22622) );
  IV U22371 ( .A(n22618), .Z(n22620) );
  XOR U22372 ( .A(n22624), .B(n22625), .Z(n22618) );
  AND U22373 ( .A(n1020), .B(n22617), .Z(n22625) );
  XNOR U22374 ( .A(n22615), .B(n22624), .Z(n22617) );
  XNOR U22375 ( .A(n22626), .B(n22627), .Z(n22615) );
  AND U22376 ( .A(n1024), .B(n22628), .Z(n22627) );
  XOR U22377 ( .A(p_input[1519]), .B(n22626), .Z(n22628) );
  XNOR U22378 ( .A(n22629), .B(n22630), .Z(n22626) );
  AND U22379 ( .A(n1028), .B(n22631), .Z(n22630) );
  XOR U22380 ( .A(n22632), .B(n22633), .Z(n22624) );
  AND U22381 ( .A(n1032), .B(n22623), .Z(n22633) );
  XNOR U22382 ( .A(n22634), .B(n22621), .Z(n22623) );
  XOR U22383 ( .A(n22635), .B(n22636), .Z(n22621) );
  AND U22384 ( .A(n1055), .B(n22637), .Z(n22636) );
  IV U22385 ( .A(n22632), .Z(n22634) );
  XOR U22386 ( .A(n22638), .B(n22639), .Z(n22632) );
  AND U22387 ( .A(n1039), .B(n22631), .Z(n22639) );
  XNOR U22388 ( .A(n22629), .B(n22638), .Z(n22631) );
  XNOR U22389 ( .A(n22640), .B(n22641), .Z(n22629) );
  AND U22390 ( .A(n1043), .B(n22642), .Z(n22641) );
  XOR U22391 ( .A(p_input[1551]), .B(n22640), .Z(n22642) );
  XNOR U22392 ( .A(n22643), .B(n22644), .Z(n22640) );
  AND U22393 ( .A(n1047), .B(n22645), .Z(n22644) );
  XOR U22394 ( .A(n22646), .B(n22647), .Z(n22638) );
  AND U22395 ( .A(n1051), .B(n22637), .Z(n22647) );
  XNOR U22396 ( .A(n22648), .B(n22635), .Z(n22637) );
  XOR U22397 ( .A(n22649), .B(n22650), .Z(n22635) );
  AND U22398 ( .A(n1074), .B(n22651), .Z(n22650) );
  IV U22399 ( .A(n22646), .Z(n22648) );
  XOR U22400 ( .A(n22652), .B(n22653), .Z(n22646) );
  AND U22401 ( .A(n1058), .B(n22645), .Z(n22653) );
  XNOR U22402 ( .A(n22643), .B(n22652), .Z(n22645) );
  XNOR U22403 ( .A(n22654), .B(n22655), .Z(n22643) );
  AND U22404 ( .A(n1062), .B(n22656), .Z(n22655) );
  XOR U22405 ( .A(p_input[1583]), .B(n22654), .Z(n22656) );
  XNOR U22406 ( .A(n22657), .B(n22658), .Z(n22654) );
  AND U22407 ( .A(n1066), .B(n22659), .Z(n22658) );
  XOR U22408 ( .A(n22660), .B(n22661), .Z(n22652) );
  AND U22409 ( .A(n1070), .B(n22651), .Z(n22661) );
  XNOR U22410 ( .A(n22662), .B(n22649), .Z(n22651) );
  XOR U22411 ( .A(n22663), .B(n22664), .Z(n22649) );
  AND U22412 ( .A(n1093), .B(n22665), .Z(n22664) );
  IV U22413 ( .A(n22660), .Z(n22662) );
  XOR U22414 ( .A(n22666), .B(n22667), .Z(n22660) );
  AND U22415 ( .A(n1077), .B(n22659), .Z(n22667) );
  XNOR U22416 ( .A(n22657), .B(n22666), .Z(n22659) );
  XNOR U22417 ( .A(n22668), .B(n22669), .Z(n22657) );
  AND U22418 ( .A(n1081), .B(n22670), .Z(n22669) );
  XOR U22419 ( .A(p_input[1615]), .B(n22668), .Z(n22670) );
  XNOR U22420 ( .A(n22671), .B(n22672), .Z(n22668) );
  AND U22421 ( .A(n1085), .B(n22673), .Z(n22672) );
  XOR U22422 ( .A(n22674), .B(n22675), .Z(n22666) );
  AND U22423 ( .A(n1089), .B(n22665), .Z(n22675) );
  XNOR U22424 ( .A(n22676), .B(n22663), .Z(n22665) );
  XOR U22425 ( .A(n22677), .B(n22678), .Z(n22663) );
  AND U22426 ( .A(n1112), .B(n22679), .Z(n22678) );
  IV U22427 ( .A(n22674), .Z(n22676) );
  XOR U22428 ( .A(n22680), .B(n22681), .Z(n22674) );
  AND U22429 ( .A(n1096), .B(n22673), .Z(n22681) );
  XNOR U22430 ( .A(n22671), .B(n22680), .Z(n22673) );
  XNOR U22431 ( .A(n22682), .B(n22683), .Z(n22671) );
  AND U22432 ( .A(n1100), .B(n22684), .Z(n22683) );
  XOR U22433 ( .A(p_input[1647]), .B(n22682), .Z(n22684) );
  XNOR U22434 ( .A(n22685), .B(n22686), .Z(n22682) );
  AND U22435 ( .A(n1104), .B(n22687), .Z(n22686) );
  XOR U22436 ( .A(n22688), .B(n22689), .Z(n22680) );
  AND U22437 ( .A(n1108), .B(n22679), .Z(n22689) );
  XNOR U22438 ( .A(n22690), .B(n22677), .Z(n22679) );
  XOR U22439 ( .A(n22691), .B(n22692), .Z(n22677) );
  AND U22440 ( .A(n1131), .B(n22693), .Z(n22692) );
  IV U22441 ( .A(n22688), .Z(n22690) );
  XOR U22442 ( .A(n22694), .B(n22695), .Z(n22688) );
  AND U22443 ( .A(n1115), .B(n22687), .Z(n22695) );
  XNOR U22444 ( .A(n22685), .B(n22694), .Z(n22687) );
  XNOR U22445 ( .A(n22696), .B(n22697), .Z(n22685) );
  AND U22446 ( .A(n1119), .B(n22698), .Z(n22697) );
  XOR U22447 ( .A(p_input[1679]), .B(n22696), .Z(n22698) );
  XNOR U22448 ( .A(n22699), .B(n22700), .Z(n22696) );
  AND U22449 ( .A(n1123), .B(n22701), .Z(n22700) );
  XOR U22450 ( .A(n22702), .B(n22703), .Z(n22694) );
  AND U22451 ( .A(n1127), .B(n22693), .Z(n22703) );
  XNOR U22452 ( .A(n22704), .B(n22691), .Z(n22693) );
  XOR U22453 ( .A(n22705), .B(n22706), .Z(n22691) );
  AND U22454 ( .A(n1150), .B(n22707), .Z(n22706) );
  IV U22455 ( .A(n22702), .Z(n22704) );
  XOR U22456 ( .A(n22708), .B(n22709), .Z(n22702) );
  AND U22457 ( .A(n1134), .B(n22701), .Z(n22709) );
  XNOR U22458 ( .A(n22699), .B(n22708), .Z(n22701) );
  XNOR U22459 ( .A(n22710), .B(n22711), .Z(n22699) );
  AND U22460 ( .A(n1138), .B(n22712), .Z(n22711) );
  XOR U22461 ( .A(p_input[1711]), .B(n22710), .Z(n22712) );
  XNOR U22462 ( .A(n22713), .B(n22714), .Z(n22710) );
  AND U22463 ( .A(n1142), .B(n22715), .Z(n22714) );
  XOR U22464 ( .A(n22716), .B(n22717), .Z(n22708) );
  AND U22465 ( .A(n1146), .B(n22707), .Z(n22717) );
  XNOR U22466 ( .A(n22718), .B(n22705), .Z(n22707) );
  XOR U22467 ( .A(n22719), .B(n22720), .Z(n22705) );
  AND U22468 ( .A(n1169), .B(n22721), .Z(n22720) );
  IV U22469 ( .A(n22716), .Z(n22718) );
  XOR U22470 ( .A(n22722), .B(n22723), .Z(n22716) );
  AND U22471 ( .A(n1153), .B(n22715), .Z(n22723) );
  XNOR U22472 ( .A(n22713), .B(n22722), .Z(n22715) );
  XNOR U22473 ( .A(n22724), .B(n22725), .Z(n22713) );
  AND U22474 ( .A(n1157), .B(n22726), .Z(n22725) );
  XOR U22475 ( .A(p_input[1743]), .B(n22724), .Z(n22726) );
  XNOR U22476 ( .A(n22727), .B(n22728), .Z(n22724) );
  AND U22477 ( .A(n1161), .B(n22729), .Z(n22728) );
  XOR U22478 ( .A(n22730), .B(n22731), .Z(n22722) );
  AND U22479 ( .A(n1165), .B(n22721), .Z(n22731) );
  XNOR U22480 ( .A(n22732), .B(n22719), .Z(n22721) );
  XOR U22481 ( .A(n22733), .B(n22734), .Z(n22719) );
  AND U22482 ( .A(n1188), .B(n22735), .Z(n22734) );
  IV U22483 ( .A(n22730), .Z(n22732) );
  XOR U22484 ( .A(n22736), .B(n22737), .Z(n22730) );
  AND U22485 ( .A(n1172), .B(n22729), .Z(n22737) );
  XNOR U22486 ( .A(n22727), .B(n22736), .Z(n22729) );
  XNOR U22487 ( .A(n22738), .B(n22739), .Z(n22727) );
  AND U22488 ( .A(n1176), .B(n22740), .Z(n22739) );
  XOR U22489 ( .A(p_input[1775]), .B(n22738), .Z(n22740) );
  XNOR U22490 ( .A(n22741), .B(n22742), .Z(n22738) );
  AND U22491 ( .A(n1180), .B(n22743), .Z(n22742) );
  XOR U22492 ( .A(n22744), .B(n22745), .Z(n22736) );
  AND U22493 ( .A(n1184), .B(n22735), .Z(n22745) );
  XNOR U22494 ( .A(n22746), .B(n22733), .Z(n22735) );
  XOR U22495 ( .A(n22747), .B(n22748), .Z(n22733) );
  AND U22496 ( .A(n1207), .B(n22749), .Z(n22748) );
  IV U22497 ( .A(n22744), .Z(n22746) );
  XOR U22498 ( .A(n22750), .B(n22751), .Z(n22744) );
  AND U22499 ( .A(n1191), .B(n22743), .Z(n22751) );
  XNOR U22500 ( .A(n22741), .B(n22750), .Z(n22743) );
  XNOR U22501 ( .A(n22752), .B(n22753), .Z(n22741) );
  AND U22502 ( .A(n1195), .B(n22754), .Z(n22753) );
  XOR U22503 ( .A(p_input[1807]), .B(n22752), .Z(n22754) );
  XNOR U22504 ( .A(n22755), .B(n22756), .Z(n22752) );
  AND U22505 ( .A(n1199), .B(n22757), .Z(n22756) );
  XOR U22506 ( .A(n22758), .B(n22759), .Z(n22750) );
  AND U22507 ( .A(n1203), .B(n22749), .Z(n22759) );
  XNOR U22508 ( .A(n22760), .B(n22747), .Z(n22749) );
  XOR U22509 ( .A(n22761), .B(n22762), .Z(n22747) );
  AND U22510 ( .A(n1226), .B(n22763), .Z(n22762) );
  IV U22511 ( .A(n22758), .Z(n22760) );
  XOR U22512 ( .A(n22764), .B(n22765), .Z(n22758) );
  AND U22513 ( .A(n1210), .B(n22757), .Z(n22765) );
  XNOR U22514 ( .A(n22755), .B(n22764), .Z(n22757) );
  XNOR U22515 ( .A(n22766), .B(n22767), .Z(n22755) );
  AND U22516 ( .A(n1214), .B(n22768), .Z(n22767) );
  XOR U22517 ( .A(p_input[1839]), .B(n22766), .Z(n22768) );
  XNOR U22518 ( .A(n22769), .B(n22770), .Z(n22766) );
  AND U22519 ( .A(n1218), .B(n22771), .Z(n22770) );
  XOR U22520 ( .A(n22772), .B(n22773), .Z(n22764) );
  AND U22521 ( .A(n1222), .B(n22763), .Z(n22773) );
  XNOR U22522 ( .A(n22774), .B(n22761), .Z(n22763) );
  XOR U22523 ( .A(n22775), .B(n22776), .Z(n22761) );
  AND U22524 ( .A(n1245), .B(n22777), .Z(n22776) );
  IV U22525 ( .A(n22772), .Z(n22774) );
  XOR U22526 ( .A(n22778), .B(n22779), .Z(n22772) );
  AND U22527 ( .A(n1229), .B(n22771), .Z(n22779) );
  XNOR U22528 ( .A(n22769), .B(n22778), .Z(n22771) );
  XNOR U22529 ( .A(n22780), .B(n22781), .Z(n22769) );
  AND U22530 ( .A(n1233), .B(n22782), .Z(n22781) );
  XOR U22531 ( .A(p_input[1871]), .B(n22780), .Z(n22782) );
  XNOR U22532 ( .A(n22783), .B(n22784), .Z(n22780) );
  AND U22533 ( .A(n1237), .B(n22785), .Z(n22784) );
  XOR U22534 ( .A(n22786), .B(n22787), .Z(n22778) );
  AND U22535 ( .A(n1241), .B(n22777), .Z(n22787) );
  XNOR U22536 ( .A(n22788), .B(n22775), .Z(n22777) );
  XOR U22537 ( .A(n22789), .B(n22790), .Z(n22775) );
  AND U22538 ( .A(n1264), .B(n22791), .Z(n22790) );
  IV U22539 ( .A(n22786), .Z(n22788) );
  XOR U22540 ( .A(n22792), .B(n22793), .Z(n22786) );
  AND U22541 ( .A(n1248), .B(n22785), .Z(n22793) );
  XNOR U22542 ( .A(n22783), .B(n22792), .Z(n22785) );
  XNOR U22543 ( .A(n22794), .B(n22795), .Z(n22783) );
  AND U22544 ( .A(n1252), .B(n22796), .Z(n22795) );
  XOR U22545 ( .A(p_input[1903]), .B(n22794), .Z(n22796) );
  XNOR U22546 ( .A(n22797), .B(n22798), .Z(n22794) );
  AND U22547 ( .A(n1256), .B(n22799), .Z(n22798) );
  XOR U22548 ( .A(n22800), .B(n22801), .Z(n22792) );
  AND U22549 ( .A(n1260), .B(n22791), .Z(n22801) );
  XNOR U22550 ( .A(n22802), .B(n22789), .Z(n22791) );
  XOR U22551 ( .A(n22803), .B(n22804), .Z(n22789) );
  AND U22552 ( .A(n1282), .B(n22805), .Z(n22804) );
  IV U22553 ( .A(n22800), .Z(n22802) );
  XOR U22554 ( .A(n22806), .B(n22807), .Z(n22800) );
  AND U22555 ( .A(n1267), .B(n22799), .Z(n22807) );
  XNOR U22556 ( .A(n22797), .B(n22806), .Z(n22799) );
  XNOR U22557 ( .A(n22808), .B(n22809), .Z(n22797) );
  AND U22558 ( .A(n1271), .B(n22810), .Z(n22809) );
  XOR U22559 ( .A(p_input[1935]), .B(n22808), .Z(n22810) );
  XOR U22560 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n22811), 
        .Z(n22808) );
  AND U22561 ( .A(n1274), .B(n22812), .Z(n22811) );
  XOR U22562 ( .A(n22813), .B(n22814), .Z(n22806) );
  AND U22563 ( .A(n1278), .B(n22805), .Z(n22814) );
  XNOR U22564 ( .A(n22815), .B(n22803), .Z(n22805) );
  XOR U22565 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n22816), .Z(n22803) );
  AND U22566 ( .A(n1290), .B(n22817), .Z(n22816) );
  IV U22567 ( .A(n22813), .Z(n22815) );
  XOR U22568 ( .A(n22818), .B(n22819), .Z(n22813) );
  AND U22569 ( .A(n1285), .B(n22812), .Z(n22819) );
  XOR U22570 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n22818), 
        .Z(n22812) );
  XOR U22571 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(n22820), 
        .Z(n22818) );
  AND U22572 ( .A(n1287), .B(n22817), .Z(n22820) );
  XOR U22573 ( .A(n22821), .B(n22822), .Z(n22817) );
  IV U22574 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .Z(n22822)
         );
  IV U22575 ( .A(\knn_comb_/min_val_out[0][15] ), .Z(n22821) );
  XOR U22576 ( .A(n111), .B(n22823), .Z(o[14]) );
  AND U22577 ( .A(n122), .B(n22824), .Z(n111) );
  XOR U22578 ( .A(n112), .B(n22823), .Z(n22824) );
  XOR U22579 ( .A(n22825), .B(n22826), .Z(n22823) );
  AND U22580 ( .A(n142), .B(n22827), .Z(n22826) );
  XOR U22581 ( .A(n22828), .B(n41), .Z(n112) );
  AND U22582 ( .A(n125), .B(n22829), .Z(n41) );
  XOR U22583 ( .A(n42), .B(n22828), .Z(n22829) );
  XOR U22584 ( .A(n22830), .B(n22831), .Z(n42) );
  AND U22585 ( .A(n130), .B(n22832), .Z(n22831) );
  XOR U22586 ( .A(p_input[14]), .B(n22830), .Z(n22832) );
  XNOR U22587 ( .A(n22833), .B(n22834), .Z(n22830) );
  AND U22588 ( .A(n134), .B(n22835), .Z(n22834) );
  XOR U22589 ( .A(n22836), .B(n22837), .Z(n22828) );
  AND U22590 ( .A(n138), .B(n22827), .Z(n22837) );
  XNOR U22591 ( .A(n22838), .B(n22825), .Z(n22827) );
  XOR U22592 ( .A(n22839), .B(n22840), .Z(n22825) );
  AND U22593 ( .A(n162), .B(n22841), .Z(n22840) );
  IV U22594 ( .A(n22836), .Z(n22838) );
  XOR U22595 ( .A(n22842), .B(n22843), .Z(n22836) );
  AND U22596 ( .A(n146), .B(n22835), .Z(n22843) );
  XNOR U22597 ( .A(n22833), .B(n22842), .Z(n22835) );
  XNOR U22598 ( .A(n22844), .B(n22845), .Z(n22833) );
  AND U22599 ( .A(n150), .B(n22846), .Z(n22845) );
  XOR U22600 ( .A(p_input[46]), .B(n22844), .Z(n22846) );
  XNOR U22601 ( .A(n22847), .B(n22848), .Z(n22844) );
  AND U22602 ( .A(n154), .B(n22849), .Z(n22848) );
  XOR U22603 ( .A(n22850), .B(n22851), .Z(n22842) );
  AND U22604 ( .A(n158), .B(n22841), .Z(n22851) );
  XNOR U22605 ( .A(n22852), .B(n22839), .Z(n22841) );
  XOR U22606 ( .A(n22853), .B(n22854), .Z(n22839) );
  AND U22607 ( .A(n181), .B(n22855), .Z(n22854) );
  IV U22608 ( .A(n22850), .Z(n22852) );
  XOR U22609 ( .A(n22856), .B(n22857), .Z(n22850) );
  AND U22610 ( .A(n165), .B(n22849), .Z(n22857) );
  XNOR U22611 ( .A(n22847), .B(n22856), .Z(n22849) );
  XNOR U22612 ( .A(n22858), .B(n22859), .Z(n22847) );
  AND U22613 ( .A(n169), .B(n22860), .Z(n22859) );
  XOR U22614 ( .A(p_input[78]), .B(n22858), .Z(n22860) );
  XNOR U22615 ( .A(n22861), .B(n22862), .Z(n22858) );
  AND U22616 ( .A(n173), .B(n22863), .Z(n22862) );
  XOR U22617 ( .A(n22864), .B(n22865), .Z(n22856) );
  AND U22618 ( .A(n177), .B(n22855), .Z(n22865) );
  XNOR U22619 ( .A(n22866), .B(n22853), .Z(n22855) );
  XOR U22620 ( .A(n22867), .B(n22868), .Z(n22853) );
  AND U22621 ( .A(n200), .B(n22869), .Z(n22868) );
  IV U22622 ( .A(n22864), .Z(n22866) );
  XOR U22623 ( .A(n22870), .B(n22871), .Z(n22864) );
  AND U22624 ( .A(n184), .B(n22863), .Z(n22871) );
  XNOR U22625 ( .A(n22861), .B(n22870), .Z(n22863) );
  XNOR U22626 ( .A(n22872), .B(n22873), .Z(n22861) );
  AND U22627 ( .A(n188), .B(n22874), .Z(n22873) );
  XOR U22628 ( .A(p_input[110]), .B(n22872), .Z(n22874) );
  XNOR U22629 ( .A(n22875), .B(n22876), .Z(n22872) );
  AND U22630 ( .A(n192), .B(n22877), .Z(n22876) );
  XOR U22631 ( .A(n22878), .B(n22879), .Z(n22870) );
  AND U22632 ( .A(n196), .B(n22869), .Z(n22879) );
  XNOR U22633 ( .A(n22880), .B(n22867), .Z(n22869) );
  XOR U22634 ( .A(n22881), .B(n22882), .Z(n22867) );
  AND U22635 ( .A(n219), .B(n22883), .Z(n22882) );
  IV U22636 ( .A(n22878), .Z(n22880) );
  XOR U22637 ( .A(n22884), .B(n22885), .Z(n22878) );
  AND U22638 ( .A(n203), .B(n22877), .Z(n22885) );
  XNOR U22639 ( .A(n22875), .B(n22884), .Z(n22877) );
  XNOR U22640 ( .A(n22886), .B(n22887), .Z(n22875) );
  AND U22641 ( .A(n207), .B(n22888), .Z(n22887) );
  XOR U22642 ( .A(p_input[142]), .B(n22886), .Z(n22888) );
  XNOR U22643 ( .A(n22889), .B(n22890), .Z(n22886) );
  AND U22644 ( .A(n211), .B(n22891), .Z(n22890) );
  XOR U22645 ( .A(n22892), .B(n22893), .Z(n22884) );
  AND U22646 ( .A(n215), .B(n22883), .Z(n22893) );
  XNOR U22647 ( .A(n22894), .B(n22881), .Z(n22883) );
  XOR U22648 ( .A(n22895), .B(n22896), .Z(n22881) );
  AND U22649 ( .A(n238), .B(n22897), .Z(n22896) );
  IV U22650 ( .A(n22892), .Z(n22894) );
  XOR U22651 ( .A(n22898), .B(n22899), .Z(n22892) );
  AND U22652 ( .A(n222), .B(n22891), .Z(n22899) );
  XNOR U22653 ( .A(n22889), .B(n22898), .Z(n22891) );
  XNOR U22654 ( .A(n22900), .B(n22901), .Z(n22889) );
  AND U22655 ( .A(n226), .B(n22902), .Z(n22901) );
  XOR U22656 ( .A(p_input[174]), .B(n22900), .Z(n22902) );
  XNOR U22657 ( .A(n22903), .B(n22904), .Z(n22900) );
  AND U22658 ( .A(n230), .B(n22905), .Z(n22904) );
  XOR U22659 ( .A(n22906), .B(n22907), .Z(n22898) );
  AND U22660 ( .A(n234), .B(n22897), .Z(n22907) );
  XNOR U22661 ( .A(n22908), .B(n22895), .Z(n22897) );
  XOR U22662 ( .A(n22909), .B(n22910), .Z(n22895) );
  AND U22663 ( .A(n257), .B(n22911), .Z(n22910) );
  IV U22664 ( .A(n22906), .Z(n22908) );
  XOR U22665 ( .A(n22912), .B(n22913), .Z(n22906) );
  AND U22666 ( .A(n241), .B(n22905), .Z(n22913) );
  XNOR U22667 ( .A(n22903), .B(n22912), .Z(n22905) );
  XNOR U22668 ( .A(n22914), .B(n22915), .Z(n22903) );
  AND U22669 ( .A(n245), .B(n22916), .Z(n22915) );
  XOR U22670 ( .A(p_input[206]), .B(n22914), .Z(n22916) );
  XNOR U22671 ( .A(n22917), .B(n22918), .Z(n22914) );
  AND U22672 ( .A(n249), .B(n22919), .Z(n22918) );
  XOR U22673 ( .A(n22920), .B(n22921), .Z(n22912) );
  AND U22674 ( .A(n253), .B(n22911), .Z(n22921) );
  XNOR U22675 ( .A(n22922), .B(n22909), .Z(n22911) );
  XOR U22676 ( .A(n22923), .B(n22924), .Z(n22909) );
  AND U22677 ( .A(n276), .B(n22925), .Z(n22924) );
  IV U22678 ( .A(n22920), .Z(n22922) );
  XOR U22679 ( .A(n22926), .B(n22927), .Z(n22920) );
  AND U22680 ( .A(n260), .B(n22919), .Z(n22927) );
  XNOR U22681 ( .A(n22917), .B(n22926), .Z(n22919) );
  XNOR U22682 ( .A(n22928), .B(n22929), .Z(n22917) );
  AND U22683 ( .A(n264), .B(n22930), .Z(n22929) );
  XOR U22684 ( .A(p_input[238]), .B(n22928), .Z(n22930) );
  XNOR U22685 ( .A(n22931), .B(n22932), .Z(n22928) );
  AND U22686 ( .A(n268), .B(n22933), .Z(n22932) );
  XOR U22687 ( .A(n22934), .B(n22935), .Z(n22926) );
  AND U22688 ( .A(n272), .B(n22925), .Z(n22935) );
  XNOR U22689 ( .A(n22936), .B(n22923), .Z(n22925) );
  XOR U22690 ( .A(n22937), .B(n22938), .Z(n22923) );
  AND U22691 ( .A(n295), .B(n22939), .Z(n22938) );
  IV U22692 ( .A(n22934), .Z(n22936) );
  XOR U22693 ( .A(n22940), .B(n22941), .Z(n22934) );
  AND U22694 ( .A(n279), .B(n22933), .Z(n22941) );
  XNOR U22695 ( .A(n22931), .B(n22940), .Z(n22933) );
  XNOR U22696 ( .A(n22942), .B(n22943), .Z(n22931) );
  AND U22697 ( .A(n283), .B(n22944), .Z(n22943) );
  XOR U22698 ( .A(p_input[270]), .B(n22942), .Z(n22944) );
  XNOR U22699 ( .A(n22945), .B(n22946), .Z(n22942) );
  AND U22700 ( .A(n287), .B(n22947), .Z(n22946) );
  XOR U22701 ( .A(n22948), .B(n22949), .Z(n22940) );
  AND U22702 ( .A(n291), .B(n22939), .Z(n22949) );
  XNOR U22703 ( .A(n22950), .B(n22937), .Z(n22939) );
  XOR U22704 ( .A(n22951), .B(n22952), .Z(n22937) );
  AND U22705 ( .A(n314), .B(n22953), .Z(n22952) );
  IV U22706 ( .A(n22948), .Z(n22950) );
  XOR U22707 ( .A(n22954), .B(n22955), .Z(n22948) );
  AND U22708 ( .A(n298), .B(n22947), .Z(n22955) );
  XNOR U22709 ( .A(n22945), .B(n22954), .Z(n22947) );
  XNOR U22710 ( .A(n22956), .B(n22957), .Z(n22945) );
  AND U22711 ( .A(n302), .B(n22958), .Z(n22957) );
  XOR U22712 ( .A(p_input[302]), .B(n22956), .Z(n22958) );
  XNOR U22713 ( .A(n22959), .B(n22960), .Z(n22956) );
  AND U22714 ( .A(n306), .B(n22961), .Z(n22960) );
  XOR U22715 ( .A(n22962), .B(n22963), .Z(n22954) );
  AND U22716 ( .A(n310), .B(n22953), .Z(n22963) );
  XNOR U22717 ( .A(n22964), .B(n22951), .Z(n22953) );
  XOR U22718 ( .A(n22965), .B(n22966), .Z(n22951) );
  AND U22719 ( .A(n333), .B(n22967), .Z(n22966) );
  IV U22720 ( .A(n22962), .Z(n22964) );
  XOR U22721 ( .A(n22968), .B(n22969), .Z(n22962) );
  AND U22722 ( .A(n317), .B(n22961), .Z(n22969) );
  XNOR U22723 ( .A(n22959), .B(n22968), .Z(n22961) );
  XNOR U22724 ( .A(n22970), .B(n22971), .Z(n22959) );
  AND U22725 ( .A(n321), .B(n22972), .Z(n22971) );
  XOR U22726 ( .A(p_input[334]), .B(n22970), .Z(n22972) );
  XNOR U22727 ( .A(n22973), .B(n22974), .Z(n22970) );
  AND U22728 ( .A(n325), .B(n22975), .Z(n22974) );
  XOR U22729 ( .A(n22976), .B(n22977), .Z(n22968) );
  AND U22730 ( .A(n329), .B(n22967), .Z(n22977) );
  XNOR U22731 ( .A(n22978), .B(n22965), .Z(n22967) );
  XOR U22732 ( .A(n22979), .B(n22980), .Z(n22965) );
  AND U22733 ( .A(n352), .B(n22981), .Z(n22980) );
  IV U22734 ( .A(n22976), .Z(n22978) );
  XOR U22735 ( .A(n22982), .B(n22983), .Z(n22976) );
  AND U22736 ( .A(n336), .B(n22975), .Z(n22983) );
  XNOR U22737 ( .A(n22973), .B(n22982), .Z(n22975) );
  XNOR U22738 ( .A(n22984), .B(n22985), .Z(n22973) );
  AND U22739 ( .A(n340), .B(n22986), .Z(n22985) );
  XOR U22740 ( .A(p_input[366]), .B(n22984), .Z(n22986) );
  XNOR U22741 ( .A(n22987), .B(n22988), .Z(n22984) );
  AND U22742 ( .A(n344), .B(n22989), .Z(n22988) );
  XOR U22743 ( .A(n22990), .B(n22991), .Z(n22982) );
  AND U22744 ( .A(n348), .B(n22981), .Z(n22991) );
  XNOR U22745 ( .A(n22992), .B(n22979), .Z(n22981) );
  XOR U22746 ( .A(n22993), .B(n22994), .Z(n22979) );
  AND U22747 ( .A(n371), .B(n22995), .Z(n22994) );
  IV U22748 ( .A(n22990), .Z(n22992) );
  XOR U22749 ( .A(n22996), .B(n22997), .Z(n22990) );
  AND U22750 ( .A(n355), .B(n22989), .Z(n22997) );
  XNOR U22751 ( .A(n22987), .B(n22996), .Z(n22989) );
  XNOR U22752 ( .A(n22998), .B(n22999), .Z(n22987) );
  AND U22753 ( .A(n359), .B(n23000), .Z(n22999) );
  XOR U22754 ( .A(p_input[398]), .B(n22998), .Z(n23000) );
  XNOR U22755 ( .A(n23001), .B(n23002), .Z(n22998) );
  AND U22756 ( .A(n363), .B(n23003), .Z(n23002) );
  XOR U22757 ( .A(n23004), .B(n23005), .Z(n22996) );
  AND U22758 ( .A(n367), .B(n22995), .Z(n23005) );
  XNOR U22759 ( .A(n23006), .B(n22993), .Z(n22995) );
  XOR U22760 ( .A(n23007), .B(n23008), .Z(n22993) );
  AND U22761 ( .A(n390), .B(n23009), .Z(n23008) );
  IV U22762 ( .A(n23004), .Z(n23006) );
  XOR U22763 ( .A(n23010), .B(n23011), .Z(n23004) );
  AND U22764 ( .A(n374), .B(n23003), .Z(n23011) );
  XNOR U22765 ( .A(n23001), .B(n23010), .Z(n23003) );
  XNOR U22766 ( .A(n23012), .B(n23013), .Z(n23001) );
  AND U22767 ( .A(n378), .B(n23014), .Z(n23013) );
  XOR U22768 ( .A(p_input[430]), .B(n23012), .Z(n23014) );
  XNOR U22769 ( .A(n23015), .B(n23016), .Z(n23012) );
  AND U22770 ( .A(n382), .B(n23017), .Z(n23016) );
  XOR U22771 ( .A(n23018), .B(n23019), .Z(n23010) );
  AND U22772 ( .A(n386), .B(n23009), .Z(n23019) );
  XNOR U22773 ( .A(n23020), .B(n23007), .Z(n23009) );
  XOR U22774 ( .A(n23021), .B(n23022), .Z(n23007) );
  AND U22775 ( .A(n409), .B(n23023), .Z(n23022) );
  IV U22776 ( .A(n23018), .Z(n23020) );
  XOR U22777 ( .A(n23024), .B(n23025), .Z(n23018) );
  AND U22778 ( .A(n393), .B(n23017), .Z(n23025) );
  XNOR U22779 ( .A(n23015), .B(n23024), .Z(n23017) );
  XNOR U22780 ( .A(n23026), .B(n23027), .Z(n23015) );
  AND U22781 ( .A(n397), .B(n23028), .Z(n23027) );
  XOR U22782 ( .A(p_input[462]), .B(n23026), .Z(n23028) );
  XNOR U22783 ( .A(n23029), .B(n23030), .Z(n23026) );
  AND U22784 ( .A(n401), .B(n23031), .Z(n23030) );
  XOR U22785 ( .A(n23032), .B(n23033), .Z(n23024) );
  AND U22786 ( .A(n405), .B(n23023), .Z(n23033) );
  XNOR U22787 ( .A(n23034), .B(n23021), .Z(n23023) );
  XOR U22788 ( .A(n23035), .B(n23036), .Z(n23021) );
  AND U22789 ( .A(n428), .B(n23037), .Z(n23036) );
  IV U22790 ( .A(n23032), .Z(n23034) );
  XOR U22791 ( .A(n23038), .B(n23039), .Z(n23032) );
  AND U22792 ( .A(n412), .B(n23031), .Z(n23039) );
  XNOR U22793 ( .A(n23029), .B(n23038), .Z(n23031) );
  XNOR U22794 ( .A(n23040), .B(n23041), .Z(n23029) );
  AND U22795 ( .A(n416), .B(n23042), .Z(n23041) );
  XOR U22796 ( .A(p_input[494]), .B(n23040), .Z(n23042) );
  XNOR U22797 ( .A(n23043), .B(n23044), .Z(n23040) );
  AND U22798 ( .A(n420), .B(n23045), .Z(n23044) );
  XOR U22799 ( .A(n23046), .B(n23047), .Z(n23038) );
  AND U22800 ( .A(n424), .B(n23037), .Z(n23047) );
  XNOR U22801 ( .A(n23048), .B(n23035), .Z(n23037) );
  XOR U22802 ( .A(n23049), .B(n23050), .Z(n23035) );
  AND U22803 ( .A(n447), .B(n23051), .Z(n23050) );
  IV U22804 ( .A(n23046), .Z(n23048) );
  XOR U22805 ( .A(n23052), .B(n23053), .Z(n23046) );
  AND U22806 ( .A(n431), .B(n23045), .Z(n23053) );
  XNOR U22807 ( .A(n23043), .B(n23052), .Z(n23045) );
  XNOR U22808 ( .A(n23054), .B(n23055), .Z(n23043) );
  AND U22809 ( .A(n435), .B(n23056), .Z(n23055) );
  XOR U22810 ( .A(p_input[526]), .B(n23054), .Z(n23056) );
  XNOR U22811 ( .A(n23057), .B(n23058), .Z(n23054) );
  AND U22812 ( .A(n439), .B(n23059), .Z(n23058) );
  XOR U22813 ( .A(n23060), .B(n23061), .Z(n23052) );
  AND U22814 ( .A(n443), .B(n23051), .Z(n23061) );
  XNOR U22815 ( .A(n23062), .B(n23049), .Z(n23051) );
  XOR U22816 ( .A(n23063), .B(n23064), .Z(n23049) );
  AND U22817 ( .A(n466), .B(n23065), .Z(n23064) );
  IV U22818 ( .A(n23060), .Z(n23062) );
  XOR U22819 ( .A(n23066), .B(n23067), .Z(n23060) );
  AND U22820 ( .A(n450), .B(n23059), .Z(n23067) );
  XNOR U22821 ( .A(n23057), .B(n23066), .Z(n23059) );
  XNOR U22822 ( .A(n23068), .B(n23069), .Z(n23057) );
  AND U22823 ( .A(n454), .B(n23070), .Z(n23069) );
  XOR U22824 ( .A(p_input[558]), .B(n23068), .Z(n23070) );
  XNOR U22825 ( .A(n23071), .B(n23072), .Z(n23068) );
  AND U22826 ( .A(n458), .B(n23073), .Z(n23072) );
  XOR U22827 ( .A(n23074), .B(n23075), .Z(n23066) );
  AND U22828 ( .A(n462), .B(n23065), .Z(n23075) );
  XNOR U22829 ( .A(n23076), .B(n23063), .Z(n23065) );
  XOR U22830 ( .A(n23077), .B(n23078), .Z(n23063) );
  AND U22831 ( .A(n485), .B(n23079), .Z(n23078) );
  IV U22832 ( .A(n23074), .Z(n23076) );
  XOR U22833 ( .A(n23080), .B(n23081), .Z(n23074) );
  AND U22834 ( .A(n469), .B(n23073), .Z(n23081) );
  XNOR U22835 ( .A(n23071), .B(n23080), .Z(n23073) );
  XNOR U22836 ( .A(n23082), .B(n23083), .Z(n23071) );
  AND U22837 ( .A(n473), .B(n23084), .Z(n23083) );
  XOR U22838 ( .A(p_input[590]), .B(n23082), .Z(n23084) );
  XNOR U22839 ( .A(n23085), .B(n23086), .Z(n23082) );
  AND U22840 ( .A(n477), .B(n23087), .Z(n23086) );
  XOR U22841 ( .A(n23088), .B(n23089), .Z(n23080) );
  AND U22842 ( .A(n481), .B(n23079), .Z(n23089) );
  XNOR U22843 ( .A(n23090), .B(n23077), .Z(n23079) );
  XOR U22844 ( .A(n23091), .B(n23092), .Z(n23077) );
  AND U22845 ( .A(n504), .B(n23093), .Z(n23092) );
  IV U22846 ( .A(n23088), .Z(n23090) );
  XOR U22847 ( .A(n23094), .B(n23095), .Z(n23088) );
  AND U22848 ( .A(n488), .B(n23087), .Z(n23095) );
  XNOR U22849 ( .A(n23085), .B(n23094), .Z(n23087) );
  XNOR U22850 ( .A(n23096), .B(n23097), .Z(n23085) );
  AND U22851 ( .A(n492), .B(n23098), .Z(n23097) );
  XOR U22852 ( .A(p_input[622]), .B(n23096), .Z(n23098) );
  XNOR U22853 ( .A(n23099), .B(n23100), .Z(n23096) );
  AND U22854 ( .A(n496), .B(n23101), .Z(n23100) );
  XOR U22855 ( .A(n23102), .B(n23103), .Z(n23094) );
  AND U22856 ( .A(n500), .B(n23093), .Z(n23103) );
  XNOR U22857 ( .A(n23104), .B(n23091), .Z(n23093) );
  XOR U22858 ( .A(n23105), .B(n23106), .Z(n23091) );
  AND U22859 ( .A(n523), .B(n23107), .Z(n23106) );
  IV U22860 ( .A(n23102), .Z(n23104) );
  XOR U22861 ( .A(n23108), .B(n23109), .Z(n23102) );
  AND U22862 ( .A(n507), .B(n23101), .Z(n23109) );
  XNOR U22863 ( .A(n23099), .B(n23108), .Z(n23101) );
  XNOR U22864 ( .A(n23110), .B(n23111), .Z(n23099) );
  AND U22865 ( .A(n511), .B(n23112), .Z(n23111) );
  XOR U22866 ( .A(p_input[654]), .B(n23110), .Z(n23112) );
  XNOR U22867 ( .A(n23113), .B(n23114), .Z(n23110) );
  AND U22868 ( .A(n515), .B(n23115), .Z(n23114) );
  XOR U22869 ( .A(n23116), .B(n23117), .Z(n23108) );
  AND U22870 ( .A(n519), .B(n23107), .Z(n23117) );
  XNOR U22871 ( .A(n23118), .B(n23105), .Z(n23107) );
  XOR U22872 ( .A(n23119), .B(n23120), .Z(n23105) );
  AND U22873 ( .A(n542), .B(n23121), .Z(n23120) );
  IV U22874 ( .A(n23116), .Z(n23118) );
  XOR U22875 ( .A(n23122), .B(n23123), .Z(n23116) );
  AND U22876 ( .A(n526), .B(n23115), .Z(n23123) );
  XNOR U22877 ( .A(n23113), .B(n23122), .Z(n23115) );
  XNOR U22878 ( .A(n23124), .B(n23125), .Z(n23113) );
  AND U22879 ( .A(n530), .B(n23126), .Z(n23125) );
  XOR U22880 ( .A(p_input[686]), .B(n23124), .Z(n23126) );
  XNOR U22881 ( .A(n23127), .B(n23128), .Z(n23124) );
  AND U22882 ( .A(n534), .B(n23129), .Z(n23128) );
  XOR U22883 ( .A(n23130), .B(n23131), .Z(n23122) );
  AND U22884 ( .A(n538), .B(n23121), .Z(n23131) );
  XNOR U22885 ( .A(n23132), .B(n23119), .Z(n23121) );
  XOR U22886 ( .A(n23133), .B(n23134), .Z(n23119) );
  AND U22887 ( .A(n561), .B(n23135), .Z(n23134) );
  IV U22888 ( .A(n23130), .Z(n23132) );
  XOR U22889 ( .A(n23136), .B(n23137), .Z(n23130) );
  AND U22890 ( .A(n545), .B(n23129), .Z(n23137) );
  XNOR U22891 ( .A(n23127), .B(n23136), .Z(n23129) );
  XNOR U22892 ( .A(n23138), .B(n23139), .Z(n23127) );
  AND U22893 ( .A(n549), .B(n23140), .Z(n23139) );
  XOR U22894 ( .A(p_input[718]), .B(n23138), .Z(n23140) );
  XNOR U22895 ( .A(n23141), .B(n23142), .Z(n23138) );
  AND U22896 ( .A(n553), .B(n23143), .Z(n23142) );
  XOR U22897 ( .A(n23144), .B(n23145), .Z(n23136) );
  AND U22898 ( .A(n557), .B(n23135), .Z(n23145) );
  XNOR U22899 ( .A(n23146), .B(n23133), .Z(n23135) );
  XOR U22900 ( .A(n23147), .B(n23148), .Z(n23133) );
  AND U22901 ( .A(n580), .B(n23149), .Z(n23148) );
  IV U22902 ( .A(n23144), .Z(n23146) );
  XOR U22903 ( .A(n23150), .B(n23151), .Z(n23144) );
  AND U22904 ( .A(n564), .B(n23143), .Z(n23151) );
  XNOR U22905 ( .A(n23141), .B(n23150), .Z(n23143) );
  XNOR U22906 ( .A(n23152), .B(n23153), .Z(n23141) );
  AND U22907 ( .A(n568), .B(n23154), .Z(n23153) );
  XOR U22908 ( .A(p_input[750]), .B(n23152), .Z(n23154) );
  XNOR U22909 ( .A(n23155), .B(n23156), .Z(n23152) );
  AND U22910 ( .A(n572), .B(n23157), .Z(n23156) );
  XOR U22911 ( .A(n23158), .B(n23159), .Z(n23150) );
  AND U22912 ( .A(n576), .B(n23149), .Z(n23159) );
  XNOR U22913 ( .A(n23160), .B(n23147), .Z(n23149) );
  XOR U22914 ( .A(n23161), .B(n23162), .Z(n23147) );
  AND U22915 ( .A(n599), .B(n23163), .Z(n23162) );
  IV U22916 ( .A(n23158), .Z(n23160) );
  XOR U22917 ( .A(n23164), .B(n23165), .Z(n23158) );
  AND U22918 ( .A(n583), .B(n23157), .Z(n23165) );
  XNOR U22919 ( .A(n23155), .B(n23164), .Z(n23157) );
  XNOR U22920 ( .A(n23166), .B(n23167), .Z(n23155) );
  AND U22921 ( .A(n587), .B(n23168), .Z(n23167) );
  XOR U22922 ( .A(p_input[782]), .B(n23166), .Z(n23168) );
  XNOR U22923 ( .A(n23169), .B(n23170), .Z(n23166) );
  AND U22924 ( .A(n591), .B(n23171), .Z(n23170) );
  XOR U22925 ( .A(n23172), .B(n23173), .Z(n23164) );
  AND U22926 ( .A(n595), .B(n23163), .Z(n23173) );
  XNOR U22927 ( .A(n23174), .B(n23161), .Z(n23163) );
  XOR U22928 ( .A(n23175), .B(n23176), .Z(n23161) );
  AND U22929 ( .A(n618), .B(n23177), .Z(n23176) );
  IV U22930 ( .A(n23172), .Z(n23174) );
  XOR U22931 ( .A(n23178), .B(n23179), .Z(n23172) );
  AND U22932 ( .A(n602), .B(n23171), .Z(n23179) );
  XNOR U22933 ( .A(n23169), .B(n23178), .Z(n23171) );
  XNOR U22934 ( .A(n23180), .B(n23181), .Z(n23169) );
  AND U22935 ( .A(n606), .B(n23182), .Z(n23181) );
  XOR U22936 ( .A(p_input[814]), .B(n23180), .Z(n23182) );
  XNOR U22937 ( .A(n23183), .B(n23184), .Z(n23180) );
  AND U22938 ( .A(n610), .B(n23185), .Z(n23184) );
  XOR U22939 ( .A(n23186), .B(n23187), .Z(n23178) );
  AND U22940 ( .A(n614), .B(n23177), .Z(n23187) );
  XNOR U22941 ( .A(n23188), .B(n23175), .Z(n23177) );
  XOR U22942 ( .A(n23189), .B(n23190), .Z(n23175) );
  AND U22943 ( .A(n637), .B(n23191), .Z(n23190) );
  IV U22944 ( .A(n23186), .Z(n23188) );
  XOR U22945 ( .A(n23192), .B(n23193), .Z(n23186) );
  AND U22946 ( .A(n621), .B(n23185), .Z(n23193) );
  XNOR U22947 ( .A(n23183), .B(n23192), .Z(n23185) );
  XNOR U22948 ( .A(n23194), .B(n23195), .Z(n23183) );
  AND U22949 ( .A(n625), .B(n23196), .Z(n23195) );
  XOR U22950 ( .A(p_input[846]), .B(n23194), .Z(n23196) );
  XNOR U22951 ( .A(n23197), .B(n23198), .Z(n23194) );
  AND U22952 ( .A(n629), .B(n23199), .Z(n23198) );
  XOR U22953 ( .A(n23200), .B(n23201), .Z(n23192) );
  AND U22954 ( .A(n633), .B(n23191), .Z(n23201) );
  XNOR U22955 ( .A(n23202), .B(n23189), .Z(n23191) );
  XOR U22956 ( .A(n23203), .B(n23204), .Z(n23189) );
  AND U22957 ( .A(n656), .B(n23205), .Z(n23204) );
  IV U22958 ( .A(n23200), .Z(n23202) );
  XOR U22959 ( .A(n23206), .B(n23207), .Z(n23200) );
  AND U22960 ( .A(n640), .B(n23199), .Z(n23207) );
  XNOR U22961 ( .A(n23197), .B(n23206), .Z(n23199) );
  XNOR U22962 ( .A(n23208), .B(n23209), .Z(n23197) );
  AND U22963 ( .A(n644), .B(n23210), .Z(n23209) );
  XOR U22964 ( .A(p_input[878]), .B(n23208), .Z(n23210) );
  XNOR U22965 ( .A(n23211), .B(n23212), .Z(n23208) );
  AND U22966 ( .A(n648), .B(n23213), .Z(n23212) );
  XOR U22967 ( .A(n23214), .B(n23215), .Z(n23206) );
  AND U22968 ( .A(n652), .B(n23205), .Z(n23215) );
  XNOR U22969 ( .A(n23216), .B(n23203), .Z(n23205) );
  XOR U22970 ( .A(n23217), .B(n23218), .Z(n23203) );
  AND U22971 ( .A(n675), .B(n23219), .Z(n23218) );
  IV U22972 ( .A(n23214), .Z(n23216) );
  XOR U22973 ( .A(n23220), .B(n23221), .Z(n23214) );
  AND U22974 ( .A(n659), .B(n23213), .Z(n23221) );
  XNOR U22975 ( .A(n23211), .B(n23220), .Z(n23213) );
  XNOR U22976 ( .A(n23222), .B(n23223), .Z(n23211) );
  AND U22977 ( .A(n663), .B(n23224), .Z(n23223) );
  XOR U22978 ( .A(p_input[910]), .B(n23222), .Z(n23224) );
  XNOR U22979 ( .A(n23225), .B(n23226), .Z(n23222) );
  AND U22980 ( .A(n667), .B(n23227), .Z(n23226) );
  XOR U22981 ( .A(n23228), .B(n23229), .Z(n23220) );
  AND U22982 ( .A(n671), .B(n23219), .Z(n23229) );
  XNOR U22983 ( .A(n23230), .B(n23217), .Z(n23219) );
  XOR U22984 ( .A(n23231), .B(n23232), .Z(n23217) );
  AND U22985 ( .A(n694), .B(n23233), .Z(n23232) );
  IV U22986 ( .A(n23228), .Z(n23230) );
  XOR U22987 ( .A(n23234), .B(n23235), .Z(n23228) );
  AND U22988 ( .A(n678), .B(n23227), .Z(n23235) );
  XNOR U22989 ( .A(n23225), .B(n23234), .Z(n23227) );
  XNOR U22990 ( .A(n23236), .B(n23237), .Z(n23225) );
  AND U22991 ( .A(n682), .B(n23238), .Z(n23237) );
  XOR U22992 ( .A(p_input[942]), .B(n23236), .Z(n23238) );
  XNOR U22993 ( .A(n23239), .B(n23240), .Z(n23236) );
  AND U22994 ( .A(n686), .B(n23241), .Z(n23240) );
  XOR U22995 ( .A(n23242), .B(n23243), .Z(n23234) );
  AND U22996 ( .A(n690), .B(n23233), .Z(n23243) );
  XNOR U22997 ( .A(n23244), .B(n23231), .Z(n23233) );
  XOR U22998 ( .A(n23245), .B(n23246), .Z(n23231) );
  AND U22999 ( .A(n713), .B(n23247), .Z(n23246) );
  IV U23000 ( .A(n23242), .Z(n23244) );
  XOR U23001 ( .A(n23248), .B(n23249), .Z(n23242) );
  AND U23002 ( .A(n697), .B(n23241), .Z(n23249) );
  XNOR U23003 ( .A(n23239), .B(n23248), .Z(n23241) );
  XNOR U23004 ( .A(n23250), .B(n23251), .Z(n23239) );
  AND U23005 ( .A(n701), .B(n23252), .Z(n23251) );
  XOR U23006 ( .A(p_input[974]), .B(n23250), .Z(n23252) );
  XNOR U23007 ( .A(n23253), .B(n23254), .Z(n23250) );
  AND U23008 ( .A(n705), .B(n23255), .Z(n23254) );
  XOR U23009 ( .A(n23256), .B(n23257), .Z(n23248) );
  AND U23010 ( .A(n709), .B(n23247), .Z(n23257) );
  XNOR U23011 ( .A(n23258), .B(n23245), .Z(n23247) );
  XOR U23012 ( .A(n23259), .B(n23260), .Z(n23245) );
  AND U23013 ( .A(n732), .B(n23261), .Z(n23260) );
  IV U23014 ( .A(n23256), .Z(n23258) );
  XOR U23015 ( .A(n23262), .B(n23263), .Z(n23256) );
  AND U23016 ( .A(n716), .B(n23255), .Z(n23263) );
  XNOR U23017 ( .A(n23253), .B(n23262), .Z(n23255) );
  XNOR U23018 ( .A(n23264), .B(n23265), .Z(n23253) );
  AND U23019 ( .A(n720), .B(n23266), .Z(n23265) );
  XOR U23020 ( .A(p_input[1006]), .B(n23264), .Z(n23266) );
  XNOR U23021 ( .A(n23267), .B(n23268), .Z(n23264) );
  AND U23022 ( .A(n724), .B(n23269), .Z(n23268) );
  XOR U23023 ( .A(n23270), .B(n23271), .Z(n23262) );
  AND U23024 ( .A(n728), .B(n23261), .Z(n23271) );
  XNOR U23025 ( .A(n23272), .B(n23259), .Z(n23261) );
  XOR U23026 ( .A(n23273), .B(n23274), .Z(n23259) );
  AND U23027 ( .A(n751), .B(n23275), .Z(n23274) );
  IV U23028 ( .A(n23270), .Z(n23272) );
  XOR U23029 ( .A(n23276), .B(n23277), .Z(n23270) );
  AND U23030 ( .A(n735), .B(n23269), .Z(n23277) );
  XNOR U23031 ( .A(n23267), .B(n23276), .Z(n23269) );
  XNOR U23032 ( .A(n23278), .B(n23279), .Z(n23267) );
  AND U23033 ( .A(n739), .B(n23280), .Z(n23279) );
  XOR U23034 ( .A(p_input[1038]), .B(n23278), .Z(n23280) );
  XNOR U23035 ( .A(n23281), .B(n23282), .Z(n23278) );
  AND U23036 ( .A(n743), .B(n23283), .Z(n23282) );
  XOR U23037 ( .A(n23284), .B(n23285), .Z(n23276) );
  AND U23038 ( .A(n747), .B(n23275), .Z(n23285) );
  XNOR U23039 ( .A(n23286), .B(n23273), .Z(n23275) );
  XOR U23040 ( .A(n23287), .B(n23288), .Z(n23273) );
  AND U23041 ( .A(n770), .B(n23289), .Z(n23288) );
  IV U23042 ( .A(n23284), .Z(n23286) );
  XOR U23043 ( .A(n23290), .B(n23291), .Z(n23284) );
  AND U23044 ( .A(n754), .B(n23283), .Z(n23291) );
  XNOR U23045 ( .A(n23281), .B(n23290), .Z(n23283) );
  XNOR U23046 ( .A(n23292), .B(n23293), .Z(n23281) );
  AND U23047 ( .A(n758), .B(n23294), .Z(n23293) );
  XOR U23048 ( .A(p_input[1070]), .B(n23292), .Z(n23294) );
  XNOR U23049 ( .A(n23295), .B(n23296), .Z(n23292) );
  AND U23050 ( .A(n762), .B(n23297), .Z(n23296) );
  XOR U23051 ( .A(n23298), .B(n23299), .Z(n23290) );
  AND U23052 ( .A(n766), .B(n23289), .Z(n23299) );
  XNOR U23053 ( .A(n23300), .B(n23287), .Z(n23289) );
  XOR U23054 ( .A(n23301), .B(n23302), .Z(n23287) );
  AND U23055 ( .A(n789), .B(n23303), .Z(n23302) );
  IV U23056 ( .A(n23298), .Z(n23300) );
  XOR U23057 ( .A(n23304), .B(n23305), .Z(n23298) );
  AND U23058 ( .A(n773), .B(n23297), .Z(n23305) );
  XNOR U23059 ( .A(n23295), .B(n23304), .Z(n23297) );
  XNOR U23060 ( .A(n23306), .B(n23307), .Z(n23295) );
  AND U23061 ( .A(n777), .B(n23308), .Z(n23307) );
  XOR U23062 ( .A(p_input[1102]), .B(n23306), .Z(n23308) );
  XNOR U23063 ( .A(n23309), .B(n23310), .Z(n23306) );
  AND U23064 ( .A(n781), .B(n23311), .Z(n23310) );
  XOR U23065 ( .A(n23312), .B(n23313), .Z(n23304) );
  AND U23066 ( .A(n785), .B(n23303), .Z(n23313) );
  XNOR U23067 ( .A(n23314), .B(n23301), .Z(n23303) );
  XOR U23068 ( .A(n23315), .B(n23316), .Z(n23301) );
  AND U23069 ( .A(n808), .B(n23317), .Z(n23316) );
  IV U23070 ( .A(n23312), .Z(n23314) );
  XOR U23071 ( .A(n23318), .B(n23319), .Z(n23312) );
  AND U23072 ( .A(n792), .B(n23311), .Z(n23319) );
  XNOR U23073 ( .A(n23309), .B(n23318), .Z(n23311) );
  XNOR U23074 ( .A(n23320), .B(n23321), .Z(n23309) );
  AND U23075 ( .A(n796), .B(n23322), .Z(n23321) );
  XOR U23076 ( .A(p_input[1134]), .B(n23320), .Z(n23322) );
  XNOR U23077 ( .A(n23323), .B(n23324), .Z(n23320) );
  AND U23078 ( .A(n800), .B(n23325), .Z(n23324) );
  XOR U23079 ( .A(n23326), .B(n23327), .Z(n23318) );
  AND U23080 ( .A(n804), .B(n23317), .Z(n23327) );
  XNOR U23081 ( .A(n23328), .B(n23315), .Z(n23317) );
  XOR U23082 ( .A(n23329), .B(n23330), .Z(n23315) );
  AND U23083 ( .A(n827), .B(n23331), .Z(n23330) );
  IV U23084 ( .A(n23326), .Z(n23328) );
  XOR U23085 ( .A(n23332), .B(n23333), .Z(n23326) );
  AND U23086 ( .A(n811), .B(n23325), .Z(n23333) );
  XNOR U23087 ( .A(n23323), .B(n23332), .Z(n23325) );
  XNOR U23088 ( .A(n23334), .B(n23335), .Z(n23323) );
  AND U23089 ( .A(n815), .B(n23336), .Z(n23335) );
  XOR U23090 ( .A(p_input[1166]), .B(n23334), .Z(n23336) );
  XNOR U23091 ( .A(n23337), .B(n23338), .Z(n23334) );
  AND U23092 ( .A(n819), .B(n23339), .Z(n23338) );
  XOR U23093 ( .A(n23340), .B(n23341), .Z(n23332) );
  AND U23094 ( .A(n823), .B(n23331), .Z(n23341) );
  XNOR U23095 ( .A(n23342), .B(n23329), .Z(n23331) );
  XOR U23096 ( .A(n23343), .B(n23344), .Z(n23329) );
  AND U23097 ( .A(n846), .B(n23345), .Z(n23344) );
  IV U23098 ( .A(n23340), .Z(n23342) );
  XOR U23099 ( .A(n23346), .B(n23347), .Z(n23340) );
  AND U23100 ( .A(n830), .B(n23339), .Z(n23347) );
  XNOR U23101 ( .A(n23337), .B(n23346), .Z(n23339) );
  XNOR U23102 ( .A(n23348), .B(n23349), .Z(n23337) );
  AND U23103 ( .A(n834), .B(n23350), .Z(n23349) );
  XOR U23104 ( .A(p_input[1198]), .B(n23348), .Z(n23350) );
  XNOR U23105 ( .A(n23351), .B(n23352), .Z(n23348) );
  AND U23106 ( .A(n838), .B(n23353), .Z(n23352) );
  XOR U23107 ( .A(n23354), .B(n23355), .Z(n23346) );
  AND U23108 ( .A(n842), .B(n23345), .Z(n23355) );
  XNOR U23109 ( .A(n23356), .B(n23343), .Z(n23345) );
  XOR U23110 ( .A(n23357), .B(n23358), .Z(n23343) );
  AND U23111 ( .A(n865), .B(n23359), .Z(n23358) );
  IV U23112 ( .A(n23354), .Z(n23356) );
  XOR U23113 ( .A(n23360), .B(n23361), .Z(n23354) );
  AND U23114 ( .A(n849), .B(n23353), .Z(n23361) );
  XNOR U23115 ( .A(n23351), .B(n23360), .Z(n23353) );
  XNOR U23116 ( .A(n23362), .B(n23363), .Z(n23351) );
  AND U23117 ( .A(n853), .B(n23364), .Z(n23363) );
  XOR U23118 ( .A(p_input[1230]), .B(n23362), .Z(n23364) );
  XNOR U23119 ( .A(n23365), .B(n23366), .Z(n23362) );
  AND U23120 ( .A(n857), .B(n23367), .Z(n23366) );
  XOR U23121 ( .A(n23368), .B(n23369), .Z(n23360) );
  AND U23122 ( .A(n861), .B(n23359), .Z(n23369) );
  XNOR U23123 ( .A(n23370), .B(n23357), .Z(n23359) );
  XOR U23124 ( .A(n23371), .B(n23372), .Z(n23357) );
  AND U23125 ( .A(n884), .B(n23373), .Z(n23372) );
  IV U23126 ( .A(n23368), .Z(n23370) );
  XOR U23127 ( .A(n23374), .B(n23375), .Z(n23368) );
  AND U23128 ( .A(n868), .B(n23367), .Z(n23375) );
  XNOR U23129 ( .A(n23365), .B(n23374), .Z(n23367) );
  XNOR U23130 ( .A(n23376), .B(n23377), .Z(n23365) );
  AND U23131 ( .A(n872), .B(n23378), .Z(n23377) );
  XOR U23132 ( .A(p_input[1262]), .B(n23376), .Z(n23378) );
  XNOR U23133 ( .A(n23379), .B(n23380), .Z(n23376) );
  AND U23134 ( .A(n876), .B(n23381), .Z(n23380) );
  XOR U23135 ( .A(n23382), .B(n23383), .Z(n23374) );
  AND U23136 ( .A(n880), .B(n23373), .Z(n23383) );
  XNOR U23137 ( .A(n23384), .B(n23371), .Z(n23373) );
  XOR U23138 ( .A(n23385), .B(n23386), .Z(n23371) );
  AND U23139 ( .A(n903), .B(n23387), .Z(n23386) );
  IV U23140 ( .A(n23382), .Z(n23384) );
  XOR U23141 ( .A(n23388), .B(n23389), .Z(n23382) );
  AND U23142 ( .A(n887), .B(n23381), .Z(n23389) );
  XNOR U23143 ( .A(n23379), .B(n23388), .Z(n23381) );
  XNOR U23144 ( .A(n23390), .B(n23391), .Z(n23379) );
  AND U23145 ( .A(n891), .B(n23392), .Z(n23391) );
  XOR U23146 ( .A(p_input[1294]), .B(n23390), .Z(n23392) );
  XNOR U23147 ( .A(n23393), .B(n23394), .Z(n23390) );
  AND U23148 ( .A(n895), .B(n23395), .Z(n23394) );
  XOR U23149 ( .A(n23396), .B(n23397), .Z(n23388) );
  AND U23150 ( .A(n899), .B(n23387), .Z(n23397) );
  XNOR U23151 ( .A(n23398), .B(n23385), .Z(n23387) );
  XOR U23152 ( .A(n23399), .B(n23400), .Z(n23385) );
  AND U23153 ( .A(n922), .B(n23401), .Z(n23400) );
  IV U23154 ( .A(n23396), .Z(n23398) );
  XOR U23155 ( .A(n23402), .B(n23403), .Z(n23396) );
  AND U23156 ( .A(n906), .B(n23395), .Z(n23403) );
  XNOR U23157 ( .A(n23393), .B(n23402), .Z(n23395) );
  XNOR U23158 ( .A(n23404), .B(n23405), .Z(n23393) );
  AND U23159 ( .A(n910), .B(n23406), .Z(n23405) );
  XOR U23160 ( .A(p_input[1326]), .B(n23404), .Z(n23406) );
  XNOR U23161 ( .A(n23407), .B(n23408), .Z(n23404) );
  AND U23162 ( .A(n914), .B(n23409), .Z(n23408) );
  XOR U23163 ( .A(n23410), .B(n23411), .Z(n23402) );
  AND U23164 ( .A(n918), .B(n23401), .Z(n23411) );
  XNOR U23165 ( .A(n23412), .B(n23399), .Z(n23401) );
  XOR U23166 ( .A(n23413), .B(n23414), .Z(n23399) );
  AND U23167 ( .A(n941), .B(n23415), .Z(n23414) );
  IV U23168 ( .A(n23410), .Z(n23412) );
  XOR U23169 ( .A(n23416), .B(n23417), .Z(n23410) );
  AND U23170 ( .A(n925), .B(n23409), .Z(n23417) );
  XNOR U23171 ( .A(n23407), .B(n23416), .Z(n23409) );
  XNOR U23172 ( .A(n23418), .B(n23419), .Z(n23407) );
  AND U23173 ( .A(n929), .B(n23420), .Z(n23419) );
  XOR U23174 ( .A(p_input[1358]), .B(n23418), .Z(n23420) );
  XNOR U23175 ( .A(n23421), .B(n23422), .Z(n23418) );
  AND U23176 ( .A(n933), .B(n23423), .Z(n23422) );
  XOR U23177 ( .A(n23424), .B(n23425), .Z(n23416) );
  AND U23178 ( .A(n937), .B(n23415), .Z(n23425) );
  XNOR U23179 ( .A(n23426), .B(n23413), .Z(n23415) );
  XOR U23180 ( .A(n23427), .B(n23428), .Z(n23413) );
  AND U23181 ( .A(n960), .B(n23429), .Z(n23428) );
  IV U23182 ( .A(n23424), .Z(n23426) );
  XOR U23183 ( .A(n23430), .B(n23431), .Z(n23424) );
  AND U23184 ( .A(n944), .B(n23423), .Z(n23431) );
  XNOR U23185 ( .A(n23421), .B(n23430), .Z(n23423) );
  XNOR U23186 ( .A(n23432), .B(n23433), .Z(n23421) );
  AND U23187 ( .A(n948), .B(n23434), .Z(n23433) );
  XOR U23188 ( .A(p_input[1390]), .B(n23432), .Z(n23434) );
  XNOR U23189 ( .A(n23435), .B(n23436), .Z(n23432) );
  AND U23190 ( .A(n952), .B(n23437), .Z(n23436) );
  XOR U23191 ( .A(n23438), .B(n23439), .Z(n23430) );
  AND U23192 ( .A(n956), .B(n23429), .Z(n23439) );
  XNOR U23193 ( .A(n23440), .B(n23427), .Z(n23429) );
  XOR U23194 ( .A(n23441), .B(n23442), .Z(n23427) );
  AND U23195 ( .A(n979), .B(n23443), .Z(n23442) );
  IV U23196 ( .A(n23438), .Z(n23440) );
  XOR U23197 ( .A(n23444), .B(n23445), .Z(n23438) );
  AND U23198 ( .A(n963), .B(n23437), .Z(n23445) );
  XNOR U23199 ( .A(n23435), .B(n23444), .Z(n23437) );
  XNOR U23200 ( .A(n23446), .B(n23447), .Z(n23435) );
  AND U23201 ( .A(n967), .B(n23448), .Z(n23447) );
  XOR U23202 ( .A(p_input[1422]), .B(n23446), .Z(n23448) );
  XNOR U23203 ( .A(n23449), .B(n23450), .Z(n23446) );
  AND U23204 ( .A(n971), .B(n23451), .Z(n23450) );
  XOR U23205 ( .A(n23452), .B(n23453), .Z(n23444) );
  AND U23206 ( .A(n975), .B(n23443), .Z(n23453) );
  XNOR U23207 ( .A(n23454), .B(n23441), .Z(n23443) );
  XOR U23208 ( .A(n23455), .B(n23456), .Z(n23441) );
  AND U23209 ( .A(n998), .B(n23457), .Z(n23456) );
  IV U23210 ( .A(n23452), .Z(n23454) );
  XOR U23211 ( .A(n23458), .B(n23459), .Z(n23452) );
  AND U23212 ( .A(n982), .B(n23451), .Z(n23459) );
  XNOR U23213 ( .A(n23449), .B(n23458), .Z(n23451) );
  XNOR U23214 ( .A(n23460), .B(n23461), .Z(n23449) );
  AND U23215 ( .A(n986), .B(n23462), .Z(n23461) );
  XOR U23216 ( .A(p_input[1454]), .B(n23460), .Z(n23462) );
  XNOR U23217 ( .A(n23463), .B(n23464), .Z(n23460) );
  AND U23218 ( .A(n990), .B(n23465), .Z(n23464) );
  XOR U23219 ( .A(n23466), .B(n23467), .Z(n23458) );
  AND U23220 ( .A(n994), .B(n23457), .Z(n23467) );
  XNOR U23221 ( .A(n23468), .B(n23455), .Z(n23457) );
  XOR U23222 ( .A(n23469), .B(n23470), .Z(n23455) );
  AND U23223 ( .A(n1017), .B(n23471), .Z(n23470) );
  IV U23224 ( .A(n23466), .Z(n23468) );
  XOR U23225 ( .A(n23472), .B(n23473), .Z(n23466) );
  AND U23226 ( .A(n1001), .B(n23465), .Z(n23473) );
  XNOR U23227 ( .A(n23463), .B(n23472), .Z(n23465) );
  XNOR U23228 ( .A(n23474), .B(n23475), .Z(n23463) );
  AND U23229 ( .A(n1005), .B(n23476), .Z(n23475) );
  XOR U23230 ( .A(p_input[1486]), .B(n23474), .Z(n23476) );
  XNOR U23231 ( .A(n23477), .B(n23478), .Z(n23474) );
  AND U23232 ( .A(n1009), .B(n23479), .Z(n23478) );
  XOR U23233 ( .A(n23480), .B(n23481), .Z(n23472) );
  AND U23234 ( .A(n1013), .B(n23471), .Z(n23481) );
  XNOR U23235 ( .A(n23482), .B(n23469), .Z(n23471) );
  XOR U23236 ( .A(n23483), .B(n23484), .Z(n23469) );
  AND U23237 ( .A(n1036), .B(n23485), .Z(n23484) );
  IV U23238 ( .A(n23480), .Z(n23482) );
  XOR U23239 ( .A(n23486), .B(n23487), .Z(n23480) );
  AND U23240 ( .A(n1020), .B(n23479), .Z(n23487) );
  XNOR U23241 ( .A(n23477), .B(n23486), .Z(n23479) );
  XNOR U23242 ( .A(n23488), .B(n23489), .Z(n23477) );
  AND U23243 ( .A(n1024), .B(n23490), .Z(n23489) );
  XOR U23244 ( .A(p_input[1518]), .B(n23488), .Z(n23490) );
  XNOR U23245 ( .A(n23491), .B(n23492), .Z(n23488) );
  AND U23246 ( .A(n1028), .B(n23493), .Z(n23492) );
  XOR U23247 ( .A(n23494), .B(n23495), .Z(n23486) );
  AND U23248 ( .A(n1032), .B(n23485), .Z(n23495) );
  XNOR U23249 ( .A(n23496), .B(n23483), .Z(n23485) );
  XOR U23250 ( .A(n23497), .B(n23498), .Z(n23483) );
  AND U23251 ( .A(n1055), .B(n23499), .Z(n23498) );
  IV U23252 ( .A(n23494), .Z(n23496) );
  XOR U23253 ( .A(n23500), .B(n23501), .Z(n23494) );
  AND U23254 ( .A(n1039), .B(n23493), .Z(n23501) );
  XNOR U23255 ( .A(n23491), .B(n23500), .Z(n23493) );
  XNOR U23256 ( .A(n23502), .B(n23503), .Z(n23491) );
  AND U23257 ( .A(n1043), .B(n23504), .Z(n23503) );
  XOR U23258 ( .A(p_input[1550]), .B(n23502), .Z(n23504) );
  XNOR U23259 ( .A(n23505), .B(n23506), .Z(n23502) );
  AND U23260 ( .A(n1047), .B(n23507), .Z(n23506) );
  XOR U23261 ( .A(n23508), .B(n23509), .Z(n23500) );
  AND U23262 ( .A(n1051), .B(n23499), .Z(n23509) );
  XNOR U23263 ( .A(n23510), .B(n23497), .Z(n23499) );
  XOR U23264 ( .A(n23511), .B(n23512), .Z(n23497) );
  AND U23265 ( .A(n1074), .B(n23513), .Z(n23512) );
  IV U23266 ( .A(n23508), .Z(n23510) );
  XOR U23267 ( .A(n23514), .B(n23515), .Z(n23508) );
  AND U23268 ( .A(n1058), .B(n23507), .Z(n23515) );
  XNOR U23269 ( .A(n23505), .B(n23514), .Z(n23507) );
  XNOR U23270 ( .A(n23516), .B(n23517), .Z(n23505) );
  AND U23271 ( .A(n1062), .B(n23518), .Z(n23517) );
  XOR U23272 ( .A(p_input[1582]), .B(n23516), .Z(n23518) );
  XNOR U23273 ( .A(n23519), .B(n23520), .Z(n23516) );
  AND U23274 ( .A(n1066), .B(n23521), .Z(n23520) );
  XOR U23275 ( .A(n23522), .B(n23523), .Z(n23514) );
  AND U23276 ( .A(n1070), .B(n23513), .Z(n23523) );
  XNOR U23277 ( .A(n23524), .B(n23511), .Z(n23513) );
  XOR U23278 ( .A(n23525), .B(n23526), .Z(n23511) );
  AND U23279 ( .A(n1093), .B(n23527), .Z(n23526) );
  IV U23280 ( .A(n23522), .Z(n23524) );
  XOR U23281 ( .A(n23528), .B(n23529), .Z(n23522) );
  AND U23282 ( .A(n1077), .B(n23521), .Z(n23529) );
  XNOR U23283 ( .A(n23519), .B(n23528), .Z(n23521) );
  XNOR U23284 ( .A(n23530), .B(n23531), .Z(n23519) );
  AND U23285 ( .A(n1081), .B(n23532), .Z(n23531) );
  XOR U23286 ( .A(p_input[1614]), .B(n23530), .Z(n23532) );
  XNOR U23287 ( .A(n23533), .B(n23534), .Z(n23530) );
  AND U23288 ( .A(n1085), .B(n23535), .Z(n23534) );
  XOR U23289 ( .A(n23536), .B(n23537), .Z(n23528) );
  AND U23290 ( .A(n1089), .B(n23527), .Z(n23537) );
  XNOR U23291 ( .A(n23538), .B(n23525), .Z(n23527) );
  XOR U23292 ( .A(n23539), .B(n23540), .Z(n23525) );
  AND U23293 ( .A(n1112), .B(n23541), .Z(n23540) );
  IV U23294 ( .A(n23536), .Z(n23538) );
  XOR U23295 ( .A(n23542), .B(n23543), .Z(n23536) );
  AND U23296 ( .A(n1096), .B(n23535), .Z(n23543) );
  XNOR U23297 ( .A(n23533), .B(n23542), .Z(n23535) );
  XNOR U23298 ( .A(n23544), .B(n23545), .Z(n23533) );
  AND U23299 ( .A(n1100), .B(n23546), .Z(n23545) );
  XOR U23300 ( .A(p_input[1646]), .B(n23544), .Z(n23546) );
  XNOR U23301 ( .A(n23547), .B(n23548), .Z(n23544) );
  AND U23302 ( .A(n1104), .B(n23549), .Z(n23548) );
  XOR U23303 ( .A(n23550), .B(n23551), .Z(n23542) );
  AND U23304 ( .A(n1108), .B(n23541), .Z(n23551) );
  XNOR U23305 ( .A(n23552), .B(n23539), .Z(n23541) );
  XOR U23306 ( .A(n23553), .B(n23554), .Z(n23539) );
  AND U23307 ( .A(n1131), .B(n23555), .Z(n23554) );
  IV U23308 ( .A(n23550), .Z(n23552) );
  XOR U23309 ( .A(n23556), .B(n23557), .Z(n23550) );
  AND U23310 ( .A(n1115), .B(n23549), .Z(n23557) );
  XNOR U23311 ( .A(n23547), .B(n23556), .Z(n23549) );
  XNOR U23312 ( .A(n23558), .B(n23559), .Z(n23547) );
  AND U23313 ( .A(n1119), .B(n23560), .Z(n23559) );
  XOR U23314 ( .A(p_input[1678]), .B(n23558), .Z(n23560) );
  XNOR U23315 ( .A(n23561), .B(n23562), .Z(n23558) );
  AND U23316 ( .A(n1123), .B(n23563), .Z(n23562) );
  XOR U23317 ( .A(n23564), .B(n23565), .Z(n23556) );
  AND U23318 ( .A(n1127), .B(n23555), .Z(n23565) );
  XNOR U23319 ( .A(n23566), .B(n23553), .Z(n23555) );
  XOR U23320 ( .A(n23567), .B(n23568), .Z(n23553) );
  AND U23321 ( .A(n1150), .B(n23569), .Z(n23568) );
  IV U23322 ( .A(n23564), .Z(n23566) );
  XOR U23323 ( .A(n23570), .B(n23571), .Z(n23564) );
  AND U23324 ( .A(n1134), .B(n23563), .Z(n23571) );
  XNOR U23325 ( .A(n23561), .B(n23570), .Z(n23563) );
  XNOR U23326 ( .A(n23572), .B(n23573), .Z(n23561) );
  AND U23327 ( .A(n1138), .B(n23574), .Z(n23573) );
  XOR U23328 ( .A(p_input[1710]), .B(n23572), .Z(n23574) );
  XNOR U23329 ( .A(n23575), .B(n23576), .Z(n23572) );
  AND U23330 ( .A(n1142), .B(n23577), .Z(n23576) );
  XOR U23331 ( .A(n23578), .B(n23579), .Z(n23570) );
  AND U23332 ( .A(n1146), .B(n23569), .Z(n23579) );
  XNOR U23333 ( .A(n23580), .B(n23567), .Z(n23569) );
  XOR U23334 ( .A(n23581), .B(n23582), .Z(n23567) );
  AND U23335 ( .A(n1169), .B(n23583), .Z(n23582) );
  IV U23336 ( .A(n23578), .Z(n23580) );
  XOR U23337 ( .A(n23584), .B(n23585), .Z(n23578) );
  AND U23338 ( .A(n1153), .B(n23577), .Z(n23585) );
  XNOR U23339 ( .A(n23575), .B(n23584), .Z(n23577) );
  XNOR U23340 ( .A(n23586), .B(n23587), .Z(n23575) );
  AND U23341 ( .A(n1157), .B(n23588), .Z(n23587) );
  XOR U23342 ( .A(p_input[1742]), .B(n23586), .Z(n23588) );
  XNOR U23343 ( .A(n23589), .B(n23590), .Z(n23586) );
  AND U23344 ( .A(n1161), .B(n23591), .Z(n23590) );
  XOR U23345 ( .A(n23592), .B(n23593), .Z(n23584) );
  AND U23346 ( .A(n1165), .B(n23583), .Z(n23593) );
  XNOR U23347 ( .A(n23594), .B(n23581), .Z(n23583) );
  XOR U23348 ( .A(n23595), .B(n23596), .Z(n23581) );
  AND U23349 ( .A(n1188), .B(n23597), .Z(n23596) );
  IV U23350 ( .A(n23592), .Z(n23594) );
  XOR U23351 ( .A(n23598), .B(n23599), .Z(n23592) );
  AND U23352 ( .A(n1172), .B(n23591), .Z(n23599) );
  XNOR U23353 ( .A(n23589), .B(n23598), .Z(n23591) );
  XNOR U23354 ( .A(n23600), .B(n23601), .Z(n23589) );
  AND U23355 ( .A(n1176), .B(n23602), .Z(n23601) );
  XOR U23356 ( .A(p_input[1774]), .B(n23600), .Z(n23602) );
  XNOR U23357 ( .A(n23603), .B(n23604), .Z(n23600) );
  AND U23358 ( .A(n1180), .B(n23605), .Z(n23604) );
  XOR U23359 ( .A(n23606), .B(n23607), .Z(n23598) );
  AND U23360 ( .A(n1184), .B(n23597), .Z(n23607) );
  XNOR U23361 ( .A(n23608), .B(n23595), .Z(n23597) );
  XOR U23362 ( .A(n23609), .B(n23610), .Z(n23595) );
  AND U23363 ( .A(n1207), .B(n23611), .Z(n23610) );
  IV U23364 ( .A(n23606), .Z(n23608) );
  XOR U23365 ( .A(n23612), .B(n23613), .Z(n23606) );
  AND U23366 ( .A(n1191), .B(n23605), .Z(n23613) );
  XNOR U23367 ( .A(n23603), .B(n23612), .Z(n23605) );
  XNOR U23368 ( .A(n23614), .B(n23615), .Z(n23603) );
  AND U23369 ( .A(n1195), .B(n23616), .Z(n23615) );
  XOR U23370 ( .A(p_input[1806]), .B(n23614), .Z(n23616) );
  XNOR U23371 ( .A(n23617), .B(n23618), .Z(n23614) );
  AND U23372 ( .A(n1199), .B(n23619), .Z(n23618) );
  XOR U23373 ( .A(n23620), .B(n23621), .Z(n23612) );
  AND U23374 ( .A(n1203), .B(n23611), .Z(n23621) );
  XNOR U23375 ( .A(n23622), .B(n23609), .Z(n23611) );
  XOR U23376 ( .A(n23623), .B(n23624), .Z(n23609) );
  AND U23377 ( .A(n1226), .B(n23625), .Z(n23624) );
  IV U23378 ( .A(n23620), .Z(n23622) );
  XOR U23379 ( .A(n23626), .B(n23627), .Z(n23620) );
  AND U23380 ( .A(n1210), .B(n23619), .Z(n23627) );
  XNOR U23381 ( .A(n23617), .B(n23626), .Z(n23619) );
  XNOR U23382 ( .A(n23628), .B(n23629), .Z(n23617) );
  AND U23383 ( .A(n1214), .B(n23630), .Z(n23629) );
  XOR U23384 ( .A(p_input[1838]), .B(n23628), .Z(n23630) );
  XNOR U23385 ( .A(n23631), .B(n23632), .Z(n23628) );
  AND U23386 ( .A(n1218), .B(n23633), .Z(n23632) );
  XOR U23387 ( .A(n23634), .B(n23635), .Z(n23626) );
  AND U23388 ( .A(n1222), .B(n23625), .Z(n23635) );
  XNOR U23389 ( .A(n23636), .B(n23623), .Z(n23625) );
  XOR U23390 ( .A(n23637), .B(n23638), .Z(n23623) );
  AND U23391 ( .A(n1245), .B(n23639), .Z(n23638) );
  IV U23392 ( .A(n23634), .Z(n23636) );
  XOR U23393 ( .A(n23640), .B(n23641), .Z(n23634) );
  AND U23394 ( .A(n1229), .B(n23633), .Z(n23641) );
  XNOR U23395 ( .A(n23631), .B(n23640), .Z(n23633) );
  XNOR U23396 ( .A(n23642), .B(n23643), .Z(n23631) );
  AND U23397 ( .A(n1233), .B(n23644), .Z(n23643) );
  XOR U23398 ( .A(p_input[1870]), .B(n23642), .Z(n23644) );
  XNOR U23399 ( .A(n23645), .B(n23646), .Z(n23642) );
  AND U23400 ( .A(n1237), .B(n23647), .Z(n23646) );
  XOR U23401 ( .A(n23648), .B(n23649), .Z(n23640) );
  AND U23402 ( .A(n1241), .B(n23639), .Z(n23649) );
  XNOR U23403 ( .A(n23650), .B(n23637), .Z(n23639) );
  XOR U23404 ( .A(n23651), .B(n23652), .Z(n23637) );
  AND U23405 ( .A(n1264), .B(n23653), .Z(n23652) );
  IV U23406 ( .A(n23648), .Z(n23650) );
  XOR U23407 ( .A(n23654), .B(n23655), .Z(n23648) );
  AND U23408 ( .A(n1248), .B(n23647), .Z(n23655) );
  XNOR U23409 ( .A(n23645), .B(n23654), .Z(n23647) );
  XNOR U23410 ( .A(n23656), .B(n23657), .Z(n23645) );
  AND U23411 ( .A(n1252), .B(n23658), .Z(n23657) );
  XOR U23412 ( .A(p_input[1902]), .B(n23656), .Z(n23658) );
  XNOR U23413 ( .A(n23659), .B(n23660), .Z(n23656) );
  AND U23414 ( .A(n1256), .B(n23661), .Z(n23660) );
  XOR U23415 ( .A(n23662), .B(n23663), .Z(n23654) );
  AND U23416 ( .A(n1260), .B(n23653), .Z(n23663) );
  XNOR U23417 ( .A(n23664), .B(n23651), .Z(n23653) );
  XOR U23418 ( .A(n23665), .B(n23666), .Z(n23651) );
  AND U23419 ( .A(n1282), .B(n23667), .Z(n23666) );
  IV U23420 ( .A(n23662), .Z(n23664) );
  XOR U23421 ( .A(n23668), .B(n23669), .Z(n23662) );
  AND U23422 ( .A(n1267), .B(n23661), .Z(n23669) );
  XNOR U23423 ( .A(n23659), .B(n23668), .Z(n23661) );
  XNOR U23424 ( .A(n23670), .B(n23671), .Z(n23659) );
  AND U23425 ( .A(n1271), .B(n23672), .Z(n23671) );
  XOR U23426 ( .A(p_input[1934]), .B(n23670), .Z(n23672) );
  XOR U23427 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n23673), 
        .Z(n23670) );
  AND U23428 ( .A(n1274), .B(n23674), .Z(n23673) );
  XOR U23429 ( .A(n23675), .B(n23676), .Z(n23668) );
  AND U23430 ( .A(n1278), .B(n23667), .Z(n23676) );
  XNOR U23431 ( .A(n23677), .B(n23665), .Z(n23667) );
  XOR U23432 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n23678), .Z(n23665) );
  AND U23433 ( .A(n1290), .B(n23679), .Z(n23678) );
  IV U23434 ( .A(n23675), .Z(n23677) );
  XOR U23435 ( .A(n23680), .B(n23681), .Z(n23675) );
  AND U23436 ( .A(n1285), .B(n23674), .Z(n23681) );
  XOR U23437 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n23680), 
        .Z(n23674) );
  XOR U23438 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(n23682), 
        .Z(n23680) );
  AND U23439 ( .A(n1287), .B(n23679), .Z(n23682) );
  XOR U23440 ( .A(\knn_comb_/min_val_out[0][14] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n23679) );
  XOR U23441 ( .A(n113), .B(n23683), .Z(o[13]) );
  AND U23442 ( .A(n122), .B(n23684), .Z(n113) );
  XOR U23443 ( .A(n114), .B(n23683), .Z(n23684) );
  XOR U23444 ( .A(n23685), .B(n23686), .Z(n23683) );
  AND U23445 ( .A(n142), .B(n23687), .Z(n23686) );
  XOR U23446 ( .A(n23688), .B(n43), .Z(n114) );
  AND U23447 ( .A(n125), .B(n23689), .Z(n43) );
  XOR U23448 ( .A(n44), .B(n23688), .Z(n23689) );
  XOR U23449 ( .A(n23690), .B(n23691), .Z(n44) );
  AND U23450 ( .A(n130), .B(n23692), .Z(n23691) );
  XOR U23451 ( .A(p_input[13]), .B(n23690), .Z(n23692) );
  XNOR U23452 ( .A(n23693), .B(n23694), .Z(n23690) );
  AND U23453 ( .A(n134), .B(n23695), .Z(n23694) );
  XOR U23454 ( .A(n23696), .B(n23697), .Z(n23688) );
  AND U23455 ( .A(n138), .B(n23687), .Z(n23697) );
  XNOR U23456 ( .A(n23698), .B(n23685), .Z(n23687) );
  XOR U23457 ( .A(n23699), .B(n23700), .Z(n23685) );
  AND U23458 ( .A(n162), .B(n23701), .Z(n23700) );
  IV U23459 ( .A(n23696), .Z(n23698) );
  XOR U23460 ( .A(n23702), .B(n23703), .Z(n23696) );
  AND U23461 ( .A(n146), .B(n23695), .Z(n23703) );
  XNOR U23462 ( .A(n23693), .B(n23702), .Z(n23695) );
  XNOR U23463 ( .A(n23704), .B(n23705), .Z(n23693) );
  AND U23464 ( .A(n150), .B(n23706), .Z(n23705) );
  XOR U23465 ( .A(p_input[45]), .B(n23704), .Z(n23706) );
  XNOR U23466 ( .A(n23707), .B(n23708), .Z(n23704) );
  AND U23467 ( .A(n154), .B(n23709), .Z(n23708) );
  XOR U23468 ( .A(n23710), .B(n23711), .Z(n23702) );
  AND U23469 ( .A(n158), .B(n23701), .Z(n23711) );
  XNOR U23470 ( .A(n23712), .B(n23699), .Z(n23701) );
  XOR U23471 ( .A(n23713), .B(n23714), .Z(n23699) );
  AND U23472 ( .A(n181), .B(n23715), .Z(n23714) );
  IV U23473 ( .A(n23710), .Z(n23712) );
  XOR U23474 ( .A(n23716), .B(n23717), .Z(n23710) );
  AND U23475 ( .A(n165), .B(n23709), .Z(n23717) );
  XNOR U23476 ( .A(n23707), .B(n23716), .Z(n23709) );
  XNOR U23477 ( .A(n23718), .B(n23719), .Z(n23707) );
  AND U23478 ( .A(n169), .B(n23720), .Z(n23719) );
  XOR U23479 ( .A(p_input[77]), .B(n23718), .Z(n23720) );
  XNOR U23480 ( .A(n23721), .B(n23722), .Z(n23718) );
  AND U23481 ( .A(n173), .B(n23723), .Z(n23722) );
  XOR U23482 ( .A(n23724), .B(n23725), .Z(n23716) );
  AND U23483 ( .A(n177), .B(n23715), .Z(n23725) );
  XNOR U23484 ( .A(n23726), .B(n23713), .Z(n23715) );
  XOR U23485 ( .A(n23727), .B(n23728), .Z(n23713) );
  AND U23486 ( .A(n200), .B(n23729), .Z(n23728) );
  IV U23487 ( .A(n23724), .Z(n23726) );
  XOR U23488 ( .A(n23730), .B(n23731), .Z(n23724) );
  AND U23489 ( .A(n184), .B(n23723), .Z(n23731) );
  XNOR U23490 ( .A(n23721), .B(n23730), .Z(n23723) );
  XNOR U23491 ( .A(n23732), .B(n23733), .Z(n23721) );
  AND U23492 ( .A(n188), .B(n23734), .Z(n23733) );
  XOR U23493 ( .A(p_input[109]), .B(n23732), .Z(n23734) );
  XNOR U23494 ( .A(n23735), .B(n23736), .Z(n23732) );
  AND U23495 ( .A(n192), .B(n23737), .Z(n23736) );
  XOR U23496 ( .A(n23738), .B(n23739), .Z(n23730) );
  AND U23497 ( .A(n196), .B(n23729), .Z(n23739) );
  XNOR U23498 ( .A(n23740), .B(n23727), .Z(n23729) );
  XOR U23499 ( .A(n23741), .B(n23742), .Z(n23727) );
  AND U23500 ( .A(n219), .B(n23743), .Z(n23742) );
  IV U23501 ( .A(n23738), .Z(n23740) );
  XOR U23502 ( .A(n23744), .B(n23745), .Z(n23738) );
  AND U23503 ( .A(n203), .B(n23737), .Z(n23745) );
  XNOR U23504 ( .A(n23735), .B(n23744), .Z(n23737) );
  XNOR U23505 ( .A(n23746), .B(n23747), .Z(n23735) );
  AND U23506 ( .A(n207), .B(n23748), .Z(n23747) );
  XOR U23507 ( .A(p_input[141]), .B(n23746), .Z(n23748) );
  XNOR U23508 ( .A(n23749), .B(n23750), .Z(n23746) );
  AND U23509 ( .A(n211), .B(n23751), .Z(n23750) );
  XOR U23510 ( .A(n23752), .B(n23753), .Z(n23744) );
  AND U23511 ( .A(n215), .B(n23743), .Z(n23753) );
  XNOR U23512 ( .A(n23754), .B(n23741), .Z(n23743) );
  XOR U23513 ( .A(n23755), .B(n23756), .Z(n23741) );
  AND U23514 ( .A(n238), .B(n23757), .Z(n23756) );
  IV U23515 ( .A(n23752), .Z(n23754) );
  XOR U23516 ( .A(n23758), .B(n23759), .Z(n23752) );
  AND U23517 ( .A(n222), .B(n23751), .Z(n23759) );
  XNOR U23518 ( .A(n23749), .B(n23758), .Z(n23751) );
  XNOR U23519 ( .A(n23760), .B(n23761), .Z(n23749) );
  AND U23520 ( .A(n226), .B(n23762), .Z(n23761) );
  XOR U23521 ( .A(p_input[173]), .B(n23760), .Z(n23762) );
  XNOR U23522 ( .A(n23763), .B(n23764), .Z(n23760) );
  AND U23523 ( .A(n230), .B(n23765), .Z(n23764) );
  XOR U23524 ( .A(n23766), .B(n23767), .Z(n23758) );
  AND U23525 ( .A(n234), .B(n23757), .Z(n23767) );
  XNOR U23526 ( .A(n23768), .B(n23755), .Z(n23757) );
  XOR U23527 ( .A(n23769), .B(n23770), .Z(n23755) );
  AND U23528 ( .A(n257), .B(n23771), .Z(n23770) );
  IV U23529 ( .A(n23766), .Z(n23768) );
  XOR U23530 ( .A(n23772), .B(n23773), .Z(n23766) );
  AND U23531 ( .A(n241), .B(n23765), .Z(n23773) );
  XNOR U23532 ( .A(n23763), .B(n23772), .Z(n23765) );
  XNOR U23533 ( .A(n23774), .B(n23775), .Z(n23763) );
  AND U23534 ( .A(n245), .B(n23776), .Z(n23775) );
  XOR U23535 ( .A(p_input[205]), .B(n23774), .Z(n23776) );
  XNOR U23536 ( .A(n23777), .B(n23778), .Z(n23774) );
  AND U23537 ( .A(n249), .B(n23779), .Z(n23778) );
  XOR U23538 ( .A(n23780), .B(n23781), .Z(n23772) );
  AND U23539 ( .A(n253), .B(n23771), .Z(n23781) );
  XNOR U23540 ( .A(n23782), .B(n23769), .Z(n23771) );
  XOR U23541 ( .A(n23783), .B(n23784), .Z(n23769) );
  AND U23542 ( .A(n276), .B(n23785), .Z(n23784) );
  IV U23543 ( .A(n23780), .Z(n23782) );
  XOR U23544 ( .A(n23786), .B(n23787), .Z(n23780) );
  AND U23545 ( .A(n260), .B(n23779), .Z(n23787) );
  XNOR U23546 ( .A(n23777), .B(n23786), .Z(n23779) );
  XNOR U23547 ( .A(n23788), .B(n23789), .Z(n23777) );
  AND U23548 ( .A(n264), .B(n23790), .Z(n23789) );
  XOR U23549 ( .A(p_input[237]), .B(n23788), .Z(n23790) );
  XNOR U23550 ( .A(n23791), .B(n23792), .Z(n23788) );
  AND U23551 ( .A(n268), .B(n23793), .Z(n23792) );
  XOR U23552 ( .A(n23794), .B(n23795), .Z(n23786) );
  AND U23553 ( .A(n272), .B(n23785), .Z(n23795) );
  XNOR U23554 ( .A(n23796), .B(n23783), .Z(n23785) );
  XOR U23555 ( .A(n23797), .B(n23798), .Z(n23783) );
  AND U23556 ( .A(n295), .B(n23799), .Z(n23798) );
  IV U23557 ( .A(n23794), .Z(n23796) );
  XOR U23558 ( .A(n23800), .B(n23801), .Z(n23794) );
  AND U23559 ( .A(n279), .B(n23793), .Z(n23801) );
  XNOR U23560 ( .A(n23791), .B(n23800), .Z(n23793) );
  XNOR U23561 ( .A(n23802), .B(n23803), .Z(n23791) );
  AND U23562 ( .A(n283), .B(n23804), .Z(n23803) );
  XOR U23563 ( .A(p_input[269]), .B(n23802), .Z(n23804) );
  XNOR U23564 ( .A(n23805), .B(n23806), .Z(n23802) );
  AND U23565 ( .A(n287), .B(n23807), .Z(n23806) );
  XOR U23566 ( .A(n23808), .B(n23809), .Z(n23800) );
  AND U23567 ( .A(n291), .B(n23799), .Z(n23809) );
  XNOR U23568 ( .A(n23810), .B(n23797), .Z(n23799) );
  XOR U23569 ( .A(n23811), .B(n23812), .Z(n23797) );
  AND U23570 ( .A(n314), .B(n23813), .Z(n23812) );
  IV U23571 ( .A(n23808), .Z(n23810) );
  XOR U23572 ( .A(n23814), .B(n23815), .Z(n23808) );
  AND U23573 ( .A(n298), .B(n23807), .Z(n23815) );
  XNOR U23574 ( .A(n23805), .B(n23814), .Z(n23807) );
  XNOR U23575 ( .A(n23816), .B(n23817), .Z(n23805) );
  AND U23576 ( .A(n302), .B(n23818), .Z(n23817) );
  XOR U23577 ( .A(p_input[301]), .B(n23816), .Z(n23818) );
  XNOR U23578 ( .A(n23819), .B(n23820), .Z(n23816) );
  AND U23579 ( .A(n306), .B(n23821), .Z(n23820) );
  XOR U23580 ( .A(n23822), .B(n23823), .Z(n23814) );
  AND U23581 ( .A(n310), .B(n23813), .Z(n23823) );
  XNOR U23582 ( .A(n23824), .B(n23811), .Z(n23813) );
  XOR U23583 ( .A(n23825), .B(n23826), .Z(n23811) );
  AND U23584 ( .A(n333), .B(n23827), .Z(n23826) );
  IV U23585 ( .A(n23822), .Z(n23824) );
  XOR U23586 ( .A(n23828), .B(n23829), .Z(n23822) );
  AND U23587 ( .A(n317), .B(n23821), .Z(n23829) );
  XNOR U23588 ( .A(n23819), .B(n23828), .Z(n23821) );
  XNOR U23589 ( .A(n23830), .B(n23831), .Z(n23819) );
  AND U23590 ( .A(n321), .B(n23832), .Z(n23831) );
  XOR U23591 ( .A(p_input[333]), .B(n23830), .Z(n23832) );
  XNOR U23592 ( .A(n23833), .B(n23834), .Z(n23830) );
  AND U23593 ( .A(n325), .B(n23835), .Z(n23834) );
  XOR U23594 ( .A(n23836), .B(n23837), .Z(n23828) );
  AND U23595 ( .A(n329), .B(n23827), .Z(n23837) );
  XNOR U23596 ( .A(n23838), .B(n23825), .Z(n23827) );
  XOR U23597 ( .A(n23839), .B(n23840), .Z(n23825) );
  AND U23598 ( .A(n352), .B(n23841), .Z(n23840) );
  IV U23599 ( .A(n23836), .Z(n23838) );
  XOR U23600 ( .A(n23842), .B(n23843), .Z(n23836) );
  AND U23601 ( .A(n336), .B(n23835), .Z(n23843) );
  XNOR U23602 ( .A(n23833), .B(n23842), .Z(n23835) );
  XNOR U23603 ( .A(n23844), .B(n23845), .Z(n23833) );
  AND U23604 ( .A(n340), .B(n23846), .Z(n23845) );
  XOR U23605 ( .A(p_input[365]), .B(n23844), .Z(n23846) );
  XNOR U23606 ( .A(n23847), .B(n23848), .Z(n23844) );
  AND U23607 ( .A(n344), .B(n23849), .Z(n23848) );
  XOR U23608 ( .A(n23850), .B(n23851), .Z(n23842) );
  AND U23609 ( .A(n348), .B(n23841), .Z(n23851) );
  XNOR U23610 ( .A(n23852), .B(n23839), .Z(n23841) );
  XOR U23611 ( .A(n23853), .B(n23854), .Z(n23839) );
  AND U23612 ( .A(n371), .B(n23855), .Z(n23854) );
  IV U23613 ( .A(n23850), .Z(n23852) );
  XOR U23614 ( .A(n23856), .B(n23857), .Z(n23850) );
  AND U23615 ( .A(n355), .B(n23849), .Z(n23857) );
  XNOR U23616 ( .A(n23847), .B(n23856), .Z(n23849) );
  XNOR U23617 ( .A(n23858), .B(n23859), .Z(n23847) );
  AND U23618 ( .A(n359), .B(n23860), .Z(n23859) );
  XOR U23619 ( .A(p_input[397]), .B(n23858), .Z(n23860) );
  XNOR U23620 ( .A(n23861), .B(n23862), .Z(n23858) );
  AND U23621 ( .A(n363), .B(n23863), .Z(n23862) );
  XOR U23622 ( .A(n23864), .B(n23865), .Z(n23856) );
  AND U23623 ( .A(n367), .B(n23855), .Z(n23865) );
  XNOR U23624 ( .A(n23866), .B(n23853), .Z(n23855) );
  XOR U23625 ( .A(n23867), .B(n23868), .Z(n23853) );
  AND U23626 ( .A(n390), .B(n23869), .Z(n23868) );
  IV U23627 ( .A(n23864), .Z(n23866) );
  XOR U23628 ( .A(n23870), .B(n23871), .Z(n23864) );
  AND U23629 ( .A(n374), .B(n23863), .Z(n23871) );
  XNOR U23630 ( .A(n23861), .B(n23870), .Z(n23863) );
  XNOR U23631 ( .A(n23872), .B(n23873), .Z(n23861) );
  AND U23632 ( .A(n378), .B(n23874), .Z(n23873) );
  XOR U23633 ( .A(p_input[429]), .B(n23872), .Z(n23874) );
  XNOR U23634 ( .A(n23875), .B(n23876), .Z(n23872) );
  AND U23635 ( .A(n382), .B(n23877), .Z(n23876) );
  XOR U23636 ( .A(n23878), .B(n23879), .Z(n23870) );
  AND U23637 ( .A(n386), .B(n23869), .Z(n23879) );
  XNOR U23638 ( .A(n23880), .B(n23867), .Z(n23869) );
  XOR U23639 ( .A(n23881), .B(n23882), .Z(n23867) );
  AND U23640 ( .A(n409), .B(n23883), .Z(n23882) );
  IV U23641 ( .A(n23878), .Z(n23880) );
  XOR U23642 ( .A(n23884), .B(n23885), .Z(n23878) );
  AND U23643 ( .A(n393), .B(n23877), .Z(n23885) );
  XNOR U23644 ( .A(n23875), .B(n23884), .Z(n23877) );
  XNOR U23645 ( .A(n23886), .B(n23887), .Z(n23875) );
  AND U23646 ( .A(n397), .B(n23888), .Z(n23887) );
  XOR U23647 ( .A(p_input[461]), .B(n23886), .Z(n23888) );
  XNOR U23648 ( .A(n23889), .B(n23890), .Z(n23886) );
  AND U23649 ( .A(n401), .B(n23891), .Z(n23890) );
  XOR U23650 ( .A(n23892), .B(n23893), .Z(n23884) );
  AND U23651 ( .A(n405), .B(n23883), .Z(n23893) );
  XNOR U23652 ( .A(n23894), .B(n23881), .Z(n23883) );
  XOR U23653 ( .A(n23895), .B(n23896), .Z(n23881) );
  AND U23654 ( .A(n428), .B(n23897), .Z(n23896) );
  IV U23655 ( .A(n23892), .Z(n23894) );
  XOR U23656 ( .A(n23898), .B(n23899), .Z(n23892) );
  AND U23657 ( .A(n412), .B(n23891), .Z(n23899) );
  XNOR U23658 ( .A(n23889), .B(n23898), .Z(n23891) );
  XNOR U23659 ( .A(n23900), .B(n23901), .Z(n23889) );
  AND U23660 ( .A(n416), .B(n23902), .Z(n23901) );
  XOR U23661 ( .A(p_input[493]), .B(n23900), .Z(n23902) );
  XNOR U23662 ( .A(n23903), .B(n23904), .Z(n23900) );
  AND U23663 ( .A(n420), .B(n23905), .Z(n23904) );
  XOR U23664 ( .A(n23906), .B(n23907), .Z(n23898) );
  AND U23665 ( .A(n424), .B(n23897), .Z(n23907) );
  XNOR U23666 ( .A(n23908), .B(n23895), .Z(n23897) );
  XOR U23667 ( .A(n23909), .B(n23910), .Z(n23895) );
  AND U23668 ( .A(n447), .B(n23911), .Z(n23910) );
  IV U23669 ( .A(n23906), .Z(n23908) );
  XOR U23670 ( .A(n23912), .B(n23913), .Z(n23906) );
  AND U23671 ( .A(n431), .B(n23905), .Z(n23913) );
  XNOR U23672 ( .A(n23903), .B(n23912), .Z(n23905) );
  XNOR U23673 ( .A(n23914), .B(n23915), .Z(n23903) );
  AND U23674 ( .A(n435), .B(n23916), .Z(n23915) );
  XOR U23675 ( .A(p_input[525]), .B(n23914), .Z(n23916) );
  XNOR U23676 ( .A(n23917), .B(n23918), .Z(n23914) );
  AND U23677 ( .A(n439), .B(n23919), .Z(n23918) );
  XOR U23678 ( .A(n23920), .B(n23921), .Z(n23912) );
  AND U23679 ( .A(n443), .B(n23911), .Z(n23921) );
  XNOR U23680 ( .A(n23922), .B(n23909), .Z(n23911) );
  XOR U23681 ( .A(n23923), .B(n23924), .Z(n23909) );
  AND U23682 ( .A(n466), .B(n23925), .Z(n23924) );
  IV U23683 ( .A(n23920), .Z(n23922) );
  XOR U23684 ( .A(n23926), .B(n23927), .Z(n23920) );
  AND U23685 ( .A(n450), .B(n23919), .Z(n23927) );
  XNOR U23686 ( .A(n23917), .B(n23926), .Z(n23919) );
  XNOR U23687 ( .A(n23928), .B(n23929), .Z(n23917) );
  AND U23688 ( .A(n454), .B(n23930), .Z(n23929) );
  XOR U23689 ( .A(p_input[557]), .B(n23928), .Z(n23930) );
  XNOR U23690 ( .A(n23931), .B(n23932), .Z(n23928) );
  AND U23691 ( .A(n458), .B(n23933), .Z(n23932) );
  XOR U23692 ( .A(n23934), .B(n23935), .Z(n23926) );
  AND U23693 ( .A(n462), .B(n23925), .Z(n23935) );
  XNOR U23694 ( .A(n23936), .B(n23923), .Z(n23925) );
  XOR U23695 ( .A(n23937), .B(n23938), .Z(n23923) );
  AND U23696 ( .A(n485), .B(n23939), .Z(n23938) );
  IV U23697 ( .A(n23934), .Z(n23936) );
  XOR U23698 ( .A(n23940), .B(n23941), .Z(n23934) );
  AND U23699 ( .A(n469), .B(n23933), .Z(n23941) );
  XNOR U23700 ( .A(n23931), .B(n23940), .Z(n23933) );
  XNOR U23701 ( .A(n23942), .B(n23943), .Z(n23931) );
  AND U23702 ( .A(n473), .B(n23944), .Z(n23943) );
  XOR U23703 ( .A(p_input[589]), .B(n23942), .Z(n23944) );
  XNOR U23704 ( .A(n23945), .B(n23946), .Z(n23942) );
  AND U23705 ( .A(n477), .B(n23947), .Z(n23946) );
  XOR U23706 ( .A(n23948), .B(n23949), .Z(n23940) );
  AND U23707 ( .A(n481), .B(n23939), .Z(n23949) );
  XNOR U23708 ( .A(n23950), .B(n23937), .Z(n23939) );
  XOR U23709 ( .A(n23951), .B(n23952), .Z(n23937) );
  AND U23710 ( .A(n504), .B(n23953), .Z(n23952) );
  IV U23711 ( .A(n23948), .Z(n23950) );
  XOR U23712 ( .A(n23954), .B(n23955), .Z(n23948) );
  AND U23713 ( .A(n488), .B(n23947), .Z(n23955) );
  XNOR U23714 ( .A(n23945), .B(n23954), .Z(n23947) );
  XNOR U23715 ( .A(n23956), .B(n23957), .Z(n23945) );
  AND U23716 ( .A(n492), .B(n23958), .Z(n23957) );
  XOR U23717 ( .A(p_input[621]), .B(n23956), .Z(n23958) );
  XNOR U23718 ( .A(n23959), .B(n23960), .Z(n23956) );
  AND U23719 ( .A(n496), .B(n23961), .Z(n23960) );
  XOR U23720 ( .A(n23962), .B(n23963), .Z(n23954) );
  AND U23721 ( .A(n500), .B(n23953), .Z(n23963) );
  XNOR U23722 ( .A(n23964), .B(n23951), .Z(n23953) );
  XOR U23723 ( .A(n23965), .B(n23966), .Z(n23951) );
  AND U23724 ( .A(n523), .B(n23967), .Z(n23966) );
  IV U23725 ( .A(n23962), .Z(n23964) );
  XOR U23726 ( .A(n23968), .B(n23969), .Z(n23962) );
  AND U23727 ( .A(n507), .B(n23961), .Z(n23969) );
  XNOR U23728 ( .A(n23959), .B(n23968), .Z(n23961) );
  XNOR U23729 ( .A(n23970), .B(n23971), .Z(n23959) );
  AND U23730 ( .A(n511), .B(n23972), .Z(n23971) );
  XOR U23731 ( .A(p_input[653]), .B(n23970), .Z(n23972) );
  XNOR U23732 ( .A(n23973), .B(n23974), .Z(n23970) );
  AND U23733 ( .A(n515), .B(n23975), .Z(n23974) );
  XOR U23734 ( .A(n23976), .B(n23977), .Z(n23968) );
  AND U23735 ( .A(n519), .B(n23967), .Z(n23977) );
  XNOR U23736 ( .A(n23978), .B(n23965), .Z(n23967) );
  XOR U23737 ( .A(n23979), .B(n23980), .Z(n23965) );
  AND U23738 ( .A(n542), .B(n23981), .Z(n23980) );
  IV U23739 ( .A(n23976), .Z(n23978) );
  XOR U23740 ( .A(n23982), .B(n23983), .Z(n23976) );
  AND U23741 ( .A(n526), .B(n23975), .Z(n23983) );
  XNOR U23742 ( .A(n23973), .B(n23982), .Z(n23975) );
  XNOR U23743 ( .A(n23984), .B(n23985), .Z(n23973) );
  AND U23744 ( .A(n530), .B(n23986), .Z(n23985) );
  XOR U23745 ( .A(p_input[685]), .B(n23984), .Z(n23986) );
  XNOR U23746 ( .A(n23987), .B(n23988), .Z(n23984) );
  AND U23747 ( .A(n534), .B(n23989), .Z(n23988) );
  XOR U23748 ( .A(n23990), .B(n23991), .Z(n23982) );
  AND U23749 ( .A(n538), .B(n23981), .Z(n23991) );
  XNOR U23750 ( .A(n23992), .B(n23979), .Z(n23981) );
  XOR U23751 ( .A(n23993), .B(n23994), .Z(n23979) );
  AND U23752 ( .A(n561), .B(n23995), .Z(n23994) );
  IV U23753 ( .A(n23990), .Z(n23992) );
  XOR U23754 ( .A(n23996), .B(n23997), .Z(n23990) );
  AND U23755 ( .A(n545), .B(n23989), .Z(n23997) );
  XNOR U23756 ( .A(n23987), .B(n23996), .Z(n23989) );
  XNOR U23757 ( .A(n23998), .B(n23999), .Z(n23987) );
  AND U23758 ( .A(n549), .B(n24000), .Z(n23999) );
  XOR U23759 ( .A(p_input[717]), .B(n23998), .Z(n24000) );
  XNOR U23760 ( .A(n24001), .B(n24002), .Z(n23998) );
  AND U23761 ( .A(n553), .B(n24003), .Z(n24002) );
  XOR U23762 ( .A(n24004), .B(n24005), .Z(n23996) );
  AND U23763 ( .A(n557), .B(n23995), .Z(n24005) );
  XNOR U23764 ( .A(n24006), .B(n23993), .Z(n23995) );
  XOR U23765 ( .A(n24007), .B(n24008), .Z(n23993) );
  AND U23766 ( .A(n580), .B(n24009), .Z(n24008) );
  IV U23767 ( .A(n24004), .Z(n24006) );
  XOR U23768 ( .A(n24010), .B(n24011), .Z(n24004) );
  AND U23769 ( .A(n564), .B(n24003), .Z(n24011) );
  XNOR U23770 ( .A(n24001), .B(n24010), .Z(n24003) );
  XNOR U23771 ( .A(n24012), .B(n24013), .Z(n24001) );
  AND U23772 ( .A(n568), .B(n24014), .Z(n24013) );
  XOR U23773 ( .A(p_input[749]), .B(n24012), .Z(n24014) );
  XNOR U23774 ( .A(n24015), .B(n24016), .Z(n24012) );
  AND U23775 ( .A(n572), .B(n24017), .Z(n24016) );
  XOR U23776 ( .A(n24018), .B(n24019), .Z(n24010) );
  AND U23777 ( .A(n576), .B(n24009), .Z(n24019) );
  XNOR U23778 ( .A(n24020), .B(n24007), .Z(n24009) );
  XOR U23779 ( .A(n24021), .B(n24022), .Z(n24007) );
  AND U23780 ( .A(n599), .B(n24023), .Z(n24022) );
  IV U23781 ( .A(n24018), .Z(n24020) );
  XOR U23782 ( .A(n24024), .B(n24025), .Z(n24018) );
  AND U23783 ( .A(n583), .B(n24017), .Z(n24025) );
  XNOR U23784 ( .A(n24015), .B(n24024), .Z(n24017) );
  XNOR U23785 ( .A(n24026), .B(n24027), .Z(n24015) );
  AND U23786 ( .A(n587), .B(n24028), .Z(n24027) );
  XOR U23787 ( .A(p_input[781]), .B(n24026), .Z(n24028) );
  XNOR U23788 ( .A(n24029), .B(n24030), .Z(n24026) );
  AND U23789 ( .A(n591), .B(n24031), .Z(n24030) );
  XOR U23790 ( .A(n24032), .B(n24033), .Z(n24024) );
  AND U23791 ( .A(n595), .B(n24023), .Z(n24033) );
  XNOR U23792 ( .A(n24034), .B(n24021), .Z(n24023) );
  XOR U23793 ( .A(n24035), .B(n24036), .Z(n24021) );
  AND U23794 ( .A(n618), .B(n24037), .Z(n24036) );
  IV U23795 ( .A(n24032), .Z(n24034) );
  XOR U23796 ( .A(n24038), .B(n24039), .Z(n24032) );
  AND U23797 ( .A(n602), .B(n24031), .Z(n24039) );
  XNOR U23798 ( .A(n24029), .B(n24038), .Z(n24031) );
  XNOR U23799 ( .A(n24040), .B(n24041), .Z(n24029) );
  AND U23800 ( .A(n606), .B(n24042), .Z(n24041) );
  XOR U23801 ( .A(p_input[813]), .B(n24040), .Z(n24042) );
  XNOR U23802 ( .A(n24043), .B(n24044), .Z(n24040) );
  AND U23803 ( .A(n610), .B(n24045), .Z(n24044) );
  XOR U23804 ( .A(n24046), .B(n24047), .Z(n24038) );
  AND U23805 ( .A(n614), .B(n24037), .Z(n24047) );
  XNOR U23806 ( .A(n24048), .B(n24035), .Z(n24037) );
  XOR U23807 ( .A(n24049), .B(n24050), .Z(n24035) );
  AND U23808 ( .A(n637), .B(n24051), .Z(n24050) );
  IV U23809 ( .A(n24046), .Z(n24048) );
  XOR U23810 ( .A(n24052), .B(n24053), .Z(n24046) );
  AND U23811 ( .A(n621), .B(n24045), .Z(n24053) );
  XNOR U23812 ( .A(n24043), .B(n24052), .Z(n24045) );
  XNOR U23813 ( .A(n24054), .B(n24055), .Z(n24043) );
  AND U23814 ( .A(n625), .B(n24056), .Z(n24055) );
  XOR U23815 ( .A(p_input[845]), .B(n24054), .Z(n24056) );
  XNOR U23816 ( .A(n24057), .B(n24058), .Z(n24054) );
  AND U23817 ( .A(n629), .B(n24059), .Z(n24058) );
  XOR U23818 ( .A(n24060), .B(n24061), .Z(n24052) );
  AND U23819 ( .A(n633), .B(n24051), .Z(n24061) );
  XNOR U23820 ( .A(n24062), .B(n24049), .Z(n24051) );
  XOR U23821 ( .A(n24063), .B(n24064), .Z(n24049) );
  AND U23822 ( .A(n656), .B(n24065), .Z(n24064) );
  IV U23823 ( .A(n24060), .Z(n24062) );
  XOR U23824 ( .A(n24066), .B(n24067), .Z(n24060) );
  AND U23825 ( .A(n640), .B(n24059), .Z(n24067) );
  XNOR U23826 ( .A(n24057), .B(n24066), .Z(n24059) );
  XNOR U23827 ( .A(n24068), .B(n24069), .Z(n24057) );
  AND U23828 ( .A(n644), .B(n24070), .Z(n24069) );
  XOR U23829 ( .A(p_input[877]), .B(n24068), .Z(n24070) );
  XNOR U23830 ( .A(n24071), .B(n24072), .Z(n24068) );
  AND U23831 ( .A(n648), .B(n24073), .Z(n24072) );
  XOR U23832 ( .A(n24074), .B(n24075), .Z(n24066) );
  AND U23833 ( .A(n652), .B(n24065), .Z(n24075) );
  XNOR U23834 ( .A(n24076), .B(n24063), .Z(n24065) );
  XOR U23835 ( .A(n24077), .B(n24078), .Z(n24063) );
  AND U23836 ( .A(n675), .B(n24079), .Z(n24078) );
  IV U23837 ( .A(n24074), .Z(n24076) );
  XOR U23838 ( .A(n24080), .B(n24081), .Z(n24074) );
  AND U23839 ( .A(n659), .B(n24073), .Z(n24081) );
  XNOR U23840 ( .A(n24071), .B(n24080), .Z(n24073) );
  XNOR U23841 ( .A(n24082), .B(n24083), .Z(n24071) );
  AND U23842 ( .A(n663), .B(n24084), .Z(n24083) );
  XOR U23843 ( .A(p_input[909]), .B(n24082), .Z(n24084) );
  XNOR U23844 ( .A(n24085), .B(n24086), .Z(n24082) );
  AND U23845 ( .A(n667), .B(n24087), .Z(n24086) );
  XOR U23846 ( .A(n24088), .B(n24089), .Z(n24080) );
  AND U23847 ( .A(n671), .B(n24079), .Z(n24089) );
  XNOR U23848 ( .A(n24090), .B(n24077), .Z(n24079) );
  XOR U23849 ( .A(n24091), .B(n24092), .Z(n24077) );
  AND U23850 ( .A(n694), .B(n24093), .Z(n24092) );
  IV U23851 ( .A(n24088), .Z(n24090) );
  XOR U23852 ( .A(n24094), .B(n24095), .Z(n24088) );
  AND U23853 ( .A(n678), .B(n24087), .Z(n24095) );
  XNOR U23854 ( .A(n24085), .B(n24094), .Z(n24087) );
  XNOR U23855 ( .A(n24096), .B(n24097), .Z(n24085) );
  AND U23856 ( .A(n682), .B(n24098), .Z(n24097) );
  XOR U23857 ( .A(p_input[941]), .B(n24096), .Z(n24098) );
  XNOR U23858 ( .A(n24099), .B(n24100), .Z(n24096) );
  AND U23859 ( .A(n686), .B(n24101), .Z(n24100) );
  XOR U23860 ( .A(n24102), .B(n24103), .Z(n24094) );
  AND U23861 ( .A(n690), .B(n24093), .Z(n24103) );
  XNOR U23862 ( .A(n24104), .B(n24091), .Z(n24093) );
  XOR U23863 ( .A(n24105), .B(n24106), .Z(n24091) );
  AND U23864 ( .A(n713), .B(n24107), .Z(n24106) );
  IV U23865 ( .A(n24102), .Z(n24104) );
  XOR U23866 ( .A(n24108), .B(n24109), .Z(n24102) );
  AND U23867 ( .A(n697), .B(n24101), .Z(n24109) );
  XNOR U23868 ( .A(n24099), .B(n24108), .Z(n24101) );
  XNOR U23869 ( .A(n24110), .B(n24111), .Z(n24099) );
  AND U23870 ( .A(n701), .B(n24112), .Z(n24111) );
  XOR U23871 ( .A(p_input[973]), .B(n24110), .Z(n24112) );
  XNOR U23872 ( .A(n24113), .B(n24114), .Z(n24110) );
  AND U23873 ( .A(n705), .B(n24115), .Z(n24114) );
  XOR U23874 ( .A(n24116), .B(n24117), .Z(n24108) );
  AND U23875 ( .A(n709), .B(n24107), .Z(n24117) );
  XNOR U23876 ( .A(n24118), .B(n24105), .Z(n24107) );
  XOR U23877 ( .A(n24119), .B(n24120), .Z(n24105) );
  AND U23878 ( .A(n732), .B(n24121), .Z(n24120) );
  IV U23879 ( .A(n24116), .Z(n24118) );
  XOR U23880 ( .A(n24122), .B(n24123), .Z(n24116) );
  AND U23881 ( .A(n716), .B(n24115), .Z(n24123) );
  XNOR U23882 ( .A(n24113), .B(n24122), .Z(n24115) );
  XNOR U23883 ( .A(n24124), .B(n24125), .Z(n24113) );
  AND U23884 ( .A(n720), .B(n24126), .Z(n24125) );
  XOR U23885 ( .A(p_input[1005]), .B(n24124), .Z(n24126) );
  XNOR U23886 ( .A(n24127), .B(n24128), .Z(n24124) );
  AND U23887 ( .A(n724), .B(n24129), .Z(n24128) );
  XOR U23888 ( .A(n24130), .B(n24131), .Z(n24122) );
  AND U23889 ( .A(n728), .B(n24121), .Z(n24131) );
  XNOR U23890 ( .A(n24132), .B(n24119), .Z(n24121) );
  XOR U23891 ( .A(n24133), .B(n24134), .Z(n24119) );
  AND U23892 ( .A(n751), .B(n24135), .Z(n24134) );
  IV U23893 ( .A(n24130), .Z(n24132) );
  XOR U23894 ( .A(n24136), .B(n24137), .Z(n24130) );
  AND U23895 ( .A(n735), .B(n24129), .Z(n24137) );
  XNOR U23896 ( .A(n24127), .B(n24136), .Z(n24129) );
  XNOR U23897 ( .A(n24138), .B(n24139), .Z(n24127) );
  AND U23898 ( .A(n739), .B(n24140), .Z(n24139) );
  XOR U23899 ( .A(p_input[1037]), .B(n24138), .Z(n24140) );
  XNOR U23900 ( .A(n24141), .B(n24142), .Z(n24138) );
  AND U23901 ( .A(n743), .B(n24143), .Z(n24142) );
  XOR U23902 ( .A(n24144), .B(n24145), .Z(n24136) );
  AND U23903 ( .A(n747), .B(n24135), .Z(n24145) );
  XNOR U23904 ( .A(n24146), .B(n24133), .Z(n24135) );
  XOR U23905 ( .A(n24147), .B(n24148), .Z(n24133) );
  AND U23906 ( .A(n770), .B(n24149), .Z(n24148) );
  IV U23907 ( .A(n24144), .Z(n24146) );
  XOR U23908 ( .A(n24150), .B(n24151), .Z(n24144) );
  AND U23909 ( .A(n754), .B(n24143), .Z(n24151) );
  XNOR U23910 ( .A(n24141), .B(n24150), .Z(n24143) );
  XNOR U23911 ( .A(n24152), .B(n24153), .Z(n24141) );
  AND U23912 ( .A(n758), .B(n24154), .Z(n24153) );
  XOR U23913 ( .A(p_input[1069]), .B(n24152), .Z(n24154) );
  XNOR U23914 ( .A(n24155), .B(n24156), .Z(n24152) );
  AND U23915 ( .A(n762), .B(n24157), .Z(n24156) );
  XOR U23916 ( .A(n24158), .B(n24159), .Z(n24150) );
  AND U23917 ( .A(n766), .B(n24149), .Z(n24159) );
  XNOR U23918 ( .A(n24160), .B(n24147), .Z(n24149) );
  XOR U23919 ( .A(n24161), .B(n24162), .Z(n24147) );
  AND U23920 ( .A(n789), .B(n24163), .Z(n24162) );
  IV U23921 ( .A(n24158), .Z(n24160) );
  XOR U23922 ( .A(n24164), .B(n24165), .Z(n24158) );
  AND U23923 ( .A(n773), .B(n24157), .Z(n24165) );
  XNOR U23924 ( .A(n24155), .B(n24164), .Z(n24157) );
  XNOR U23925 ( .A(n24166), .B(n24167), .Z(n24155) );
  AND U23926 ( .A(n777), .B(n24168), .Z(n24167) );
  XOR U23927 ( .A(p_input[1101]), .B(n24166), .Z(n24168) );
  XNOR U23928 ( .A(n24169), .B(n24170), .Z(n24166) );
  AND U23929 ( .A(n781), .B(n24171), .Z(n24170) );
  XOR U23930 ( .A(n24172), .B(n24173), .Z(n24164) );
  AND U23931 ( .A(n785), .B(n24163), .Z(n24173) );
  XNOR U23932 ( .A(n24174), .B(n24161), .Z(n24163) );
  XOR U23933 ( .A(n24175), .B(n24176), .Z(n24161) );
  AND U23934 ( .A(n808), .B(n24177), .Z(n24176) );
  IV U23935 ( .A(n24172), .Z(n24174) );
  XOR U23936 ( .A(n24178), .B(n24179), .Z(n24172) );
  AND U23937 ( .A(n792), .B(n24171), .Z(n24179) );
  XNOR U23938 ( .A(n24169), .B(n24178), .Z(n24171) );
  XNOR U23939 ( .A(n24180), .B(n24181), .Z(n24169) );
  AND U23940 ( .A(n796), .B(n24182), .Z(n24181) );
  XOR U23941 ( .A(p_input[1133]), .B(n24180), .Z(n24182) );
  XNOR U23942 ( .A(n24183), .B(n24184), .Z(n24180) );
  AND U23943 ( .A(n800), .B(n24185), .Z(n24184) );
  XOR U23944 ( .A(n24186), .B(n24187), .Z(n24178) );
  AND U23945 ( .A(n804), .B(n24177), .Z(n24187) );
  XNOR U23946 ( .A(n24188), .B(n24175), .Z(n24177) );
  XOR U23947 ( .A(n24189), .B(n24190), .Z(n24175) );
  AND U23948 ( .A(n827), .B(n24191), .Z(n24190) );
  IV U23949 ( .A(n24186), .Z(n24188) );
  XOR U23950 ( .A(n24192), .B(n24193), .Z(n24186) );
  AND U23951 ( .A(n811), .B(n24185), .Z(n24193) );
  XNOR U23952 ( .A(n24183), .B(n24192), .Z(n24185) );
  XNOR U23953 ( .A(n24194), .B(n24195), .Z(n24183) );
  AND U23954 ( .A(n815), .B(n24196), .Z(n24195) );
  XOR U23955 ( .A(p_input[1165]), .B(n24194), .Z(n24196) );
  XNOR U23956 ( .A(n24197), .B(n24198), .Z(n24194) );
  AND U23957 ( .A(n819), .B(n24199), .Z(n24198) );
  XOR U23958 ( .A(n24200), .B(n24201), .Z(n24192) );
  AND U23959 ( .A(n823), .B(n24191), .Z(n24201) );
  XNOR U23960 ( .A(n24202), .B(n24189), .Z(n24191) );
  XOR U23961 ( .A(n24203), .B(n24204), .Z(n24189) );
  AND U23962 ( .A(n846), .B(n24205), .Z(n24204) );
  IV U23963 ( .A(n24200), .Z(n24202) );
  XOR U23964 ( .A(n24206), .B(n24207), .Z(n24200) );
  AND U23965 ( .A(n830), .B(n24199), .Z(n24207) );
  XNOR U23966 ( .A(n24197), .B(n24206), .Z(n24199) );
  XNOR U23967 ( .A(n24208), .B(n24209), .Z(n24197) );
  AND U23968 ( .A(n834), .B(n24210), .Z(n24209) );
  XOR U23969 ( .A(p_input[1197]), .B(n24208), .Z(n24210) );
  XNOR U23970 ( .A(n24211), .B(n24212), .Z(n24208) );
  AND U23971 ( .A(n838), .B(n24213), .Z(n24212) );
  XOR U23972 ( .A(n24214), .B(n24215), .Z(n24206) );
  AND U23973 ( .A(n842), .B(n24205), .Z(n24215) );
  XNOR U23974 ( .A(n24216), .B(n24203), .Z(n24205) );
  XOR U23975 ( .A(n24217), .B(n24218), .Z(n24203) );
  AND U23976 ( .A(n865), .B(n24219), .Z(n24218) );
  IV U23977 ( .A(n24214), .Z(n24216) );
  XOR U23978 ( .A(n24220), .B(n24221), .Z(n24214) );
  AND U23979 ( .A(n849), .B(n24213), .Z(n24221) );
  XNOR U23980 ( .A(n24211), .B(n24220), .Z(n24213) );
  XNOR U23981 ( .A(n24222), .B(n24223), .Z(n24211) );
  AND U23982 ( .A(n853), .B(n24224), .Z(n24223) );
  XOR U23983 ( .A(p_input[1229]), .B(n24222), .Z(n24224) );
  XNOR U23984 ( .A(n24225), .B(n24226), .Z(n24222) );
  AND U23985 ( .A(n857), .B(n24227), .Z(n24226) );
  XOR U23986 ( .A(n24228), .B(n24229), .Z(n24220) );
  AND U23987 ( .A(n861), .B(n24219), .Z(n24229) );
  XNOR U23988 ( .A(n24230), .B(n24217), .Z(n24219) );
  XOR U23989 ( .A(n24231), .B(n24232), .Z(n24217) );
  AND U23990 ( .A(n884), .B(n24233), .Z(n24232) );
  IV U23991 ( .A(n24228), .Z(n24230) );
  XOR U23992 ( .A(n24234), .B(n24235), .Z(n24228) );
  AND U23993 ( .A(n868), .B(n24227), .Z(n24235) );
  XNOR U23994 ( .A(n24225), .B(n24234), .Z(n24227) );
  XNOR U23995 ( .A(n24236), .B(n24237), .Z(n24225) );
  AND U23996 ( .A(n872), .B(n24238), .Z(n24237) );
  XOR U23997 ( .A(p_input[1261]), .B(n24236), .Z(n24238) );
  XNOR U23998 ( .A(n24239), .B(n24240), .Z(n24236) );
  AND U23999 ( .A(n876), .B(n24241), .Z(n24240) );
  XOR U24000 ( .A(n24242), .B(n24243), .Z(n24234) );
  AND U24001 ( .A(n880), .B(n24233), .Z(n24243) );
  XNOR U24002 ( .A(n24244), .B(n24231), .Z(n24233) );
  XOR U24003 ( .A(n24245), .B(n24246), .Z(n24231) );
  AND U24004 ( .A(n903), .B(n24247), .Z(n24246) );
  IV U24005 ( .A(n24242), .Z(n24244) );
  XOR U24006 ( .A(n24248), .B(n24249), .Z(n24242) );
  AND U24007 ( .A(n887), .B(n24241), .Z(n24249) );
  XNOR U24008 ( .A(n24239), .B(n24248), .Z(n24241) );
  XNOR U24009 ( .A(n24250), .B(n24251), .Z(n24239) );
  AND U24010 ( .A(n891), .B(n24252), .Z(n24251) );
  XOR U24011 ( .A(p_input[1293]), .B(n24250), .Z(n24252) );
  XNOR U24012 ( .A(n24253), .B(n24254), .Z(n24250) );
  AND U24013 ( .A(n895), .B(n24255), .Z(n24254) );
  XOR U24014 ( .A(n24256), .B(n24257), .Z(n24248) );
  AND U24015 ( .A(n899), .B(n24247), .Z(n24257) );
  XNOR U24016 ( .A(n24258), .B(n24245), .Z(n24247) );
  XOR U24017 ( .A(n24259), .B(n24260), .Z(n24245) );
  AND U24018 ( .A(n922), .B(n24261), .Z(n24260) );
  IV U24019 ( .A(n24256), .Z(n24258) );
  XOR U24020 ( .A(n24262), .B(n24263), .Z(n24256) );
  AND U24021 ( .A(n906), .B(n24255), .Z(n24263) );
  XNOR U24022 ( .A(n24253), .B(n24262), .Z(n24255) );
  XNOR U24023 ( .A(n24264), .B(n24265), .Z(n24253) );
  AND U24024 ( .A(n910), .B(n24266), .Z(n24265) );
  XOR U24025 ( .A(p_input[1325]), .B(n24264), .Z(n24266) );
  XNOR U24026 ( .A(n24267), .B(n24268), .Z(n24264) );
  AND U24027 ( .A(n914), .B(n24269), .Z(n24268) );
  XOR U24028 ( .A(n24270), .B(n24271), .Z(n24262) );
  AND U24029 ( .A(n918), .B(n24261), .Z(n24271) );
  XNOR U24030 ( .A(n24272), .B(n24259), .Z(n24261) );
  XOR U24031 ( .A(n24273), .B(n24274), .Z(n24259) );
  AND U24032 ( .A(n941), .B(n24275), .Z(n24274) );
  IV U24033 ( .A(n24270), .Z(n24272) );
  XOR U24034 ( .A(n24276), .B(n24277), .Z(n24270) );
  AND U24035 ( .A(n925), .B(n24269), .Z(n24277) );
  XNOR U24036 ( .A(n24267), .B(n24276), .Z(n24269) );
  XNOR U24037 ( .A(n24278), .B(n24279), .Z(n24267) );
  AND U24038 ( .A(n929), .B(n24280), .Z(n24279) );
  XOR U24039 ( .A(p_input[1357]), .B(n24278), .Z(n24280) );
  XNOR U24040 ( .A(n24281), .B(n24282), .Z(n24278) );
  AND U24041 ( .A(n933), .B(n24283), .Z(n24282) );
  XOR U24042 ( .A(n24284), .B(n24285), .Z(n24276) );
  AND U24043 ( .A(n937), .B(n24275), .Z(n24285) );
  XNOR U24044 ( .A(n24286), .B(n24273), .Z(n24275) );
  XOR U24045 ( .A(n24287), .B(n24288), .Z(n24273) );
  AND U24046 ( .A(n960), .B(n24289), .Z(n24288) );
  IV U24047 ( .A(n24284), .Z(n24286) );
  XOR U24048 ( .A(n24290), .B(n24291), .Z(n24284) );
  AND U24049 ( .A(n944), .B(n24283), .Z(n24291) );
  XNOR U24050 ( .A(n24281), .B(n24290), .Z(n24283) );
  XNOR U24051 ( .A(n24292), .B(n24293), .Z(n24281) );
  AND U24052 ( .A(n948), .B(n24294), .Z(n24293) );
  XOR U24053 ( .A(p_input[1389]), .B(n24292), .Z(n24294) );
  XNOR U24054 ( .A(n24295), .B(n24296), .Z(n24292) );
  AND U24055 ( .A(n952), .B(n24297), .Z(n24296) );
  XOR U24056 ( .A(n24298), .B(n24299), .Z(n24290) );
  AND U24057 ( .A(n956), .B(n24289), .Z(n24299) );
  XNOR U24058 ( .A(n24300), .B(n24287), .Z(n24289) );
  XOR U24059 ( .A(n24301), .B(n24302), .Z(n24287) );
  AND U24060 ( .A(n979), .B(n24303), .Z(n24302) );
  IV U24061 ( .A(n24298), .Z(n24300) );
  XOR U24062 ( .A(n24304), .B(n24305), .Z(n24298) );
  AND U24063 ( .A(n963), .B(n24297), .Z(n24305) );
  XNOR U24064 ( .A(n24295), .B(n24304), .Z(n24297) );
  XNOR U24065 ( .A(n24306), .B(n24307), .Z(n24295) );
  AND U24066 ( .A(n967), .B(n24308), .Z(n24307) );
  XOR U24067 ( .A(p_input[1421]), .B(n24306), .Z(n24308) );
  XNOR U24068 ( .A(n24309), .B(n24310), .Z(n24306) );
  AND U24069 ( .A(n971), .B(n24311), .Z(n24310) );
  XOR U24070 ( .A(n24312), .B(n24313), .Z(n24304) );
  AND U24071 ( .A(n975), .B(n24303), .Z(n24313) );
  XNOR U24072 ( .A(n24314), .B(n24301), .Z(n24303) );
  XOR U24073 ( .A(n24315), .B(n24316), .Z(n24301) );
  AND U24074 ( .A(n998), .B(n24317), .Z(n24316) );
  IV U24075 ( .A(n24312), .Z(n24314) );
  XOR U24076 ( .A(n24318), .B(n24319), .Z(n24312) );
  AND U24077 ( .A(n982), .B(n24311), .Z(n24319) );
  XNOR U24078 ( .A(n24309), .B(n24318), .Z(n24311) );
  XNOR U24079 ( .A(n24320), .B(n24321), .Z(n24309) );
  AND U24080 ( .A(n986), .B(n24322), .Z(n24321) );
  XOR U24081 ( .A(p_input[1453]), .B(n24320), .Z(n24322) );
  XNOR U24082 ( .A(n24323), .B(n24324), .Z(n24320) );
  AND U24083 ( .A(n990), .B(n24325), .Z(n24324) );
  XOR U24084 ( .A(n24326), .B(n24327), .Z(n24318) );
  AND U24085 ( .A(n994), .B(n24317), .Z(n24327) );
  XNOR U24086 ( .A(n24328), .B(n24315), .Z(n24317) );
  XOR U24087 ( .A(n24329), .B(n24330), .Z(n24315) );
  AND U24088 ( .A(n1017), .B(n24331), .Z(n24330) );
  IV U24089 ( .A(n24326), .Z(n24328) );
  XOR U24090 ( .A(n24332), .B(n24333), .Z(n24326) );
  AND U24091 ( .A(n1001), .B(n24325), .Z(n24333) );
  XNOR U24092 ( .A(n24323), .B(n24332), .Z(n24325) );
  XNOR U24093 ( .A(n24334), .B(n24335), .Z(n24323) );
  AND U24094 ( .A(n1005), .B(n24336), .Z(n24335) );
  XOR U24095 ( .A(p_input[1485]), .B(n24334), .Z(n24336) );
  XNOR U24096 ( .A(n24337), .B(n24338), .Z(n24334) );
  AND U24097 ( .A(n1009), .B(n24339), .Z(n24338) );
  XOR U24098 ( .A(n24340), .B(n24341), .Z(n24332) );
  AND U24099 ( .A(n1013), .B(n24331), .Z(n24341) );
  XNOR U24100 ( .A(n24342), .B(n24329), .Z(n24331) );
  XOR U24101 ( .A(n24343), .B(n24344), .Z(n24329) );
  AND U24102 ( .A(n1036), .B(n24345), .Z(n24344) );
  IV U24103 ( .A(n24340), .Z(n24342) );
  XOR U24104 ( .A(n24346), .B(n24347), .Z(n24340) );
  AND U24105 ( .A(n1020), .B(n24339), .Z(n24347) );
  XNOR U24106 ( .A(n24337), .B(n24346), .Z(n24339) );
  XNOR U24107 ( .A(n24348), .B(n24349), .Z(n24337) );
  AND U24108 ( .A(n1024), .B(n24350), .Z(n24349) );
  XOR U24109 ( .A(p_input[1517]), .B(n24348), .Z(n24350) );
  XNOR U24110 ( .A(n24351), .B(n24352), .Z(n24348) );
  AND U24111 ( .A(n1028), .B(n24353), .Z(n24352) );
  XOR U24112 ( .A(n24354), .B(n24355), .Z(n24346) );
  AND U24113 ( .A(n1032), .B(n24345), .Z(n24355) );
  XNOR U24114 ( .A(n24356), .B(n24343), .Z(n24345) );
  XOR U24115 ( .A(n24357), .B(n24358), .Z(n24343) );
  AND U24116 ( .A(n1055), .B(n24359), .Z(n24358) );
  IV U24117 ( .A(n24354), .Z(n24356) );
  XOR U24118 ( .A(n24360), .B(n24361), .Z(n24354) );
  AND U24119 ( .A(n1039), .B(n24353), .Z(n24361) );
  XNOR U24120 ( .A(n24351), .B(n24360), .Z(n24353) );
  XNOR U24121 ( .A(n24362), .B(n24363), .Z(n24351) );
  AND U24122 ( .A(n1043), .B(n24364), .Z(n24363) );
  XOR U24123 ( .A(p_input[1549]), .B(n24362), .Z(n24364) );
  XNOR U24124 ( .A(n24365), .B(n24366), .Z(n24362) );
  AND U24125 ( .A(n1047), .B(n24367), .Z(n24366) );
  XOR U24126 ( .A(n24368), .B(n24369), .Z(n24360) );
  AND U24127 ( .A(n1051), .B(n24359), .Z(n24369) );
  XNOR U24128 ( .A(n24370), .B(n24357), .Z(n24359) );
  XOR U24129 ( .A(n24371), .B(n24372), .Z(n24357) );
  AND U24130 ( .A(n1074), .B(n24373), .Z(n24372) );
  IV U24131 ( .A(n24368), .Z(n24370) );
  XOR U24132 ( .A(n24374), .B(n24375), .Z(n24368) );
  AND U24133 ( .A(n1058), .B(n24367), .Z(n24375) );
  XNOR U24134 ( .A(n24365), .B(n24374), .Z(n24367) );
  XNOR U24135 ( .A(n24376), .B(n24377), .Z(n24365) );
  AND U24136 ( .A(n1062), .B(n24378), .Z(n24377) );
  XOR U24137 ( .A(p_input[1581]), .B(n24376), .Z(n24378) );
  XNOR U24138 ( .A(n24379), .B(n24380), .Z(n24376) );
  AND U24139 ( .A(n1066), .B(n24381), .Z(n24380) );
  XOR U24140 ( .A(n24382), .B(n24383), .Z(n24374) );
  AND U24141 ( .A(n1070), .B(n24373), .Z(n24383) );
  XNOR U24142 ( .A(n24384), .B(n24371), .Z(n24373) );
  XOR U24143 ( .A(n24385), .B(n24386), .Z(n24371) );
  AND U24144 ( .A(n1093), .B(n24387), .Z(n24386) );
  IV U24145 ( .A(n24382), .Z(n24384) );
  XOR U24146 ( .A(n24388), .B(n24389), .Z(n24382) );
  AND U24147 ( .A(n1077), .B(n24381), .Z(n24389) );
  XNOR U24148 ( .A(n24379), .B(n24388), .Z(n24381) );
  XNOR U24149 ( .A(n24390), .B(n24391), .Z(n24379) );
  AND U24150 ( .A(n1081), .B(n24392), .Z(n24391) );
  XOR U24151 ( .A(p_input[1613]), .B(n24390), .Z(n24392) );
  XNOR U24152 ( .A(n24393), .B(n24394), .Z(n24390) );
  AND U24153 ( .A(n1085), .B(n24395), .Z(n24394) );
  XOR U24154 ( .A(n24396), .B(n24397), .Z(n24388) );
  AND U24155 ( .A(n1089), .B(n24387), .Z(n24397) );
  XNOR U24156 ( .A(n24398), .B(n24385), .Z(n24387) );
  XOR U24157 ( .A(n24399), .B(n24400), .Z(n24385) );
  AND U24158 ( .A(n1112), .B(n24401), .Z(n24400) );
  IV U24159 ( .A(n24396), .Z(n24398) );
  XOR U24160 ( .A(n24402), .B(n24403), .Z(n24396) );
  AND U24161 ( .A(n1096), .B(n24395), .Z(n24403) );
  XNOR U24162 ( .A(n24393), .B(n24402), .Z(n24395) );
  XNOR U24163 ( .A(n24404), .B(n24405), .Z(n24393) );
  AND U24164 ( .A(n1100), .B(n24406), .Z(n24405) );
  XOR U24165 ( .A(p_input[1645]), .B(n24404), .Z(n24406) );
  XNOR U24166 ( .A(n24407), .B(n24408), .Z(n24404) );
  AND U24167 ( .A(n1104), .B(n24409), .Z(n24408) );
  XOR U24168 ( .A(n24410), .B(n24411), .Z(n24402) );
  AND U24169 ( .A(n1108), .B(n24401), .Z(n24411) );
  XNOR U24170 ( .A(n24412), .B(n24399), .Z(n24401) );
  XOR U24171 ( .A(n24413), .B(n24414), .Z(n24399) );
  AND U24172 ( .A(n1131), .B(n24415), .Z(n24414) );
  IV U24173 ( .A(n24410), .Z(n24412) );
  XOR U24174 ( .A(n24416), .B(n24417), .Z(n24410) );
  AND U24175 ( .A(n1115), .B(n24409), .Z(n24417) );
  XNOR U24176 ( .A(n24407), .B(n24416), .Z(n24409) );
  XNOR U24177 ( .A(n24418), .B(n24419), .Z(n24407) );
  AND U24178 ( .A(n1119), .B(n24420), .Z(n24419) );
  XOR U24179 ( .A(p_input[1677]), .B(n24418), .Z(n24420) );
  XNOR U24180 ( .A(n24421), .B(n24422), .Z(n24418) );
  AND U24181 ( .A(n1123), .B(n24423), .Z(n24422) );
  XOR U24182 ( .A(n24424), .B(n24425), .Z(n24416) );
  AND U24183 ( .A(n1127), .B(n24415), .Z(n24425) );
  XNOR U24184 ( .A(n24426), .B(n24413), .Z(n24415) );
  XOR U24185 ( .A(n24427), .B(n24428), .Z(n24413) );
  AND U24186 ( .A(n1150), .B(n24429), .Z(n24428) );
  IV U24187 ( .A(n24424), .Z(n24426) );
  XOR U24188 ( .A(n24430), .B(n24431), .Z(n24424) );
  AND U24189 ( .A(n1134), .B(n24423), .Z(n24431) );
  XNOR U24190 ( .A(n24421), .B(n24430), .Z(n24423) );
  XNOR U24191 ( .A(n24432), .B(n24433), .Z(n24421) );
  AND U24192 ( .A(n1138), .B(n24434), .Z(n24433) );
  XOR U24193 ( .A(p_input[1709]), .B(n24432), .Z(n24434) );
  XNOR U24194 ( .A(n24435), .B(n24436), .Z(n24432) );
  AND U24195 ( .A(n1142), .B(n24437), .Z(n24436) );
  XOR U24196 ( .A(n24438), .B(n24439), .Z(n24430) );
  AND U24197 ( .A(n1146), .B(n24429), .Z(n24439) );
  XNOR U24198 ( .A(n24440), .B(n24427), .Z(n24429) );
  XOR U24199 ( .A(n24441), .B(n24442), .Z(n24427) );
  AND U24200 ( .A(n1169), .B(n24443), .Z(n24442) );
  IV U24201 ( .A(n24438), .Z(n24440) );
  XOR U24202 ( .A(n24444), .B(n24445), .Z(n24438) );
  AND U24203 ( .A(n1153), .B(n24437), .Z(n24445) );
  XNOR U24204 ( .A(n24435), .B(n24444), .Z(n24437) );
  XNOR U24205 ( .A(n24446), .B(n24447), .Z(n24435) );
  AND U24206 ( .A(n1157), .B(n24448), .Z(n24447) );
  XOR U24207 ( .A(p_input[1741]), .B(n24446), .Z(n24448) );
  XNOR U24208 ( .A(n24449), .B(n24450), .Z(n24446) );
  AND U24209 ( .A(n1161), .B(n24451), .Z(n24450) );
  XOR U24210 ( .A(n24452), .B(n24453), .Z(n24444) );
  AND U24211 ( .A(n1165), .B(n24443), .Z(n24453) );
  XNOR U24212 ( .A(n24454), .B(n24441), .Z(n24443) );
  XOR U24213 ( .A(n24455), .B(n24456), .Z(n24441) );
  AND U24214 ( .A(n1188), .B(n24457), .Z(n24456) );
  IV U24215 ( .A(n24452), .Z(n24454) );
  XOR U24216 ( .A(n24458), .B(n24459), .Z(n24452) );
  AND U24217 ( .A(n1172), .B(n24451), .Z(n24459) );
  XNOR U24218 ( .A(n24449), .B(n24458), .Z(n24451) );
  XNOR U24219 ( .A(n24460), .B(n24461), .Z(n24449) );
  AND U24220 ( .A(n1176), .B(n24462), .Z(n24461) );
  XOR U24221 ( .A(p_input[1773]), .B(n24460), .Z(n24462) );
  XNOR U24222 ( .A(n24463), .B(n24464), .Z(n24460) );
  AND U24223 ( .A(n1180), .B(n24465), .Z(n24464) );
  XOR U24224 ( .A(n24466), .B(n24467), .Z(n24458) );
  AND U24225 ( .A(n1184), .B(n24457), .Z(n24467) );
  XNOR U24226 ( .A(n24468), .B(n24455), .Z(n24457) );
  XOR U24227 ( .A(n24469), .B(n24470), .Z(n24455) );
  AND U24228 ( .A(n1207), .B(n24471), .Z(n24470) );
  IV U24229 ( .A(n24466), .Z(n24468) );
  XOR U24230 ( .A(n24472), .B(n24473), .Z(n24466) );
  AND U24231 ( .A(n1191), .B(n24465), .Z(n24473) );
  XNOR U24232 ( .A(n24463), .B(n24472), .Z(n24465) );
  XNOR U24233 ( .A(n24474), .B(n24475), .Z(n24463) );
  AND U24234 ( .A(n1195), .B(n24476), .Z(n24475) );
  XOR U24235 ( .A(p_input[1805]), .B(n24474), .Z(n24476) );
  XNOR U24236 ( .A(n24477), .B(n24478), .Z(n24474) );
  AND U24237 ( .A(n1199), .B(n24479), .Z(n24478) );
  XOR U24238 ( .A(n24480), .B(n24481), .Z(n24472) );
  AND U24239 ( .A(n1203), .B(n24471), .Z(n24481) );
  XNOR U24240 ( .A(n24482), .B(n24469), .Z(n24471) );
  XOR U24241 ( .A(n24483), .B(n24484), .Z(n24469) );
  AND U24242 ( .A(n1226), .B(n24485), .Z(n24484) );
  IV U24243 ( .A(n24480), .Z(n24482) );
  XOR U24244 ( .A(n24486), .B(n24487), .Z(n24480) );
  AND U24245 ( .A(n1210), .B(n24479), .Z(n24487) );
  XNOR U24246 ( .A(n24477), .B(n24486), .Z(n24479) );
  XNOR U24247 ( .A(n24488), .B(n24489), .Z(n24477) );
  AND U24248 ( .A(n1214), .B(n24490), .Z(n24489) );
  XOR U24249 ( .A(p_input[1837]), .B(n24488), .Z(n24490) );
  XNOR U24250 ( .A(n24491), .B(n24492), .Z(n24488) );
  AND U24251 ( .A(n1218), .B(n24493), .Z(n24492) );
  XOR U24252 ( .A(n24494), .B(n24495), .Z(n24486) );
  AND U24253 ( .A(n1222), .B(n24485), .Z(n24495) );
  XNOR U24254 ( .A(n24496), .B(n24483), .Z(n24485) );
  XOR U24255 ( .A(n24497), .B(n24498), .Z(n24483) );
  AND U24256 ( .A(n1245), .B(n24499), .Z(n24498) );
  IV U24257 ( .A(n24494), .Z(n24496) );
  XOR U24258 ( .A(n24500), .B(n24501), .Z(n24494) );
  AND U24259 ( .A(n1229), .B(n24493), .Z(n24501) );
  XNOR U24260 ( .A(n24491), .B(n24500), .Z(n24493) );
  XNOR U24261 ( .A(n24502), .B(n24503), .Z(n24491) );
  AND U24262 ( .A(n1233), .B(n24504), .Z(n24503) );
  XOR U24263 ( .A(p_input[1869]), .B(n24502), .Z(n24504) );
  XNOR U24264 ( .A(n24505), .B(n24506), .Z(n24502) );
  AND U24265 ( .A(n1237), .B(n24507), .Z(n24506) );
  XOR U24266 ( .A(n24508), .B(n24509), .Z(n24500) );
  AND U24267 ( .A(n1241), .B(n24499), .Z(n24509) );
  XNOR U24268 ( .A(n24510), .B(n24497), .Z(n24499) );
  XOR U24269 ( .A(n24511), .B(n24512), .Z(n24497) );
  AND U24270 ( .A(n1264), .B(n24513), .Z(n24512) );
  IV U24271 ( .A(n24508), .Z(n24510) );
  XOR U24272 ( .A(n24514), .B(n24515), .Z(n24508) );
  AND U24273 ( .A(n1248), .B(n24507), .Z(n24515) );
  XNOR U24274 ( .A(n24505), .B(n24514), .Z(n24507) );
  XNOR U24275 ( .A(n24516), .B(n24517), .Z(n24505) );
  AND U24276 ( .A(n1252), .B(n24518), .Z(n24517) );
  XOR U24277 ( .A(p_input[1901]), .B(n24516), .Z(n24518) );
  XNOR U24278 ( .A(n24519), .B(n24520), .Z(n24516) );
  AND U24279 ( .A(n1256), .B(n24521), .Z(n24520) );
  XOR U24280 ( .A(n24522), .B(n24523), .Z(n24514) );
  AND U24281 ( .A(n1260), .B(n24513), .Z(n24523) );
  XNOR U24282 ( .A(n24524), .B(n24511), .Z(n24513) );
  XOR U24283 ( .A(n24525), .B(n24526), .Z(n24511) );
  AND U24284 ( .A(n1282), .B(n24527), .Z(n24526) );
  IV U24285 ( .A(n24522), .Z(n24524) );
  XOR U24286 ( .A(n24528), .B(n24529), .Z(n24522) );
  AND U24287 ( .A(n1267), .B(n24521), .Z(n24529) );
  XNOR U24288 ( .A(n24519), .B(n24528), .Z(n24521) );
  XNOR U24289 ( .A(n24530), .B(n24531), .Z(n24519) );
  AND U24290 ( .A(n1271), .B(n24532), .Z(n24531) );
  XOR U24291 ( .A(p_input[1933]), .B(n24530), .Z(n24532) );
  XOR U24292 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(n24533), 
        .Z(n24530) );
  AND U24293 ( .A(n1274), .B(n24534), .Z(n24533) );
  XOR U24294 ( .A(n24535), .B(n24536), .Z(n24528) );
  AND U24295 ( .A(n1278), .B(n24527), .Z(n24536) );
  XNOR U24296 ( .A(n24537), .B(n24525), .Z(n24527) );
  XOR U24297 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n24538), .Z(n24525) );
  AND U24298 ( .A(n1290), .B(n24539), .Z(n24538) );
  IV U24299 ( .A(n24535), .Z(n24537) );
  XOR U24300 ( .A(n24540), .B(n24541), .Z(n24535) );
  AND U24301 ( .A(n1285), .B(n24534), .Z(n24541) );
  XOR U24302 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(n24540), 
        .Z(n24534) );
  XOR U24303 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(n24542), 
        .Z(n24540) );
  AND U24304 ( .A(n1287), .B(n24539), .Z(n24542) );
  XOR U24305 ( .A(\knn_comb_/min_val_out[0][13] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n24539) );
  XOR U24306 ( .A(n115), .B(n24543), .Z(o[12]) );
  AND U24307 ( .A(n122), .B(n24544), .Z(n115) );
  XOR U24308 ( .A(n116), .B(n24543), .Z(n24544) );
  XOR U24309 ( .A(n24545), .B(n24546), .Z(n24543) );
  AND U24310 ( .A(n142), .B(n24547), .Z(n24546) );
  XOR U24311 ( .A(n24548), .B(n45), .Z(n116) );
  AND U24312 ( .A(n125), .B(n24549), .Z(n45) );
  XOR U24313 ( .A(n46), .B(n24548), .Z(n24549) );
  XOR U24314 ( .A(n24550), .B(n24551), .Z(n46) );
  AND U24315 ( .A(n130), .B(n24552), .Z(n24551) );
  XOR U24316 ( .A(p_input[12]), .B(n24550), .Z(n24552) );
  XNOR U24317 ( .A(n24553), .B(n24554), .Z(n24550) );
  AND U24318 ( .A(n134), .B(n24555), .Z(n24554) );
  XOR U24319 ( .A(n24556), .B(n24557), .Z(n24548) );
  AND U24320 ( .A(n138), .B(n24547), .Z(n24557) );
  XNOR U24321 ( .A(n24558), .B(n24545), .Z(n24547) );
  XOR U24322 ( .A(n24559), .B(n24560), .Z(n24545) );
  AND U24323 ( .A(n162), .B(n24561), .Z(n24560) );
  IV U24324 ( .A(n24556), .Z(n24558) );
  XOR U24325 ( .A(n24562), .B(n24563), .Z(n24556) );
  AND U24326 ( .A(n146), .B(n24555), .Z(n24563) );
  XNOR U24327 ( .A(n24553), .B(n24562), .Z(n24555) );
  XNOR U24328 ( .A(n24564), .B(n24565), .Z(n24553) );
  AND U24329 ( .A(n150), .B(n24566), .Z(n24565) );
  XOR U24330 ( .A(p_input[44]), .B(n24564), .Z(n24566) );
  XNOR U24331 ( .A(n24567), .B(n24568), .Z(n24564) );
  AND U24332 ( .A(n154), .B(n24569), .Z(n24568) );
  XOR U24333 ( .A(n24570), .B(n24571), .Z(n24562) );
  AND U24334 ( .A(n158), .B(n24561), .Z(n24571) );
  XNOR U24335 ( .A(n24572), .B(n24559), .Z(n24561) );
  XOR U24336 ( .A(n24573), .B(n24574), .Z(n24559) );
  AND U24337 ( .A(n181), .B(n24575), .Z(n24574) );
  IV U24338 ( .A(n24570), .Z(n24572) );
  XOR U24339 ( .A(n24576), .B(n24577), .Z(n24570) );
  AND U24340 ( .A(n165), .B(n24569), .Z(n24577) );
  XNOR U24341 ( .A(n24567), .B(n24576), .Z(n24569) );
  XNOR U24342 ( .A(n24578), .B(n24579), .Z(n24567) );
  AND U24343 ( .A(n169), .B(n24580), .Z(n24579) );
  XOR U24344 ( .A(p_input[76]), .B(n24578), .Z(n24580) );
  XNOR U24345 ( .A(n24581), .B(n24582), .Z(n24578) );
  AND U24346 ( .A(n173), .B(n24583), .Z(n24582) );
  XOR U24347 ( .A(n24584), .B(n24585), .Z(n24576) );
  AND U24348 ( .A(n177), .B(n24575), .Z(n24585) );
  XNOR U24349 ( .A(n24586), .B(n24573), .Z(n24575) );
  XOR U24350 ( .A(n24587), .B(n24588), .Z(n24573) );
  AND U24351 ( .A(n200), .B(n24589), .Z(n24588) );
  IV U24352 ( .A(n24584), .Z(n24586) );
  XOR U24353 ( .A(n24590), .B(n24591), .Z(n24584) );
  AND U24354 ( .A(n184), .B(n24583), .Z(n24591) );
  XNOR U24355 ( .A(n24581), .B(n24590), .Z(n24583) );
  XNOR U24356 ( .A(n24592), .B(n24593), .Z(n24581) );
  AND U24357 ( .A(n188), .B(n24594), .Z(n24593) );
  XOR U24358 ( .A(p_input[108]), .B(n24592), .Z(n24594) );
  XNOR U24359 ( .A(n24595), .B(n24596), .Z(n24592) );
  AND U24360 ( .A(n192), .B(n24597), .Z(n24596) );
  XOR U24361 ( .A(n24598), .B(n24599), .Z(n24590) );
  AND U24362 ( .A(n196), .B(n24589), .Z(n24599) );
  XNOR U24363 ( .A(n24600), .B(n24587), .Z(n24589) );
  XOR U24364 ( .A(n24601), .B(n24602), .Z(n24587) );
  AND U24365 ( .A(n219), .B(n24603), .Z(n24602) );
  IV U24366 ( .A(n24598), .Z(n24600) );
  XOR U24367 ( .A(n24604), .B(n24605), .Z(n24598) );
  AND U24368 ( .A(n203), .B(n24597), .Z(n24605) );
  XNOR U24369 ( .A(n24595), .B(n24604), .Z(n24597) );
  XNOR U24370 ( .A(n24606), .B(n24607), .Z(n24595) );
  AND U24371 ( .A(n207), .B(n24608), .Z(n24607) );
  XOR U24372 ( .A(p_input[140]), .B(n24606), .Z(n24608) );
  XNOR U24373 ( .A(n24609), .B(n24610), .Z(n24606) );
  AND U24374 ( .A(n211), .B(n24611), .Z(n24610) );
  XOR U24375 ( .A(n24612), .B(n24613), .Z(n24604) );
  AND U24376 ( .A(n215), .B(n24603), .Z(n24613) );
  XNOR U24377 ( .A(n24614), .B(n24601), .Z(n24603) );
  XOR U24378 ( .A(n24615), .B(n24616), .Z(n24601) );
  AND U24379 ( .A(n238), .B(n24617), .Z(n24616) );
  IV U24380 ( .A(n24612), .Z(n24614) );
  XOR U24381 ( .A(n24618), .B(n24619), .Z(n24612) );
  AND U24382 ( .A(n222), .B(n24611), .Z(n24619) );
  XNOR U24383 ( .A(n24609), .B(n24618), .Z(n24611) );
  XNOR U24384 ( .A(n24620), .B(n24621), .Z(n24609) );
  AND U24385 ( .A(n226), .B(n24622), .Z(n24621) );
  XOR U24386 ( .A(p_input[172]), .B(n24620), .Z(n24622) );
  XNOR U24387 ( .A(n24623), .B(n24624), .Z(n24620) );
  AND U24388 ( .A(n230), .B(n24625), .Z(n24624) );
  XOR U24389 ( .A(n24626), .B(n24627), .Z(n24618) );
  AND U24390 ( .A(n234), .B(n24617), .Z(n24627) );
  XNOR U24391 ( .A(n24628), .B(n24615), .Z(n24617) );
  XOR U24392 ( .A(n24629), .B(n24630), .Z(n24615) );
  AND U24393 ( .A(n257), .B(n24631), .Z(n24630) );
  IV U24394 ( .A(n24626), .Z(n24628) );
  XOR U24395 ( .A(n24632), .B(n24633), .Z(n24626) );
  AND U24396 ( .A(n241), .B(n24625), .Z(n24633) );
  XNOR U24397 ( .A(n24623), .B(n24632), .Z(n24625) );
  XNOR U24398 ( .A(n24634), .B(n24635), .Z(n24623) );
  AND U24399 ( .A(n245), .B(n24636), .Z(n24635) );
  XOR U24400 ( .A(p_input[204]), .B(n24634), .Z(n24636) );
  XNOR U24401 ( .A(n24637), .B(n24638), .Z(n24634) );
  AND U24402 ( .A(n249), .B(n24639), .Z(n24638) );
  XOR U24403 ( .A(n24640), .B(n24641), .Z(n24632) );
  AND U24404 ( .A(n253), .B(n24631), .Z(n24641) );
  XNOR U24405 ( .A(n24642), .B(n24629), .Z(n24631) );
  XOR U24406 ( .A(n24643), .B(n24644), .Z(n24629) );
  AND U24407 ( .A(n276), .B(n24645), .Z(n24644) );
  IV U24408 ( .A(n24640), .Z(n24642) );
  XOR U24409 ( .A(n24646), .B(n24647), .Z(n24640) );
  AND U24410 ( .A(n260), .B(n24639), .Z(n24647) );
  XNOR U24411 ( .A(n24637), .B(n24646), .Z(n24639) );
  XNOR U24412 ( .A(n24648), .B(n24649), .Z(n24637) );
  AND U24413 ( .A(n264), .B(n24650), .Z(n24649) );
  XOR U24414 ( .A(p_input[236]), .B(n24648), .Z(n24650) );
  XNOR U24415 ( .A(n24651), .B(n24652), .Z(n24648) );
  AND U24416 ( .A(n268), .B(n24653), .Z(n24652) );
  XOR U24417 ( .A(n24654), .B(n24655), .Z(n24646) );
  AND U24418 ( .A(n272), .B(n24645), .Z(n24655) );
  XNOR U24419 ( .A(n24656), .B(n24643), .Z(n24645) );
  XOR U24420 ( .A(n24657), .B(n24658), .Z(n24643) );
  AND U24421 ( .A(n295), .B(n24659), .Z(n24658) );
  IV U24422 ( .A(n24654), .Z(n24656) );
  XOR U24423 ( .A(n24660), .B(n24661), .Z(n24654) );
  AND U24424 ( .A(n279), .B(n24653), .Z(n24661) );
  XNOR U24425 ( .A(n24651), .B(n24660), .Z(n24653) );
  XNOR U24426 ( .A(n24662), .B(n24663), .Z(n24651) );
  AND U24427 ( .A(n283), .B(n24664), .Z(n24663) );
  XOR U24428 ( .A(p_input[268]), .B(n24662), .Z(n24664) );
  XNOR U24429 ( .A(n24665), .B(n24666), .Z(n24662) );
  AND U24430 ( .A(n287), .B(n24667), .Z(n24666) );
  XOR U24431 ( .A(n24668), .B(n24669), .Z(n24660) );
  AND U24432 ( .A(n291), .B(n24659), .Z(n24669) );
  XNOR U24433 ( .A(n24670), .B(n24657), .Z(n24659) );
  XOR U24434 ( .A(n24671), .B(n24672), .Z(n24657) );
  AND U24435 ( .A(n314), .B(n24673), .Z(n24672) );
  IV U24436 ( .A(n24668), .Z(n24670) );
  XOR U24437 ( .A(n24674), .B(n24675), .Z(n24668) );
  AND U24438 ( .A(n298), .B(n24667), .Z(n24675) );
  XNOR U24439 ( .A(n24665), .B(n24674), .Z(n24667) );
  XNOR U24440 ( .A(n24676), .B(n24677), .Z(n24665) );
  AND U24441 ( .A(n302), .B(n24678), .Z(n24677) );
  XOR U24442 ( .A(p_input[300]), .B(n24676), .Z(n24678) );
  XNOR U24443 ( .A(n24679), .B(n24680), .Z(n24676) );
  AND U24444 ( .A(n306), .B(n24681), .Z(n24680) );
  XOR U24445 ( .A(n24682), .B(n24683), .Z(n24674) );
  AND U24446 ( .A(n310), .B(n24673), .Z(n24683) );
  XNOR U24447 ( .A(n24684), .B(n24671), .Z(n24673) );
  XOR U24448 ( .A(n24685), .B(n24686), .Z(n24671) );
  AND U24449 ( .A(n333), .B(n24687), .Z(n24686) );
  IV U24450 ( .A(n24682), .Z(n24684) );
  XOR U24451 ( .A(n24688), .B(n24689), .Z(n24682) );
  AND U24452 ( .A(n317), .B(n24681), .Z(n24689) );
  XNOR U24453 ( .A(n24679), .B(n24688), .Z(n24681) );
  XNOR U24454 ( .A(n24690), .B(n24691), .Z(n24679) );
  AND U24455 ( .A(n321), .B(n24692), .Z(n24691) );
  XOR U24456 ( .A(p_input[332]), .B(n24690), .Z(n24692) );
  XNOR U24457 ( .A(n24693), .B(n24694), .Z(n24690) );
  AND U24458 ( .A(n325), .B(n24695), .Z(n24694) );
  XOR U24459 ( .A(n24696), .B(n24697), .Z(n24688) );
  AND U24460 ( .A(n329), .B(n24687), .Z(n24697) );
  XNOR U24461 ( .A(n24698), .B(n24685), .Z(n24687) );
  XOR U24462 ( .A(n24699), .B(n24700), .Z(n24685) );
  AND U24463 ( .A(n352), .B(n24701), .Z(n24700) );
  IV U24464 ( .A(n24696), .Z(n24698) );
  XOR U24465 ( .A(n24702), .B(n24703), .Z(n24696) );
  AND U24466 ( .A(n336), .B(n24695), .Z(n24703) );
  XNOR U24467 ( .A(n24693), .B(n24702), .Z(n24695) );
  XNOR U24468 ( .A(n24704), .B(n24705), .Z(n24693) );
  AND U24469 ( .A(n340), .B(n24706), .Z(n24705) );
  XOR U24470 ( .A(p_input[364]), .B(n24704), .Z(n24706) );
  XNOR U24471 ( .A(n24707), .B(n24708), .Z(n24704) );
  AND U24472 ( .A(n344), .B(n24709), .Z(n24708) );
  XOR U24473 ( .A(n24710), .B(n24711), .Z(n24702) );
  AND U24474 ( .A(n348), .B(n24701), .Z(n24711) );
  XNOR U24475 ( .A(n24712), .B(n24699), .Z(n24701) );
  XOR U24476 ( .A(n24713), .B(n24714), .Z(n24699) );
  AND U24477 ( .A(n371), .B(n24715), .Z(n24714) );
  IV U24478 ( .A(n24710), .Z(n24712) );
  XOR U24479 ( .A(n24716), .B(n24717), .Z(n24710) );
  AND U24480 ( .A(n355), .B(n24709), .Z(n24717) );
  XNOR U24481 ( .A(n24707), .B(n24716), .Z(n24709) );
  XNOR U24482 ( .A(n24718), .B(n24719), .Z(n24707) );
  AND U24483 ( .A(n359), .B(n24720), .Z(n24719) );
  XOR U24484 ( .A(p_input[396]), .B(n24718), .Z(n24720) );
  XNOR U24485 ( .A(n24721), .B(n24722), .Z(n24718) );
  AND U24486 ( .A(n363), .B(n24723), .Z(n24722) );
  XOR U24487 ( .A(n24724), .B(n24725), .Z(n24716) );
  AND U24488 ( .A(n367), .B(n24715), .Z(n24725) );
  XNOR U24489 ( .A(n24726), .B(n24713), .Z(n24715) );
  XOR U24490 ( .A(n24727), .B(n24728), .Z(n24713) );
  AND U24491 ( .A(n390), .B(n24729), .Z(n24728) );
  IV U24492 ( .A(n24724), .Z(n24726) );
  XOR U24493 ( .A(n24730), .B(n24731), .Z(n24724) );
  AND U24494 ( .A(n374), .B(n24723), .Z(n24731) );
  XNOR U24495 ( .A(n24721), .B(n24730), .Z(n24723) );
  XNOR U24496 ( .A(n24732), .B(n24733), .Z(n24721) );
  AND U24497 ( .A(n378), .B(n24734), .Z(n24733) );
  XOR U24498 ( .A(p_input[428]), .B(n24732), .Z(n24734) );
  XNOR U24499 ( .A(n24735), .B(n24736), .Z(n24732) );
  AND U24500 ( .A(n382), .B(n24737), .Z(n24736) );
  XOR U24501 ( .A(n24738), .B(n24739), .Z(n24730) );
  AND U24502 ( .A(n386), .B(n24729), .Z(n24739) );
  XNOR U24503 ( .A(n24740), .B(n24727), .Z(n24729) );
  XOR U24504 ( .A(n24741), .B(n24742), .Z(n24727) );
  AND U24505 ( .A(n409), .B(n24743), .Z(n24742) );
  IV U24506 ( .A(n24738), .Z(n24740) );
  XOR U24507 ( .A(n24744), .B(n24745), .Z(n24738) );
  AND U24508 ( .A(n393), .B(n24737), .Z(n24745) );
  XNOR U24509 ( .A(n24735), .B(n24744), .Z(n24737) );
  XNOR U24510 ( .A(n24746), .B(n24747), .Z(n24735) );
  AND U24511 ( .A(n397), .B(n24748), .Z(n24747) );
  XOR U24512 ( .A(p_input[460]), .B(n24746), .Z(n24748) );
  XNOR U24513 ( .A(n24749), .B(n24750), .Z(n24746) );
  AND U24514 ( .A(n401), .B(n24751), .Z(n24750) );
  XOR U24515 ( .A(n24752), .B(n24753), .Z(n24744) );
  AND U24516 ( .A(n405), .B(n24743), .Z(n24753) );
  XNOR U24517 ( .A(n24754), .B(n24741), .Z(n24743) );
  XOR U24518 ( .A(n24755), .B(n24756), .Z(n24741) );
  AND U24519 ( .A(n428), .B(n24757), .Z(n24756) );
  IV U24520 ( .A(n24752), .Z(n24754) );
  XOR U24521 ( .A(n24758), .B(n24759), .Z(n24752) );
  AND U24522 ( .A(n412), .B(n24751), .Z(n24759) );
  XNOR U24523 ( .A(n24749), .B(n24758), .Z(n24751) );
  XNOR U24524 ( .A(n24760), .B(n24761), .Z(n24749) );
  AND U24525 ( .A(n416), .B(n24762), .Z(n24761) );
  XOR U24526 ( .A(p_input[492]), .B(n24760), .Z(n24762) );
  XNOR U24527 ( .A(n24763), .B(n24764), .Z(n24760) );
  AND U24528 ( .A(n420), .B(n24765), .Z(n24764) );
  XOR U24529 ( .A(n24766), .B(n24767), .Z(n24758) );
  AND U24530 ( .A(n424), .B(n24757), .Z(n24767) );
  XNOR U24531 ( .A(n24768), .B(n24755), .Z(n24757) );
  XOR U24532 ( .A(n24769), .B(n24770), .Z(n24755) );
  AND U24533 ( .A(n447), .B(n24771), .Z(n24770) );
  IV U24534 ( .A(n24766), .Z(n24768) );
  XOR U24535 ( .A(n24772), .B(n24773), .Z(n24766) );
  AND U24536 ( .A(n431), .B(n24765), .Z(n24773) );
  XNOR U24537 ( .A(n24763), .B(n24772), .Z(n24765) );
  XNOR U24538 ( .A(n24774), .B(n24775), .Z(n24763) );
  AND U24539 ( .A(n435), .B(n24776), .Z(n24775) );
  XOR U24540 ( .A(p_input[524]), .B(n24774), .Z(n24776) );
  XNOR U24541 ( .A(n24777), .B(n24778), .Z(n24774) );
  AND U24542 ( .A(n439), .B(n24779), .Z(n24778) );
  XOR U24543 ( .A(n24780), .B(n24781), .Z(n24772) );
  AND U24544 ( .A(n443), .B(n24771), .Z(n24781) );
  XNOR U24545 ( .A(n24782), .B(n24769), .Z(n24771) );
  XOR U24546 ( .A(n24783), .B(n24784), .Z(n24769) );
  AND U24547 ( .A(n466), .B(n24785), .Z(n24784) );
  IV U24548 ( .A(n24780), .Z(n24782) );
  XOR U24549 ( .A(n24786), .B(n24787), .Z(n24780) );
  AND U24550 ( .A(n450), .B(n24779), .Z(n24787) );
  XNOR U24551 ( .A(n24777), .B(n24786), .Z(n24779) );
  XNOR U24552 ( .A(n24788), .B(n24789), .Z(n24777) );
  AND U24553 ( .A(n454), .B(n24790), .Z(n24789) );
  XOR U24554 ( .A(p_input[556]), .B(n24788), .Z(n24790) );
  XNOR U24555 ( .A(n24791), .B(n24792), .Z(n24788) );
  AND U24556 ( .A(n458), .B(n24793), .Z(n24792) );
  XOR U24557 ( .A(n24794), .B(n24795), .Z(n24786) );
  AND U24558 ( .A(n462), .B(n24785), .Z(n24795) );
  XNOR U24559 ( .A(n24796), .B(n24783), .Z(n24785) );
  XOR U24560 ( .A(n24797), .B(n24798), .Z(n24783) );
  AND U24561 ( .A(n485), .B(n24799), .Z(n24798) );
  IV U24562 ( .A(n24794), .Z(n24796) );
  XOR U24563 ( .A(n24800), .B(n24801), .Z(n24794) );
  AND U24564 ( .A(n469), .B(n24793), .Z(n24801) );
  XNOR U24565 ( .A(n24791), .B(n24800), .Z(n24793) );
  XNOR U24566 ( .A(n24802), .B(n24803), .Z(n24791) );
  AND U24567 ( .A(n473), .B(n24804), .Z(n24803) );
  XOR U24568 ( .A(p_input[588]), .B(n24802), .Z(n24804) );
  XNOR U24569 ( .A(n24805), .B(n24806), .Z(n24802) );
  AND U24570 ( .A(n477), .B(n24807), .Z(n24806) );
  XOR U24571 ( .A(n24808), .B(n24809), .Z(n24800) );
  AND U24572 ( .A(n481), .B(n24799), .Z(n24809) );
  XNOR U24573 ( .A(n24810), .B(n24797), .Z(n24799) );
  XOR U24574 ( .A(n24811), .B(n24812), .Z(n24797) );
  AND U24575 ( .A(n504), .B(n24813), .Z(n24812) );
  IV U24576 ( .A(n24808), .Z(n24810) );
  XOR U24577 ( .A(n24814), .B(n24815), .Z(n24808) );
  AND U24578 ( .A(n488), .B(n24807), .Z(n24815) );
  XNOR U24579 ( .A(n24805), .B(n24814), .Z(n24807) );
  XNOR U24580 ( .A(n24816), .B(n24817), .Z(n24805) );
  AND U24581 ( .A(n492), .B(n24818), .Z(n24817) );
  XOR U24582 ( .A(p_input[620]), .B(n24816), .Z(n24818) );
  XNOR U24583 ( .A(n24819), .B(n24820), .Z(n24816) );
  AND U24584 ( .A(n496), .B(n24821), .Z(n24820) );
  XOR U24585 ( .A(n24822), .B(n24823), .Z(n24814) );
  AND U24586 ( .A(n500), .B(n24813), .Z(n24823) );
  XNOR U24587 ( .A(n24824), .B(n24811), .Z(n24813) );
  XOR U24588 ( .A(n24825), .B(n24826), .Z(n24811) );
  AND U24589 ( .A(n523), .B(n24827), .Z(n24826) );
  IV U24590 ( .A(n24822), .Z(n24824) );
  XOR U24591 ( .A(n24828), .B(n24829), .Z(n24822) );
  AND U24592 ( .A(n507), .B(n24821), .Z(n24829) );
  XNOR U24593 ( .A(n24819), .B(n24828), .Z(n24821) );
  XNOR U24594 ( .A(n24830), .B(n24831), .Z(n24819) );
  AND U24595 ( .A(n511), .B(n24832), .Z(n24831) );
  XOR U24596 ( .A(p_input[652]), .B(n24830), .Z(n24832) );
  XNOR U24597 ( .A(n24833), .B(n24834), .Z(n24830) );
  AND U24598 ( .A(n515), .B(n24835), .Z(n24834) );
  XOR U24599 ( .A(n24836), .B(n24837), .Z(n24828) );
  AND U24600 ( .A(n519), .B(n24827), .Z(n24837) );
  XNOR U24601 ( .A(n24838), .B(n24825), .Z(n24827) );
  XOR U24602 ( .A(n24839), .B(n24840), .Z(n24825) );
  AND U24603 ( .A(n542), .B(n24841), .Z(n24840) );
  IV U24604 ( .A(n24836), .Z(n24838) );
  XOR U24605 ( .A(n24842), .B(n24843), .Z(n24836) );
  AND U24606 ( .A(n526), .B(n24835), .Z(n24843) );
  XNOR U24607 ( .A(n24833), .B(n24842), .Z(n24835) );
  XNOR U24608 ( .A(n24844), .B(n24845), .Z(n24833) );
  AND U24609 ( .A(n530), .B(n24846), .Z(n24845) );
  XOR U24610 ( .A(p_input[684]), .B(n24844), .Z(n24846) );
  XNOR U24611 ( .A(n24847), .B(n24848), .Z(n24844) );
  AND U24612 ( .A(n534), .B(n24849), .Z(n24848) );
  XOR U24613 ( .A(n24850), .B(n24851), .Z(n24842) );
  AND U24614 ( .A(n538), .B(n24841), .Z(n24851) );
  XNOR U24615 ( .A(n24852), .B(n24839), .Z(n24841) );
  XOR U24616 ( .A(n24853), .B(n24854), .Z(n24839) );
  AND U24617 ( .A(n561), .B(n24855), .Z(n24854) );
  IV U24618 ( .A(n24850), .Z(n24852) );
  XOR U24619 ( .A(n24856), .B(n24857), .Z(n24850) );
  AND U24620 ( .A(n545), .B(n24849), .Z(n24857) );
  XNOR U24621 ( .A(n24847), .B(n24856), .Z(n24849) );
  XNOR U24622 ( .A(n24858), .B(n24859), .Z(n24847) );
  AND U24623 ( .A(n549), .B(n24860), .Z(n24859) );
  XOR U24624 ( .A(p_input[716]), .B(n24858), .Z(n24860) );
  XNOR U24625 ( .A(n24861), .B(n24862), .Z(n24858) );
  AND U24626 ( .A(n553), .B(n24863), .Z(n24862) );
  XOR U24627 ( .A(n24864), .B(n24865), .Z(n24856) );
  AND U24628 ( .A(n557), .B(n24855), .Z(n24865) );
  XNOR U24629 ( .A(n24866), .B(n24853), .Z(n24855) );
  XOR U24630 ( .A(n24867), .B(n24868), .Z(n24853) );
  AND U24631 ( .A(n580), .B(n24869), .Z(n24868) );
  IV U24632 ( .A(n24864), .Z(n24866) );
  XOR U24633 ( .A(n24870), .B(n24871), .Z(n24864) );
  AND U24634 ( .A(n564), .B(n24863), .Z(n24871) );
  XNOR U24635 ( .A(n24861), .B(n24870), .Z(n24863) );
  XNOR U24636 ( .A(n24872), .B(n24873), .Z(n24861) );
  AND U24637 ( .A(n568), .B(n24874), .Z(n24873) );
  XOR U24638 ( .A(p_input[748]), .B(n24872), .Z(n24874) );
  XNOR U24639 ( .A(n24875), .B(n24876), .Z(n24872) );
  AND U24640 ( .A(n572), .B(n24877), .Z(n24876) );
  XOR U24641 ( .A(n24878), .B(n24879), .Z(n24870) );
  AND U24642 ( .A(n576), .B(n24869), .Z(n24879) );
  XNOR U24643 ( .A(n24880), .B(n24867), .Z(n24869) );
  XOR U24644 ( .A(n24881), .B(n24882), .Z(n24867) );
  AND U24645 ( .A(n599), .B(n24883), .Z(n24882) );
  IV U24646 ( .A(n24878), .Z(n24880) );
  XOR U24647 ( .A(n24884), .B(n24885), .Z(n24878) );
  AND U24648 ( .A(n583), .B(n24877), .Z(n24885) );
  XNOR U24649 ( .A(n24875), .B(n24884), .Z(n24877) );
  XNOR U24650 ( .A(n24886), .B(n24887), .Z(n24875) );
  AND U24651 ( .A(n587), .B(n24888), .Z(n24887) );
  XOR U24652 ( .A(p_input[780]), .B(n24886), .Z(n24888) );
  XNOR U24653 ( .A(n24889), .B(n24890), .Z(n24886) );
  AND U24654 ( .A(n591), .B(n24891), .Z(n24890) );
  XOR U24655 ( .A(n24892), .B(n24893), .Z(n24884) );
  AND U24656 ( .A(n595), .B(n24883), .Z(n24893) );
  XNOR U24657 ( .A(n24894), .B(n24881), .Z(n24883) );
  XOR U24658 ( .A(n24895), .B(n24896), .Z(n24881) );
  AND U24659 ( .A(n618), .B(n24897), .Z(n24896) );
  IV U24660 ( .A(n24892), .Z(n24894) );
  XOR U24661 ( .A(n24898), .B(n24899), .Z(n24892) );
  AND U24662 ( .A(n602), .B(n24891), .Z(n24899) );
  XNOR U24663 ( .A(n24889), .B(n24898), .Z(n24891) );
  XNOR U24664 ( .A(n24900), .B(n24901), .Z(n24889) );
  AND U24665 ( .A(n606), .B(n24902), .Z(n24901) );
  XOR U24666 ( .A(p_input[812]), .B(n24900), .Z(n24902) );
  XNOR U24667 ( .A(n24903), .B(n24904), .Z(n24900) );
  AND U24668 ( .A(n610), .B(n24905), .Z(n24904) );
  XOR U24669 ( .A(n24906), .B(n24907), .Z(n24898) );
  AND U24670 ( .A(n614), .B(n24897), .Z(n24907) );
  XNOR U24671 ( .A(n24908), .B(n24895), .Z(n24897) );
  XOR U24672 ( .A(n24909), .B(n24910), .Z(n24895) );
  AND U24673 ( .A(n637), .B(n24911), .Z(n24910) );
  IV U24674 ( .A(n24906), .Z(n24908) );
  XOR U24675 ( .A(n24912), .B(n24913), .Z(n24906) );
  AND U24676 ( .A(n621), .B(n24905), .Z(n24913) );
  XNOR U24677 ( .A(n24903), .B(n24912), .Z(n24905) );
  XNOR U24678 ( .A(n24914), .B(n24915), .Z(n24903) );
  AND U24679 ( .A(n625), .B(n24916), .Z(n24915) );
  XOR U24680 ( .A(p_input[844]), .B(n24914), .Z(n24916) );
  XNOR U24681 ( .A(n24917), .B(n24918), .Z(n24914) );
  AND U24682 ( .A(n629), .B(n24919), .Z(n24918) );
  XOR U24683 ( .A(n24920), .B(n24921), .Z(n24912) );
  AND U24684 ( .A(n633), .B(n24911), .Z(n24921) );
  XNOR U24685 ( .A(n24922), .B(n24909), .Z(n24911) );
  XOR U24686 ( .A(n24923), .B(n24924), .Z(n24909) );
  AND U24687 ( .A(n656), .B(n24925), .Z(n24924) );
  IV U24688 ( .A(n24920), .Z(n24922) );
  XOR U24689 ( .A(n24926), .B(n24927), .Z(n24920) );
  AND U24690 ( .A(n640), .B(n24919), .Z(n24927) );
  XNOR U24691 ( .A(n24917), .B(n24926), .Z(n24919) );
  XNOR U24692 ( .A(n24928), .B(n24929), .Z(n24917) );
  AND U24693 ( .A(n644), .B(n24930), .Z(n24929) );
  XOR U24694 ( .A(p_input[876]), .B(n24928), .Z(n24930) );
  XNOR U24695 ( .A(n24931), .B(n24932), .Z(n24928) );
  AND U24696 ( .A(n648), .B(n24933), .Z(n24932) );
  XOR U24697 ( .A(n24934), .B(n24935), .Z(n24926) );
  AND U24698 ( .A(n652), .B(n24925), .Z(n24935) );
  XNOR U24699 ( .A(n24936), .B(n24923), .Z(n24925) );
  XOR U24700 ( .A(n24937), .B(n24938), .Z(n24923) );
  AND U24701 ( .A(n675), .B(n24939), .Z(n24938) );
  IV U24702 ( .A(n24934), .Z(n24936) );
  XOR U24703 ( .A(n24940), .B(n24941), .Z(n24934) );
  AND U24704 ( .A(n659), .B(n24933), .Z(n24941) );
  XNOR U24705 ( .A(n24931), .B(n24940), .Z(n24933) );
  XNOR U24706 ( .A(n24942), .B(n24943), .Z(n24931) );
  AND U24707 ( .A(n663), .B(n24944), .Z(n24943) );
  XOR U24708 ( .A(p_input[908]), .B(n24942), .Z(n24944) );
  XNOR U24709 ( .A(n24945), .B(n24946), .Z(n24942) );
  AND U24710 ( .A(n667), .B(n24947), .Z(n24946) );
  XOR U24711 ( .A(n24948), .B(n24949), .Z(n24940) );
  AND U24712 ( .A(n671), .B(n24939), .Z(n24949) );
  XNOR U24713 ( .A(n24950), .B(n24937), .Z(n24939) );
  XOR U24714 ( .A(n24951), .B(n24952), .Z(n24937) );
  AND U24715 ( .A(n694), .B(n24953), .Z(n24952) );
  IV U24716 ( .A(n24948), .Z(n24950) );
  XOR U24717 ( .A(n24954), .B(n24955), .Z(n24948) );
  AND U24718 ( .A(n678), .B(n24947), .Z(n24955) );
  XNOR U24719 ( .A(n24945), .B(n24954), .Z(n24947) );
  XNOR U24720 ( .A(n24956), .B(n24957), .Z(n24945) );
  AND U24721 ( .A(n682), .B(n24958), .Z(n24957) );
  XOR U24722 ( .A(p_input[940]), .B(n24956), .Z(n24958) );
  XNOR U24723 ( .A(n24959), .B(n24960), .Z(n24956) );
  AND U24724 ( .A(n686), .B(n24961), .Z(n24960) );
  XOR U24725 ( .A(n24962), .B(n24963), .Z(n24954) );
  AND U24726 ( .A(n690), .B(n24953), .Z(n24963) );
  XNOR U24727 ( .A(n24964), .B(n24951), .Z(n24953) );
  XOR U24728 ( .A(n24965), .B(n24966), .Z(n24951) );
  AND U24729 ( .A(n713), .B(n24967), .Z(n24966) );
  IV U24730 ( .A(n24962), .Z(n24964) );
  XOR U24731 ( .A(n24968), .B(n24969), .Z(n24962) );
  AND U24732 ( .A(n697), .B(n24961), .Z(n24969) );
  XNOR U24733 ( .A(n24959), .B(n24968), .Z(n24961) );
  XNOR U24734 ( .A(n24970), .B(n24971), .Z(n24959) );
  AND U24735 ( .A(n701), .B(n24972), .Z(n24971) );
  XOR U24736 ( .A(p_input[972]), .B(n24970), .Z(n24972) );
  XNOR U24737 ( .A(n24973), .B(n24974), .Z(n24970) );
  AND U24738 ( .A(n705), .B(n24975), .Z(n24974) );
  XOR U24739 ( .A(n24976), .B(n24977), .Z(n24968) );
  AND U24740 ( .A(n709), .B(n24967), .Z(n24977) );
  XNOR U24741 ( .A(n24978), .B(n24965), .Z(n24967) );
  XOR U24742 ( .A(n24979), .B(n24980), .Z(n24965) );
  AND U24743 ( .A(n732), .B(n24981), .Z(n24980) );
  IV U24744 ( .A(n24976), .Z(n24978) );
  XOR U24745 ( .A(n24982), .B(n24983), .Z(n24976) );
  AND U24746 ( .A(n716), .B(n24975), .Z(n24983) );
  XNOR U24747 ( .A(n24973), .B(n24982), .Z(n24975) );
  XNOR U24748 ( .A(n24984), .B(n24985), .Z(n24973) );
  AND U24749 ( .A(n720), .B(n24986), .Z(n24985) );
  XOR U24750 ( .A(p_input[1004]), .B(n24984), .Z(n24986) );
  XNOR U24751 ( .A(n24987), .B(n24988), .Z(n24984) );
  AND U24752 ( .A(n724), .B(n24989), .Z(n24988) );
  XOR U24753 ( .A(n24990), .B(n24991), .Z(n24982) );
  AND U24754 ( .A(n728), .B(n24981), .Z(n24991) );
  XNOR U24755 ( .A(n24992), .B(n24979), .Z(n24981) );
  XOR U24756 ( .A(n24993), .B(n24994), .Z(n24979) );
  AND U24757 ( .A(n751), .B(n24995), .Z(n24994) );
  IV U24758 ( .A(n24990), .Z(n24992) );
  XOR U24759 ( .A(n24996), .B(n24997), .Z(n24990) );
  AND U24760 ( .A(n735), .B(n24989), .Z(n24997) );
  XNOR U24761 ( .A(n24987), .B(n24996), .Z(n24989) );
  XNOR U24762 ( .A(n24998), .B(n24999), .Z(n24987) );
  AND U24763 ( .A(n739), .B(n25000), .Z(n24999) );
  XOR U24764 ( .A(p_input[1036]), .B(n24998), .Z(n25000) );
  XNOR U24765 ( .A(n25001), .B(n25002), .Z(n24998) );
  AND U24766 ( .A(n743), .B(n25003), .Z(n25002) );
  XOR U24767 ( .A(n25004), .B(n25005), .Z(n24996) );
  AND U24768 ( .A(n747), .B(n24995), .Z(n25005) );
  XNOR U24769 ( .A(n25006), .B(n24993), .Z(n24995) );
  XOR U24770 ( .A(n25007), .B(n25008), .Z(n24993) );
  AND U24771 ( .A(n770), .B(n25009), .Z(n25008) );
  IV U24772 ( .A(n25004), .Z(n25006) );
  XOR U24773 ( .A(n25010), .B(n25011), .Z(n25004) );
  AND U24774 ( .A(n754), .B(n25003), .Z(n25011) );
  XNOR U24775 ( .A(n25001), .B(n25010), .Z(n25003) );
  XNOR U24776 ( .A(n25012), .B(n25013), .Z(n25001) );
  AND U24777 ( .A(n758), .B(n25014), .Z(n25013) );
  XOR U24778 ( .A(p_input[1068]), .B(n25012), .Z(n25014) );
  XNOR U24779 ( .A(n25015), .B(n25016), .Z(n25012) );
  AND U24780 ( .A(n762), .B(n25017), .Z(n25016) );
  XOR U24781 ( .A(n25018), .B(n25019), .Z(n25010) );
  AND U24782 ( .A(n766), .B(n25009), .Z(n25019) );
  XNOR U24783 ( .A(n25020), .B(n25007), .Z(n25009) );
  XOR U24784 ( .A(n25021), .B(n25022), .Z(n25007) );
  AND U24785 ( .A(n789), .B(n25023), .Z(n25022) );
  IV U24786 ( .A(n25018), .Z(n25020) );
  XOR U24787 ( .A(n25024), .B(n25025), .Z(n25018) );
  AND U24788 ( .A(n773), .B(n25017), .Z(n25025) );
  XNOR U24789 ( .A(n25015), .B(n25024), .Z(n25017) );
  XNOR U24790 ( .A(n25026), .B(n25027), .Z(n25015) );
  AND U24791 ( .A(n777), .B(n25028), .Z(n25027) );
  XOR U24792 ( .A(p_input[1100]), .B(n25026), .Z(n25028) );
  XNOR U24793 ( .A(n25029), .B(n25030), .Z(n25026) );
  AND U24794 ( .A(n781), .B(n25031), .Z(n25030) );
  XOR U24795 ( .A(n25032), .B(n25033), .Z(n25024) );
  AND U24796 ( .A(n785), .B(n25023), .Z(n25033) );
  XNOR U24797 ( .A(n25034), .B(n25021), .Z(n25023) );
  XOR U24798 ( .A(n25035), .B(n25036), .Z(n25021) );
  AND U24799 ( .A(n808), .B(n25037), .Z(n25036) );
  IV U24800 ( .A(n25032), .Z(n25034) );
  XOR U24801 ( .A(n25038), .B(n25039), .Z(n25032) );
  AND U24802 ( .A(n792), .B(n25031), .Z(n25039) );
  XNOR U24803 ( .A(n25029), .B(n25038), .Z(n25031) );
  XNOR U24804 ( .A(n25040), .B(n25041), .Z(n25029) );
  AND U24805 ( .A(n796), .B(n25042), .Z(n25041) );
  XOR U24806 ( .A(p_input[1132]), .B(n25040), .Z(n25042) );
  XNOR U24807 ( .A(n25043), .B(n25044), .Z(n25040) );
  AND U24808 ( .A(n800), .B(n25045), .Z(n25044) );
  XOR U24809 ( .A(n25046), .B(n25047), .Z(n25038) );
  AND U24810 ( .A(n804), .B(n25037), .Z(n25047) );
  XNOR U24811 ( .A(n25048), .B(n25035), .Z(n25037) );
  XOR U24812 ( .A(n25049), .B(n25050), .Z(n25035) );
  AND U24813 ( .A(n827), .B(n25051), .Z(n25050) );
  IV U24814 ( .A(n25046), .Z(n25048) );
  XOR U24815 ( .A(n25052), .B(n25053), .Z(n25046) );
  AND U24816 ( .A(n811), .B(n25045), .Z(n25053) );
  XNOR U24817 ( .A(n25043), .B(n25052), .Z(n25045) );
  XNOR U24818 ( .A(n25054), .B(n25055), .Z(n25043) );
  AND U24819 ( .A(n815), .B(n25056), .Z(n25055) );
  XOR U24820 ( .A(p_input[1164]), .B(n25054), .Z(n25056) );
  XNOR U24821 ( .A(n25057), .B(n25058), .Z(n25054) );
  AND U24822 ( .A(n819), .B(n25059), .Z(n25058) );
  XOR U24823 ( .A(n25060), .B(n25061), .Z(n25052) );
  AND U24824 ( .A(n823), .B(n25051), .Z(n25061) );
  XNOR U24825 ( .A(n25062), .B(n25049), .Z(n25051) );
  XOR U24826 ( .A(n25063), .B(n25064), .Z(n25049) );
  AND U24827 ( .A(n846), .B(n25065), .Z(n25064) );
  IV U24828 ( .A(n25060), .Z(n25062) );
  XOR U24829 ( .A(n25066), .B(n25067), .Z(n25060) );
  AND U24830 ( .A(n830), .B(n25059), .Z(n25067) );
  XNOR U24831 ( .A(n25057), .B(n25066), .Z(n25059) );
  XNOR U24832 ( .A(n25068), .B(n25069), .Z(n25057) );
  AND U24833 ( .A(n834), .B(n25070), .Z(n25069) );
  XOR U24834 ( .A(p_input[1196]), .B(n25068), .Z(n25070) );
  XNOR U24835 ( .A(n25071), .B(n25072), .Z(n25068) );
  AND U24836 ( .A(n838), .B(n25073), .Z(n25072) );
  XOR U24837 ( .A(n25074), .B(n25075), .Z(n25066) );
  AND U24838 ( .A(n842), .B(n25065), .Z(n25075) );
  XNOR U24839 ( .A(n25076), .B(n25063), .Z(n25065) );
  XOR U24840 ( .A(n25077), .B(n25078), .Z(n25063) );
  AND U24841 ( .A(n865), .B(n25079), .Z(n25078) );
  IV U24842 ( .A(n25074), .Z(n25076) );
  XOR U24843 ( .A(n25080), .B(n25081), .Z(n25074) );
  AND U24844 ( .A(n849), .B(n25073), .Z(n25081) );
  XNOR U24845 ( .A(n25071), .B(n25080), .Z(n25073) );
  XNOR U24846 ( .A(n25082), .B(n25083), .Z(n25071) );
  AND U24847 ( .A(n853), .B(n25084), .Z(n25083) );
  XOR U24848 ( .A(p_input[1228]), .B(n25082), .Z(n25084) );
  XNOR U24849 ( .A(n25085), .B(n25086), .Z(n25082) );
  AND U24850 ( .A(n857), .B(n25087), .Z(n25086) );
  XOR U24851 ( .A(n25088), .B(n25089), .Z(n25080) );
  AND U24852 ( .A(n861), .B(n25079), .Z(n25089) );
  XNOR U24853 ( .A(n25090), .B(n25077), .Z(n25079) );
  XOR U24854 ( .A(n25091), .B(n25092), .Z(n25077) );
  AND U24855 ( .A(n884), .B(n25093), .Z(n25092) );
  IV U24856 ( .A(n25088), .Z(n25090) );
  XOR U24857 ( .A(n25094), .B(n25095), .Z(n25088) );
  AND U24858 ( .A(n868), .B(n25087), .Z(n25095) );
  XNOR U24859 ( .A(n25085), .B(n25094), .Z(n25087) );
  XNOR U24860 ( .A(n25096), .B(n25097), .Z(n25085) );
  AND U24861 ( .A(n872), .B(n25098), .Z(n25097) );
  XOR U24862 ( .A(p_input[1260]), .B(n25096), .Z(n25098) );
  XNOR U24863 ( .A(n25099), .B(n25100), .Z(n25096) );
  AND U24864 ( .A(n876), .B(n25101), .Z(n25100) );
  XOR U24865 ( .A(n25102), .B(n25103), .Z(n25094) );
  AND U24866 ( .A(n880), .B(n25093), .Z(n25103) );
  XNOR U24867 ( .A(n25104), .B(n25091), .Z(n25093) );
  XOR U24868 ( .A(n25105), .B(n25106), .Z(n25091) );
  AND U24869 ( .A(n903), .B(n25107), .Z(n25106) );
  IV U24870 ( .A(n25102), .Z(n25104) );
  XOR U24871 ( .A(n25108), .B(n25109), .Z(n25102) );
  AND U24872 ( .A(n887), .B(n25101), .Z(n25109) );
  XNOR U24873 ( .A(n25099), .B(n25108), .Z(n25101) );
  XNOR U24874 ( .A(n25110), .B(n25111), .Z(n25099) );
  AND U24875 ( .A(n891), .B(n25112), .Z(n25111) );
  XOR U24876 ( .A(p_input[1292]), .B(n25110), .Z(n25112) );
  XNOR U24877 ( .A(n25113), .B(n25114), .Z(n25110) );
  AND U24878 ( .A(n895), .B(n25115), .Z(n25114) );
  XOR U24879 ( .A(n25116), .B(n25117), .Z(n25108) );
  AND U24880 ( .A(n899), .B(n25107), .Z(n25117) );
  XNOR U24881 ( .A(n25118), .B(n25105), .Z(n25107) );
  XOR U24882 ( .A(n25119), .B(n25120), .Z(n25105) );
  AND U24883 ( .A(n922), .B(n25121), .Z(n25120) );
  IV U24884 ( .A(n25116), .Z(n25118) );
  XOR U24885 ( .A(n25122), .B(n25123), .Z(n25116) );
  AND U24886 ( .A(n906), .B(n25115), .Z(n25123) );
  XNOR U24887 ( .A(n25113), .B(n25122), .Z(n25115) );
  XNOR U24888 ( .A(n25124), .B(n25125), .Z(n25113) );
  AND U24889 ( .A(n910), .B(n25126), .Z(n25125) );
  XOR U24890 ( .A(p_input[1324]), .B(n25124), .Z(n25126) );
  XNOR U24891 ( .A(n25127), .B(n25128), .Z(n25124) );
  AND U24892 ( .A(n914), .B(n25129), .Z(n25128) );
  XOR U24893 ( .A(n25130), .B(n25131), .Z(n25122) );
  AND U24894 ( .A(n918), .B(n25121), .Z(n25131) );
  XNOR U24895 ( .A(n25132), .B(n25119), .Z(n25121) );
  XOR U24896 ( .A(n25133), .B(n25134), .Z(n25119) );
  AND U24897 ( .A(n941), .B(n25135), .Z(n25134) );
  IV U24898 ( .A(n25130), .Z(n25132) );
  XOR U24899 ( .A(n25136), .B(n25137), .Z(n25130) );
  AND U24900 ( .A(n925), .B(n25129), .Z(n25137) );
  XNOR U24901 ( .A(n25127), .B(n25136), .Z(n25129) );
  XNOR U24902 ( .A(n25138), .B(n25139), .Z(n25127) );
  AND U24903 ( .A(n929), .B(n25140), .Z(n25139) );
  XOR U24904 ( .A(p_input[1356]), .B(n25138), .Z(n25140) );
  XNOR U24905 ( .A(n25141), .B(n25142), .Z(n25138) );
  AND U24906 ( .A(n933), .B(n25143), .Z(n25142) );
  XOR U24907 ( .A(n25144), .B(n25145), .Z(n25136) );
  AND U24908 ( .A(n937), .B(n25135), .Z(n25145) );
  XNOR U24909 ( .A(n25146), .B(n25133), .Z(n25135) );
  XOR U24910 ( .A(n25147), .B(n25148), .Z(n25133) );
  AND U24911 ( .A(n960), .B(n25149), .Z(n25148) );
  IV U24912 ( .A(n25144), .Z(n25146) );
  XOR U24913 ( .A(n25150), .B(n25151), .Z(n25144) );
  AND U24914 ( .A(n944), .B(n25143), .Z(n25151) );
  XNOR U24915 ( .A(n25141), .B(n25150), .Z(n25143) );
  XNOR U24916 ( .A(n25152), .B(n25153), .Z(n25141) );
  AND U24917 ( .A(n948), .B(n25154), .Z(n25153) );
  XOR U24918 ( .A(p_input[1388]), .B(n25152), .Z(n25154) );
  XNOR U24919 ( .A(n25155), .B(n25156), .Z(n25152) );
  AND U24920 ( .A(n952), .B(n25157), .Z(n25156) );
  XOR U24921 ( .A(n25158), .B(n25159), .Z(n25150) );
  AND U24922 ( .A(n956), .B(n25149), .Z(n25159) );
  XNOR U24923 ( .A(n25160), .B(n25147), .Z(n25149) );
  XOR U24924 ( .A(n25161), .B(n25162), .Z(n25147) );
  AND U24925 ( .A(n979), .B(n25163), .Z(n25162) );
  IV U24926 ( .A(n25158), .Z(n25160) );
  XOR U24927 ( .A(n25164), .B(n25165), .Z(n25158) );
  AND U24928 ( .A(n963), .B(n25157), .Z(n25165) );
  XNOR U24929 ( .A(n25155), .B(n25164), .Z(n25157) );
  XNOR U24930 ( .A(n25166), .B(n25167), .Z(n25155) );
  AND U24931 ( .A(n967), .B(n25168), .Z(n25167) );
  XOR U24932 ( .A(p_input[1420]), .B(n25166), .Z(n25168) );
  XNOR U24933 ( .A(n25169), .B(n25170), .Z(n25166) );
  AND U24934 ( .A(n971), .B(n25171), .Z(n25170) );
  XOR U24935 ( .A(n25172), .B(n25173), .Z(n25164) );
  AND U24936 ( .A(n975), .B(n25163), .Z(n25173) );
  XNOR U24937 ( .A(n25174), .B(n25161), .Z(n25163) );
  XOR U24938 ( .A(n25175), .B(n25176), .Z(n25161) );
  AND U24939 ( .A(n998), .B(n25177), .Z(n25176) );
  IV U24940 ( .A(n25172), .Z(n25174) );
  XOR U24941 ( .A(n25178), .B(n25179), .Z(n25172) );
  AND U24942 ( .A(n982), .B(n25171), .Z(n25179) );
  XNOR U24943 ( .A(n25169), .B(n25178), .Z(n25171) );
  XNOR U24944 ( .A(n25180), .B(n25181), .Z(n25169) );
  AND U24945 ( .A(n986), .B(n25182), .Z(n25181) );
  XOR U24946 ( .A(p_input[1452]), .B(n25180), .Z(n25182) );
  XNOR U24947 ( .A(n25183), .B(n25184), .Z(n25180) );
  AND U24948 ( .A(n990), .B(n25185), .Z(n25184) );
  XOR U24949 ( .A(n25186), .B(n25187), .Z(n25178) );
  AND U24950 ( .A(n994), .B(n25177), .Z(n25187) );
  XNOR U24951 ( .A(n25188), .B(n25175), .Z(n25177) );
  XOR U24952 ( .A(n25189), .B(n25190), .Z(n25175) );
  AND U24953 ( .A(n1017), .B(n25191), .Z(n25190) );
  IV U24954 ( .A(n25186), .Z(n25188) );
  XOR U24955 ( .A(n25192), .B(n25193), .Z(n25186) );
  AND U24956 ( .A(n1001), .B(n25185), .Z(n25193) );
  XNOR U24957 ( .A(n25183), .B(n25192), .Z(n25185) );
  XNOR U24958 ( .A(n25194), .B(n25195), .Z(n25183) );
  AND U24959 ( .A(n1005), .B(n25196), .Z(n25195) );
  XOR U24960 ( .A(p_input[1484]), .B(n25194), .Z(n25196) );
  XNOR U24961 ( .A(n25197), .B(n25198), .Z(n25194) );
  AND U24962 ( .A(n1009), .B(n25199), .Z(n25198) );
  XOR U24963 ( .A(n25200), .B(n25201), .Z(n25192) );
  AND U24964 ( .A(n1013), .B(n25191), .Z(n25201) );
  XNOR U24965 ( .A(n25202), .B(n25189), .Z(n25191) );
  XOR U24966 ( .A(n25203), .B(n25204), .Z(n25189) );
  AND U24967 ( .A(n1036), .B(n25205), .Z(n25204) );
  IV U24968 ( .A(n25200), .Z(n25202) );
  XOR U24969 ( .A(n25206), .B(n25207), .Z(n25200) );
  AND U24970 ( .A(n1020), .B(n25199), .Z(n25207) );
  XNOR U24971 ( .A(n25197), .B(n25206), .Z(n25199) );
  XNOR U24972 ( .A(n25208), .B(n25209), .Z(n25197) );
  AND U24973 ( .A(n1024), .B(n25210), .Z(n25209) );
  XOR U24974 ( .A(p_input[1516]), .B(n25208), .Z(n25210) );
  XNOR U24975 ( .A(n25211), .B(n25212), .Z(n25208) );
  AND U24976 ( .A(n1028), .B(n25213), .Z(n25212) );
  XOR U24977 ( .A(n25214), .B(n25215), .Z(n25206) );
  AND U24978 ( .A(n1032), .B(n25205), .Z(n25215) );
  XNOR U24979 ( .A(n25216), .B(n25203), .Z(n25205) );
  XOR U24980 ( .A(n25217), .B(n25218), .Z(n25203) );
  AND U24981 ( .A(n1055), .B(n25219), .Z(n25218) );
  IV U24982 ( .A(n25214), .Z(n25216) );
  XOR U24983 ( .A(n25220), .B(n25221), .Z(n25214) );
  AND U24984 ( .A(n1039), .B(n25213), .Z(n25221) );
  XNOR U24985 ( .A(n25211), .B(n25220), .Z(n25213) );
  XNOR U24986 ( .A(n25222), .B(n25223), .Z(n25211) );
  AND U24987 ( .A(n1043), .B(n25224), .Z(n25223) );
  XOR U24988 ( .A(p_input[1548]), .B(n25222), .Z(n25224) );
  XNOR U24989 ( .A(n25225), .B(n25226), .Z(n25222) );
  AND U24990 ( .A(n1047), .B(n25227), .Z(n25226) );
  XOR U24991 ( .A(n25228), .B(n25229), .Z(n25220) );
  AND U24992 ( .A(n1051), .B(n25219), .Z(n25229) );
  XNOR U24993 ( .A(n25230), .B(n25217), .Z(n25219) );
  XOR U24994 ( .A(n25231), .B(n25232), .Z(n25217) );
  AND U24995 ( .A(n1074), .B(n25233), .Z(n25232) );
  IV U24996 ( .A(n25228), .Z(n25230) );
  XOR U24997 ( .A(n25234), .B(n25235), .Z(n25228) );
  AND U24998 ( .A(n1058), .B(n25227), .Z(n25235) );
  XNOR U24999 ( .A(n25225), .B(n25234), .Z(n25227) );
  XNOR U25000 ( .A(n25236), .B(n25237), .Z(n25225) );
  AND U25001 ( .A(n1062), .B(n25238), .Z(n25237) );
  XOR U25002 ( .A(p_input[1580]), .B(n25236), .Z(n25238) );
  XNOR U25003 ( .A(n25239), .B(n25240), .Z(n25236) );
  AND U25004 ( .A(n1066), .B(n25241), .Z(n25240) );
  XOR U25005 ( .A(n25242), .B(n25243), .Z(n25234) );
  AND U25006 ( .A(n1070), .B(n25233), .Z(n25243) );
  XNOR U25007 ( .A(n25244), .B(n25231), .Z(n25233) );
  XOR U25008 ( .A(n25245), .B(n25246), .Z(n25231) );
  AND U25009 ( .A(n1093), .B(n25247), .Z(n25246) );
  IV U25010 ( .A(n25242), .Z(n25244) );
  XOR U25011 ( .A(n25248), .B(n25249), .Z(n25242) );
  AND U25012 ( .A(n1077), .B(n25241), .Z(n25249) );
  XNOR U25013 ( .A(n25239), .B(n25248), .Z(n25241) );
  XNOR U25014 ( .A(n25250), .B(n25251), .Z(n25239) );
  AND U25015 ( .A(n1081), .B(n25252), .Z(n25251) );
  XOR U25016 ( .A(p_input[1612]), .B(n25250), .Z(n25252) );
  XNOR U25017 ( .A(n25253), .B(n25254), .Z(n25250) );
  AND U25018 ( .A(n1085), .B(n25255), .Z(n25254) );
  XOR U25019 ( .A(n25256), .B(n25257), .Z(n25248) );
  AND U25020 ( .A(n1089), .B(n25247), .Z(n25257) );
  XNOR U25021 ( .A(n25258), .B(n25245), .Z(n25247) );
  XOR U25022 ( .A(n25259), .B(n25260), .Z(n25245) );
  AND U25023 ( .A(n1112), .B(n25261), .Z(n25260) );
  IV U25024 ( .A(n25256), .Z(n25258) );
  XOR U25025 ( .A(n25262), .B(n25263), .Z(n25256) );
  AND U25026 ( .A(n1096), .B(n25255), .Z(n25263) );
  XNOR U25027 ( .A(n25253), .B(n25262), .Z(n25255) );
  XNOR U25028 ( .A(n25264), .B(n25265), .Z(n25253) );
  AND U25029 ( .A(n1100), .B(n25266), .Z(n25265) );
  XOR U25030 ( .A(p_input[1644]), .B(n25264), .Z(n25266) );
  XNOR U25031 ( .A(n25267), .B(n25268), .Z(n25264) );
  AND U25032 ( .A(n1104), .B(n25269), .Z(n25268) );
  XOR U25033 ( .A(n25270), .B(n25271), .Z(n25262) );
  AND U25034 ( .A(n1108), .B(n25261), .Z(n25271) );
  XNOR U25035 ( .A(n25272), .B(n25259), .Z(n25261) );
  XOR U25036 ( .A(n25273), .B(n25274), .Z(n25259) );
  AND U25037 ( .A(n1131), .B(n25275), .Z(n25274) );
  IV U25038 ( .A(n25270), .Z(n25272) );
  XOR U25039 ( .A(n25276), .B(n25277), .Z(n25270) );
  AND U25040 ( .A(n1115), .B(n25269), .Z(n25277) );
  XNOR U25041 ( .A(n25267), .B(n25276), .Z(n25269) );
  XNOR U25042 ( .A(n25278), .B(n25279), .Z(n25267) );
  AND U25043 ( .A(n1119), .B(n25280), .Z(n25279) );
  XOR U25044 ( .A(p_input[1676]), .B(n25278), .Z(n25280) );
  XNOR U25045 ( .A(n25281), .B(n25282), .Z(n25278) );
  AND U25046 ( .A(n1123), .B(n25283), .Z(n25282) );
  XOR U25047 ( .A(n25284), .B(n25285), .Z(n25276) );
  AND U25048 ( .A(n1127), .B(n25275), .Z(n25285) );
  XNOR U25049 ( .A(n25286), .B(n25273), .Z(n25275) );
  XOR U25050 ( .A(n25287), .B(n25288), .Z(n25273) );
  AND U25051 ( .A(n1150), .B(n25289), .Z(n25288) );
  IV U25052 ( .A(n25284), .Z(n25286) );
  XOR U25053 ( .A(n25290), .B(n25291), .Z(n25284) );
  AND U25054 ( .A(n1134), .B(n25283), .Z(n25291) );
  XNOR U25055 ( .A(n25281), .B(n25290), .Z(n25283) );
  XNOR U25056 ( .A(n25292), .B(n25293), .Z(n25281) );
  AND U25057 ( .A(n1138), .B(n25294), .Z(n25293) );
  XOR U25058 ( .A(p_input[1708]), .B(n25292), .Z(n25294) );
  XNOR U25059 ( .A(n25295), .B(n25296), .Z(n25292) );
  AND U25060 ( .A(n1142), .B(n25297), .Z(n25296) );
  XOR U25061 ( .A(n25298), .B(n25299), .Z(n25290) );
  AND U25062 ( .A(n1146), .B(n25289), .Z(n25299) );
  XNOR U25063 ( .A(n25300), .B(n25287), .Z(n25289) );
  XOR U25064 ( .A(n25301), .B(n25302), .Z(n25287) );
  AND U25065 ( .A(n1169), .B(n25303), .Z(n25302) );
  IV U25066 ( .A(n25298), .Z(n25300) );
  XOR U25067 ( .A(n25304), .B(n25305), .Z(n25298) );
  AND U25068 ( .A(n1153), .B(n25297), .Z(n25305) );
  XNOR U25069 ( .A(n25295), .B(n25304), .Z(n25297) );
  XNOR U25070 ( .A(n25306), .B(n25307), .Z(n25295) );
  AND U25071 ( .A(n1157), .B(n25308), .Z(n25307) );
  XOR U25072 ( .A(p_input[1740]), .B(n25306), .Z(n25308) );
  XNOR U25073 ( .A(n25309), .B(n25310), .Z(n25306) );
  AND U25074 ( .A(n1161), .B(n25311), .Z(n25310) );
  XOR U25075 ( .A(n25312), .B(n25313), .Z(n25304) );
  AND U25076 ( .A(n1165), .B(n25303), .Z(n25313) );
  XNOR U25077 ( .A(n25314), .B(n25301), .Z(n25303) );
  XOR U25078 ( .A(n25315), .B(n25316), .Z(n25301) );
  AND U25079 ( .A(n1188), .B(n25317), .Z(n25316) );
  IV U25080 ( .A(n25312), .Z(n25314) );
  XOR U25081 ( .A(n25318), .B(n25319), .Z(n25312) );
  AND U25082 ( .A(n1172), .B(n25311), .Z(n25319) );
  XNOR U25083 ( .A(n25309), .B(n25318), .Z(n25311) );
  XNOR U25084 ( .A(n25320), .B(n25321), .Z(n25309) );
  AND U25085 ( .A(n1176), .B(n25322), .Z(n25321) );
  XOR U25086 ( .A(p_input[1772]), .B(n25320), .Z(n25322) );
  XNOR U25087 ( .A(n25323), .B(n25324), .Z(n25320) );
  AND U25088 ( .A(n1180), .B(n25325), .Z(n25324) );
  XOR U25089 ( .A(n25326), .B(n25327), .Z(n25318) );
  AND U25090 ( .A(n1184), .B(n25317), .Z(n25327) );
  XNOR U25091 ( .A(n25328), .B(n25315), .Z(n25317) );
  XOR U25092 ( .A(n25329), .B(n25330), .Z(n25315) );
  AND U25093 ( .A(n1207), .B(n25331), .Z(n25330) );
  IV U25094 ( .A(n25326), .Z(n25328) );
  XOR U25095 ( .A(n25332), .B(n25333), .Z(n25326) );
  AND U25096 ( .A(n1191), .B(n25325), .Z(n25333) );
  XNOR U25097 ( .A(n25323), .B(n25332), .Z(n25325) );
  XNOR U25098 ( .A(n25334), .B(n25335), .Z(n25323) );
  AND U25099 ( .A(n1195), .B(n25336), .Z(n25335) );
  XOR U25100 ( .A(p_input[1804]), .B(n25334), .Z(n25336) );
  XNOR U25101 ( .A(n25337), .B(n25338), .Z(n25334) );
  AND U25102 ( .A(n1199), .B(n25339), .Z(n25338) );
  XOR U25103 ( .A(n25340), .B(n25341), .Z(n25332) );
  AND U25104 ( .A(n1203), .B(n25331), .Z(n25341) );
  XNOR U25105 ( .A(n25342), .B(n25329), .Z(n25331) );
  XOR U25106 ( .A(n25343), .B(n25344), .Z(n25329) );
  AND U25107 ( .A(n1226), .B(n25345), .Z(n25344) );
  IV U25108 ( .A(n25340), .Z(n25342) );
  XOR U25109 ( .A(n25346), .B(n25347), .Z(n25340) );
  AND U25110 ( .A(n1210), .B(n25339), .Z(n25347) );
  XNOR U25111 ( .A(n25337), .B(n25346), .Z(n25339) );
  XNOR U25112 ( .A(n25348), .B(n25349), .Z(n25337) );
  AND U25113 ( .A(n1214), .B(n25350), .Z(n25349) );
  XOR U25114 ( .A(p_input[1836]), .B(n25348), .Z(n25350) );
  XNOR U25115 ( .A(n25351), .B(n25352), .Z(n25348) );
  AND U25116 ( .A(n1218), .B(n25353), .Z(n25352) );
  XOR U25117 ( .A(n25354), .B(n25355), .Z(n25346) );
  AND U25118 ( .A(n1222), .B(n25345), .Z(n25355) );
  XNOR U25119 ( .A(n25356), .B(n25343), .Z(n25345) );
  XOR U25120 ( .A(n25357), .B(n25358), .Z(n25343) );
  AND U25121 ( .A(n1245), .B(n25359), .Z(n25358) );
  IV U25122 ( .A(n25354), .Z(n25356) );
  XOR U25123 ( .A(n25360), .B(n25361), .Z(n25354) );
  AND U25124 ( .A(n1229), .B(n25353), .Z(n25361) );
  XNOR U25125 ( .A(n25351), .B(n25360), .Z(n25353) );
  XNOR U25126 ( .A(n25362), .B(n25363), .Z(n25351) );
  AND U25127 ( .A(n1233), .B(n25364), .Z(n25363) );
  XOR U25128 ( .A(p_input[1868]), .B(n25362), .Z(n25364) );
  XNOR U25129 ( .A(n25365), .B(n25366), .Z(n25362) );
  AND U25130 ( .A(n1237), .B(n25367), .Z(n25366) );
  XOR U25131 ( .A(n25368), .B(n25369), .Z(n25360) );
  AND U25132 ( .A(n1241), .B(n25359), .Z(n25369) );
  XNOR U25133 ( .A(n25370), .B(n25357), .Z(n25359) );
  XOR U25134 ( .A(n25371), .B(n25372), .Z(n25357) );
  AND U25135 ( .A(n1264), .B(n25373), .Z(n25372) );
  IV U25136 ( .A(n25368), .Z(n25370) );
  XOR U25137 ( .A(n25374), .B(n25375), .Z(n25368) );
  AND U25138 ( .A(n1248), .B(n25367), .Z(n25375) );
  XNOR U25139 ( .A(n25365), .B(n25374), .Z(n25367) );
  XNOR U25140 ( .A(n25376), .B(n25377), .Z(n25365) );
  AND U25141 ( .A(n1252), .B(n25378), .Z(n25377) );
  XOR U25142 ( .A(p_input[1900]), .B(n25376), .Z(n25378) );
  XNOR U25143 ( .A(n25379), .B(n25380), .Z(n25376) );
  AND U25144 ( .A(n1256), .B(n25381), .Z(n25380) );
  XOR U25145 ( .A(n25382), .B(n25383), .Z(n25374) );
  AND U25146 ( .A(n1260), .B(n25373), .Z(n25383) );
  XNOR U25147 ( .A(n25384), .B(n25371), .Z(n25373) );
  XOR U25148 ( .A(n25385), .B(n25386), .Z(n25371) );
  AND U25149 ( .A(n1282), .B(n25387), .Z(n25386) );
  IV U25150 ( .A(n25382), .Z(n25384) );
  XOR U25151 ( .A(n25388), .B(n25389), .Z(n25382) );
  AND U25152 ( .A(n1267), .B(n25381), .Z(n25389) );
  XNOR U25153 ( .A(n25379), .B(n25388), .Z(n25381) );
  XNOR U25154 ( .A(n25390), .B(n25391), .Z(n25379) );
  AND U25155 ( .A(n1271), .B(n25392), .Z(n25391) );
  XOR U25156 ( .A(p_input[1932]), .B(n25390), .Z(n25392) );
  XOR U25157 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n25393), 
        .Z(n25390) );
  AND U25158 ( .A(n1274), .B(n25394), .Z(n25393) );
  XOR U25159 ( .A(n25395), .B(n25396), .Z(n25388) );
  AND U25160 ( .A(n1278), .B(n25387), .Z(n25396) );
  XNOR U25161 ( .A(n25397), .B(n25385), .Z(n25387) );
  XOR U25162 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n25398), .Z(n25385) );
  AND U25163 ( .A(n1290), .B(n25399), .Z(n25398) );
  IV U25164 ( .A(n25395), .Z(n25397) );
  XOR U25165 ( .A(n25400), .B(n25401), .Z(n25395) );
  AND U25166 ( .A(n1285), .B(n25394), .Z(n25401) );
  XOR U25167 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n25400), 
        .Z(n25394) );
  XOR U25168 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(n25402), 
        .Z(n25400) );
  AND U25169 ( .A(n1287), .B(n25399), .Z(n25402) );
  XOR U25170 ( .A(n25403), .B(n25404), .Z(n25399) );
  IV U25171 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n25404)
         );
  IV U25172 ( .A(\knn_comb_/min_val_out[0][12] ), .Z(n25403) );
  XOR U25173 ( .A(n117), .B(n25405), .Z(o[11]) );
  AND U25174 ( .A(n122), .B(n25406), .Z(n117) );
  XOR U25175 ( .A(n118), .B(n25405), .Z(n25406) );
  XOR U25176 ( .A(n25407), .B(n25408), .Z(n25405) );
  AND U25177 ( .A(n142), .B(n25409), .Z(n25408) );
  XOR U25178 ( .A(n25410), .B(n47), .Z(n118) );
  AND U25179 ( .A(n125), .B(n25411), .Z(n47) );
  XOR U25180 ( .A(n48), .B(n25410), .Z(n25411) );
  XOR U25181 ( .A(n25412), .B(n25413), .Z(n48) );
  AND U25182 ( .A(n130), .B(n25414), .Z(n25413) );
  XOR U25183 ( .A(p_input[11]), .B(n25412), .Z(n25414) );
  XNOR U25184 ( .A(n25415), .B(n25416), .Z(n25412) );
  AND U25185 ( .A(n134), .B(n25417), .Z(n25416) );
  XOR U25186 ( .A(n25418), .B(n25419), .Z(n25410) );
  AND U25187 ( .A(n138), .B(n25409), .Z(n25419) );
  XNOR U25188 ( .A(n25420), .B(n25407), .Z(n25409) );
  XOR U25189 ( .A(n25421), .B(n25422), .Z(n25407) );
  AND U25190 ( .A(n162), .B(n25423), .Z(n25422) );
  IV U25191 ( .A(n25418), .Z(n25420) );
  XOR U25192 ( .A(n25424), .B(n25425), .Z(n25418) );
  AND U25193 ( .A(n146), .B(n25417), .Z(n25425) );
  XNOR U25194 ( .A(n25415), .B(n25424), .Z(n25417) );
  XNOR U25195 ( .A(n25426), .B(n25427), .Z(n25415) );
  AND U25196 ( .A(n150), .B(n25428), .Z(n25427) );
  XOR U25197 ( .A(p_input[43]), .B(n25426), .Z(n25428) );
  XNOR U25198 ( .A(n25429), .B(n25430), .Z(n25426) );
  AND U25199 ( .A(n154), .B(n25431), .Z(n25430) );
  XOR U25200 ( .A(n25432), .B(n25433), .Z(n25424) );
  AND U25201 ( .A(n158), .B(n25423), .Z(n25433) );
  XNOR U25202 ( .A(n25434), .B(n25421), .Z(n25423) );
  XOR U25203 ( .A(n25435), .B(n25436), .Z(n25421) );
  AND U25204 ( .A(n181), .B(n25437), .Z(n25436) );
  IV U25205 ( .A(n25432), .Z(n25434) );
  XOR U25206 ( .A(n25438), .B(n25439), .Z(n25432) );
  AND U25207 ( .A(n165), .B(n25431), .Z(n25439) );
  XNOR U25208 ( .A(n25429), .B(n25438), .Z(n25431) );
  XNOR U25209 ( .A(n25440), .B(n25441), .Z(n25429) );
  AND U25210 ( .A(n169), .B(n25442), .Z(n25441) );
  XOR U25211 ( .A(p_input[75]), .B(n25440), .Z(n25442) );
  XNOR U25212 ( .A(n25443), .B(n25444), .Z(n25440) );
  AND U25213 ( .A(n173), .B(n25445), .Z(n25444) );
  XOR U25214 ( .A(n25446), .B(n25447), .Z(n25438) );
  AND U25215 ( .A(n177), .B(n25437), .Z(n25447) );
  XNOR U25216 ( .A(n25448), .B(n25435), .Z(n25437) );
  XOR U25217 ( .A(n25449), .B(n25450), .Z(n25435) );
  AND U25218 ( .A(n200), .B(n25451), .Z(n25450) );
  IV U25219 ( .A(n25446), .Z(n25448) );
  XOR U25220 ( .A(n25452), .B(n25453), .Z(n25446) );
  AND U25221 ( .A(n184), .B(n25445), .Z(n25453) );
  XNOR U25222 ( .A(n25443), .B(n25452), .Z(n25445) );
  XNOR U25223 ( .A(n25454), .B(n25455), .Z(n25443) );
  AND U25224 ( .A(n188), .B(n25456), .Z(n25455) );
  XOR U25225 ( .A(p_input[107]), .B(n25454), .Z(n25456) );
  XNOR U25226 ( .A(n25457), .B(n25458), .Z(n25454) );
  AND U25227 ( .A(n192), .B(n25459), .Z(n25458) );
  XOR U25228 ( .A(n25460), .B(n25461), .Z(n25452) );
  AND U25229 ( .A(n196), .B(n25451), .Z(n25461) );
  XNOR U25230 ( .A(n25462), .B(n25449), .Z(n25451) );
  XOR U25231 ( .A(n25463), .B(n25464), .Z(n25449) );
  AND U25232 ( .A(n219), .B(n25465), .Z(n25464) );
  IV U25233 ( .A(n25460), .Z(n25462) );
  XOR U25234 ( .A(n25466), .B(n25467), .Z(n25460) );
  AND U25235 ( .A(n203), .B(n25459), .Z(n25467) );
  XNOR U25236 ( .A(n25457), .B(n25466), .Z(n25459) );
  XNOR U25237 ( .A(n25468), .B(n25469), .Z(n25457) );
  AND U25238 ( .A(n207), .B(n25470), .Z(n25469) );
  XOR U25239 ( .A(p_input[139]), .B(n25468), .Z(n25470) );
  XNOR U25240 ( .A(n25471), .B(n25472), .Z(n25468) );
  AND U25241 ( .A(n211), .B(n25473), .Z(n25472) );
  XOR U25242 ( .A(n25474), .B(n25475), .Z(n25466) );
  AND U25243 ( .A(n215), .B(n25465), .Z(n25475) );
  XNOR U25244 ( .A(n25476), .B(n25463), .Z(n25465) );
  XOR U25245 ( .A(n25477), .B(n25478), .Z(n25463) );
  AND U25246 ( .A(n238), .B(n25479), .Z(n25478) );
  IV U25247 ( .A(n25474), .Z(n25476) );
  XOR U25248 ( .A(n25480), .B(n25481), .Z(n25474) );
  AND U25249 ( .A(n222), .B(n25473), .Z(n25481) );
  XNOR U25250 ( .A(n25471), .B(n25480), .Z(n25473) );
  XNOR U25251 ( .A(n25482), .B(n25483), .Z(n25471) );
  AND U25252 ( .A(n226), .B(n25484), .Z(n25483) );
  XOR U25253 ( .A(p_input[171]), .B(n25482), .Z(n25484) );
  XNOR U25254 ( .A(n25485), .B(n25486), .Z(n25482) );
  AND U25255 ( .A(n230), .B(n25487), .Z(n25486) );
  XOR U25256 ( .A(n25488), .B(n25489), .Z(n25480) );
  AND U25257 ( .A(n234), .B(n25479), .Z(n25489) );
  XNOR U25258 ( .A(n25490), .B(n25477), .Z(n25479) );
  XOR U25259 ( .A(n25491), .B(n25492), .Z(n25477) );
  AND U25260 ( .A(n257), .B(n25493), .Z(n25492) );
  IV U25261 ( .A(n25488), .Z(n25490) );
  XOR U25262 ( .A(n25494), .B(n25495), .Z(n25488) );
  AND U25263 ( .A(n241), .B(n25487), .Z(n25495) );
  XNOR U25264 ( .A(n25485), .B(n25494), .Z(n25487) );
  XNOR U25265 ( .A(n25496), .B(n25497), .Z(n25485) );
  AND U25266 ( .A(n245), .B(n25498), .Z(n25497) );
  XOR U25267 ( .A(p_input[203]), .B(n25496), .Z(n25498) );
  XNOR U25268 ( .A(n25499), .B(n25500), .Z(n25496) );
  AND U25269 ( .A(n249), .B(n25501), .Z(n25500) );
  XOR U25270 ( .A(n25502), .B(n25503), .Z(n25494) );
  AND U25271 ( .A(n253), .B(n25493), .Z(n25503) );
  XNOR U25272 ( .A(n25504), .B(n25491), .Z(n25493) );
  XOR U25273 ( .A(n25505), .B(n25506), .Z(n25491) );
  AND U25274 ( .A(n276), .B(n25507), .Z(n25506) );
  IV U25275 ( .A(n25502), .Z(n25504) );
  XOR U25276 ( .A(n25508), .B(n25509), .Z(n25502) );
  AND U25277 ( .A(n260), .B(n25501), .Z(n25509) );
  XNOR U25278 ( .A(n25499), .B(n25508), .Z(n25501) );
  XNOR U25279 ( .A(n25510), .B(n25511), .Z(n25499) );
  AND U25280 ( .A(n264), .B(n25512), .Z(n25511) );
  XOR U25281 ( .A(p_input[235]), .B(n25510), .Z(n25512) );
  XNOR U25282 ( .A(n25513), .B(n25514), .Z(n25510) );
  AND U25283 ( .A(n268), .B(n25515), .Z(n25514) );
  XOR U25284 ( .A(n25516), .B(n25517), .Z(n25508) );
  AND U25285 ( .A(n272), .B(n25507), .Z(n25517) );
  XNOR U25286 ( .A(n25518), .B(n25505), .Z(n25507) );
  XOR U25287 ( .A(n25519), .B(n25520), .Z(n25505) );
  AND U25288 ( .A(n295), .B(n25521), .Z(n25520) );
  IV U25289 ( .A(n25516), .Z(n25518) );
  XOR U25290 ( .A(n25522), .B(n25523), .Z(n25516) );
  AND U25291 ( .A(n279), .B(n25515), .Z(n25523) );
  XNOR U25292 ( .A(n25513), .B(n25522), .Z(n25515) );
  XNOR U25293 ( .A(n25524), .B(n25525), .Z(n25513) );
  AND U25294 ( .A(n283), .B(n25526), .Z(n25525) );
  XOR U25295 ( .A(p_input[267]), .B(n25524), .Z(n25526) );
  XNOR U25296 ( .A(n25527), .B(n25528), .Z(n25524) );
  AND U25297 ( .A(n287), .B(n25529), .Z(n25528) );
  XOR U25298 ( .A(n25530), .B(n25531), .Z(n25522) );
  AND U25299 ( .A(n291), .B(n25521), .Z(n25531) );
  XNOR U25300 ( .A(n25532), .B(n25519), .Z(n25521) );
  XOR U25301 ( .A(n25533), .B(n25534), .Z(n25519) );
  AND U25302 ( .A(n314), .B(n25535), .Z(n25534) );
  IV U25303 ( .A(n25530), .Z(n25532) );
  XOR U25304 ( .A(n25536), .B(n25537), .Z(n25530) );
  AND U25305 ( .A(n298), .B(n25529), .Z(n25537) );
  XNOR U25306 ( .A(n25527), .B(n25536), .Z(n25529) );
  XNOR U25307 ( .A(n25538), .B(n25539), .Z(n25527) );
  AND U25308 ( .A(n302), .B(n25540), .Z(n25539) );
  XOR U25309 ( .A(p_input[299]), .B(n25538), .Z(n25540) );
  XNOR U25310 ( .A(n25541), .B(n25542), .Z(n25538) );
  AND U25311 ( .A(n306), .B(n25543), .Z(n25542) );
  XOR U25312 ( .A(n25544), .B(n25545), .Z(n25536) );
  AND U25313 ( .A(n310), .B(n25535), .Z(n25545) );
  XNOR U25314 ( .A(n25546), .B(n25533), .Z(n25535) );
  XOR U25315 ( .A(n25547), .B(n25548), .Z(n25533) );
  AND U25316 ( .A(n333), .B(n25549), .Z(n25548) );
  IV U25317 ( .A(n25544), .Z(n25546) );
  XOR U25318 ( .A(n25550), .B(n25551), .Z(n25544) );
  AND U25319 ( .A(n317), .B(n25543), .Z(n25551) );
  XNOR U25320 ( .A(n25541), .B(n25550), .Z(n25543) );
  XNOR U25321 ( .A(n25552), .B(n25553), .Z(n25541) );
  AND U25322 ( .A(n321), .B(n25554), .Z(n25553) );
  XOR U25323 ( .A(p_input[331]), .B(n25552), .Z(n25554) );
  XNOR U25324 ( .A(n25555), .B(n25556), .Z(n25552) );
  AND U25325 ( .A(n325), .B(n25557), .Z(n25556) );
  XOR U25326 ( .A(n25558), .B(n25559), .Z(n25550) );
  AND U25327 ( .A(n329), .B(n25549), .Z(n25559) );
  XNOR U25328 ( .A(n25560), .B(n25547), .Z(n25549) );
  XOR U25329 ( .A(n25561), .B(n25562), .Z(n25547) );
  AND U25330 ( .A(n352), .B(n25563), .Z(n25562) );
  IV U25331 ( .A(n25558), .Z(n25560) );
  XOR U25332 ( .A(n25564), .B(n25565), .Z(n25558) );
  AND U25333 ( .A(n336), .B(n25557), .Z(n25565) );
  XNOR U25334 ( .A(n25555), .B(n25564), .Z(n25557) );
  XNOR U25335 ( .A(n25566), .B(n25567), .Z(n25555) );
  AND U25336 ( .A(n340), .B(n25568), .Z(n25567) );
  XOR U25337 ( .A(p_input[363]), .B(n25566), .Z(n25568) );
  XNOR U25338 ( .A(n25569), .B(n25570), .Z(n25566) );
  AND U25339 ( .A(n344), .B(n25571), .Z(n25570) );
  XOR U25340 ( .A(n25572), .B(n25573), .Z(n25564) );
  AND U25341 ( .A(n348), .B(n25563), .Z(n25573) );
  XNOR U25342 ( .A(n25574), .B(n25561), .Z(n25563) );
  XOR U25343 ( .A(n25575), .B(n25576), .Z(n25561) );
  AND U25344 ( .A(n371), .B(n25577), .Z(n25576) );
  IV U25345 ( .A(n25572), .Z(n25574) );
  XOR U25346 ( .A(n25578), .B(n25579), .Z(n25572) );
  AND U25347 ( .A(n355), .B(n25571), .Z(n25579) );
  XNOR U25348 ( .A(n25569), .B(n25578), .Z(n25571) );
  XNOR U25349 ( .A(n25580), .B(n25581), .Z(n25569) );
  AND U25350 ( .A(n359), .B(n25582), .Z(n25581) );
  XOR U25351 ( .A(p_input[395]), .B(n25580), .Z(n25582) );
  XNOR U25352 ( .A(n25583), .B(n25584), .Z(n25580) );
  AND U25353 ( .A(n363), .B(n25585), .Z(n25584) );
  XOR U25354 ( .A(n25586), .B(n25587), .Z(n25578) );
  AND U25355 ( .A(n367), .B(n25577), .Z(n25587) );
  XNOR U25356 ( .A(n25588), .B(n25575), .Z(n25577) );
  XOR U25357 ( .A(n25589), .B(n25590), .Z(n25575) );
  AND U25358 ( .A(n390), .B(n25591), .Z(n25590) );
  IV U25359 ( .A(n25586), .Z(n25588) );
  XOR U25360 ( .A(n25592), .B(n25593), .Z(n25586) );
  AND U25361 ( .A(n374), .B(n25585), .Z(n25593) );
  XNOR U25362 ( .A(n25583), .B(n25592), .Z(n25585) );
  XNOR U25363 ( .A(n25594), .B(n25595), .Z(n25583) );
  AND U25364 ( .A(n378), .B(n25596), .Z(n25595) );
  XOR U25365 ( .A(p_input[427]), .B(n25594), .Z(n25596) );
  XNOR U25366 ( .A(n25597), .B(n25598), .Z(n25594) );
  AND U25367 ( .A(n382), .B(n25599), .Z(n25598) );
  XOR U25368 ( .A(n25600), .B(n25601), .Z(n25592) );
  AND U25369 ( .A(n386), .B(n25591), .Z(n25601) );
  XNOR U25370 ( .A(n25602), .B(n25589), .Z(n25591) );
  XOR U25371 ( .A(n25603), .B(n25604), .Z(n25589) );
  AND U25372 ( .A(n409), .B(n25605), .Z(n25604) );
  IV U25373 ( .A(n25600), .Z(n25602) );
  XOR U25374 ( .A(n25606), .B(n25607), .Z(n25600) );
  AND U25375 ( .A(n393), .B(n25599), .Z(n25607) );
  XNOR U25376 ( .A(n25597), .B(n25606), .Z(n25599) );
  XNOR U25377 ( .A(n25608), .B(n25609), .Z(n25597) );
  AND U25378 ( .A(n397), .B(n25610), .Z(n25609) );
  XOR U25379 ( .A(p_input[459]), .B(n25608), .Z(n25610) );
  XNOR U25380 ( .A(n25611), .B(n25612), .Z(n25608) );
  AND U25381 ( .A(n401), .B(n25613), .Z(n25612) );
  XOR U25382 ( .A(n25614), .B(n25615), .Z(n25606) );
  AND U25383 ( .A(n405), .B(n25605), .Z(n25615) );
  XNOR U25384 ( .A(n25616), .B(n25603), .Z(n25605) );
  XOR U25385 ( .A(n25617), .B(n25618), .Z(n25603) );
  AND U25386 ( .A(n428), .B(n25619), .Z(n25618) );
  IV U25387 ( .A(n25614), .Z(n25616) );
  XOR U25388 ( .A(n25620), .B(n25621), .Z(n25614) );
  AND U25389 ( .A(n412), .B(n25613), .Z(n25621) );
  XNOR U25390 ( .A(n25611), .B(n25620), .Z(n25613) );
  XNOR U25391 ( .A(n25622), .B(n25623), .Z(n25611) );
  AND U25392 ( .A(n416), .B(n25624), .Z(n25623) );
  XOR U25393 ( .A(p_input[491]), .B(n25622), .Z(n25624) );
  XNOR U25394 ( .A(n25625), .B(n25626), .Z(n25622) );
  AND U25395 ( .A(n420), .B(n25627), .Z(n25626) );
  XOR U25396 ( .A(n25628), .B(n25629), .Z(n25620) );
  AND U25397 ( .A(n424), .B(n25619), .Z(n25629) );
  XNOR U25398 ( .A(n25630), .B(n25617), .Z(n25619) );
  XOR U25399 ( .A(n25631), .B(n25632), .Z(n25617) );
  AND U25400 ( .A(n447), .B(n25633), .Z(n25632) );
  IV U25401 ( .A(n25628), .Z(n25630) );
  XOR U25402 ( .A(n25634), .B(n25635), .Z(n25628) );
  AND U25403 ( .A(n431), .B(n25627), .Z(n25635) );
  XNOR U25404 ( .A(n25625), .B(n25634), .Z(n25627) );
  XNOR U25405 ( .A(n25636), .B(n25637), .Z(n25625) );
  AND U25406 ( .A(n435), .B(n25638), .Z(n25637) );
  XOR U25407 ( .A(p_input[523]), .B(n25636), .Z(n25638) );
  XNOR U25408 ( .A(n25639), .B(n25640), .Z(n25636) );
  AND U25409 ( .A(n439), .B(n25641), .Z(n25640) );
  XOR U25410 ( .A(n25642), .B(n25643), .Z(n25634) );
  AND U25411 ( .A(n443), .B(n25633), .Z(n25643) );
  XNOR U25412 ( .A(n25644), .B(n25631), .Z(n25633) );
  XOR U25413 ( .A(n25645), .B(n25646), .Z(n25631) );
  AND U25414 ( .A(n466), .B(n25647), .Z(n25646) );
  IV U25415 ( .A(n25642), .Z(n25644) );
  XOR U25416 ( .A(n25648), .B(n25649), .Z(n25642) );
  AND U25417 ( .A(n450), .B(n25641), .Z(n25649) );
  XNOR U25418 ( .A(n25639), .B(n25648), .Z(n25641) );
  XNOR U25419 ( .A(n25650), .B(n25651), .Z(n25639) );
  AND U25420 ( .A(n454), .B(n25652), .Z(n25651) );
  XOR U25421 ( .A(p_input[555]), .B(n25650), .Z(n25652) );
  XNOR U25422 ( .A(n25653), .B(n25654), .Z(n25650) );
  AND U25423 ( .A(n458), .B(n25655), .Z(n25654) );
  XOR U25424 ( .A(n25656), .B(n25657), .Z(n25648) );
  AND U25425 ( .A(n462), .B(n25647), .Z(n25657) );
  XNOR U25426 ( .A(n25658), .B(n25645), .Z(n25647) );
  XOR U25427 ( .A(n25659), .B(n25660), .Z(n25645) );
  AND U25428 ( .A(n485), .B(n25661), .Z(n25660) );
  IV U25429 ( .A(n25656), .Z(n25658) );
  XOR U25430 ( .A(n25662), .B(n25663), .Z(n25656) );
  AND U25431 ( .A(n469), .B(n25655), .Z(n25663) );
  XNOR U25432 ( .A(n25653), .B(n25662), .Z(n25655) );
  XNOR U25433 ( .A(n25664), .B(n25665), .Z(n25653) );
  AND U25434 ( .A(n473), .B(n25666), .Z(n25665) );
  XOR U25435 ( .A(p_input[587]), .B(n25664), .Z(n25666) );
  XNOR U25436 ( .A(n25667), .B(n25668), .Z(n25664) );
  AND U25437 ( .A(n477), .B(n25669), .Z(n25668) );
  XOR U25438 ( .A(n25670), .B(n25671), .Z(n25662) );
  AND U25439 ( .A(n481), .B(n25661), .Z(n25671) );
  XNOR U25440 ( .A(n25672), .B(n25659), .Z(n25661) );
  XOR U25441 ( .A(n25673), .B(n25674), .Z(n25659) );
  AND U25442 ( .A(n504), .B(n25675), .Z(n25674) );
  IV U25443 ( .A(n25670), .Z(n25672) );
  XOR U25444 ( .A(n25676), .B(n25677), .Z(n25670) );
  AND U25445 ( .A(n488), .B(n25669), .Z(n25677) );
  XNOR U25446 ( .A(n25667), .B(n25676), .Z(n25669) );
  XNOR U25447 ( .A(n25678), .B(n25679), .Z(n25667) );
  AND U25448 ( .A(n492), .B(n25680), .Z(n25679) );
  XOR U25449 ( .A(p_input[619]), .B(n25678), .Z(n25680) );
  XNOR U25450 ( .A(n25681), .B(n25682), .Z(n25678) );
  AND U25451 ( .A(n496), .B(n25683), .Z(n25682) );
  XOR U25452 ( .A(n25684), .B(n25685), .Z(n25676) );
  AND U25453 ( .A(n500), .B(n25675), .Z(n25685) );
  XNOR U25454 ( .A(n25686), .B(n25673), .Z(n25675) );
  XOR U25455 ( .A(n25687), .B(n25688), .Z(n25673) );
  AND U25456 ( .A(n523), .B(n25689), .Z(n25688) );
  IV U25457 ( .A(n25684), .Z(n25686) );
  XOR U25458 ( .A(n25690), .B(n25691), .Z(n25684) );
  AND U25459 ( .A(n507), .B(n25683), .Z(n25691) );
  XNOR U25460 ( .A(n25681), .B(n25690), .Z(n25683) );
  XNOR U25461 ( .A(n25692), .B(n25693), .Z(n25681) );
  AND U25462 ( .A(n511), .B(n25694), .Z(n25693) );
  XOR U25463 ( .A(p_input[651]), .B(n25692), .Z(n25694) );
  XNOR U25464 ( .A(n25695), .B(n25696), .Z(n25692) );
  AND U25465 ( .A(n515), .B(n25697), .Z(n25696) );
  XOR U25466 ( .A(n25698), .B(n25699), .Z(n25690) );
  AND U25467 ( .A(n519), .B(n25689), .Z(n25699) );
  XNOR U25468 ( .A(n25700), .B(n25687), .Z(n25689) );
  XOR U25469 ( .A(n25701), .B(n25702), .Z(n25687) );
  AND U25470 ( .A(n542), .B(n25703), .Z(n25702) );
  IV U25471 ( .A(n25698), .Z(n25700) );
  XOR U25472 ( .A(n25704), .B(n25705), .Z(n25698) );
  AND U25473 ( .A(n526), .B(n25697), .Z(n25705) );
  XNOR U25474 ( .A(n25695), .B(n25704), .Z(n25697) );
  XNOR U25475 ( .A(n25706), .B(n25707), .Z(n25695) );
  AND U25476 ( .A(n530), .B(n25708), .Z(n25707) );
  XOR U25477 ( .A(p_input[683]), .B(n25706), .Z(n25708) );
  XNOR U25478 ( .A(n25709), .B(n25710), .Z(n25706) );
  AND U25479 ( .A(n534), .B(n25711), .Z(n25710) );
  XOR U25480 ( .A(n25712), .B(n25713), .Z(n25704) );
  AND U25481 ( .A(n538), .B(n25703), .Z(n25713) );
  XNOR U25482 ( .A(n25714), .B(n25701), .Z(n25703) );
  XOR U25483 ( .A(n25715), .B(n25716), .Z(n25701) );
  AND U25484 ( .A(n561), .B(n25717), .Z(n25716) );
  IV U25485 ( .A(n25712), .Z(n25714) );
  XOR U25486 ( .A(n25718), .B(n25719), .Z(n25712) );
  AND U25487 ( .A(n545), .B(n25711), .Z(n25719) );
  XNOR U25488 ( .A(n25709), .B(n25718), .Z(n25711) );
  XNOR U25489 ( .A(n25720), .B(n25721), .Z(n25709) );
  AND U25490 ( .A(n549), .B(n25722), .Z(n25721) );
  XOR U25491 ( .A(p_input[715]), .B(n25720), .Z(n25722) );
  XNOR U25492 ( .A(n25723), .B(n25724), .Z(n25720) );
  AND U25493 ( .A(n553), .B(n25725), .Z(n25724) );
  XOR U25494 ( .A(n25726), .B(n25727), .Z(n25718) );
  AND U25495 ( .A(n557), .B(n25717), .Z(n25727) );
  XNOR U25496 ( .A(n25728), .B(n25715), .Z(n25717) );
  XOR U25497 ( .A(n25729), .B(n25730), .Z(n25715) );
  AND U25498 ( .A(n580), .B(n25731), .Z(n25730) );
  IV U25499 ( .A(n25726), .Z(n25728) );
  XOR U25500 ( .A(n25732), .B(n25733), .Z(n25726) );
  AND U25501 ( .A(n564), .B(n25725), .Z(n25733) );
  XNOR U25502 ( .A(n25723), .B(n25732), .Z(n25725) );
  XNOR U25503 ( .A(n25734), .B(n25735), .Z(n25723) );
  AND U25504 ( .A(n568), .B(n25736), .Z(n25735) );
  XOR U25505 ( .A(p_input[747]), .B(n25734), .Z(n25736) );
  XNOR U25506 ( .A(n25737), .B(n25738), .Z(n25734) );
  AND U25507 ( .A(n572), .B(n25739), .Z(n25738) );
  XOR U25508 ( .A(n25740), .B(n25741), .Z(n25732) );
  AND U25509 ( .A(n576), .B(n25731), .Z(n25741) );
  XNOR U25510 ( .A(n25742), .B(n25729), .Z(n25731) );
  XOR U25511 ( .A(n25743), .B(n25744), .Z(n25729) );
  AND U25512 ( .A(n599), .B(n25745), .Z(n25744) );
  IV U25513 ( .A(n25740), .Z(n25742) );
  XOR U25514 ( .A(n25746), .B(n25747), .Z(n25740) );
  AND U25515 ( .A(n583), .B(n25739), .Z(n25747) );
  XNOR U25516 ( .A(n25737), .B(n25746), .Z(n25739) );
  XNOR U25517 ( .A(n25748), .B(n25749), .Z(n25737) );
  AND U25518 ( .A(n587), .B(n25750), .Z(n25749) );
  XOR U25519 ( .A(p_input[779]), .B(n25748), .Z(n25750) );
  XNOR U25520 ( .A(n25751), .B(n25752), .Z(n25748) );
  AND U25521 ( .A(n591), .B(n25753), .Z(n25752) );
  XOR U25522 ( .A(n25754), .B(n25755), .Z(n25746) );
  AND U25523 ( .A(n595), .B(n25745), .Z(n25755) );
  XNOR U25524 ( .A(n25756), .B(n25743), .Z(n25745) );
  XOR U25525 ( .A(n25757), .B(n25758), .Z(n25743) );
  AND U25526 ( .A(n618), .B(n25759), .Z(n25758) );
  IV U25527 ( .A(n25754), .Z(n25756) );
  XOR U25528 ( .A(n25760), .B(n25761), .Z(n25754) );
  AND U25529 ( .A(n602), .B(n25753), .Z(n25761) );
  XNOR U25530 ( .A(n25751), .B(n25760), .Z(n25753) );
  XNOR U25531 ( .A(n25762), .B(n25763), .Z(n25751) );
  AND U25532 ( .A(n606), .B(n25764), .Z(n25763) );
  XOR U25533 ( .A(p_input[811]), .B(n25762), .Z(n25764) );
  XNOR U25534 ( .A(n25765), .B(n25766), .Z(n25762) );
  AND U25535 ( .A(n610), .B(n25767), .Z(n25766) );
  XOR U25536 ( .A(n25768), .B(n25769), .Z(n25760) );
  AND U25537 ( .A(n614), .B(n25759), .Z(n25769) );
  XNOR U25538 ( .A(n25770), .B(n25757), .Z(n25759) );
  XOR U25539 ( .A(n25771), .B(n25772), .Z(n25757) );
  AND U25540 ( .A(n637), .B(n25773), .Z(n25772) );
  IV U25541 ( .A(n25768), .Z(n25770) );
  XOR U25542 ( .A(n25774), .B(n25775), .Z(n25768) );
  AND U25543 ( .A(n621), .B(n25767), .Z(n25775) );
  XNOR U25544 ( .A(n25765), .B(n25774), .Z(n25767) );
  XNOR U25545 ( .A(n25776), .B(n25777), .Z(n25765) );
  AND U25546 ( .A(n625), .B(n25778), .Z(n25777) );
  XOR U25547 ( .A(p_input[843]), .B(n25776), .Z(n25778) );
  XNOR U25548 ( .A(n25779), .B(n25780), .Z(n25776) );
  AND U25549 ( .A(n629), .B(n25781), .Z(n25780) );
  XOR U25550 ( .A(n25782), .B(n25783), .Z(n25774) );
  AND U25551 ( .A(n633), .B(n25773), .Z(n25783) );
  XNOR U25552 ( .A(n25784), .B(n25771), .Z(n25773) );
  XOR U25553 ( .A(n25785), .B(n25786), .Z(n25771) );
  AND U25554 ( .A(n656), .B(n25787), .Z(n25786) );
  IV U25555 ( .A(n25782), .Z(n25784) );
  XOR U25556 ( .A(n25788), .B(n25789), .Z(n25782) );
  AND U25557 ( .A(n640), .B(n25781), .Z(n25789) );
  XNOR U25558 ( .A(n25779), .B(n25788), .Z(n25781) );
  XNOR U25559 ( .A(n25790), .B(n25791), .Z(n25779) );
  AND U25560 ( .A(n644), .B(n25792), .Z(n25791) );
  XOR U25561 ( .A(p_input[875]), .B(n25790), .Z(n25792) );
  XNOR U25562 ( .A(n25793), .B(n25794), .Z(n25790) );
  AND U25563 ( .A(n648), .B(n25795), .Z(n25794) );
  XOR U25564 ( .A(n25796), .B(n25797), .Z(n25788) );
  AND U25565 ( .A(n652), .B(n25787), .Z(n25797) );
  XNOR U25566 ( .A(n25798), .B(n25785), .Z(n25787) );
  XOR U25567 ( .A(n25799), .B(n25800), .Z(n25785) );
  AND U25568 ( .A(n675), .B(n25801), .Z(n25800) );
  IV U25569 ( .A(n25796), .Z(n25798) );
  XOR U25570 ( .A(n25802), .B(n25803), .Z(n25796) );
  AND U25571 ( .A(n659), .B(n25795), .Z(n25803) );
  XNOR U25572 ( .A(n25793), .B(n25802), .Z(n25795) );
  XNOR U25573 ( .A(n25804), .B(n25805), .Z(n25793) );
  AND U25574 ( .A(n663), .B(n25806), .Z(n25805) );
  XOR U25575 ( .A(p_input[907]), .B(n25804), .Z(n25806) );
  XNOR U25576 ( .A(n25807), .B(n25808), .Z(n25804) );
  AND U25577 ( .A(n667), .B(n25809), .Z(n25808) );
  XOR U25578 ( .A(n25810), .B(n25811), .Z(n25802) );
  AND U25579 ( .A(n671), .B(n25801), .Z(n25811) );
  XNOR U25580 ( .A(n25812), .B(n25799), .Z(n25801) );
  XOR U25581 ( .A(n25813), .B(n25814), .Z(n25799) );
  AND U25582 ( .A(n694), .B(n25815), .Z(n25814) );
  IV U25583 ( .A(n25810), .Z(n25812) );
  XOR U25584 ( .A(n25816), .B(n25817), .Z(n25810) );
  AND U25585 ( .A(n678), .B(n25809), .Z(n25817) );
  XNOR U25586 ( .A(n25807), .B(n25816), .Z(n25809) );
  XNOR U25587 ( .A(n25818), .B(n25819), .Z(n25807) );
  AND U25588 ( .A(n682), .B(n25820), .Z(n25819) );
  XOR U25589 ( .A(p_input[939]), .B(n25818), .Z(n25820) );
  XNOR U25590 ( .A(n25821), .B(n25822), .Z(n25818) );
  AND U25591 ( .A(n686), .B(n25823), .Z(n25822) );
  XOR U25592 ( .A(n25824), .B(n25825), .Z(n25816) );
  AND U25593 ( .A(n690), .B(n25815), .Z(n25825) );
  XNOR U25594 ( .A(n25826), .B(n25813), .Z(n25815) );
  XOR U25595 ( .A(n25827), .B(n25828), .Z(n25813) );
  AND U25596 ( .A(n713), .B(n25829), .Z(n25828) );
  IV U25597 ( .A(n25824), .Z(n25826) );
  XOR U25598 ( .A(n25830), .B(n25831), .Z(n25824) );
  AND U25599 ( .A(n697), .B(n25823), .Z(n25831) );
  XNOR U25600 ( .A(n25821), .B(n25830), .Z(n25823) );
  XNOR U25601 ( .A(n25832), .B(n25833), .Z(n25821) );
  AND U25602 ( .A(n701), .B(n25834), .Z(n25833) );
  XOR U25603 ( .A(p_input[971]), .B(n25832), .Z(n25834) );
  XNOR U25604 ( .A(n25835), .B(n25836), .Z(n25832) );
  AND U25605 ( .A(n705), .B(n25837), .Z(n25836) );
  XOR U25606 ( .A(n25838), .B(n25839), .Z(n25830) );
  AND U25607 ( .A(n709), .B(n25829), .Z(n25839) );
  XNOR U25608 ( .A(n25840), .B(n25827), .Z(n25829) );
  XOR U25609 ( .A(n25841), .B(n25842), .Z(n25827) );
  AND U25610 ( .A(n732), .B(n25843), .Z(n25842) );
  IV U25611 ( .A(n25838), .Z(n25840) );
  XOR U25612 ( .A(n25844), .B(n25845), .Z(n25838) );
  AND U25613 ( .A(n716), .B(n25837), .Z(n25845) );
  XNOR U25614 ( .A(n25835), .B(n25844), .Z(n25837) );
  XNOR U25615 ( .A(n25846), .B(n25847), .Z(n25835) );
  AND U25616 ( .A(n720), .B(n25848), .Z(n25847) );
  XOR U25617 ( .A(p_input[1003]), .B(n25846), .Z(n25848) );
  XNOR U25618 ( .A(n25849), .B(n25850), .Z(n25846) );
  AND U25619 ( .A(n724), .B(n25851), .Z(n25850) );
  XOR U25620 ( .A(n25852), .B(n25853), .Z(n25844) );
  AND U25621 ( .A(n728), .B(n25843), .Z(n25853) );
  XNOR U25622 ( .A(n25854), .B(n25841), .Z(n25843) );
  XOR U25623 ( .A(n25855), .B(n25856), .Z(n25841) );
  AND U25624 ( .A(n751), .B(n25857), .Z(n25856) );
  IV U25625 ( .A(n25852), .Z(n25854) );
  XOR U25626 ( .A(n25858), .B(n25859), .Z(n25852) );
  AND U25627 ( .A(n735), .B(n25851), .Z(n25859) );
  XNOR U25628 ( .A(n25849), .B(n25858), .Z(n25851) );
  XNOR U25629 ( .A(n25860), .B(n25861), .Z(n25849) );
  AND U25630 ( .A(n739), .B(n25862), .Z(n25861) );
  XOR U25631 ( .A(p_input[1035]), .B(n25860), .Z(n25862) );
  XNOR U25632 ( .A(n25863), .B(n25864), .Z(n25860) );
  AND U25633 ( .A(n743), .B(n25865), .Z(n25864) );
  XOR U25634 ( .A(n25866), .B(n25867), .Z(n25858) );
  AND U25635 ( .A(n747), .B(n25857), .Z(n25867) );
  XNOR U25636 ( .A(n25868), .B(n25855), .Z(n25857) );
  XOR U25637 ( .A(n25869), .B(n25870), .Z(n25855) );
  AND U25638 ( .A(n770), .B(n25871), .Z(n25870) );
  IV U25639 ( .A(n25866), .Z(n25868) );
  XOR U25640 ( .A(n25872), .B(n25873), .Z(n25866) );
  AND U25641 ( .A(n754), .B(n25865), .Z(n25873) );
  XNOR U25642 ( .A(n25863), .B(n25872), .Z(n25865) );
  XNOR U25643 ( .A(n25874), .B(n25875), .Z(n25863) );
  AND U25644 ( .A(n758), .B(n25876), .Z(n25875) );
  XOR U25645 ( .A(p_input[1067]), .B(n25874), .Z(n25876) );
  XNOR U25646 ( .A(n25877), .B(n25878), .Z(n25874) );
  AND U25647 ( .A(n762), .B(n25879), .Z(n25878) );
  XOR U25648 ( .A(n25880), .B(n25881), .Z(n25872) );
  AND U25649 ( .A(n766), .B(n25871), .Z(n25881) );
  XNOR U25650 ( .A(n25882), .B(n25869), .Z(n25871) );
  XOR U25651 ( .A(n25883), .B(n25884), .Z(n25869) );
  AND U25652 ( .A(n789), .B(n25885), .Z(n25884) );
  IV U25653 ( .A(n25880), .Z(n25882) );
  XOR U25654 ( .A(n25886), .B(n25887), .Z(n25880) );
  AND U25655 ( .A(n773), .B(n25879), .Z(n25887) );
  XNOR U25656 ( .A(n25877), .B(n25886), .Z(n25879) );
  XNOR U25657 ( .A(n25888), .B(n25889), .Z(n25877) );
  AND U25658 ( .A(n777), .B(n25890), .Z(n25889) );
  XOR U25659 ( .A(p_input[1099]), .B(n25888), .Z(n25890) );
  XNOR U25660 ( .A(n25891), .B(n25892), .Z(n25888) );
  AND U25661 ( .A(n781), .B(n25893), .Z(n25892) );
  XOR U25662 ( .A(n25894), .B(n25895), .Z(n25886) );
  AND U25663 ( .A(n785), .B(n25885), .Z(n25895) );
  XNOR U25664 ( .A(n25896), .B(n25883), .Z(n25885) );
  XOR U25665 ( .A(n25897), .B(n25898), .Z(n25883) );
  AND U25666 ( .A(n808), .B(n25899), .Z(n25898) );
  IV U25667 ( .A(n25894), .Z(n25896) );
  XOR U25668 ( .A(n25900), .B(n25901), .Z(n25894) );
  AND U25669 ( .A(n792), .B(n25893), .Z(n25901) );
  XNOR U25670 ( .A(n25891), .B(n25900), .Z(n25893) );
  XNOR U25671 ( .A(n25902), .B(n25903), .Z(n25891) );
  AND U25672 ( .A(n796), .B(n25904), .Z(n25903) );
  XOR U25673 ( .A(p_input[1131]), .B(n25902), .Z(n25904) );
  XNOR U25674 ( .A(n25905), .B(n25906), .Z(n25902) );
  AND U25675 ( .A(n800), .B(n25907), .Z(n25906) );
  XOR U25676 ( .A(n25908), .B(n25909), .Z(n25900) );
  AND U25677 ( .A(n804), .B(n25899), .Z(n25909) );
  XNOR U25678 ( .A(n25910), .B(n25897), .Z(n25899) );
  XOR U25679 ( .A(n25911), .B(n25912), .Z(n25897) );
  AND U25680 ( .A(n827), .B(n25913), .Z(n25912) );
  IV U25681 ( .A(n25908), .Z(n25910) );
  XOR U25682 ( .A(n25914), .B(n25915), .Z(n25908) );
  AND U25683 ( .A(n811), .B(n25907), .Z(n25915) );
  XNOR U25684 ( .A(n25905), .B(n25914), .Z(n25907) );
  XNOR U25685 ( .A(n25916), .B(n25917), .Z(n25905) );
  AND U25686 ( .A(n815), .B(n25918), .Z(n25917) );
  XOR U25687 ( .A(p_input[1163]), .B(n25916), .Z(n25918) );
  XNOR U25688 ( .A(n25919), .B(n25920), .Z(n25916) );
  AND U25689 ( .A(n819), .B(n25921), .Z(n25920) );
  XOR U25690 ( .A(n25922), .B(n25923), .Z(n25914) );
  AND U25691 ( .A(n823), .B(n25913), .Z(n25923) );
  XNOR U25692 ( .A(n25924), .B(n25911), .Z(n25913) );
  XOR U25693 ( .A(n25925), .B(n25926), .Z(n25911) );
  AND U25694 ( .A(n846), .B(n25927), .Z(n25926) );
  IV U25695 ( .A(n25922), .Z(n25924) );
  XOR U25696 ( .A(n25928), .B(n25929), .Z(n25922) );
  AND U25697 ( .A(n830), .B(n25921), .Z(n25929) );
  XNOR U25698 ( .A(n25919), .B(n25928), .Z(n25921) );
  XNOR U25699 ( .A(n25930), .B(n25931), .Z(n25919) );
  AND U25700 ( .A(n834), .B(n25932), .Z(n25931) );
  XOR U25701 ( .A(p_input[1195]), .B(n25930), .Z(n25932) );
  XNOR U25702 ( .A(n25933), .B(n25934), .Z(n25930) );
  AND U25703 ( .A(n838), .B(n25935), .Z(n25934) );
  XOR U25704 ( .A(n25936), .B(n25937), .Z(n25928) );
  AND U25705 ( .A(n842), .B(n25927), .Z(n25937) );
  XNOR U25706 ( .A(n25938), .B(n25925), .Z(n25927) );
  XOR U25707 ( .A(n25939), .B(n25940), .Z(n25925) );
  AND U25708 ( .A(n865), .B(n25941), .Z(n25940) );
  IV U25709 ( .A(n25936), .Z(n25938) );
  XOR U25710 ( .A(n25942), .B(n25943), .Z(n25936) );
  AND U25711 ( .A(n849), .B(n25935), .Z(n25943) );
  XNOR U25712 ( .A(n25933), .B(n25942), .Z(n25935) );
  XNOR U25713 ( .A(n25944), .B(n25945), .Z(n25933) );
  AND U25714 ( .A(n853), .B(n25946), .Z(n25945) );
  XOR U25715 ( .A(p_input[1227]), .B(n25944), .Z(n25946) );
  XNOR U25716 ( .A(n25947), .B(n25948), .Z(n25944) );
  AND U25717 ( .A(n857), .B(n25949), .Z(n25948) );
  XOR U25718 ( .A(n25950), .B(n25951), .Z(n25942) );
  AND U25719 ( .A(n861), .B(n25941), .Z(n25951) );
  XNOR U25720 ( .A(n25952), .B(n25939), .Z(n25941) );
  XOR U25721 ( .A(n25953), .B(n25954), .Z(n25939) );
  AND U25722 ( .A(n884), .B(n25955), .Z(n25954) );
  IV U25723 ( .A(n25950), .Z(n25952) );
  XOR U25724 ( .A(n25956), .B(n25957), .Z(n25950) );
  AND U25725 ( .A(n868), .B(n25949), .Z(n25957) );
  XNOR U25726 ( .A(n25947), .B(n25956), .Z(n25949) );
  XNOR U25727 ( .A(n25958), .B(n25959), .Z(n25947) );
  AND U25728 ( .A(n872), .B(n25960), .Z(n25959) );
  XOR U25729 ( .A(p_input[1259]), .B(n25958), .Z(n25960) );
  XNOR U25730 ( .A(n25961), .B(n25962), .Z(n25958) );
  AND U25731 ( .A(n876), .B(n25963), .Z(n25962) );
  XOR U25732 ( .A(n25964), .B(n25965), .Z(n25956) );
  AND U25733 ( .A(n880), .B(n25955), .Z(n25965) );
  XNOR U25734 ( .A(n25966), .B(n25953), .Z(n25955) );
  XOR U25735 ( .A(n25967), .B(n25968), .Z(n25953) );
  AND U25736 ( .A(n903), .B(n25969), .Z(n25968) );
  IV U25737 ( .A(n25964), .Z(n25966) );
  XOR U25738 ( .A(n25970), .B(n25971), .Z(n25964) );
  AND U25739 ( .A(n887), .B(n25963), .Z(n25971) );
  XNOR U25740 ( .A(n25961), .B(n25970), .Z(n25963) );
  XNOR U25741 ( .A(n25972), .B(n25973), .Z(n25961) );
  AND U25742 ( .A(n891), .B(n25974), .Z(n25973) );
  XOR U25743 ( .A(p_input[1291]), .B(n25972), .Z(n25974) );
  XNOR U25744 ( .A(n25975), .B(n25976), .Z(n25972) );
  AND U25745 ( .A(n895), .B(n25977), .Z(n25976) );
  XOR U25746 ( .A(n25978), .B(n25979), .Z(n25970) );
  AND U25747 ( .A(n899), .B(n25969), .Z(n25979) );
  XNOR U25748 ( .A(n25980), .B(n25967), .Z(n25969) );
  XOR U25749 ( .A(n25981), .B(n25982), .Z(n25967) );
  AND U25750 ( .A(n922), .B(n25983), .Z(n25982) );
  IV U25751 ( .A(n25978), .Z(n25980) );
  XOR U25752 ( .A(n25984), .B(n25985), .Z(n25978) );
  AND U25753 ( .A(n906), .B(n25977), .Z(n25985) );
  XNOR U25754 ( .A(n25975), .B(n25984), .Z(n25977) );
  XNOR U25755 ( .A(n25986), .B(n25987), .Z(n25975) );
  AND U25756 ( .A(n910), .B(n25988), .Z(n25987) );
  XOR U25757 ( .A(p_input[1323]), .B(n25986), .Z(n25988) );
  XNOR U25758 ( .A(n25989), .B(n25990), .Z(n25986) );
  AND U25759 ( .A(n914), .B(n25991), .Z(n25990) );
  XOR U25760 ( .A(n25992), .B(n25993), .Z(n25984) );
  AND U25761 ( .A(n918), .B(n25983), .Z(n25993) );
  XNOR U25762 ( .A(n25994), .B(n25981), .Z(n25983) );
  XOR U25763 ( .A(n25995), .B(n25996), .Z(n25981) );
  AND U25764 ( .A(n941), .B(n25997), .Z(n25996) );
  IV U25765 ( .A(n25992), .Z(n25994) );
  XOR U25766 ( .A(n25998), .B(n25999), .Z(n25992) );
  AND U25767 ( .A(n925), .B(n25991), .Z(n25999) );
  XNOR U25768 ( .A(n25989), .B(n25998), .Z(n25991) );
  XNOR U25769 ( .A(n26000), .B(n26001), .Z(n25989) );
  AND U25770 ( .A(n929), .B(n26002), .Z(n26001) );
  XOR U25771 ( .A(p_input[1355]), .B(n26000), .Z(n26002) );
  XNOR U25772 ( .A(n26003), .B(n26004), .Z(n26000) );
  AND U25773 ( .A(n933), .B(n26005), .Z(n26004) );
  XOR U25774 ( .A(n26006), .B(n26007), .Z(n25998) );
  AND U25775 ( .A(n937), .B(n25997), .Z(n26007) );
  XNOR U25776 ( .A(n26008), .B(n25995), .Z(n25997) );
  XOR U25777 ( .A(n26009), .B(n26010), .Z(n25995) );
  AND U25778 ( .A(n960), .B(n26011), .Z(n26010) );
  IV U25779 ( .A(n26006), .Z(n26008) );
  XOR U25780 ( .A(n26012), .B(n26013), .Z(n26006) );
  AND U25781 ( .A(n944), .B(n26005), .Z(n26013) );
  XNOR U25782 ( .A(n26003), .B(n26012), .Z(n26005) );
  XNOR U25783 ( .A(n26014), .B(n26015), .Z(n26003) );
  AND U25784 ( .A(n948), .B(n26016), .Z(n26015) );
  XOR U25785 ( .A(p_input[1387]), .B(n26014), .Z(n26016) );
  XNOR U25786 ( .A(n26017), .B(n26018), .Z(n26014) );
  AND U25787 ( .A(n952), .B(n26019), .Z(n26018) );
  XOR U25788 ( .A(n26020), .B(n26021), .Z(n26012) );
  AND U25789 ( .A(n956), .B(n26011), .Z(n26021) );
  XNOR U25790 ( .A(n26022), .B(n26009), .Z(n26011) );
  XOR U25791 ( .A(n26023), .B(n26024), .Z(n26009) );
  AND U25792 ( .A(n979), .B(n26025), .Z(n26024) );
  IV U25793 ( .A(n26020), .Z(n26022) );
  XOR U25794 ( .A(n26026), .B(n26027), .Z(n26020) );
  AND U25795 ( .A(n963), .B(n26019), .Z(n26027) );
  XNOR U25796 ( .A(n26017), .B(n26026), .Z(n26019) );
  XNOR U25797 ( .A(n26028), .B(n26029), .Z(n26017) );
  AND U25798 ( .A(n967), .B(n26030), .Z(n26029) );
  XOR U25799 ( .A(p_input[1419]), .B(n26028), .Z(n26030) );
  XNOR U25800 ( .A(n26031), .B(n26032), .Z(n26028) );
  AND U25801 ( .A(n971), .B(n26033), .Z(n26032) );
  XOR U25802 ( .A(n26034), .B(n26035), .Z(n26026) );
  AND U25803 ( .A(n975), .B(n26025), .Z(n26035) );
  XNOR U25804 ( .A(n26036), .B(n26023), .Z(n26025) );
  XOR U25805 ( .A(n26037), .B(n26038), .Z(n26023) );
  AND U25806 ( .A(n998), .B(n26039), .Z(n26038) );
  IV U25807 ( .A(n26034), .Z(n26036) );
  XOR U25808 ( .A(n26040), .B(n26041), .Z(n26034) );
  AND U25809 ( .A(n982), .B(n26033), .Z(n26041) );
  XNOR U25810 ( .A(n26031), .B(n26040), .Z(n26033) );
  XNOR U25811 ( .A(n26042), .B(n26043), .Z(n26031) );
  AND U25812 ( .A(n986), .B(n26044), .Z(n26043) );
  XOR U25813 ( .A(p_input[1451]), .B(n26042), .Z(n26044) );
  XNOR U25814 ( .A(n26045), .B(n26046), .Z(n26042) );
  AND U25815 ( .A(n990), .B(n26047), .Z(n26046) );
  XOR U25816 ( .A(n26048), .B(n26049), .Z(n26040) );
  AND U25817 ( .A(n994), .B(n26039), .Z(n26049) );
  XNOR U25818 ( .A(n26050), .B(n26037), .Z(n26039) );
  XOR U25819 ( .A(n26051), .B(n26052), .Z(n26037) );
  AND U25820 ( .A(n1017), .B(n26053), .Z(n26052) );
  IV U25821 ( .A(n26048), .Z(n26050) );
  XOR U25822 ( .A(n26054), .B(n26055), .Z(n26048) );
  AND U25823 ( .A(n1001), .B(n26047), .Z(n26055) );
  XNOR U25824 ( .A(n26045), .B(n26054), .Z(n26047) );
  XNOR U25825 ( .A(n26056), .B(n26057), .Z(n26045) );
  AND U25826 ( .A(n1005), .B(n26058), .Z(n26057) );
  XOR U25827 ( .A(p_input[1483]), .B(n26056), .Z(n26058) );
  XNOR U25828 ( .A(n26059), .B(n26060), .Z(n26056) );
  AND U25829 ( .A(n1009), .B(n26061), .Z(n26060) );
  XOR U25830 ( .A(n26062), .B(n26063), .Z(n26054) );
  AND U25831 ( .A(n1013), .B(n26053), .Z(n26063) );
  XNOR U25832 ( .A(n26064), .B(n26051), .Z(n26053) );
  XOR U25833 ( .A(n26065), .B(n26066), .Z(n26051) );
  AND U25834 ( .A(n1036), .B(n26067), .Z(n26066) );
  IV U25835 ( .A(n26062), .Z(n26064) );
  XOR U25836 ( .A(n26068), .B(n26069), .Z(n26062) );
  AND U25837 ( .A(n1020), .B(n26061), .Z(n26069) );
  XNOR U25838 ( .A(n26059), .B(n26068), .Z(n26061) );
  XNOR U25839 ( .A(n26070), .B(n26071), .Z(n26059) );
  AND U25840 ( .A(n1024), .B(n26072), .Z(n26071) );
  XOR U25841 ( .A(p_input[1515]), .B(n26070), .Z(n26072) );
  XNOR U25842 ( .A(n26073), .B(n26074), .Z(n26070) );
  AND U25843 ( .A(n1028), .B(n26075), .Z(n26074) );
  XOR U25844 ( .A(n26076), .B(n26077), .Z(n26068) );
  AND U25845 ( .A(n1032), .B(n26067), .Z(n26077) );
  XNOR U25846 ( .A(n26078), .B(n26065), .Z(n26067) );
  XOR U25847 ( .A(n26079), .B(n26080), .Z(n26065) );
  AND U25848 ( .A(n1055), .B(n26081), .Z(n26080) );
  IV U25849 ( .A(n26076), .Z(n26078) );
  XOR U25850 ( .A(n26082), .B(n26083), .Z(n26076) );
  AND U25851 ( .A(n1039), .B(n26075), .Z(n26083) );
  XNOR U25852 ( .A(n26073), .B(n26082), .Z(n26075) );
  XNOR U25853 ( .A(n26084), .B(n26085), .Z(n26073) );
  AND U25854 ( .A(n1043), .B(n26086), .Z(n26085) );
  XOR U25855 ( .A(p_input[1547]), .B(n26084), .Z(n26086) );
  XNOR U25856 ( .A(n26087), .B(n26088), .Z(n26084) );
  AND U25857 ( .A(n1047), .B(n26089), .Z(n26088) );
  XOR U25858 ( .A(n26090), .B(n26091), .Z(n26082) );
  AND U25859 ( .A(n1051), .B(n26081), .Z(n26091) );
  XNOR U25860 ( .A(n26092), .B(n26079), .Z(n26081) );
  XOR U25861 ( .A(n26093), .B(n26094), .Z(n26079) );
  AND U25862 ( .A(n1074), .B(n26095), .Z(n26094) );
  IV U25863 ( .A(n26090), .Z(n26092) );
  XOR U25864 ( .A(n26096), .B(n26097), .Z(n26090) );
  AND U25865 ( .A(n1058), .B(n26089), .Z(n26097) );
  XNOR U25866 ( .A(n26087), .B(n26096), .Z(n26089) );
  XNOR U25867 ( .A(n26098), .B(n26099), .Z(n26087) );
  AND U25868 ( .A(n1062), .B(n26100), .Z(n26099) );
  XOR U25869 ( .A(p_input[1579]), .B(n26098), .Z(n26100) );
  XNOR U25870 ( .A(n26101), .B(n26102), .Z(n26098) );
  AND U25871 ( .A(n1066), .B(n26103), .Z(n26102) );
  XOR U25872 ( .A(n26104), .B(n26105), .Z(n26096) );
  AND U25873 ( .A(n1070), .B(n26095), .Z(n26105) );
  XNOR U25874 ( .A(n26106), .B(n26093), .Z(n26095) );
  XOR U25875 ( .A(n26107), .B(n26108), .Z(n26093) );
  AND U25876 ( .A(n1093), .B(n26109), .Z(n26108) );
  IV U25877 ( .A(n26104), .Z(n26106) );
  XOR U25878 ( .A(n26110), .B(n26111), .Z(n26104) );
  AND U25879 ( .A(n1077), .B(n26103), .Z(n26111) );
  XNOR U25880 ( .A(n26101), .B(n26110), .Z(n26103) );
  XNOR U25881 ( .A(n26112), .B(n26113), .Z(n26101) );
  AND U25882 ( .A(n1081), .B(n26114), .Z(n26113) );
  XOR U25883 ( .A(p_input[1611]), .B(n26112), .Z(n26114) );
  XNOR U25884 ( .A(n26115), .B(n26116), .Z(n26112) );
  AND U25885 ( .A(n1085), .B(n26117), .Z(n26116) );
  XOR U25886 ( .A(n26118), .B(n26119), .Z(n26110) );
  AND U25887 ( .A(n1089), .B(n26109), .Z(n26119) );
  XNOR U25888 ( .A(n26120), .B(n26107), .Z(n26109) );
  XOR U25889 ( .A(n26121), .B(n26122), .Z(n26107) );
  AND U25890 ( .A(n1112), .B(n26123), .Z(n26122) );
  IV U25891 ( .A(n26118), .Z(n26120) );
  XOR U25892 ( .A(n26124), .B(n26125), .Z(n26118) );
  AND U25893 ( .A(n1096), .B(n26117), .Z(n26125) );
  XNOR U25894 ( .A(n26115), .B(n26124), .Z(n26117) );
  XNOR U25895 ( .A(n26126), .B(n26127), .Z(n26115) );
  AND U25896 ( .A(n1100), .B(n26128), .Z(n26127) );
  XOR U25897 ( .A(p_input[1643]), .B(n26126), .Z(n26128) );
  XNOR U25898 ( .A(n26129), .B(n26130), .Z(n26126) );
  AND U25899 ( .A(n1104), .B(n26131), .Z(n26130) );
  XOR U25900 ( .A(n26132), .B(n26133), .Z(n26124) );
  AND U25901 ( .A(n1108), .B(n26123), .Z(n26133) );
  XNOR U25902 ( .A(n26134), .B(n26121), .Z(n26123) );
  XOR U25903 ( .A(n26135), .B(n26136), .Z(n26121) );
  AND U25904 ( .A(n1131), .B(n26137), .Z(n26136) );
  IV U25905 ( .A(n26132), .Z(n26134) );
  XOR U25906 ( .A(n26138), .B(n26139), .Z(n26132) );
  AND U25907 ( .A(n1115), .B(n26131), .Z(n26139) );
  XNOR U25908 ( .A(n26129), .B(n26138), .Z(n26131) );
  XNOR U25909 ( .A(n26140), .B(n26141), .Z(n26129) );
  AND U25910 ( .A(n1119), .B(n26142), .Z(n26141) );
  XOR U25911 ( .A(p_input[1675]), .B(n26140), .Z(n26142) );
  XNOR U25912 ( .A(n26143), .B(n26144), .Z(n26140) );
  AND U25913 ( .A(n1123), .B(n26145), .Z(n26144) );
  XOR U25914 ( .A(n26146), .B(n26147), .Z(n26138) );
  AND U25915 ( .A(n1127), .B(n26137), .Z(n26147) );
  XNOR U25916 ( .A(n26148), .B(n26135), .Z(n26137) );
  XOR U25917 ( .A(n26149), .B(n26150), .Z(n26135) );
  AND U25918 ( .A(n1150), .B(n26151), .Z(n26150) );
  IV U25919 ( .A(n26146), .Z(n26148) );
  XOR U25920 ( .A(n26152), .B(n26153), .Z(n26146) );
  AND U25921 ( .A(n1134), .B(n26145), .Z(n26153) );
  XNOR U25922 ( .A(n26143), .B(n26152), .Z(n26145) );
  XNOR U25923 ( .A(n26154), .B(n26155), .Z(n26143) );
  AND U25924 ( .A(n1138), .B(n26156), .Z(n26155) );
  XOR U25925 ( .A(p_input[1707]), .B(n26154), .Z(n26156) );
  XNOR U25926 ( .A(n26157), .B(n26158), .Z(n26154) );
  AND U25927 ( .A(n1142), .B(n26159), .Z(n26158) );
  XOR U25928 ( .A(n26160), .B(n26161), .Z(n26152) );
  AND U25929 ( .A(n1146), .B(n26151), .Z(n26161) );
  XNOR U25930 ( .A(n26162), .B(n26149), .Z(n26151) );
  XOR U25931 ( .A(n26163), .B(n26164), .Z(n26149) );
  AND U25932 ( .A(n1169), .B(n26165), .Z(n26164) );
  IV U25933 ( .A(n26160), .Z(n26162) );
  XOR U25934 ( .A(n26166), .B(n26167), .Z(n26160) );
  AND U25935 ( .A(n1153), .B(n26159), .Z(n26167) );
  XNOR U25936 ( .A(n26157), .B(n26166), .Z(n26159) );
  XNOR U25937 ( .A(n26168), .B(n26169), .Z(n26157) );
  AND U25938 ( .A(n1157), .B(n26170), .Z(n26169) );
  XOR U25939 ( .A(p_input[1739]), .B(n26168), .Z(n26170) );
  XNOR U25940 ( .A(n26171), .B(n26172), .Z(n26168) );
  AND U25941 ( .A(n1161), .B(n26173), .Z(n26172) );
  XOR U25942 ( .A(n26174), .B(n26175), .Z(n26166) );
  AND U25943 ( .A(n1165), .B(n26165), .Z(n26175) );
  XNOR U25944 ( .A(n26176), .B(n26163), .Z(n26165) );
  XOR U25945 ( .A(n26177), .B(n26178), .Z(n26163) );
  AND U25946 ( .A(n1188), .B(n26179), .Z(n26178) );
  IV U25947 ( .A(n26174), .Z(n26176) );
  XOR U25948 ( .A(n26180), .B(n26181), .Z(n26174) );
  AND U25949 ( .A(n1172), .B(n26173), .Z(n26181) );
  XNOR U25950 ( .A(n26171), .B(n26180), .Z(n26173) );
  XNOR U25951 ( .A(n26182), .B(n26183), .Z(n26171) );
  AND U25952 ( .A(n1176), .B(n26184), .Z(n26183) );
  XOR U25953 ( .A(p_input[1771]), .B(n26182), .Z(n26184) );
  XNOR U25954 ( .A(n26185), .B(n26186), .Z(n26182) );
  AND U25955 ( .A(n1180), .B(n26187), .Z(n26186) );
  XOR U25956 ( .A(n26188), .B(n26189), .Z(n26180) );
  AND U25957 ( .A(n1184), .B(n26179), .Z(n26189) );
  XNOR U25958 ( .A(n26190), .B(n26177), .Z(n26179) );
  XOR U25959 ( .A(n26191), .B(n26192), .Z(n26177) );
  AND U25960 ( .A(n1207), .B(n26193), .Z(n26192) );
  IV U25961 ( .A(n26188), .Z(n26190) );
  XOR U25962 ( .A(n26194), .B(n26195), .Z(n26188) );
  AND U25963 ( .A(n1191), .B(n26187), .Z(n26195) );
  XNOR U25964 ( .A(n26185), .B(n26194), .Z(n26187) );
  XNOR U25965 ( .A(n26196), .B(n26197), .Z(n26185) );
  AND U25966 ( .A(n1195), .B(n26198), .Z(n26197) );
  XOR U25967 ( .A(p_input[1803]), .B(n26196), .Z(n26198) );
  XNOR U25968 ( .A(n26199), .B(n26200), .Z(n26196) );
  AND U25969 ( .A(n1199), .B(n26201), .Z(n26200) );
  XOR U25970 ( .A(n26202), .B(n26203), .Z(n26194) );
  AND U25971 ( .A(n1203), .B(n26193), .Z(n26203) );
  XNOR U25972 ( .A(n26204), .B(n26191), .Z(n26193) );
  XOR U25973 ( .A(n26205), .B(n26206), .Z(n26191) );
  AND U25974 ( .A(n1226), .B(n26207), .Z(n26206) );
  IV U25975 ( .A(n26202), .Z(n26204) );
  XOR U25976 ( .A(n26208), .B(n26209), .Z(n26202) );
  AND U25977 ( .A(n1210), .B(n26201), .Z(n26209) );
  XNOR U25978 ( .A(n26199), .B(n26208), .Z(n26201) );
  XNOR U25979 ( .A(n26210), .B(n26211), .Z(n26199) );
  AND U25980 ( .A(n1214), .B(n26212), .Z(n26211) );
  XOR U25981 ( .A(p_input[1835]), .B(n26210), .Z(n26212) );
  XNOR U25982 ( .A(n26213), .B(n26214), .Z(n26210) );
  AND U25983 ( .A(n1218), .B(n26215), .Z(n26214) );
  XOR U25984 ( .A(n26216), .B(n26217), .Z(n26208) );
  AND U25985 ( .A(n1222), .B(n26207), .Z(n26217) );
  XNOR U25986 ( .A(n26218), .B(n26205), .Z(n26207) );
  XOR U25987 ( .A(n26219), .B(n26220), .Z(n26205) );
  AND U25988 ( .A(n1245), .B(n26221), .Z(n26220) );
  IV U25989 ( .A(n26216), .Z(n26218) );
  XOR U25990 ( .A(n26222), .B(n26223), .Z(n26216) );
  AND U25991 ( .A(n1229), .B(n26215), .Z(n26223) );
  XNOR U25992 ( .A(n26213), .B(n26222), .Z(n26215) );
  XNOR U25993 ( .A(n26224), .B(n26225), .Z(n26213) );
  AND U25994 ( .A(n1233), .B(n26226), .Z(n26225) );
  XOR U25995 ( .A(p_input[1867]), .B(n26224), .Z(n26226) );
  XNOR U25996 ( .A(n26227), .B(n26228), .Z(n26224) );
  AND U25997 ( .A(n1237), .B(n26229), .Z(n26228) );
  XOR U25998 ( .A(n26230), .B(n26231), .Z(n26222) );
  AND U25999 ( .A(n1241), .B(n26221), .Z(n26231) );
  XNOR U26000 ( .A(n26232), .B(n26219), .Z(n26221) );
  XOR U26001 ( .A(n26233), .B(n26234), .Z(n26219) );
  AND U26002 ( .A(n1264), .B(n26235), .Z(n26234) );
  IV U26003 ( .A(n26230), .Z(n26232) );
  XOR U26004 ( .A(n26236), .B(n26237), .Z(n26230) );
  AND U26005 ( .A(n1248), .B(n26229), .Z(n26237) );
  XNOR U26006 ( .A(n26227), .B(n26236), .Z(n26229) );
  XNOR U26007 ( .A(n26238), .B(n26239), .Z(n26227) );
  AND U26008 ( .A(n1252), .B(n26240), .Z(n26239) );
  XOR U26009 ( .A(p_input[1899]), .B(n26238), .Z(n26240) );
  XNOR U26010 ( .A(n26241), .B(n26242), .Z(n26238) );
  AND U26011 ( .A(n1256), .B(n26243), .Z(n26242) );
  XOR U26012 ( .A(n26244), .B(n26245), .Z(n26236) );
  AND U26013 ( .A(n1260), .B(n26235), .Z(n26245) );
  XNOR U26014 ( .A(n26246), .B(n26233), .Z(n26235) );
  XOR U26015 ( .A(n26247), .B(n26248), .Z(n26233) );
  AND U26016 ( .A(n1282), .B(n26249), .Z(n26248) );
  IV U26017 ( .A(n26244), .Z(n26246) );
  XOR U26018 ( .A(n26250), .B(n26251), .Z(n26244) );
  AND U26019 ( .A(n1267), .B(n26243), .Z(n26251) );
  XNOR U26020 ( .A(n26241), .B(n26250), .Z(n26243) );
  XNOR U26021 ( .A(n26252), .B(n26253), .Z(n26241) );
  AND U26022 ( .A(n1271), .B(n26254), .Z(n26253) );
  XOR U26023 ( .A(p_input[1931]), .B(n26252), .Z(n26254) );
  XOR U26024 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n26255), 
        .Z(n26252) );
  AND U26025 ( .A(n1274), .B(n26256), .Z(n26255) );
  XOR U26026 ( .A(n26257), .B(n26258), .Z(n26250) );
  AND U26027 ( .A(n1278), .B(n26249), .Z(n26258) );
  XNOR U26028 ( .A(n26259), .B(n26247), .Z(n26249) );
  XOR U26029 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n26260), .Z(n26247) );
  AND U26030 ( .A(n1290), .B(n26261), .Z(n26260) );
  IV U26031 ( .A(n26257), .Z(n26259) );
  XOR U26032 ( .A(n26262), .B(n26263), .Z(n26257) );
  AND U26033 ( .A(n1285), .B(n26256), .Z(n26263) );
  XOR U26034 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n26262), 
        .Z(n26256) );
  XOR U26035 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n26264), 
        .Z(n26262) );
  AND U26036 ( .A(n1287), .B(n26261), .Z(n26264) );
  XOR U26037 ( .A(\knn_comb_/min_val_out[0][11] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n26261) );
  XOR U26038 ( .A(n119), .B(n26265), .Z(o[10]) );
  AND U26039 ( .A(n122), .B(n26266), .Z(n119) );
  XOR U26040 ( .A(n120), .B(n26265), .Z(n26266) );
  XOR U26041 ( .A(n26267), .B(n26268), .Z(n26265) );
  AND U26042 ( .A(n142), .B(n26269), .Z(n26268) );
  XOR U26043 ( .A(n26270), .B(n49), .Z(n120) );
  AND U26044 ( .A(n125), .B(n26271), .Z(n49) );
  XOR U26045 ( .A(n50), .B(n26270), .Z(n26271) );
  XOR U26046 ( .A(n26272), .B(n26273), .Z(n50) );
  AND U26047 ( .A(n130), .B(n26274), .Z(n26273) );
  XOR U26048 ( .A(p_input[10]), .B(n26272), .Z(n26274) );
  XNOR U26049 ( .A(n26275), .B(n26276), .Z(n26272) );
  AND U26050 ( .A(n134), .B(n26277), .Z(n26276) );
  XOR U26051 ( .A(n26278), .B(n26279), .Z(n26270) );
  AND U26052 ( .A(n138), .B(n26269), .Z(n26279) );
  XNOR U26053 ( .A(n26280), .B(n26267), .Z(n26269) );
  XOR U26054 ( .A(n26281), .B(n26282), .Z(n26267) );
  AND U26055 ( .A(n162), .B(n26283), .Z(n26282) );
  IV U26056 ( .A(n26278), .Z(n26280) );
  XOR U26057 ( .A(n26284), .B(n26285), .Z(n26278) );
  AND U26058 ( .A(n146), .B(n26277), .Z(n26285) );
  XNOR U26059 ( .A(n26275), .B(n26284), .Z(n26277) );
  XNOR U26060 ( .A(n26286), .B(n26287), .Z(n26275) );
  AND U26061 ( .A(n150), .B(n26288), .Z(n26287) );
  XOR U26062 ( .A(p_input[42]), .B(n26286), .Z(n26288) );
  XNOR U26063 ( .A(n26289), .B(n26290), .Z(n26286) );
  AND U26064 ( .A(n154), .B(n26291), .Z(n26290) );
  XOR U26065 ( .A(n26292), .B(n26293), .Z(n26284) );
  AND U26066 ( .A(n158), .B(n26283), .Z(n26293) );
  XNOR U26067 ( .A(n26294), .B(n26281), .Z(n26283) );
  XOR U26068 ( .A(n26295), .B(n26296), .Z(n26281) );
  AND U26069 ( .A(n181), .B(n26297), .Z(n26296) );
  IV U26070 ( .A(n26292), .Z(n26294) );
  XOR U26071 ( .A(n26298), .B(n26299), .Z(n26292) );
  AND U26072 ( .A(n165), .B(n26291), .Z(n26299) );
  XNOR U26073 ( .A(n26289), .B(n26298), .Z(n26291) );
  XNOR U26074 ( .A(n26300), .B(n26301), .Z(n26289) );
  AND U26075 ( .A(n169), .B(n26302), .Z(n26301) );
  XOR U26076 ( .A(p_input[74]), .B(n26300), .Z(n26302) );
  XNOR U26077 ( .A(n26303), .B(n26304), .Z(n26300) );
  AND U26078 ( .A(n173), .B(n26305), .Z(n26304) );
  XOR U26079 ( .A(n26306), .B(n26307), .Z(n26298) );
  AND U26080 ( .A(n177), .B(n26297), .Z(n26307) );
  XNOR U26081 ( .A(n26308), .B(n26295), .Z(n26297) );
  XOR U26082 ( .A(n26309), .B(n26310), .Z(n26295) );
  AND U26083 ( .A(n200), .B(n26311), .Z(n26310) );
  IV U26084 ( .A(n26306), .Z(n26308) );
  XOR U26085 ( .A(n26312), .B(n26313), .Z(n26306) );
  AND U26086 ( .A(n184), .B(n26305), .Z(n26313) );
  XNOR U26087 ( .A(n26303), .B(n26312), .Z(n26305) );
  XNOR U26088 ( .A(n26314), .B(n26315), .Z(n26303) );
  AND U26089 ( .A(n188), .B(n26316), .Z(n26315) );
  XOR U26090 ( .A(p_input[106]), .B(n26314), .Z(n26316) );
  XNOR U26091 ( .A(n26317), .B(n26318), .Z(n26314) );
  AND U26092 ( .A(n192), .B(n26319), .Z(n26318) );
  XOR U26093 ( .A(n26320), .B(n26321), .Z(n26312) );
  AND U26094 ( .A(n196), .B(n26311), .Z(n26321) );
  XNOR U26095 ( .A(n26322), .B(n26309), .Z(n26311) );
  XOR U26096 ( .A(n26323), .B(n26324), .Z(n26309) );
  AND U26097 ( .A(n219), .B(n26325), .Z(n26324) );
  IV U26098 ( .A(n26320), .Z(n26322) );
  XOR U26099 ( .A(n26326), .B(n26327), .Z(n26320) );
  AND U26100 ( .A(n203), .B(n26319), .Z(n26327) );
  XNOR U26101 ( .A(n26317), .B(n26326), .Z(n26319) );
  XNOR U26102 ( .A(n26328), .B(n26329), .Z(n26317) );
  AND U26103 ( .A(n207), .B(n26330), .Z(n26329) );
  XOR U26104 ( .A(p_input[138]), .B(n26328), .Z(n26330) );
  XNOR U26105 ( .A(n26331), .B(n26332), .Z(n26328) );
  AND U26106 ( .A(n211), .B(n26333), .Z(n26332) );
  XOR U26107 ( .A(n26334), .B(n26335), .Z(n26326) );
  AND U26108 ( .A(n215), .B(n26325), .Z(n26335) );
  XNOR U26109 ( .A(n26336), .B(n26323), .Z(n26325) );
  XOR U26110 ( .A(n26337), .B(n26338), .Z(n26323) );
  AND U26111 ( .A(n238), .B(n26339), .Z(n26338) );
  IV U26112 ( .A(n26334), .Z(n26336) );
  XOR U26113 ( .A(n26340), .B(n26341), .Z(n26334) );
  AND U26114 ( .A(n222), .B(n26333), .Z(n26341) );
  XNOR U26115 ( .A(n26331), .B(n26340), .Z(n26333) );
  XNOR U26116 ( .A(n26342), .B(n26343), .Z(n26331) );
  AND U26117 ( .A(n226), .B(n26344), .Z(n26343) );
  XOR U26118 ( .A(p_input[170]), .B(n26342), .Z(n26344) );
  XNOR U26119 ( .A(n26345), .B(n26346), .Z(n26342) );
  AND U26120 ( .A(n230), .B(n26347), .Z(n26346) );
  XOR U26121 ( .A(n26348), .B(n26349), .Z(n26340) );
  AND U26122 ( .A(n234), .B(n26339), .Z(n26349) );
  XNOR U26123 ( .A(n26350), .B(n26337), .Z(n26339) );
  XOR U26124 ( .A(n26351), .B(n26352), .Z(n26337) );
  AND U26125 ( .A(n257), .B(n26353), .Z(n26352) );
  IV U26126 ( .A(n26348), .Z(n26350) );
  XOR U26127 ( .A(n26354), .B(n26355), .Z(n26348) );
  AND U26128 ( .A(n241), .B(n26347), .Z(n26355) );
  XNOR U26129 ( .A(n26345), .B(n26354), .Z(n26347) );
  XNOR U26130 ( .A(n26356), .B(n26357), .Z(n26345) );
  AND U26131 ( .A(n245), .B(n26358), .Z(n26357) );
  XOR U26132 ( .A(p_input[202]), .B(n26356), .Z(n26358) );
  XNOR U26133 ( .A(n26359), .B(n26360), .Z(n26356) );
  AND U26134 ( .A(n249), .B(n26361), .Z(n26360) );
  XOR U26135 ( .A(n26362), .B(n26363), .Z(n26354) );
  AND U26136 ( .A(n253), .B(n26353), .Z(n26363) );
  XNOR U26137 ( .A(n26364), .B(n26351), .Z(n26353) );
  XOR U26138 ( .A(n26365), .B(n26366), .Z(n26351) );
  AND U26139 ( .A(n276), .B(n26367), .Z(n26366) );
  IV U26140 ( .A(n26362), .Z(n26364) );
  XOR U26141 ( .A(n26368), .B(n26369), .Z(n26362) );
  AND U26142 ( .A(n260), .B(n26361), .Z(n26369) );
  XNOR U26143 ( .A(n26359), .B(n26368), .Z(n26361) );
  XNOR U26144 ( .A(n26370), .B(n26371), .Z(n26359) );
  AND U26145 ( .A(n264), .B(n26372), .Z(n26371) );
  XOR U26146 ( .A(p_input[234]), .B(n26370), .Z(n26372) );
  XNOR U26147 ( .A(n26373), .B(n26374), .Z(n26370) );
  AND U26148 ( .A(n268), .B(n26375), .Z(n26374) );
  XOR U26149 ( .A(n26376), .B(n26377), .Z(n26368) );
  AND U26150 ( .A(n272), .B(n26367), .Z(n26377) );
  XNOR U26151 ( .A(n26378), .B(n26365), .Z(n26367) );
  XOR U26152 ( .A(n26379), .B(n26380), .Z(n26365) );
  AND U26153 ( .A(n295), .B(n26381), .Z(n26380) );
  IV U26154 ( .A(n26376), .Z(n26378) );
  XOR U26155 ( .A(n26382), .B(n26383), .Z(n26376) );
  AND U26156 ( .A(n279), .B(n26375), .Z(n26383) );
  XNOR U26157 ( .A(n26373), .B(n26382), .Z(n26375) );
  XNOR U26158 ( .A(n26384), .B(n26385), .Z(n26373) );
  AND U26159 ( .A(n283), .B(n26386), .Z(n26385) );
  XOR U26160 ( .A(p_input[266]), .B(n26384), .Z(n26386) );
  XNOR U26161 ( .A(n26387), .B(n26388), .Z(n26384) );
  AND U26162 ( .A(n287), .B(n26389), .Z(n26388) );
  XOR U26163 ( .A(n26390), .B(n26391), .Z(n26382) );
  AND U26164 ( .A(n291), .B(n26381), .Z(n26391) );
  XNOR U26165 ( .A(n26392), .B(n26379), .Z(n26381) );
  XOR U26166 ( .A(n26393), .B(n26394), .Z(n26379) );
  AND U26167 ( .A(n314), .B(n26395), .Z(n26394) );
  IV U26168 ( .A(n26390), .Z(n26392) );
  XOR U26169 ( .A(n26396), .B(n26397), .Z(n26390) );
  AND U26170 ( .A(n298), .B(n26389), .Z(n26397) );
  XNOR U26171 ( .A(n26387), .B(n26396), .Z(n26389) );
  XNOR U26172 ( .A(n26398), .B(n26399), .Z(n26387) );
  AND U26173 ( .A(n302), .B(n26400), .Z(n26399) );
  XOR U26174 ( .A(p_input[298]), .B(n26398), .Z(n26400) );
  XNOR U26175 ( .A(n26401), .B(n26402), .Z(n26398) );
  AND U26176 ( .A(n306), .B(n26403), .Z(n26402) );
  XOR U26177 ( .A(n26404), .B(n26405), .Z(n26396) );
  AND U26178 ( .A(n310), .B(n26395), .Z(n26405) );
  XNOR U26179 ( .A(n26406), .B(n26393), .Z(n26395) );
  XOR U26180 ( .A(n26407), .B(n26408), .Z(n26393) );
  AND U26181 ( .A(n333), .B(n26409), .Z(n26408) );
  IV U26182 ( .A(n26404), .Z(n26406) );
  XOR U26183 ( .A(n26410), .B(n26411), .Z(n26404) );
  AND U26184 ( .A(n317), .B(n26403), .Z(n26411) );
  XNOR U26185 ( .A(n26401), .B(n26410), .Z(n26403) );
  XNOR U26186 ( .A(n26412), .B(n26413), .Z(n26401) );
  AND U26187 ( .A(n321), .B(n26414), .Z(n26413) );
  XOR U26188 ( .A(p_input[330]), .B(n26412), .Z(n26414) );
  XNOR U26189 ( .A(n26415), .B(n26416), .Z(n26412) );
  AND U26190 ( .A(n325), .B(n26417), .Z(n26416) );
  XOR U26191 ( .A(n26418), .B(n26419), .Z(n26410) );
  AND U26192 ( .A(n329), .B(n26409), .Z(n26419) );
  XNOR U26193 ( .A(n26420), .B(n26407), .Z(n26409) );
  XOR U26194 ( .A(n26421), .B(n26422), .Z(n26407) );
  AND U26195 ( .A(n352), .B(n26423), .Z(n26422) );
  IV U26196 ( .A(n26418), .Z(n26420) );
  XOR U26197 ( .A(n26424), .B(n26425), .Z(n26418) );
  AND U26198 ( .A(n336), .B(n26417), .Z(n26425) );
  XNOR U26199 ( .A(n26415), .B(n26424), .Z(n26417) );
  XNOR U26200 ( .A(n26426), .B(n26427), .Z(n26415) );
  AND U26201 ( .A(n340), .B(n26428), .Z(n26427) );
  XOR U26202 ( .A(p_input[362]), .B(n26426), .Z(n26428) );
  XNOR U26203 ( .A(n26429), .B(n26430), .Z(n26426) );
  AND U26204 ( .A(n344), .B(n26431), .Z(n26430) );
  XOR U26205 ( .A(n26432), .B(n26433), .Z(n26424) );
  AND U26206 ( .A(n348), .B(n26423), .Z(n26433) );
  XNOR U26207 ( .A(n26434), .B(n26421), .Z(n26423) );
  XOR U26208 ( .A(n26435), .B(n26436), .Z(n26421) );
  AND U26209 ( .A(n371), .B(n26437), .Z(n26436) );
  IV U26210 ( .A(n26432), .Z(n26434) );
  XOR U26211 ( .A(n26438), .B(n26439), .Z(n26432) );
  AND U26212 ( .A(n355), .B(n26431), .Z(n26439) );
  XNOR U26213 ( .A(n26429), .B(n26438), .Z(n26431) );
  XNOR U26214 ( .A(n26440), .B(n26441), .Z(n26429) );
  AND U26215 ( .A(n359), .B(n26442), .Z(n26441) );
  XOR U26216 ( .A(p_input[394]), .B(n26440), .Z(n26442) );
  XNOR U26217 ( .A(n26443), .B(n26444), .Z(n26440) );
  AND U26218 ( .A(n363), .B(n26445), .Z(n26444) );
  XOR U26219 ( .A(n26446), .B(n26447), .Z(n26438) );
  AND U26220 ( .A(n367), .B(n26437), .Z(n26447) );
  XNOR U26221 ( .A(n26448), .B(n26435), .Z(n26437) );
  XOR U26222 ( .A(n26449), .B(n26450), .Z(n26435) );
  AND U26223 ( .A(n390), .B(n26451), .Z(n26450) );
  IV U26224 ( .A(n26446), .Z(n26448) );
  XOR U26225 ( .A(n26452), .B(n26453), .Z(n26446) );
  AND U26226 ( .A(n374), .B(n26445), .Z(n26453) );
  XNOR U26227 ( .A(n26443), .B(n26452), .Z(n26445) );
  XNOR U26228 ( .A(n26454), .B(n26455), .Z(n26443) );
  AND U26229 ( .A(n378), .B(n26456), .Z(n26455) );
  XOR U26230 ( .A(p_input[426]), .B(n26454), .Z(n26456) );
  XNOR U26231 ( .A(n26457), .B(n26458), .Z(n26454) );
  AND U26232 ( .A(n382), .B(n26459), .Z(n26458) );
  XOR U26233 ( .A(n26460), .B(n26461), .Z(n26452) );
  AND U26234 ( .A(n386), .B(n26451), .Z(n26461) );
  XNOR U26235 ( .A(n26462), .B(n26449), .Z(n26451) );
  XOR U26236 ( .A(n26463), .B(n26464), .Z(n26449) );
  AND U26237 ( .A(n409), .B(n26465), .Z(n26464) );
  IV U26238 ( .A(n26460), .Z(n26462) );
  XOR U26239 ( .A(n26466), .B(n26467), .Z(n26460) );
  AND U26240 ( .A(n393), .B(n26459), .Z(n26467) );
  XNOR U26241 ( .A(n26457), .B(n26466), .Z(n26459) );
  XNOR U26242 ( .A(n26468), .B(n26469), .Z(n26457) );
  AND U26243 ( .A(n397), .B(n26470), .Z(n26469) );
  XOR U26244 ( .A(p_input[458]), .B(n26468), .Z(n26470) );
  XNOR U26245 ( .A(n26471), .B(n26472), .Z(n26468) );
  AND U26246 ( .A(n401), .B(n26473), .Z(n26472) );
  XOR U26247 ( .A(n26474), .B(n26475), .Z(n26466) );
  AND U26248 ( .A(n405), .B(n26465), .Z(n26475) );
  XNOR U26249 ( .A(n26476), .B(n26463), .Z(n26465) );
  XOR U26250 ( .A(n26477), .B(n26478), .Z(n26463) );
  AND U26251 ( .A(n428), .B(n26479), .Z(n26478) );
  IV U26252 ( .A(n26474), .Z(n26476) );
  XOR U26253 ( .A(n26480), .B(n26481), .Z(n26474) );
  AND U26254 ( .A(n412), .B(n26473), .Z(n26481) );
  XNOR U26255 ( .A(n26471), .B(n26480), .Z(n26473) );
  XNOR U26256 ( .A(n26482), .B(n26483), .Z(n26471) );
  AND U26257 ( .A(n416), .B(n26484), .Z(n26483) );
  XOR U26258 ( .A(p_input[490]), .B(n26482), .Z(n26484) );
  XNOR U26259 ( .A(n26485), .B(n26486), .Z(n26482) );
  AND U26260 ( .A(n420), .B(n26487), .Z(n26486) );
  XOR U26261 ( .A(n26488), .B(n26489), .Z(n26480) );
  AND U26262 ( .A(n424), .B(n26479), .Z(n26489) );
  XNOR U26263 ( .A(n26490), .B(n26477), .Z(n26479) );
  XOR U26264 ( .A(n26491), .B(n26492), .Z(n26477) );
  AND U26265 ( .A(n447), .B(n26493), .Z(n26492) );
  IV U26266 ( .A(n26488), .Z(n26490) );
  XOR U26267 ( .A(n26494), .B(n26495), .Z(n26488) );
  AND U26268 ( .A(n431), .B(n26487), .Z(n26495) );
  XNOR U26269 ( .A(n26485), .B(n26494), .Z(n26487) );
  XNOR U26270 ( .A(n26496), .B(n26497), .Z(n26485) );
  AND U26271 ( .A(n435), .B(n26498), .Z(n26497) );
  XOR U26272 ( .A(p_input[522]), .B(n26496), .Z(n26498) );
  XNOR U26273 ( .A(n26499), .B(n26500), .Z(n26496) );
  AND U26274 ( .A(n439), .B(n26501), .Z(n26500) );
  XOR U26275 ( .A(n26502), .B(n26503), .Z(n26494) );
  AND U26276 ( .A(n443), .B(n26493), .Z(n26503) );
  XNOR U26277 ( .A(n26504), .B(n26491), .Z(n26493) );
  XOR U26278 ( .A(n26505), .B(n26506), .Z(n26491) );
  AND U26279 ( .A(n466), .B(n26507), .Z(n26506) );
  IV U26280 ( .A(n26502), .Z(n26504) );
  XOR U26281 ( .A(n26508), .B(n26509), .Z(n26502) );
  AND U26282 ( .A(n450), .B(n26501), .Z(n26509) );
  XNOR U26283 ( .A(n26499), .B(n26508), .Z(n26501) );
  XNOR U26284 ( .A(n26510), .B(n26511), .Z(n26499) );
  AND U26285 ( .A(n454), .B(n26512), .Z(n26511) );
  XOR U26286 ( .A(p_input[554]), .B(n26510), .Z(n26512) );
  XNOR U26287 ( .A(n26513), .B(n26514), .Z(n26510) );
  AND U26288 ( .A(n458), .B(n26515), .Z(n26514) );
  XOR U26289 ( .A(n26516), .B(n26517), .Z(n26508) );
  AND U26290 ( .A(n462), .B(n26507), .Z(n26517) );
  XNOR U26291 ( .A(n26518), .B(n26505), .Z(n26507) );
  XOR U26292 ( .A(n26519), .B(n26520), .Z(n26505) );
  AND U26293 ( .A(n485), .B(n26521), .Z(n26520) );
  IV U26294 ( .A(n26516), .Z(n26518) );
  XOR U26295 ( .A(n26522), .B(n26523), .Z(n26516) );
  AND U26296 ( .A(n469), .B(n26515), .Z(n26523) );
  XNOR U26297 ( .A(n26513), .B(n26522), .Z(n26515) );
  XNOR U26298 ( .A(n26524), .B(n26525), .Z(n26513) );
  AND U26299 ( .A(n473), .B(n26526), .Z(n26525) );
  XOR U26300 ( .A(p_input[586]), .B(n26524), .Z(n26526) );
  XNOR U26301 ( .A(n26527), .B(n26528), .Z(n26524) );
  AND U26302 ( .A(n477), .B(n26529), .Z(n26528) );
  XOR U26303 ( .A(n26530), .B(n26531), .Z(n26522) );
  AND U26304 ( .A(n481), .B(n26521), .Z(n26531) );
  XNOR U26305 ( .A(n26532), .B(n26519), .Z(n26521) );
  XOR U26306 ( .A(n26533), .B(n26534), .Z(n26519) );
  AND U26307 ( .A(n504), .B(n26535), .Z(n26534) );
  IV U26308 ( .A(n26530), .Z(n26532) );
  XOR U26309 ( .A(n26536), .B(n26537), .Z(n26530) );
  AND U26310 ( .A(n488), .B(n26529), .Z(n26537) );
  XNOR U26311 ( .A(n26527), .B(n26536), .Z(n26529) );
  XNOR U26312 ( .A(n26538), .B(n26539), .Z(n26527) );
  AND U26313 ( .A(n492), .B(n26540), .Z(n26539) );
  XOR U26314 ( .A(p_input[618]), .B(n26538), .Z(n26540) );
  XNOR U26315 ( .A(n26541), .B(n26542), .Z(n26538) );
  AND U26316 ( .A(n496), .B(n26543), .Z(n26542) );
  XOR U26317 ( .A(n26544), .B(n26545), .Z(n26536) );
  AND U26318 ( .A(n500), .B(n26535), .Z(n26545) );
  XNOR U26319 ( .A(n26546), .B(n26533), .Z(n26535) );
  XOR U26320 ( .A(n26547), .B(n26548), .Z(n26533) );
  AND U26321 ( .A(n523), .B(n26549), .Z(n26548) );
  IV U26322 ( .A(n26544), .Z(n26546) );
  XOR U26323 ( .A(n26550), .B(n26551), .Z(n26544) );
  AND U26324 ( .A(n507), .B(n26543), .Z(n26551) );
  XNOR U26325 ( .A(n26541), .B(n26550), .Z(n26543) );
  XNOR U26326 ( .A(n26552), .B(n26553), .Z(n26541) );
  AND U26327 ( .A(n511), .B(n26554), .Z(n26553) );
  XOR U26328 ( .A(p_input[650]), .B(n26552), .Z(n26554) );
  XNOR U26329 ( .A(n26555), .B(n26556), .Z(n26552) );
  AND U26330 ( .A(n515), .B(n26557), .Z(n26556) );
  XOR U26331 ( .A(n26558), .B(n26559), .Z(n26550) );
  AND U26332 ( .A(n519), .B(n26549), .Z(n26559) );
  XNOR U26333 ( .A(n26560), .B(n26547), .Z(n26549) );
  XOR U26334 ( .A(n26561), .B(n26562), .Z(n26547) );
  AND U26335 ( .A(n542), .B(n26563), .Z(n26562) );
  IV U26336 ( .A(n26558), .Z(n26560) );
  XOR U26337 ( .A(n26564), .B(n26565), .Z(n26558) );
  AND U26338 ( .A(n526), .B(n26557), .Z(n26565) );
  XNOR U26339 ( .A(n26555), .B(n26564), .Z(n26557) );
  XNOR U26340 ( .A(n26566), .B(n26567), .Z(n26555) );
  AND U26341 ( .A(n530), .B(n26568), .Z(n26567) );
  XOR U26342 ( .A(p_input[682]), .B(n26566), .Z(n26568) );
  XNOR U26343 ( .A(n26569), .B(n26570), .Z(n26566) );
  AND U26344 ( .A(n534), .B(n26571), .Z(n26570) );
  XOR U26345 ( .A(n26572), .B(n26573), .Z(n26564) );
  AND U26346 ( .A(n538), .B(n26563), .Z(n26573) );
  XNOR U26347 ( .A(n26574), .B(n26561), .Z(n26563) );
  XOR U26348 ( .A(n26575), .B(n26576), .Z(n26561) );
  AND U26349 ( .A(n561), .B(n26577), .Z(n26576) );
  IV U26350 ( .A(n26572), .Z(n26574) );
  XOR U26351 ( .A(n26578), .B(n26579), .Z(n26572) );
  AND U26352 ( .A(n545), .B(n26571), .Z(n26579) );
  XNOR U26353 ( .A(n26569), .B(n26578), .Z(n26571) );
  XNOR U26354 ( .A(n26580), .B(n26581), .Z(n26569) );
  AND U26355 ( .A(n549), .B(n26582), .Z(n26581) );
  XOR U26356 ( .A(p_input[714]), .B(n26580), .Z(n26582) );
  XNOR U26357 ( .A(n26583), .B(n26584), .Z(n26580) );
  AND U26358 ( .A(n553), .B(n26585), .Z(n26584) );
  XOR U26359 ( .A(n26586), .B(n26587), .Z(n26578) );
  AND U26360 ( .A(n557), .B(n26577), .Z(n26587) );
  XNOR U26361 ( .A(n26588), .B(n26575), .Z(n26577) );
  XOR U26362 ( .A(n26589), .B(n26590), .Z(n26575) );
  AND U26363 ( .A(n580), .B(n26591), .Z(n26590) );
  IV U26364 ( .A(n26586), .Z(n26588) );
  XOR U26365 ( .A(n26592), .B(n26593), .Z(n26586) );
  AND U26366 ( .A(n564), .B(n26585), .Z(n26593) );
  XNOR U26367 ( .A(n26583), .B(n26592), .Z(n26585) );
  XNOR U26368 ( .A(n26594), .B(n26595), .Z(n26583) );
  AND U26369 ( .A(n568), .B(n26596), .Z(n26595) );
  XOR U26370 ( .A(p_input[746]), .B(n26594), .Z(n26596) );
  XNOR U26371 ( .A(n26597), .B(n26598), .Z(n26594) );
  AND U26372 ( .A(n572), .B(n26599), .Z(n26598) );
  XOR U26373 ( .A(n26600), .B(n26601), .Z(n26592) );
  AND U26374 ( .A(n576), .B(n26591), .Z(n26601) );
  XNOR U26375 ( .A(n26602), .B(n26589), .Z(n26591) );
  XOR U26376 ( .A(n26603), .B(n26604), .Z(n26589) );
  AND U26377 ( .A(n599), .B(n26605), .Z(n26604) );
  IV U26378 ( .A(n26600), .Z(n26602) );
  XOR U26379 ( .A(n26606), .B(n26607), .Z(n26600) );
  AND U26380 ( .A(n583), .B(n26599), .Z(n26607) );
  XNOR U26381 ( .A(n26597), .B(n26606), .Z(n26599) );
  XNOR U26382 ( .A(n26608), .B(n26609), .Z(n26597) );
  AND U26383 ( .A(n587), .B(n26610), .Z(n26609) );
  XOR U26384 ( .A(p_input[778]), .B(n26608), .Z(n26610) );
  XNOR U26385 ( .A(n26611), .B(n26612), .Z(n26608) );
  AND U26386 ( .A(n591), .B(n26613), .Z(n26612) );
  XOR U26387 ( .A(n26614), .B(n26615), .Z(n26606) );
  AND U26388 ( .A(n595), .B(n26605), .Z(n26615) );
  XNOR U26389 ( .A(n26616), .B(n26603), .Z(n26605) );
  XOR U26390 ( .A(n26617), .B(n26618), .Z(n26603) );
  AND U26391 ( .A(n618), .B(n26619), .Z(n26618) );
  IV U26392 ( .A(n26614), .Z(n26616) );
  XOR U26393 ( .A(n26620), .B(n26621), .Z(n26614) );
  AND U26394 ( .A(n602), .B(n26613), .Z(n26621) );
  XNOR U26395 ( .A(n26611), .B(n26620), .Z(n26613) );
  XNOR U26396 ( .A(n26622), .B(n26623), .Z(n26611) );
  AND U26397 ( .A(n606), .B(n26624), .Z(n26623) );
  XOR U26398 ( .A(p_input[810]), .B(n26622), .Z(n26624) );
  XNOR U26399 ( .A(n26625), .B(n26626), .Z(n26622) );
  AND U26400 ( .A(n610), .B(n26627), .Z(n26626) );
  XOR U26401 ( .A(n26628), .B(n26629), .Z(n26620) );
  AND U26402 ( .A(n614), .B(n26619), .Z(n26629) );
  XNOR U26403 ( .A(n26630), .B(n26617), .Z(n26619) );
  XOR U26404 ( .A(n26631), .B(n26632), .Z(n26617) );
  AND U26405 ( .A(n637), .B(n26633), .Z(n26632) );
  IV U26406 ( .A(n26628), .Z(n26630) );
  XOR U26407 ( .A(n26634), .B(n26635), .Z(n26628) );
  AND U26408 ( .A(n621), .B(n26627), .Z(n26635) );
  XNOR U26409 ( .A(n26625), .B(n26634), .Z(n26627) );
  XNOR U26410 ( .A(n26636), .B(n26637), .Z(n26625) );
  AND U26411 ( .A(n625), .B(n26638), .Z(n26637) );
  XOR U26412 ( .A(p_input[842]), .B(n26636), .Z(n26638) );
  XNOR U26413 ( .A(n26639), .B(n26640), .Z(n26636) );
  AND U26414 ( .A(n629), .B(n26641), .Z(n26640) );
  XOR U26415 ( .A(n26642), .B(n26643), .Z(n26634) );
  AND U26416 ( .A(n633), .B(n26633), .Z(n26643) );
  XNOR U26417 ( .A(n26644), .B(n26631), .Z(n26633) );
  XOR U26418 ( .A(n26645), .B(n26646), .Z(n26631) );
  AND U26419 ( .A(n656), .B(n26647), .Z(n26646) );
  IV U26420 ( .A(n26642), .Z(n26644) );
  XOR U26421 ( .A(n26648), .B(n26649), .Z(n26642) );
  AND U26422 ( .A(n640), .B(n26641), .Z(n26649) );
  XNOR U26423 ( .A(n26639), .B(n26648), .Z(n26641) );
  XNOR U26424 ( .A(n26650), .B(n26651), .Z(n26639) );
  AND U26425 ( .A(n644), .B(n26652), .Z(n26651) );
  XOR U26426 ( .A(p_input[874]), .B(n26650), .Z(n26652) );
  XNOR U26427 ( .A(n26653), .B(n26654), .Z(n26650) );
  AND U26428 ( .A(n648), .B(n26655), .Z(n26654) );
  XOR U26429 ( .A(n26656), .B(n26657), .Z(n26648) );
  AND U26430 ( .A(n652), .B(n26647), .Z(n26657) );
  XNOR U26431 ( .A(n26658), .B(n26645), .Z(n26647) );
  XOR U26432 ( .A(n26659), .B(n26660), .Z(n26645) );
  AND U26433 ( .A(n675), .B(n26661), .Z(n26660) );
  IV U26434 ( .A(n26656), .Z(n26658) );
  XOR U26435 ( .A(n26662), .B(n26663), .Z(n26656) );
  AND U26436 ( .A(n659), .B(n26655), .Z(n26663) );
  XNOR U26437 ( .A(n26653), .B(n26662), .Z(n26655) );
  XNOR U26438 ( .A(n26664), .B(n26665), .Z(n26653) );
  AND U26439 ( .A(n663), .B(n26666), .Z(n26665) );
  XOR U26440 ( .A(p_input[906]), .B(n26664), .Z(n26666) );
  XNOR U26441 ( .A(n26667), .B(n26668), .Z(n26664) );
  AND U26442 ( .A(n667), .B(n26669), .Z(n26668) );
  XOR U26443 ( .A(n26670), .B(n26671), .Z(n26662) );
  AND U26444 ( .A(n671), .B(n26661), .Z(n26671) );
  XNOR U26445 ( .A(n26672), .B(n26659), .Z(n26661) );
  XOR U26446 ( .A(n26673), .B(n26674), .Z(n26659) );
  AND U26447 ( .A(n694), .B(n26675), .Z(n26674) );
  IV U26448 ( .A(n26670), .Z(n26672) );
  XOR U26449 ( .A(n26676), .B(n26677), .Z(n26670) );
  AND U26450 ( .A(n678), .B(n26669), .Z(n26677) );
  XNOR U26451 ( .A(n26667), .B(n26676), .Z(n26669) );
  XNOR U26452 ( .A(n26678), .B(n26679), .Z(n26667) );
  AND U26453 ( .A(n682), .B(n26680), .Z(n26679) );
  XOR U26454 ( .A(p_input[938]), .B(n26678), .Z(n26680) );
  XNOR U26455 ( .A(n26681), .B(n26682), .Z(n26678) );
  AND U26456 ( .A(n686), .B(n26683), .Z(n26682) );
  XOR U26457 ( .A(n26684), .B(n26685), .Z(n26676) );
  AND U26458 ( .A(n690), .B(n26675), .Z(n26685) );
  XNOR U26459 ( .A(n26686), .B(n26673), .Z(n26675) );
  XOR U26460 ( .A(n26687), .B(n26688), .Z(n26673) );
  AND U26461 ( .A(n713), .B(n26689), .Z(n26688) );
  IV U26462 ( .A(n26684), .Z(n26686) );
  XOR U26463 ( .A(n26690), .B(n26691), .Z(n26684) );
  AND U26464 ( .A(n697), .B(n26683), .Z(n26691) );
  XNOR U26465 ( .A(n26681), .B(n26690), .Z(n26683) );
  XNOR U26466 ( .A(n26692), .B(n26693), .Z(n26681) );
  AND U26467 ( .A(n701), .B(n26694), .Z(n26693) );
  XOR U26468 ( .A(p_input[970]), .B(n26692), .Z(n26694) );
  XNOR U26469 ( .A(n26695), .B(n26696), .Z(n26692) );
  AND U26470 ( .A(n705), .B(n26697), .Z(n26696) );
  XOR U26471 ( .A(n26698), .B(n26699), .Z(n26690) );
  AND U26472 ( .A(n709), .B(n26689), .Z(n26699) );
  XNOR U26473 ( .A(n26700), .B(n26687), .Z(n26689) );
  XOR U26474 ( .A(n26701), .B(n26702), .Z(n26687) );
  AND U26475 ( .A(n732), .B(n26703), .Z(n26702) );
  IV U26476 ( .A(n26698), .Z(n26700) );
  XOR U26477 ( .A(n26704), .B(n26705), .Z(n26698) );
  AND U26478 ( .A(n716), .B(n26697), .Z(n26705) );
  XNOR U26479 ( .A(n26695), .B(n26704), .Z(n26697) );
  XNOR U26480 ( .A(n26706), .B(n26707), .Z(n26695) );
  AND U26481 ( .A(n720), .B(n26708), .Z(n26707) );
  XOR U26482 ( .A(p_input[1002]), .B(n26706), .Z(n26708) );
  XNOR U26483 ( .A(n26709), .B(n26710), .Z(n26706) );
  AND U26484 ( .A(n724), .B(n26711), .Z(n26710) );
  XOR U26485 ( .A(n26712), .B(n26713), .Z(n26704) );
  AND U26486 ( .A(n728), .B(n26703), .Z(n26713) );
  XNOR U26487 ( .A(n26714), .B(n26701), .Z(n26703) );
  XOR U26488 ( .A(n26715), .B(n26716), .Z(n26701) );
  AND U26489 ( .A(n751), .B(n26717), .Z(n26716) );
  IV U26490 ( .A(n26712), .Z(n26714) );
  XOR U26491 ( .A(n26718), .B(n26719), .Z(n26712) );
  AND U26492 ( .A(n735), .B(n26711), .Z(n26719) );
  XNOR U26493 ( .A(n26709), .B(n26718), .Z(n26711) );
  XNOR U26494 ( .A(n26720), .B(n26721), .Z(n26709) );
  AND U26495 ( .A(n739), .B(n26722), .Z(n26721) );
  XOR U26496 ( .A(p_input[1034]), .B(n26720), .Z(n26722) );
  XNOR U26497 ( .A(n26723), .B(n26724), .Z(n26720) );
  AND U26498 ( .A(n743), .B(n26725), .Z(n26724) );
  XOR U26499 ( .A(n26726), .B(n26727), .Z(n26718) );
  AND U26500 ( .A(n747), .B(n26717), .Z(n26727) );
  XNOR U26501 ( .A(n26728), .B(n26715), .Z(n26717) );
  XOR U26502 ( .A(n26729), .B(n26730), .Z(n26715) );
  AND U26503 ( .A(n770), .B(n26731), .Z(n26730) );
  IV U26504 ( .A(n26726), .Z(n26728) );
  XOR U26505 ( .A(n26732), .B(n26733), .Z(n26726) );
  AND U26506 ( .A(n754), .B(n26725), .Z(n26733) );
  XNOR U26507 ( .A(n26723), .B(n26732), .Z(n26725) );
  XNOR U26508 ( .A(n26734), .B(n26735), .Z(n26723) );
  AND U26509 ( .A(n758), .B(n26736), .Z(n26735) );
  XOR U26510 ( .A(p_input[1066]), .B(n26734), .Z(n26736) );
  XNOR U26511 ( .A(n26737), .B(n26738), .Z(n26734) );
  AND U26512 ( .A(n762), .B(n26739), .Z(n26738) );
  XOR U26513 ( .A(n26740), .B(n26741), .Z(n26732) );
  AND U26514 ( .A(n766), .B(n26731), .Z(n26741) );
  XNOR U26515 ( .A(n26742), .B(n26729), .Z(n26731) );
  XOR U26516 ( .A(n26743), .B(n26744), .Z(n26729) );
  AND U26517 ( .A(n789), .B(n26745), .Z(n26744) );
  IV U26518 ( .A(n26740), .Z(n26742) );
  XOR U26519 ( .A(n26746), .B(n26747), .Z(n26740) );
  AND U26520 ( .A(n773), .B(n26739), .Z(n26747) );
  XNOR U26521 ( .A(n26737), .B(n26746), .Z(n26739) );
  XNOR U26522 ( .A(n26748), .B(n26749), .Z(n26737) );
  AND U26523 ( .A(n777), .B(n26750), .Z(n26749) );
  XOR U26524 ( .A(p_input[1098]), .B(n26748), .Z(n26750) );
  XNOR U26525 ( .A(n26751), .B(n26752), .Z(n26748) );
  AND U26526 ( .A(n781), .B(n26753), .Z(n26752) );
  XOR U26527 ( .A(n26754), .B(n26755), .Z(n26746) );
  AND U26528 ( .A(n785), .B(n26745), .Z(n26755) );
  XNOR U26529 ( .A(n26756), .B(n26743), .Z(n26745) );
  XOR U26530 ( .A(n26757), .B(n26758), .Z(n26743) );
  AND U26531 ( .A(n808), .B(n26759), .Z(n26758) );
  IV U26532 ( .A(n26754), .Z(n26756) );
  XOR U26533 ( .A(n26760), .B(n26761), .Z(n26754) );
  AND U26534 ( .A(n792), .B(n26753), .Z(n26761) );
  XNOR U26535 ( .A(n26751), .B(n26760), .Z(n26753) );
  XNOR U26536 ( .A(n26762), .B(n26763), .Z(n26751) );
  AND U26537 ( .A(n796), .B(n26764), .Z(n26763) );
  XOR U26538 ( .A(p_input[1130]), .B(n26762), .Z(n26764) );
  XNOR U26539 ( .A(n26765), .B(n26766), .Z(n26762) );
  AND U26540 ( .A(n800), .B(n26767), .Z(n26766) );
  XOR U26541 ( .A(n26768), .B(n26769), .Z(n26760) );
  AND U26542 ( .A(n804), .B(n26759), .Z(n26769) );
  XNOR U26543 ( .A(n26770), .B(n26757), .Z(n26759) );
  XOR U26544 ( .A(n26771), .B(n26772), .Z(n26757) );
  AND U26545 ( .A(n827), .B(n26773), .Z(n26772) );
  IV U26546 ( .A(n26768), .Z(n26770) );
  XOR U26547 ( .A(n26774), .B(n26775), .Z(n26768) );
  AND U26548 ( .A(n811), .B(n26767), .Z(n26775) );
  XNOR U26549 ( .A(n26765), .B(n26774), .Z(n26767) );
  XNOR U26550 ( .A(n26776), .B(n26777), .Z(n26765) );
  AND U26551 ( .A(n815), .B(n26778), .Z(n26777) );
  XOR U26552 ( .A(p_input[1162]), .B(n26776), .Z(n26778) );
  XNOR U26553 ( .A(n26779), .B(n26780), .Z(n26776) );
  AND U26554 ( .A(n819), .B(n26781), .Z(n26780) );
  XOR U26555 ( .A(n26782), .B(n26783), .Z(n26774) );
  AND U26556 ( .A(n823), .B(n26773), .Z(n26783) );
  XNOR U26557 ( .A(n26784), .B(n26771), .Z(n26773) );
  XOR U26558 ( .A(n26785), .B(n26786), .Z(n26771) );
  AND U26559 ( .A(n846), .B(n26787), .Z(n26786) );
  IV U26560 ( .A(n26782), .Z(n26784) );
  XOR U26561 ( .A(n26788), .B(n26789), .Z(n26782) );
  AND U26562 ( .A(n830), .B(n26781), .Z(n26789) );
  XNOR U26563 ( .A(n26779), .B(n26788), .Z(n26781) );
  XNOR U26564 ( .A(n26790), .B(n26791), .Z(n26779) );
  AND U26565 ( .A(n834), .B(n26792), .Z(n26791) );
  XOR U26566 ( .A(p_input[1194]), .B(n26790), .Z(n26792) );
  XNOR U26567 ( .A(n26793), .B(n26794), .Z(n26790) );
  AND U26568 ( .A(n838), .B(n26795), .Z(n26794) );
  XOR U26569 ( .A(n26796), .B(n26797), .Z(n26788) );
  AND U26570 ( .A(n842), .B(n26787), .Z(n26797) );
  XNOR U26571 ( .A(n26798), .B(n26785), .Z(n26787) );
  XOR U26572 ( .A(n26799), .B(n26800), .Z(n26785) );
  AND U26573 ( .A(n865), .B(n26801), .Z(n26800) );
  IV U26574 ( .A(n26796), .Z(n26798) );
  XOR U26575 ( .A(n26802), .B(n26803), .Z(n26796) );
  AND U26576 ( .A(n849), .B(n26795), .Z(n26803) );
  XNOR U26577 ( .A(n26793), .B(n26802), .Z(n26795) );
  XNOR U26578 ( .A(n26804), .B(n26805), .Z(n26793) );
  AND U26579 ( .A(n853), .B(n26806), .Z(n26805) );
  XOR U26580 ( .A(p_input[1226]), .B(n26804), .Z(n26806) );
  XNOR U26581 ( .A(n26807), .B(n26808), .Z(n26804) );
  AND U26582 ( .A(n857), .B(n26809), .Z(n26808) );
  XOR U26583 ( .A(n26810), .B(n26811), .Z(n26802) );
  AND U26584 ( .A(n861), .B(n26801), .Z(n26811) );
  XNOR U26585 ( .A(n26812), .B(n26799), .Z(n26801) );
  XOR U26586 ( .A(n26813), .B(n26814), .Z(n26799) );
  AND U26587 ( .A(n884), .B(n26815), .Z(n26814) );
  IV U26588 ( .A(n26810), .Z(n26812) );
  XOR U26589 ( .A(n26816), .B(n26817), .Z(n26810) );
  AND U26590 ( .A(n868), .B(n26809), .Z(n26817) );
  XNOR U26591 ( .A(n26807), .B(n26816), .Z(n26809) );
  XNOR U26592 ( .A(n26818), .B(n26819), .Z(n26807) );
  AND U26593 ( .A(n872), .B(n26820), .Z(n26819) );
  XOR U26594 ( .A(p_input[1258]), .B(n26818), .Z(n26820) );
  XNOR U26595 ( .A(n26821), .B(n26822), .Z(n26818) );
  AND U26596 ( .A(n876), .B(n26823), .Z(n26822) );
  XOR U26597 ( .A(n26824), .B(n26825), .Z(n26816) );
  AND U26598 ( .A(n880), .B(n26815), .Z(n26825) );
  XNOR U26599 ( .A(n26826), .B(n26813), .Z(n26815) );
  XOR U26600 ( .A(n26827), .B(n26828), .Z(n26813) );
  AND U26601 ( .A(n903), .B(n26829), .Z(n26828) );
  IV U26602 ( .A(n26824), .Z(n26826) );
  XOR U26603 ( .A(n26830), .B(n26831), .Z(n26824) );
  AND U26604 ( .A(n887), .B(n26823), .Z(n26831) );
  XNOR U26605 ( .A(n26821), .B(n26830), .Z(n26823) );
  XNOR U26606 ( .A(n26832), .B(n26833), .Z(n26821) );
  AND U26607 ( .A(n891), .B(n26834), .Z(n26833) );
  XOR U26608 ( .A(p_input[1290]), .B(n26832), .Z(n26834) );
  XNOR U26609 ( .A(n26835), .B(n26836), .Z(n26832) );
  AND U26610 ( .A(n895), .B(n26837), .Z(n26836) );
  XOR U26611 ( .A(n26838), .B(n26839), .Z(n26830) );
  AND U26612 ( .A(n899), .B(n26829), .Z(n26839) );
  XNOR U26613 ( .A(n26840), .B(n26827), .Z(n26829) );
  XOR U26614 ( .A(n26841), .B(n26842), .Z(n26827) );
  AND U26615 ( .A(n922), .B(n26843), .Z(n26842) );
  IV U26616 ( .A(n26838), .Z(n26840) );
  XOR U26617 ( .A(n26844), .B(n26845), .Z(n26838) );
  AND U26618 ( .A(n906), .B(n26837), .Z(n26845) );
  XNOR U26619 ( .A(n26835), .B(n26844), .Z(n26837) );
  XNOR U26620 ( .A(n26846), .B(n26847), .Z(n26835) );
  AND U26621 ( .A(n910), .B(n26848), .Z(n26847) );
  XOR U26622 ( .A(p_input[1322]), .B(n26846), .Z(n26848) );
  XNOR U26623 ( .A(n26849), .B(n26850), .Z(n26846) );
  AND U26624 ( .A(n914), .B(n26851), .Z(n26850) );
  XOR U26625 ( .A(n26852), .B(n26853), .Z(n26844) );
  AND U26626 ( .A(n918), .B(n26843), .Z(n26853) );
  XNOR U26627 ( .A(n26854), .B(n26841), .Z(n26843) );
  XOR U26628 ( .A(n26855), .B(n26856), .Z(n26841) );
  AND U26629 ( .A(n941), .B(n26857), .Z(n26856) );
  IV U26630 ( .A(n26852), .Z(n26854) );
  XOR U26631 ( .A(n26858), .B(n26859), .Z(n26852) );
  AND U26632 ( .A(n925), .B(n26851), .Z(n26859) );
  XNOR U26633 ( .A(n26849), .B(n26858), .Z(n26851) );
  XNOR U26634 ( .A(n26860), .B(n26861), .Z(n26849) );
  AND U26635 ( .A(n929), .B(n26862), .Z(n26861) );
  XOR U26636 ( .A(p_input[1354]), .B(n26860), .Z(n26862) );
  XNOR U26637 ( .A(n26863), .B(n26864), .Z(n26860) );
  AND U26638 ( .A(n933), .B(n26865), .Z(n26864) );
  XOR U26639 ( .A(n26866), .B(n26867), .Z(n26858) );
  AND U26640 ( .A(n937), .B(n26857), .Z(n26867) );
  XNOR U26641 ( .A(n26868), .B(n26855), .Z(n26857) );
  XOR U26642 ( .A(n26869), .B(n26870), .Z(n26855) );
  AND U26643 ( .A(n960), .B(n26871), .Z(n26870) );
  IV U26644 ( .A(n26866), .Z(n26868) );
  XOR U26645 ( .A(n26872), .B(n26873), .Z(n26866) );
  AND U26646 ( .A(n944), .B(n26865), .Z(n26873) );
  XNOR U26647 ( .A(n26863), .B(n26872), .Z(n26865) );
  XNOR U26648 ( .A(n26874), .B(n26875), .Z(n26863) );
  AND U26649 ( .A(n948), .B(n26876), .Z(n26875) );
  XOR U26650 ( .A(p_input[1386]), .B(n26874), .Z(n26876) );
  XNOR U26651 ( .A(n26877), .B(n26878), .Z(n26874) );
  AND U26652 ( .A(n952), .B(n26879), .Z(n26878) );
  XOR U26653 ( .A(n26880), .B(n26881), .Z(n26872) );
  AND U26654 ( .A(n956), .B(n26871), .Z(n26881) );
  XNOR U26655 ( .A(n26882), .B(n26869), .Z(n26871) );
  XOR U26656 ( .A(n26883), .B(n26884), .Z(n26869) );
  AND U26657 ( .A(n979), .B(n26885), .Z(n26884) );
  IV U26658 ( .A(n26880), .Z(n26882) );
  XOR U26659 ( .A(n26886), .B(n26887), .Z(n26880) );
  AND U26660 ( .A(n963), .B(n26879), .Z(n26887) );
  XNOR U26661 ( .A(n26877), .B(n26886), .Z(n26879) );
  XNOR U26662 ( .A(n26888), .B(n26889), .Z(n26877) );
  AND U26663 ( .A(n967), .B(n26890), .Z(n26889) );
  XOR U26664 ( .A(p_input[1418]), .B(n26888), .Z(n26890) );
  XNOR U26665 ( .A(n26891), .B(n26892), .Z(n26888) );
  AND U26666 ( .A(n971), .B(n26893), .Z(n26892) );
  XOR U26667 ( .A(n26894), .B(n26895), .Z(n26886) );
  AND U26668 ( .A(n975), .B(n26885), .Z(n26895) );
  XNOR U26669 ( .A(n26896), .B(n26883), .Z(n26885) );
  XOR U26670 ( .A(n26897), .B(n26898), .Z(n26883) );
  AND U26671 ( .A(n998), .B(n26899), .Z(n26898) );
  IV U26672 ( .A(n26894), .Z(n26896) );
  XOR U26673 ( .A(n26900), .B(n26901), .Z(n26894) );
  AND U26674 ( .A(n982), .B(n26893), .Z(n26901) );
  XNOR U26675 ( .A(n26891), .B(n26900), .Z(n26893) );
  XNOR U26676 ( .A(n26902), .B(n26903), .Z(n26891) );
  AND U26677 ( .A(n986), .B(n26904), .Z(n26903) );
  XOR U26678 ( .A(p_input[1450]), .B(n26902), .Z(n26904) );
  XNOR U26679 ( .A(n26905), .B(n26906), .Z(n26902) );
  AND U26680 ( .A(n990), .B(n26907), .Z(n26906) );
  XOR U26681 ( .A(n26908), .B(n26909), .Z(n26900) );
  AND U26682 ( .A(n994), .B(n26899), .Z(n26909) );
  XNOR U26683 ( .A(n26910), .B(n26897), .Z(n26899) );
  XOR U26684 ( .A(n26911), .B(n26912), .Z(n26897) );
  AND U26685 ( .A(n1017), .B(n26913), .Z(n26912) );
  IV U26686 ( .A(n26908), .Z(n26910) );
  XOR U26687 ( .A(n26914), .B(n26915), .Z(n26908) );
  AND U26688 ( .A(n1001), .B(n26907), .Z(n26915) );
  XNOR U26689 ( .A(n26905), .B(n26914), .Z(n26907) );
  XNOR U26690 ( .A(n26916), .B(n26917), .Z(n26905) );
  AND U26691 ( .A(n1005), .B(n26918), .Z(n26917) );
  XOR U26692 ( .A(p_input[1482]), .B(n26916), .Z(n26918) );
  XNOR U26693 ( .A(n26919), .B(n26920), .Z(n26916) );
  AND U26694 ( .A(n1009), .B(n26921), .Z(n26920) );
  XOR U26695 ( .A(n26922), .B(n26923), .Z(n26914) );
  AND U26696 ( .A(n1013), .B(n26913), .Z(n26923) );
  XNOR U26697 ( .A(n26924), .B(n26911), .Z(n26913) );
  XOR U26698 ( .A(n26925), .B(n26926), .Z(n26911) );
  AND U26699 ( .A(n1036), .B(n26927), .Z(n26926) );
  IV U26700 ( .A(n26922), .Z(n26924) );
  XOR U26701 ( .A(n26928), .B(n26929), .Z(n26922) );
  AND U26702 ( .A(n1020), .B(n26921), .Z(n26929) );
  XNOR U26703 ( .A(n26919), .B(n26928), .Z(n26921) );
  XNOR U26704 ( .A(n26930), .B(n26931), .Z(n26919) );
  AND U26705 ( .A(n1024), .B(n26932), .Z(n26931) );
  XOR U26706 ( .A(p_input[1514]), .B(n26930), .Z(n26932) );
  XNOR U26707 ( .A(n26933), .B(n26934), .Z(n26930) );
  AND U26708 ( .A(n1028), .B(n26935), .Z(n26934) );
  XOR U26709 ( .A(n26936), .B(n26937), .Z(n26928) );
  AND U26710 ( .A(n1032), .B(n26927), .Z(n26937) );
  XNOR U26711 ( .A(n26938), .B(n26925), .Z(n26927) );
  XOR U26712 ( .A(n26939), .B(n26940), .Z(n26925) );
  AND U26713 ( .A(n1055), .B(n26941), .Z(n26940) );
  IV U26714 ( .A(n26936), .Z(n26938) );
  XOR U26715 ( .A(n26942), .B(n26943), .Z(n26936) );
  AND U26716 ( .A(n1039), .B(n26935), .Z(n26943) );
  XNOR U26717 ( .A(n26933), .B(n26942), .Z(n26935) );
  XNOR U26718 ( .A(n26944), .B(n26945), .Z(n26933) );
  AND U26719 ( .A(n1043), .B(n26946), .Z(n26945) );
  XOR U26720 ( .A(p_input[1546]), .B(n26944), .Z(n26946) );
  XNOR U26721 ( .A(n26947), .B(n26948), .Z(n26944) );
  AND U26722 ( .A(n1047), .B(n26949), .Z(n26948) );
  XOR U26723 ( .A(n26950), .B(n26951), .Z(n26942) );
  AND U26724 ( .A(n1051), .B(n26941), .Z(n26951) );
  XNOR U26725 ( .A(n26952), .B(n26939), .Z(n26941) );
  XOR U26726 ( .A(n26953), .B(n26954), .Z(n26939) );
  AND U26727 ( .A(n1074), .B(n26955), .Z(n26954) );
  IV U26728 ( .A(n26950), .Z(n26952) );
  XOR U26729 ( .A(n26956), .B(n26957), .Z(n26950) );
  AND U26730 ( .A(n1058), .B(n26949), .Z(n26957) );
  XNOR U26731 ( .A(n26947), .B(n26956), .Z(n26949) );
  XNOR U26732 ( .A(n26958), .B(n26959), .Z(n26947) );
  AND U26733 ( .A(n1062), .B(n26960), .Z(n26959) );
  XOR U26734 ( .A(p_input[1578]), .B(n26958), .Z(n26960) );
  XNOR U26735 ( .A(n26961), .B(n26962), .Z(n26958) );
  AND U26736 ( .A(n1066), .B(n26963), .Z(n26962) );
  XOR U26737 ( .A(n26964), .B(n26965), .Z(n26956) );
  AND U26738 ( .A(n1070), .B(n26955), .Z(n26965) );
  XNOR U26739 ( .A(n26966), .B(n26953), .Z(n26955) );
  XOR U26740 ( .A(n26967), .B(n26968), .Z(n26953) );
  AND U26741 ( .A(n1093), .B(n26969), .Z(n26968) );
  IV U26742 ( .A(n26964), .Z(n26966) );
  XOR U26743 ( .A(n26970), .B(n26971), .Z(n26964) );
  AND U26744 ( .A(n1077), .B(n26963), .Z(n26971) );
  XNOR U26745 ( .A(n26961), .B(n26970), .Z(n26963) );
  XNOR U26746 ( .A(n26972), .B(n26973), .Z(n26961) );
  AND U26747 ( .A(n1081), .B(n26974), .Z(n26973) );
  XOR U26748 ( .A(p_input[1610]), .B(n26972), .Z(n26974) );
  XNOR U26749 ( .A(n26975), .B(n26976), .Z(n26972) );
  AND U26750 ( .A(n1085), .B(n26977), .Z(n26976) );
  XOR U26751 ( .A(n26978), .B(n26979), .Z(n26970) );
  AND U26752 ( .A(n1089), .B(n26969), .Z(n26979) );
  XNOR U26753 ( .A(n26980), .B(n26967), .Z(n26969) );
  XOR U26754 ( .A(n26981), .B(n26982), .Z(n26967) );
  AND U26755 ( .A(n1112), .B(n26983), .Z(n26982) );
  IV U26756 ( .A(n26978), .Z(n26980) );
  XOR U26757 ( .A(n26984), .B(n26985), .Z(n26978) );
  AND U26758 ( .A(n1096), .B(n26977), .Z(n26985) );
  XNOR U26759 ( .A(n26975), .B(n26984), .Z(n26977) );
  XNOR U26760 ( .A(n26986), .B(n26987), .Z(n26975) );
  AND U26761 ( .A(n1100), .B(n26988), .Z(n26987) );
  XOR U26762 ( .A(p_input[1642]), .B(n26986), .Z(n26988) );
  XNOR U26763 ( .A(n26989), .B(n26990), .Z(n26986) );
  AND U26764 ( .A(n1104), .B(n26991), .Z(n26990) );
  XOR U26765 ( .A(n26992), .B(n26993), .Z(n26984) );
  AND U26766 ( .A(n1108), .B(n26983), .Z(n26993) );
  XNOR U26767 ( .A(n26994), .B(n26981), .Z(n26983) );
  XOR U26768 ( .A(n26995), .B(n26996), .Z(n26981) );
  AND U26769 ( .A(n1131), .B(n26997), .Z(n26996) );
  IV U26770 ( .A(n26992), .Z(n26994) );
  XOR U26771 ( .A(n26998), .B(n26999), .Z(n26992) );
  AND U26772 ( .A(n1115), .B(n26991), .Z(n26999) );
  XNOR U26773 ( .A(n26989), .B(n26998), .Z(n26991) );
  XNOR U26774 ( .A(n27000), .B(n27001), .Z(n26989) );
  AND U26775 ( .A(n1119), .B(n27002), .Z(n27001) );
  XOR U26776 ( .A(p_input[1674]), .B(n27000), .Z(n27002) );
  XNOR U26777 ( .A(n27003), .B(n27004), .Z(n27000) );
  AND U26778 ( .A(n1123), .B(n27005), .Z(n27004) );
  XOR U26779 ( .A(n27006), .B(n27007), .Z(n26998) );
  AND U26780 ( .A(n1127), .B(n26997), .Z(n27007) );
  XNOR U26781 ( .A(n27008), .B(n26995), .Z(n26997) );
  XOR U26782 ( .A(n27009), .B(n27010), .Z(n26995) );
  AND U26783 ( .A(n1150), .B(n27011), .Z(n27010) );
  IV U26784 ( .A(n27006), .Z(n27008) );
  XOR U26785 ( .A(n27012), .B(n27013), .Z(n27006) );
  AND U26786 ( .A(n1134), .B(n27005), .Z(n27013) );
  XNOR U26787 ( .A(n27003), .B(n27012), .Z(n27005) );
  XNOR U26788 ( .A(n27014), .B(n27015), .Z(n27003) );
  AND U26789 ( .A(n1138), .B(n27016), .Z(n27015) );
  XOR U26790 ( .A(p_input[1706]), .B(n27014), .Z(n27016) );
  XNOR U26791 ( .A(n27017), .B(n27018), .Z(n27014) );
  AND U26792 ( .A(n1142), .B(n27019), .Z(n27018) );
  XOR U26793 ( .A(n27020), .B(n27021), .Z(n27012) );
  AND U26794 ( .A(n1146), .B(n27011), .Z(n27021) );
  XNOR U26795 ( .A(n27022), .B(n27009), .Z(n27011) );
  XOR U26796 ( .A(n27023), .B(n27024), .Z(n27009) );
  AND U26797 ( .A(n1169), .B(n27025), .Z(n27024) );
  IV U26798 ( .A(n27020), .Z(n27022) );
  XOR U26799 ( .A(n27026), .B(n27027), .Z(n27020) );
  AND U26800 ( .A(n1153), .B(n27019), .Z(n27027) );
  XNOR U26801 ( .A(n27017), .B(n27026), .Z(n27019) );
  XNOR U26802 ( .A(n27028), .B(n27029), .Z(n27017) );
  AND U26803 ( .A(n1157), .B(n27030), .Z(n27029) );
  XOR U26804 ( .A(p_input[1738]), .B(n27028), .Z(n27030) );
  XNOR U26805 ( .A(n27031), .B(n27032), .Z(n27028) );
  AND U26806 ( .A(n1161), .B(n27033), .Z(n27032) );
  XOR U26807 ( .A(n27034), .B(n27035), .Z(n27026) );
  AND U26808 ( .A(n1165), .B(n27025), .Z(n27035) );
  XNOR U26809 ( .A(n27036), .B(n27023), .Z(n27025) );
  XOR U26810 ( .A(n27037), .B(n27038), .Z(n27023) );
  AND U26811 ( .A(n1188), .B(n27039), .Z(n27038) );
  IV U26812 ( .A(n27034), .Z(n27036) );
  XOR U26813 ( .A(n27040), .B(n27041), .Z(n27034) );
  AND U26814 ( .A(n1172), .B(n27033), .Z(n27041) );
  XNOR U26815 ( .A(n27031), .B(n27040), .Z(n27033) );
  XNOR U26816 ( .A(n27042), .B(n27043), .Z(n27031) );
  AND U26817 ( .A(n1176), .B(n27044), .Z(n27043) );
  XOR U26818 ( .A(p_input[1770]), .B(n27042), .Z(n27044) );
  XNOR U26819 ( .A(n27045), .B(n27046), .Z(n27042) );
  AND U26820 ( .A(n1180), .B(n27047), .Z(n27046) );
  XOR U26821 ( .A(n27048), .B(n27049), .Z(n27040) );
  AND U26822 ( .A(n1184), .B(n27039), .Z(n27049) );
  XNOR U26823 ( .A(n27050), .B(n27037), .Z(n27039) );
  XOR U26824 ( .A(n27051), .B(n27052), .Z(n27037) );
  AND U26825 ( .A(n1207), .B(n27053), .Z(n27052) );
  IV U26826 ( .A(n27048), .Z(n27050) );
  XOR U26827 ( .A(n27054), .B(n27055), .Z(n27048) );
  AND U26828 ( .A(n1191), .B(n27047), .Z(n27055) );
  XNOR U26829 ( .A(n27045), .B(n27054), .Z(n27047) );
  XNOR U26830 ( .A(n27056), .B(n27057), .Z(n27045) );
  AND U26831 ( .A(n1195), .B(n27058), .Z(n27057) );
  XOR U26832 ( .A(p_input[1802]), .B(n27056), .Z(n27058) );
  XNOR U26833 ( .A(n27059), .B(n27060), .Z(n27056) );
  AND U26834 ( .A(n1199), .B(n27061), .Z(n27060) );
  XOR U26835 ( .A(n27062), .B(n27063), .Z(n27054) );
  AND U26836 ( .A(n1203), .B(n27053), .Z(n27063) );
  XNOR U26837 ( .A(n27064), .B(n27051), .Z(n27053) );
  XOR U26838 ( .A(n27065), .B(n27066), .Z(n27051) );
  AND U26839 ( .A(n1226), .B(n27067), .Z(n27066) );
  IV U26840 ( .A(n27062), .Z(n27064) );
  XOR U26841 ( .A(n27068), .B(n27069), .Z(n27062) );
  AND U26842 ( .A(n1210), .B(n27061), .Z(n27069) );
  XNOR U26843 ( .A(n27059), .B(n27068), .Z(n27061) );
  XNOR U26844 ( .A(n27070), .B(n27071), .Z(n27059) );
  AND U26845 ( .A(n1214), .B(n27072), .Z(n27071) );
  XOR U26846 ( .A(p_input[1834]), .B(n27070), .Z(n27072) );
  XNOR U26847 ( .A(n27073), .B(n27074), .Z(n27070) );
  AND U26848 ( .A(n1218), .B(n27075), .Z(n27074) );
  XOR U26849 ( .A(n27076), .B(n27077), .Z(n27068) );
  AND U26850 ( .A(n1222), .B(n27067), .Z(n27077) );
  XNOR U26851 ( .A(n27078), .B(n27065), .Z(n27067) );
  XOR U26852 ( .A(n27079), .B(n27080), .Z(n27065) );
  AND U26853 ( .A(n1245), .B(n27081), .Z(n27080) );
  IV U26854 ( .A(n27076), .Z(n27078) );
  XOR U26855 ( .A(n27082), .B(n27083), .Z(n27076) );
  AND U26856 ( .A(n1229), .B(n27075), .Z(n27083) );
  XNOR U26857 ( .A(n27073), .B(n27082), .Z(n27075) );
  XNOR U26858 ( .A(n27084), .B(n27085), .Z(n27073) );
  AND U26859 ( .A(n1233), .B(n27086), .Z(n27085) );
  XOR U26860 ( .A(p_input[1866]), .B(n27084), .Z(n27086) );
  XNOR U26861 ( .A(n27087), .B(n27088), .Z(n27084) );
  AND U26862 ( .A(n1237), .B(n27089), .Z(n27088) );
  XOR U26863 ( .A(n27090), .B(n27091), .Z(n27082) );
  AND U26864 ( .A(n1241), .B(n27081), .Z(n27091) );
  XNOR U26865 ( .A(n27092), .B(n27079), .Z(n27081) );
  XOR U26866 ( .A(n27093), .B(n27094), .Z(n27079) );
  AND U26867 ( .A(n1264), .B(n27095), .Z(n27094) );
  IV U26868 ( .A(n27090), .Z(n27092) );
  XOR U26869 ( .A(n27096), .B(n27097), .Z(n27090) );
  AND U26870 ( .A(n1248), .B(n27089), .Z(n27097) );
  XNOR U26871 ( .A(n27087), .B(n27096), .Z(n27089) );
  XNOR U26872 ( .A(n27098), .B(n27099), .Z(n27087) );
  AND U26873 ( .A(n1252), .B(n27100), .Z(n27099) );
  XOR U26874 ( .A(p_input[1898]), .B(n27098), .Z(n27100) );
  XNOR U26875 ( .A(n27101), .B(n27102), .Z(n27098) );
  AND U26876 ( .A(n1256), .B(n27103), .Z(n27102) );
  XOR U26877 ( .A(n27104), .B(n27105), .Z(n27096) );
  AND U26878 ( .A(n1260), .B(n27095), .Z(n27105) );
  XNOR U26879 ( .A(n27106), .B(n27093), .Z(n27095) );
  XOR U26880 ( .A(n27107), .B(n27108), .Z(n27093) );
  AND U26881 ( .A(n1282), .B(n27109), .Z(n27108) );
  IV U26882 ( .A(n27104), .Z(n27106) );
  XOR U26883 ( .A(n27110), .B(n27111), .Z(n27104) );
  AND U26884 ( .A(n1267), .B(n27103), .Z(n27111) );
  XNOR U26885 ( .A(n27101), .B(n27110), .Z(n27103) );
  XNOR U26886 ( .A(n27112), .B(n27113), .Z(n27101) );
  AND U26887 ( .A(n1271), .B(n27114), .Z(n27113) );
  XOR U26888 ( .A(p_input[1930]), .B(n27112), .Z(n27114) );
  XOR U26889 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n27115), 
        .Z(n27112) );
  AND U26890 ( .A(n1274), .B(n27116), .Z(n27115) );
  XOR U26891 ( .A(n27117), .B(n27118), .Z(n27110) );
  AND U26892 ( .A(n1278), .B(n27109), .Z(n27118) );
  XNOR U26893 ( .A(n27119), .B(n27107), .Z(n27109) );
  XOR U26894 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n27120), .Z(n27107) );
  AND U26895 ( .A(n1290), .B(n27121), .Z(n27120) );
  IV U26896 ( .A(n27117), .Z(n27119) );
  XOR U26897 ( .A(n27122), .B(n27123), .Z(n27117) );
  AND U26898 ( .A(n1285), .B(n27116), .Z(n27123) );
  XOR U26899 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n27122), 
        .Z(n27116) );
  XOR U26900 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(n27124), 
        .Z(n27122) );
  AND U26901 ( .A(n1287), .B(n27121), .Z(n27124) );
  XOR U26902 ( .A(\knn_comb_/min_val_out[0][10] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n27121) );
  XOR U26903 ( .A(n6467), .B(n27125), .Z(o[0]) );
  AND U26904 ( .A(n122), .B(n27126), .Z(n6467) );
  XOR U26905 ( .A(n6468), .B(n27125), .Z(n27126) );
  XOR U26906 ( .A(n27127), .B(n27128), .Z(n27125) );
  AND U26907 ( .A(n142), .B(n27129), .Z(n27128) );
  XOR U26908 ( .A(n27130), .B(n71), .Z(n6468) );
  AND U26909 ( .A(n125), .B(n27131), .Z(n71) );
  XOR U26910 ( .A(n72), .B(n27130), .Z(n27131) );
  XOR U26911 ( .A(n27132), .B(n27133), .Z(n72) );
  AND U26912 ( .A(n130), .B(n27134), .Z(n27133) );
  XOR U26913 ( .A(p_input[0]), .B(n27132), .Z(n27134) );
  XNOR U26914 ( .A(n27135), .B(n27136), .Z(n27132) );
  AND U26915 ( .A(n134), .B(n27137), .Z(n27136) );
  XOR U26916 ( .A(n27138), .B(n27139), .Z(n27130) );
  AND U26917 ( .A(n138), .B(n27129), .Z(n27139) );
  XNOR U26918 ( .A(n27140), .B(n27127), .Z(n27129) );
  XOR U26919 ( .A(n27141), .B(n27142), .Z(n27127) );
  AND U26920 ( .A(n162), .B(n27143), .Z(n27142) );
  IV U26921 ( .A(n27138), .Z(n27140) );
  XOR U26922 ( .A(n27144), .B(n27145), .Z(n27138) );
  AND U26923 ( .A(n146), .B(n27137), .Z(n27145) );
  XNOR U26924 ( .A(n27135), .B(n27144), .Z(n27137) );
  XNOR U26925 ( .A(n27146), .B(n27147), .Z(n27135) );
  AND U26926 ( .A(n150), .B(n27148), .Z(n27147) );
  XOR U26927 ( .A(p_input[32]), .B(n27146), .Z(n27148) );
  XNOR U26928 ( .A(n27149), .B(n27150), .Z(n27146) );
  AND U26929 ( .A(n154), .B(n27151), .Z(n27150) );
  XOR U26930 ( .A(n27152), .B(n27153), .Z(n27144) );
  AND U26931 ( .A(n158), .B(n27143), .Z(n27153) );
  XNOR U26932 ( .A(n27154), .B(n27141), .Z(n27143) );
  XOR U26933 ( .A(n27155), .B(n27156), .Z(n27141) );
  AND U26934 ( .A(n181), .B(n27157), .Z(n27156) );
  IV U26935 ( .A(n27152), .Z(n27154) );
  XOR U26936 ( .A(n27158), .B(n27159), .Z(n27152) );
  AND U26937 ( .A(n165), .B(n27151), .Z(n27159) );
  XNOR U26938 ( .A(n27149), .B(n27158), .Z(n27151) );
  XNOR U26939 ( .A(n27160), .B(n27161), .Z(n27149) );
  AND U26940 ( .A(n169), .B(n27162), .Z(n27161) );
  XOR U26941 ( .A(p_input[64]), .B(n27160), .Z(n27162) );
  XNOR U26942 ( .A(n27163), .B(n27164), .Z(n27160) );
  AND U26943 ( .A(n173), .B(n27165), .Z(n27164) );
  XOR U26944 ( .A(n27166), .B(n27167), .Z(n27158) );
  AND U26945 ( .A(n177), .B(n27157), .Z(n27167) );
  XNOR U26946 ( .A(n27168), .B(n27155), .Z(n27157) );
  XOR U26947 ( .A(n27169), .B(n27170), .Z(n27155) );
  AND U26948 ( .A(n200), .B(n27171), .Z(n27170) );
  IV U26949 ( .A(n27166), .Z(n27168) );
  XOR U26950 ( .A(n27172), .B(n27173), .Z(n27166) );
  AND U26951 ( .A(n184), .B(n27165), .Z(n27173) );
  XNOR U26952 ( .A(n27163), .B(n27172), .Z(n27165) );
  XNOR U26953 ( .A(n27174), .B(n27175), .Z(n27163) );
  AND U26954 ( .A(n188), .B(n27176), .Z(n27175) );
  XOR U26955 ( .A(p_input[96]), .B(n27174), .Z(n27176) );
  XNOR U26956 ( .A(n27177), .B(n27178), .Z(n27174) );
  AND U26957 ( .A(n192), .B(n27179), .Z(n27178) );
  XOR U26958 ( .A(n27180), .B(n27181), .Z(n27172) );
  AND U26959 ( .A(n196), .B(n27171), .Z(n27181) );
  XNOR U26960 ( .A(n27182), .B(n27169), .Z(n27171) );
  XOR U26961 ( .A(n27183), .B(n27184), .Z(n27169) );
  AND U26962 ( .A(n219), .B(n27185), .Z(n27184) );
  IV U26963 ( .A(n27180), .Z(n27182) );
  XOR U26964 ( .A(n27186), .B(n27187), .Z(n27180) );
  AND U26965 ( .A(n203), .B(n27179), .Z(n27187) );
  XNOR U26966 ( .A(n27177), .B(n27186), .Z(n27179) );
  XNOR U26967 ( .A(n27188), .B(n27189), .Z(n27177) );
  AND U26968 ( .A(n207), .B(n27190), .Z(n27189) );
  XOR U26969 ( .A(p_input[128]), .B(n27188), .Z(n27190) );
  XNOR U26970 ( .A(n27191), .B(n27192), .Z(n27188) );
  AND U26971 ( .A(n211), .B(n27193), .Z(n27192) );
  XOR U26972 ( .A(n27194), .B(n27195), .Z(n27186) );
  AND U26973 ( .A(n215), .B(n27185), .Z(n27195) );
  XNOR U26974 ( .A(n27196), .B(n27183), .Z(n27185) );
  XOR U26975 ( .A(n27197), .B(n27198), .Z(n27183) );
  AND U26976 ( .A(n238), .B(n27199), .Z(n27198) );
  IV U26977 ( .A(n27194), .Z(n27196) );
  XOR U26978 ( .A(n27200), .B(n27201), .Z(n27194) );
  AND U26979 ( .A(n222), .B(n27193), .Z(n27201) );
  XNOR U26980 ( .A(n27191), .B(n27200), .Z(n27193) );
  XNOR U26981 ( .A(n27202), .B(n27203), .Z(n27191) );
  AND U26982 ( .A(n226), .B(n27204), .Z(n27203) );
  XOR U26983 ( .A(p_input[160]), .B(n27202), .Z(n27204) );
  XNOR U26984 ( .A(n27205), .B(n27206), .Z(n27202) );
  AND U26985 ( .A(n230), .B(n27207), .Z(n27206) );
  XOR U26986 ( .A(n27208), .B(n27209), .Z(n27200) );
  AND U26987 ( .A(n234), .B(n27199), .Z(n27209) );
  XNOR U26988 ( .A(n27210), .B(n27197), .Z(n27199) );
  XOR U26989 ( .A(n27211), .B(n27212), .Z(n27197) );
  AND U26990 ( .A(n257), .B(n27213), .Z(n27212) );
  IV U26991 ( .A(n27208), .Z(n27210) );
  XOR U26992 ( .A(n27214), .B(n27215), .Z(n27208) );
  AND U26993 ( .A(n241), .B(n27207), .Z(n27215) );
  XNOR U26994 ( .A(n27205), .B(n27214), .Z(n27207) );
  XNOR U26995 ( .A(n27216), .B(n27217), .Z(n27205) );
  AND U26996 ( .A(n245), .B(n27218), .Z(n27217) );
  XOR U26997 ( .A(p_input[192]), .B(n27216), .Z(n27218) );
  XNOR U26998 ( .A(n27219), .B(n27220), .Z(n27216) );
  AND U26999 ( .A(n249), .B(n27221), .Z(n27220) );
  XOR U27000 ( .A(n27222), .B(n27223), .Z(n27214) );
  AND U27001 ( .A(n253), .B(n27213), .Z(n27223) );
  XNOR U27002 ( .A(n27224), .B(n27211), .Z(n27213) );
  XOR U27003 ( .A(n27225), .B(n27226), .Z(n27211) );
  AND U27004 ( .A(n276), .B(n27227), .Z(n27226) );
  IV U27005 ( .A(n27222), .Z(n27224) );
  XOR U27006 ( .A(n27228), .B(n27229), .Z(n27222) );
  AND U27007 ( .A(n260), .B(n27221), .Z(n27229) );
  XNOR U27008 ( .A(n27219), .B(n27228), .Z(n27221) );
  XNOR U27009 ( .A(n27230), .B(n27231), .Z(n27219) );
  AND U27010 ( .A(n264), .B(n27232), .Z(n27231) );
  XOR U27011 ( .A(p_input[224]), .B(n27230), .Z(n27232) );
  XNOR U27012 ( .A(n27233), .B(n27234), .Z(n27230) );
  AND U27013 ( .A(n268), .B(n27235), .Z(n27234) );
  XOR U27014 ( .A(n27236), .B(n27237), .Z(n27228) );
  AND U27015 ( .A(n272), .B(n27227), .Z(n27237) );
  XNOR U27016 ( .A(n27238), .B(n27225), .Z(n27227) );
  XOR U27017 ( .A(n27239), .B(n27240), .Z(n27225) );
  AND U27018 ( .A(n295), .B(n27241), .Z(n27240) );
  IV U27019 ( .A(n27236), .Z(n27238) );
  XOR U27020 ( .A(n27242), .B(n27243), .Z(n27236) );
  AND U27021 ( .A(n279), .B(n27235), .Z(n27243) );
  XNOR U27022 ( .A(n27233), .B(n27242), .Z(n27235) );
  XNOR U27023 ( .A(n27244), .B(n27245), .Z(n27233) );
  AND U27024 ( .A(n283), .B(n27246), .Z(n27245) );
  XOR U27025 ( .A(p_input[256]), .B(n27244), .Z(n27246) );
  XNOR U27026 ( .A(n27247), .B(n27248), .Z(n27244) );
  AND U27027 ( .A(n287), .B(n27249), .Z(n27248) );
  XOR U27028 ( .A(n27250), .B(n27251), .Z(n27242) );
  AND U27029 ( .A(n291), .B(n27241), .Z(n27251) );
  XNOR U27030 ( .A(n27252), .B(n27239), .Z(n27241) );
  XOR U27031 ( .A(n27253), .B(n27254), .Z(n27239) );
  AND U27032 ( .A(n314), .B(n27255), .Z(n27254) );
  IV U27033 ( .A(n27250), .Z(n27252) );
  XOR U27034 ( .A(n27256), .B(n27257), .Z(n27250) );
  AND U27035 ( .A(n298), .B(n27249), .Z(n27257) );
  XNOR U27036 ( .A(n27247), .B(n27256), .Z(n27249) );
  XNOR U27037 ( .A(n27258), .B(n27259), .Z(n27247) );
  AND U27038 ( .A(n302), .B(n27260), .Z(n27259) );
  XOR U27039 ( .A(p_input[288]), .B(n27258), .Z(n27260) );
  XNOR U27040 ( .A(n27261), .B(n27262), .Z(n27258) );
  AND U27041 ( .A(n306), .B(n27263), .Z(n27262) );
  XOR U27042 ( .A(n27264), .B(n27265), .Z(n27256) );
  AND U27043 ( .A(n310), .B(n27255), .Z(n27265) );
  XNOR U27044 ( .A(n27266), .B(n27253), .Z(n27255) );
  XOR U27045 ( .A(n27267), .B(n27268), .Z(n27253) );
  AND U27046 ( .A(n333), .B(n27269), .Z(n27268) );
  IV U27047 ( .A(n27264), .Z(n27266) );
  XOR U27048 ( .A(n27270), .B(n27271), .Z(n27264) );
  AND U27049 ( .A(n317), .B(n27263), .Z(n27271) );
  XNOR U27050 ( .A(n27261), .B(n27270), .Z(n27263) );
  XNOR U27051 ( .A(n27272), .B(n27273), .Z(n27261) );
  AND U27052 ( .A(n321), .B(n27274), .Z(n27273) );
  XOR U27053 ( .A(p_input[320]), .B(n27272), .Z(n27274) );
  XNOR U27054 ( .A(n27275), .B(n27276), .Z(n27272) );
  AND U27055 ( .A(n325), .B(n27277), .Z(n27276) );
  XOR U27056 ( .A(n27278), .B(n27279), .Z(n27270) );
  AND U27057 ( .A(n329), .B(n27269), .Z(n27279) );
  XNOR U27058 ( .A(n27280), .B(n27267), .Z(n27269) );
  XOR U27059 ( .A(n27281), .B(n27282), .Z(n27267) );
  AND U27060 ( .A(n352), .B(n27283), .Z(n27282) );
  IV U27061 ( .A(n27278), .Z(n27280) );
  XOR U27062 ( .A(n27284), .B(n27285), .Z(n27278) );
  AND U27063 ( .A(n336), .B(n27277), .Z(n27285) );
  XNOR U27064 ( .A(n27275), .B(n27284), .Z(n27277) );
  XNOR U27065 ( .A(n27286), .B(n27287), .Z(n27275) );
  AND U27066 ( .A(n340), .B(n27288), .Z(n27287) );
  XOR U27067 ( .A(p_input[352]), .B(n27286), .Z(n27288) );
  XNOR U27068 ( .A(n27289), .B(n27290), .Z(n27286) );
  AND U27069 ( .A(n344), .B(n27291), .Z(n27290) );
  XOR U27070 ( .A(n27292), .B(n27293), .Z(n27284) );
  AND U27071 ( .A(n348), .B(n27283), .Z(n27293) );
  XNOR U27072 ( .A(n27294), .B(n27281), .Z(n27283) );
  XOR U27073 ( .A(n27295), .B(n27296), .Z(n27281) );
  AND U27074 ( .A(n371), .B(n27297), .Z(n27296) );
  IV U27075 ( .A(n27292), .Z(n27294) );
  XOR U27076 ( .A(n27298), .B(n27299), .Z(n27292) );
  AND U27077 ( .A(n355), .B(n27291), .Z(n27299) );
  XNOR U27078 ( .A(n27289), .B(n27298), .Z(n27291) );
  XNOR U27079 ( .A(n27300), .B(n27301), .Z(n27289) );
  AND U27080 ( .A(n359), .B(n27302), .Z(n27301) );
  XOR U27081 ( .A(p_input[384]), .B(n27300), .Z(n27302) );
  XNOR U27082 ( .A(n27303), .B(n27304), .Z(n27300) );
  AND U27083 ( .A(n363), .B(n27305), .Z(n27304) );
  XOR U27084 ( .A(n27306), .B(n27307), .Z(n27298) );
  AND U27085 ( .A(n367), .B(n27297), .Z(n27307) );
  XNOR U27086 ( .A(n27308), .B(n27295), .Z(n27297) );
  XOR U27087 ( .A(n27309), .B(n27310), .Z(n27295) );
  AND U27088 ( .A(n390), .B(n27311), .Z(n27310) );
  IV U27089 ( .A(n27306), .Z(n27308) );
  XOR U27090 ( .A(n27312), .B(n27313), .Z(n27306) );
  AND U27091 ( .A(n374), .B(n27305), .Z(n27313) );
  XNOR U27092 ( .A(n27303), .B(n27312), .Z(n27305) );
  XNOR U27093 ( .A(n27314), .B(n27315), .Z(n27303) );
  AND U27094 ( .A(n378), .B(n27316), .Z(n27315) );
  XOR U27095 ( .A(p_input[416]), .B(n27314), .Z(n27316) );
  XNOR U27096 ( .A(n27317), .B(n27318), .Z(n27314) );
  AND U27097 ( .A(n382), .B(n27319), .Z(n27318) );
  XOR U27098 ( .A(n27320), .B(n27321), .Z(n27312) );
  AND U27099 ( .A(n386), .B(n27311), .Z(n27321) );
  XNOR U27100 ( .A(n27322), .B(n27309), .Z(n27311) );
  XOR U27101 ( .A(n27323), .B(n27324), .Z(n27309) );
  AND U27102 ( .A(n409), .B(n27325), .Z(n27324) );
  IV U27103 ( .A(n27320), .Z(n27322) );
  XOR U27104 ( .A(n27326), .B(n27327), .Z(n27320) );
  AND U27105 ( .A(n393), .B(n27319), .Z(n27327) );
  XNOR U27106 ( .A(n27317), .B(n27326), .Z(n27319) );
  XNOR U27107 ( .A(n27328), .B(n27329), .Z(n27317) );
  AND U27108 ( .A(n397), .B(n27330), .Z(n27329) );
  XOR U27109 ( .A(p_input[448]), .B(n27328), .Z(n27330) );
  XNOR U27110 ( .A(n27331), .B(n27332), .Z(n27328) );
  AND U27111 ( .A(n401), .B(n27333), .Z(n27332) );
  XOR U27112 ( .A(n27334), .B(n27335), .Z(n27326) );
  AND U27113 ( .A(n405), .B(n27325), .Z(n27335) );
  XNOR U27114 ( .A(n27336), .B(n27323), .Z(n27325) );
  XOR U27115 ( .A(n27337), .B(n27338), .Z(n27323) );
  AND U27116 ( .A(n428), .B(n27339), .Z(n27338) );
  IV U27117 ( .A(n27334), .Z(n27336) );
  XOR U27118 ( .A(n27340), .B(n27341), .Z(n27334) );
  AND U27119 ( .A(n412), .B(n27333), .Z(n27341) );
  XNOR U27120 ( .A(n27331), .B(n27340), .Z(n27333) );
  XNOR U27121 ( .A(n27342), .B(n27343), .Z(n27331) );
  AND U27122 ( .A(n416), .B(n27344), .Z(n27343) );
  XOR U27123 ( .A(p_input[480]), .B(n27342), .Z(n27344) );
  XNOR U27124 ( .A(n27345), .B(n27346), .Z(n27342) );
  AND U27125 ( .A(n420), .B(n27347), .Z(n27346) );
  XOR U27126 ( .A(n27348), .B(n27349), .Z(n27340) );
  AND U27127 ( .A(n424), .B(n27339), .Z(n27349) );
  XNOR U27128 ( .A(n27350), .B(n27337), .Z(n27339) );
  XOR U27129 ( .A(n27351), .B(n27352), .Z(n27337) );
  AND U27130 ( .A(n447), .B(n27353), .Z(n27352) );
  IV U27131 ( .A(n27348), .Z(n27350) );
  XOR U27132 ( .A(n27354), .B(n27355), .Z(n27348) );
  AND U27133 ( .A(n431), .B(n27347), .Z(n27355) );
  XNOR U27134 ( .A(n27345), .B(n27354), .Z(n27347) );
  XNOR U27135 ( .A(n27356), .B(n27357), .Z(n27345) );
  AND U27136 ( .A(n435), .B(n27358), .Z(n27357) );
  XOR U27137 ( .A(p_input[512]), .B(n27356), .Z(n27358) );
  XNOR U27138 ( .A(n27359), .B(n27360), .Z(n27356) );
  AND U27139 ( .A(n439), .B(n27361), .Z(n27360) );
  XOR U27140 ( .A(n27362), .B(n27363), .Z(n27354) );
  AND U27141 ( .A(n443), .B(n27353), .Z(n27363) );
  XNOR U27142 ( .A(n27364), .B(n27351), .Z(n27353) );
  XOR U27143 ( .A(n27365), .B(n27366), .Z(n27351) );
  AND U27144 ( .A(n466), .B(n27367), .Z(n27366) );
  IV U27145 ( .A(n27362), .Z(n27364) );
  XOR U27146 ( .A(n27368), .B(n27369), .Z(n27362) );
  AND U27147 ( .A(n450), .B(n27361), .Z(n27369) );
  XNOR U27148 ( .A(n27359), .B(n27368), .Z(n27361) );
  XNOR U27149 ( .A(n27370), .B(n27371), .Z(n27359) );
  AND U27150 ( .A(n454), .B(n27372), .Z(n27371) );
  XOR U27151 ( .A(p_input[544]), .B(n27370), .Z(n27372) );
  XNOR U27152 ( .A(n27373), .B(n27374), .Z(n27370) );
  AND U27153 ( .A(n458), .B(n27375), .Z(n27374) );
  XOR U27154 ( .A(n27376), .B(n27377), .Z(n27368) );
  AND U27155 ( .A(n462), .B(n27367), .Z(n27377) );
  XNOR U27156 ( .A(n27378), .B(n27365), .Z(n27367) );
  XOR U27157 ( .A(n27379), .B(n27380), .Z(n27365) );
  AND U27158 ( .A(n485), .B(n27381), .Z(n27380) );
  IV U27159 ( .A(n27376), .Z(n27378) );
  XOR U27160 ( .A(n27382), .B(n27383), .Z(n27376) );
  AND U27161 ( .A(n469), .B(n27375), .Z(n27383) );
  XNOR U27162 ( .A(n27373), .B(n27382), .Z(n27375) );
  XNOR U27163 ( .A(n27384), .B(n27385), .Z(n27373) );
  AND U27164 ( .A(n473), .B(n27386), .Z(n27385) );
  XOR U27165 ( .A(p_input[576]), .B(n27384), .Z(n27386) );
  XNOR U27166 ( .A(n27387), .B(n27388), .Z(n27384) );
  AND U27167 ( .A(n477), .B(n27389), .Z(n27388) );
  XOR U27168 ( .A(n27390), .B(n27391), .Z(n27382) );
  AND U27169 ( .A(n481), .B(n27381), .Z(n27391) );
  XNOR U27170 ( .A(n27392), .B(n27379), .Z(n27381) );
  XOR U27171 ( .A(n27393), .B(n27394), .Z(n27379) );
  AND U27172 ( .A(n504), .B(n27395), .Z(n27394) );
  IV U27173 ( .A(n27390), .Z(n27392) );
  XOR U27174 ( .A(n27396), .B(n27397), .Z(n27390) );
  AND U27175 ( .A(n488), .B(n27389), .Z(n27397) );
  XNOR U27176 ( .A(n27387), .B(n27396), .Z(n27389) );
  XNOR U27177 ( .A(n27398), .B(n27399), .Z(n27387) );
  AND U27178 ( .A(n492), .B(n27400), .Z(n27399) );
  XOR U27179 ( .A(p_input[608]), .B(n27398), .Z(n27400) );
  XNOR U27180 ( .A(n27401), .B(n27402), .Z(n27398) );
  AND U27181 ( .A(n496), .B(n27403), .Z(n27402) );
  XOR U27182 ( .A(n27404), .B(n27405), .Z(n27396) );
  AND U27183 ( .A(n500), .B(n27395), .Z(n27405) );
  XNOR U27184 ( .A(n27406), .B(n27393), .Z(n27395) );
  XOR U27185 ( .A(n27407), .B(n27408), .Z(n27393) );
  AND U27186 ( .A(n523), .B(n27409), .Z(n27408) );
  IV U27187 ( .A(n27404), .Z(n27406) );
  XOR U27188 ( .A(n27410), .B(n27411), .Z(n27404) );
  AND U27189 ( .A(n507), .B(n27403), .Z(n27411) );
  XNOR U27190 ( .A(n27401), .B(n27410), .Z(n27403) );
  XNOR U27191 ( .A(n27412), .B(n27413), .Z(n27401) );
  AND U27192 ( .A(n511), .B(n27414), .Z(n27413) );
  XOR U27193 ( .A(p_input[640]), .B(n27412), .Z(n27414) );
  XNOR U27194 ( .A(n27415), .B(n27416), .Z(n27412) );
  AND U27195 ( .A(n515), .B(n27417), .Z(n27416) );
  XOR U27196 ( .A(n27418), .B(n27419), .Z(n27410) );
  AND U27197 ( .A(n519), .B(n27409), .Z(n27419) );
  XNOR U27198 ( .A(n27420), .B(n27407), .Z(n27409) );
  XOR U27199 ( .A(n27421), .B(n27422), .Z(n27407) );
  AND U27200 ( .A(n542), .B(n27423), .Z(n27422) );
  IV U27201 ( .A(n27418), .Z(n27420) );
  XOR U27202 ( .A(n27424), .B(n27425), .Z(n27418) );
  AND U27203 ( .A(n526), .B(n27417), .Z(n27425) );
  XNOR U27204 ( .A(n27415), .B(n27424), .Z(n27417) );
  XNOR U27205 ( .A(n27426), .B(n27427), .Z(n27415) );
  AND U27206 ( .A(n530), .B(n27428), .Z(n27427) );
  XOR U27207 ( .A(p_input[672]), .B(n27426), .Z(n27428) );
  XNOR U27208 ( .A(n27429), .B(n27430), .Z(n27426) );
  AND U27209 ( .A(n534), .B(n27431), .Z(n27430) );
  XOR U27210 ( .A(n27432), .B(n27433), .Z(n27424) );
  AND U27211 ( .A(n538), .B(n27423), .Z(n27433) );
  XNOR U27212 ( .A(n27434), .B(n27421), .Z(n27423) );
  XOR U27213 ( .A(n27435), .B(n27436), .Z(n27421) );
  AND U27214 ( .A(n561), .B(n27437), .Z(n27436) );
  IV U27215 ( .A(n27432), .Z(n27434) );
  XOR U27216 ( .A(n27438), .B(n27439), .Z(n27432) );
  AND U27217 ( .A(n545), .B(n27431), .Z(n27439) );
  XNOR U27218 ( .A(n27429), .B(n27438), .Z(n27431) );
  XNOR U27219 ( .A(n27440), .B(n27441), .Z(n27429) );
  AND U27220 ( .A(n549), .B(n27442), .Z(n27441) );
  XOR U27221 ( .A(p_input[704]), .B(n27440), .Z(n27442) );
  XNOR U27222 ( .A(n27443), .B(n27444), .Z(n27440) );
  AND U27223 ( .A(n553), .B(n27445), .Z(n27444) );
  XOR U27224 ( .A(n27446), .B(n27447), .Z(n27438) );
  AND U27225 ( .A(n557), .B(n27437), .Z(n27447) );
  XNOR U27226 ( .A(n27448), .B(n27435), .Z(n27437) );
  XOR U27227 ( .A(n27449), .B(n27450), .Z(n27435) );
  AND U27228 ( .A(n580), .B(n27451), .Z(n27450) );
  IV U27229 ( .A(n27446), .Z(n27448) );
  XOR U27230 ( .A(n27452), .B(n27453), .Z(n27446) );
  AND U27231 ( .A(n564), .B(n27445), .Z(n27453) );
  XNOR U27232 ( .A(n27443), .B(n27452), .Z(n27445) );
  XNOR U27233 ( .A(n27454), .B(n27455), .Z(n27443) );
  AND U27234 ( .A(n568), .B(n27456), .Z(n27455) );
  XOR U27235 ( .A(p_input[736]), .B(n27454), .Z(n27456) );
  XNOR U27236 ( .A(n27457), .B(n27458), .Z(n27454) );
  AND U27237 ( .A(n572), .B(n27459), .Z(n27458) );
  XOR U27238 ( .A(n27460), .B(n27461), .Z(n27452) );
  AND U27239 ( .A(n576), .B(n27451), .Z(n27461) );
  XNOR U27240 ( .A(n27462), .B(n27449), .Z(n27451) );
  XOR U27241 ( .A(n27463), .B(n27464), .Z(n27449) );
  AND U27242 ( .A(n599), .B(n27465), .Z(n27464) );
  IV U27243 ( .A(n27460), .Z(n27462) );
  XOR U27244 ( .A(n27466), .B(n27467), .Z(n27460) );
  AND U27245 ( .A(n583), .B(n27459), .Z(n27467) );
  XNOR U27246 ( .A(n27457), .B(n27466), .Z(n27459) );
  XNOR U27247 ( .A(n27468), .B(n27469), .Z(n27457) );
  AND U27248 ( .A(n587), .B(n27470), .Z(n27469) );
  XOR U27249 ( .A(p_input[768]), .B(n27468), .Z(n27470) );
  XNOR U27250 ( .A(n27471), .B(n27472), .Z(n27468) );
  AND U27251 ( .A(n591), .B(n27473), .Z(n27472) );
  XOR U27252 ( .A(n27474), .B(n27475), .Z(n27466) );
  AND U27253 ( .A(n595), .B(n27465), .Z(n27475) );
  XNOR U27254 ( .A(n27476), .B(n27463), .Z(n27465) );
  XOR U27255 ( .A(n27477), .B(n27478), .Z(n27463) );
  AND U27256 ( .A(n618), .B(n27479), .Z(n27478) );
  IV U27257 ( .A(n27474), .Z(n27476) );
  XOR U27258 ( .A(n27480), .B(n27481), .Z(n27474) );
  AND U27259 ( .A(n602), .B(n27473), .Z(n27481) );
  XNOR U27260 ( .A(n27471), .B(n27480), .Z(n27473) );
  XNOR U27261 ( .A(n27482), .B(n27483), .Z(n27471) );
  AND U27262 ( .A(n606), .B(n27484), .Z(n27483) );
  XOR U27263 ( .A(p_input[800]), .B(n27482), .Z(n27484) );
  XNOR U27264 ( .A(n27485), .B(n27486), .Z(n27482) );
  AND U27265 ( .A(n610), .B(n27487), .Z(n27486) );
  XOR U27266 ( .A(n27488), .B(n27489), .Z(n27480) );
  AND U27267 ( .A(n614), .B(n27479), .Z(n27489) );
  XNOR U27268 ( .A(n27490), .B(n27477), .Z(n27479) );
  XOR U27269 ( .A(n27491), .B(n27492), .Z(n27477) );
  AND U27270 ( .A(n637), .B(n27493), .Z(n27492) );
  IV U27271 ( .A(n27488), .Z(n27490) );
  XOR U27272 ( .A(n27494), .B(n27495), .Z(n27488) );
  AND U27273 ( .A(n621), .B(n27487), .Z(n27495) );
  XNOR U27274 ( .A(n27485), .B(n27494), .Z(n27487) );
  XNOR U27275 ( .A(n27496), .B(n27497), .Z(n27485) );
  AND U27276 ( .A(n625), .B(n27498), .Z(n27497) );
  XOR U27277 ( .A(p_input[832]), .B(n27496), .Z(n27498) );
  XNOR U27278 ( .A(n27499), .B(n27500), .Z(n27496) );
  AND U27279 ( .A(n629), .B(n27501), .Z(n27500) );
  XOR U27280 ( .A(n27502), .B(n27503), .Z(n27494) );
  AND U27281 ( .A(n633), .B(n27493), .Z(n27503) );
  XNOR U27282 ( .A(n27504), .B(n27491), .Z(n27493) );
  XOR U27283 ( .A(n27505), .B(n27506), .Z(n27491) );
  AND U27284 ( .A(n656), .B(n27507), .Z(n27506) );
  IV U27285 ( .A(n27502), .Z(n27504) );
  XOR U27286 ( .A(n27508), .B(n27509), .Z(n27502) );
  AND U27287 ( .A(n640), .B(n27501), .Z(n27509) );
  XNOR U27288 ( .A(n27499), .B(n27508), .Z(n27501) );
  XNOR U27289 ( .A(n27510), .B(n27511), .Z(n27499) );
  AND U27290 ( .A(n644), .B(n27512), .Z(n27511) );
  XOR U27291 ( .A(p_input[864]), .B(n27510), .Z(n27512) );
  XNOR U27292 ( .A(n27513), .B(n27514), .Z(n27510) );
  AND U27293 ( .A(n648), .B(n27515), .Z(n27514) );
  XOR U27294 ( .A(n27516), .B(n27517), .Z(n27508) );
  AND U27295 ( .A(n652), .B(n27507), .Z(n27517) );
  XNOR U27296 ( .A(n27518), .B(n27505), .Z(n27507) );
  XOR U27297 ( .A(n27519), .B(n27520), .Z(n27505) );
  AND U27298 ( .A(n675), .B(n27521), .Z(n27520) );
  IV U27299 ( .A(n27516), .Z(n27518) );
  XOR U27300 ( .A(n27522), .B(n27523), .Z(n27516) );
  AND U27301 ( .A(n659), .B(n27515), .Z(n27523) );
  XNOR U27302 ( .A(n27513), .B(n27522), .Z(n27515) );
  XNOR U27303 ( .A(n27524), .B(n27525), .Z(n27513) );
  AND U27304 ( .A(n663), .B(n27526), .Z(n27525) );
  XOR U27305 ( .A(p_input[896]), .B(n27524), .Z(n27526) );
  XNOR U27306 ( .A(n27527), .B(n27528), .Z(n27524) );
  AND U27307 ( .A(n667), .B(n27529), .Z(n27528) );
  XOR U27308 ( .A(n27530), .B(n27531), .Z(n27522) );
  AND U27309 ( .A(n671), .B(n27521), .Z(n27531) );
  XNOR U27310 ( .A(n27532), .B(n27519), .Z(n27521) );
  XOR U27311 ( .A(n27533), .B(n27534), .Z(n27519) );
  AND U27312 ( .A(n694), .B(n27535), .Z(n27534) );
  IV U27313 ( .A(n27530), .Z(n27532) );
  XOR U27314 ( .A(n27536), .B(n27537), .Z(n27530) );
  AND U27315 ( .A(n678), .B(n27529), .Z(n27537) );
  XNOR U27316 ( .A(n27527), .B(n27536), .Z(n27529) );
  XNOR U27317 ( .A(n27538), .B(n27539), .Z(n27527) );
  AND U27318 ( .A(n682), .B(n27540), .Z(n27539) );
  XOR U27319 ( .A(p_input[928]), .B(n27538), .Z(n27540) );
  XNOR U27320 ( .A(n27541), .B(n27542), .Z(n27538) );
  AND U27321 ( .A(n686), .B(n27543), .Z(n27542) );
  XOR U27322 ( .A(n27544), .B(n27545), .Z(n27536) );
  AND U27323 ( .A(n690), .B(n27535), .Z(n27545) );
  XNOR U27324 ( .A(n27546), .B(n27533), .Z(n27535) );
  XOR U27325 ( .A(n27547), .B(n27548), .Z(n27533) );
  AND U27326 ( .A(n713), .B(n27549), .Z(n27548) );
  IV U27327 ( .A(n27544), .Z(n27546) );
  XOR U27328 ( .A(n27550), .B(n27551), .Z(n27544) );
  AND U27329 ( .A(n697), .B(n27543), .Z(n27551) );
  XNOR U27330 ( .A(n27541), .B(n27550), .Z(n27543) );
  XNOR U27331 ( .A(n27552), .B(n27553), .Z(n27541) );
  AND U27332 ( .A(n701), .B(n27554), .Z(n27553) );
  XOR U27333 ( .A(p_input[960]), .B(n27552), .Z(n27554) );
  XNOR U27334 ( .A(n27555), .B(n27556), .Z(n27552) );
  AND U27335 ( .A(n705), .B(n27557), .Z(n27556) );
  XOR U27336 ( .A(n27558), .B(n27559), .Z(n27550) );
  AND U27337 ( .A(n709), .B(n27549), .Z(n27559) );
  XNOR U27338 ( .A(n27560), .B(n27547), .Z(n27549) );
  XOR U27339 ( .A(n27561), .B(n27562), .Z(n27547) );
  AND U27340 ( .A(n732), .B(n27563), .Z(n27562) );
  IV U27341 ( .A(n27558), .Z(n27560) );
  XOR U27342 ( .A(n27564), .B(n27565), .Z(n27558) );
  AND U27343 ( .A(n716), .B(n27557), .Z(n27565) );
  XNOR U27344 ( .A(n27555), .B(n27564), .Z(n27557) );
  XNOR U27345 ( .A(n27566), .B(n27567), .Z(n27555) );
  AND U27346 ( .A(n720), .B(n27568), .Z(n27567) );
  XOR U27347 ( .A(p_input[992]), .B(n27566), .Z(n27568) );
  XNOR U27348 ( .A(n27569), .B(n27570), .Z(n27566) );
  AND U27349 ( .A(n724), .B(n27571), .Z(n27570) );
  XOR U27350 ( .A(n27572), .B(n27573), .Z(n27564) );
  AND U27351 ( .A(n728), .B(n27563), .Z(n27573) );
  XNOR U27352 ( .A(n27574), .B(n27561), .Z(n27563) );
  XOR U27353 ( .A(n27575), .B(n27576), .Z(n27561) );
  AND U27354 ( .A(n751), .B(n27577), .Z(n27576) );
  IV U27355 ( .A(n27572), .Z(n27574) );
  XOR U27356 ( .A(n27578), .B(n27579), .Z(n27572) );
  AND U27357 ( .A(n735), .B(n27571), .Z(n27579) );
  XNOR U27358 ( .A(n27569), .B(n27578), .Z(n27571) );
  XNOR U27359 ( .A(n27580), .B(n27581), .Z(n27569) );
  AND U27360 ( .A(n739), .B(n27582), .Z(n27581) );
  XOR U27361 ( .A(p_input[1024]), .B(n27580), .Z(n27582) );
  XNOR U27362 ( .A(n27583), .B(n27584), .Z(n27580) );
  AND U27363 ( .A(n743), .B(n27585), .Z(n27584) );
  XOR U27364 ( .A(n27586), .B(n27587), .Z(n27578) );
  AND U27365 ( .A(n747), .B(n27577), .Z(n27587) );
  XNOR U27366 ( .A(n27588), .B(n27575), .Z(n27577) );
  XOR U27367 ( .A(n27589), .B(n27590), .Z(n27575) );
  AND U27368 ( .A(n770), .B(n27591), .Z(n27590) );
  IV U27369 ( .A(n27586), .Z(n27588) );
  XOR U27370 ( .A(n27592), .B(n27593), .Z(n27586) );
  AND U27371 ( .A(n754), .B(n27585), .Z(n27593) );
  XNOR U27372 ( .A(n27583), .B(n27592), .Z(n27585) );
  XNOR U27373 ( .A(n27594), .B(n27595), .Z(n27583) );
  AND U27374 ( .A(n758), .B(n27596), .Z(n27595) );
  XOR U27375 ( .A(p_input[1056]), .B(n27594), .Z(n27596) );
  XNOR U27376 ( .A(n27597), .B(n27598), .Z(n27594) );
  AND U27377 ( .A(n762), .B(n27599), .Z(n27598) );
  XOR U27378 ( .A(n27600), .B(n27601), .Z(n27592) );
  AND U27379 ( .A(n766), .B(n27591), .Z(n27601) );
  XNOR U27380 ( .A(n27602), .B(n27589), .Z(n27591) );
  XOR U27381 ( .A(n27603), .B(n27604), .Z(n27589) );
  AND U27382 ( .A(n789), .B(n27605), .Z(n27604) );
  IV U27383 ( .A(n27600), .Z(n27602) );
  XOR U27384 ( .A(n27606), .B(n27607), .Z(n27600) );
  AND U27385 ( .A(n773), .B(n27599), .Z(n27607) );
  XNOR U27386 ( .A(n27597), .B(n27606), .Z(n27599) );
  XNOR U27387 ( .A(n27608), .B(n27609), .Z(n27597) );
  AND U27388 ( .A(n777), .B(n27610), .Z(n27609) );
  XOR U27389 ( .A(p_input[1088]), .B(n27608), .Z(n27610) );
  XNOR U27390 ( .A(n27611), .B(n27612), .Z(n27608) );
  AND U27391 ( .A(n781), .B(n27613), .Z(n27612) );
  XOR U27392 ( .A(n27614), .B(n27615), .Z(n27606) );
  AND U27393 ( .A(n785), .B(n27605), .Z(n27615) );
  XNOR U27394 ( .A(n27616), .B(n27603), .Z(n27605) );
  XOR U27395 ( .A(n27617), .B(n27618), .Z(n27603) );
  AND U27396 ( .A(n808), .B(n27619), .Z(n27618) );
  IV U27397 ( .A(n27614), .Z(n27616) );
  XOR U27398 ( .A(n27620), .B(n27621), .Z(n27614) );
  AND U27399 ( .A(n792), .B(n27613), .Z(n27621) );
  XNOR U27400 ( .A(n27611), .B(n27620), .Z(n27613) );
  XNOR U27401 ( .A(n27622), .B(n27623), .Z(n27611) );
  AND U27402 ( .A(n796), .B(n27624), .Z(n27623) );
  XOR U27403 ( .A(p_input[1120]), .B(n27622), .Z(n27624) );
  XNOR U27404 ( .A(n27625), .B(n27626), .Z(n27622) );
  AND U27405 ( .A(n800), .B(n27627), .Z(n27626) );
  XOR U27406 ( .A(n27628), .B(n27629), .Z(n27620) );
  AND U27407 ( .A(n804), .B(n27619), .Z(n27629) );
  XNOR U27408 ( .A(n27630), .B(n27617), .Z(n27619) );
  XOR U27409 ( .A(n27631), .B(n27632), .Z(n27617) );
  AND U27410 ( .A(n827), .B(n27633), .Z(n27632) );
  IV U27411 ( .A(n27628), .Z(n27630) );
  XOR U27412 ( .A(n27634), .B(n27635), .Z(n27628) );
  AND U27413 ( .A(n811), .B(n27627), .Z(n27635) );
  XNOR U27414 ( .A(n27625), .B(n27634), .Z(n27627) );
  XNOR U27415 ( .A(n27636), .B(n27637), .Z(n27625) );
  AND U27416 ( .A(n815), .B(n27638), .Z(n27637) );
  XOR U27417 ( .A(p_input[1152]), .B(n27636), .Z(n27638) );
  XNOR U27418 ( .A(n27639), .B(n27640), .Z(n27636) );
  AND U27419 ( .A(n819), .B(n27641), .Z(n27640) );
  XOR U27420 ( .A(n27642), .B(n27643), .Z(n27634) );
  AND U27421 ( .A(n823), .B(n27633), .Z(n27643) );
  XNOR U27422 ( .A(n27644), .B(n27631), .Z(n27633) );
  XOR U27423 ( .A(n27645), .B(n27646), .Z(n27631) );
  AND U27424 ( .A(n846), .B(n27647), .Z(n27646) );
  IV U27425 ( .A(n27642), .Z(n27644) );
  XOR U27426 ( .A(n27648), .B(n27649), .Z(n27642) );
  AND U27427 ( .A(n830), .B(n27641), .Z(n27649) );
  XNOR U27428 ( .A(n27639), .B(n27648), .Z(n27641) );
  XNOR U27429 ( .A(n27650), .B(n27651), .Z(n27639) );
  AND U27430 ( .A(n834), .B(n27652), .Z(n27651) );
  XOR U27431 ( .A(p_input[1184]), .B(n27650), .Z(n27652) );
  XNOR U27432 ( .A(n27653), .B(n27654), .Z(n27650) );
  AND U27433 ( .A(n838), .B(n27655), .Z(n27654) );
  XOR U27434 ( .A(n27656), .B(n27657), .Z(n27648) );
  AND U27435 ( .A(n842), .B(n27647), .Z(n27657) );
  XNOR U27436 ( .A(n27658), .B(n27645), .Z(n27647) );
  XOR U27437 ( .A(n27659), .B(n27660), .Z(n27645) );
  AND U27438 ( .A(n865), .B(n27661), .Z(n27660) );
  IV U27439 ( .A(n27656), .Z(n27658) );
  XOR U27440 ( .A(n27662), .B(n27663), .Z(n27656) );
  AND U27441 ( .A(n849), .B(n27655), .Z(n27663) );
  XNOR U27442 ( .A(n27653), .B(n27662), .Z(n27655) );
  XNOR U27443 ( .A(n27664), .B(n27665), .Z(n27653) );
  AND U27444 ( .A(n853), .B(n27666), .Z(n27665) );
  XOR U27445 ( .A(p_input[1216]), .B(n27664), .Z(n27666) );
  XNOR U27446 ( .A(n27667), .B(n27668), .Z(n27664) );
  AND U27447 ( .A(n857), .B(n27669), .Z(n27668) );
  XOR U27448 ( .A(n27670), .B(n27671), .Z(n27662) );
  AND U27449 ( .A(n861), .B(n27661), .Z(n27671) );
  XNOR U27450 ( .A(n27672), .B(n27659), .Z(n27661) );
  XOR U27451 ( .A(n27673), .B(n27674), .Z(n27659) );
  AND U27452 ( .A(n884), .B(n27675), .Z(n27674) );
  IV U27453 ( .A(n27670), .Z(n27672) );
  XOR U27454 ( .A(n27676), .B(n27677), .Z(n27670) );
  AND U27455 ( .A(n868), .B(n27669), .Z(n27677) );
  XNOR U27456 ( .A(n27667), .B(n27676), .Z(n27669) );
  XNOR U27457 ( .A(n27678), .B(n27679), .Z(n27667) );
  AND U27458 ( .A(n872), .B(n27680), .Z(n27679) );
  XOR U27459 ( .A(p_input[1248]), .B(n27678), .Z(n27680) );
  XNOR U27460 ( .A(n27681), .B(n27682), .Z(n27678) );
  AND U27461 ( .A(n876), .B(n27683), .Z(n27682) );
  XOR U27462 ( .A(n27684), .B(n27685), .Z(n27676) );
  AND U27463 ( .A(n880), .B(n27675), .Z(n27685) );
  XNOR U27464 ( .A(n27686), .B(n27673), .Z(n27675) );
  XOR U27465 ( .A(n27687), .B(n27688), .Z(n27673) );
  AND U27466 ( .A(n903), .B(n27689), .Z(n27688) );
  IV U27467 ( .A(n27684), .Z(n27686) );
  XOR U27468 ( .A(n27690), .B(n27691), .Z(n27684) );
  AND U27469 ( .A(n887), .B(n27683), .Z(n27691) );
  XNOR U27470 ( .A(n27681), .B(n27690), .Z(n27683) );
  XNOR U27471 ( .A(n27692), .B(n27693), .Z(n27681) );
  AND U27472 ( .A(n891), .B(n27694), .Z(n27693) );
  XOR U27473 ( .A(p_input[1280]), .B(n27692), .Z(n27694) );
  XNOR U27474 ( .A(n27695), .B(n27696), .Z(n27692) );
  AND U27475 ( .A(n895), .B(n27697), .Z(n27696) );
  XOR U27476 ( .A(n27698), .B(n27699), .Z(n27690) );
  AND U27477 ( .A(n899), .B(n27689), .Z(n27699) );
  XNOR U27478 ( .A(n27700), .B(n27687), .Z(n27689) );
  XOR U27479 ( .A(n27701), .B(n27702), .Z(n27687) );
  AND U27480 ( .A(n922), .B(n27703), .Z(n27702) );
  IV U27481 ( .A(n27698), .Z(n27700) );
  XOR U27482 ( .A(n27704), .B(n27705), .Z(n27698) );
  AND U27483 ( .A(n906), .B(n27697), .Z(n27705) );
  XNOR U27484 ( .A(n27695), .B(n27704), .Z(n27697) );
  XNOR U27485 ( .A(n27706), .B(n27707), .Z(n27695) );
  AND U27486 ( .A(n910), .B(n27708), .Z(n27707) );
  XOR U27487 ( .A(p_input[1312]), .B(n27706), .Z(n27708) );
  XNOR U27488 ( .A(n27709), .B(n27710), .Z(n27706) );
  AND U27489 ( .A(n914), .B(n27711), .Z(n27710) );
  XOR U27490 ( .A(n27712), .B(n27713), .Z(n27704) );
  AND U27491 ( .A(n918), .B(n27703), .Z(n27713) );
  XNOR U27492 ( .A(n27714), .B(n27701), .Z(n27703) );
  XOR U27493 ( .A(n27715), .B(n27716), .Z(n27701) );
  AND U27494 ( .A(n941), .B(n27717), .Z(n27716) );
  IV U27495 ( .A(n27712), .Z(n27714) );
  XOR U27496 ( .A(n27718), .B(n27719), .Z(n27712) );
  AND U27497 ( .A(n925), .B(n27711), .Z(n27719) );
  XNOR U27498 ( .A(n27709), .B(n27718), .Z(n27711) );
  XNOR U27499 ( .A(n27720), .B(n27721), .Z(n27709) );
  AND U27500 ( .A(n929), .B(n27722), .Z(n27721) );
  XOR U27501 ( .A(p_input[1344]), .B(n27720), .Z(n27722) );
  XNOR U27502 ( .A(n27723), .B(n27724), .Z(n27720) );
  AND U27503 ( .A(n933), .B(n27725), .Z(n27724) );
  XOR U27504 ( .A(n27726), .B(n27727), .Z(n27718) );
  AND U27505 ( .A(n937), .B(n27717), .Z(n27727) );
  XNOR U27506 ( .A(n27728), .B(n27715), .Z(n27717) );
  XOR U27507 ( .A(n27729), .B(n27730), .Z(n27715) );
  AND U27508 ( .A(n960), .B(n27731), .Z(n27730) );
  IV U27509 ( .A(n27726), .Z(n27728) );
  XOR U27510 ( .A(n27732), .B(n27733), .Z(n27726) );
  AND U27511 ( .A(n944), .B(n27725), .Z(n27733) );
  XNOR U27512 ( .A(n27723), .B(n27732), .Z(n27725) );
  XNOR U27513 ( .A(n27734), .B(n27735), .Z(n27723) );
  AND U27514 ( .A(n948), .B(n27736), .Z(n27735) );
  XOR U27515 ( .A(p_input[1376]), .B(n27734), .Z(n27736) );
  XNOR U27516 ( .A(n27737), .B(n27738), .Z(n27734) );
  AND U27517 ( .A(n952), .B(n27739), .Z(n27738) );
  XOR U27518 ( .A(n27740), .B(n27741), .Z(n27732) );
  AND U27519 ( .A(n956), .B(n27731), .Z(n27741) );
  XNOR U27520 ( .A(n27742), .B(n27729), .Z(n27731) );
  XOR U27521 ( .A(n27743), .B(n27744), .Z(n27729) );
  AND U27522 ( .A(n979), .B(n27745), .Z(n27744) );
  IV U27523 ( .A(n27740), .Z(n27742) );
  XOR U27524 ( .A(n27746), .B(n27747), .Z(n27740) );
  AND U27525 ( .A(n963), .B(n27739), .Z(n27747) );
  XNOR U27526 ( .A(n27737), .B(n27746), .Z(n27739) );
  XNOR U27527 ( .A(n27748), .B(n27749), .Z(n27737) );
  AND U27528 ( .A(n967), .B(n27750), .Z(n27749) );
  XOR U27529 ( .A(p_input[1408]), .B(n27748), .Z(n27750) );
  XNOR U27530 ( .A(n27751), .B(n27752), .Z(n27748) );
  AND U27531 ( .A(n971), .B(n27753), .Z(n27752) );
  XOR U27532 ( .A(n27754), .B(n27755), .Z(n27746) );
  AND U27533 ( .A(n975), .B(n27745), .Z(n27755) );
  XNOR U27534 ( .A(n27756), .B(n27743), .Z(n27745) );
  XOR U27535 ( .A(n27757), .B(n27758), .Z(n27743) );
  AND U27536 ( .A(n998), .B(n27759), .Z(n27758) );
  IV U27537 ( .A(n27754), .Z(n27756) );
  XOR U27538 ( .A(n27760), .B(n27761), .Z(n27754) );
  AND U27539 ( .A(n982), .B(n27753), .Z(n27761) );
  XNOR U27540 ( .A(n27751), .B(n27760), .Z(n27753) );
  XNOR U27541 ( .A(n27762), .B(n27763), .Z(n27751) );
  AND U27542 ( .A(n986), .B(n27764), .Z(n27763) );
  XOR U27543 ( .A(p_input[1440]), .B(n27762), .Z(n27764) );
  XNOR U27544 ( .A(n27765), .B(n27766), .Z(n27762) );
  AND U27545 ( .A(n990), .B(n27767), .Z(n27766) );
  XOR U27546 ( .A(n27768), .B(n27769), .Z(n27760) );
  AND U27547 ( .A(n994), .B(n27759), .Z(n27769) );
  XNOR U27548 ( .A(n27770), .B(n27757), .Z(n27759) );
  XOR U27549 ( .A(n27771), .B(n27772), .Z(n27757) );
  AND U27550 ( .A(n1017), .B(n27773), .Z(n27772) );
  IV U27551 ( .A(n27768), .Z(n27770) );
  XOR U27552 ( .A(n27774), .B(n27775), .Z(n27768) );
  AND U27553 ( .A(n1001), .B(n27767), .Z(n27775) );
  XNOR U27554 ( .A(n27765), .B(n27774), .Z(n27767) );
  XNOR U27555 ( .A(n27776), .B(n27777), .Z(n27765) );
  AND U27556 ( .A(n1005), .B(n27778), .Z(n27777) );
  XOR U27557 ( .A(p_input[1472]), .B(n27776), .Z(n27778) );
  XNOR U27558 ( .A(n27779), .B(n27780), .Z(n27776) );
  AND U27559 ( .A(n1009), .B(n27781), .Z(n27780) );
  XOR U27560 ( .A(n27782), .B(n27783), .Z(n27774) );
  AND U27561 ( .A(n1013), .B(n27773), .Z(n27783) );
  XNOR U27562 ( .A(n27784), .B(n27771), .Z(n27773) );
  XOR U27563 ( .A(n27785), .B(n27786), .Z(n27771) );
  AND U27564 ( .A(n1036), .B(n27787), .Z(n27786) );
  IV U27565 ( .A(n27782), .Z(n27784) );
  XOR U27566 ( .A(n27788), .B(n27789), .Z(n27782) );
  AND U27567 ( .A(n1020), .B(n27781), .Z(n27789) );
  XNOR U27568 ( .A(n27779), .B(n27788), .Z(n27781) );
  XNOR U27569 ( .A(n27790), .B(n27791), .Z(n27779) );
  AND U27570 ( .A(n1024), .B(n27792), .Z(n27791) );
  XOR U27571 ( .A(p_input[1504]), .B(n27790), .Z(n27792) );
  XNOR U27572 ( .A(n27793), .B(n27794), .Z(n27790) );
  AND U27573 ( .A(n1028), .B(n27795), .Z(n27794) );
  XOR U27574 ( .A(n27796), .B(n27797), .Z(n27788) );
  AND U27575 ( .A(n1032), .B(n27787), .Z(n27797) );
  XNOR U27576 ( .A(n27798), .B(n27785), .Z(n27787) );
  XOR U27577 ( .A(n27799), .B(n27800), .Z(n27785) );
  AND U27578 ( .A(n1055), .B(n27801), .Z(n27800) );
  IV U27579 ( .A(n27796), .Z(n27798) );
  XOR U27580 ( .A(n27802), .B(n27803), .Z(n27796) );
  AND U27581 ( .A(n1039), .B(n27795), .Z(n27803) );
  XNOR U27582 ( .A(n27793), .B(n27802), .Z(n27795) );
  XNOR U27583 ( .A(n27804), .B(n27805), .Z(n27793) );
  AND U27584 ( .A(n1043), .B(n27806), .Z(n27805) );
  XOR U27585 ( .A(p_input[1536]), .B(n27804), .Z(n27806) );
  XNOR U27586 ( .A(n27807), .B(n27808), .Z(n27804) );
  AND U27587 ( .A(n1047), .B(n27809), .Z(n27808) );
  XOR U27588 ( .A(n27810), .B(n27811), .Z(n27802) );
  AND U27589 ( .A(n1051), .B(n27801), .Z(n27811) );
  XNOR U27590 ( .A(n27812), .B(n27799), .Z(n27801) );
  XOR U27591 ( .A(n27813), .B(n27814), .Z(n27799) );
  AND U27592 ( .A(n1074), .B(n27815), .Z(n27814) );
  IV U27593 ( .A(n27810), .Z(n27812) );
  XOR U27594 ( .A(n27816), .B(n27817), .Z(n27810) );
  AND U27595 ( .A(n1058), .B(n27809), .Z(n27817) );
  XNOR U27596 ( .A(n27807), .B(n27816), .Z(n27809) );
  XNOR U27597 ( .A(n27818), .B(n27819), .Z(n27807) );
  AND U27598 ( .A(n1062), .B(n27820), .Z(n27819) );
  XOR U27599 ( .A(p_input[1568]), .B(n27818), .Z(n27820) );
  XNOR U27600 ( .A(n27821), .B(n27822), .Z(n27818) );
  AND U27601 ( .A(n1066), .B(n27823), .Z(n27822) );
  XOR U27602 ( .A(n27824), .B(n27825), .Z(n27816) );
  AND U27603 ( .A(n1070), .B(n27815), .Z(n27825) );
  XNOR U27604 ( .A(n27826), .B(n27813), .Z(n27815) );
  XOR U27605 ( .A(n27827), .B(n27828), .Z(n27813) );
  AND U27606 ( .A(n1093), .B(n27829), .Z(n27828) );
  IV U27607 ( .A(n27824), .Z(n27826) );
  XOR U27608 ( .A(n27830), .B(n27831), .Z(n27824) );
  AND U27609 ( .A(n1077), .B(n27823), .Z(n27831) );
  XNOR U27610 ( .A(n27821), .B(n27830), .Z(n27823) );
  XNOR U27611 ( .A(n27832), .B(n27833), .Z(n27821) );
  AND U27612 ( .A(n1081), .B(n27834), .Z(n27833) );
  XOR U27613 ( .A(p_input[1600]), .B(n27832), .Z(n27834) );
  XNOR U27614 ( .A(n27835), .B(n27836), .Z(n27832) );
  AND U27615 ( .A(n1085), .B(n27837), .Z(n27836) );
  XOR U27616 ( .A(n27838), .B(n27839), .Z(n27830) );
  AND U27617 ( .A(n1089), .B(n27829), .Z(n27839) );
  XNOR U27618 ( .A(n27840), .B(n27827), .Z(n27829) );
  XOR U27619 ( .A(n27841), .B(n27842), .Z(n27827) );
  AND U27620 ( .A(n1112), .B(n27843), .Z(n27842) );
  IV U27621 ( .A(n27838), .Z(n27840) );
  XOR U27622 ( .A(n27844), .B(n27845), .Z(n27838) );
  AND U27623 ( .A(n1096), .B(n27837), .Z(n27845) );
  XNOR U27624 ( .A(n27835), .B(n27844), .Z(n27837) );
  XNOR U27625 ( .A(n27846), .B(n27847), .Z(n27835) );
  AND U27626 ( .A(n1100), .B(n27848), .Z(n27847) );
  XOR U27627 ( .A(p_input[1632]), .B(n27846), .Z(n27848) );
  XNOR U27628 ( .A(n27849), .B(n27850), .Z(n27846) );
  AND U27629 ( .A(n1104), .B(n27851), .Z(n27850) );
  XOR U27630 ( .A(n27852), .B(n27853), .Z(n27844) );
  AND U27631 ( .A(n1108), .B(n27843), .Z(n27853) );
  XNOR U27632 ( .A(n27854), .B(n27841), .Z(n27843) );
  XOR U27633 ( .A(n27855), .B(n27856), .Z(n27841) );
  AND U27634 ( .A(n1131), .B(n27857), .Z(n27856) );
  IV U27635 ( .A(n27852), .Z(n27854) );
  XOR U27636 ( .A(n27858), .B(n27859), .Z(n27852) );
  AND U27637 ( .A(n1115), .B(n27851), .Z(n27859) );
  XNOR U27638 ( .A(n27849), .B(n27858), .Z(n27851) );
  XNOR U27639 ( .A(n27860), .B(n27861), .Z(n27849) );
  AND U27640 ( .A(n1119), .B(n27862), .Z(n27861) );
  XOR U27641 ( .A(p_input[1664]), .B(n27860), .Z(n27862) );
  XNOR U27642 ( .A(n27863), .B(n27864), .Z(n27860) );
  AND U27643 ( .A(n1123), .B(n27865), .Z(n27864) );
  XOR U27644 ( .A(n27866), .B(n27867), .Z(n27858) );
  AND U27645 ( .A(n1127), .B(n27857), .Z(n27867) );
  XNOR U27646 ( .A(n27868), .B(n27855), .Z(n27857) );
  XOR U27647 ( .A(n27869), .B(n27870), .Z(n27855) );
  AND U27648 ( .A(n1150), .B(n27871), .Z(n27870) );
  IV U27649 ( .A(n27866), .Z(n27868) );
  XOR U27650 ( .A(n27872), .B(n27873), .Z(n27866) );
  AND U27651 ( .A(n1134), .B(n27865), .Z(n27873) );
  XNOR U27652 ( .A(n27863), .B(n27872), .Z(n27865) );
  XNOR U27653 ( .A(n27874), .B(n27875), .Z(n27863) );
  AND U27654 ( .A(n1138), .B(n27876), .Z(n27875) );
  XOR U27655 ( .A(p_input[1696]), .B(n27874), .Z(n27876) );
  XNOR U27656 ( .A(n27877), .B(n27878), .Z(n27874) );
  AND U27657 ( .A(n1142), .B(n27879), .Z(n27878) );
  XOR U27658 ( .A(n27880), .B(n27881), .Z(n27872) );
  AND U27659 ( .A(n1146), .B(n27871), .Z(n27881) );
  XNOR U27660 ( .A(n27882), .B(n27869), .Z(n27871) );
  XOR U27661 ( .A(n27883), .B(n27884), .Z(n27869) );
  AND U27662 ( .A(n1169), .B(n27885), .Z(n27884) );
  IV U27663 ( .A(n27880), .Z(n27882) );
  XOR U27664 ( .A(n27886), .B(n27887), .Z(n27880) );
  AND U27665 ( .A(n1153), .B(n27879), .Z(n27887) );
  XNOR U27666 ( .A(n27877), .B(n27886), .Z(n27879) );
  XNOR U27667 ( .A(n27888), .B(n27889), .Z(n27877) );
  AND U27668 ( .A(n1157), .B(n27890), .Z(n27889) );
  XOR U27669 ( .A(p_input[1728]), .B(n27888), .Z(n27890) );
  XNOR U27670 ( .A(n27891), .B(n27892), .Z(n27888) );
  AND U27671 ( .A(n1161), .B(n27893), .Z(n27892) );
  XOR U27672 ( .A(n27894), .B(n27895), .Z(n27886) );
  AND U27673 ( .A(n1165), .B(n27885), .Z(n27895) );
  XNOR U27674 ( .A(n27896), .B(n27883), .Z(n27885) );
  XOR U27675 ( .A(n27897), .B(n27898), .Z(n27883) );
  AND U27676 ( .A(n1188), .B(n27899), .Z(n27898) );
  IV U27677 ( .A(n27894), .Z(n27896) );
  XOR U27678 ( .A(n27900), .B(n27901), .Z(n27894) );
  AND U27679 ( .A(n1172), .B(n27893), .Z(n27901) );
  XNOR U27680 ( .A(n27891), .B(n27900), .Z(n27893) );
  XNOR U27681 ( .A(n27902), .B(n27903), .Z(n27891) );
  AND U27682 ( .A(n1176), .B(n27904), .Z(n27903) );
  XOR U27683 ( .A(p_input[1760]), .B(n27902), .Z(n27904) );
  XNOR U27684 ( .A(n27905), .B(n27906), .Z(n27902) );
  AND U27685 ( .A(n1180), .B(n27907), .Z(n27906) );
  XOR U27686 ( .A(n27908), .B(n27909), .Z(n27900) );
  AND U27687 ( .A(n1184), .B(n27899), .Z(n27909) );
  XNOR U27688 ( .A(n27910), .B(n27897), .Z(n27899) );
  XOR U27689 ( .A(n27911), .B(n27912), .Z(n27897) );
  AND U27690 ( .A(n1207), .B(n27913), .Z(n27912) );
  IV U27691 ( .A(n27908), .Z(n27910) );
  XOR U27692 ( .A(n27914), .B(n27915), .Z(n27908) );
  AND U27693 ( .A(n1191), .B(n27907), .Z(n27915) );
  XNOR U27694 ( .A(n27905), .B(n27914), .Z(n27907) );
  XNOR U27695 ( .A(n27916), .B(n27917), .Z(n27905) );
  AND U27696 ( .A(n1195), .B(n27918), .Z(n27917) );
  XOR U27697 ( .A(p_input[1792]), .B(n27916), .Z(n27918) );
  XNOR U27698 ( .A(n27919), .B(n27920), .Z(n27916) );
  AND U27699 ( .A(n1199), .B(n27921), .Z(n27920) );
  XOR U27700 ( .A(n27922), .B(n27923), .Z(n27914) );
  AND U27701 ( .A(n1203), .B(n27913), .Z(n27923) );
  XNOR U27702 ( .A(n27924), .B(n27911), .Z(n27913) );
  XOR U27703 ( .A(n27925), .B(n27926), .Z(n27911) );
  AND U27704 ( .A(n1226), .B(n27927), .Z(n27926) );
  IV U27705 ( .A(n27922), .Z(n27924) );
  XOR U27706 ( .A(n27928), .B(n27929), .Z(n27922) );
  AND U27707 ( .A(n1210), .B(n27921), .Z(n27929) );
  XNOR U27708 ( .A(n27919), .B(n27928), .Z(n27921) );
  XNOR U27709 ( .A(n27930), .B(n27931), .Z(n27919) );
  AND U27710 ( .A(n1214), .B(n27932), .Z(n27931) );
  XOR U27711 ( .A(p_input[1824]), .B(n27930), .Z(n27932) );
  XNOR U27712 ( .A(n27933), .B(n27934), .Z(n27930) );
  AND U27713 ( .A(n1218), .B(n27935), .Z(n27934) );
  XOR U27714 ( .A(n27936), .B(n27937), .Z(n27928) );
  AND U27715 ( .A(n1222), .B(n27927), .Z(n27937) );
  XNOR U27716 ( .A(n27938), .B(n27925), .Z(n27927) );
  XOR U27717 ( .A(n27939), .B(n27940), .Z(n27925) );
  AND U27718 ( .A(n1245), .B(n27941), .Z(n27940) );
  IV U27719 ( .A(n27936), .Z(n27938) );
  XOR U27720 ( .A(n27942), .B(n27943), .Z(n27936) );
  AND U27721 ( .A(n1229), .B(n27935), .Z(n27943) );
  XNOR U27722 ( .A(n27933), .B(n27942), .Z(n27935) );
  XNOR U27723 ( .A(n27944), .B(n27945), .Z(n27933) );
  AND U27724 ( .A(n1233), .B(n27946), .Z(n27945) );
  XOR U27725 ( .A(p_input[1856]), .B(n27944), .Z(n27946) );
  XNOR U27726 ( .A(n27947), .B(n27948), .Z(n27944) );
  AND U27727 ( .A(n1237), .B(n27949), .Z(n27948) );
  XOR U27728 ( .A(n27950), .B(n27951), .Z(n27942) );
  AND U27729 ( .A(n1241), .B(n27941), .Z(n27951) );
  XNOR U27730 ( .A(n27952), .B(n27939), .Z(n27941) );
  XOR U27731 ( .A(n27953), .B(n27954), .Z(n27939) );
  AND U27732 ( .A(n1264), .B(n27955), .Z(n27954) );
  IV U27733 ( .A(n27950), .Z(n27952) );
  XOR U27734 ( .A(n27956), .B(n27957), .Z(n27950) );
  AND U27735 ( .A(n1248), .B(n27949), .Z(n27957) );
  XNOR U27736 ( .A(n27947), .B(n27956), .Z(n27949) );
  XNOR U27737 ( .A(n27958), .B(n27959), .Z(n27947) );
  AND U27738 ( .A(n1252), .B(n27960), .Z(n27959) );
  XOR U27739 ( .A(p_input[1888]), .B(n27958), .Z(n27960) );
  XNOR U27740 ( .A(n27961), .B(n27962), .Z(n27958) );
  AND U27741 ( .A(n1256), .B(n27963), .Z(n27962) );
  XOR U27742 ( .A(n27964), .B(n27965), .Z(n27956) );
  AND U27743 ( .A(n1260), .B(n27955), .Z(n27965) );
  XNOR U27744 ( .A(n27966), .B(n27953), .Z(n27955) );
  XOR U27745 ( .A(n27967), .B(n27968), .Z(n27953) );
  AND U27746 ( .A(n1282), .B(n27969), .Z(n27968) );
  IV U27747 ( .A(n27964), .Z(n27966) );
  XOR U27748 ( .A(n27970), .B(n27971), .Z(n27964) );
  AND U27749 ( .A(n1267), .B(n27963), .Z(n27971) );
  XNOR U27750 ( .A(n27961), .B(n27970), .Z(n27963) );
  XNOR U27751 ( .A(n27972), .B(n27973), .Z(n27961) );
  AND U27752 ( .A(n1271), .B(n27974), .Z(n27973) );
  XOR U27753 ( .A(p_input[1920]), .B(n27972), .Z(n27974) );
  XOR U27754 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(n27975), 
        .Z(n27972) );
  AND U27755 ( .A(n1274), .B(n27976), .Z(n27975) );
  XOR U27756 ( .A(n27977), .B(n27978), .Z(n27970) );
  AND U27757 ( .A(n1278), .B(n27969), .Z(n27978) );
  XNOR U27758 ( .A(n27979), .B(n27967), .Z(n27969) );
  XOR U27759 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n27980), .Z(n27967) );
  AND U27760 ( .A(n1290), .B(n27981), .Z(n27980) );
  IV U27761 ( .A(n27977), .Z(n27979) );
  XOR U27762 ( .A(n27982), .B(n27983), .Z(n27977) );
  AND U27763 ( .A(n1285), .B(n27976), .Z(n27983) );
  XOR U27764 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(n27982), 
        .Z(n27976) );
  XOR U27765 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(n27984), 
        .Z(n27982) );
  AND U27766 ( .A(n1287), .B(n27981), .Z(n27984) );
  XOR U27767 ( .A(\knn_comb_/min_val_out[0][0] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n27981) );
  XNOR U27768 ( .A(n27985), .B(n27986), .Z(n122) );
  AND U27769 ( .A(n27987), .B(n27988), .Z(n27986) );
  XNOR U27770 ( .A(n27985), .B(n27989), .Z(n27988) );
  XOR U27771 ( .A(n27990), .B(n27991), .Z(n27989) );
  AND U27772 ( .A(n125), .B(n27992), .Z(n27991) );
  XNOR U27773 ( .A(n27990), .B(n27993), .Z(n27992) );
  IV U27774 ( .A(n27994), .Z(n27990) );
  XNOR U27775 ( .A(n27985), .B(n27995), .Z(n27987) );
  XOR U27776 ( .A(n27996), .B(n27997), .Z(n27995) );
  AND U27777 ( .A(n142), .B(n27998), .Z(n27997) );
  XOR U27778 ( .A(n27999), .B(n28000), .Z(n27985) );
  AND U27779 ( .A(n28001), .B(n28002), .Z(n28000) );
  XOR U27780 ( .A(n28003), .B(n27999), .Z(n28002) );
  XNOR U27781 ( .A(n28004), .B(n28005), .Z(n28003) );
  AND U27782 ( .A(n125), .B(n28006), .Z(n28005) );
  XNOR U27783 ( .A(n28007), .B(n28004), .Z(n28006) );
  XNOR U27784 ( .A(n27999), .B(n28008), .Z(n28001) );
  XOR U27785 ( .A(n28009), .B(n28010), .Z(n28008) );
  AND U27786 ( .A(n142), .B(n28011), .Z(n28010) );
  XOR U27787 ( .A(n28012), .B(n28013), .Z(n27999) );
  AND U27788 ( .A(n28014), .B(n28015), .Z(n28013) );
  XOR U27789 ( .A(n28016), .B(n28012), .Z(n28015) );
  XNOR U27790 ( .A(n28017), .B(n28018), .Z(n28016) );
  AND U27791 ( .A(n125), .B(n28019), .Z(n28018) );
  XNOR U27792 ( .A(n28020), .B(n28017), .Z(n28019) );
  XNOR U27793 ( .A(n28012), .B(n28021), .Z(n28014) );
  XOR U27794 ( .A(n28022), .B(n28023), .Z(n28021) );
  AND U27795 ( .A(n142), .B(n28024), .Z(n28023) );
  XOR U27796 ( .A(n28025), .B(n28026), .Z(n28012) );
  AND U27797 ( .A(n28027), .B(n28028), .Z(n28026) );
  XOR U27798 ( .A(n28029), .B(n28025), .Z(n28028) );
  XNOR U27799 ( .A(n28030), .B(n28031), .Z(n28029) );
  AND U27800 ( .A(n125), .B(n28032), .Z(n28031) );
  XNOR U27801 ( .A(n28033), .B(n28030), .Z(n28032) );
  XNOR U27802 ( .A(n28025), .B(n28034), .Z(n28027) );
  XOR U27803 ( .A(n28035), .B(n28036), .Z(n28034) );
  AND U27804 ( .A(n142), .B(n28037), .Z(n28036) );
  XOR U27805 ( .A(n28038), .B(n28039), .Z(n28025) );
  AND U27806 ( .A(n28040), .B(n28041), .Z(n28039) );
  XOR U27807 ( .A(n28038), .B(n28042), .Z(n28041) );
  XOR U27808 ( .A(n28043), .B(n28044), .Z(n28042) );
  AND U27809 ( .A(n125), .B(n28045), .Z(n28044) );
  XOR U27810 ( .A(n28046), .B(n28043), .Z(n28045) );
  XNOR U27811 ( .A(n28047), .B(n28038), .Z(n28040) );
  XNOR U27812 ( .A(n28048), .B(n28049), .Z(n28047) );
  AND U27813 ( .A(n142), .B(n28050), .Z(n28049) );
  AND U27814 ( .A(n28051), .B(n28052), .Z(n28038) );
  XNOR U27815 ( .A(n28053), .B(n28054), .Z(n28052) );
  AND U27816 ( .A(n125), .B(n28055), .Z(n28054) );
  XNOR U27817 ( .A(n28056), .B(n28053), .Z(n28055) );
  XNOR U27818 ( .A(n28057), .B(n28058), .Z(n125) );
  AND U27819 ( .A(n28059), .B(n28060), .Z(n28058) );
  XOR U27820 ( .A(n27993), .B(n28057), .Z(n28060) );
  XOR U27821 ( .A(n28061), .B(n28062), .Z(n27993) );
  AND U27822 ( .A(n130), .B(n28063), .Z(n28062) );
  XOR U27823 ( .A(n28064), .B(n28061), .Z(n28063) );
  XNOR U27824 ( .A(n27994), .B(n28057), .Z(n28059) );
  XOR U27825 ( .A(n28065), .B(n28066), .Z(n27994) );
  AND U27826 ( .A(n138), .B(n27998), .Z(n28066) );
  XOR U27827 ( .A(n27996), .B(n28065), .Z(n27998) );
  XOR U27828 ( .A(n28067), .B(n28068), .Z(n28057) );
  AND U27829 ( .A(n28069), .B(n28070), .Z(n28068) );
  XOR U27830 ( .A(n28007), .B(n28067), .Z(n28070) );
  XOR U27831 ( .A(n28071), .B(n28072), .Z(n28007) );
  AND U27832 ( .A(n130), .B(n28073), .Z(n28072) );
  XOR U27833 ( .A(n28074), .B(n28071), .Z(n28073) );
  XOR U27834 ( .A(n28067), .B(n28004), .Z(n28069) );
  XOR U27835 ( .A(n28075), .B(n28076), .Z(n28004) );
  AND U27836 ( .A(n138), .B(n28011), .Z(n28076) );
  XOR U27837 ( .A(n28075), .B(n28077), .Z(n28011) );
  XOR U27838 ( .A(n28078), .B(n28079), .Z(n28067) );
  AND U27839 ( .A(n28080), .B(n28081), .Z(n28079) );
  XOR U27840 ( .A(n28020), .B(n28078), .Z(n28081) );
  XOR U27841 ( .A(n28082), .B(n28083), .Z(n28020) );
  AND U27842 ( .A(n130), .B(n28084), .Z(n28083) );
  XNOR U27843 ( .A(n28085), .B(n28082), .Z(n28084) );
  XOR U27844 ( .A(n28078), .B(n28017), .Z(n28080) );
  XOR U27845 ( .A(n28086), .B(n28087), .Z(n28017) );
  AND U27846 ( .A(n138), .B(n28024), .Z(n28087) );
  XOR U27847 ( .A(n28086), .B(n28088), .Z(n28024) );
  XOR U27848 ( .A(n28089), .B(n28090), .Z(n28078) );
  AND U27849 ( .A(n28091), .B(n28092), .Z(n28090) );
  XOR U27850 ( .A(n28033), .B(n28089), .Z(n28092) );
  XOR U27851 ( .A(n28093), .B(n28094), .Z(n28033) );
  AND U27852 ( .A(n130), .B(n28095), .Z(n28094) );
  XOR U27853 ( .A(n28096), .B(n28093), .Z(n28095) );
  XOR U27854 ( .A(n28089), .B(n28030), .Z(n28091) );
  XOR U27855 ( .A(n28097), .B(n28098), .Z(n28030) );
  AND U27856 ( .A(n138), .B(n28037), .Z(n28098) );
  XOR U27857 ( .A(n28097), .B(n28099), .Z(n28037) );
  XOR U27858 ( .A(n28100), .B(n28101), .Z(n28089) );
  AND U27859 ( .A(n28102), .B(n28103), .Z(n28101) );
  XOR U27860 ( .A(n28100), .B(n28046), .Z(n28103) );
  XOR U27861 ( .A(n28104), .B(n28105), .Z(n28046) );
  AND U27862 ( .A(n130), .B(n28106), .Z(n28105) );
  XNOR U27863 ( .A(n28107), .B(n28104), .Z(n28106) );
  XNOR U27864 ( .A(n28043), .B(n28100), .Z(n28102) );
  XNOR U27865 ( .A(n28108), .B(n28109), .Z(n28043) );
  AND U27866 ( .A(n138), .B(n28050), .Z(n28109) );
  XOR U27867 ( .A(n28108), .B(n28048), .Z(n28050) );
  AND U27868 ( .A(n28053), .B(n28056), .Z(n28100) );
  XOR U27869 ( .A(n28110), .B(n28111), .Z(n28056) );
  AND U27870 ( .A(n130), .B(n28112), .Z(n28111) );
  XNOR U27871 ( .A(n28113), .B(n28114), .Z(n28112) );
  XNOR U27872 ( .A(n28115), .B(n28116), .Z(n130) );
  AND U27873 ( .A(n28117), .B(n28118), .Z(n28116) );
  XOR U27874 ( .A(n28064), .B(n28115), .Z(n28118) );
  AND U27875 ( .A(n28119), .B(n28120), .Z(n28064) );
  XNOR U27876 ( .A(n28061), .B(n28115), .Z(n28117) );
  XNOR U27877 ( .A(n28121), .B(n28122), .Z(n28061) );
  AND U27878 ( .A(n134), .B(n28123), .Z(n28122) );
  XNOR U27879 ( .A(n28124), .B(n28125), .Z(n28123) );
  XOR U27880 ( .A(n28126), .B(n28127), .Z(n28115) );
  AND U27881 ( .A(n28128), .B(n28129), .Z(n28127) );
  XNOR U27882 ( .A(n28126), .B(n28119), .Z(n28129) );
  IV U27883 ( .A(n28074), .Z(n28119) );
  XOR U27884 ( .A(n28130), .B(n28131), .Z(n28074) );
  XOR U27885 ( .A(n28132), .B(n28120), .Z(n28131) );
  AND U27886 ( .A(n28085), .B(n28133), .Z(n28120) );
  AND U27887 ( .A(n28134), .B(n28135), .Z(n28132) );
  XOR U27888 ( .A(n28136), .B(n28130), .Z(n28134) );
  XNOR U27889 ( .A(n28071), .B(n28126), .Z(n28128) );
  XNOR U27890 ( .A(n28137), .B(n28138), .Z(n28071) );
  AND U27891 ( .A(n134), .B(n28139), .Z(n28138) );
  XNOR U27892 ( .A(n28140), .B(n28141), .Z(n28139) );
  XOR U27893 ( .A(n28142), .B(n28143), .Z(n28126) );
  AND U27894 ( .A(n28144), .B(n28145), .Z(n28143) );
  XNOR U27895 ( .A(n28142), .B(n28085), .Z(n28145) );
  XOR U27896 ( .A(n28146), .B(n28135), .Z(n28085) );
  XNOR U27897 ( .A(n28147), .B(n28130), .Z(n28135) );
  XOR U27898 ( .A(n28148), .B(n28149), .Z(n28130) );
  AND U27899 ( .A(n28150), .B(n28151), .Z(n28149) );
  XOR U27900 ( .A(n28152), .B(n28148), .Z(n28150) );
  XNOR U27901 ( .A(n28153), .B(n28154), .Z(n28147) );
  AND U27902 ( .A(n28155), .B(n28156), .Z(n28154) );
  XOR U27903 ( .A(n28153), .B(n28157), .Z(n28155) );
  XNOR U27904 ( .A(n28136), .B(n28133), .Z(n28146) );
  AND U27905 ( .A(n28158), .B(n28159), .Z(n28133) );
  XOR U27906 ( .A(n28160), .B(n28161), .Z(n28136) );
  AND U27907 ( .A(n28162), .B(n28163), .Z(n28161) );
  XOR U27908 ( .A(n28160), .B(n28164), .Z(n28162) );
  XNOR U27909 ( .A(n28082), .B(n28142), .Z(n28144) );
  XNOR U27910 ( .A(n28165), .B(n28166), .Z(n28082) );
  AND U27911 ( .A(n134), .B(n28167), .Z(n28166) );
  XNOR U27912 ( .A(n28168), .B(n28169), .Z(n28167) );
  XOR U27913 ( .A(n28170), .B(n28171), .Z(n28142) );
  AND U27914 ( .A(n28172), .B(n28173), .Z(n28171) );
  XNOR U27915 ( .A(n28170), .B(n28158), .Z(n28173) );
  IV U27916 ( .A(n28096), .Z(n28158) );
  XNOR U27917 ( .A(n28174), .B(n28151), .Z(n28096) );
  XNOR U27918 ( .A(n28175), .B(n28157), .Z(n28151) );
  XOR U27919 ( .A(n28176), .B(n28177), .Z(n28157) );
  AND U27920 ( .A(n28178), .B(n28179), .Z(n28177) );
  XOR U27921 ( .A(n28176), .B(n28180), .Z(n28178) );
  XNOR U27922 ( .A(n28156), .B(n28148), .Z(n28175) );
  XOR U27923 ( .A(n28181), .B(n28182), .Z(n28148) );
  AND U27924 ( .A(n28183), .B(n28184), .Z(n28182) );
  XNOR U27925 ( .A(n28185), .B(n28181), .Z(n28183) );
  XNOR U27926 ( .A(n28186), .B(n28153), .Z(n28156) );
  XOR U27927 ( .A(n28187), .B(n28188), .Z(n28153) );
  AND U27928 ( .A(n28189), .B(n28190), .Z(n28188) );
  XOR U27929 ( .A(n28187), .B(n28191), .Z(n28189) );
  XNOR U27930 ( .A(n28192), .B(n28193), .Z(n28186) );
  AND U27931 ( .A(n28194), .B(n28195), .Z(n28193) );
  XNOR U27932 ( .A(n28192), .B(n28196), .Z(n28194) );
  XNOR U27933 ( .A(n28152), .B(n28159), .Z(n28174) );
  AND U27934 ( .A(n28107), .B(n28197), .Z(n28159) );
  XOR U27935 ( .A(n28164), .B(n28163), .Z(n28152) );
  XNOR U27936 ( .A(n28198), .B(n28160), .Z(n28163) );
  XOR U27937 ( .A(n28199), .B(n28200), .Z(n28160) );
  AND U27938 ( .A(n28201), .B(n28202), .Z(n28200) );
  XOR U27939 ( .A(n28199), .B(n28203), .Z(n28201) );
  XNOR U27940 ( .A(n28204), .B(n28205), .Z(n28198) );
  AND U27941 ( .A(n28206), .B(n28207), .Z(n28205) );
  XOR U27942 ( .A(n28204), .B(n28208), .Z(n28206) );
  XOR U27943 ( .A(n28209), .B(n28210), .Z(n28164) );
  AND U27944 ( .A(n28211), .B(n28212), .Z(n28210) );
  XOR U27945 ( .A(n28209), .B(n28213), .Z(n28211) );
  XNOR U27946 ( .A(n28093), .B(n28170), .Z(n28172) );
  XNOR U27947 ( .A(n28214), .B(n28215), .Z(n28093) );
  AND U27948 ( .A(n134), .B(n28216), .Z(n28215) );
  XNOR U27949 ( .A(n28217), .B(n28218), .Z(n28216) );
  XOR U27950 ( .A(n28219), .B(n28220), .Z(n28170) );
  AND U27951 ( .A(n28221), .B(n28222), .Z(n28220) );
  XNOR U27952 ( .A(n28219), .B(n28107), .Z(n28222) );
  XOR U27953 ( .A(n28223), .B(n28184), .Z(n28107) );
  XNOR U27954 ( .A(n28224), .B(n28191), .Z(n28184) );
  XOR U27955 ( .A(n28180), .B(n28179), .Z(n28191) );
  XNOR U27956 ( .A(n28225), .B(n28176), .Z(n28179) );
  XOR U27957 ( .A(n28226), .B(n28227), .Z(n28176) );
  AND U27958 ( .A(n28228), .B(n28229), .Z(n28227) );
  XNOR U27959 ( .A(n28230), .B(n28231), .Z(n28228) );
  IV U27960 ( .A(n28226), .Z(n28230) );
  XNOR U27961 ( .A(n28232), .B(n28233), .Z(n28225) );
  NOR U27962 ( .A(n28234), .B(n28235), .Z(n28233) );
  XNOR U27963 ( .A(n28232), .B(n28236), .Z(n28234) );
  XOR U27964 ( .A(n28237), .B(n28238), .Z(n28180) );
  NOR U27965 ( .A(n28239), .B(n28240), .Z(n28238) );
  XNOR U27966 ( .A(n28237), .B(n28241), .Z(n28239) );
  XNOR U27967 ( .A(n28190), .B(n28181), .Z(n28224) );
  XOR U27968 ( .A(n28242), .B(n28243), .Z(n28181) );
  NOR U27969 ( .A(n28244), .B(n28245), .Z(n28243) );
  XOR U27970 ( .A(n28246), .B(n28247), .Z(n28244) );
  XOR U27971 ( .A(n28248), .B(n28196), .Z(n28190) );
  XNOR U27972 ( .A(n28249), .B(n28250), .Z(n28196) );
  NOR U27973 ( .A(n28251), .B(n28252), .Z(n28250) );
  XNOR U27974 ( .A(n28249), .B(n28253), .Z(n28251) );
  XNOR U27975 ( .A(n28195), .B(n28187), .Z(n28248) );
  XOR U27976 ( .A(n28254), .B(n28255), .Z(n28187) );
  AND U27977 ( .A(n28256), .B(n28257), .Z(n28255) );
  XOR U27978 ( .A(n28254), .B(n28258), .Z(n28256) );
  XNOR U27979 ( .A(n28259), .B(n28192), .Z(n28195) );
  XOR U27980 ( .A(n28260), .B(n28261), .Z(n28192) );
  AND U27981 ( .A(n28262), .B(n28263), .Z(n28261) );
  XOR U27982 ( .A(n28260), .B(n28264), .Z(n28262) );
  XNOR U27983 ( .A(n28265), .B(n28266), .Z(n28259) );
  NOR U27984 ( .A(n28267), .B(n28268), .Z(n28266) );
  XOR U27985 ( .A(n28265), .B(n28269), .Z(n28267) );
  XOR U27986 ( .A(n28185), .B(n28197), .Z(n28223) );
  NOR U27987 ( .A(n28113), .B(n28270), .Z(n28197) );
  XNOR U27988 ( .A(n28203), .B(n28202), .Z(n28185) );
  XNOR U27989 ( .A(n28271), .B(n28208), .Z(n28202) );
  XNOR U27990 ( .A(n28272), .B(n28273), .Z(n28208) );
  NOR U27991 ( .A(n28274), .B(n28275), .Z(n28273) );
  XOR U27992 ( .A(n28272), .B(n28276), .Z(n28274) );
  XNOR U27993 ( .A(n28207), .B(n28199), .Z(n28271) );
  XOR U27994 ( .A(n28277), .B(n28278), .Z(n28199) );
  AND U27995 ( .A(n28279), .B(n28280), .Z(n28278) );
  XNOR U27996 ( .A(n28277), .B(n28281), .Z(n28279) );
  XNOR U27997 ( .A(n28282), .B(n28204), .Z(n28207) );
  XOR U27998 ( .A(n28283), .B(n28284), .Z(n28204) );
  AND U27999 ( .A(n28285), .B(n28286), .Z(n28284) );
  XNOR U28000 ( .A(n28287), .B(n28288), .Z(n28285) );
  IV U28001 ( .A(n28283), .Z(n28287) );
  XNOR U28002 ( .A(n28289), .B(n28290), .Z(n28282) );
  NOR U28003 ( .A(n28291), .B(n28292), .Z(n28290) );
  XNOR U28004 ( .A(n28289), .B(n28293), .Z(n28291) );
  XOR U28005 ( .A(n28213), .B(n28212), .Z(n28203) );
  XNOR U28006 ( .A(n28294), .B(n28209), .Z(n28212) );
  XOR U28007 ( .A(n28295), .B(n28296), .Z(n28209) );
  AND U28008 ( .A(n28297), .B(n28298), .Z(n28296) );
  XOR U28009 ( .A(n28295), .B(n28299), .Z(n28297) );
  XNOR U28010 ( .A(n28300), .B(n28301), .Z(n28294) );
  NOR U28011 ( .A(n28302), .B(n28303), .Z(n28301) );
  XNOR U28012 ( .A(n28300), .B(n28304), .Z(n28302) );
  XOR U28013 ( .A(n28305), .B(n28306), .Z(n28213) );
  NOR U28014 ( .A(n28307), .B(n28308), .Z(n28306) );
  XNOR U28015 ( .A(n28305), .B(n28309), .Z(n28307) );
  XNOR U28016 ( .A(n28104), .B(n28219), .Z(n28221) );
  XNOR U28017 ( .A(n28310), .B(n28311), .Z(n28104) );
  AND U28018 ( .A(n134), .B(n28312), .Z(n28311) );
  XNOR U28019 ( .A(n28313), .B(n28314), .Z(n28312) );
  AND U28020 ( .A(n28114), .B(n28113), .Z(n28219) );
  XOR U28021 ( .A(n28315), .B(n28270), .Z(n28113) );
  XNOR U28022 ( .A(p_input[0]), .B(p_input[2048]), .Z(n28270) );
  XOR U28023 ( .A(n28247), .B(n28245), .Z(n28315) );
  XOR U28024 ( .A(n28316), .B(n28258), .Z(n28245) );
  XOR U28025 ( .A(n28231), .B(n28229), .Z(n28258) );
  XNOR U28026 ( .A(n28317), .B(n28236), .Z(n28229) );
  XOR U28027 ( .A(p_input[2072]), .B(p_input[24]), .Z(n28236) );
  XOR U28028 ( .A(n28226), .B(n28235), .Z(n28317) );
  XOR U28029 ( .A(n28318), .B(n28232), .Z(n28235) );
  XOR U28030 ( .A(p_input[2070]), .B(p_input[22]), .Z(n28232) );
  XNOR U28031 ( .A(p_input[2071]), .B(p_input[23]), .Z(n28318) );
  XOR U28032 ( .A(p_input[18]), .B(p_input[2066]), .Z(n28226) );
  XNOR U28033 ( .A(n28241), .B(n28240), .Z(n28231) );
  XOR U28034 ( .A(n28319), .B(n28237), .Z(n28240) );
  XOR U28035 ( .A(p_input[19]), .B(p_input[2067]), .Z(n28237) );
  XNOR U28036 ( .A(p_input[2068]), .B(p_input[20]), .Z(n28319) );
  XOR U28037 ( .A(p_input[2069]), .B(p_input[21]), .Z(n28241) );
  XOR U28038 ( .A(n28257), .B(n28246), .Z(n28316) );
  IV U28039 ( .A(n28242), .Z(n28246) );
  XOR U28040 ( .A(p_input[1]), .B(p_input[2049]), .Z(n28242) );
  XNOR U28041 ( .A(n28320), .B(n28264), .Z(n28257) );
  XNOR U28042 ( .A(n28253), .B(n28252), .Z(n28264) );
  XOR U28043 ( .A(n28321), .B(n28249), .Z(n28252) );
  XNOR U28044 ( .A(n28322), .B(p_input[26]), .Z(n28249) );
  XNOR U28045 ( .A(p_input[2075]), .B(p_input[27]), .Z(n28321) );
  XOR U28046 ( .A(p_input[2076]), .B(p_input[28]), .Z(n28253) );
  XOR U28047 ( .A(n28263), .B(n28323), .Z(n28320) );
  IV U28048 ( .A(n28254), .Z(n28323) );
  XOR U28049 ( .A(p_input[17]), .B(p_input[2065]), .Z(n28254) );
  XOR U28050 ( .A(n28324), .B(n28269), .Z(n28263) );
  XNOR U28051 ( .A(p_input[2079]), .B(p_input[31]), .Z(n28269) );
  XOR U28052 ( .A(n28260), .B(n28268), .Z(n28324) );
  XOR U28053 ( .A(n28325), .B(n28265), .Z(n28268) );
  XOR U28054 ( .A(p_input[2077]), .B(p_input[29]), .Z(n28265) );
  XNOR U28055 ( .A(p_input[2078]), .B(p_input[30]), .Z(n28325) );
  XNOR U28056 ( .A(n28326), .B(p_input[25]), .Z(n28260) );
  XNOR U28057 ( .A(n28281), .B(n28280), .Z(n28247) );
  XNOR U28058 ( .A(n28327), .B(n28288), .Z(n28280) );
  XNOR U28059 ( .A(n28276), .B(n28275), .Z(n28288) );
  XNOR U28060 ( .A(n28328), .B(n28272), .Z(n28275) );
  XNOR U28061 ( .A(p_input[11]), .B(p_input[2059]), .Z(n28272) );
  XOR U28062 ( .A(p_input[12]), .B(n28329), .Z(n28328) );
  XOR U28063 ( .A(p_input[13]), .B(p_input[2061]), .Z(n28276) );
  XNOR U28064 ( .A(n28286), .B(n28277), .Z(n28327) );
  XNOR U28065 ( .A(n28330), .B(p_input[2]), .Z(n28277) );
  XNOR U28066 ( .A(n28331), .B(n28293), .Z(n28286) );
  XNOR U28067 ( .A(p_input[16]), .B(n28332), .Z(n28293) );
  XOR U28068 ( .A(n28283), .B(n28292), .Z(n28331) );
  XOR U28069 ( .A(n28333), .B(n28289), .Z(n28292) );
  XOR U28070 ( .A(p_input[14]), .B(p_input[2062]), .Z(n28289) );
  XOR U28071 ( .A(p_input[15]), .B(n28334), .Z(n28333) );
  XOR U28072 ( .A(p_input[10]), .B(p_input[2058]), .Z(n28283) );
  XNOR U28073 ( .A(n28299), .B(n28298), .Z(n28281) );
  XNOR U28074 ( .A(n28335), .B(n28304), .Z(n28298) );
  XOR U28075 ( .A(p_input[2057]), .B(p_input[9]), .Z(n28304) );
  XOR U28076 ( .A(n28295), .B(n28303), .Z(n28335) );
  XOR U28077 ( .A(n28336), .B(n28300), .Z(n28303) );
  XOR U28078 ( .A(p_input[2055]), .B(p_input[7]), .Z(n28300) );
  XNOR U28079 ( .A(p_input[2056]), .B(p_input[8]), .Z(n28336) );
  XNOR U28080 ( .A(n28337), .B(p_input[3]), .Z(n28295) );
  XNOR U28081 ( .A(n28309), .B(n28308), .Z(n28299) );
  XOR U28082 ( .A(n28338), .B(n28305), .Z(n28308) );
  XOR U28083 ( .A(p_input[2052]), .B(p_input[4]), .Z(n28305) );
  XNOR U28084 ( .A(p_input[2053]), .B(p_input[5]), .Z(n28338) );
  XOR U28085 ( .A(p_input[2054]), .B(p_input[6]), .Z(n28309) );
  IV U28086 ( .A(n28110), .Z(n28114) );
  XOR U28087 ( .A(n28339), .B(n28340), .Z(n28110) );
  AND U28088 ( .A(n134), .B(n28341), .Z(n28340) );
  XNOR U28089 ( .A(n28342), .B(n28343), .Z(n134) );
  AND U28090 ( .A(n28344), .B(n28345), .Z(n28343) );
  XOR U28091 ( .A(n28125), .B(n28342), .Z(n28345) );
  XNOR U28092 ( .A(n28346), .B(n28342), .Z(n28344) );
  XOR U28093 ( .A(n28347), .B(n28348), .Z(n28342) );
  AND U28094 ( .A(n28349), .B(n28350), .Z(n28348) );
  XOR U28095 ( .A(n28140), .B(n28347), .Z(n28350) );
  XOR U28096 ( .A(n28347), .B(n28141), .Z(n28349) );
  XOR U28097 ( .A(n28351), .B(n28352), .Z(n28347) );
  AND U28098 ( .A(n28353), .B(n28354), .Z(n28352) );
  XOR U28099 ( .A(n28168), .B(n28351), .Z(n28354) );
  XOR U28100 ( .A(n28351), .B(n28169), .Z(n28353) );
  XOR U28101 ( .A(n28355), .B(n28356), .Z(n28351) );
  AND U28102 ( .A(n28357), .B(n28358), .Z(n28356) );
  XOR U28103 ( .A(n28217), .B(n28355), .Z(n28358) );
  XOR U28104 ( .A(n28355), .B(n28218), .Z(n28357) );
  XOR U28105 ( .A(n28359), .B(n28360), .Z(n28355) );
  AND U28106 ( .A(n28361), .B(n28362), .Z(n28360) );
  XOR U28107 ( .A(n28359), .B(n28313), .Z(n28362) );
  XNOR U28108 ( .A(n28363), .B(n28364), .Z(n28053) );
  AND U28109 ( .A(n138), .B(n28365), .Z(n28364) );
  XNOR U28110 ( .A(n28366), .B(n28367), .Z(n138) );
  AND U28111 ( .A(n28368), .B(n28369), .Z(n28367) );
  XOR U28112 ( .A(n28366), .B(n28065), .Z(n28369) );
  XNOR U28113 ( .A(n28366), .B(n27996), .Z(n28368) );
  XOR U28114 ( .A(n28370), .B(n28371), .Z(n28366) );
  AND U28115 ( .A(n28372), .B(n28373), .Z(n28371) );
  XNOR U28116 ( .A(n28075), .B(n28370), .Z(n28373) );
  XOR U28117 ( .A(n28370), .B(n28077), .Z(n28372) );
  XOR U28118 ( .A(n28374), .B(n28375), .Z(n28370) );
  AND U28119 ( .A(n28376), .B(n28377), .Z(n28375) );
  XNOR U28120 ( .A(n28086), .B(n28374), .Z(n28377) );
  XOR U28121 ( .A(n28374), .B(n28088), .Z(n28376) );
  IV U28122 ( .A(n28022), .Z(n28088) );
  XOR U28123 ( .A(n28378), .B(n28379), .Z(n28374) );
  AND U28124 ( .A(n28380), .B(n28381), .Z(n28379) );
  XOR U28125 ( .A(n28378), .B(n28099), .Z(n28380) );
  XOR U28126 ( .A(n28382), .B(n28383), .Z(n28051) );
  AND U28127 ( .A(n142), .B(n28365), .Z(n28383) );
  XNOR U28128 ( .A(n28363), .B(n28382), .Z(n28365) );
  XNOR U28129 ( .A(n28384), .B(n28385), .Z(n142) );
  AND U28130 ( .A(n28386), .B(n28387), .Z(n28385) );
  XNOR U28131 ( .A(n28388), .B(n28384), .Z(n28387) );
  IV U28132 ( .A(n28065), .Z(n28388) );
  XOR U28133 ( .A(n28346), .B(n28389), .Z(n28065) );
  AND U28134 ( .A(n146), .B(n28390), .Z(n28389) );
  XOR U28135 ( .A(n28124), .B(n28121), .Z(n28390) );
  IV U28136 ( .A(n28346), .Z(n28124) );
  XNOR U28137 ( .A(n27996), .B(n28384), .Z(n28386) );
  XOR U28138 ( .A(n28391), .B(n28392), .Z(n27996) );
  AND U28139 ( .A(n162), .B(n28393), .Z(n28392) );
  XOR U28140 ( .A(n28394), .B(n28395), .Z(n28384) );
  AND U28141 ( .A(n28396), .B(n28397), .Z(n28395) );
  XNOR U28142 ( .A(n28394), .B(n28075), .Z(n28397) );
  XOR U28143 ( .A(n28141), .B(n28398), .Z(n28075) );
  AND U28144 ( .A(n146), .B(n28399), .Z(n28398) );
  XOR U28145 ( .A(n28137), .B(n28141), .Z(n28399) );
  XNOR U28146 ( .A(n28009), .B(n28394), .Z(n28396) );
  IV U28147 ( .A(n28077), .Z(n28009) );
  XOR U28148 ( .A(n28400), .B(n28401), .Z(n28077) );
  AND U28149 ( .A(n162), .B(n28402), .Z(n28401) );
  XOR U28150 ( .A(n28403), .B(n28404), .Z(n28394) );
  AND U28151 ( .A(n28405), .B(n28406), .Z(n28404) );
  XNOR U28152 ( .A(n28403), .B(n28086), .Z(n28406) );
  XOR U28153 ( .A(n28169), .B(n28407), .Z(n28086) );
  AND U28154 ( .A(n146), .B(n28408), .Z(n28407) );
  XOR U28155 ( .A(n28165), .B(n28169), .Z(n28408) );
  XNOR U28156 ( .A(n28022), .B(n28403), .Z(n28405) );
  XNOR U28157 ( .A(n28409), .B(n28410), .Z(n28022) );
  AND U28158 ( .A(n162), .B(n28411), .Z(n28410) );
  XOR U28159 ( .A(n28378), .B(n28412), .Z(n28403) );
  AND U28160 ( .A(n28413), .B(n28381), .Z(n28412) );
  XNOR U28161 ( .A(n28097), .B(n28378), .Z(n28381) );
  XOR U28162 ( .A(n28218), .B(n28414), .Z(n28097) );
  AND U28163 ( .A(n146), .B(n28415), .Z(n28414) );
  XOR U28164 ( .A(n28214), .B(n28218), .Z(n28415) );
  XNOR U28165 ( .A(n28035), .B(n28378), .Z(n28413) );
  IV U28166 ( .A(n28099), .Z(n28035) );
  XOR U28167 ( .A(n28416), .B(n28417), .Z(n28099) );
  AND U28168 ( .A(n162), .B(n28418), .Z(n28417) );
  XOR U28169 ( .A(n28419), .B(n28420), .Z(n28378) );
  AND U28170 ( .A(n28421), .B(n28422), .Z(n28420) );
  XNOR U28171 ( .A(n28419), .B(n28108), .Z(n28422) );
  XOR U28172 ( .A(n28314), .B(n28423), .Z(n28108) );
  AND U28173 ( .A(n146), .B(n28424), .Z(n28423) );
  XOR U28174 ( .A(n28310), .B(n28314), .Z(n28424) );
  XNOR U28175 ( .A(n28425), .B(n28419), .Z(n28421) );
  IV U28176 ( .A(n28048), .Z(n28425) );
  XOR U28177 ( .A(n28426), .B(n28427), .Z(n28048) );
  AND U28178 ( .A(n162), .B(n28428), .Z(n28427) );
  AND U28179 ( .A(n28382), .B(n28363), .Z(n28419) );
  XNOR U28180 ( .A(n28429), .B(n28430), .Z(n28363) );
  AND U28181 ( .A(n146), .B(n28341), .Z(n28430) );
  XNOR U28182 ( .A(n28339), .B(n28429), .Z(n28341) );
  XNOR U28183 ( .A(n28431), .B(n28432), .Z(n146) );
  AND U28184 ( .A(n28433), .B(n28434), .Z(n28432) );
  XNOR U28185 ( .A(n28431), .B(n28121), .Z(n28434) );
  IV U28186 ( .A(n28125), .Z(n28121) );
  XOR U28187 ( .A(n28435), .B(n28436), .Z(n28125) );
  AND U28188 ( .A(n150), .B(n28437), .Z(n28436) );
  XOR U28189 ( .A(n28438), .B(n28435), .Z(n28437) );
  XNOR U28190 ( .A(n28431), .B(n28346), .Z(n28433) );
  XOR U28191 ( .A(n28439), .B(n28440), .Z(n28346) );
  AND U28192 ( .A(n158), .B(n28393), .Z(n28440) );
  XOR U28193 ( .A(n28391), .B(n28439), .Z(n28393) );
  XOR U28194 ( .A(n28441), .B(n28442), .Z(n28431) );
  AND U28195 ( .A(n28443), .B(n28444), .Z(n28442) );
  XNOR U28196 ( .A(n28441), .B(n28137), .Z(n28444) );
  IV U28197 ( .A(n28140), .Z(n28137) );
  XOR U28198 ( .A(n28445), .B(n28446), .Z(n28140) );
  AND U28199 ( .A(n150), .B(n28447), .Z(n28446) );
  XOR U28200 ( .A(n28448), .B(n28445), .Z(n28447) );
  XOR U28201 ( .A(n28141), .B(n28441), .Z(n28443) );
  XOR U28202 ( .A(n28449), .B(n28450), .Z(n28141) );
  AND U28203 ( .A(n158), .B(n28402), .Z(n28450) );
  XOR U28204 ( .A(n28449), .B(n28400), .Z(n28402) );
  XOR U28205 ( .A(n28451), .B(n28452), .Z(n28441) );
  AND U28206 ( .A(n28453), .B(n28454), .Z(n28452) );
  XNOR U28207 ( .A(n28451), .B(n28165), .Z(n28454) );
  IV U28208 ( .A(n28168), .Z(n28165) );
  XOR U28209 ( .A(n28455), .B(n28456), .Z(n28168) );
  AND U28210 ( .A(n150), .B(n28457), .Z(n28456) );
  XNOR U28211 ( .A(n28458), .B(n28455), .Z(n28457) );
  XOR U28212 ( .A(n28169), .B(n28451), .Z(n28453) );
  XOR U28213 ( .A(n28459), .B(n28460), .Z(n28169) );
  AND U28214 ( .A(n158), .B(n28411), .Z(n28460) );
  XOR U28215 ( .A(n28459), .B(n28409), .Z(n28411) );
  XOR U28216 ( .A(n28461), .B(n28462), .Z(n28451) );
  AND U28217 ( .A(n28463), .B(n28464), .Z(n28462) );
  XNOR U28218 ( .A(n28461), .B(n28214), .Z(n28464) );
  IV U28219 ( .A(n28217), .Z(n28214) );
  XOR U28220 ( .A(n28465), .B(n28466), .Z(n28217) );
  AND U28221 ( .A(n150), .B(n28467), .Z(n28466) );
  XOR U28222 ( .A(n28468), .B(n28465), .Z(n28467) );
  XOR U28223 ( .A(n28218), .B(n28461), .Z(n28463) );
  XOR U28224 ( .A(n28469), .B(n28470), .Z(n28218) );
  AND U28225 ( .A(n158), .B(n28418), .Z(n28470) );
  XOR U28226 ( .A(n28469), .B(n28416), .Z(n28418) );
  XOR U28227 ( .A(n28359), .B(n28471), .Z(n28461) );
  AND U28228 ( .A(n28361), .B(n28472), .Z(n28471) );
  XNOR U28229 ( .A(n28359), .B(n28310), .Z(n28472) );
  IV U28230 ( .A(n28313), .Z(n28310) );
  XOR U28231 ( .A(n28473), .B(n28474), .Z(n28313) );
  AND U28232 ( .A(n150), .B(n28475), .Z(n28474) );
  XNOR U28233 ( .A(n28476), .B(n28473), .Z(n28475) );
  XOR U28234 ( .A(n28314), .B(n28359), .Z(n28361) );
  XOR U28235 ( .A(n28477), .B(n28478), .Z(n28314) );
  AND U28236 ( .A(n158), .B(n28428), .Z(n28478) );
  XOR U28237 ( .A(n28477), .B(n28426), .Z(n28428) );
  AND U28238 ( .A(n28429), .B(n28339), .Z(n28359) );
  XNOR U28239 ( .A(n28479), .B(n28480), .Z(n28339) );
  AND U28240 ( .A(n150), .B(n28481), .Z(n28480) );
  XNOR U28241 ( .A(n28482), .B(n28479), .Z(n28481) );
  XNOR U28242 ( .A(n28483), .B(n28484), .Z(n150) );
  AND U28243 ( .A(n28485), .B(n28486), .Z(n28484) );
  XOR U28244 ( .A(n28438), .B(n28483), .Z(n28486) );
  AND U28245 ( .A(n28487), .B(n28488), .Z(n28438) );
  XNOR U28246 ( .A(n28435), .B(n28483), .Z(n28485) );
  XNOR U28247 ( .A(n28489), .B(n28490), .Z(n28435) );
  AND U28248 ( .A(n154), .B(n28491), .Z(n28490) );
  XNOR U28249 ( .A(n28492), .B(n28493), .Z(n28491) );
  XOR U28250 ( .A(n28494), .B(n28495), .Z(n28483) );
  AND U28251 ( .A(n28496), .B(n28497), .Z(n28495) );
  XNOR U28252 ( .A(n28494), .B(n28487), .Z(n28497) );
  IV U28253 ( .A(n28448), .Z(n28487) );
  XOR U28254 ( .A(n28498), .B(n28499), .Z(n28448) );
  XOR U28255 ( .A(n28500), .B(n28488), .Z(n28499) );
  AND U28256 ( .A(n28458), .B(n28501), .Z(n28488) );
  AND U28257 ( .A(n28502), .B(n28503), .Z(n28500) );
  XOR U28258 ( .A(n28504), .B(n28498), .Z(n28502) );
  XNOR U28259 ( .A(n28445), .B(n28494), .Z(n28496) );
  XNOR U28260 ( .A(n28505), .B(n28506), .Z(n28445) );
  AND U28261 ( .A(n154), .B(n28507), .Z(n28506) );
  XNOR U28262 ( .A(n28508), .B(n28509), .Z(n28507) );
  XOR U28263 ( .A(n28510), .B(n28511), .Z(n28494) );
  AND U28264 ( .A(n28512), .B(n28513), .Z(n28511) );
  XNOR U28265 ( .A(n28510), .B(n28458), .Z(n28513) );
  XOR U28266 ( .A(n28514), .B(n28503), .Z(n28458) );
  XNOR U28267 ( .A(n28515), .B(n28498), .Z(n28503) );
  XOR U28268 ( .A(n28516), .B(n28517), .Z(n28498) );
  AND U28269 ( .A(n28518), .B(n28519), .Z(n28517) );
  XOR U28270 ( .A(n28520), .B(n28516), .Z(n28518) );
  XNOR U28271 ( .A(n28521), .B(n28522), .Z(n28515) );
  AND U28272 ( .A(n28523), .B(n28524), .Z(n28522) );
  XOR U28273 ( .A(n28521), .B(n28525), .Z(n28523) );
  XNOR U28274 ( .A(n28504), .B(n28501), .Z(n28514) );
  AND U28275 ( .A(n28526), .B(n28527), .Z(n28501) );
  XOR U28276 ( .A(n28528), .B(n28529), .Z(n28504) );
  AND U28277 ( .A(n28530), .B(n28531), .Z(n28529) );
  XOR U28278 ( .A(n28528), .B(n28532), .Z(n28530) );
  XNOR U28279 ( .A(n28455), .B(n28510), .Z(n28512) );
  XNOR U28280 ( .A(n28533), .B(n28534), .Z(n28455) );
  AND U28281 ( .A(n154), .B(n28535), .Z(n28534) );
  XNOR U28282 ( .A(n28536), .B(n28537), .Z(n28535) );
  XOR U28283 ( .A(n28538), .B(n28539), .Z(n28510) );
  AND U28284 ( .A(n28540), .B(n28541), .Z(n28539) );
  XNOR U28285 ( .A(n28538), .B(n28526), .Z(n28541) );
  IV U28286 ( .A(n28468), .Z(n28526) );
  XNOR U28287 ( .A(n28542), .B(n28519), .Z(n28468) );
  XNOR U28288 ( .A(n28543), .B(n28525), .Z(n28519) );
  XOR U28289 ( .A(n28544), .B(n28545), .Z(n28525) );
  AND U28290 ( .A(n28546), .B(n28547), .Z(n28545) );
  XOR U28291 ( .A(n28544), .B(n28548), .Z(n28546) );
  XNOR U28292 ( .A(n28524), .B(n28516), .Z(n28543) );
  XOR U28293 ( .A(n28549), .B(n28550), .Z(n28516) );
  AND U28294 ( .A(n28551), .B(n28552), .Z(n28550) );
  XNOR U28295 ( .A(n28553), .B(n28549), .Z(n28551) );
  XNOR U28296 ( .A(n28554), .B(n28521), .Z(n28524) );
  XOR U28297 ( .A(n28555), .B(n28556), .Z(n28521) );
  AND U28298 ( .A(n28557), .B(n28558), .Z(n28556) );
  XOR U28299 ( .A(n28555), .B(n28559), .Z(n28557) );
  XNOR U28300 ( .A(n28560), .B(n28561), .Z(n28554) );
  AND U28301 ( .A(n28562), .B(n28563), .Z(n28561) );
  XNOR U28302 ( .A(n28560), .B(n28564), .Z(n28562) );
  XNOR U28303 ( .A(n28520), .B(n28527), .Z(n28542) );
  AND U28304 ( .A(n28476), .B(n28565), .Z(n28527) );
  XOR U28305 ( .A(n28532), .B(n28531), .Z(n28520) );
  XNOR U28306 ( .A(n28566), .B(n28528), .Z(n28531) );
  XOR U28307 ( .A(n28567), .B(n28568), .Z(n28528) );
  AND U28308 ( .A(n28569), .B(n28570), .Z(n28568) );
  XOR U28309 ( .A(n28567), .B(n28571), .Z(n28569) );
  XNOR U28310 ( .A(n28572), .B(n28573), .Z(n28566) );
  AND U28311 ( .A(n28574), .B(n28575), .Z(n28573) );
  XOR U28312 ( .A(n28572), .B(n28576), .Z(n28574) );
  XOR U28313 ( .A(n28577), .B(n28578), .Z(n28532) );
  AND U28314 ( .A(n28579), .B(n28580), .Z(n28578) );
  XOR U28315 ( .A(n28577), .B(n28581), .Z(n28579) );
  XNOR U28316 ( .A(n28465), .B(n28538), .Z(n28540) );
  XNOR U28317 ( .A(n28582), .B(n28583), .Z(n28465) );
  AND U28318 ( .A(n154), .B(n28584), .Z(n28583) );
  XNOR U28319 ( .A(n28585), .B(n28586), .Z(n28584) );
  XOR U28320 ( .A(n28587), .B(n28588), .Z(n28538) );
  AND U28321 ( .A(n28589), .B(n28590), .Z(n28588) );
  XNOR U28322 ( .A(n28587), .B(n28476), .Z(n28590) );
  XOR U28323 ( .A(n28591), .B(n28552), .Z(n28476) );
  XNOR U28324 ( .A(n28592), .B(n28559), .Z(n28552) );
  XOR U28325 ( .A(n28548), .B(n28547), .Z(n28559) );
  XNOR U28326 ( .A(n28593), .B(n28544), .Z(n28547) );
  XOR U28327 ( .A(n28594), .B(n28595), .Z(n28544) );
  AND U28328 ( .A(n28596), .B(n28597), .Z(n28595) );
  XOR U28329 ( .A(n28594), .B(n28598), .Z(n28596) );
  XNOR U28330 ( .A(n28599), .B(n28600), .Z(n28593) );
  NOR U28331 ( .A(n28601), .B(n28602), .Z(n28600) );
  XNOR U28332 ( .A(n28599), .B(n28603), .Z(n28601) );
  XOR U28333 ( .A(n28604), .B(n28605), .Z(n28548) );
  NOR U28334 ( .A(n28606), .B(n28607), .Z(n28605) );
  XNOR U28335 ( .A(n28604), .B(n28608), .Z(n28606) );
  XNOR U28336 ( .A(n28558), .B(n28549), .Z(n28592) );
  XOR U28337 ( .A(n28609), .B(n28610), .Z(n28549) );
  NOR U28338 ( .A(n28611), .B(n28612), .Z(n28610) );
  XNOR U28339 ( .A(n28609), .B(n28613), .Z(n28611) );
  XOR U28340 ( .A(n28614), .B(n28564), .Z(n28558) );
  XNOR U28341 ( .A(n28615), .B(n28616), .Z(n28564) );
  NOR U28342 ( .A(n28617), .B(n28618), .Z(n28616) );
  XNOR U28343 ( .A(n28615), .B(n28619), .Z(n28617) );
  XNOR U28344 ( .A(n28563), .B(n28555), .Z(n28614) );
  XOR U28345 ( .A(n28620), .B(n28621), .Z(n28555) );
  AND U28346 ( .A(n28622), .B(n28623), .Z(n28621) );
  XOR U28347 ( .A(n28620), .B(n28624), .Z(n28622) );
  XNOR U28348 ( .A(n28625), .B(n28560), .Z(n28563) );
  XOR U28349 ( .A(n28626), .B(n28627), .Z(n28560) );
  AND U28350 ( .A(n28628), .B(n28629), .Z(n28627) );
  XOR U28351 ( .A(n28626), .B(n28630), .Z(n28628) );
  XNOR U28352 ( .A(n28631), .B(n28632), .Z(n28625) );
  NOR U28353 ( .A(n28633), .B(n28634), .Z(n28632) );
  XOR U28354 ( .A(n28631), .B(n28635), .Z(n28633) );
  XOR U28355 ( .A(n28553), .B(n28565), .Z(n28591) );
  NOR U28356 ( .A(n28482), .B(n28636), .Z(n28565) );
  XNOR U28357 ( .A(n28571), .B(n28570), .Z(n28553) );
  XNOR U28358 ( .A(n28637), .B(n28576), .Z(n28570) );
  XOR U28359 ( .A(n28638), .B(n28639), .Z(n28576) );
  NOR U28360 ( .A(n28640), .B(n28641), .Z(n28639) );
  XNOR U28361 ( .A(n28638), .B(n28642), .Z(n28640) );
  XNOR U28362 ( .A(n28575), .B(n28567), .Z(n28637) );
  XOR U28363 ( .A(n28643), .B(n28644), .Z(n28567) );
  AND U28364 ( .A(n28645), .B(n28646), .Z(n28644) );
  XNOR U28365 ( .A(n28643), .B(n28647), .Z(n28645) );
  XNOR U28366 ( .A(n28648), .B(n28572), .Z(n28575) );
  XOR U28367 ( .A(n28649), .B(n28650), .Z(n28572) );
  AND U28368 ( .A(n28651), .B(n28652), .Z(n28650) );
  XOR U28369 ( .A(n28649), .B(n28653), .Z(n28651) );
  XNOR U28370 ( .A(n28654), .B(n28655), .Z(n28648) );
  NOR U28371 ( .A(n28656), .B(n28657), .Z(n28655) );
  XOR U28372 ( .A(n28654), .B(n28658), .Z(n28656) );
  XOR U28373 ( .A(n28581), .B(n28580), .Z(n28571) );
  XNOR U28374 ( .A(n28659), .B(n28577), .Z(n28580) );
  XOR U28375 ( .A(n28660), .B(n28661), .Z(n28577) );
  AND U28376 ( .A(n28662), .B(n28663), .Z(n28661) );
  XOR U28377 ( .A(n28660), .B(n28664), .Z(n28662) );
  XNOR U28378 ( .A(n28665), .B(n28666), .Z(n28659) );
  NOR U28379 ( .A(n28667), .B(n28668), .Z(n28666) );
  XNOR U28380 ( .A(n28665), .B(n28669), .Z(n28667) );
  XOR U28381 ( .A(n28670), .B(n28671), .Z(n28581) );
  NOR U28382 ( .A(n28672), .B(n28673), .Z(n28671) );
  XNOR U28383 ( .A(n28670), .B(n28674), .Z(n28672) );
  XNOR U28384 ( .A(n28473), .B(n28587), .Z(n28589) );
  XNOR U28385 ( .A(n28675), .B(n28676), .Z(n28473) );
  AND U28386 ( .A(n154), .B(n28677), .Z(n28676) );
  XNOR U28387 ( .A(n28678), .B(n28679), .Z(n28677) );
  AND U28388 ( .A(n28479), .B(n28482), .Z(n28587) );
  XOR U28389 ( .A(n28680), .B(n28636), .Z(n28482) );
  XNOR U28390 ( .A(p_input[2048]), .B(p_input[32]), .Z(n28636) );
  XOR U28391 ( .A(n28613), .B(n28612), .Z(n28680) );
  XOR U28392 ( .A(n28681), .B(n28624), .Z(n28612) );
  XOR U28393 ( .A(n28598), .B(n28597), .Z(n28624) );
  XNOR U28394 ( .A(n28682), .B(n28603), .Z(n28597) );
  XOR U28395 ( .A(p_input[2072]), .B(p_input[56]), .Z(n28603) );
  XOR U28396 ( .A(n28594), .B(n28602), .Z(n28682) );
  XOR U28397 ( .A(n28683), .B(n28599), .Z(n28602) );
  XOR U28398 ( .A(p_input[2070]), .B(p_input[54]), .Z(n28599) );
  XNOR U28399 ( .A(p_input[2071]), .B(p_input[55]), .Z(n28683) );
  XNOR U28400 ( .A(n28684), .B(p_input[50]), .Z(n28594) );
  XNOR U28401 ( .A(n28608), .B(n28607), .Z(n28598) );
  XOR U28402 ( .A(n28685), .B(n28604), .Z(n28607) );
  XOR U28403 ( .A(p_input[2067]), .B(p_input[51]), .Z(n28604) );
  XNOR U28404 ( .A(p_input[2068]), .B(p_input[52]), .Z(n28685) );
  XOR U28405 ( .A(p_input[2069]), .B(p_input[53]), .Z(n28608) );
  XNOR U28406 ( .A(n28623), .B(n28609), .Z(n28681) );
  XNOR U28407 ( .A(n28686), .B(p_input[33]), .Z(n28609) );
  XNOR U28408 ( .A(n28687), .B(n28630), .Z(n28623) );
  XNOR U28409 ( .A(n28619), .B(n28618), .Z(n28630) );
  XOR U28410 ( .A(n28688), .B(n28615), .Z(n28618) );
  XNOR U28411 ( .A(n28322), .B(p_input[58]), .Z(n28615) );
  XNOR U28412 ( .A(p_input[2075]), .B(p_input[59]), .Z(n28688) );
  XOR U28413 ( .A(p_input[2076]), .B(p_input[60]), .Z(n28619) );
  XNOR U28414 ( .A(n28629), .B(n28620), .Z(n28687) );
  XNOR U28415 ( .A(n28689), .B(p_input[49]), .Z(n28620) );
  XOR U28416 ( .A(n28690), .B(n28635), .Z(n28629) );
  XNOR U28417 ( .A(p_input[2079]), .B(p_input[63]), .Z(n28635) );
  XOR U28418 ( .A(n28626), .B(n28634), .Z(n28690) );
  XOR U28419 ( .A(n28691), .B(n28631), .Z(n28634) );
  XOR U28420 ( .A(p_input[2077]), .B(p_input[61]), .Z(n28631) );
  XNOR U28421 ( .A(p_input[2078]), .B(p_input[62]), .Z(n28691) );
  XNOR U28422 ( .A(n28326), .B(p_input[57]), .Z(n28626) );
  XNOR U28423 ( .A(n28647), .B(n28646), .Z(n28613) );
  XNOR U28424 ( .A(n28692), .B(n28653), .Z(n28646) );
  XNOR U28425 ( .A(n28642), .B(n28641), .Z(n28653) );
  XOR U28426 ( .A(n28693), .B(n28638), .Z(n28641) );
  XNOR U28427 ( .A(n28694), .B(p_input[43]), .Z(n28638) );
  XNOR U28428 ( .A(p_input[2060]), .B(p_input[44]), .Z(n28693) );
  XOR U28429 ( .A(p_input[2061]), .B(p_input[45]), .Z(n28642) );
  XNOR U28430 ( .A(n28652), .B(n28643), .Z(n28692) );
  XNOR U28431 ( .A(n28330), .B(p_input[34]), .Z(n28643) );
  XOR U28432 ( .A(n28695), .B(n28658), .Z(n28652) );
  XNOR U28433 ( .A(p_input[2064]), .B(p_input[48]), .Z(n28658) );
  XOR U28434 ( .A(n28649), .B(n28657), .Z(n28695) );
  XOR U28435 ( .A(n28696), .B(n28654), .Z(n28657) );
  XOR U28436 ( .A(p_input[2062]), .B(p_input[46]), .Z(n28654) );
  XNOR U28437 ( .A(p_input[2063]), .B(p_input[47]), .Z(n28696) );
  XNOR U28438 ( .A(n28697), .B(p_input[42]), .Z(n28649) );
  XNOR U28439 ( .A(n28664), .B(n28663), .Z(n28647) );
  XNOR U28440 ( .A(n28698), .B(n28669), .Z(n28663) );
  XOR U28441 ( .A(p_input[2057]), .B(p_input[41]), .Z(n28669) );
  XOR U28442 ( .A(n28660), .B(n28668), .Z(n28698) );
  XOR U28443 ( .A(n28699), .B(n28665), .Z(n28668) );
  XOR U28444 ( .A(p_input[2055]), .B(p_input[39]), .Z(n28665) );
  XNOR U28445 ( .A(p_input[2056]), .B(p_input[40]), .Z(n28699) );
  XNOR U28446 ( .A(n28337), .B(p_input[35]), .Z(n28660) );
  XNOR U28447 ( .A(n28674), .B(n28673), .Z(n28664) );
  XOR U28448 ( .A(n28700), .B(n28670), .Z(n28673) );
  XOR U28449 ( .A(p_input[2052]), .B(p_input[36]), .Z(n28670) );
  XNOR U28450 ( .A(p_input[2053]), .B(p_input[37]), .Z(n28700) );
  XOR U28451 ( .A(p_input[2054]), .B(p_input[38]), .Z(n28674) );
  XNOR U28452 ( .A(n28701), .B(n28702), .Z(n28479) );
  AND U28453 ( .A(n154), .B(n28703), .Z(n28702) );
  XNOR U28454 ( .A(n28704), .B(n28705), .Z(n154) );
  AND U28455 ( .A(n28706), .B(n28707), .Z(n28705) );
  XOR U28456 ( .A(n28493), .B(n28704), .Z(n28707) );
  XNOR U28457 ( .A(n28708), .B(n28704), .Z(n28706) );
  XOR U28458 ( .A(n28709), .B(n28710), .Z(n28704) );
  AND U28459 ( .A(n28711), .B(n28712), .Z(n28710) );
  XOR U28460 ( .A(n28508), .B(n28709), .Z(n28712) );
  XOR U28461 ( .A(n28709), .B(n28509), .Z(n28711) );
  XOR U28462 ( .A(n28713), .B(n28714), .Z(n28709) );
  AND U28463 ( .A(n28715), .B(n28716), .Z(n28714) );
  XOR U28464 ( .A(n28536), .B(n28713), .Z(n28716) );
  XOR U28465 ( .A(n28713), .B(n28537), .Z(n28715) );
  XOR U28466 ( .A(n28717), .B(n28718), .Z(n28713) );
  AND U28467 ( .A(n28719), .B(n28720), .Z(n28718) );
  XOR U28468 ( .A(n28585), .B(n28717), .Z(n28720) );
  XOR U28469 ( .A(n28717), .B(n28586), .Z(n28719) );
  XOR U28470 ( .A(n28721), .B(n28722), .Z(n28717) );
  AND U28471 ( .A(n28723), .B(n28724), .Z(n28722) );
  XOR U28472 ( .A(n28721), .B(n28678), .Z(n28724) );
  XNOR U28473 ( .A(n28725), .B(n28726), .Z(n28429) );
  AND U28474 ( .A(n158), .B(n28727), .Z(n28726) );
  XNOR U28475 ( .A(n28728), .B(n28729), .Z(n158) );
  AND U28476 ( .A(n28730), .B(n28731), .Z(n28729) );
  XOR U28477 ( .A(n28728), .B(n28439), .Z(n28731) );
  XNOR U28478 ( .A(n28728), .B(n28391), .Z(n28730) );
  XOR U28479 ( .A(n28732), .B(n28733), .Z(n28728) );
  AND U28480 ( .A(n28734), .B(n28735), .Z(n28733) );
  XNOR U28481 ( .A(n28449), .B(n28732), .Z(n28735) );
  XOR U28482 ( .A(n28732), .B(n28400), .Z(n28734) );
  XOR U28483 ( .A(n28736), .B(n28737), .Z(n28732) );
  AND U28484 ( .A(n28738), .B(n28739), .Z(n28737) );
  XNOR U28485 ( .A(n28459), .B(n28736), .Z(n28739) );
  XOR U28486 ( .A(n28736), .B(n28409), .Z(n28738) );
  XOR U28487 ( .A(n28740), .B(n28741), .Z(n28736) );
  AND U28488 ( .A(n28742), .B(n28743), .Z(n28741) );
  XOR U28489 ( .A(n28740), .B(n28416), .Z(n28742) );
  XOR U28490 ( .A(n28744), .B(n28745), .Z(n28382) );
  AND U28491 ( .A(n162), .B(n28727), .Z(n28745) );
  XNOR U28492 ( .A(n28725), .B(n28744), .Z(n28727) );
  XNOR U28493 ( .A(n28746), .B(n28747), .Z(n162) );
  AND U28494 ( .A(n28748), .B(n28749), .Z(n28747) );
  XNOR U28495 ( .A(n28750), .B(n28746), .Z(n28749) );
  IV U28496 ( .A(n28439), .Z(n28750) );
  XOR U28497 ( .A(n28708), .B(n28751), .Z(n28439) );
  AND U28498 ( .A(n165), .B(n28752), .Z(n28751) );
  XOR U28499 ( .A(n28492), .B(n28489), .Z(n28752) );
  IV U28500 ( .A(n28708), .Z(n28492) );
  XNOR U28501 ( .A(n28391), .B(n28746), .Z(n28748) );
  XOR U28502 ( .A(n28753), .B(n28754), .Z(n28391) );
  AND U28503 ( .A(n181), .B(n28755), .Z(n28754) );
  XOR U28504 ( .A(n28756), .B(n28757), .Z(n28746) );
  AND U28505 ( .A(n28758), .B(n28759), .Z(n28757) );
  XNOR U28506 ( .A(n28756), .B(n28449), .Z(n28759) );
  XOR U28507 ( .A(n28509), .B(n28760), .Z(n28449) );
  AND U28508 ( .A(n165), .B(n28761), .Z(n28760) );
  XOR U28509 ( .A(n28505), .B(n28509), .Z(n28761) );
  XNOR U28510 ( .A(n28762), .B(n28756), .Z(n28758) );
  IV U28511 ( .A(n28400), .Z(n28762) );
  XOR U28512 ( .A(n28763), .B(n28764), .Z(n28400) );
  AND U28513 ( .A(n181), .B(n28765), .Z(n28764) );
  XOR U28514 ( .A(n28766), .B(n28767), .Z(n28756) );
  AND U28515 ( .A(n28768), .B(n28769), .Z(n28767) );
  XNOR U28516 ( .A(n28766), .B(n28459), .Z(n28769) );
  XOR U28517 ( .A(n28537), .B(n28770), .Z(n28459) );
  AND U28518 ( .A(n165), .B(n28771), .Z(n28770) );
  XOR U28519 ( .A(n28533), .B(n28537), .Z(n28771) );
  XOR U28520 ( .A(n28409), .B(n28766), .Z(n28768) );
  XOR U28521 ( .A(n28772), .B(n28773), .Z(n28409) );
  AND U28522 ( .A(n181), .B(n28774), .Z(n28773) );
  XOR U28523 ( .A(n28740), .B(n28775), .Z(n28766) );
  AND U28524 ( .A(n28776), .B(n28743), .Z(n28775) );
  XNOR U28525 ( .A(n28469), .B(n28740), .Z(n28743) );
  XOR U28526 ( .A(n28586), .B(n28777), .Z(n28469) );
  AND U28527 ( .A(n165), .B(n28778), .Z(n28777) );
  XOR U28528 ( .A(n28582), .B(n28586), .Z(n28778) );
  XNOR U28529 ( .A(n28779), .B(n28740), .Z(n28776) );
  IV U28530 ( .A(n28416), .Z(n28779) );
  XOR U28531 ( .A(n28780), .B(n28781), .Z(n28416) );
  AND U28532 ( .A(n181), .B(n28782), .Z(n28781) );
  XOR U28533 ( .A(n28783), .B(n28784), .Z(n28740) );
  AND U28534 ( .A(n28785), .B(n28786), .Z(n28784) );
  XNOR U28535 ( .A(n28783), .B(n28477), .Z(n28786) );
  XOR U28536 ( .A(n28679), .B(n28787), .Z(n28477) );
  AND U28537 ( .A(n165), .B(n28788), .Z(n28787) );
  XOR U28538 ( .A(n28675), .B(n28679), .Z(n28788) );
  XNOR U28539 ( .A(n28789), .B(n28783), .Z(n28785) );
  IV U28540 ( .A(n28426), .Z(n28789) );
  XOR U28541 ( .A(n28790), .B(n28791), .Z(n28426) );
  AND U28542 ( .A(n181), .B(n28792), .Z(n28791) );
  AND U28543 ( .A(n28744), .B(n28725), .Z(n28783) );
  XNOR U28544 ( .A(n28793), .B(n28794), .Z(n28725) );
  AND U28545 ( .A(n165), .B(n28703), .Z(n28794) );
  XNOR U28546 ( .A(n28701), .B(n28793), .Z(n28703) );
  XNOR U28547 ( .A(n28795), .B(n28796), .Z(n165) );
  AND U28548 ( .A(n28797), .B(n28798), .Z(n28796) );
  XNOR U28549 ( .A(n28795), .B(n28489), .Z(n28798) );
  IV U28550 ( .A(n28493), .Z(n28489) );
  XOR U28551 ( .A(n28799), .B(n28800), .Z(n28493) );
  AND U28552 ( .A(n169), .B(n28801), .Z(n28800) );
  XOR U28553 ( .A(n28802), .B(n28799), .Z(n28801) );
  XNOR U28554 ( .A(n28795), .B(n28708), .Z(n28797) );
  XOR U28555 ( .A(n28803), .B(n28804), .Z(n28708) );
  AND U28556 ( .A(n177), .B(n28755), .Z(n28804) );
  XOR U28557 ( .A(n28753), .B(n28803), .Z(n28755) );
  XOR U28558 ( .A(n28805), .B(n28806), .Z(n28795) );
  AND U28559 ( .A(n28807), .B(n28808), .Z(n28806) );
  XNOR U28560 ( .A(n28805), .B(n28505), .Z(n28808) );
  IV U28561 ( .A(n28508), .Z(n28505) );
  XOR U28562 ( .A(n28809), .B(n28810), .Z(n28508) );
  AND U28563 ( .A(n169), .B(n28811), .Z(n28810) );
  XOR U28564 ( .A(n28812), .B(n28809), .Z(n28811) );
  XOR U28565 ( .A(n28509), .B(n28805), .Z(n28807) );
  XOR U28566 ( .A(n28813), .B(n28814), .Z(n28509) );
  AND U28567 ( .A(n177), .B(n28765), .Z(n28814) );
  XOR U28568 ( .A(n28813), .B(n28763), .Z(n28765) );
  XOR U28569 ( .A(n28815), .B(n28816), .Z(n28805) );
  AND U28570 ( .A(n28817), .B(n28818), .Z(n28816) );
  XNOR U28571 ( .A(n28815), .B(n28533), .Z(n28818) );
  IV U28572 ( .A(n28536), .Z(n28533) );
  XOR U28573 ( .A(n28819), .B(n28820), .Z(n28536) );
  AND U28574 ( .A(n169), .B(n28821), .Z(n28820) );
  XNOR U28575 ( .A(n28822), .B(n28819), .Z(n28821) );
  XOR U28576 ( .A(n28537), .B(n28815), .Z(n28817) );
  XOR U28577 ( .A(n28823), .B(n28824), .Z(n28537) );
  AND U28578 ( .A(n177), .B(n28774), .Z(n28824) );
  XOR U28579 ( .A(n28823), .B(n28772), .Z(n28774) );
  XOR U28580 ( .A(n28825), .B(n28826), .Z(n28815) );
  AND U28581 ( .A(n28827), .B(n28828), .Z(n28826) );
  XNOR U28582 ( .A(n28825), .B(n28582), .Z(n28828) );
  IV U28583 ( .A(n28585), .Z(n28582) );
  XOR U28584 ( .A(n28829), .B(n28830), .Z(n28585) );
  AND U28585 ( .A(n169), .B(n28831), .Z(n28830) );
  XOR U28586 ( .A(n28832), .B(n28829), .Z(n28831) );
  XOR U28587 ( .A(n28586), .B(n28825), .Z(n28827) );
  XOR U28588 ( .A(n28833), .B(n28834), .Z(n28586) );
  AND U28589 ( .A(n177), .B(n28782), .Z(n28834) );
  XOR U28590 ( .A(n28833), .B(n28780), .Z(n28782) );
  XOR U28591 ( .A(n28721), .B(n28835), .Z(n28825) );
  AND U28592 ( .A(n28723), .B(n28836), .Z(n28835) );
  XNOR U28593 ( .A(n28721), .B(n28675), .Z(n28836) );
  IV U28594 ( .A(n28678), .Z(n28675) );
  XOR U28595 ( .A(n28837), .B(n28838), .Z(n28678) );
  AND U28596 ( .A(n169), .B(n28839), .Z(n28838) );
  XNOR U28597 ( .A(n28840), .B(n28837), .Z(n28839) );
  XOR U28598 ( .A(n28679), .B(n28721), .Z(n28723) );
  XOR U28599 ( .A(n28841), .B(n28842), .Z(n28679) );
  AND U28600 ( .A(n177), .B(n28792), .Z(n28842) );
  XOR U28601 ( .A(n28841), .B(n28790), .Z(n28792) );
  AND U28602 ( .A(n28793), .B(n28701), .Z(n28721) );
  XNOR U28603 ( .A(n28843), .B(n28844), .Z(n28701) );
  AND U28604 ( .A(n169), .B(n28845), .Z(n28844) );
  XNOR U28605 ( .A(n28846), .B(n28843), .Z(n28845) );
  XNOR U28606 ( .A(n28847), .B(n28848), .Z(n169) );
  AND U28607 ( .A(n28849), .B(n28850), .Z(n28848) );
  XOR U28608 ( .A(n28802), .B(n28847), .Z(n28850) );
  AND U28609 ( .A(n28851), .B(n28852), .Z(n28802) );
  XNOR U28610 ( .A(n28799), .B(n28847), .Z(n28849) );
  XNOR U28611 ( .A(n28853), .B(n28854), .Z(n28799) );
  AND U28612 ( .A(n173), .B(n28855), .Z(n28854) );
  XNOR U28613 ( .A(n28856), .B(n28857), .Z(n28855) );
  XOR U28614 ( .A(n28858), .B(n28859), .Z(n28847) );
  AND U28615 ( .A(n28860), .B(n28861), .Z(n28859) );
  XNOR U28616 ( .A(n28858), .B(n28851), .Z(n28861) );
  IV U28617 ( .A(n28812), .Z(n28851) );
  XOR U28618 ( .A(n28862), .B(n28863), .Z(n28812) );
  XOR U28619 ( .A(n28864), .B(n28852), .Z(n28863) );
  AND U28620 ( .A(n28822), .B(n28865), .Z(n28852) );
  AND U28621 ( .A(n28866), .B(n28867), .Z(n28864) );
  XOR U28622 ( .A(n28868), .B(n28862), .Z(n28866) );
  XNOR U28623 ( .A(n28809), .B(n28858), .Z(n28860) );
  XNOR U28624 ( .A(n28869), .B(n28870), .Z(n28809) );
  AND U28625 ( .A(n173), .B(n28871), .Z(n28870) );
  XNOR U28626 ( .A(n28872), .B(n28873), .Z(n28871) );
  XOR U28627 ( .A(n28874), .B(n28875), .Z(n28858) );
  AND U28628 ( .A(n28876), .B(n28877), .Z(n28875) );
  XNOR U28629 ( .A(n28874), .B(n28822), .Z(n28877) );
  XOR U28630 ( .A(n28878), .B(n28867), .Z(n28822) );
  XNOR U28631 ( .A(n28879), .B(n28862), .Z(n28867) );
  XOR U28632 ( .A(n28880), .B(n28881), .Z(n28862) );
  AND U28633 ( .A(n28882), .B(n28883), .Z(n28881) );
  XOR U28634 ( .A(n28884), .B(n28880), .Z(n28882) );
  XNOR U28635 ( .A(n28885), .B(n28886), .Z(n28879) );
  AND U28636 ( .A(n28887), .B(n28888), .Z(n28886) );
  XOR U28637 ( .A(n28885), .B(n28889), .Z(n28887) );
  XNOR U28638 ( .A(n28868), .B(n28865), .Z(n28878) );
  AND U28639 ( .A(n28890), .B(n28891), .Z(n28865) );
  XOR U28640 ( .A(n28892), .B(n28893), .Z(n28868) );
  AND U28641 ( .A(n28894), .B(n28895), .Z(n28893) );
  XOR U28642 ( .A(n28892), .B(n28896), .Z(n28894) );
  XNOR U28643 ( .A(n28819), .B(n28874), .Z(n28876) );
  XNOR U28644 ( .A(n28897), .B(n28898), .Z(n28819) );
  AND U28645 ( .A(n173), .B(n28899), .Z(n28898) );
  XNOR U28646 ( .A(n28900), .B(n28901), .Z(n28899) );
  XOR U28647 ( .A(n28902), .B(n28903), .Z(n28874) );
  AND U28648 ( .A(n28904), .B(n28905), .Z(n28903) );
  XNOR U28649 ( .A(n28902), .B(n28890), .Z(n28905) );
  IV U28650 ( .A(n28832), .Z(n28890) );
  XNOR U28651 ( .A(n28906), .B(n28883), .Z(n28832) );
  XNOR U28652 ( .A(n28907), .B(n28889), .Z(n28883) );
  XOR U28653 ( .A(n28908), .B(n28909), .Z(n28889) );
  AND U28654 ( .A(n28910), .B(n28911), .Z(n28909) );
  XOR U28655 ( .A(n28908), .B(n28912), .Z(n28910) );
  XNOR U28656 ( .A(n28888), .B(n28880), .Z(n28907) );
  XOR U28657 ( .A(n28913), .B(n28914), .Z(n28880) );
  AND U28658 ( .A(n28915), .B(n28916), .Z(n28914) );
  XNOR U28659 ( .A(n28917), .B(n28913), .Z(n28915) );
  XNOR U28660 ( .A(n28918), .B(n28885), .Z(n28888) );
  XOR U28661 ( .A(n28919), .B(n28920), .Z(n28885) );
  AND U28662 ( .A(n28921), .B(n28922), .Z(n28920) );
  XOR U28663 ( .A(n28919), .B(n28923), .Z(n28921) );
  XNOR U28664 ( .A(n28924), .B(n28925), .Z(n28918) );
  AND U28665 ( .A(n28926), .B(n28927), .Z(n28925) );
  XNOR U28666 ( .A(n28924), .B(n28928), .Z(n28926) );
  XNOR U28667 ( .A(n28884), .B(n28891), .Z(n28906) );
  AND U28668 ( .A(n28840), .B(n28929), .Z(n28891) );
  XOR U28669 ( .A(n28896), .B(n28895), .Z(n28884) );
  XNOR U28670 ( .A(n28930), .B(n28892), .Z(n28895) );
  XOR U28671 ( .A(n28931), .B(n28932), .Z(n28892) );
  AND U28672 ( .A(n28933), .B(n28934), .Z(n28932) );
  XOR U28673 ( .A(n28931), .B(n28935), .Z(n28933) );
  XNOR U28674 ( .A(n28936), .B(n28937), .Z(n28930) );
  AND U28675 ( .A(n28938), .B(n28939), .Z(n28937) );
  XOR U28676 ( .A(n28936), .B(n28940), .Z(n28938) );
  XOR U28677 ( .A(n28941), .B(n28942), .Z(n28896) );
  AND U28678 ( .A(n28943), .B(n28944), .Z(n28942) );
  XOR U28679 ( .A(n28941), .B(n28945), .Z(n28943) );
  XNOR U28680 ( .A(n28829), .B(n28902), .Z(n28904) );
  XNOR U28681 ( .A(n28946), .B(n28947), .Z(n28829) );
  AND U28682 ( .A(n173), .B(n28948), .Z(n28947) );
  XNOR U28683 ( .A(n28949), .B(n28950), .Z(n28948) );
  XOR U28684 ( .A(n28951), .B(n28952), .Z(n28902) );
  AND U28685 ( .A(n28953), .B(n28954), .Z(n28952) );
  XNOR U28686 ( .A(n28951), .B(n28840), .Z(n28954) );
  XOR U28687 ( .A(n28955), .B(n28916), .Z(n28840) );
  XNOR U28688 ( .A(n28956), .B(n28923), .Z(n28916) );
  XOR U28689 ( .A(n28912), .B(n28911), .Z(n28923) );
  XNOR U28690 ( .A(n28957), .B(n28908), .Z(n28911) );
  XOR U28691 ( .A(n28958), .B(n28959), .Z(n28908) );
  AND U28692 ( .A(n28960), .B(n28961), .Z(n28959) );
  XOR U28693 ( .A(n28958), .B(n28962), .Z(n28960) );
  XNOR U28694 ( .A(n28963), .B(n28964), .Z(n28957) );
  NOR U28695 ( .A(n28965), .B(n28966), .Z(n28964) );
  XNOR U28696 ( .A(n28963), .B(n28967), .Z(n28965) );
  XOR U28697 ( .A(n28968), .B(n28969), .Z(n28912) );
  NOR U28698 ( .A(n28970), .B(n28971), .Z(n28969) );
  XNOR U28699 ( .A(n28968), .B(n28972), .Z(n28970) );
  XNOR U28700 ( .A(n28922), .B(n28913), .Z(n28956) );
  XOR U28701 ( .A(n28973), .B(n28974), .Z(n28913) );
  NOR U28702 ( .A(n28975), .B(n28976), .Z(n28974) );
  XNOR U28703 ( .A(n28973), .B(n28977), .Z(n28975) );
  XOR U28704 ( .A(n28978), .B(n28928), .Z(n28922) );
  XNOR U28705 ( .A(n28979), .B(n28980), .Z(n28928) );
  NOR U28706 ( .A(n28981), .B(n28982), .Z(n28980) );
  XNOR U28707 ( .A(n28979), .B(n28983), .Z(n28981) );
  XNOR U28708 ( .A(n28927), .B(n28919), .Z(n28978) );
  XOR U28709 ( .A(n28984), .B(n28985), .Z(n28919) );
  AND U28710 ( .A(n28986), .B(n28987), .Z(n28985) );
  XOR U28711 ( .A(n28984), .B(n28988), .Z(n28986) );
  XNOR U28712 ( .A(n28989), .B(n28924), .Z(n28927) );
  XOR U28713 ( .A(n28990), .B(n28991), .Z(n28924) );
  AND U28714 ( .A(n28992), .B(n28993), .Z(n28991) );
  XOR U28715 ( .A(n28990), .B(n28994), .Z(n28992) );
  XNOR U28716 ( .A(n28995), .B(n28996), .Z(n28989) );
  NOR U28717 ( .A(n28997), .B(n28998), .Z(n28996) );
  XOR U28718 ( .A(n28995), .B(n28999), .Z(n28997) );
  XOR U28719 ( .A(n28917), .B(n28929), .Z(n28955) );
  NOR U28720 ( .A(n28846), .B(n29000), .Z(n28929) );
  XNOR U28721 ( .A(n28935), .B(n28934), .Z(n28917) );
  XNOR U28722 ( .A(n29001), .B(n28940), .Z(n28934) );
  XOR U28723 ( .A(n29002), .B(n29003), .Z(n28940) );
  NOR U28724 ( .A(n29004), .B(n29005), .Z(n29003) );
  XNOR U28725 ( .A(n29002), .B(n29006), .Z(n29004) );
  XNOR U28726 ( .A(n28939), .B(n28931), .Z(n29001) );
  XOR U28727 ( .A(n29007), .B(n29008), .Z(n28931) );
  AND U28728 ( .A(n29009), .B(n29010), .Z(n29008) );
  XNOR U28729 ( .A(n29007), .B(n29011), .Z(n29009) );
  XNOR U28730 ( .A(n29012), .B(n28936), .Z(n28939) );
  XOR U28731 ( .A(n29013), .B(n29014), .Z(n28936) );
  AND U28732 ( .A(n29015), .B(n29016), .Z(n29014) );
  XOR U28733 ( .A(n29013), .B(n29017), .Z(n29015) );
  XNOR U28734 ( .A(n29018), .B(n29019), .Z(n29012) );
  NOR U28735 ( .A(n29020), .B(n29021), .Z(n29019) );
  XOR U28736 ( .A(n29018), .B(n29022), .Z(n29020) );
  XOR U28737 ( .A(n28945), .B(n28944), .Z(n28935) );
  XNOR U28738 ( .A(n29023), .B(n28941), .Z(n28944) );
  XOR U28739 ( .A(n29024), .B(n29025), .Z(n28941) );
  AND U28740 ( .A(n29026), .B(n29027), .Z(n29025) );
  XOR U28741 ( .A(n29024), .B(n29028), .Z(n29026) );
  XNOR U28742 ( .A(n29029), .B(n29030), .Z(n29023) );
  NOR U28743 ( .A(n29031), .B(n29032), .Z(n29030) );
  XNOR U28744 ( .A(n29029), .B(n29033), .Z(n29031) );
  XOR U28745 ( .A(n29034), .B(n29035), .Z(n28945) );
  NOR U28746 ( .A(n29036), .B(n29037), .Z(n29035) );
  XNOR U28747 ( .A(n29034), .B(n29038), .Z(n29036) );
  XNOR U28748 ( .A(n28837), .B(n28951), .Z(n28953) );
  XNOR U28749 ( .A(n29039), .B(n29040), .Z(n28837) );
  AND U28750 ( .A(n173), .B(n29041), .Z(n29040) );
  XNOR U28751 ( .A(n29042), .B(n29043), .Z(n29041) );
  AND U28752 ( .A(n28843), .B(n28846), .Z(n28951) );
  XOR U28753 ( .A(n29044), .B(n29000), .Z(n28846) );
  XNOR U28754 ( .A(p_input[2048]), .B(p_input[64]), .Z(n29000) );
  XOR U28755 ( .A(n28977), .B(n28976), .Z(n29044) );
  XOR U28756 ( .A(n29045), .B(n28988), .Z(n28976) );
  XOR U28757 ( .A(n28962), .B(n28961), .Z(n28988) );
  XNOR U28758 ( .A(n29046), .B(n28967), .Z(n28961) );
  XOR U28759 ( .A(p_input[2072]), .B(p_input[88]), .Z(n28967) );
  XOR U28760 ( .A(n28958), .B(n28966), .Z(n29046) );
  XOR U28761 ( .A(n29047), .B(n28963), .Z(n28966) );
  XOR U28762 ( .A(p_input[2070]), .B(p_input[86]), .Z(n28963) );
  XNOR U28763 ( .A(p_input[2071]), .B(p_input[87]), .Z(n29047) );
  XNOR U28764 ( .A(n28684), .B(p_input[82]), .Z(n28958) );
  XNOR U28765 ( .A(n28972), .B(n28971), .Z(n28962) );
  XOR U28766 ( .A(n29048), .B(n28968), .Z(n28971) );
  XOR U28767 ( .A(p_input[2067]), .B(p_input[83]), .Z(n28968) );
  XNOR U28768 ( .A(p_input[2068]), .B(p_input[84]), .Z(n29048) );
  XOR U28769 ( .A(p_input[2069]), .B(p_input[85]), .Z(n28972) );
  XNOR U28770 ( .A(n28987), .B(n28973), .Z(n29045) );
  XNOR U28771 ( .A(n28686), .B(p_input[65]), .Z(n28973) );
  XNOR U28772 ( .A(n29049), .B(n28994), .Z(n28987) );
  XNOR U28773 ( .A(n28983), .B(n28982), .Z(n28994) );
  XOR U28774 ( .A(n29050), .B(n28979), .Z(n28982) );
  XNOR U28775 ( .A(n28322), .B(p_input[90]), .Z(n28979) );
  XNOR U28776 ( .A(p_input[2075]), .B(p_input[91]), .Z(n29050) );
  XOR U28777 ( .A(p_input[2076]), .B(p_input[92]), .Z(n28983) );
  XNOR U28778 ( .A(n28993), .B(n28984), .Z(n29049) );
  XNOR U28779 ( .A(n28689), .B(p_input[81]), .Z(n28984) );
  XOR U28780 ( .A(n29051), .B(n28999), .Z(n28993) );
  XNOR U28781 ( .A(p_input[2079]), .B(p_input[95]), .Z(n28999) );
  XOR U28782 ( .A(n28990), .B(n28998), .Z(n29051) );
  XOR U28783 ( .A(n29052), .B(n28995), .Z(n28998) );
  XOR U28784 ( .A(p_input[2077]), .B(p_input[93]), .Z(n28995) );
  XNOR U28785 ( .A(p_input[2078]), .B(p_input[94]), .Z(n29052) );
  XNOR U28786 ( .A(n28326), .B(p_input[89]), .Z(n28990) );
  XNOR U28787 ( .A(n29011), .B(n29010), .Z(n28977) );
  XNOR U28788 ( .A(n29053), .B(n29017), .Z(n29010) );
  XNOR U28789 ( .A(n29006), .B(n29005), .Z(n29017) );
  XOR U28790 ( .A(n29054), .B(n29002), .Z(n29005) );
  XNOR U28791 ( .A(n28694), .B(p_input[75]), .Z(n29002) );
  XNOR U28792 ( .A(p_input[2060]), .B(p_input[76]), .Z(n29054) );
  XOR U28793 ( .A(p_input[2061]), .B(p_input[77]), .Z(n29006) );
  XNOR U28794 ( .A(n29016), .B(n29007), .Z(n29053) );
  XNOR U28795 ( .A(n28330), .B(p_input[66]), .Z(n29007) );
  XOR U28796 ( .A(n29055), .B(n29022), .Z(n29016) );
  XNOR U28797 ( .A(p_input[2064]), .B(p_input[80]), .Z(n29022) );
  XOR U28798 ( .A(n29013), .B(n29021), .Z(n29055) );
  XOR U28799 ( .A(n29056), .B(n29018), .Z(n29021) );
  XOR U28800 ( .A(p_input[2062]), .B(p_input[78]), .Z(n29018) );
  XNOR U28801 ( .A(p_input[2063]), .B(p_input[79]), .Z(n29056) );
  XNOR U28802 ( .A(n28697), .B(p_input[74]), .Z(n29013) );
  XNOR U28803 ( .A(n29028), .B(n29027), .Z(n29011) );
  XNOR U28804 ( .A(n29057), .B(n29033), .Z(n29027) );
  XOR U28805 ( .A(p_input[2057]), .B(p_input[73]), .Z(n29033) );
  XOR U28806 ( .A(n29024), .B(n29032), .Z(n29057) );
  XOR U28807 ( .A(n29058), .B(n29029), .Z(n29032) );
  XOR U28808 ( .A(p_input[2055]), .B(p_input[71]), .Z(n29029) );
  XNOR U28809 ( .A(p_input[2056]), .B(p_input[72]), .Z(n29058) );
  XNOR U28810 ( .A(n28337), .B(p_input[67]), .Z(n29024) );
  XNOR U28811 ( .A(n29038), .B(n29037), .Z(n29028) );
  XOR U28812 ( .A(n29059), .B(n29034), .Z(n29037) );
  XOR U28813 ( .A(p_input[2052]), .B(p_input[68]), .Z(n29034) );
  XNOR U28814 ( .A(p_input[2053]), .B(p_input[69]), .Z(n29059) );
  XOR U28815 ( .A(p_input[2054]), .B(p_input[70]), .Z(n29038) );
  XNOR U28816 ( .A(n29060), .B(n29061), .Z(n28843) );
  AND U28817 ( .A(n173), .B(n29062), .Z(n29061) );
  XNOR U28818 ( .A(n29063), .B(n29064), .Z(n173) );
  AND U28819 ( .A(n29065), .B(n29066), .Z(n29064) );
  XOR U28820 ( .A(n28857), .B(n29063), .Z(n29066) );
  XNOR U28821 ( .A(n29067), .B(n29063), .Z(n29065) );
  XOR U28822 ( .A(n29068), .B(n29069), .Z(n29063) );
  AND U28823 ( .A(n29070), .B(n29071), .Z(n29069) );
  XOR U28824 ( .A(n28872), .B(n29068), .Z(n29071) );
  XOR U28825 ( .A(n29068), .B(n28873), .Z(n29070) );
  XOR U28826 ( .A(n29072), .B(n29073), .Z(n29068) );
  AND U28827 ( .A(n29074), .B(n29075), .Z(n29073) );
  XOR U28828 ( .A(n28900), .B(n29072), .Z(n29075) );
  XOR U28829 ( .A(n29072), .B(n28901), .Z(n29074) );
  XOR U28830 ( .A(n29076), .B(n29077), .Z(n29072) );
  AND U28831 ( .A(n29078), .B(n29079), .Z(n29077) );
  XOR U28832 ( .A(n28949), .B(n29076), .Z(n29079) );
  XOR U28833 ( .A(n29076), .B(n28950), .Z(n29078) );
  XOR U28834 ( .A(n29080), .B(n29081), .Z(n29076) );
  AND U28835 ( .A(n29082), .B(n29083), .Z(n29081) );
  XOR U28836 ( .A(n29080), .B(n29042), .Z(n29083) );
  XNOR U28837 ( .A(n29084), .B(n29085), .Z(n28793) );
  AND U28838 ( .A(n177), .B(n29086), .Z(n29085) );
  XNOR U28839 ( .A(n29087), .B(n29088), .Z(n177) );
  AND U28840 ( .A(n29089), .B(n29090), .Z(n29088) );
  XOR U28841 ( .A(n29087), .B(n28803), .Z(n29090) );
  XNOR U28842 ( .A(n29087), .B(n28753), .Z(n29089) );
  XOR U28843 ( .A(n29091), .B(n29092), .Z(n29087) );
  AND U28844 ( .A(n29093), .B(n29094), .Z(n29092) );
  XNOR U28845 ( .A(n28813), .B(n29091), .Z(n29094) );
  XOR U28846 ( .A(n29091), .B(n28763), .Z(n29093) );
  XOR U28847 ( .A(n29095), .B(n29096), .Z(n29091) );
  AND U28848 ( .A(n29097), .B(n29098), .Z(n29096) );
  XNOR U28849 ( .A(n28823), .B(n29095), .Z(n29098) );
  XOR U28850 ( .A(n29095), .B(n28772), .Z(n29097) );
  XOR U28851 ( .A(n29099), .B(n29100), .Z(n29095) );
  AND U28852 ( .A(n29101), .B(n29102), .Z(n29100) );
  XOR U28853 ( .A(n29099), .B(n28780), .Z(n29101) );
  XOR U28854 ( .A(n29103), .B(n29104), .Z(n28744) );
  AND U28855 ( .A(n181), .B(n29086), .Z(n29104) );
  XNOR U28856 ( .A(n29084), .B(n29103), .Z(n29086) );
  XNOR U28857 ( .A(n29105), .B(n29106), .Z(n181) );
  AND U28858 ( .A(n29107), .B(n29108), .Z(n29106) );
  XNOR U28859 ( .A(n29109), .B(n29105), .Z(n29108) );
  IV U28860 ( .A(n28803), .Z(n29109) );
  XOR U28861 ( .A(n29067), .B(n29110), .Z(n28803) );
  AND U28862 ( .A(n184), .B(n29111), .Z(n29110) );
  XOR U28863 ( .A(n28856), .B(n28853), .Z(n29111) );
  IV U28864 ( .A(n29067), .Z(n28856) );
  XNOR U28865 ( .A(n28753), .B(n29105), .Z(n29107) );
  XOR U28866 ( .A(n29112), .B(n29113), .Z(n28753) );
  AND U28867 ( .A(n200), .B(n29114), .Z(n29113) );
  XOR U28868 ( .A(n29115), .B(n29116), .Z(n29105) );
  AND U28869 ( .A(n29117), .B(n29118), .Z(n29116) );
  XNOR U28870 ( .A(n29115), .B(n28813), .Z(n29118) );
  XOR U28871 ( .A(n28873), .B(n29119), .Z(n28813) );
  AND U28872 ( .A(n184), .B(n29120), .Z(n29119) );
  XOR U28873 ( .A(n28869), .B(n28873), .Z(n29120) );
  XNOR U28874 ( .A(n29121), .B(n29115), .Z(n29117) );
  IV U28875 ( .A(n28763), .Z(n29121) );
  XOR U28876 ( .A(n29122), .B(n29123), .Z(n28763) );
  AND U28877 ( .A(n200), .B(n29124), .Z(n29123) );
  XOR U28878 ( .A(n29125), .B(n29126), .Z(n29115) );
  AND U28879 ( .A(n29127), .B(n29128), .Z(n29126) );
  XNOR U28880 ( .A(n29125), .B(n28823), .Z(n29128) );
  XOR U28881 ( .A(n28901), .B(n29129), .Z(n28823) );
  AND U28882 ( .A(n184), .B(n29130), .Z(n29129) );
  XOR U28883 ( .A(n28897), .B(n28901), .Z(n29130) );
  XOR U28884 ( .A(n28772), .B(n29125), .Z(n29127) );
  XOR U28885 ( .A(n29131), .B(n29132), .Z(n28772) );
  AND U28886 ( .A(n200), .B(n29133), .Z(n29132) );
  XOR U28887 ( .A(n29099), .B(n29134), .Z(n29125) );
  AND U28888 ( .A(n29135), .B(n29102), .Z(n29134) );
  XNOR U28889 ( .A(n28833), .B(n29099), .Z(n29102) );
  XOR U28890 ( .A(n28950), .B(n29136), .Z(n28833) );
  AND U28891 ( .A(n184), .B(n29137), .Z(n29136) );
  XOR U28892 ( .A(n28946), .B(n28950), .Z(n29137) );
  XNOR U28893 ( .A(n29138), .B(n29099), .Z(n29135) );
  IV U28894 ( .A(n28780), .Z(n29138) );
  XOR U28895 ( .A(n29139), .B(n29140), .Z(n28780) );
  AND U28896 ( .A(n200), .B(n29141), .Z(n29140) );
  XOR U28897 ( .A(n29142), .B(n29143), .Z(n29099) );
  AND U28898 ( .A(n29144), .B(n29145), .Z(n29143) );
  XNOR U28899 ( .A(n29142), .B(n28841), .Z(n29145) );
  XOR U28900 ( .A(n29043), .B(n29146), .Z(n28841) );
  AND U28901 ( .A(n184), .B(n29147), .Z(n29146) );
  XOR U28902 ( .A(n29039), .B(n29043), .Z(n29147) );
  XNOR U28903 ( .A(n29148), .B(n29142), .Z(n29144) );
  IV U28904 ( .A(n28790), .Z(n29148) );
  XOR U28905 ( .A(n29149), .B(n29150), .Z(n28790) );
  AND U28906 ( .A(n200), .B(n29151), .Z(n29150) );
  AND U28907 ( .A(n29103), .B(n29084), .Z(n29142) );
  XNOR U28908 ( .A(n29152), .B(n29153), .Z(n29084) );
  AND U28909 ( .A(n184), .B(n29062), .Z(n29153) );
  XNOR U28910 ( .A(n29060), .B(n29152), .Z(n29062) );
  XNOR U28911 ( .A(n29154), .B(n29155), .Z(n184) );
  AND U28912 ( .A(n29156), .B(n29157), .Z(n29155) );
  XNOR U28913 ( .A(n29154), .B(n28853), .Z(n29157) );
  IV U28914 ( .A(n28857), .Z(n28853) );
  XOR U28915 ( .A(n29158), .B(n29159), .Z(n28857) );
  AND U28916 ( .A(n188), .B(n29160), .Z(n29159) );
  XOR U28917 ( .A(n29161), .B(n29158), .Z(n29160) );
  XNOR U28918 ( .A(n29154), .B(n29067), .Z(n29156) );
  XOR U28919 ( .A(n29162), .B(n29163), .Z(n29067) );
  AND U28920 ( .A(n196), .B(n29114), .Z(n29163) );
  XOR U28921 ( .A(n29112), .B(n29162), .Z(n29114) );
  XOR U28922 ( .A(n29164), .B(n29165), .Z(n29154) );
  AND U28923 ( .A(n29166), .B(n29167), .Z(n29165) );
  XNOR U28924 ( .A(n29164), .B(n28869), .Z(n29167) );
  IV U28925 ( .A(n28872), .Z(n28869) );
  XOR U28926 ( .A(n29168), .B(n29169), .Z(n28872) );
  AND U28927 ( .A(n188), .B(n29170), .Z(n29169) );
  XOR U28928 ( .A(n29171), .B(n29168), .Z(n29170) );
  XOR U28929 ( .A(n28873), .B(n29164), .Z(n29166) );
  XOR U28930 ( .A(n29172), .B(n29173), .Z(n28873) );
  AND U28931 ( .A(n196), .B(n29124), .Z(n29173) );
  XOR U28932 ( .A(n29172), .B(n29122), .Z(n29124) );
  XOR U28933 ( .A(n29174), .B(n29175), .Z(n29164) );
  AND U28934 ( .A(n29176), .B(n29177), .Z(n29175) );
  XNOR U28935 ( .A(n29174), .B(n28897), .Z(n29177) );
  IV U28936 ( .A(n28900), .Z(n28897) );
  XOR U28937 ( .A(n29178), .B(n29179), .Z(n28900) );
  AND U28938 ( .A(n188), .B(n29180), .Z(n29179) );
  XNOR U28939 ( .A(n29181), .B(n29178), .Z(n29180) );
  XOR U28940 ( .A(n28901), .B(n29174), .Z(n29176) );
  XOR U28941 ( .A(n29182), .B(n29183), .Z(n28901) );
  AND U28942 ( .A(n196), .B(n29133), .Z(n29183) );
  XOR U28943 ( .A(n29182), .B(n29131), .Z(n29133) );
  XOR U28944 ( .A(n29184), .B(n29185), .Z(n29174) );
  AND U28945 ( .A(n29186), .B(n29187), .Z(n29185) );
  XNOR U28946 ( .A(n29184), .B(n28946), .Z(n29187) );
  IV U28947 ( .A(n28949), .Z(n28946) );
  XOR U28948 ( .A(n29188), .B(n29189), .Z(n28949) );
  AND U28949 ( .A(n188), .B(n29190), .Z(n29189) );
  XOR U28950 ( .A(n29191), .B(n29188), .Z(n29190) );
  XOR U28951 ( .A(n28950), .B(n29184), .Z(n29186) );
  XOR U28952 ( .A(n29192), .B(n29193), .Z(n28950) );
  AND U28953 ( .A(n196), .B(n29141), .Z(n29193) );
  XOR U28954 ( .A(n29192), .B(n29139), .Z(n29141) );
  XOR U28955 ( .A(n29080), .B(n29194), .Z(n29184) );
  AND U28956 ( .A(n29082), .B(n29195), .Z(n29194) );
  XNOR U28957 ( .A(n29080), .B(n29039), .Z(n29195) );
  IV U28958 ( .A(n29042), .Z(n29039) );
  XOR U28959 ( .A(n29196), .B(n29197), .Z(n29042) );
  AND U28960 ( .A(n188), .B(n29198), .Z(n29197) );
  XNOR U28961 ( .A(n29199), .B(n29196), .Z(n29198) );
  XOR U28962 ( .A(n29043), .B(n29080), .Z(n29082) );
  XOR U28963 ( .A(n29200), .B(n29201), .Z(n29043) );
  AND U28964 ( .A(n196), .B(n29151), .Z(n29201) );
  XOR U28965 ( .A(n29200), .B(n29149), .Z(n29151) );
  AND U28966 ( .A(n29152), .B(n29060), .Z(n29080) );
  XNOR U28967 ( .A(n29202), .B(n29203), .Z(n29060) );
  AND U28968 ( .A(n188), .B(n29204), .Z(n29203) );
  XNOR U28969 ( .A(n29205), .B(n29202), .Z(n29204) );
  XNOR U28970 ( .A(n29206), .B(n29207), .Z(n188) );
  AND U28971 ( .A(n29208), .B(n29209), .Z(n29207) );
  XOR U28972 ( .A(n29161), .B(n29206), .Z(n29209) );
  AND U28973 ( .A(n29210), .B(n29211), .Z(n29161) );
  XNOR U28974 ( .A(n29158), .B(n29206), .Z(n29208) );
  XNOR U28975 ( .A(n29212), .B(n29213), .Z(n29158) );
  AND U28976 ( .A(n192), .B(n29214), .Z(n29213) );
  XNOR U28977 ( .A(n29215), .B(n29216), .Z(n29214) );
  XOR U28978 ( .A(n29217), .B(n29218), .Z(n29206) );
  AND U28979 ( .A(n29219), .B(n29220), .Z(n29218) );
  XNOR U28980 ( .A(n29217), .B(n29210), .Z(n29220) );
  IV U28981 ( .A(n29171), .Z(n29210) );
  XOR U28982 ( .A(n29221), .B(n29222), .Z(n29171) );
  XOR U28983 ( .A(n29223), .B(n29211), .Z(n29222) );
  AND U28984 ( .A(n29181), .B(n29224), .Z(n29211) );
  AND U28985 ( .A(n29225), .B(n29226), .Z(n29223) );
  XOR U28986 ( .A(n29227), .B(n29221), .Z(n29225) );
  XNOR U28987 ( .A(n29168), .B(n29217), .Z(n29219) );
  XNOR U28988 ( .A(n29228), .B(n29229), .Z(n29168) );
  AND U28989 ( .A(n192), .B(n29230), .Z(n29229) );
  XNOR U28990 ( .A(n29231), .B(n29232), .Z(n29230) );
  XOR U28991 ( .A(n29233), .B(n29234), .Z(n29217) );
  AND U28992 ( .A(n29235), .B(n29236), .Z(n29234) );
  XNOR U28993 ( .A(n29233), .B(n29181), .Z(n29236) );
  XOR U28994 ( .A(n29237), .B(n29226), .Z(n29181) );
  XNOR U28995 ( .A(n29238), .B(n29221), .Z(n29226) );
  XOR U28996 ( .A(n29239), .B(n29240), .Z(n29221) );
  AND U28997 ( .A(n29241), .B(n29242), .Z(n29240) );
  XOR U28998 ( .A(n29243), .B(n29239), .Z(n29241) );
  XNOR U28999 ( .A(n29244), .B(n29245), .Z(n29238) );
  AND U29000 ( .A(n29246), .B(n29247), .Z(n29245) );
  XOR U29001 ( .A(n29244), .B(n29248), .Z(n29246) );
  XNOR U29002 ( .A(n29227), .B(n29224), .Z(n29237) );
  AND U29003 ( .A(n29249), .B(n29250), .Z(n29224) );
  XOR U29004 ( .A(n29251), .B(n29252), .Z(n29227) );
  AND U29005 ( .A(n29253), .B(n29254), .Z(n29252) );
  XOR U29006 ( .A(n29251), .B(n29255), .Z(n29253) );
  XNOR U29007 ( .A(n29178), .B(n29233), .Z(n29235) );
  XNOR U29008 ( .A(n29256), .B(n29257), .Z(n29178) );
  AND U29009 ( .A(n192), .B(n29258), .Z(n29257) );
  XNOR U29010 ( .A(n29259), .B(n29260), .Z(n29258) );
  XOR U29011 ( .A(n29261), .B(n29262), .Z(n29233) );
  AND U29012 ( .A(n29263), .B(n29264), .Z(n29262) );
  XNOR U29013 ( .A(n29261), .B(n29249), .Z(n29264) );
  IV U29014 ( .A(n29191), .Z(n29249) );
  XNOR U29015 ( .A(n29265), .B(n29242), .Z(n29191) );
  XNOR U29016 ( .A(n29266), .B(n29248), .Z(n29242) );
  XOR U29017 ( .A(n29267), .B(n29268), .Z(n29248) );
  AND U29018 ( .A(n29269), .B(n29270), .Z(n29268) );
  XOR U29019 ( .A(n29267), .B(n29271), .Z(n29269) );
  XNOR U29020 ( .A(n29247), .B(n29239), .Z(n29266) );
  XOR U29021 ( .A(n29272), .B(n29273), .Z(n29239) );
  AND U29022 ( .A(n29274), .B(n29275), .Z(n29273) );
  XNOR U29023 ( .A(n29276), .B(n29272), .Z(n29274) );
  XNOR U29024 ( .A(n29277), .B(n29244), .Z(n29247) );
  XOR U29025 ( .A(n29278), .B(n29279), .Z(n29244) );
  AND U29026 ( .A(n29280), .B(n29281), .Z(n29279) );
  XOR U29027 ( .A(n29278), .B(n29282), .Z(n29280) );
  XNOR U29028 ( .A(n29283), .B(n29284), .Z(n29277) );
  AND U29029 ( .A(n29285), .B(n29286), .Z(n29284) );
  XNOR U29030 ( .A(n29283), .B(n29287), .Z(n29285) );
  XNOR U29031 ( .A(n29243), .B(n29250), .Z(n29265) );
  AND U29032 ( .A(n29199), .B(n29288), .Z(n29250) );
  XOR U29033 ( .A(n29255), .B(n29254), .Z(n29243) );
  XNOR U29034 ( .A(n29289), .B(n29251), .Z(n29254) );
  XOR U29035 ( .A(n29290), .B(n29291), .Z(n29251) );
  AND U29036 ( .A(n29292), .B(n29293), .Z(n29291) );
  XOR U29037 ( .A(n29290), .B(n29294), .Z(n29292) );
  XNOR U29038 ( .A(n29295), .B(n29296), .Z(n29289) );
  AND U29039 ( .A(n29297), .B(n29298), .Z(n29296) );
  XOR U29040 ( .A(n29295), .B(n29299), .Z(n29297) );
  XOR U29041 ( .A(n29300), .B(n29301), .Z(n29255) );
  AND U29042 ( .A(n29302), .B(n29303), .Z(n29301) );
  XOR U29043 ( .A(n29300), .B(n29304), .Z(n29302) );
  XNOR U29044 ( .A(n29188), .B(n29261), .Z(n29263) );
  XNOR U29045 ( .A(n29305), .B(n29306), .Z(n29188) );
  AND U29046 ( .A(n192), .B(n29307), .Z(n29306) );
  XNOR U29047 ( .A(n29308), .B(n29309), .Z(n29307) );
  XOR U29048 ( .A(n29310), .B(n29311), .Z(n29261) );
  AND U29049 ( .A(n29312), .B(n29313), .Z(n29311) );
  XNOR U29050 ( .A(n29310), .B(n29199), .Z(n29313) );
  XOR U29051 ( .A(n29314), .B(n29275), .Z(n29199) );
  XNOR U29052 ( .A(n29315), .B(n29282), .Z(n29275) );
  XOR U29053 ( .A(n29271), .B(n29270), .Z(n29282) );
  XNOR U29054 ( .A(n29316), .B(n29267), .Z(n29270) );
  XOR U29055 ( .A(n29317), .B(n29318), .Z(n29267) );
  AND U29056 ( .A(n29319), .B(n29320), .Z(n29318) );
  XNOR U29057 ( .A(n29321), .B(n29322), .Z(n29319) );
  IV U29058 ( .A(n29317), .Z(n29321) );
  XNOR U29059 ( .A(n29323), .B(n29324), .Z(n29316) );
  NOR U29060 ( .A(n29325), .B(n29326), .Z(n29324) );
  XNOR U29061 ( .A(n29323), .B(n29327), .Z(n29325) );
  XOR U29062 ( .A(n29328), .B(n29329), .Z(n29271) );
  NOR U29063 ( .A(n29330), .B(n29331), .Z(n29329) );
  XNOR U29064 ( .A(n29328), .B(n29332), .Z(n29330) );
  XNOR U29065 ( .A(n29281), .B(n29272), .Z(n29315) );
  XOR U29066 ( .A(n29333), .B(n29334), .Z(n29272) );
  AND U29067 ( .A(n29335), .B(n29336), .Z(n29334) );
  XOR U29068 ( .A(n29333), .B(n29337), .Z(n29335) );
  XOR U29069 ( .A(n29338), .B(n29287), .Z(n29281) );
  XOR U29070 ( .A(n29339), .B(n29340), .Z(n29287) );
  NOR U29071 ( .A(n29341), .B(n29342), .Z(n29340) );
  XOR U29072 ( .A(n29339), .B(n29343), .Z(n29341) );
  XNOR U29073 ( .A(n29286), .B(n29278), .Z(n29338) );
  XOR U29074 ( .A(n29344), .B(n29345), .Z(n29278) );
  AND U29075 ( .A(n29346), .B(n29347), .Z(n29345) );
  XOR U29076 ( .A(n29344), .B(n29348), .Z(n29346) );
  XNOR U29077 ( .A(n29349), .B(n29283), .Z(n29286) );
  XOR U29078 ( .A(n29350), .B(n29351), .Z(n29283) );
  AND U29079 ( .A(n29352), .B(n29353), .Z(n29351) );
  XNOR U29080 ( .A(n29354), .B(n29355), .Z(n29352) );
  IV U29081 ( .A(n29350), .Z(n29354) );
  XNOR U29082 ( .A(n29356), .B(n29357), .Z(n29349) );
  NOR U29083 ( .A(n29358), .B(n29359), .Z(n29357) );
  XNOR U29084 ( .A(n29356), .B(n29360), .Z(n29358) );
  XOR U29085 ( .A(n29276), .B(n29288), .Z(n29314) );
  NOR U29086 ( .A(n29205), .B(n29361), .Z(n29288) );
  XNOR U29087 ( .A(n29294), .B(n29293), .Z(n29276) );
  XNOR U29088 ( .A(n29362), .B(n29299), .Z(n29293) );
  XNOR U29089 ( .A(n29363), .B(n29364), .Z(n29299) );
  NOR U29090 ( .A(n29365), .B(n29366), .Z(n29364) );
  XOR U29091 ( .A(n29363), .B(n29367), .Z(n29365) );
  XNOR U29092 ( .A(n29298), .B(n29290), .Z(n29362) );
  XOR U29093 ( .A(n29368), .B(n29369), .Z(n29290) );
  AND U29094 ( .A(n29370), .B(n29371), .Z(n29369) );
  XOR U29095 ( .A(n29368), .B(n29372), .Z(n29370) );
  XNOR U29096 ( .A(n29373), .B(n29295), .Z(n29298) );
  XOR U29097 ( .A(n29374), .B(n29375), .Z(n29295) );
  AND U29098 ( .A(n29376), .B(n29377), .Z(n29375) );
  XNOR U29099 ( .A(n29378), .B(n29379), .Z(n29376) );
  IV U29100 ( .A(n29374), .Z(n29378) );
  XNOR U29101 ( .A(n29380), .B(n29381), .Z(n29373) );
  NOR U29102 ( .A(n29382), .B(n29383), .Z(n29381) );
  XNOR U29103 ( .A(n29380), .B(n29384), .Z(n29382) );
  XOR U29104 ( .A(n29304), .B(n29303), .Z(n29294) );
  XNOR U29105 ( .A(n29385), .B(n29300), .Z(n29303) );
  XOR U29106 ( .A(n29386), .B(n29387), .Z(n29300) );
  AND U29107 ( .A(n29388), .B(n29389), .Z(n29387) );
  XOR U29108 ( .A(n29386), .B(n29390), .Z(n29388) );
  XNOR U29109 ( .A(n29391), .B(n29392), .Z(n29385) );
  NOR U29110 ( .A(n29393), .B(n29394), .Z(n29392) );
  XNOR U29111 ( .A(n29391), .B(n29395), .Z(n29393) );
  XOR U29112 ( .A(n29396), .B(n29397), .Z(n29304) );
  NOR U29113 ( .A(n29398), .B(n29399), .Z(n29397) );
  XNOR U29114 ( .A(n29396), .B(n29400), .Z(n29398) );
  XNOR U29115 ( .A(n29196), .B(n29310), .Z(n29312) );
  XNOR U29116 ( .A(n29401), .B(n29402), .Z(n29196) );
  AND U29117 ( .A(n192), .B(n29403), .Z(n29402) );
  XNOR U29118 ( .A(n29404), .B(n29405), .Z(n29403) );
  AND U29119 ( .A(n29202), .B(n29205), .Z(n29310) );
  XOR U29120 ( .A(n29406), .B(n29361), .Z(n29205) );
  XNOR U29121 ( .A(p_input[2048]), .B(p_input[96]), .Z(n29361) );
  XNOR U29122 ( .A(n29337), .B(n29336), .Z(n29406) );
  XNOR U29123 ( .A(n29407), .B(n29348), .Z(n29336) );
  XOR U29124 ( .A(n29322), .B(n29320), .Z(n29348) );
  XNOR U29125 ( .A(n29408), .B(n29327), .Z(n29320) );
  XOR U29126 ( .A(p_input[120]), .B(p_input[2072]), .Z(n29327) );
  XOR U29127 ( .A(n29317), .B(n29326), .Z(n29408) );
  XOR U29128 ( .A(n29409), .B(n29323), .Z(n29326) );
  XOR U29129 ( .A(p_input[118]), .B(p_input[2070]), .Z(n29323) );
  XOR U29130 ( .A(p_input[119]), .B(n29410), .Z(n29409) );
  XOR U29131 ( .A(p_input[114]), .B(p_input[2066]), .Z(n29317) );
  XNOR U29132 ( .A(n29332), .B(n29331), .Z(n29322) );
  XOR U29133 ( .A(n29411), .B(n29328), .Z(n29331) );
  XOR U29134 ( .A(p_input[115]), .B(p_input[2067]), .Z(n29328) );
  XOR U29135 ( .A(p_input[116]), .B(n29412), .Z(n29411) );
  XOR U29136 ( .A(p_input[117]), .B(p_input[2069]), .Z(n29332) );
  XNOR U29137 ( .A(n29347), .B(n29333), .Z(n29407) );
  XNOR U29138 ( .A(n28686), .B(p_input[97]), .Z(n29333) );
  XNOR U29139 ( .A(n29413), .B(n29355), .Z(n29347) );
  XNOR U29140 ( .A(n29343), .B(n29342), .Z(n29355) );
  XNOR U29141 ( .A(n29414), .B(n29339), .Z(n29342) );
  XNOR U29142 ( .A(p_input[122]), .B(p_input[2074]), .Z(n29339) );
  XOR U29143 ( .A(p_input[123]), .B(n29415), .Z(n29414) );
  XOR U29144 ( .A(p_input[124]), .B(p_input[2076]), .Z(n29343) );
  XOR U29145 ( .A(n29353), .B(n29416), .Z(n29413) );
  IV U29146 ( .A(n29344), .Z(n29416) );
  XOR U29147 ( .A(p_input[113]), .B(p_input[2065]), .Z(n29344) );
  XNOR U29148 ( .A(n29417), .B(n29360), .Z(n29353) );
  XNOR U29149 ( .A(p_input[127]), .B(n29418), .Z(n29360) );
  XOR U29150 ( .A(n29350), .B(n29359), .Z(n29417) );
  XOR U29151 ( .A(n29419), .B(n29356), .Z(n29359) );
  XOR U29152 ( .A(p_input[125]), .B(p_input[2077]), .Z(n29356) );
  XOR U29153 ( .A(p_input[126]), .B(n29420), .Z(n29419) );
  XOR U29154 ( .A(p_input[121]), .B(p_input[2073]), .Z(n29350) );
  XOR U29155 ( .A(n29372), .B(n29371), .Z(n29337) );
  XNOR U29156 ( .A(n29421), .B(n29379), .Z(n29371) );
  XNOR U29157 ( .A(n29367), .B(n29366), .Z(n29379) );
  XNOR U29158 ( .A(n29422), .B(n29363), .Z(n29366) );
  XNOR U29159 ( .A(p_input[107]), .B(p_input[2059]), .Z(n29363) );
  XOR U29160 ( .A(p_input[108]), .B(n28329), .Z(n29422) );
  XOR U29161 ( .A(p_input[109]), .B(p_input[2061]), .Z(n29367) );
  XNOR U29162 ( .A(n29377), .B(n29368), .Z(n29421) );
  XNOR U29163 ( .A(n28330), .B(p_input[98]), .Z(n29368) );
  XNOR U29164 ( .A(n29423), .B(n29384), .Z(n29377) );
  XNOR U29165 ( .A(p_input[112]), .B(n28332), .Z(n29384) );
  XOR U29166 ( .A(n29374), .B(n29383), .Z(n29423) );
  XOR U29167 ( .A(n29424), .B(n29380), .Z(n29383) );
  XOR U29168 ( .A(p_input[110]), .B(p_input[2062]), .Z(n29380) );
  XOR U29169 ( .A(p_input[111]), .B(n28334), .Z(n29424) );
  XOR U29170 ( .A(p_input[106]), .B(p_input[2058]), .Z(n29374) );
  XOR U29171 ( .A(n29390), .B(n29389), .Z(n29372) );
  XNOR U29172 ( .A(n29425), .B(n29395), .Z(n29389) );
  XOR U29173 ( .A(p_input[105]), .B(p_input[2057]), .Z(n29395) );
  XOR U29174 ( .A(n29386), .B(n29394), .Z(n29425) );
  XOR U29175 ( .A(n29426), .B(n29391), .Z(n29394) );
  XOR U29176 ( .A(p_input[103]), .B(p_input[2055]), .Z(n29391) );
  XOR U29177 ( .A(p_input[104]), .B(n29427), .Z(n29426) );
  XNOR U29178 ( .A(n28337), .B(p_input[99]), .Z(n29386) );
  XNOR U29179 ( .A(n29400), .B(n29399), .Z(n29390) );
  XOR U29180 ( .A(n29428), .B(n29396), .Z(n29399) );
  XOR U29181 ( .A(p_input[100]), .B(p_input[2052]), .Z(n29396) );
  XOR U29182 ( .A(p_input[101]), .B(n29429), .Z(n29428) );
  XOR U29183 ( .A(p_input[102]), .B(p_input[2054]), .Z(n29400) );
  XNOR U29184 ( .A(n29430), .B(n29431), .Z(n29202) );
  AND U29185 ( .A(n192), .B(n29432), .Z(n29431) );
  XNOR U29186 ( .A(n29433), .B(n29434), .Z(n192) );
  AND U29187 ( .A(n29435), .B(n29436), .Z(n29434) );
  XOR U29188 ( .A(n29216), .B(n29433), .Z(n29436) );
  XNOR U29189 ( .A(n29437), .B(n29433), .Z(n29435) );
  XOR U29190 ( .A(n29438), .B(n29439), .Z(n29433) );
  AND U29191 ( .A(n29440), .B(n29441), .Z(n29439) );
  XOR U29192 ( .A(n29231), .B(n29438), .Z(n29441) );
  XOR U29193 ( .A(n29438), .B(n29232), .Z(n29440) );
  XOR U29194 ( .A(n29442), .B(n29443), .Z(n29438) );
  AND U29195 ( .A(n29444), .B(n29445), .Z(n29443) );
  XOR U29196 ( .A(n29259), .B(n29442), .Z(n29445) );
  XOR U29197 ( .A(n29442), .B(n29260), .Z(n29444) );
  XOR U29198 ( .A(n29446), .B(n29447), .Z(n29442) );
  AND U29199 ( .A(n29448), .B(n29449), .Z(n29447) );
  XOR U29200 ( .A(n29308), .B(n29446), .Z(n29449) );
  XOR U29201 ( .A(n29446), .B(n29309), .Z(n29448) );
  XOR U29202 ( .A(n29450), .B(n29451), .Z(n29446) );
  AND U29203 ( .A(n29452), .B(n29453), .Z(n29451) );
  XOR U29204 ( .A(n29450), .B(n29404), .Z(n29453) );
  XNOR U29205 ( .A(n29454), .B(n29455), .Z(n29152) );
  AND U29206 ( .A(n196), .B(n29456), .Z(n29455) );
  XNOR U29207 ( .A(n29457), .B(n29458), .Z(n196) );
  AND U29208 ( .A(n29459), .B(n29460), .Z(n29458) );
  XOR U29209 ( .A(n29457), .B(n29162), .Z(n29460) );
  XNOR U29210 ( .A(n29457), .B(n29112), .Z(n29459) );
  XOR U29211 ( .A(n29461), .B(n29462), .Z(n29457) );
  AND U29212 ( .A(n29463), .B(n29464), .Z(n29462) );
  XNOR U29213 ( .A(n29172), .B(n29461), .Z(n29464) );
  XOR U29214 ( .A(n29461), .B(n29122), .Z(n29463) );
  XOR U29215 ( .A(n29465), .B(n29466), .Z(n29461) );
  AND U29216 ( .A(n29467), .B(n29468), .Z(n29466) );
  XNOR U29217 ( .A(n29182), .B(n29465), .Z(n29468) );
  XOR U29218 ( .A(n29465), .B(n29131), .Z(n29467) );
  XOR U29219 ( .A(n29469), .B(n29470), .Z(n29465) );
  AND U29220 ( .A(n29471), .B(n29472), .Z(n29470) );
  XOR U29221 ( .A(n29469), .B(n29139), .Z(n29471) );
  XOR U29222 ( .A(n29473), .B(n29474), .Z(n29103) );
  AND U29223 ( .A(n200), .B(n29456), .Z(n29474) );
  XNOR U29224 ( .A(n29454), .B(n29473), .Z(n29456) );
  XNOR U29225 ( .A(n29475), .B(n29476), .Z(n200) );
  AND U29226 ( .A(n29477), .B(n29478), .Z(n29476) );
  XNOR U29227 ( .A(n29479), .B(n29475), .Z(n29478) );
  IV U29228 ( .A(n29162), .Z(n29479) );
  XOR U29229 ( .A(n29437), .B(n29480), .Z(n29162) );
  AND U29230 ( .A(n203), .B(n29481), .Z(n29480) );
  XOR U29231 ( .A(n29215), .B(n29212), .Z(n29481) );
  IV U29232 ( .A(n29437), .Z(n29215) );
  XNOR U29233 ( .A(n29112), .B(n29475), .Z(n29477) );
  XOR U29234 ( .A(n29482), .B(n29483), .Z(n29112) );
  AND U29235 ( .A(n219), .B(n29484), .Z(n29483) );
  XOR U29236 ( .A(n29485), .B(n29486), .Z(n29475) );
  AND U29237 ( .A(n29487), .B(n29488), .Z(n29486) );
  XNOR U29238 ( .A(n29485), .B(n29172), .Z(n29488) );
  XOR U29239 ( .A(n29232), .B(n29489), .Z(n29172) );
  AND U29240 ( .A(n203), .B(n29490), .Z(n29489) );
  XOR U29241 ( .A(n29228), .B(n29232), .Z(n29490) );
  XNOR U29242 ( .A(n29491), .B(n29485), .Z(n29487) );
  IV U29243 ( .A(n29122), .Z(n29491) );
  XOR U29244 ( .A(n29492), .B(n29493), .Z(n29122) );
  AND U29245 ( .A(n219), .B(n29494), .Z(n29493) );
  XOR U29246 ( .A(n29495), .B(n29496), .Z(n29485) );
  AND U29247 ( .A(n29497), .B(n29498), .Z(n29496) );
  XNOR U29248 ( .A(n29495), .B(n29182), .Z(n29498) );
  XOR U29249 ( .A(n29260), .B(n29499), .Z(n29182) );
  AND U29250 ( .A(n203), .B(n29500), .Z(n29499) );
  XOR U29251 ( .A(n29256), .B(n29260), .Z(n29500) );
  XOR U29252 ( .A(n29131), .B(n29495), .Z(n29497) );
  XOR U29253 ( .A(n29501), .B(n29502), .Z(n29131) );
  AND U29254 ( .A(n219), .B(n29503), .Z(n29502) );
  XOR U29255 ( .A(n29469), .B(n29504), .Z(n29495) );
  AND U29256 ( .A(n29505), .B(n29472), .Z(n29504) );
  XNOR U29257 ( .A(n29192), .B(n29469), .Z(n29472) );
  XOR U29258 ( .A(n29309), .B(n29506), .Z(n29192) );
  AND U29259 ( .A(n203), .B(n29507), .Z(n29506) );
  XOR U29260 ( .A(n29305), .B(n29309), .Z(n29507) );
  XNOR U29261 ( .A(n29508), .B(n29469), .Z(n29505) );
  IV U29262 ( .A(n29139), .Z(n29508) );
  XOR U29263 ( .A(n29509), .B(n29510), .Z(n29139) );
  AND U29264 ( .A(n219), .B(n29511), .Z(n29510) );
  XOR U29265 ( .A(n29512), .B(n29513), .Z(n29469) );
  AND U29266 ( .A(n29514), .B(n29515), .Z(n29513) );
  XNOR U29267 ( .A(n29512), .B(n29200), .Z(n29515) );
  XOR U29268 ( .A(n29405), .B(n29516), .Z(n29200) );
  AND U29269 ( .A(n203), .B(n29517), .Z(n29516) );
  XOR U29270 ( .A(n29401), .B(n29405), .Z(n29517) );
  XNOR U29271 ( .A(n29518), .B(n29512), .Z(n29514) );
  IV U29272 ( .A(n29149), .Z(n29518) );
  XOR U29273 ( .A(n29519), .B(n29520), .Z(n29149) );
  AND U29274 ( .A(n219), .B(n29521), .Z(n29520) );
  AND U29275 ( .A(n29473), .B(n29454), .Z(n29512) );
  XNOR U29276 ( .A(n29522), .B(n29523), .Z(n29454) );
  AND U29277 ( .A(n203), .B(n29432), .Z(n29523) );
  XNOR U29278 ( .A(n29430), .B(n29522), .Z(n29432) );
  XNOR U29279 ( .A(n29524), .B(n29525), .Z(n203) );
  AND U29280 ( .A(n29526), .B(n29527), .Z(n29525) );
  XNOR U29281 ( .A(n29524), .B(n29212), .Z(n29527) );
  IV U29282 ( .A(n29216), .Z(n29212) );
  XOR U29283 ( .A(n29528), .B(n29529), .Z(n29216) );
  AND U29284 ( .A(n207), .B(n29530), .Z(n29529) );
  XOR U29285 ( .A(n29531), .B(n29528), .Z(n29530) );
  XNOR U29286 ( .A(n29524), .B(n29437), .Z(n29526) );
  XOR U29287 ( .A(n29532), .B(n29533), .Z(n29437) );
  AND U29288 ( .A(n215), .B(n29484), .Z(n29533) );
  XOR U29289 ( .A(n29482), .B(n29532), .Z(n29484) );
  XOR U29290 ( .A(n29534), .B(n29535), .Z(n29524) );
  AND U29291 ( .A(n29536), .B(n29537), .Z(n29535) );
  XNOR U29292 ( .A(n29534), .B(n29228), .Z(n29537) );
  IV U29293 ( .A(n29231), .Z(n29228) );
  XOR U29294 ( .A(n29538), .B(n29539), .Z(n29231) );
  AND U29295 ( .A(n207), .B(n29540), .Z(n29539) );
  XOR U29296 ( .A(n29541), .B(n29538), .Z(n29540) );
  XOR U29297 ( .A(n29232), .B(n29534), .Z(n29536) );
  XOR U29298 ( .A(n29542), .B(n29543), .Z(n29232) );
  AND U29299 ( .A(n215), .B(n29494), .Z(n29543) );
  XOR U29300 ( .A(n29542), .B(n29492), .Z(n29494) );
  XOR U29301 ( .A(n29544), .B(n29545), .Z(n29534) );
  AND U29302 ( .A(n29546), .B(n29547), .Z(n29545) );
  XNOR U29303 ( .A(n29544), .B(n29256), .Z(n29547) );
  IV U29304 ( .A(n29259), .Z(n29256) );
  XOR U29305 ( .A(n29548), .B(n29549), .Z(n29259) );
  AND U29306 ( .A(n207), .B(n29550), .Z(n29549) );
  XNOR U29307 ( .A(n29551), .B(n29548), .Z(n29550) );
  XOR U29308 ( .A(n29260), .B(n29544), .Z(n29546) );
  XOR U29309 ( .A(n29552), .B(n29553), .Z(n29260) );
  AND U29310 ( .A(n215), .B(n29503), .Z(n29553) );
  XOR U29311 ( .A(n29552), .B(n29501), .Z(n29503) );
  XOR U29312 ( .A(n29554), .B(n29555), .Z(n29544) );
  AND U29313 ( .A(n29556), .B(n29557), .Z(n29555) );
  XNOR U29314 ( .A(n29554), .B(n29305), .Z(n29557) );
  IV U29315 ( .A(n29308), .Z(n29305) );
  XOR U29316 ( .A(n29558), .B(n29559), .Z(n29308) );
  AND U29317 ( .A(n207), .B(n29560), .Z(n29559) );
  XOR U29318 ( .A(n29561), .B(n29558), .Z(n29560) );
  XOR U29319 ( .A(n29309), .B(n29554), .Z(n29556) );
  XOR U29320 ( .A(n29562), .B(n29563), .Z(n29309) );
  AND U29321 ( .A(n215), .B(n29511), .Z(n29563) );
  XOR U29322 ( .A(n29562), .B(n29509), .Z(n29511) );
  XOR U29323 ( .A(n29450), .B(n29564), .Z(n29554) );
  AND U29324 ( .A(n29452), .B(n29565), .Z(n29564) );
  XNOR U29325 ( .A(n29450), .B(n29401), .Z(n29565) );
  IV U29326 ( .A(n29404), .Z(n29401) );
  XOR U29327 ( .A(n29566), .B(n29567), .Z(n29404) );
  AND U29328 ( .A(n207), .B(n29568), .Z(n29567) );
  XNOR U29329 ( .A(n29569), .B(n29566), .Z(n29568) );
  XOR U29330 ( .A(n29405), .B(n29450), .Z(n29452) );
  XOR U29331 ( .A(n29570), .B(n29571), .Z(n29405) );
  AND U29332 ( .A(n215), .B(n29521), .Z(n29571) );
  XOR U29333 ( .A(n29570), .B(n29519), .Z(n29521) );
  AND U29334 ( .A(n29522), .B(n29430), .Z(n29450) );
  XNOR U29335 ( .A(n29572), .B(n29573), .Z(n29430) );
  AND U29336 ( .A(n207), .B(n29574), .Z(n29573) );
  XNOR U29337 ( .A(n29575), .B(n29572), .Z(n29574) );
  XNOR U29338 ( .A(n29576), .B(n29577), .Z(n207) );
  AND U29339 ( .A(n29578), .B(n29579), .Z(n29577) );
  XOR U29340 ( .A(n29531), .B(n29576), .Z(n29579) );
  AND U29341 ( .A(n29580), .B(n29581), .Z(n29531) );
  XNOR U29342 ( .A(n29528), .B(n29576), .Z(n29578) );
  XNOR U29343 ( .A(n29582), .B(n29583), .Z(n29528) );
  AND U29344 ( .A(n211), .B(n29584), .Z(n29583) );
  XNOR U29345 ( .A(n29585), .B(n29586), .Z(n29584) );
  XOR U29346 ( .A(n29587), .B(n29588), .Z(n29576) );
  AND U29347 ( .A(n29589), .B(n29590), .Z(n29588) );
  XNOR U29348 ( .A(n29587), .B(n29580), .Z(n29590) );
  IV U29349 ( .A(n29541), .Z(n29580) );
  XOR U29350 ( .A(n29591), .B(n29592), .Z(n29541) );
  XOR U29351 ( .A(n29593), .B(n29581), .Z(n29592) );
  AND U29352 ( .A(n29551), .B(n29594), .Z(n29581) );
  AND U29353 ( .A(n29595), .B(n29596), .Z(n29593) );
  XOR U29354 ( .A(n29597), .B(n29591), .Z(n29595) );
  XNOR U29355 ( .A(n29538), .B(n29587), .Z(n29589) );
  XNOR U29356 ( .A(n29598), .B(n29599), .Z(n29538) );
  AND U29357 ( .A(n211), .B(n29600), .Z(n29599) );
  XNOR U29358 ( .A(n29601), .B(n29602), .Z(n29600) );
  XOR U29359 ( .A(n29603), .B(n29604), .Z(n29587) );
  AND U29360 ( .A(n29605), .B(n29606), .Z(n29604) );
  XNOR U29361 ( .A(n29603), .B(n29551), .Z(n29606) );
  XOR U29362 ( .A(n29607), .B(n29596), .Z(n29551) );
  XNOR U29363 ( .A(n29608), .B(n29591), .Z(n29596) );
  XOR U29364 ( .A(n29609), .B(n29610), .Z(n29591) );
  AND U29365 ( .A(n29611), .B(n29612), .Z(n29610) );
  XOR U29366 ( .A(n29613), .B(n29609), .Z(n29611) );
  XNOR U29367 ( .A(n29614), .B(n29615), .Z(n29608) );
  AND U29368 ( .A(n29616), .B(n29617), .Z(n29615) );
  XOR U29369 ( .A(n29614), .B(n29618), .Z(n29616) );
  XNOR U29370 ( .A(n29597), .B(n29594), .Z(n29607) );
  AND U29371 ( .A(n29619), .B(n29620), .Z(n29594) );
  XOR U29372 ( .A(n29621), .B(n29622), .Z(n29597) );
  AND U29373 ( .A(n29623), .B(n29624), .Z(n29622) );
  XOR U29374 ( .A(n29621), .B(n29625), .Z(n29623) );
  XNOR U29375 ( .A(n29548), .B(n29603), .Z(n29605) );
  XNOR U29376 ( .A(n29626), .B(n29627), .Z(n29548) );
  AND U29377 ( .A(n211), .B(n29628), .Z(n29627) );
  XNOR U29378 ( .A(n29629), .B(n29630), .Z(n29628) );
  XOR U29379 ( .A(n29631), .B(n29632), .Z(n29603) );
  AND U29380 ( .A(n29633), .B(n29634), .Z(n29632) );
  XNOR U29381 ( .A(n29631), .B(n29619), .Z(n29634) );
  IV U29382 ( .A(n29561), .Z(n29619) );
  XNOR U29383 ( .A(n29635), .B(n29612), .Z(n29561) );
  XNOR U29384 ( .A(n29636), .B(n29618), .Z(n29612) );
  XOR U29385 ( .A(n29637), .B(n29638), .Z(n29618) );
  AND U29386 ( .A(n29639), .B(n29640), .Z(n29638) );
  XOR U29387 ( .A(n29637), .B(n29641), .Z(n29639) );
  XNOR U29388 ( .A(n29617), .B(n29609), .Z(n29636) );
  XOR U29389 ( .A(n29642), .B(n29643), .Z(n29609) );
  AND U29390 ( .A(n29644), .B(n29645), .Z(n29643) );
  XNOR U29391 ( .A(n29646), .B(n29642), .Z(n29644) );
  XNOR U29392 ( .A(n29647), .B(n29614), .Z(n29617) );
  XOR U29393 ( .A(n29648), .B(n29649), .Z(n29614) );
  AND U29394 ( .A(n29650), .B(n29651), .Z(n29649) );
  XOR U29395 ( .A(n29648), .B(n29652), .Z(n29650) );
  XNOR U29396 ( .A(n29653), .B(n29654), .Z(n29647) );
  AND U29397 ( .A(n29655), .B(n29656), .Z(n29654) );
  XNOR U29398 ( .A(n29653), .B(n29657), .Z(n29655) );
  XNOR U29399 ( .A(n29613), .B(n29620), .Z(n29635) );
  AND U29400 ( .A(n29569), .B(n29658), .Z(n29620) );
  XOR U29401 ( .A(n29625), .B(n29624), .Z(n29613) );
  XNOR U29402 ( .A(n29659), .B(n29621), .Z(n29624) );
  XOR U29403 ( .A(n29660), .B(n29661), .Z(n29621) );
  AND U29404 ( .A(n29662), .B(n29663), .Z(n29661) );
  XOR U29405 ( .A(n29660), .B(n29664), .Z(n29662) );
  XNOR U29406 ( .A(n29665), .B(n29666), .Z(n29659) );
  AND U29407 ( .A(n29667), .B(n29668), .Z(n29666) );
  XOR U29408 ( .A(n29665), .B(n29669), .Z(n29667) );
  XOR U29409 ( .A(n29670), .B(n29671), .Z(n29625) );
  AND U29410 ( .A(n29672), .B(n29673), .Z(n29671) );
  XOR U29411 ( .A(n29670), .B(n29674), .Z(n29672) );
  XNOR U29412 ( .A(n29558), .B(n29631), .Z(n29633) );
  XNOR U29413 ( .A(n29675), .B(n29676), .Z(n29558) );
  AND U29414 ( .A(n211), .B(n29677), .Z(n29676) );
  XNOR U29415 ( .A(n29678), .B(n29679), .Z(n29677) );
  XOR U29416 ( .A(n29680), .B(n29681), .Z(n29631) );
  AND U29417 ( .A(n29682), .B(n29683), .Z(n29681) );
  XNOR U29418 ( .A(n29680), .B(n29569), .Z(n29683) );
  XOR U29419 ( .A(n29684), .B(n29645), .Z(n29569) );
  XNOR U29420 ( .A(n29685), .B(n29652), .Z(n29645) );
  XOR U29421 ( .A(n29641), .B(n29640), .Z(n29652) );
  XNOR U29422 ( .A(n29686), .B(n29637), .Z(n29640) );
  XOR U29423 ( .A(n29687), .B(n29688), .Z(n29637) );
  AND U29424 ( .A(n29689), .B(n29690), .Z(n29688) );
  XNOR U29425 ( .A(n29691), .B(n29692), .Z(n29689) );
  IV U29426 ( .A(n29687), .Z(n29691) );
  XNOR U29427 ( .A(n29693), .B(n29694), .Z(n29686) );
  NOR U29428 ( .A(n29695), .B(n29696), .Z(n29694) );
  XNOR U29429 ( .A(n29693), .B(n29697), .Z(n29695) );
  XOR U29430 ( .A(n29698), .B(n29699), .Z(n29641) );
  NOR U29431 ( .A(n29700), .B(n29701), .Z(n29699) );
  XNOR U29432 ( .A(n29698), .B(n29702), .Z(n29700) );
  XNOR U29433 ( .A(n29651), .B(n29642), .Z(n29685) );
  XOR U29434 ( .A(n29703), .B(n29704), .Z(n29642) );
  AND U29435 ( .A(n29705), .B(n29706), .Z(n29704) );
  XOR U29436 ( .A(n29703), .B(n29707), .Z(n29705) );
  XOR U29437 ( .A(n29708), .B(n29657), .Z(n29651) );
  XOR U29438 ( .A(n29709), .B(n29710), .Z(n29657) );
  NOR U29439 ( .A(n29711), .B(n29712), .Z(n29710) );
  XOR U29440 ( .A(n29709), .B(n29713), .Z(n29711) );
  XNOR U29441 ( .A(n29656), .B(n29648), .Z(n29708) );
  XOR U29442 ( .A(n29714), .B(n29715), .Z(n29648) );
  AND U29443 ( .A(n29716), .B(n29717), .Z(n29715) );
  XOR U29444 ( .A(n29714), .B(n29718), .Z(n29716) );
  XNOR U29445 ( .A(n29719), .B(n29653), .Z(n29656) );
  XOR U29446 ( .A(n29720), .B(n29721), .Z(n29653) );
  AND U29447 ( .A(n29722), .B(n29723), .Z(n29721) );
  XNOR U29448 ( .A(n29724), .B(n29725), .Z(n29722) );
  IV U29449 ( .A(n29720), .Z(n29724) );
  XNOR U29450 ( .A(n29726), .B(n29727), .Z(n29719) );
  NOR U29451 ( .A(n29728), .B(n29729), .Z(n29727) );
  XNOR U29452 ( .A(n29726), .B(n29730), .Z(n29728) );
  XOR U29453 ( .A(n29646), .B(n29658), .Z(n29684) );
  NOR U29454 ( .A(n29575), .B(n29731), .Z(n29658) );
  XNOR U29455 ( .A(n29664), .B(n29663), .Z(n29646) );
  XNOR U29456 ( .A(n29732), .B(n29669), .Z(n29663) );
  XNOR U29457 ( .A(n29733), .B(n29734), .Z(n29669) );
  NOR U29458 ( .A(n29735), .B(n29736), .Z(n29734) );
  XOR U29459 ( .A(n29733), .B(n29737), .Z(n29735) );
  XNOR U29460 ( .A(n29668), .B(n29660), .Z(n29732) );
  XOR U29461 ( .A(n29738), .B(n29739), .Z(n29660) );
  AND U29462 ( .A(n29740), .B(n29741), .Z(n29739) );
  XOR U29463 ( .A(n29738), .B(n29742), .Z(n29740) );
  XNOR U29464 ( .A(n29743), .B(n29665), .Z(n29668) );
  XOR U29465 ( .A(n29744), .B(n29745), .Z(n29665) );
  AND U29466 ( .A(n29746), .B(n29747), .Z(n29745) );
  XNOR U29467 ( .A(n29748), .B(n29749), .Z(n29746) );
  IV U29468 ( .A(n29744), .Z(n29748) );
  XNOR U29469 ( .A(n29750), .B(n29751), .Z(n29743) );
  NOR U29470 ( .A(n29752), .B(n29753), .Z(n29751) );
  XNOR U29471 ( .A(n29750), .B(n29754), .Z(n29752) );
  XOR U29472 ( .A(n29674), .B(n29673), .Z(n29664) );
  XNOR U29473 ( .A(n29755), .B(n29670), .Z(n29673) );
  XOR U29474 ( .A(n29756), .B(n29757), .Z(n29670) );
  AND U29475 ( .A(n29758), .B(n29759), .Z(n29757) );
  XNOR U29476 ( .A(n29760), .B(n29761), .Z(n29758) );
  IV U29477 ( .A(n29756), .Z(n29760) );
  XNOR U29478 ( .A(n29762), .B(n29763), .Z(n29755) );
  NOR U29479 ( .A(n29764), .B(n29765), .Z(n29763) );
  XNOR U29480 ( .A(n29762), .B(n29766), .Z(n29764) );
  XOR U29481 ( .A(n29767), .B(n29768), .Z(n29674) );
  NOR U29482 ( .A(n29769), .B(n29770), .Z(n29768) );
  XNOR U29483 ( .A(n29767), .B(n29771), .Z(n29769) );
  XNOR U29484 ( .A(n29566), .B(n29680), .Z(n29682) );
  XNOR U29485 ( .A(n29772), .B(n29773), .Z(n29566) );
  AND U29486 ( .A(n211), .B(n29774), .Z(n29773) );
  XNOR U29487 ( .A(n29775), .B(n29776), .Z(n29774) );
  AND U29488 ( .A(n29572), .B(n29575), .Z(n29680) );
  XOR U29489 ( .A(n29777), .B(n29731), .Z(n29575) );
  XNOR U29490 ( .A(p_input[128]), .B(p_input[2048]), .Z(n29731) );
  XNOR U29491 ( .A(n29707), .B(n29706), .Z(n29777) );
  XNOR U29492 ( .A(n29778), .B(n29718), .Z(n29706) );
  XOR U29493 ( .A(n29692), .B(n29690), .Z(n29718) );
  XNOR U29494 ( .A(n29779), .B(n29697), .Z(n29690) );
  XOR U29495 ( .A(p_input[152]), .B(p_input[2072]), .Z(n29697) );
  XOR U29496 ( .A(n29687), .B(n29696), .Z(n29779) );
  XOR U29497 ( .A(n29780), .B(n29693), .Z(n29696) );
  XOR U29498 ( .A(p_input[150]), .B(p_input[2070]), .Z(n29693) );
  XOR U29499 ( .A(p_input[151]), .B(n29410), .Z(n29780) );
  XOR U29500 ( .A(p_input[146]), .B(p_input[2066]), .Z(n29687) );
  XNOR U29501 ( .A(n29702), .B(n29701), .Z(n29692) );
  XOR U29502 ( .A(n29781), .B(n29698), .Z(n29701) );
  XOR U29503 ( .A(p_input[147]), .B(p_input[2067]), .Z(n29698) );
  XOR U29504 ( .A(p_input[148]), .B(n29412), .Z(n29781) );
  XOR U29505 ( .A(p_input[149]), .B(p_input[2069]), .Z(n29702) );
  XOR U29506 ( .A(n29717), .B(n29782), .Z(n29778) );
  IV U29507 ( .A(n29703), .Z(n29782) );
  XOR U29508 ( .A(p_input[129]), .B(p_input[2049]), .Z(n29703) );
  XNOR U29509 ( .A(n29783), .B(n29725), .Z(n29717) );
  XNOR U29510 ( .A(n29713), .B(n29712), .Z(n29725) );
  XNOR U29511 ( .A(n29784), .B(n29709), .Z(n29712) );
  XNOR U29512 ( .A(p_input[154]), .B(p_input[2074]), .Z(n29709) );
  XOR U29513 ( .A(p_input[155]), .B(n29415), .Z(n29784) );
  XOR U29514 ( .A(p_input[156]), .B(p_input[2076]), .Z(n29713) );
  XOR U29515 ( .A(n29723), .B(n29785), .Z(n29783) );
  IV U29516 ( .A(n29714), .Z(n29785) );
  XOR U29517 ( .A(p_input[145]), .B(p_input[2065]), .Z(n29714) );
  XNOR U29518 ( .A(n29786), .B(n29730), .Z(n29723) );
  XNOR U29519 ( .A(p_input[159]), .B(n29418), .Z(n29730) );
  XOR U29520 ( .A(n29720), .B(n29729), .Z(n29786) );
  XOR U29521 ( .A(n29787), .B(n29726), .Z(n29729) );
  XOR U29522 ( .A(p_input[157]), .B(p_input[2077]), .Z(n29726) );
  XOR U29523 ( .A(p_input[158]), .B(n29420), .Z(n29787) );
  XOR U29524 ( .A(p_input[153]), .B(p_input[2073]), .Z(n29720) );
  XOR U29525 ( .A(n29742), .B(n29741), .Z(n29707) );
  XNOR U29526 ( .A(n29788), .B(n29749), .Z(n29741) );
  XNOR U29527 ( .A(n29737), .B(n29736), .Z(n29749) );
  XNOR U29528 ( .A(n29789), .B(n29733), .Z(n29736) );
  XNOR U29529 ( .A(p_input[139]), .B(p_input[2059]), .Z(n29733) );
  XOR U29530 ( .A(p_input[140]), .B(n28329), .Z(n29789) );
  XOR U29531 ( .A(p_input[141]), .B(p_input[2061]), .Z(n29737) );
  XOR U29532 ( .A(n29747), .B(n29790), .Z(n29788) );
  IV U29533 ( .A(n29738), .Z(n29790) );
  XOR U29534 ( .A(p_input[130]), .B(p_input[2050]), .Z(n29738) );
  XNOR U29535 ( .A(n29791), .B(n29754), .Z(n29747) );
  XNOR U29536 ( .A(p_input[144]), .B(n28332), .Z(n29754) );
  XOR U29537 ( .A(n29744), .B(n29753), .Z(n29791) );
  XOR U29538 ( .A(n29792), .B(n29750), .Z(n29753) );
  XOR U29539 ( .A(p_input[142]), .B(p_input[2062]), .Z(n29750) );
  XOR U29540 ( .A(p_input[143]), .B(n28334), .Z(n29792) );
  XOR U29541 ( .A(p_input[138]), .B(p_input[2058]), .Z(n29744) );
  XOR U29542 ( .A(n29761), .B(n29759), .Z(n29742) );
  XNOR U29543 ( .A(n29793), .B(n29766), .Z(n29759) );
  XOR U29544 ( .A(p_input[137]), .B(p_input[2057]), .Z(n29766) );
  XOR U29545 ( .A(n29756), .B(n29765), .Z(n29793) );
  XOR U29546 ( .A(n29794), .B(n29762), .Z(n29765) );
  XOR U29547 ( .A(p_input[135]), .B(p_input[2055]), .Z(n29762) );
  XOR U29548 ( .A(p_input[136]), .B(n29427), .Z(n29794) );
  XOR U29549 ( .A(p_input[131]), .B(p_input[2051]), .Z(n29756) );
  XNOR U29550 ( .A(n29771), .B(n29770), .Z(n29761) );
  XOR U29551 ( .A(n29795), .B(n29767), .Z(n29770) );
  XOR U29552 ( .A(p_input[132]), .B(p_input[2052]), .Z(n29767) );
  XOR U29553 ( .A(p_input[133]), .B(n29429), .Z(n29795) );
  XOR U29554 ( .A(p_input[134]), .B(p_input[2054]), .Z(n29771) );
  XNOR U29555 ( .A(n29796), .B(n29797), .Z(n29572) );
  AND U29556 ( .A(n211), .B(n29798), .Z(n29797) );
  XNOR U29557 ( .A(n29799), .B(n29800), .Z(n211) );
  AND U29558 ( .A(n29801), .B(n29802), .Z(n29800) );
  XOR U29559 ( .A(n29586), .B(n29799), .Z(n29802) );
  XNOR U29560 ( .A(n29803), .B(n29799), .Z(n29801) );
  XOR U29561 ( .A(n29804), .B(n29805), .Z(n29799) );
  AND U29562 ( .A(n29806), .B(n29807), .Z(n29805) );
  XOR U29563 ( .A(n29601), .B(n29804), .Z(n29807) );
  XOR U29564 ( .A(n29804), .B(n29602), .Z(n29806) );
  XOR U29565 ( .A(n29808), .B(n29809), .Z(n29804) );
  AND U29566 ( .A(n29810), .B(n29811), .Z(n29809) );
  XOR U29567 ( .A(n29629), .B(n29808), .Z(n29811) );
  XOR U29568 ( .A(n29808), .B(n29630), .Z(n29810) );
  XOR U29569 ( .A(n29812), .B(n29813), .Z(n29808) );
  AND U29570 ( .A(n29814), .B(n29815), .Z(n29813) );
  XOR U29571 ( .A(n29678), .B(n29812), .Z(n29815) );
  XOR U29572 ( .A(n29812), .B(n29679), .Z(n29814) );
  XOR U29573 ( .A(n29816), .B(n29817), .Z(n29812) );
  AND U29574 ( .A(n29818), .B(n29819), .Z(n29817) );
  XOR U29575 ( .A(n29816), .B(n29775), .Z(n29819) );
  XNOR U29576 ( .A(n29820), .B(n29821), .Z(n29522) );
  AND U29577 ( .A(n215), .B(n29822), .Z(n29821) );
  XNOR U29578 ( .A(n29823), .B(n29824), .Z(n215) );
  AND U29579 ( .A(n29825), .B(n29826), .Z(n29824) );
  XOR U29580 ( .A(n29823), .B(n29532), .Z(n29826) );
  XNOR U29581 ( .A(n29823), .B(n29482), .Z(n29825) );
  XOR U29582 ( .A(n29827), .B(n29828), .Z(n29823) );
  AND U29583 ( .A(n29829), .B(n29830), .Z(n29828) );
  XNOR U29584 ( .A(n29542), .B(n29827), .Z(n29830) );
  XOR U29585 ( .A(n29827), .B(n29492), .Z(n29829) );
  XOR U29586 ( .A(n29831), .B(n29832), .Z(n29827) );
  AND U29587 ( .A(n29833), .B(n29834), .Z(n29832) );
  XNOR U29588 ( .A(n29552), .B(n29831), .Z(n29834) );
  XOR U29589 ( .A(n29831), .B(n29501), .Z(n29833) );
  XOR U29590 ( .A(n29835), .B(n29836), .Z(n29831) );
  AND U29591 ( .A(n29837), .B(n29838), .Z(n29836) );
  XOR U29592 ( .A(n29835), .B(n29509), .Z(n29837) );
  XOR U29593 ( .A(n29839), .B(n29840), .Z(n29473) );
  AND U29594 ( .A(n219), .B(n29822), .Z(n29840) );
  XNOR U29595 ( .A(n29820), .B(n29839), .Z(n29822) );
  XNOR U29596 ( .A(n29841), .B(n29842), .Z(n219) );
  AND U29597 ( .A(n29843), .B(n29844), .Z(n29842) );
  XNOR U29598 ( .A(n29845), .B(n29841), .Z(n29844) );
  IV U29599 ( .A(n29532), .Z(n29845) );
  XOR U29600 ( .A(n29803), .B(n29846), .Z(n29532) );
  AND U29601 ( .A(n222), .B(n29847), .Z(n29846) );
  XOR U29602 ( .A(n29585), .B(n29582), .Z(n29847) );
  IV U29603 ( .A(n29803), .Z(n29585) );
  XNOR U29604 ( .A(n29482), .B(n29841), .Z(n29843) );
  XOR U29605 ( .A(n29848), .B(n29849), .Z(n29482) );
  AND U29606 ( .A(n238), .B(n29850), .Z(n29849) );
  XOR U29607 ( .A(n29851), .B(n29852), .Z(n29841) );
  AND U29608 ( .A(n29853), .B(n29854), .Z(n29852) );
  XNOR U29609 ( .A(n29851), .B(n29542), .Z(n29854) );
  XOR U29610 ( .A(n29602), .B(n29855), .Z(n29542) );
  AND U29611 ( .A(n222), .B(n29856), .Z(n29855) );
  XOR U29612 ( .A(n29598), .B(n29602), .Z(n29856) );
  XNOR U29613 ( .A(n29857), .B(n29851), .Z(n29853) );
  IV U29614 ( .A(n29492), .Z(n29857) );
  XOR U29615 ( .A(n29858), .B(n29859), .Z(n29492) );
  AND U29616 ( .A(n238), .B(n29860), .Z(n29859) );
  XOR U29617 ( .A(n29861), .B(n29862), .Z(n29851) );
  AND U29618 ( .A(n29863), .B(n29864), .Z(n29862) );
  XNOR U29619 ( .A(n29861), .B(n29552), .Z(n29864) );
  XOR U29620 ( .A(n29630), .B(n29865), .Z(n29552) );
  AND U29621 ( .A(n222), .B(n29866), .Z(n29865) );
  XOR U29622 ( .A(n29626), .B(n29630), .Z(n29866) );
  XOR U29623 ( .A(n29501), .B(n29861), .Z(n29863) );
  XOR U29624 ( .A(n29867), .B(n29868), .Z(n29501) );
  AND U29625 ( .A(n238), .B(n29869), .Z(n29868) );
  XOR U29626 ( .A(n29835), .B(n29870), .Z(n29861) );
  AND U29627 ( .A(n29871), .B(n29838), .Z(n29870) );
  XNOR U29628 ( .A(n29562), .B(n29835), .Z(n29838) );
  XOR U29629 ( .A(n29679), .B(n29872), .Z(n29562) );
  AND U29630 ( .A(n222), .B(n29873), .Z(n29872) );
  XOR U29631 ( .A(n29675), .B(n29679), .Z(n29873) );
  XNOR U29632 ( .A(n29874), .B(n29835), .Z(n29871) );
  IV U29633 ( .A(n29509), .Z(n29874) );
  XOR U29634 ( .A(n29875), .B(n29876), .Z(n29509) );
  AND U29635 ( .A(n238), .B(n29877), .Z(n29876) );
  XOR U29636 ( .A(n29878), .B(n29879), .Z(n29835) );
  AND U29637 ( .A(n29880), .B(n29881), .Z(n29879) );
  XNOR U29638 ( .A(n29878), .B(n29570), .Z(n29881) );
  XOR U29639 ( .A(n29776), .B(n29882), .Z(n29570) );
  AND U29640 ( .A(n222), .B(n29883), .Z(n29882) );
  XOR U29641 ( .A(n29772), .B(n29776), .Z(n29883) );
  XNOR U29642 ( .A(n29884), .B(n29878), .Z(n29880) );
  IV U29643 ( .A(n29519), .Z(n29884) );
  XOR U29644 ( .A(n29885), .B(n29886), .Z(n29519) );
  AND U29645 ( .A(n238), .B(n29887), .Z(n29886) );
  AND U29646 ( .A(n29839), .B(n29820), .Z(n29878) );
  XNOR U29647 ( .A(n29888), .B(n29889), .Z(n29820) );
  AND U29648 ( .A(n222), .B(n29798), .Z(n29889) );
  XNOR U29649 ( .A(n29796), .B(n29888), .Z(n29798) );
  XNOR U29650 ( .A(n29890), .B(n29891), .Z(n222) );
  AND U29651 ( .A(n29892), .B(n29893), .Z(n29891) );
  XNOR U29652 ( .A(n29890), .B(n29582), .Z(n29893) );
  IV U29653 ( .A(n29586), .Z(n29582) );
  XOR U29654 ( .A(n29894), .B(n29895), .Z(n29586) );
  AND U29655 ( .A(n226), .B(n29896), .Z(n29895) );
  XOR U29656 ( .A(n29897), .B(n29894), .Z(n29896) );
  XNOR U29657 ( .A(n29890), .B(n29803), .Z(n29892) );
  XOR U29658 ( .A(n29898), .B(n29899), .Z(n29803) );
  AND U29659 ( .A(n234), .B(n29850), .Z(n29899) );
  XOR U29660 ( .A(n29848), .B(n29898), .Z(n29850) );
  XOR U29661 ( .A(n29900), .B(n29901), .Z(n29890) );
  AND U29662 ( .A(n29902), .B(n29903), .Z(n29901) );
  XNOR U29663 ( .A(n29900), .B(n29598), .Z(n29903) );
  IV U29664 ( .A(n29601), .Z(n29598) );
  XOR U29665 ( .A(n29904), .B(n29905), .Z(n29601) );
  AND U29666 ( .A(n226), .B(n29906), .Z(n29905) );
  XOR U29667 ( .A(n29907), .B(n29904), .Z(n29906) );
  XOR U29668 ( .A(n29602), .B(n29900), .Z(n29902) );
  XOR U29669 ( .A(n29908), .B(n29909), .Z(n29602) );
  AND U29670 ( .A(n234), .B(n29860), .Z(n29909) );
  XOR U29671 ( .A(n29908), .B(n29858), .Z(n29860) );
  XOR U29672 ( .A(n29910), .B(n29911), .Z(n29900) );
  AND U29673 ( .A(n29912), .B(n29913), .Z(n29911) );
  XNOR U29674 ( .A(n29910), .B(n29626), .Z(n29913) );
  IV U29675 ( .A(n29629), .Z(n29626) );
  XOR U29676 ( .A(n29914), .B(n29915), .Z(n29629) );
  AND U29677 ( .A(n226), .B(n29916), .Z(n29915) );
  XNOR U29678 ( .A(n29917), .B(n29914), .Z(n29916) );
  XOR U29679 ( .A(n29630), .B(n29910), .Z(n29912) );
  XOR U29680 ( .A(n29918), .B(n29919), .Z(n29630) );
  AND U29681 ( .A(n234), .B(n29869), .Z(n29919) );
  XOR U29682 ( .A(n29918), .B(n29867), .Z(n29869) );
  XOR U29683 ( .A(n29920), .B(n29921), .Z(n29910) );
  AND U29684 ( .A(n29922), .B(n29923), .Z(n29921) );
  XNOR U29685 ( .A(n29920), .B(n29675), .Z(n29923) );
  IV U29686 ( .A(n29678), .Z(n29675) );
  XOR U29687 ( .A(n29924), .B(n29925), .Z(n29678) );
  AND U29688 ( .A(n226), .B(n29926), .Z(n29925) );
  XOR U29689 ( .A(n29927), .B(n29924), .Z(n29926) );
  XOR U29690 ( .A(n29679), .B(n29920), .Z(n29922) );
  XOR U29691 ( .A(n29928), .B(n29929), .Z(n29679) );
  AND U29692 ( .A(n234), .B(n29877), .Z(n29929) );
  XOR U29693 ( .A(n29928), .B(n29875), .Z(n29877) );
  XOR U29694 ( .A(n29816), .B(n29930), .Z(n29920) );
  AND U29695 ( .A(n29818), .B(n29931), .Z(n29930) );
  XNOR U29696 ( .A(n29816), .B(n29772), .Z(n29931) );
  IV U29697 ( .A(n29775), .Z(n29772) );
  XOR U29698 ( .A(n29932), .B(n29933), .Z(n29775) );
  AND U29699 ( .A(n226), .B(n29934), .Z(n29933) );
  XNOR U29700 ( .A(n29935), .B(n29932), .Z(n29934) );
  XOR U29701 ( .A(n29776), .B(n29816), .Z(n29818) );
  XOR U29702 ( .A(n29936), .B(n29937), .Z(n29776) );
  AND U29703 ( .A(n234), .B(n29887), .Z(n29937) );
  XOR U29704 ( .A(n29936), .B(n29885), .Z(n29887) );
  AND U29705 ( .A(n29888), .B(n29796), .Z(n29816) );
  XNOR U29706 ( .A(n29938), .B(n29939), .Z(n29796) );
  AND U29707 ( .A(n226), .B(n29940), .Z(n29939) );
  XNOR U29708 ( .A(n29941), .B(n29938), .Z(n29940) );
  XNOR U29709 ( .A(n29942), .B(n29943), .Z(n226) );
  AND U29710 ( .A(n29944), .B(n29945), .Z(n29943) );
  XOR U29711 ( .A(n29897), .B(n29942), .Z(n29945) );
  AND U29712 ( .A(n29946), .B(n29947), .Z(n29897) );
  XNOR U29713 ( .A(n29894), .B(n29942), .Z(n29944) );
  XNOR U29714 ( .A(n29948), .B(n29949), .Z(n29894) );
  AND U29715 ( .A(n230), .B(n29950), .Z(n29949) );
  XNOR U29716 ( .A(n29951), .B(n29952), .Z(n29950) );
  XOR U29717 ( .A(n29953), .B(n29954), .Z(n29942) );
  AND U29718 ( .A(n29955), .B(n29956), .Z(n29954) );
  XNOR U29719 ( .A(n29953), .B(n29946), .Z(n29956) );
  IV U29720 ( .A(n29907), .Z(n29946) );
  XOR U29721 ( .A(n29957), .B(n29958), .Z(n29907) );
  XOR U29722 ( .A(n29959), .B(n29947), .Z(n29958) );
  AND U29723 ( .A(n29917), .B(n29960), .Z(n29947) );
  AND U29724 ( .A(n29961), .B(n29962), .Z(n29959) );
  XOR U29725 ( .A(n29963), .B(n29957), .Z(n29961) );
  XNOR U29726 ( .A(n29904), .B(n29953), .Z(n29955) );
  XNOR U29727 ( .A(n29964), .B(n29965), .Z(n29904) );
  AND U29728 ( .A(n230), .B(n29966), .Z(n29965) );
  XNOR U29729 ( .A(n29967), .B(n29968), .Z(n29966) );
  XOR U29730 ( .A(n29969), .B(n29970), .Z(n29953) );
  AND U29731 ( .A(n29971), .B(n29972), .Z(n29970) );
  XNOR U29732 ( .A(n29969), .B(n29917), .Z(n29972) );
  XOR U29733 ( .A(n29973), .B(n29962), .Z(n29917) );
  XNOR U29734 ( .A(n29974), .B(n29957), .Z(n29962) );
  XOR U29735 ( .A(n29975), .B(n29976), .Z(n29957) );
  AND U29736 ( .A(n29977), .B(n29978), .Z(n29976) );
  XOR U29737 ( .A(n29979), .B(n29975), .Z(n29977) );
  XNOR U29738 ( .A(n29980), .B(n29981), .Z(n29974) );
  AND U29739 ( .A(n29982), .B(n29983), .Z(n29981) );
  XOR U29740 ( .A(n29980), .B(n29984), .Z(n29982) );
  XNOR U29741 ( .A(n29963), .B(n29960), .Z(n29973) );
  AND U29742 ( .A(n29985), .B(n29986), .Z(n29960) );
  XOR U29743 ( .A(n29987), .B(n29988), .Z(n29963) );
  AND U29744 ( .A(n29989), .B(n29990), .Z(n29988) );
  XOR U29745 ( .A(n29987), .B(n29991), .Z(n29989) );
  XNOR U29746 ( .A(n29914), .B(n29969), .Z(n29971) );
  XNOR U29747 ( .A(n29992), .B(n29993), .Z(n29914) );
  AND U29748 ( .A(n230), .B(n29994), .Z(n29993) );
  XNOR U29749 ( .A(n29995), .B(n29996), .Z(n29994) );
  XOR U29750 ( .A(n29997), .B(n29998), .Z(n29969) );
  AND U29751 ( .A(n29999), .B(n30000), .Z(n29998) );
  XNOR U29752 ( .A(n29997), .B(n29985), .Z(n30000) );
  IV U29753 ( .A(n29927), .Z(n29985) );
  XNOR U29754 ( .A(n30001), .B(n29978), .Z(n29927) );
  XNOR U29755 ( .A(n30002), .B(n29984), .Z(n29978) );
  XOR U29756 ( .A(n30003), .B(n30004), .Z(n29984) );
  AND U29757 ( .A(n30005), .B(n30006), .Z(n30004) );
  XOR U29758 ( .A(n30003), .B(n30007), .Z(n30005) );
  XNOR U29759 ( .A(n29983), .B(n29975), .Z(n30002) );
  XOR U29760 ( .A(n30008), .B(n30009), .Z(n29975) );
  AND U29761 ( .A(n30010), .B(n30011), .Z(n30009) );
  XNOR U29762 ( .A(n30012), .B(n30008), .Z(n30010) );
  XNOR U29763 ( .A(n30013), .B(n29980), .Z(n29983) );
  XOR U29764 ( .A(n30014), .B(n30015), .Z(n29980) );
  AND U29765 ( .A(n30016), .B(n30017), .Z(n30015) );
  XOR U29766 ( .A(n30014), .B(n30018), .Z(n30016) );
  XNOR U29767 ( .A(n30019), .B(n30020), .Z(n30013) );
  AND U29768 ( .A(n30021), .B(n30022), .Z(n30020) );
  XNOR U29769 ( .A(n30019), .B(n30023), .Z(n30021) );
  XNOR U29770 ( .A(n29979), .B(n29986), .Z(n30001) );
  AND U29771 ( .A(n29935), .B(n30024), .Z(n29986) );
  XOR U29772 ( .A(n29991), .B(n29990), .Z(n29979) );
  XNOR U29773 ( .A(n30025), .B(n29987), .Z(n29990) );
  XOR U29774 ( .A(n30026), .B(n30027), .Z(n29987) );
  AND U29775 ( .A(n30028), .B(n30029), .Z(n30027) );
  XOR U29776 ( .A(n30026), .B(n30030), .Z(n30028) );
  XNOR U29777 ( .A(n30031), .B(n30032), .Z(n30025) );
  AND U29778 ( .A(n30033), .B(n30034), .Z(n30032) );
  XOR U29779 ( .A(n30031), .B(n30035), .Z(n30033) );
  XOR U29780 ( .A(n30036), .B(n30037), .Z(n29991) );
  AND U29781 ( .A(n30038), .B(n30039), .Z(n30037) );
  XOR U29782 ( .A(n30036), .B(n30040), .Z(n30038) );
  XNOR U29783 ( .A(n29924), .B(n29997), .Z(n29999) );
  XNOR U29784 ( .A(n30041), .B(n30042), .Z(n29924) );
  AND U29785 ( .A(n230), .B(n30043), .Z(n30042) );
  XNOR U29786 ( .A(n30044), .B(n30045), .Z(n30043) );
  XOR U29787 ( .A(n30046), .B(n30047), .Z(n29997) );
  AND U29788 ( .A(n30048), .B(n30049), .Z(n30047) );
  XNOR U29789 ( .A(n30046), .B(n29935), .Z(n30049) );
  XOR U29790 ( .A(n30050), .B(n30011), .Z(n29935) );
  XNOR U29791 ( .A(n30051), .B(n30018), .Z(n30011) );
  XOR U29792 ( .A(n30007), .B(n30006), .Z(n30018) );
  XNOR U29793 ( .A(n30052), .B(n30003), .Z(n30006) );
  XOR U29794 ( .A(n30053), .B(n30054), .Z(n30003) );
  AND U29795 ( .A(n30055), .B(n30056), .Z(n30054) );
  XNOR U29796 ( .A(n30057), .B(n30058), .Z(n30055) );
  IV U29797 ( .A(n30053), .Z(n30057) );
  XNOR U29798 ( .A(n30059), .B(n30060), .Z(n30052) );
  NOR U29799 ( .A(n30061), .B(n30062), .Z(n30060) );
  XNOR U29800 ( .A(n30059), .B(n30063), .Z(n30061) );
  XOR U29801 ( .A(n30064), .B(n30065), .Z(n30007) );
  NOR U29802 ( .A(n30066), .B(n30067), .Z(n30065) );
  XNOR U29803 ( .A(n30064), .B(n30068), .Z(n30066) );
  XNOR U29804 ( .A(n30017), .B(n30008), .Z(n30051) );
  XOR U29805 ( .A(n30069), .B(n30070), .Z(n30008) );
  AND U29806 ( .A(n30071), .B(n30072), .Z(n30070) );
  XOR U29807 ( .A(n30069), .B(n30073), .Z(n30071) );
  XOR U29808 ( .A(n30074), .B(n30023), .Z(n30017) );
  XOR U29809 ( .A(n30075), .B(n30076), .Z(n30023) );
  NOR U29810 ( .A(n30077), .B(n30078), .Z(n30076) );
  XOR U29811 ( .A(n30075), .B(n30079), .Z(n30077) );
  XNOR U29812 ( .A(n30022), .B(n30014), .Z(n30074) );
  XOR U29813 ( .A(n30080), .B(n30081), .Z(n30014) );
  AND U29814 ( .A(n30082), .B(n30083), .Z(n30081) );
  XOR U29815 ( .A(n30080), .B(n30084), .Z(n30082) );
  XNOR U29816 ( .A(n30085), .B(n30019), .Z(n30022) );
  XOR U29817 ( .A(n30086), .B(n30087), .Z(n30019) );
  AND U29818 ( .A(n30088), .B(n30089), .Z(n30087) );
  XNOR U29819 ( .A(n30090), .B(n30091), .Z(n30088) );
  IV U29820 ( .A(n30086), .Z(n30090) );
  XNOR U29821 ( .A(n30092), .B(n30093), .Z(n30085) );
  NOR U29822 ( .A(n30094), .B(n30095), .Z(n30093) );
  XNOR U29823 ( .A(n30092), .B(n30096), .Z(n30094) );
  XOR U29824 ( .A(n30012), .B(n30024), .Z(n30050) );
  NOR U29825 ( .A(n29941), .B(n30097), .Z(n30024) );
  XNOR U29826 ( .A(n30030), .B(n30029), .Z(n30012) );
  XNOR U29827 ( .A(n30098), .B(n30035), .Z(n30029) );
  XNOR U29828 ( .A(n30099), .B(n30100), .Z(n30035) );
  NOR U29829 ( .A(n30101), .B(n30102), .Z(n30100) );
  XOR U29830 ( .A(n30099), .B(n30103), .Z(n30101) );
  XNOR U29831 ( .A(n30034), .B(n30026), .Z(n30098) );
  XOR U29832 ( .A(n30104), .B(n30105), .Z(n30026) );
  AND U29833 ( .A(n30106), .B(n30107), .Z(n30105) );
  XOR U29834 ( .A(n30104), .B(n30108), .Z(n30106) );
  XNOR U29835 ( .A(n30109), .B(n30031), .Z(n30034) );
  XOR U29836 ( .A(n30110), .B(n30111), .Z(n30031) );
  AND U29837 ( .A(n30112), .B(n30113), .Z(n30111) );
  XNOR U29838 ( .A(n30114), .B(n30115), .Z(n30112) );
  IV U29839 ( .A(n30110), .Z(n30114) );
  XNOR U29840 ( .A(n30116), .B(n30117), .Z(n30109) );
  NOR U29841 ( .A(n30118), .B(n30119), .Z(n30117) );
  XNOR U29842 ( .A(n30116), .B(n30120), .Z(n30118) );
  XOR U29843 ( .A(n30040), .B(n30039), .Z(n30030) );
  XNOR U29844 ( .A(n30121), .B(n30036), .Z(n30039) );
  XOR U29845 ( .A(n30122), .B(n30123), .Z(n30036) );
  AND U29846 ( .A(n30124), .B(n30125), .Z(n30123) );
  XNOR U29847 ( .A(n30126), .B(n30127), .Z(n30124) );
  IV U29848 ( .A(n30122), .Z(n30126) );
  XNOR U29849 ( .A(n30128), .B(n30129), .Z(n30121) );
  NOR U29850 ( .A(n30130), .B(n30131), .Z(n30129) );
  XNOR U29851 ( .A(n30128), .B(n30132), .Z(n30130) );
  XOR U29852 ( .A(n30133), .B(n30134), .Z(n30040) );
  NOR U29853 ( .A(n30135), .B(n30136), .Z(n30134) );
  XNOR U29854 ( .A(n30133), .B(n30137), .Z(n30135) );
  XNOR U29855 ( .A(n29932), .B(n30046), .Z(n30048) );
  XNOR U29856 ( .A(n30138), .B(n30139), .Z(n29932) );
  AND U29857 ( .A(n230), .B(n30140), .Z(n30139) );
  XNOR U29858 ( .A(n30141), .B(n30142), .Z(n30140) );
  AND U29859 ( .A(n29938), .B(n29941), .Z(n30046) );
  XOR U29860 ( .A(n30143), .B(n30097), .Z(n29941) );
  XNOR U29861 ( .A(p_input[160]), .B(p_input[2048]), .Z(n30097) );
  XNOR U29862 ( .A(n30073), .B(n30072), .Z(n30143) );
  XNOR U29863 ( .A(n30144), .B(n30084), .Z(n30072) );
  XOR U29864 ( .A(n30058), .B(n30056), .Z(n30084) );
  XNOR U29865 ( .A(n30145), .B(n30063), .Z(n30056) );
  XOR U29866 ( .A(p_input[184]), .B(p_input[2072]), .Z(n30063) );
  XOR U29867 ( .A(n30053), .B(n30062), .Z(n30145) );
  XOR U29868 ( .A(n30146), .B(n30059), .Z(n30062) );
  XOR U29869 ( .A(p_input[182]), .B(p_input[2070]), .Z(n30059) );
  XOR U29870 ( .A(p_input[183]), .B(n29410), .Z(n30146) );
  XOR U29871 ( .A(p_input[178]), .B(p_input[2066]), .Z(n30053) );
  XNOR U29872 ( .A(n30068), .B(n30067), .Z(n30058) );
  XOR U29873 ( .A(n30147), .B(n30064), .Z(n30067) );
  XOR U29874 ( .A(p_input[179]), .B(p_input[2067]), .Z(n30064) );
  XOR U29875 ( .A(p_input[180]), .B(n29412), .Z(n30147) );
  XOR U29876 ( .A(p_input[181]), .B(p_input[2069]), .Z(n30068) );
  XOR U29877 ( .A(n30083), .B(n30148), .Z(n30144) );
  IV U29878 ( .A(n30069), .Z(n30148) );
  XOR U29879 ( .A(p_input[161]), .B(p_input[2049]), .Z(n30069) );
  XNOR U29880 ( .A(n30149), .B(n30091), .Z(n30083) );
  XNOR U29881 ( .A(n30079), .B(n30078), .Z(n30091) );
  XNOR U29882 ( .A(n30150), .B(n30075), .Z(n30078) );
  XNOR U29883 ( .A(p_input[186]), .B(p_input[2074]), .Z(n30075) );
  XOR U29884 ( .A(p_input[187]), .B(n29415), .Z(n30150) );
  XOR U29885 ( .A(p_input[188]), .B(p_input[2076]), .Z(n30079) );
  XOR U29886 ( .A(n30089), .B(n30151), .Z(n30149) );
  IV U29887 ( .A(n30080), .Z(n30151) );
  XOR U29888 ( .A(p_input[177]), .B(p_input[2065]), .Z(n30080) );
  XNOR U29889 ( .A(n30152), .B(n30096), .Z(n30089) );
  XNOR U29890 ( .A(p_input[191]), .B(n29418), .Z(n30096) );
  XOR U29891 ( .A(n30086), .B(n30095), .Z(n30152) );
  XOR U29892 ( .A(n30153), .B(n30092), .Z(n30095) );
  XOR U29893 ( .A(p_input[189]), .B(p_input[2077]), .Z(n30092) );
  XOR U29894 ( .A(p_input[190]), .B(n29420), .Z(n30153) );
  XOR U29895 ( .A(p_input[185]), .B(p_input[2073]), .Z(n30086) );
  XOR U29896 ( .A(n30108), .B(n30107), .Z(n30073) );
  XNOR U29897 ( .A(n30154), .B(n30115), .Z(n30107) );
  XNOR U29898 ( .A(n30103), .B(n30102), .Z(n30115) );
  XNOR U29899 ( .A(n30155), .B(n30099), .Z(n30102) );
  XNOR U29900 ( .A(p_input[171]), .B(p_input[2059]), .Z(n30099) );
  XOR U29901 ( .A(p_input[172]), .B(n28329), .Z(n30155) );
  XOR U29902 ( .A(p_input[173]), .B(p_input[2061]), .Z(n30103) );
  XOR U29903 ( .A(n30113), .B(n30156), .Z(n30154) );
  IV U29904 ( .A(n30104), .Z(n30156) );
  XOR U29905 ( .A(p_input[162]), .B(p_input[2050]), .Z(n30104) );
  XNOR U29906 ( .A(n30157), .B(n30120), .Z(n30113) );
  XNOR U29907 ( .A(p_input[176]), .B(n28332), .Z(n30120) );
  XOR U29908 ( .A(n30110), .B(n30119), .Z(n30157) );
  XOR U29909 ( .A(n30158), .B(n30116), .Z(n30119) );
  XOR U29910 ( .A(p_input[174]), .B(p_input[2062]), .Z(n30116) );
  XOR U29911 ( .A(p_input[175]), .B(n28334), .Z(n30158) );
  XOR U29912 ( .A(p_input[170]), .B(p_input[2058]), .Z(n30110) );
  XOR U29913 ( .A(n30127), .B(n30125), .Z(n30108) );
  XNOR U29914 ( .A(n30159), .B(n30132), .Z(n30125) );
  XOR U29915 ( .A(p_input[169]), .B(p_input[2057]), .Z(n30132) );
  XOR U29916 ( .A(n30122), .B(n30131), .Z(n30159) );
  XOR U29917 ( .A(n30160), .B(n30128), .Z(n30131) );
  XOR U29918 ( .A(p_input[167]), .B(p_input[2055]), .Z(n30128) );
  XOR U29919 ( .A(p_input[168]), .B(n29427), .Z(n30160) );
  XOR U29920 ( .A(p_input[163]), .B(p_input[2051]), .Z(n30122) );
  XNOR U29921 ( .A(n30137), .B(n30136), .Z(n30127) );
  XOR U29922 ( .A(n30161), .B(n30133), .Z(n30136) );
  XOR U29923 ( .A(p_input[164]), .B(p_input[2052]), .Z(n30133) );
  XOR U29924 ( .A(p_input[165]), .B(n29429), .Z(n30161) );
  XOR U29925 ( .A(p_input[166]), .B(p_input[2054]), .Z(n30137) );
  XNOR U29926 ( .A(n30162), .B(n30163), .Z(n29938) );
  AND U29927 ( .A(n230), .B(n30164), .Z(n30163) );
  XNOR U29928 ( .A(n30165), .B(n30166), .Z(n230) );
  AND U29929 ( .A(n30167), .B(n30168), .Z(n30166) );
  XOR U29930 ( .A(n29952), .B(n30165), .Z(n30168) );
  XNOR U29931 ( .A(n30169), .B(n30165), .Z(n30167) );
  XOR U29932 ( .A(n30170), .B(n30171), .Z(n30165) );
  AND U29933 ( .A(n30172), .B(n30173), .Z(n30171) );
  XOR U29934 ( .A(n29967), .B(n30170), .Z(n30173) );
  XOR U29935 ( .A(n30170), .B(n29968), .Z(n30172) );
  XOR U29936 ( .A(n30174), .B(n30175), .Z(n30170) );
  AND U29937 ( .A(n30176), .B(n30177), .Z(n30175) );
  XOR U29938 ( .A(n29995), .B(n30174), .Z(n30177) );
  XOR U29939 ( .A(n30174), .B(n29996), .Z(n30176) );
  XOR U29940 ( .A(n30178), .B(n30179), .Z(n30174) );
  AND U29941 ( .A(n30180), .B(n30181), .Z(n30179) );
  XOR U29942 ( .A(n30044), .B(n30178), .Z(n30181) );
  XOR U29943 ( .A(n30178), .B(n30045), .Z(n30180) );
  XOR U29944 ( .A(n30182), .B(n30183), .Z(n30178) );
  AND U29945 ( .A(n30184), .B(n30185), .Z(n30183) );
  XOR U29946 ( .A(n30182), .B(n30141), .Z(n30185) );
  XNOR U29947 ( .A(n30186), .B(n30187), .Z(n29888) );
  AND U29948 ( .A(n234), .B(n30188), .Z(n30187) );
  XNOR U29949 ( .A(n30189), .B(n30190), .Z(n234) );
  AND U29950 ( .A(n30191), .B(n30192), .Z(n30190) );
  XOR U29951 ( .A(n30189), .B(n29898), .Z(n30192) );
  XNOR U29952 ( .A(n30189), .B(n29848), .Z(n30191) );
  XOR U29953 ( .A(n30193), .B(n30194), .Z(n30189) );
  AND U29954 ( .A(n30195), .B(n30196), .Z(n30194) );
  XNOR U29955 ( .A(n29908), .B(n30193), .Z(n30196) );
  XOR U29956 ( .A(n30193), .B(n29858), .Z(n30195) );
  XOR U29957 ( .A(n30197), .B(n30198), .Z(n30193) );
  AND U29958 ( .A(n30199), .B(n30200), .Z(n30198) );
  XNOR U29959 ( .A(n29918), .B(n30197), .Z(n30200) );
  XOR U29960 ( .A(n30197), .B(n29867), .Z(n30199) );
  XOR U29961 ( .A(n30201), .B(n30202), .Z(n30197) );
  AND U29962 ( .A(n30203), .B(n30204), .Z(n30202) );
  XOR U29963 ( .A(n30201), .B(n29875), .Z(n30203) );
  XOR U29964 ( .A(n30205), .B(n30206), .Z(n29839) );
  AND U29965 ( .A(n238), .B(n30188), .Z(n30206) );
  XNOR U29966 ( .A(n30186), .B(n30205), .Z(n30188) );
  XNOR U29967 ( .A(n30207), .B(n30208), .Z(n238) );
  AND U29968 ( .A(n30209), .B(n30210), .Z(n30208) );
  XNOR U29969 ( .A(n30211), .B(n30207), .Z(n30210) );
  IV U29970 ( .A(n29898), .Z(n30211) );
  XOR U29971 ( .A(n30169), .B(n30212), .Z(n29898) );
  AND U29972 ( .A(n241), .B(n30213), .Z(n30212) );
  XOR U29973 ( .A(n29951), .B(n29948), .Z(n30213) );
  IV U29974 ( .A(n30169), .Z(n29951) );
  XNOR U29975 ( .A(n29848), .B(n30207), .Z(n30209) );
  XOR U29976 ( .A(n30214), .B(n30215), .Z(n29848) );
  AND U29977 ( .A(n257), .B(n30216), .Z(n30215) );
  XOR U29978 ( .A(n30217), .B(n30218), .Z(n30207) );
  AND U29979 ( .A(n30219), .B(n30220), .Z(n30218) );
  XNOR U29980 ( .A(n30217), .B(n29908), .Z(n30220) );
  XOR U29981 ( .A(n29968), .B(n30221), .Z(n29908) );
  AND U29982 ( .A(n241), .B(n30222), .Z(n30221) );
  XOR U29983 ( .A(n29964), .B(n29968), .Z(n30222) );
  XNOR U29984 ( .A(n30223), .B(n30217), .Z(n30219) );
  IV U29985 ( .A(n29858), .Z(n30223) );
  XOR U29986 ( .A(n30224), .B(n30225), .Z(n29858) );
  AND U29987 ( .A(n257), .B(n30226), .Z(n30225) );
  XOR U29988 ( .A(n30227), .B(n30228), .Z(n30217) );
  AND U29989 ( .A(n30229), .B(n30230), .Z(n30228) );
  XNOR U29990 ( .A(n30227), .B(n29918), .Z(n30230) );
  XOR U29991 ( .A(n29996), .B(n30231), .Z(n29918) );
  AND U29992 ( .A(n241), .B(n30232), .Z(n30231) );
  XOR U29993 ( .A(n29992), .B(n29996), .Z(n30232) );
  XOR U29994 ( .A(n29867), .B(n30227), .Z(n30229) );
  XOR U29995 ( .A(n30233), .B(n30234), .Z(n29867) );
  AND U29996 ( .A(n257), .B(n30235), .Z(n30234) );
  XOR U29997 ( .A(n30201), .B(n30236), .Z(n30227) );
  AND U29998 ( .A(n30237), .B(n30204), .Z(n30236) );
  XNOR U29999 ( .A(n29928), .B(n30201), .Z(n30204) );
  XOR U30000 ( .A(n30045), .B(n30238), .Z(n29928) );
  AND U30001 ( .A(n241), .B(n30239), .Z(n30238) );
  XOR U30002 ( .A(n30041), .B(n30045), .Z(n30239) );
  XNOR U30003 ( .A(n30240), .B(n30201), .Z(n30237) );
  IV U30004 ( .A(n29875), .Z(n30240) );
  XOR U30005 ( .A(n30241), .B(n30242), .Z(n29875) );
  AND U30006 ( .A(n257), .B(n30243), .Z(n30242) );
  XOR U30007 ( .A(n30244), .B(n30245), .Z(n30201) );
  AND U30008 ( .A(n30246), .B(n30247), .Z(n30245) );
  XNOR U30009 ( .A(n30244), .B(n29936), .Z(n30247) );
  XOR U30010 ( .A(n30142), .B(n30248), .Z(n29936) );
  AND U30011 ( .A(n241), .B(n30249), .Z(n30248) );
  XOR U30012 ( .A(n30138), .B(n30142), .Z(n30249) );
  XNOR U30013 ( .A(n30250), .B(n30244), .Z(n30246) );
  IV U30014 ( .A(n29885), .Z(n30250) );
  XOR U30015 ( .A(n30251), .B(n30252), .Z(n29885) );
  AND U30016 ( .A(n257), .B(n30253), .Z(n30252) );
  AND U30017 ( .A(n30205), .B(n30186), .Z(n30244) );
  XNOR U30018 ( .A(n30254), .B(n30255), .Z(n30186) );
  AND U30019 ( .A(n241), .B(n30164), .Z(n30255) );
  XNOR U30020 ( .A(n30162), .B(n30254), .Z(n30164) );
  XNOR U30021 ( .A(n30256), .B(n30257), .Z(n241) );
  AND U30022 ( .A(n30258), .B(n30259), .Z(n30257) );
  XNOR U30023 ( .A(n30256), .B(n29948), .Z(n30259) );
  IV U30024 ( .A(n29952), .Z(n29948) );
  XOR U30025 ( .A(n30260), .B(n30261), .Z(n29952) );
  AND U30026 ( .A(n245), .B(n30262), .Z(n30261) );
  XOR U30027 ( .A(n30263), .B(n30260), .Z(n30262) );
  XNOR U30028 ( .A(n30256), .B(n30169), .Z(n30258) );
  XOR U30029 ( .A(n30264), .B(n30265), .Z(n30169) );
  AND U30030 ( .A(n253), .B(n30216), .Z(n30265) );
  XOR U30031 ( .A(n30214), .B(n30264), .Z(n30216) );
  XOR U30032 ( .A(n30266), .B(n30267), .Z(n30256) );
  AND U30033 ( .A(n30268), .B(n30269), .Z(n30267) );
  XNOR U30034 ( .A(n30266), .B(n29964), .Z(n30269) );
  IV U30035 ( .A(n29967), .Z(n29964) );
  XOR U30036 ( .A(n30270), .B(n30271), .Z(n29967) );
  AND U30037 ( .A(n245), .B(n30272), .Z(n30271) );
  XOR U30038 ( .A(n30273), .B(n30270), .Z(n30272) );
  XOR U30039 ( .A(n29968), .B(n30266), .Z(n30268) );
  XOR U30040 ( .A(n30274), .B(n30275), .Z(n29968) );
  AND U30041 ( .A(n253), .B(n30226), .Z(n30275) );
  XOR U30042 ( .A(n30274), .B(n30224), .Z(n30226) );
  XOR U30043 ( .A(n30276), .B(n30277), .Z(n30266) );
  AND U30044 ( .A(n30278), .B(n30279), .Z(n30277) );
  XNOR U30045 ( .A(n30276), .B(n29992), .Z(n30279) );
  IV U30046 ( .A(n29995), .Z(n29992) );
  XOR U30047 ( .A(n30280), .B(n30281), .Z(n29995) );
  AND U30048 ( .A(n245), .B(n30282), .Z(n30281) );
  XNOR U30049 ( .A(n30283), .B(n30280), .Z(n30282) );
  XOR U30050 ( .A(n29996), .B(n30276), .Z(n30278) );
  XOR U30051 ( .A(n30284), .B(n30285), .Z(n29996) );
  AND U30052 ( .A(n253), .B(n30235), .Z(n30285) );
  XOR U30053 ( .A(n30284), .B(n30233), .Z(n30235) );
  XOR U30054 ( .A(n30286), .B(n30287), .Z(n30276) );
  AND U30055 ( .A(n30288), .B(n30289), .Z(n30287) );
  XNOR U30056 ( .A(n30286), .B(n30041), .Z(n30289) );
  IV U30057 ( .A(n30044), .Z(n30041) );
  XOR U30058 ( .A(n30290), .B(n30291), .Z(n30044) );
  AND U30059 ( .A(n245), .B(n30292), .Z(n30291) );
  XOR U30060 ( .A(n30293), .B(n30290), .Z(n30292) );
  XOR U30061 ( .A(n30045), .B(n30286), .Z(n30288) );
  XOR U30062 ( .A(n30294), .B(n30295), .Z(n30045) );
  AND U30063 ( .A(n253), .B(n30243), .Z(n30295) );
  XOR U30064 ( .A(n30294), .B(n30241), .Z(n30243) );
  XOR U30065 ( .A(n30182), .B(n30296), .Z(n30286) );
  AND U30066 ( .A(n30184), .B(n30297), .Z(n30296) );
  XNOR U30067 ( .A(n30182), .B(n30138), .Z(n30297) );
  IV U30068 ( .A(n30141), .Z(n30138) );
  XOR U30069 ( .A(n30298), .B(n30299), .Z(n30141) );
  AND U30070 ( .A(n245), .B(n30300), .Z(n30299) );
  XNOR U30071 ( .A(n30301), .B(n30298), .Z(n30300) );
  XOR U30072 ( .A(n30142), .B(n30182), .Z(n30184) );
  XOR U30073 ( .A(n30302), .B(n30303), .Z(n30142) );
  AND U30074 ( .A(n253), .B(n30253), .Z(n30303) );
  XOR U30075 ( .A(n30302), .B(n30251), .Z(n30253) );
  AND U30076 ( .A(n30254), .B(n30162), .Z(n30182) );
  XNOR U30077 ( .A(n30304), .B(n30305), .Z(n30162) );
  AND U30078 ( .A(n245), .B(n30306), .Z(n30305) );
  XNOR U30079 ( .A(n30307), .B(n30304), .Z(n30306) );
  XNOR U30080 ( .A(n30308), .B(n30309), .Z(n245) );
  AND U30081 ( .A(n30310), .B(n30311), .Z(n30309) );
  XOR U30082 ( .A(n30263), .B(n30308), .Z(n30311) );
  AND U30083 ( .A(n30312), .B(n30313), .Z(n30263) );
  XNOR U30084 ( .A(n30260), .B(n30308), .Z(n30310) );
  XNOR U30085 ( .A(n30314), .B(n30315), .Z(n30260) );
  AND U30086 ( .A(n249), .B(n30316), .Z(n30315) );
  XNOR U30087 ( .A(n30317), .B(n30318), .Z(n30316) );
  XOR U30088 ( .A(n30319), .B(n30320), .Z(n30308) );
  AND U30089 ( .A(n30321), .B(n30322), .Z(n30320) );
  XNOR U30090 ( .A(n30319), .B(n30312), .Z(n30322) );
  IV U30091 ( .A(n30273), .Z(n30312) );
  XOR U30092 ( .A(n30323), .B(n30324), .Z(n30273) );
  XOR U30093 ( .A(n30325), .B(n30313), .Z(n30324) );
  AND U30094 ( .A(n30283), .B(n30326), .Z(n30313) );
  AND U30095 ( .A(n30327), .B(n30328), .Z(n30325) );
  XOR U30096 ( .A(n30329), .B(n30323), .Z(n30327) );
  XNOR U30097 ( .A(n30270), .B(n30319), .Z(n30321) );
  XNOR U30098 ( .A(n30330), .B(n30331), .Z(n30270) );
  AND U30099 ( .A(n249), .B(n30332), .Z(n30331) );
  XNOR U30100 ( .A(n30333), .B(n30334), .Z(n30332) );
  XOR U30101 ( .A(n30335), .B(n30336), .Z(n30319) );
  AND U30102 ( .A(n30337), .B(n30338), .Z(n30336) );
  XNOR U30103 ( .A(n30335), .B(n30283), .Z(n30338) );
  XOR U30104 ( .A(n30339), .B(n30328), .Z(n30283) );
  XNOR U30105 ( .A(n30340), .B(n30323), .Z(n30328) );
  XOR U30106 ( .A(n30341), .B(n30342), .Z(n30323) );
  AND U30107 ( .A(n30343), .B(n30344), .Z(n30342) );
  XOR U30108 ( .A(n30345), .B(n30341), .Z(n30343) );
  XNOR U30109 ( .A(n30346), .B(n30347), .Z(n30340) );
  AND U30110 ( .A(n30348), .B(n30349), .Z(n30347) );
  XOR U30111 ( .A(n30346), .B(n30350), .Z(n30348) );
  XNOR U30112 ( .A(n30329), .B(n30326), .Z(n30339) );
  AND U30113 ( .A(n30351), .B(n30352), .Z(n30326) );
  XOR U30114 ( .A(n30353), .B(n30354), .Z(n30329) );
  AND U30115 ( .A(n30355), .B(n30356), .Z(n30354) );
  XOR U30116 ( .A(n30353), .B(n30357), .Z(n30355) );
  XNOR U30117 ( .A(n30280), .B(n30335), .Z(n30337) );
  XNOR U30118 ( .A(n30358), .B(n30359), .Z(n30280) );
  AND U30119 ( .A(n249), .B(n30360), .Z(n30359) );
  XNOR U30120 ( .A(n30361), .B(n30362), .Z(n30360) );
  XOR U30121 ( .A(n30363), .B(n30364), .Z(n30335) );
  AND U30122 ( .A(n30365), .B(n30366), .Z(n30364) );
  XNOR U30123 ( .A(n30363), .B(n30351), .Z(n30366) );
  IV U30124 ( .A(n30293), .Z(n30351) );
  XNOR U30125 ( .A(n30367), .B(n30344), .Z(n30293) );
  XNOR U30126 ( .A(n30368), .B(n30350), .Z(n30344) );
  XOR U30127 ( .A(n30369), .B(n30370), .Z(n30350) );
  AND U30128 ( .A(n30371), .B(n30372), .Z(n30370) );
  XOR U30129 ( .A(n30369), .B(n30373), .Z(n30371) );
  XNOR U30130 ( .A(n30349), .B(n30341), .Z(n30368) );
  XOR U30131 ( .A(n30374), .B(n30375), .Z(n30341) );
  AND U30132 ( .A(n30376), .B(n30377), .Z(n30375) );
  XNOR U30133 ( .A(n30378), .B(n30374), .Z(n30376) );
  XNOR U30134 ( .A(n30379), .B(n30346), .Z(n30349) );
  XOR U30135 ( .A(n30380), .B(n30381), .Z(n30346) );
  AND U30136 ( .A(n30382), .B(n30383), .Z(n30381) );
  XOR U30137 ( .A(n30380), .B(n30384), .Z(n30382) );
  XNOR U30138 ( .A(n30385), .B(n30386), .Z(n30379) );
  AND U30139 ( .A(n30387), .B(n30388), .Z(n30386) );
  XNOR U30140 ( .A(n30385), .B(n30389), .Z(n30387) );
  XNOR U30141 ( .A(n30345), .B(n30352), .Z(n30367) );
  AND U30142 ( .A(n30301), .B(n30390), .Z(n30352) );
  XOR U30143 ( .A(n30357), .B(n30356), .Z(n30345) );
  XNOR U30144 ( .A(n30391), .B(n30353), .Z(n30356) );
  XOR U30145 ( .A(n30392), .B(n30393), .Z(n30353) );
  AND U30146 ( .A(n30394), .B(n30395), .Z(n30393) );
  XOR U30147 ( .A(n30392), .B(n30396), .Z(n30394) );
  XNOR U30148 ( .A(n30397), .B(n30398), .Z(n30391) );
  AND U30149 ( .A(n30399), .B(n30400), .Z(n30398) );
  XOR U30150 ( .A(n30397), .B(n30401), .Z(n30399) );
  XOR U30151 ( .A(n30402), .B(n30403), .Z(n30357) );
  AND U30152 ( .A(n30404), .B(n30405), .Z(n30403) );
  XOR U30153 ( .A(n30402), .B(n30406), .Z(n30404) );
  XNOR U30154 ( .A(n30290), .B(n30363), .Z(n30365) );
  XNOR U30155 ( .A(n30407), .B(n30408), .Z(n30290) );
  AND U30156 ( .A(n249), .B(n30409), .Z(n30408) );
  XNOR U30157 ( .A(n30410), .B(n30411), .Z(n30409) );
  XOR U30158 ( .A(n30412), .B(n30413), .Z(n30363) );
  AND U30159 ( .A(n30414), .B(n30415), .Z(n30413) );
  XNOR U30160 ( .A(n30412), .B(n30301), .Z(n30415) );
  XOR U30161 ( .A(n30416), .B(n30377), .Z(n30301) );
  XNOR U30162 ( .A(n30417), .B(n30384), .Z(n30377) );
  XOR U30163 ( .A(n30373), .B(n30372), .Z(n30384) );
  XNOR U30164 ( .A(n30418), .B(n30369), .Z(n30372) );
  XOR U30165 ( .A(n30419), .B(n30420), .Z(n30369) );
  AND U30166 ( .A(n30421), .B(n30422), .Z(n30420) );
  XOR U30167 ( .A(n30419), .B(n30423), .Z(n30421) );
  XNOR U30168 ( .A(n30424), .B(n30425), .Z(n30418) );
  NOR U30169 ( .A(n30426), .B(n30427), .Z(n30425) );
  XNOR U30170 ( .A(n30424), .B(n30428), .Z(n30426) );
  XOR U30171 ( .A(n30429), .B(n30430), .Z(n30373) );
  NOR U30172 ( .A(n30431), .B(n30432), .Z(n30430) );
  XNOR U30173 ( .A(n30429), .B(n30433), .Z(n30431) );
  XNOR U30174 ( .A(n30383), .B(n30374), .Z(n30417) );
  XOR U30175 ( .A(n30434), .B(n30435), .Z(n30374) );
  NOR U30176 ( .A(n30436), .B(n30437), .Z(n30435) );
  XOR U30177 ( .A(n30438), .B(n30439), .Z(n30436) );
  XOR U30178 ( .A(n30440), .B(n30389), .Z(n30383) );
  XNOR U30179 ( .A(n30441), .B(n30442), .Z(n30389) );
  NOR U30180 ( .A(n30443), .B(n30444), .Z(n30442) );
  XNOR U30181 ( .A(n30441), .B(n30445), .Z(n30443) );
  XNOR U30182 ( .A(n30388), .B(n30380), .Z(n30440) );
  XOR U30183 ( .A(n30446), .B(n30447), .Z(n30380) );
  AND U30184 ( .A(n30448), .B(n30449), .Z(n30447) );
  XOR U30185 ( .A(n30446), .B(n30450), .Z(n30448) );
  XNOR U30186 ( .A(n30451), .B(n30385), .Z(n30388) );
  XOR U30187 ( .A(n30452), .B(n30453), .Z(n30385) );
  AND U30188 ( .A(n30454), .B(n30455), .Z(n30453) );
  XOR U30189 ( .A(n30452), .B(n30456), .Z(n30454) );
  XNOR U30190 ( .A(n30457), .B(n30458), .Z(n30451) );
  NOR U30191 ( .A(n30459), .B(n30460), .Z(n30458) );
  XOR U30192 ( .A(n30457), .B(n30461), .Z(n30459) );
  XOR U30193 ( .A(n30378), .B(n30390), .Z(n30416) );
  NOR U30194 ( .A(n30307), .B(n30462), .Z(n30390) );
  XNOR U30195 ( .A(n30396), .B(n30395), .Z(n30378) );
  XNOR U30196 ( .A(n30463), .B(n30401), .Z(n30395) );
  XNOR U30197 ( .A(n30464), .B(n30465), .Z(n30401) );
  NOR U30198 ( .A(n30466), .B(n30467), .Z(n30465) );
  XOR U30199 ( .A(n30464), .B(n30468), .Z(n30466) );
  XNOR U30200 ( .A(n30400), .B(n30392), .Z(n30463) );
  XOR U30201 ( .A(n30469), .B(n30470), .Z(n30392) );
  AND U30202 ( .A(n30471), .B(n30472), .Z(n30470) );
  XOR U30203 ( .A(n30469), .B(n30473), .Z(n30471) );
  XNOR U30204 ( .A(n30474), .B(n30397), .Z(n30400) );
  XOR U30205 ( .A(n30475), .B(n30476), .Z(n30397) );
  AND U30206 ( .A(n30477), .B(n30478), .Z(n30476) );
  XNOR U30207 ( .A(n30479), .B(n30480), .Z(n30477) );
  IV U30208 ( .A(n30475), .Z(n30479) );
  XNOR U30209 ( .A(n30481), .B(n30482), .Z(n30474) );
  NOR U30210 ( .A(n30483), .B(n30484), .Z(n30482) );
  XOR U30211 ( .A(n30481), .B(n30485), .Z(n30483) );
  XOR U30212 ( .A(n30406), .B(n30405), .Z(n30396) );
  XNOR U30213 ( .A(n30486), .B(n30402), .Z(n30405) );
  XOR U30214 ( .A(n30487), .B(n30488), .Z(n30402) );
  AND U30215 ( .A(n30489), .B(n30490), .Z(n30488) );
  XNOR U30216 ( .A(n30491), .B(n30492), .Z(n30489) );
  IV U30217 ( .A(n30487), .Z(n30491) );
  XNOR U30218 ( .A(n30493), .B(n30494), .Z(n30486) );
  NOR U30219 ( .A(n30495), .B(n30496), .Z(n30494) );
  XNOR U30220 ( .A(n30493), .B(n30497), .Z(n30495) );
  XOR U30221 ( .A(n30498), .B(n30499), .Z(n30406) );
  NOR U30222 ( .A(n30500), .B(n30501), .Z(n30499) );
  XNOR U30223 ( .A(n30498), .B(n30502), .Z(n30500) );
  XNOR U30224 ( .A(n30298), .B(n30412), .Z(n30414) );
  XNOR U30225 ( .A(n30503), .B(n30504), .Z(n30298) );
  AND U30226 ( .A(n249), .B(n30505), .Z(n30504) );
  XNOR U30227 ( .A(n30506), .B(n30507), .Z(n30505) );
  AND U30228 ( .A(n30304), .B(n30307), .Z(n30412) );
  XOR U30229 ( .A(n30508), .B(n30462), .Z(n30307) );
  XNOR U30230 ( .A(p_input[192]), .B(p_input[2048]), .Z(n30462) );
  XOR U30231 ( .A(n30439), .B(n30437), .Z(n30508) );
  XOR U30232 ( .A(n30509), .B(n30450), .Z(n30437) );
  XOR U30233 ( .A(n30423), .B(n30422), .Z(n30450) );
  XNOR U30234 ( .A(n30510), .B(n30428), .Z(n30422) );
  XOR U30235 ( .A(p_input[2072]), .B(p_input[216]), .Z(n30428) );
  XOR U30236 ( .A(n30419), .B(n30427), .Z(n30510) );
  XOR U30237 ( .A(n30511), .B(n30424), .Z(n30427) );
  XOR U30238 ( .A(p_input[2070]), .B(p_input[214]), .Z(n30424) );
  XNOR U30239 ( .A(p_input[2071]), .B(p_input[215]), .Z(n30511) );
  XNOR U30240 ( .A(n28684), .B(p_input[210]), .Z(n30419) );
  XNOR U30241 ( .A(n30433), .B(n30432), .Z(n30423) );
  XOR U30242 ( .A(n30512), .B(n30429), .Z(n30432) );
  XOR U30243 ( .A(p_input[2067]), .B(p_input[211]), .Z(n30429) );
  XNOR U30244 ( .A(p_input[2068]), .B(p_input[212]), .Z(n30512) );
  XOR U30245 ( .A(p_input[2069]), .B(p_input[213]), .Z(n30433) );
  XOR U30246 ( .A(n30449), .B(n30438), .Z(n30509) );
  IV U30247 ( .A(n30434), .Z(n30438) );
  XOR U30248 ( .A(p_input[193]), .B(p_input[2049]), .Z(n30434) );
  XNOR U30249 ( .A(n30513), .B(n30456), .Z(n30449) );
  XNOR U30250 ( .A(n30445), .B(n30444), .Z(n30456) );
  XOR U30251 ( .A(n30514), .B(n30441), .Z(n30444) );
  XNOR U30252 ( .A(n28322), .B(p_input[218]), .Z(n30441) );
  XNOR U30253 ( .A(p_input[2075]), .B(p_input[219]), .Z(n30514) );
  XOR U30254 ( .A(p_input[2076]), .B(p_input[220]), .Z(n30445) );
  XNOR U30255 ( .A(n30455), .B(n30446), .Z(n30513) );
  XNOR U30256 ( .A(n28689), .B(p_input[209]), .Z(n30446) );
  XOR U30257 ( .A(n30515), .B(n30461), .Z(n30455) );
  XNOR U30258 ( .A(p_input[2079]), .B(p_input[223]), .Z(n30461) );
  XOR U30259 ( .A(n30452), .B(n30460), .Z(n30515) );
  XOR U30260 ( .A(n30516), .B(n30457), .Z(n30460) );
  XOR U30261 ( .A(p_input[2077]), .B(p_input[221]), .Z(n30457) );
  XNOR U30262 ( .A(p_input[2078]), .B(p_input[222]), .Z(n30516) );
  XNOR U30263 ( .A(n28326), .B(p_input[217]), .Z(n30452) );
  XOR U30264 ( .A(n30473), .B(n30472), .Z(n30439) );
  XNOR U30265 ( .A(n30517), .B(n30480), .Z(n30472) );
  XNOR U30266 ( .A(n30468), .B(n30467), .Z(n30480) );
  XNOR U30267 ( .A(n30518), .B(n30464), .Z(n30467) );
  XNOR U30268 ( .A(p_input[203]), .B(p_input[2059]), .Z(n30464) );
  XOR U30269 ( .A(p_input[204]), .B(n28329), .Z(n30518) );
  XOR U30270 ( .A(p_input[205]), .B(p_input[2061]), .Z(n30468) );
  XOR U30271 ( .A(n30478), .B(n30519), .Z(n30517) );
  IV U30272 ( .A(n30469), .Z(n30519) );
  XOR U30273 ( .A(p_input[194]), .B(p_input[2050]), .Z(n30469) );
  XOR U30274 ( .A(n30520), .B(n30485), .Z(n30478) );
  XNOR U30275 ( .A(p_input[2064]), .B(p_input[208]), .Z(n30485) );
  XOR U30276 ( .A(n30475), .B(n30484), .Z(n30520) );
  XOR U30277 ( .A(n30521), .B(n30481), .Z(n30484) );
  XOR U30278 ( .A(p_input[2062]), .B(p_input[206]), .Z(n30481) );
  XNOR U30279 ( .A(p_input[2063]), .B(p_input[207]), .Z(n30521) );
  XOR U30280 ( .A(p_input[202]), .B(p_input[2058]), .Z(n30475) );
  XOR U30281 ( .A(n30492), .B(n30490), .Z(n30473) );
  XNOR U30282 ( .A(n30522), .B(n30497), .Z(n30490) );
  XOR U30283 ( .A(p_input[201]), .B(p_input[2057]), .Z(n30497) );
  XOR U30284 ( .A(n30487), .B(n30496), .Z(n30522) );
  XOR U30285 ( .A(n30523), .B(n30493), .Z(n30496) );
  XOR U30286 ( .A(p_input[199]), .B(p_input[2055]), .Z(n30493) );
  XOR U30287 ( .A(p_input[200]), .B(n29427), .Z(n30523) );
  XOR U30288 ( .A(p_input[195]), .B(p_input[2051]), .Z(n30487) );
  XNOR U30289 ( .A(n30502), .B(n30501), .Z(n30492) );
  XOR U30290 ( .A(n30524), .B(n30498), .Z(n30501) );
  XOR U30291 ( .A(p_input[196]), .B(p_input[2052]), .Z(n30498) );
  XOR U30292 ( .A(p_input[197]), .B(n29429), .Z(n30524) );
  XOR U30293 ( .A(p_input[198]), .B(p_input[2054]), .Z(n30502) );
  XNOR U30294 ( .A(n30525), .B(n30526), .Z(n30304) );
  AND U30295 ( .A(n249), .B(n30527), .Z(n30526) );
  XNOR U30296 ( .A(n30528), .B(n30529), .Z(n249) );
  AND U30297 ( .A(n30530), .B(n30531), .Z(n30529) );
  XOR U30298 ( .A(n30318), .B(n30528), .Z(n30531) );
  XNOR U30299 ( .A(n30532), .B(n30528), .Z(n30530) );
  XOR U30300 ( .A(n30533), .B(n30534), .Z(n30528) );
  AND U30301 ( .A(n30535), .B(n30536), .Z(n30534) );
  XOR U30302 ( .A(n30333), .B(n30533), .Z(n30536) );
  XOR U30303 ( .A(n30533), .B(n30334), .Z(n30535) );
  XOR U30304 ( .A(n30537), .B(n30538), .Z(n30533) );
  AND U30305 ( .A(n30539), .B(n30540), .Z(n30538) );
  XOR U30306 ( .A(n30361), .B(n30537), .Z(n30540) );
  XOR U30307 ( .A(n30537), .B(n30362), .Z(n30539) );
  XOR U30308 ( .A(n30541), .B(n30542), .Z(n30537) );
  AND U30309 ( .A(n30543), .B(n30544), .Z(n30542) );
  XOR U30310 ( .A(n30410), .B(n30541), .Z(n30544) );
  XOR U30311 ( .A(n30541), .B(n30411), .Z(n30543) );
  XOR U30312 ( .A(n30545), .B(n30546), .Z(n30541) );
  AND U30313 ( .A(n30547), .B(n30548), .Z(n30546) );
  XOR U30314 ( .A(n30545), .B(n30506), .Z(n30548) );
  XNOR U30315 ( .A(n30549), .B(n30550), .Z(n30254) );
  AND U30316 ( .A(n253), .B(n30551), .Z(n30550) );
  XNOR U30317 ( .A(n30552), .B(n30553), .Z(n253) );
  AND U30318 ( .A(n30554), .B(n30555), .Z(n30553) );
  XOR U30319 ( .A(n30552), .B(n30264), .Z(n30555) );
  XNOR U30320 ( .A(n30552), .B(n30214), .Z(n30554) );
  XOR U30321 ( .A(n30556), .B(n30557), .Z(n30552) );
  AND U30322 ( .A(n30558), .B(n30559), .Z(n30557) );
  XNOR U30323 ( .A(n30274), .B(n30556), .Z(n30559) );
  XOR U30324 ( .A(n30556), .B(n30224), .Z(n30558) );
  XOR U30325 ( .A(n30560), .B(n30561), .Z(n30556) );
  AND U30326 ( .A(n30562), .B(n30563), .Z(n30561) );
  XNOR U30327 ( .A(n30284), .B(n30560), .Z(n30563) );
  XOR U30328 ( .A(n30560), .B(n30233), .Z(n30562) );
  XOR U30329 ( .A(n30564), .B(n30565), .Z(n30560) );
  AND U30330 ( .A(n30566), .B(n30567), .Z(n30565) );
  XOR U30331 ( .A(n30564), .B(n30241), .Z(n30566) );
  XOR U30332 ( .A(n30568), .B(n30569), .Z(n30205) );
  AND U30333 ( .A(n257), .B(n30551), .Z(n30569) );
  XNOR U30334 ( .A(n30549), .B(n30568), .Z(n30551) );
  XNOR U30335 ( .A(n30570), .B(n30571), .Z(n257) );
  AND U30336 ( .A(n30572), .B(n30573), .Z(n30571) );
  XNOR U30337 ( .A(n30574), .B(n30570), .Z(n30573) );
  IV U30338 ( .A(n30264), .Z(n30574) );
  XOR U30339 ( .A(n30532), .B(n30575), .Z(n30264) );
  AND U30340 ( .A(n260), .B(n30576), .Z(n30575) );
  XOR U30341 ( .A(n30317), .B(n30314), .Z(n30576) );
  IV U30342 ( .A(n30532), .Z(n30317) );
  XNOR U30343 ( .A(n30214), .B(n30570), .Z(n30572) );
  XOR U30344 ( .A(n30577), .B(n30578), .Z(n30214) );
  AND U30345 ( .A(n276), .B(n30579), .Z(n30578) );
  XOR U30346 ( .A(n30580), .B(n30581), .Z(n30570) );
  AND U30347 ( .A(n30582), .B(n30583), .Z(n30581) );
  XNOR U30348 ( .A(n30580), .B(n30274), .Z(n30583) );
  XOR U30349 ( .A(n30334), .B(n30584), .Z(n30274) );
  AND U30350 ( .A(n260), .B(n30585), .Z(n30584) );
  XOR U30351 ( .A(n30330), .B(n30334), .Z(n30585) );
  XNOR U30352 ( .A(n30586), .B(n30580), .Z(n30582) );
  IV U30353 ( .A(n30224), .Z(n30586) );
  XOR U30354 ( .A(n30587), .B(n30588), .Z(n30224) );
  AND U30355 ( .A(n276), .B(n30589), .Z(n30588) );
  XOR U30356 ( .A(n30590), .B(n30591), .Z(n30580) );
  AND U30357 ( .A(n30592), .B(n30593), .Z(n30591) );
  XNOR U30358 ( .A(n30590), .B(n30284), .Z(n30593) );
  XOR U30359 ( .A(n30362), .B(n30594), .Z(n30284) );
  AND U30360 ( .A(n260), .B(n30595), .Z(n30594) );
  XOR U30361 ( .A(n30358), .B(n30362), .Z(n30595) );
  XOR U30362 ( .A(n30233), .B(n30590), .Z(n30592) );
  XOR U30363 ( .A(n30596), .B(n30597), .Z(n30233) );
  AND U30364 ( .A(n276), .B(n30598), .Z(n30597) );
  XOR U30365 ( .A(n30564), .B(n30599), .Z(n30590) );
  AND U30366 ( .A(n30600), .B(n30567), .Z(n30599) );
  XNOR U30367 ( .A(n30294), .B(n30564), .Z(n30567) );
  XOR U30368 ( .A(n30411), .B(n30601), .Z(n30294) );
  AND U30369 ( .A(n260), .B(n30602), .Z(n30601) );
  XOR U30370 ( .A(n30407), .B(n30411), .Z(n30602) );
  XNOR U30371 ( .A(n30603), .B(n30564), .Z(n30600) );
  IV U30372 ( .A(n30241), .Z(n30603) );
  XOR U30373 ( .A(n30604), .B(n30605), .Z(n30241) );
  AND U30374 ( .A(n276), .B(n30606), .Z(n30605) );
  XOR U30375 ( .A(n30607), .B(n30608), .Z(n30564) );
  AND U30376 ( .A(n30609), .B(n30610), .Z(n30608) );
  XNOR U30377 ( .A(n30607), .B(n30302), .Z(n30610) );
  XOR U30378 ( .A(n30507), .B(n30611), .Z(n30302) );
  AND U30379 ( .A(n260), .B(n30612), .Z(n30611) );
  XOR U30380 ( .A(n30503), .B(n30507), .Z(n30612) );
  XNOR U30381 ( .A(n30613), .B(n30607), .Z(n30609) );
  IV U30382 ( .A(n30251), .Z(n30613) );
  XOR U30383 ( .A(n30614), .B(n30615), .Z(n30251) );
  AND U30384 ( .A(n276), .B(n30616), .Z(n30615) );
  AND U30385 ( .A(n30568), .B(n30549), .Z(n30607) );
  XNOR U30386 ( .A(n30617), .B(n30618), .Z(n30549) );
  AND U30387 ( .A(n260), .B(n30527), .Z(n30618) );
  XNOR U30388 ( .A(n30525), .B(n30617), .Z(n30527) );
  XNOR U30389 ( .A(n30619), .B(n30620), .Z(n260) );
  AND U30390 ( .A(n30621), .B(n30622), .Z(n30620) );
  XNOR U30391 ( .A(n30619), .B(n30314), .Z(n30622) );
  IV U30392 ( .A(n30318), .Z(n30314) );
  XOR U30393 ( .A(n30623), .B(n30624), .Z(n30318) );
  AND U30394 ( .A(n264), .B(n30625), .Z(n30624) );
  XOR U30395 ( .A(n30626), .B(n30623), .Z(n30625) );
  XNOR U30396 ( .A(n30619), .B(n30532), .Z(n30621) );
  XOR U30397 ( .A(n30627), .B(n30628), .Z(n30532) );
  AND U30398 ( .A(n272), .B(n30579), .Z(n30628) );
  XOR U30399 ( .A(n30577), .B(n30627), .Z(n30579) );
  XOR U30400 ( .A(n30629), .B(n30630), .Z(n30619) );
  AND U30401 ( .A(n30631), .B(n30632), .Z(n30630) );
  XNOR U30402 ( .A(n30629), .B(n30330), .Z(n30632) );
  IV U30403 ( .A(n30333), .Z(n30330) );
  XOR U30404 ( .A(n30633), .B(n30634), .Z(n30333) );
  AND U30405 ( .A(n264), .B(n30635), .Z(n30634) );
  XOR U30406 ( .A(n30636), .B(n30633), .Z(n30635) );
  XOR U30407 ( .A(n30334), .B(n30629), .Z(n30631) );
  XOR U30408 ( .A(n30637), .B(n30638), .Z(n30334) );
  AND U30409 ( .A(n272), .B(n30589), .Z(n30638) );
  XOR U30410 ( .A(n30637), .B(n30587), .Z(n30589) );
  XOR U30411 ( .A(n30639), .B(n30640), .Z(n30629) );
  AND U30412 ( .A(n30641), .B(n30642), .Z(n30640) );
  XNOR U30413 ( .A(n30639), .B(n30358), .Z(n30642) );
  IV U30414 ( .A(n30361), .Z(n30358) );
  XOR U30415 ( .A(n30643), .B(n30644), .Z(n30361) );
  AND U30416 ( .A(n264), .B(n30645), .Z(n30644) );
  XNOR U30417 ( .A(n30646), .B(n30643), .Z(n30645) );
  XOR U30418 ( .A(n30362), .B(n30639), .Z(n30641) );
  XOR U30419 ( .A(n30647), .B(n30648), .Z(n30362) );
  AND U30420 ( .A(n272), .B(n30598), .Z(n30648) );
  XOR U30421 ( .A(n30647), .B(n30596), .Z(n30598) );
  XOR U30422 ( .A(n30649), .B(n30650), .Z(n30639) );
  AND U30423 ( .A(n30651), .B(n30652), .Z(n30650) );
  XNOR U30424 ( .A(n30649), .B(n30407), .Z(n30652) );
  IV U30425 ( .A(n30410), .Z(n30407) );
  XOR U30426 ( .A(n30653), .B(n30654), .Z(n30410) );
  AND U30427 ( .A(n264), .B(n30655), .Z(n30654) );
  XOR U30428 ( .A(n30656), .B(n30653), .Z(n30655) );
  XOR U30429 ( .A(n30411), .B(n30649), .Z(n30651) );
  XOR U30430 ( .A(n30657), .B(n30658), .Z(n30411) );
  AND U30431 ( .A(n272), .B(n30606), .Z(n30658) );
  XOR U30432 ( .A(n30657), .B(n30604), .Z(n30606) );
  XOR U30433 ( .A(n30545), .B(n30659), .Z(n30649) );
  AND U30434 ( .A(n30547), .B(n30660), .Z(n30659) );
  XNOR U30435 ( .A(n30545), .B(n30503), .Z(n30660) );
  IV U30436 ( .A(n30506), .Z(n30503) );
  XOR U30437 ( .A(n30661), .B(n30662), .Z(n30506) );
  AND U30438 ( .A(n264), .B(n30663), .Z(n30662) );
  XNOR U30439 ( .A(n30664), .B(n30661), .Z(n30663) );
  XOR U30440 ( .A(n30507), .B(n30545), .Z(n30547) );
  XOR U30441 ( .A(n30665), .B(n30666), .Z(n30507) );
  AND U30442 ( .A(n272), .B(n30616), .Z(n30666) );
  XOR U30443 ( .A(n30665), .B(n30614), .Z(n30616) );
  AND U30444 ( .A(n30617), .B(n30525), .Z(n30545) );
  XNOR U30445 ( .A(n30667), .B(n30668), .Z(n30525) );
  AND U30446 ( .A(n264), .B(n30669), .Z(n30668) );
  XNOR U30447 ( .A(n30670), .B(n30667), .Z(n30669) );
  XNOR U30448 ( .A(n30671), .B(n30672), .Z(n264) );
  AND U30449 ( .A(n30673), .B(n30674), .Z(n30672) );
  XOR U30450 ( .A(n30626), .B(n30671), .Z(n30674) );
  AND U30451 ( .A(n30675), .B(n30676), .Z(n30626) );
  XNOR U30452 ( .A(n30623), .B(n30671), .Z(n30673) );
  XNOR U30453 ( .A(n30677), .B(n30678), .Z(n30623) );
  AND U30454 ( .A(n268), .B(n30679), .Z(n30678) );
  XNOR U30455 ( .A(n30680), .B(n30681), .Z(n30679) );
  XOR U30456 ( .A(n30682), .B(n30683), .Z(n30671) );
  AND U30457 ( .A(n30684), .B(n30685), .Z(n30683) );
  XNOR U30458 ( .A(n30682), .B(n30675), .Z(n30685) );
  IV U30459 ( .A(n30636), .Z(n30675) );
  XOR U30460 ( .A(n30686), .B(n30687), .Z(n30636) );
  XOR U30461 ( .A(n30688), .B(n30676), .Z(n30687) );
  AND U30462 ( .A(n30646), .B(n30689), .Z(n30676) );
  AND U30463 ( .A(n30690), .B(n30691), .Z(n30688) );
  XOR U30464 ( .A(n30692), .B(n30686), .Z(n30690) );
  XNOR U30465 ( .A(n30633), .B(n30682), .Z(n30684) );
  XNOR U30466 ( .A(n30693), .B(n30694), .Z(n30633) );
  AND U30467 ( .A(n268), .B(n30695), .Z(n30694) );
  XNOR U30468 ( .A(n30696), .B(n30697), .Z(n30695) );
  XOR U30469 ( .A(n30698), .B(n30699), .Z(n30682) );
  AND U30470 ( .A(n30700), .B(n30701), .Z(n30699) );
  XNOR U30471 ( .A(n30698), .B(n30646), .Z(n30701) );
  XOR U30472 ( .A(n30702), .B(n30691), .Z(n30646) );
  XNOR U30473 ( .A(n30703), .B(n30686), .Z(n30691) );
  XOR U30474 ( .A(n30704), .B(n30705), .Z(n30686) );
  AND U30475 ( .A(n30706), .B(n30707), .Z(n30705) );
  XOR U30476 ( .A(n30708), .B(n30704), .Z(n30706) );
  XNOR U30477 ( .A(n30709), .B(n30710), .Z(n30703) );
  AND U30478 ( .A(n30711), .B(n30712), .Z(n30710) );
  XOR U30479 ( .A(n30709), .B(n30713), .Z(n30711) );
  XNOR U30480 ( .A(n30692), .B(n30689), .Z(n30702) );
  AND U30481 ( .A(n30714), .B(n30715), .Z(n30689) );
  XOR U30482 ( .A(n30716), .B(n30717), .Z(n30692) );
  AND U30483 ( .A(n30718), .B(n30719), .Z(n30717) );
  XOR U30484 ( .A(n30716), .B(n30720), .Z(n30718) );
  XNOR U30485 ( .A(n30643), .B(n30698), .Z(n30700) );
  XNOR U30486 ( .A(n30721), .B(n30722), .Z(n30643) );
  AND U30487 ( .A(n268), .B(n30723), .Z(n30722) );
  XNOR U30488 ( .A(n30724), .B(n30725), .Z(n30723) );
  XOR U30489 ( .A(n30726), .B(n30727), .Z(n30698) );
  AND U30490 ( .A(n30728), .B(n30729), .Z(n30727) );
  XNOR U30491 ( .A(n30726), .B(n30714), .Z(n30729) );
  IV U30492 ( .A(n30656), .Z(n30714) );
  XNOR U30493 ( .A(n30730), .B(n30707), .Z(n30656) );
  XNOR U30494 ( .A(n30731), .B(n30713), .Z(n30707) );
  XOR U30495 ( .A(n30732), .B(n30733), .Z(n30713) );
  AND U30496 ( .A(n30734), .B(n30735), .Z(n30733) );
  XOR U30497 ( .A(n30732), .B(n30736), .Z(n30734) );
  XNOR U30498 ( .A(n30712), .B(n30704), .Z(n30731) );
  XOR U30499 ( .A(n30737), .B(n30738), .Z(n30704) );
  AND U30500 ( .A(n30739), .B(n30740), .Z(n30738) );
  XNOR U30501 ( .A(n30741), .B(n30737), .Z(n30739) );
  XNOR U30502 ( .A(n30742), .B(n30709), .Z(n30712) );
  XOR U30503 ( .A(n30743), .B(n30744), .Z(n30709) );
  AND U30504 ( .A(n30745), .B(n30746), .Z(n30744) );
  XOR U30505 ( .A(n30743), .B(n30747), .Z(n30745) );
  XNOR U30506 ( .A(n30748), .B(n30749), .Z(n30742) );
  AND U30507 ( .A(n30750), .B(n30751), .Z(n30749) );
  XNOR U30508 ( .A(n30748), .B(n30752), .Z(n30750) );
  XNOR U30509 ( .A(n30708), .B(n30715), .Z(n30730) );
  AND U30510 ( .A(n30664), .B(n30753), .Z(n30715) );
  XOR U30511 ( .A(n30720), .B(n30719), .Z(n30708) );
  XNOR U30512 ( .A(n30754), .B(n30716), .Z(n30719) );
  XOR U30513 ( .A(n30755), .B(n30756), .Z(n30716) );
  AND U30514 ( .A(n30757), .B(n30758), .Z(n30756) );
  XOR U30515 ( .A(n30755), .B(n30759), .Z(n30757) );
  XNOR U30516 ( .A(n30760), .B(n30761), .Z(n30754) );
  AND U30517 ( .A(n30762), .B(n30763), .Z(n30761) );
  XOR U30518 ( .A(n30760), .B(n30764), .Z(n30762) );
  XOR U30519 ( .A(n30765), .B(n30766), .Z(n30720) );
  AND U30520 ( .A(n30767), .B(n30768), .Z(n30766) );
  XOR U30521 ( .A(n30765), .B(n30769), .Z(n30767) );
  XNOR U30522 ( .A(n30653), .B(n30726), .Z(n30728) );
  XNOR U30523 ( .A(n30770), .B(n30771), .Z(n30653) );
  AND U30524 ( .A(n268), .B(n30772), .Z(n30771) );
  XNOR U30525 ( .A(n30773), .B(n30774), .Z(n30772) );
  XOR U30526 ( .A(n30775), .B(n30776), .Z(n30726) );
  AND U30527 ( .A(n30777), .B(n30778), .Z(n30776) );
  XNOR U30528 ( .A(n30775), .B(n30664), .Z(n30778) );
  XOR U30529 ( .A(n30779), .B(n30740), .Z(n30664) );
  XNOR U30530 ( .A(n30780), .B(n30747), .Z(n30740) );
  XOR U30531 ( .A(n30736), .B(n30735), .Z(n30747) );
  XNOR U30532 ( .A(n30781), .B(n30732), .Z(n30735) );
  XOR U30533 ( .A(n30782), .B(n30783), .Z(n30732) );
  AND U30534 ( .A(n30784), .B(n30785), .Z(n30783) );
  XOR U30535 ( .A(n30782), .B(n30786), .Z(n30784) );
  XNOR U30536 ( .A(n30787), .B(n30788), .Z(n30781) );
  NOR U30537 ( .A(n30789), .B(n30790), .Z(n30788) );
  XNOR U30538 ( .A(n30787), .B(n30791), .Z(n30789) );
  XOR U30539 ( .A(n30792), .B(n30793), .Z(n30736) );
  NOR U30540 ( .A(n30794), .B(n30795), .Z(n30793) );
  XNOR U30541 ( .A(n30792), .B(n30796), .Z(n30794) );
  XNOR U30542 ( .A(n30746), .B(n30737), .Z(n30780) );
  XOR U30543 ( .A(n30797), .B(n30798), .Z(n30737) );
  NOR U30544 ( .A(n30799), .B(n30800), .Z(n30798) );
  XNOR U30545 ( .A(n30797), .B(n30801), .Z(n30799) );
  XOR U30546 ( .A(n30802), .B(n30752), .Z(n30746) );
  XNOR U30547 ( .A(n30803), .B(n30804), .Z(n30752) );
  NOR U30548 ( .A(n30805), .B(n30806), .Z(n30804) );
  XNOR U30549 ( .A(n30803), .B(n30807), .Z(n30805) );
  XNOR U30550 ( .A(n30751), .B(n30743), .Z(n30802) );
  XOR U30551 ( .A(n30808), .B(n30809), .Z(n30743) );
  AND U30552 ( .A(n30810), .B(n30811), .Z(n30809) );
  XOR U30553 ( .A(n30808), .B(n30812), .Z(n30810) );
  XNOR U30554 ( .A(n30813), .B(n30748), .Z(n30751) );
  XOR U30555 ( .A(n30814), .B(n30815), .Z(n30748) );
  AND U30556 ( .A(n30816), .B(n30817), .Z(n30815) );
  XOR U30557 ( .A(n30814), .B(n30818), .Z(n30816) );
  XNOR U30558 ( .A(n30819), .B(n30820), .Z(n30813) );
  NOR U30559 ( .A(n30821), .B(n30822), .Z(n30820) );
  XOR U30560 ( .A(n30819), .B(n30823), .Z(n30821) );
  XOR U30561 ( .A(n30741), .B(n30753), .Z(n30779) );
  NOR U30562 ( .A(n30670), .B(n30824), .Z(n30753) );
  XNOR U30563 ( .A(n30759), .B(n30758), .Z(n30741) );
  XNOR U30564 ( .A(n30825), .B(n30764), .Z(n30758) );
  XOR U30565 ( .A(n30826), .B(n30827), .Z(n30764) );
  NOR U30566 ( .A(n30828), .B(n30829), .Z(n30827) );
  XNOR U30567 ( .A(n30826), .B(n30830), .Z(n30828) );
  XNOR U30568 ( .A(n30763), .B(n30755), .Z(n30825) );
  XOR U30569 ( .A(n30831), .B(n30832), .Z(n30755) );
  AND U30570 ( .A(n30833), .B(n30834), .Z(n30832) );
  XNOR U30571 ( .A(n30831), .B(n30835), .Z(n30833) );
  XNOR U30572 ( .A(n30836), .B(n30760), .Z(n30763) );
  XOR U30573 ( .A(n30837), .B(n30838), .Z(n30760) );
  AND U30574 ( .A(n30839), .B(n30840), .Z(n30838) );
  XOR U30575 ( .A(n30837), .B(n30841), .Z(n30839) );
  XNOR U30576 ( .A(n30842), .B(n30843), .Z(n30836) );
  NOR U30577 ( .A(n30844), .B(n30845), .Z(n30843) );
  XOR U30578 ( .A(n30842), .B(n30846), .Z(n30844) );
  XOR U30579 ( .A(n30769), .B(n30768), .Z(n30759) );
  XNOR U30580 ( .A(n30847), .B(n30765), .Z(n30768) );
  XOR U30581 ( .A(n30848), .B(n30849), .Z(n30765) );
  AND U30582 ( .A(n30850), .B(n30851), .Z(n30849) );
  XOR U30583 ( .A(n30848), .B(n30852), .Z(n30850) );
  XNOR U30584 ( .A(n30853), .B(n30854), .Z(n30847) );
  NOR U30585 ( .A(n30855), .B(n30856), .Z(n30854) );
  XNOR U30586 ( .A(n30853), .B(n30857), .Z(n30855) );
  XOR U30587 ( .A(n30858), .B(n30859), .Z(n30769) );
  NOR U30588 ( .A(n30860), .B(n30861), .Z(n30859) );
  XNOR U30589 ( .A(n30858), .B(n30862), .Z(n30860) );
  XNOR U30590 ( .A(n30661), .B(n30775), .Z(n30777) );
  XNOR U30591 ( .A(n30863), .B(n30864), .Z(n30661) );
  AND U30592 ( .A(n268), .B(n30865), .Z(n30864) );
  XNOR U30593 ( .A(n30866), .B(n30867), .Z(n30865) );
  AND U30594 ( .A(n30667), .B(n30670), .Z(n30775) );
  XOR U30595 ( .A(n30868), .B(n30824), .Z(n30670) );
  XNOR U30596 ( .A(p_input[2048]), .B(p_input[224]), .Z(n30824) );
  XOR U30597 ( .A(n30801), .B(n30800), .Z(n30868) );
  XOR U30598 ( .A(n30869), .B(n30812), .Z(n30800) );
  XOR U30599 ( .A(n30786), .B(n30785), .Z(n30812) );
  XNOR U30600 ( .A(n30870), .B(n30791), .Z(n30785) );
  XOR U30601 ( .A(p_input[2072]), .B(p_input[248]), .Z(n30791) );
  XOR U30602 ( .A(n30782), .B(n30790), .Z(n30870) );
  XOR U30603 ( .A(n30871), .B(n30787), .Z(n30790) );
  XOR U30604 ( .A(p_input[2070]), .B(p_input[246]), .Z(n30787) );
  XNOR U30605 ( .A(p_input[2071]), .B(p_input[247]), .Z(n30871) );
  XNOR U30606 ( .A(n28684), .B(p_input[242]), .Z(n30782) );
  XNOR U30607 ( .A(n30796), .B(n30795), .Z(n30786) );
  XOR U30608 ( .A(n30872), .B(n30792), .Z(n30795) );
  XOR U30609 ( .A(p_input[2067]), .B(p_input[243]), .Z(n30792) );
  XNOR U30610 ( .A(p_input[2068]), .B(p_input[244]), .Z(n30872) );
  XOR U30611 ( .A(p_input[2069]), .B(p_input[245]), .Z(n30796) );
  XNOR U30612 ( .A(n30811), .B(n30797), .Z(n30869) );
  XNOR U30613 ( .A(n28686), .B(p_input[225]), .Z(n30797) );
  XNOR U30614 ( .A(n30873), .B(n30818), .Z(n30811) );
  XNOR U30615 ( .A(n30807), .B(n30806), .Z(n30818) );
  XOR U30616 ( .A(n30874), .B(n30803), .Z(n30806) );
  XNOR U30617 ( .A(n28322), .B(p_input[250]), .Z(n30803) );
  XNOR U30618 ( .A(p_input[2075]), .B(p_input[251]), .Z(n30874) );
  XOR U30619 ( .A(p_input[2076]), .B(p_input[252]), .Z(n30807) );
  XNOR U30620 ( .A(n30817), .B(n30808), .Z(n30873) );
  XNOR U30621 ( .A(n28689), .B(p_input[241]), .Z(n30808) );
  XOR U30622 ( .A(n30875), .B(n30823), .Z(n30817) );
  XNOR U30623 ( .A(p_input[2079]), .B(p_input[255]), .Z(n30823) );
  XOR U30624 ( .A(n30814), .B(n30822), .Z(n30875) );
  XOR U30625 ( .A(n30876), .B(n30819), .Z(n30822) );
  XOR U30626 ( .A(p_input[2077]), .B(p_input[253]), .Z(n30819) );
  XNOR U30627 ( .A(p_input[2078]), .B(p_input[254]), .Z(n30876) );
  XNOR U30628 ( .A(n28326), .B(p_input[249]), .Z(n30814) );
  XNOR U30629 ( .A(n30835), .B(n30834), .Z(n30801) );
  XNOR U30630 ( .A(n30877), .B(n30841), .Z(n30834) );
  XNOR U30631 ( .A(n30830), .B(n30829), .Z(n30841) );
  XOR U30632 ( .A(n30878), .B(n30826), .Z(n30829) );
  XNOR U30633 ( .A(n28694), .B(p_input[235]), .Z(n30826) );
  XNOR U30634 ( .A(p_input[2060]), .B(p_input[236]), .Z(n30878) );
  XOR U30635 ( .A(p_input[2061]), .B(p_input[237]), .Z(n30830) );
  XNOR U30636 ( .A(n30840), .B(n30831), .Z(n30877) );
  XNOR U30637 ( .A(n28330), .B(p_input[226]), .Z(n30831) );
  XOR U30638 ( .A(n30879), .B(n30846), .Z(n30840) );
  XNOR U30639 ( .A(p_input[2064]), .B(p_input[240]), .Z(n30846) );
  XOR U30640 ( .A(n30837), .B(n30845), .Z(n30879) );
  XOR U30641 ( .A(n30880), .B(n30842), .Z(n30845) );
  XOR U30642 ( .A(p_input[2062]), .B(p_input[238]), .Z(n30842) );
  XNOR U30643 ( .A(p_input[2063]), .B(p_input[239]), .Z(n30880) );
  XNOR U30644 ( .A(n28697), .B(p_input[234]), .Z(n30837) );
  XNOR U30645 ( .A(n30852), .B(n30851), .Z(n30835) );
  XNOR U30646 ( .A(n30881), .B(n30857), .Z(n30851) );
  XOR U30647 ( .A(p_input[2057]), .B(p_input[233]), .Z(n30857) );
  XOR U30648 ( .A(n30848), .B(n30856), .Z(n30881) );
  XOR U30649 ( .A(n30882), .B(n30853), .Z(n30856) );
  XOR U30650 ( .A(p_input[2055]), .B(p_input[231]), .Z(n30853) );
  XNOR U30651 ( .A(p_input[2056]), .B(p_input[232]), .Z(n30882) );
  XNOR U30652 ( .A(n28337), .B(p_input[227]), .Z(n30848) );
  XNOR U30653 ( .A(n30862), .B(n30861), .Z(n30852) );
  XOR U30654 ( .A(n30883), .B(n30858), .Z(n30861) );
  XOR U30655 ( .A(p_input[2052]), .B(p_input[228]), .Z(n30858) );
  XNOR U30656 ( .A(p_input[2053]), .B(p_input[229]), .Z(n30883) );
  XOR U30657 ( .A(p_input[2054]), .B(p_input[230]), .Z(n30862) );
  XNOR U30658 ( .A(n30884), .B(n30885), .Z(n30667) );
  AND U30659 ( .A(n268), .B(n30886), .Z(n30885) );
  XNOR U30660 ( .A(n30887), .B(n30888), .Z(n268) );
  AND U30661 ( .A(n30889), .B(n30890), .Z(n30888) );
  XOR U30662 ( .A(n30681), .B(n30887), .Z(n30890) );
  XNOR U30663 ( .A(n30891), .B(n30887), .Z(n30889) );
  XOR U30664 ( .A(n30892), .B(n30893), .Z(n30887) );
  AND U30665 ( .A(n30894), .B(n30895), .Z(n30893) );
  XOR U30666 ( .A(n30696), .B(n30892), .Z(n30895) );
  XOR U30667 ( .A(n30892), .B(n30697), .Z(n30894) );
  XOR U30668 ( .A(n30896), .B(n30897), .Z(n30892) );
  AND U30669 ( .A(n30898), .B(n30899), .Z(n30897) );
  XOR U30670 ( .A(n30724), .B(n30896), .Z(n30899) );
  XOR U30671 ( .A(n30896), .B(n30725), .Z(n30898) );
  XOR U30672 ( .A(n30900), .B(n30901), .Z(n30896) );
  AND U30673 ( .A(n30902), .B(n30903), .Z(n30901) );
  XOR U30674 ( .A(n30773), .B(n30900), .Z(n30903) );
  XOR U30675 ( .A(n30900), .B(n30774), .Z(n30902) );
  XOR U30676 ( .A(n30904), .B(n30905), .Z(n30900) );
  AND U30677 ( .A(n30906), .B(n30907), .Z(n30905) );
  XOR U30678 ( .A(n30904), .B(n30866), .Z(n30907) );
  XNOR U30679 ( .A(n30908), .B(n30909), .Z(n30617) );
  AND U30680 ( .A(n272), .B(n30910), .Z(n30909) );
  XNOR U30681 ( .A(n30911), .B(n30912), .Z(n272) );
  AND U30682 ( .A(n30913), .B(n30914), .Z(n30912) );
  XOR U30683 ( .A(n30911), .B(n30627), .Z(n30914) );
  XNOR U30684 ( .A(n30911), .B(n30577), .Z(n30913) );
  XOR U30685 ( .A(n30915), .B(n30916), .Z(n30911) );
  AND U30686 ( .A(n30917), .B(n30918), .Z(n30916) );
  XNOR U30687 ( .A(n30637), .B(n30915), .Z(n30918) );
  XOR U30688 ( .A(n30915), .B(n30587), .Z(n30917) );
  XOR U30689 ( .A(n30919), .B(n30920), .Z(n30915) );
  AND U30690 ( .A(n30921), .B(n30922), .Z(n30920) );
  XNOR U30691 ( .A(n30647), .B(n30919), .Z(n30922) );
  XOR U30692 ( .A(n30919), .B(n30596), .Z(n30921) );
  XOR U30693 ( .A(n30923), .B(n30924), .Z(n30919) );
  AND U30694 ( .A(n30925), .B(n30926), .Z(n30924) );
  XOR U30695 ( .A(n30923), .B(n30604), .Z(n30925) );
  XOR U30696 ( .A(n30927), .B(n30928), .Z(n30568) );
  AND U30697 ( .A(n276), .B(n30910), .Z(n30928) );
  XNOR U30698 ( .A(n30908), .B(n30927), .Z(n30910) );
  XNOR U30699 ( .A(n30929), .B(n30930), .Z(n276) );
  AND U30700 ( .A(n30931), .B(n30932), .Z(n30930) );
  XNOR U30701 ( .A(n30933), .B(n30929), .Z(n30932) );
  IV U30702 ( .A(n30627), .Z(n30933) );
  XOR U30703 ( .A(n30891), .B(n30934), .Z(n30627) );
  AND U30704 ( .A(n279), .B(n30935), .Z(n30934) );
  XOR U30705 ( .A(n30680), .B(n30677), .Z(n30935) );
  IV U30706 ( .A(n30891), .Z(n30680) );
  XNOR U30707 ( .A(n30577), .B(n30929), .Z(n30931) );
  XOR U30708 ( .A(n30936), .B(n30937), .Z(n30577) );
  AND U30709 ( .A(n295), .B(n30938), .Z(n30937) );
  XOR U30710 ( .A(n30939), .B(n30940), .Z(n30929) );
  AND U30711 ( .A(n30941), .B(n30942), .Z(n30940) );
  XNOR U30712 ( .A(n30939), .B(n30637), .Z(n30942) );
  XOR U30713 ( .A(n30697), .B(n30943), .Z(n30637) );
  AND U30714 ( .A(n279), .B(n30944), .Z(n30943) );
  XOR U30715 ( .A(n30693), .B(n30697), .Z(n30944) );
  XNOR U30716 ( .A(n30945), .B(n30939), .Z(n30941) );
  IV U30717 ( .A(n30587), .Z(n30945) );
  XOR U30718 ( .A(n30946), .B(n30947), .Z(n30587) );
  AND U30719 ( .A(n295), .B(n30948), .Z(n30947) );
  XOR U30720 ( .A(n30949), .B(n30950), .Z(n30939) );
  AND U30721 ( .A(n30951), .B(n30952), .Z(n30950) );
  XNOR U30722 ( .A(n30949), .B(n30647), .Z(n30952) );
  XOR U30723 ( .A(n30725), .B(n30953), .Z(n30647) );
  AND U30724 ( .A(n279), .B(n30954), .Z(n30953) );
  XOR U30725 ( .A(n30721), .B(n30725), .Z(n30954) );
  XOR U30726 ( .A(n30596), .B(n30949), .Z(n30951) );
  XOR U30727 ( .A(n30955), .B(n30956), .Z(n30596) );
  AND U30728 ( .A(n295), .B(n30957), .Z(n30956) );
  XOR U30729 ( .A(n30923), .B(n30958), .Z(n30949) );
  AND U30730 ( .A(n30959), .B(n30926), .Z(n30958) );
  XNOR U30731 ( .A(n30657), .B(n30923), .Z(n30926) );
  XOR U30732 ( .A(n30774), .B(n30960), .Z(n30657) );
  AND U30733 ( .A(n279), .B(n30961), .Z(n30960) );
  XOR U30734 ( .A(n30770), .B(n30774), .Z(n30961) );
  XNOR U30735 ( .A(n30962), .B(n30923), .Z(n30959) );
  IV U30736 ( .A(n30604), .Z(n30962) );
  XOR U30737 ( .A(n30963), .B(n30964), .Z(n30604) );
  AND U30738 ( .A(n295), .B(n30965), .Z(n30964) );
  XOR U30739 ( .A(n30966), .B(n30967), .Z(n30923) );
  AND U30740 ( .A(n30968), .B(n30969), .Z(n30967) );
  XNOR U30741 ( .A(n30966), .B(n30665), .Z(n30969) );
  XOR U30742 ( .A(n30867), .B(n30970), .Z(n30665) );
  AND U30743 ( .A(n279), .B(n30971), .Z(n30970) );
  XOR U30744 ( .A(n30863), .B(n30867), .Z(n30971) );
  XNOR U30745 ( .A(n30972), .B(n30966), .Z(n30968) );
  IV U30746 ( .A(n30614), .Z(n30972) );
  XOR U30747 ( .A(n30973), .B(n30974), .Z(n30614) );
  AND U30748 ( .A(n295), .B(n30975), .Z(n30974) );
  AND U30749 ( .A(n30927), .B(n30908), .Z(n30966) );
  XNOR U30750 ( .A(n30976), .B(n30977), .Z(n30908) );
  AND U30751 ( .A(n279), .B(n30886), .Z(n30977) );
  XNOR U30752 ( .A(n30884), .B(n30976), .Z(n30886) );
  XNOR U30753 ( .A(n30978), .B(n30979), .Z(n279) );
  AND U30754 ( .A(n30980), .B(n30981), .Z(n30979) );
  XNOR U30755 ( .A(n30978), .B(n30677), .Z(n30981) );
  IV U30756 ( .A(n30681), .Z(n30677) );
  XOR U30757 ( .A(n30982), .B(n30983), .Z(n30681) );
  AND U30758 ( .A(n283), .B(n30984), .Z(n30983) );
  XOR U30759 ( .A(n30985), .B(n30982), .Z(n30984) );
  XNOR U30760 ( .A(n30978), .B(n30891), .Z(n30980) );
  XOR U30761 ( .A(n30986), .B(n30987), .Z(n30891) );
  AND U30762 ( .A(n291), .B(n30938), .Z(n30987) );
  XOR U30763 ( .A(n30936), .B(n30986), .Z(n30938) );
  XOR U30764 ( .A(n30988), .B(n30989), .Z(n30978) );
  AND U30765 ( .A(n30990), .B(n30991), .Z(n30989) );
  XNOR U30766 ( .A(n30988), .B(n30693), .Z(n30991) );
  IV U30767 ( .A(n30696), .Z(n30693) );
  XOR U30768 ( .A(n30992), .B(n30993), .Z(n30696) );
  AND U30769 ( .A(n283), .B(n30994), .Z(n30993) );
  XOR U30770 ( .A(n30995), .B(n30992), .Z(n30994) );
  XOR U30771 ( .A(n30697), .B(n30988), .Z(n30990) );
  XOR U30772 ( .A(n30996), .B(n30997), .Z(n30697) );
  AND U30773 ( .A(n291), .B(n30948), .Z(n30997) );
  XOR U30774 ( .A(n30996), .B(n30946), .Z(n30948) );
  XOR U30775 ( .A(n30998), .B(n30999), .Z(n30988) );
  AND U30776 ( .A(n31000), .B(n31001), .Z(n30999) );
  XNOR U30777 ( .A(n30998), .B(n30721), .Z(n31001) );
  IV U30778 ( .A(n30724), .Z(n30721) );
  XOR U30779 ( .A(n31002), .B(n31003), .Z(n30724) );
  AND U30780 ( .A(n283), .B(n31004), .Z(n31003) );
  XNOR U30781 ( .A(n31005), .B(n31002), .Z(n31004) );
  XOR U30782 ( .A(n30725), .B(n30998), .Z(n31000) );
  XOR U30783 ( .A(n31006), .B(n31007), .Z(n30725) );
  AND U30784 ( .A(n291), .B(n30957), .Z(n31007) );
  XOR U30785 ( .A(n31006), .B(n30955), .Z(n30957) );
  XOR U30786 ( .A(n31008), .B(n31009), .Z(n30998) );
  AND U30787 ( .A(n31010), .B(n31011), .Z(n31009) );
  XNOR U30788 ( .A(n31008), .B(n30770), .Z(n31011) );
  IV U30789 ( .A(n30773), .Z(n30770) );
  XOR U30790 ( .A(n31012), .B(n31013), .Z(n30773) );
  AND U30791 ( .A(n283), .B(n31014), .Z(n31013) );
  XOR U30792 ( .A(n31015), .B(n31012), .Z(n31014) );
  XOR U30793 ( .A(n30774), .B(n31008), .Z(n31010) );
  XOR U30794 ( .A(n31016), .B(n31017), .Z(n30774) );
  AND U30795 ( .A(n291), .B(n30965), .Z(n31017) );
  XOR U30796 ( .A(n31016), .B(n30963), .Z(n30965) );
  XOR U30797 ( .A(n30904), .B(n31018), .Z(n31008) );
  AND U30798 ( .A(n30906), .B(n31019), .Z(n31018) );
  XNOR U30799 ( .A(n30904), .B(n30863), .Z(n31019) );
  IV U30800 ( .A(n30866), .Z(n30863) );
  XOR U30801 ( .A(n31020), .B(n31021), .Z(n30866) );
  AND U30802 ( .A(n283), .B(n31022), .Z(n31021) );
  XNOR U30803 ( .A(n31023), .B(n31020), .Z(n31022) );
  XOR U30804 ( .A(n30867), .B(n30904), .Z(n30906) );
  XOR U30805 ( .A(n31024), .B(n31025), .Z(n30867) );
  AND U30806 ( .A(n291), .B(n30975), .Z(n31025) );
  XOR U30807 ( .A(n31024), .B(n30973), .Z(n30975) );
  AND U30808 ( .A(n30976), .B(n30884), .Z(n30904) );
  XNOR U30809 ( .A(n31026), .B(n31027), .Z(n30884) );
  AND U30810 ( .A(n283), .B(n31028), .Z(n31027) );
  XNOR U30811 ( .A(n31029), .B(n31026), .Z(n31028) );
  XNOR U30812 ( .A(n31030), .B(n31031), .Z(n283) );
  AND U30813 ( .A(n31032), .B(n31033), .Z(n31031) );
  XOR U30814 ( .A(n30985), .B(n31030), .Z(n31033) );
  AND U30815 ( .A(n31034), .B(n31035), .Z(n30985) );
  XNOR U30816 ( .A(n30982), .B(n31030), .Z(n31032) );
  XNOR U30817 ( .A(n31036), .B(n31037), .Z(n30982) );
  AND U30818 ( .A(n287), .B(n31038), .Z(n31037) );
  XNOR U30819 ( .A(n31039), .B(n31040), .Z(n31038) );
  XOR U30820 ( .A(n31041), .B(n31042), .Z(n31030) );
  AND U30821 ( .A(n31043), .B(n31044), .Z(n31042) );
  XNOR U30822 ( .A(n31041), .B(n31034), .Z(n31044) );
  IV U30823 ( .A(n30995), .Z(n31034) );
  XOR U30824 ( .A(n31045), .B(n31046), .Z(n30995) );
  XOR U30825 ( .A(n31047), .B(n31035), .Z(n31046) );
  AND U30826 ( .A(n31005), .B(n31048), .Z(n31035) );
  AND U30827 ( .A(n31049), .B(n31050), .Z(n31047) );
  XOR U30828 ( .A(n31051), .B(n31045), .Z(n31049) );
  XNOR U30829 ( .A(n30992), .B(n31041), .Z(n31043) );
  XNOR U30830 ( .A(n31052), .B(n31053), .Z(n30992) );
  AND U30831 ( .A(n287), .B(n31054), .Z(n31053) );
  XNOR U30832 ( .A(n31055), .B(n31056), .Z(n31054) );
  XOR U30833 ( .A(n31057), .B(n31058), .Z(n31041) );
  AND U30834 ( .A(n31059), .B(n31060), .Z(n31058) );
  XNOR U30835 ( .A(n31057), .B(n31005), .Z(n31060) );
  XOR U30836 ( .A(n31061), .B(n31050), .Z(n31005) );
  XNOR U30837 ( .A(n31062), .B(n31045), .Z(n31050) );
  XOR U30838 ( .A(n31063), .B(n31064), .Z(n31045) );
  AND U30839 ( .A(n31065), .B(n31066), .Z(n31064) );
  XOR U30840 ( .A(n31067), .B(n31063), .Z(n31065) );
  XNOR U30841 ( .A(n31068), .B(n31069), .Z(n31062) );
  AND U30842 ( .A(n31070), .B(n31071), .Z(n31069) );
  XOR U30843 ( .A(n31068), .B(n31072), .Z(n31070) );
  XNOR U30844 ( .A(n31051), .B(n31048), .Z(n31061) );
  AND U30845 ( .A(n31073), .B(n31074), .Z(n31048) );
  XOR U30846 ( .A(n31075), .B(n31076), .Z(n31051) );
  AND U30847 ( .A(n31077), .B(n31078), .Z(n31076) );
  XOR U30848 ( .A(n31075), .B(n31079), .Z(n31077) );
  XNOR U30849 ( .A(n31002), .B(n31057), .Z(n31059) );
  XNOR U30850 ( .A(n31080), .B(n31081), .Z(n31002) );
  AND U30851 ( .A(n287), .B(n31082), .Z(n31081) );
  XNOR U30852 ( .A(n31083), .B(n31084), .Z(n31082) );
  XOR U30853 ( .A(n31085), .B(n31086), .Z(n31057) );
  AND U30854 ( .A(n31087), .B(n31088), .Z(n31086) );
  XNOR U30855 ( .A(n31085), .B(n31073), .Z(n31088) );
  IV U30856 ( .A(n31015), .Z(n31073) );
  XNOR U30857 ( .A(n31089), .B(n31066), .Z(n31015) );
  XNOR U30858 ( .A(n31090), .B(n31072), .Z(n31066) );
  XOR U30859 ( .A(n31091), .B(n31092), .Z(n31072) );
  AND U30860 ( .A(n31093), .B(n31094), .Z(n31092) );
  XOR U30861 ( .A(n31091), .B(n31095), .Z(n31093) );
  XNOR U30862 ( .A(n31071), .B(n31063), .Z(n31090) );
  XOR U30863 ( .A(n31096), .B(n31097), .Z(n31063) );
  AND U30864 ( .A(n31098), .B(n31099), .Z(n31097) );
  XNOR U30865 ( .A(n31100), .B(n31096), .Z(n31098) );
  XNOR U30866 ( .A(n31101), .B(n31068), .Z(n31071) );
  XOR U30867 ( .A(n31102), .B(n31103), .Z(n31068) );
  AND U30868 ( .A(n31104), .B(n31105), .Z(n31103) );
  XOR U30869 ( .A(n31102), .B(n31106), .Z(n31104) );
  XNOR U30870 ( .A(n31107), .B(n31108), .Z(n31101) );
  AND U30871 ( .A(n31109), .B(n31110), .Z(n31108) );
  XNOR U30872 ( .A(n31107), .B(n31111), .Z(n31109) );
  XNOR U30873 ( .A(n31067), .B(n31074), .Z(n31089) );
  AND U30874 ( .A(n31023), .B(n31112), .Z(n31074) );
  XOR U30875 ( .A(n31079), .B(n31078), .Z(n31067) );
  XNOR U30876 ( .A(n31113), .B(n31075), .Z(n31078) );
  XOR U30877 ( .A(n31114), .B(n31115), .Z(n31075) );
  AND U30878 ( .A(n31116), .B(n31117), .Z(n31115) );
  XOR U30879 ( .A(n31114), .B(n31118), .Z(n31116) );
  XNOR U30880 ( .A(n31119), .B(n31120), .Z(n31113) );
  AND U30881 ( .A(n31121), .B(n31122), .Z(n31120) );
  XOR U30882 ( .A(n31119), .B(n31123), .Z(n31121) );
  XOR U30883 ( .A(n31124), .B(n31125), .Z(n31079) );
  AND U30884 ( .A(n31126), .B(n31127), .Z(n31125) );
  XOR U30885 ( .A(n31124), .B(n31128), .Z(n31126) );
  XNOR U30886 ( .A(n31012), .B(n31085), .Z(n31087) );
  XNOR U30887 ( .A(n31129), .B(n31130), .Z(n31012) );
  AND U30888 ( .A(n287), .B(n31131), .Z(n31130) );
  XNOR U30889 ( .A(n31132), .B(n31133), .Z(n31131) );
  XOR U30890 ( .A(n31134), .B(n31135), .Z(n31085) );
  AND U30891 ( .A(n31136), .B(n31137), .Z(n31135) );
  XNOR U30892 ( .A(n31134), .B(n31023), .Z(n31137) );
  XOR U30893 ( .A(n31138), .B(n31099), .Z(n31023) );
  XNOR U30894 ( .A(n31139), .B(n31106), .Z(n31099) );
  XOR U30895 ( .A(n31095), .B(n31094), .Z(n31106) );
  XNOR U30896 ( .A(n31140), .B(n31091), .Z(n31094) );
  XOR U30897 ( .A(n31141), .B(n31142), .Z(n31091) );
  AND U30898 ( .A(n31143), .B(n31144), .Z(n31142) );
  XOR U30899 ( .A(n31141), .B(n31145), .Z(n31143) );
  XNOR U30900 ( .A(n31146), .B(n31147), .Z(n31140) );
  NOR U30901 ( .A(n31148), .B(n31149), .Z(n31147) );
  XNOR U30902 ( .A(n31146), .B(n31150), .Z(n31148) );
  XOR U30903 ( .A(n31151), .B(n31152), .Z(n31095) );
  NOR U30904 ( .A(n31153), .B(n31154), .Z(n31152) );
  XNOR U30905 ( .A(n31151), .B(n31155), .Z(n31153) );
  XNOR U30906 ( .A(n31105), .B(n31096), .Z(n31139) );
  XOR U30907 ( .A(n31156), .B(n31157), .Z(n31096) );
  NOR U30908 ( .A(n31158), .B(n31159), .Z(n31157) );
  XNOR U30909 ( .A(n31156), .B(n31160), .Z(n31158) );
  XOR U30910 ( .A(n31161), .B(n31111), .Z(n31105) );
  XNOR U30911 ( .A(n31162), .B(n31163), .Z(n31111) );
  NOR U30912 ( .A(n31164), .B(n31165), .Z(n31163) );
  XNOR U30913 ( .A(n31162), .B(n31166), .Z(n31164) );
  XNOR U30914 ( .A(n31110), .B(n31102), .Z(n31161) );
  XOR U30915 ( .A(n31167), .B(n31168), .Z(n31102) );
  AND U30916 ( .A(n31169), .B(n31170), .Z(n31168) );
  XOR U30917 ( .A(n31167), .B(n31171), .Z(n31169) );
  XNOR U30918 ( .A(n31172), .B(n31107), .Z(n31110) );
  XOR U30919 ( .A(n31173), .B(n31174), .Z(n31107) );
  AND U30920 ( .A(n31175), .B(n31176), .Z(n31174) );
  XOR U30921 ( .A(n31173), .B(n31177), .Z(n31175) );
  XNOR U30922 ( .A(n31178), .B(n31179), .Z(n31172) );
  NOR U30923 ( .A(n31180), .B(n31181), .Z(n31179) );
  XOR U30924 ( .A(n31178), .B(n31182), .Z(n31180) );
  XOR U30925 ( .A(n31100), .B(n31112), .Z(n31138) );
  NOR U30926 ( .A(n31029), .B(n31183), .Z(n31112) );
  XNOR U30927 ( .A(n31118), .B(n31117), .Z(n31100) );
  XNOR U30928 ( .A(n31184), .B(n31123), .Z(n31117) );
  XOR U30929 ( .A(n31185), .B(n31186), .Z(n31123) );
  NOR U30930 ( .A(n31187), .B(n31188), .Z(n31186) );
  XNOR U30931 ( .A(n31185), .B(n31189), .Z(n31187) );
  XNOR U30932 ( .A(n31122), .B(n31114), .Z(n31184) );
  XOR U30933 ( .A(n31190), .B(n31191), .Z(n31114) );
  AND U30934 ( .A(n31192), .B(n31193), .Z(n31191) );
  XNOR U30935 ( .A(n31190), .B(n31194), .Z(n31192) );
  XNOR U30936 ( .A(n31195), .B(n31119), .Z(n31122) );
  XOR U30937 ( .A(n31196), .B(n31197), .Z(n31119) );
  AND U30938 ( .A(n31198), .B(n31199), .Z(n31197) );
  XOR U30939 ( .A(n31196), .B(n31200), .Z(n31198) );
  XNOR U30940 ( .A(n31201), .B(n31202), .Z(n31195) );
  NOR U30941 ( .A(n31203), .B(n31204), .Z(n31202) );
  XOR U30942 ( .A(n31201), .B(n31205), .Z(n31203) );
  XOR U30943 ( .A(n31128), .B(n31127), .Z(n31118) );
  XNOR U30944 ( .A(n31206), .B(n31124), .Z(n31127) );
  XOR U30945 ( .A(n31207), .B(n31208), .Z(n31124) );
  AND U30946 ( .A(n31209), .B(n31210), .Z(n31208) );
  XOR U30947 ( .A(n31207), .B(n31211), .Z(n31209) );
  XNOR U30948 ( .A(n31212), .B(n31213), .Z(n31206) );
  NOR U30949 ( .A(n31214), .B(n31215), .Z(n31213) );
  XNOR U30950 ( .A(n31212), .B(n31216), .Z(n31214) );
  XOR U30951 ( .A(n31217), .B(n31218), .Z(n31128) );
  NOR U30952 ( .A(n31219), .B(n31220), .Z(n31218) );
  XNOR U30953 ( .A(n31217), .B(n31221), .Z(n31219) );
  XNOR U30954 ( .A(n31020), .B(n31134), .Z(n31136) );
  XNOR U30955 ( .A(n31222), .B(n31223), .Z(n31020) );
  AND U30956 ( .A(n287), .B(n31224), .Z(n31223) );
  XNOR U30957 ( .A(n31225), .B(n31226), .Z(n31224) );
  AND U30958 ( .A(n31026), .B(n31029), .Z(n31134) );
  XOR U30959 ( .A(n31227), .B(n31183), .Z(n31029) );
  XNOR U30960 ( .A(p_input[2048]), .B(p_input[256]), .Z(n31183) );
  XOR U30961 ( .A(n31160), .B(n31159), .Z(n31227) );
  XOR U30962 ( .A(n31228), .B(n31171), .Z(n31159) );
  XOR U30963 ( .A(n31145), .B(n31144), .Z(n31171) );
  XNOR U30964 ( .A(n31229), .B(n31150), .Z(n31144) );
  XOR U30965 ( .A(p_input[2072]), .B(p_input[280]), .Z(n31150) );
  XOR U30966 ( .A(n31141), .B(n31149), .Z(n31229) );
  XOR U30967 ( .A(n31230), .B(n31146), .Z(n31149) );
  XOR U30968 ( .A(p_input[2070]), .B(p_input[278]), .Z(n31146) );
  XNOR U30969 ( .A(p_input[2071]), .B(p_input[279]), .Z(n31230) );
  XNOR U30970 ( .A(n28684), .B(p_input[274]), .Z(n31141) );
  XNOR U30971 ( .A(n31155), .B(n31154), .Z(n31145) );
  XOR U30972 ( .A(n31231), .B(n31151), .Z(n31154) );
  XOR U30973 ( .A(p_input[2067]), .B(p_input[275]), .Z(n31151) );
  XNOR U30974 ( .A(p_input[2068]), .B(p_input[276]), .Z(n31231) );
  XOR U30975 ( .A(p_input[2069]), .B(p_input[277]), .Z(n31155) );
  XNOR U30976 ( .A(n31170), .B(n31156), .Z(n31228) );
  XNOR U30977 ( .A(n28686), .B(p_input[257]), .Z(n31156) );
  XNOR U30978 ( .A(n31232), .B(n31177), .Z(n31170) );
  XNOR U30979 ( .A(n31166), .B(n31165), .Z(n31177) );
  XOR U30980 ( .A(n31233), .B(n31162), .Z(n31165) );
  XNOR U30981 ( .A(n28322), .B(p_input[282]), .Z(n31162) );
  XNOR U30982 ( .A(p_input[2075]), .B(p_input[283]), .Z(n31233) );
  XOR U30983 ( .A(p_input[2076]), .B(p_input[284]), .Z(n31166) );
  XNOR U30984 ( .A(n31176), .B(n31167), .Z(n31232) );
  XNOR U30985 ( .A(n28689), .B(p_input[273]), .Z(n31167) );
  XOR U30986 ( .A(n31234), .B(n31182), .Z(n31176) );
  XNOR U30987 ( .A(p_input[2079]), .B(p_input[287]), .Z(n31182) );
  XOR U30988 ( .A(n31173), .B(n31181), .Z(n31234) );
  XOR U30989 ( .A(n31235), .B(n31178), .Z(n31181) );
  XOR U30990 ( .A(p_input[2077]), .B(p_input[285]), .Z(n31178) );
  XNOR U30991 ( .A(p_input[2078]), .B(p_input[286]), .Z(n31235) );
  XNOR U30992 ( .A(n28326), .B(p_input[281]), .Z(n31173) );
  XNOR U30993 ( .A(n31194), .B(n31193), .Z(n31160) );
  XNOR U30994 ( .A(n31236), .B(n31200), .Z(n31193) );
  XNOR U30995 ( .A(n31189), .B(n31188), .Z(n31200) );
  XOR U30996 ( .A(n31237), .B(n31185), .Z(n31188) );
  XNOR U30997 ( .A(n28694), .B(p_input[267]), .Z(n31185) );
  XNOR U30998 ( .A(p_input[2060]), .B(p_input[268]), .Z(n31237) );
  XOR U30999 ( .A(p_input[2061]), .B(p_input[269]), .Z(n31189) );
  XNOR U31000 ( .A(n31199), .B(n31190), .Z(n31236) );
  XNOR U31001 ( .A(n28330), .B(p_input[258]), .Z(n31190) );
  XOR U31002 ( .A(n31238), .B(n31205), .Z(n31199) );
  XNOR U31003 ( .A(p_input[2064]), .B(p_input[272]), .Z(n31205) );
  XOR U31004 ( .A(n31196), .B(n31204), .Z(n31238) );
  XOR U31005 ( .A(n31239), .B(n31201), .Z(n31204) );
  XOR U31006 ( .A(p_input[2062]), .B(p_input[270]), .Z(n31201) );
  XNOR U31007 ( .A(p_input[2063]), .B(p_input[271]), .Z(n31239) );
  XNOR U31008 ( .A(n28697), .B(p_input[266]), .Z(n31196) );
  XNOR U31009 ( .A(n31211), .B(n31210), .Z(n31194) );
  XNOR U31010 ( .A(n31240), .B(n31216), .Z(n31210) );
  XOR U31011 ( .A(p_input[2057]), .B(p_input[265]), .Z(n31216) );
  XOR U31012 ( .A(n31207), .B(n31215), .Z(n31240) );
  XOR U31013 ( .A(n31241), .B(n31212), .Z(n31215) );
  XOR U31014 ( .A(p_input[2055]), .B(p_input[263]), .Z(n31212) );
  XNOR U31015 ( .A(p_input[2056]), .B(p_input[264]), .Z(n31241) );
  XNOR U31016 ( .A(n28337), .B(p_input[259]), .Z(n31207) );
  XNOR U31017 ( .A(n31221), .B(n31220), .Z(n31211) );
  XOR U31018 ( .A(n31242), .B(n31217), .Z(n31220) );
  XOR U31019 ( .A(p_input[2052]), .B(p_input[260]), .Z(n31217) );
  XNOR U31020 ( .A(p_input[2053]), .B(p_input[261]), .Z(n31242) );
  XOR U31021 ( .A(p_input[2054]), .B(p_input[262]), .Z(n31221) );
  XNOR U31022 ( .A(n31243), .B(n31244), .Z(n31026) );
  AND U31023 ( .A(n287), .B(n31245), .Z(n31244) );
  XNOR U31024 ( .A(n31246), .B(n31247), .Z(n287) );
  AND U31025 ( .A(n31248), .B(n31249), .Z(n31247) );
  XOR U31026 ( .A(n31040), .B(n31246), .Z(n31249) );
  XNOR U31027 ( .A(n31250), .B(n31246), .Z(n31248) );
  XOR U31028 ( .A(n31251), .B(n31252), .Z(n31246) );
  AND U31029 ( .A(n31253), .B(n31254), .Z(n31252) );
  XOR U31030 ( .A(n31055), .B(n31251), .Z(n31254) );
  XOR U31031 ( .A(n31251), .B(n31056), .Z(n31253) );
  XOR U31032 ( .A(n31255), .B(n31256), .Z(n31251) );
  AND U31033 ( .A(n31257), .B(n31258), .Z(n31256) );
  XOR U31034 ( .A(n31083), .B(n31255), .Z(n31258) );
  XOR U31035 ( .A(n31255), .B(n31084), .Z(n31257) );
  XOR U31036 ( .A(n31259), .B(n31260), .Z(n31255) );
  AND U31037 ( .A(n31261), .B(n31262), .Z(n31260) );
  XOR U31038 ( .A(n31132), .B(n31259), .Z(n31262) );
  XOR U31039 ( .A(n31259), .B(n31133), .Z(n31261) );
  XOR U31040 ( .A(n31263), .B(n31264), .Z(n31259) );
  AND U31041 ( .A(n31265), .B(n31266), .Z(n31264) );
  XOR U31042 ( .A(n31263), .B(n31225), .Z(n31266) );
  XNOR U31043 ( .A(n31267), .B(n31268), .Z(n30976) );
  AND U31044 ( .A(n291), .B(n31269), .Z(n31268) );
  XNOR U31045 ( .A(n31270), .B(n31271), .Z(n291) );
  AND U31046 ( .A(n31272), .B(n31273), .Z(n31271) );
  XOR U31047 ( .A(n31270), .B(n30986), .Z(n31273) );
  XNOR U31048 ( .A(n31270), .B(n30936), .Z(n31272) );
  XOR U31049 ( .A(n31274), .B(n31275), .Z(n31270) );
  AND U31050 ( .A(n31276), .B(n31277), .Z(n31275) );
  XNOR U31051 ( .A(n30996), .B(n31274), .Z(n31277) );
  XOR U31052 ( .A(n31274), .B(n30946), .Z(n31276) );
  XOR U31053 ( .A(n31278), .B(n31279), .Z(n31274) );
  AND U31054 ( .A(n31280), .B(n31281), .Z(n31279) );
  XNOR U31055 ( .A(n31006), .B(n31278), .Z(n31281) );
  XOR U31056 ( .A(n31278), .B(n30955), .Z(n31280) );
  XOR U31057 ( .A(n31282), .B(n31283), .Z(n31278) );
  AND U31058 ( .A(n31284), .B(n31285), .Z(n31283) );
  XOR U31059 ( .A(n31282), .B(n30963), .Z(n31284) );
  XOR U31060 ( .A(n31286), .B(n31287), .Z(n30927) );
  AND U31061 ( .A(n295), .B(n31269), .Z(n31287) );
  XNOR U31062 ( .A(n31267), .B(n31286), .Z(n31269) );
  XNOR U31063 ( .A(n31288), .B(n31289), .Z(n295) );
  AND U31064 ( .A(n31290), .B(n31291), .Z(n31289) );
  XNOR U31065 ( .A(n31292), .B(n31288), .Z(n31291) );
  IV U31066 ( .A(n30986), .Z(n31292) );
  XOR U31067 ( .A(n31250), .B(n31293), .Z(n30986) );
  AND U31068 ( .A(n298), .B(n31294), .Z(n31293) );
  XOR U31069 ( .A(n31039), .B(n31036), .Z(n31294) );
  IV U31070 ( .A(n31250), .Z(n31039) );
  XNOR U31071 ( .A(n30936), .B(n31288), .Z(n31290) );
  XOR U31072 ( .A(n31295), .B(n31296), .Z(n30936) );
  AND U31073 ( .A(n314), .B(n31297), .Z(n31296) );
  XOR U31074 ( .A(n31298), .B(n31299), .Z(n31288) );
  AND U31075 ( .A(n31300), .B(n31301), .Z(n31299) );
  XNOR U31076 ( .A(n31298), .B(n30996), .Z(n31301) );
  XOR U31077 ( .A(n31056), .B(n31302), .Z(n30996) );
  AND U31078 ( .A(n298), .B(n31303), .Z(n31302) );
  XOR U31079 ( .A(n31052), .B(n31056), .Z(n31303) );
  XNOR U31080 ( .A(n31304), .B(n31298), .Z(n31300) );
  IV U31081 ( .A(n30946), .Z(n31304) );
  XOR U31082 ( .A(n31305), .B(n31306), .Z(n30946) );
  AND U31083 ( .A(n314), .B(n31307), .Z(n31306) );
  XOR U31084 ( .A(n31308), .B(n31309), .Z(n31298) );
  AND U31085 ( .A(n31310), .B(n31311), .Z(n31309) );
  XNOR U31086 ( .A(n31308), .B(n31006), .Z(n31311) );
  XOR U31087 ( .A(n31084), .B(n31312), .Z(n31006) );
  AND U31088 ( .A(n298), .B(n31313), .Z(n31312) );
  XOR U31089 ( .A(n31080), .B(n31084), .Z(n31313) );
  XOR U31090 ( .A(n30955), .B(n31308), .Z(n31310) );
  XOR U31091 ( .A(n31314), .B(n31315), .Z(n30955) );
  AND U31092 ( .A(n314), .B(n31316), .Z(n31315) );
  XOR U31093 ( .A(n31282), .B(n31317), .Z(n31308) );
  AND U31094 ( .A(n31318), .B(n31285), .Z(n31317) );
  XNOR U31095 ( .A(n31016), .B(n31282), .Z(n31285) );
  XOR U31096 ( .A(n31133), .B(n31319), .Z(n31016) );
  AND U31097 ( .A(n298), .B(n31320), .Z(n31319) );
  XOR U31098 ( .A(n31129), .B(n31133), .Z(n31320) );
  XNOR U31099 ( .A(n31321), .B(n31282), .Z(n31318) );
  IV U31100 ( .A(n30963), .Z(n31321) );
  XOR U31101 ( .A(n31322), .B(n31323), .Z(n30963) );
  AND U31102 ( .A(n314), .B(n31324), .Z(n31323) );
  XOR U31103 ( .A(n31325), .B(n31326), .Z(n31282) );
  AND U31104 ( .A(n31327), .B(n31328), .Z(n31326) );
  XNOR U31105 ( .A(n31325), .B(n31024), .Z(n31328) );
  XOR U31106 ( .A(n31226), .B(n31329), .Z(n31024) );
  AND U31107 ( .A(n298), .B(n31330), .Z(n31329) );
  XOR U31108 ( .A(n31222), .B(n31226), .Z(n31330) );
  XNOR U31109 ( .A(n31331), .B(n31325), .Z(n31327) );
  IV U31110 ( .A(n30973), .Z(n31331) );
  XOR U31111 ( .A(n31332), .B(n31333), .Z(n30973) );
  AND U31112 ( .A(n314), .B(n31334), .Z(n31333) );
  AND U31113 ( .A(n31286), .B(n31267), .Z(n31325) );
  XNOR U31114 ( .A(n31335), .B(n31336), .Z(n31267) );
  AND U31115 ( .A(n298), .B(n31245), .Z(n31336) );
  XNOR U31116 ( .A(n31243), .B(n31335), .Z(n31245) );
  XNOR U31117 ( .A(n31337), .B(n31338), .Z(n298) );
  AND U31118 ( .A(n31339), .B(n31340), .Z(n31338) );
  XNOR U31119 ( .A(n31337), .B(n31036), .Z(n31340) );
  IV U31120 ( .A(n31040), .Z(n31036) );
  XOR U31121 ( .A(n31341), .B(n31342), .Z(n31040) );
  AND U31122 ( .A(n302), .B(n31343), .Z(n31342) );
  XOR U31123 ( .A(n31344), .B(n31341), .Z(n31343) );
  XNOR U31124 ( .A(n31337), .B(n31250), .Z(n31339) );
  XOR U31125 ( .A(n31345), .B(n31346), .Z(n31250) );
  AND U31126 ( .A(n310), .B(n31297), .Z(n31346) );
  XOR U31127 ( .A(n31295), .B(n31345), .Z(n31297) );
  XOR U31128 ( .A(n31347), .B(n31348), .Z(n31337) );
  AND U31129 ( .A(n31349), .B(n31350), .Z(n31348) );
  XNOR U31130 ( .A(n31347), .B(n31052), .Z(n31350) );
  IV U31131 ( .A(n31055), .Z(n31052) );
  XOR U31132 ( .A(n31351), .B(n31352), .Z(n31055) );
  AND U31133 ( .A(n302), .B(n31353), .Z(n31352) );
  XOR U31134 ( .A(n31354), .B(n31351), .Z(n31353) );
  XOR U31135 ( .A(n31056), .B(n31347), .Z(n31349) );
  XOR U31136 ( .A(n31355), .B(n31356), .Z(n31056) );
  AND U31137 ( .A(n310), .B(n31307), .Z(n31356) );
  XOR U31138 ( .A(n31355), .B(n31305), .Z(n31307) );
  XOR U31139 ( .A(n31357), .B(n31358), .Z(n31347) );
  AND U31140 ( .A(n31359), .B(n31360), .Z(n31358) );
  XNOR U31141 ( .A(n31357), .B(n31080), .Z(n31360) );
  IV U31142 ( .A(n31083), .Z(n31080) );
  XOR U31143 ( .A(n31361), .B(n31362), .Z(n31083) );
  AND U31144 ( .A(n302), .B(n31363), .Z(n31362) );
  XNOR U31145 ( .A(n31364), .B(n31361), .Z(n31363) );
  XOR U31146 ( .A(n31084), .B(n31357), .Z(n31359) );
  XOR U31147 ( .A(n31365), .B(n31366), .Z(n31084) );
  AND U31148 ( .A(n310), .B(n31316), .Z(n31366) );
  XOR U31149 ( .A(n31365), .B(n31314), .Z(n31316) );
  XOR U31150 ( .A(n31367), .B(n31368), .Z(n31357) );
  AND U31151 ( .A(n31369), .B(n31370), .Z(n31368) );
  XNOR U31152 ( .A(n31367), .B(n31129), .Z(n31370) );
  IV U31153 ( .A(n31132), .Z(n31129) );
  XOR U31154 ( .A(n31371), .B(n31372), .Z(n31132) );
  AND U31155 ( .A(n302), .B(n31373), .Z(n31372) );
  XOR U31156 ( .A(n31374), .B(n31371), .Z(n31373) );
  XOR U31157 ( .A(n31133), .B(n31367), .Z(n31369) );
  XOR U31158 ( .A(n31375), .B(n31376), .Z(n31133) );
  AND U31159 ( .A(n310), .B(n31324), .Z(n31376) );
  XOR U31160 ( .A(n31375), .B(n31322), .Z(n31324) );
  XOR U31161 ( .A(n31263), .B(n31377), .Z(n31367) );
  AND U31162 ( .A(n31265), .B(n31378), .Z(n31377) );
  XNOR U31163 ( .A(n31263), .B(n31222), .Z(n31378) );
  IV U31164 ( .A(n31225), .Z(n31222) );
  XOR U31165 ( .A(n31379), .B(n31380), .Z(n31225) );
  AND U31166 ( .A(n302), .B(n31381), .Z(n31380) );
  XNOR U31167 ( .A(n31382), .B(n31379), .Z(n31381) );
  XOR U31168 ( .A(n31226), .B(n31263), .Z(n31265) );
  XOR U31169 ( .A(n31383), .B(n31384), .Z(n31226) );
  AND U31170 ( .A(n310), .B(n31334), .Z(n31384) );
  XOR U31171 ( .A(n31383), .B(n31332), .Z(n31334) );
  AND U31172 ( .A(n31335), .B(n31243), .Z(n31263) );
  XNOR U31173 ( .A(n31385), .B(n31386), .Z(n31243) );
  AND U31174 ( .A(n302), .B(n31387), .Z(n31386) );
  XNOR U31175 ( .A(n31388), .B(n31385), .Z(n31387) );
  XNOR U31176 ( .A(n31389), .B(n31390), .Z(n302) );
  AND U31177 ( .A(n31391), .B(n31392), .Z(n31390) );
  XOR U31178 ( .A(n31344), .B(n31389), .Z(n31392) );
  AND U31179 ( .A(n31393), .B(n31394), .Z(n31344) );
  XNOR U31180 ( .A(n31341), .B(n31389), .Z(n31391) );
  XNOR U31181 ( .A(n31395), .B(n31396), .Z(n31341) );
  AND U31182 ( .A(n306), .B(n31397), .Z(n31396) );
  XNOR U31183 ( .A(n31398), .B(n31399), .Z(n31397) );
  XOR U31184 ( .A(n31400), .B(n31401), .Z(n31389) );
  AND U31185 ( .A(n31402), .B(n31403), .Z(n31401) );
  XNOR U31186 ( .A(n31400), .B(n31393), .Z(n31403) );
  IV U31187 ( .A(n31354), .Z(n31393) );
  XOR U31188 ( .A(n31404), .B(n31405), .Z(n31354) );
  XOR U31189 ( .A(n31406), .B(n31394), .Z(n31405) );
  AND U31190 ( .A(n31364), .B(n31407), .Z(n31394) );
  AND U31191 ( .A(n31408), .B(n31409), .Z(n31406) );
  XOR U31192 ( .A(n31410), .B(n31404), .Z(n31408) );
  XNOR U31193 ( .A(n31351), .B(n31400), .Z(n31402) );
  XNOR U31194 ( .A(n31411), .B(n31412), .Z(n31351) );
  AND U31195 ( .A(n306), .B(n31413), .Z(n31412) );
  XNOR U31196 ( .A(n31414), .B(n31415), .Z(n31413) );
  XOR U31197 ( .A(n31416), .B(n31417), .Z(n31400) );
  AND U31198 ( .A(n31418), .B(n31419), .Z(n31417) );
  XNOR U31199 ( .A(n31416), .B(n31364), .Z(n31419) );
  XOR U31200 ( .A(n31420), .B(n31409), .Z(n31364) );
  XNOR U31201 ( .A(n31421), .B(n31404), .Z(n31409) );
  XOR U31202 ( .A(n31422), .B(n31423), .Z(n31404) );
  AND U31203 ( .A(n31424), .B(n31425), .Z(n31423) );
  XOR U31204 ( .A(n31426), .B(n31422), .Z(n31424) );
  XNOR U31205 ( .A(n31427), .B(n31428), .Z(n31421) );
  AND U31206 ( .A(n31429), .B(n31430), .Z(n31428) );
  XOR U31207 ( .A(n31427), .B(n31431), .Z(n31429) );
  XNOR U31208 ( .A(n31410), .B(n31407), .Z(n31420) );
  AND U31209 ( .A(n31432), .B(n31433), .Z(n31407) );
  XOR U31210 ( .A(n31434), .B(n31435), .Z(n31410) );
  AND U31211 ( .A(n31436), .B(n31437), .Z(n31435) );
  XOR U31212 ( .A(n31434), .B(n31438), .Z(n31436) );
  XNOR U31213 ( .A(n31361), .B(n31416), .Z(n31418) );
  XNOR U31214 ( .A(n31439), .B(n31440), .Z(n31361) );
  AND U31215 ( .A(n306), .B(n31441), .Z(n31440) );
  XNOR U31216 ( .A(n31442), .B(n31443), .Z(n31441) );
  XOR U31217 ( .A(n31444), .B(n31445), .Z(n31416) );
  AND U31218 ( .A(n31446), .B(n31447), .Z(n31445) );
  XNOR U31219 ( .A(n31444), .B(n31432), .Z(n31447) );
  IV U31220 ( .A(n31374), .Z(n31432) );
  XNOR U31221 ( .A(n31448), .B(n31425), .Z(n31374) );
  XNOR U31222 ( .A(n31449), .B(n31431), .Z(n31425) );
  XOR U31223 ( .A(n31450), .B(n31451), .Z(n31431) );
  AND U31224 ( .A(n31452), .B(n31453), .Z(n31451) );
  XOR U31225 ( .A(n31450), .B(n31454), .Z(n31452) );
  XNOR U31226 ( .A(n31430), .B(n31422), .Z(n31449) );
  XOR U31227 ( .A(n31455), .B(n31456), .Z(n31422) );
  AND U31228 ( .A(n31457), .B(n31458), .Z(n31456) );
  XNOR U31229 ( .A(n31459), .B(n31455), .Z(n31457) );
  XNOR U31230 ( .A(n31460), .B(n31427), .Z(n31430) );
  XOR U31231 ( .A(n31461), .B(n31462), .Z(n31427) );
  AND U31232 ( .A(n31463), .B(n31464), .Z(n31462) );
  XOR U31233 ( .A(n31461), .B(n31465), .Z(n31463) );
  XNOR U31234 ( .A(n31466), .B(n31467), .Z(n31460) );
  AND U31235 ( .A(n31468), .B(n31469), .Z(n31467) );
  XNOR U31236 ( .A(n31466), .B(n31470), .Z(n31468) );
  XNOR U31237 ( .A(n31426), .B(n31433), .Z(n31448) );
  AND U31238 ( .A(n31382), .B(n31471), .Z(n31433) );
  XOR U31239 ( .A(n31438), .B(n31437), .Z(n31426) );
  XNOR U31240 ( .A(n31472), .B(n31434), .Z(n31437) );
  XOR U31241 ( .A(n31473), .B(n31474), .Z(n31434) );
  AND U31242 ( .A(n31475), .B(n31476), .Z(n31474) );
  XOR U31243 ( .A(n31473), .B(n31477), .Z(n31475) );
  XNOR U31244 ( .A(n31478), .B(n31479), .Z(n31472) );
  AND U31245 ( .A(n31480), .B(n31481), .Z(n31479) );
  XOR U31246 ( .A(n31478), .B(n31482), .Z(n31480) );
  XOR U31247 ( .A(n31483), .B(n31484), .Z(n31438) );
  AND U31248 ( .A(n31485), .B(n31486), .Z(n31484) );
  XOR U31249 ( .A(n31483), .B(n31487), .Z(n31485) );
  XNOR U31250 ( .A(n31371), .B(n31444), .Z(n31446) );
  XNOR U31251 ( .A(n31488), .B(n31489), .Z(n31371) );
  AND U31252 ( .A(n306), .B(n31490), .Z(n31489) );
  XNOR U31253 ( .A(n31491), .B(n31492), .Z(n31490) );
  XOR U31254 ( .A(n31493), .B(n31494), .Z(n31444) );
  AND U31255 ( .A(n31495), .B(n31496), .Z(n31494) );
  XNOR U31256 ( .A(n31493), .B(n31382), .Z(n31496) );
  XOR U31257 ( .A(n31497), .B(n31458), .Z(n31382) );
  XNOR U31258 ( .A(n31498), .B(n31465), .Z(n31458) );
  XOR U31259 ( .A(n31454), .B(n31453), .Z(n31465) );
  XNOR U31260 ( .A(n31499), .B(n31450), .Z(n31453) );
  XOR U31261 ( .A(n31500), .B(n31501), .Z(n31450) );
  AND U31262 ( .A(n31502), .B(n31503), .Z(n31501) );
  XOR U31263 ( .A(n31500), .B(n31504), .Z(n31502) );
  XNOR U31264 ( .A(n31505), .B(n31506), .Z(n31499) );
  NOR U31265 ( .A(n31507), .B(n31508), .Z(n31506) );
  XNOR U31266 ( .A(n31505), .B(n31509), .Z(n31507) );
  XOR U31267 ( .A(n31510), .B(n31511), .Z(n31454) );
  NOR U31268 ( .A(n31512), .B(n31513), .Z(n31511) );
  XNOR U31269 ( .A(n31510), .B(n31514), .Z(n31512) );
  XNOR U31270 ( .A(n31464), .B(n31455), .Z(n31498) );
  XOR U31271 ( .A(n31515), .B(n31516), .Z(n31455) );
  NOR U31272 ( .A(n31517), .B(n31518), .Z(n31516) );
  XNOR U31273 ( .A(n31515), .B(n31519), .Z(n31517) );
  XOR U31274 ( .A(n31520), .B(n31470), .Z(n31464) );
  XNOR U31275 ( .A(n31521), .B(n31522), .Z(n31470) );
  NOR U31276 ( .A(n31523), .B(n31524), .Z(n31522) );
  XNOR U31277 ( .A(n31521), .B(n31525), .Z(n31523) );
  XNOR U31278 ( .A(n31469), .B(n31461), .Z(n31520) );
  XOR U31279 ( .A(n31526), .B(n31527), .Z(n31461) );
  AND U31280 ( .A(n31528), .B(n31529), .Z(n31527) );
  XOR U31281 ( .A(n31526), .B(n31530), .Z(n31528) );
  XNOR U31282 ( .A(n31531), .B(n31466), .Z(n31469) );
  XOR U31283 ( .A(n31532), .B(n31533), .Z(n31466) );
  AND U31284 ( .A(n31534), .B(n31535), .Z(n31533) );
  XOR U31285 ( .A(n31532), .B(n31536), .Z(n31534) );
  XNOR U31286 ( .A(n31537), .B(n31538), .Z(n31531) );
  NOR U31287 ( .A(n31539), .B(n31540), .Z(n31538) );
  XOR U31288 ( .A(n31537), .B(n31541), .Z(n31539) );
  XOR U31289 ( .A(n31459), .B(n31471), .Z(n31497) );
  NOR U31290 ( .A(n31388), .B(n31542), .Z(n31471) );
  XNOR U31291 ( .A(n31477), .B(n31476), .Z(n31459) );
  XNOR U31292 ( .A(n31543), .B(n31482), .Z(n31476) );
  XOR U31293 ( .A(n31544), .B(n31545), .Z(n31482) );
  NOR U31294 ( .A(n31546), .B(n31547), .Z(n31545) );
  XNOR U31295 ( .A(n31544), .B(n31548), .Z(n31546) );
  XNOR U31296 ( .A(n31481), .B(n31473), .Z(n31543) );
  XOR U31297 ( .A(n31549), .B(n31550), .Z(n31473) );
  AND U31298 ( .A(n31551), .B(n31552), .Z(n31550) );
  XNOR U31299 ( .A(n31549), .B(n31553), .Z(n31551) );
  XNOR U31300 ( .A(n31554), .B(n31478), .Z(n31481) );
  XOR U31301 ( .A(n31555), .B(n31556), .Z(n31478) );
  AND U31302 ( .A(n31557), .B(n31558), .Z(n31556) );
  XOR U31303 ( .A(n31555), .B(n31559), .Z(n31557) );
  XNOR U31304 ( .A(n31560), .B(n31561), .Z(n31554) );
  NOR U31305 ( .A(n31562), .B(n31563), .Z(n31561) );
  XOR U31306 ( .A(n31560), .B(n31564), .Z(n31562) );
  XOR U31307 ( .A(n31487), .B(n31486), .Z(n31477) );
  XNOR U31308 ( .A(n31565), .B(n31483), .Z(n31486) );
  XOR U31309 ( .A(n31566), .B(n31567), .Z(n31483) );
  AND U31310 ( .A(n31568), .B(n31569), .Z(n31567) );
  XOR U31311 ( .A(n31566), .B(n31570), .Z(n31568) );
  XNOR U31312 ( .A(n31571), .B(n31572), .Z(n31565) );
  NOR U31313 ( .A(n31573), .B(n31574), .Z(n31572) );
  XNOR U31314 ( .A(n31571), .B(n31575), .Z(n31573) );
  XOR U31315 ( .A(n31576), .B(n31577), .Z(n31487) );
  NOR U31316 ( .A(n31578), .B(n31579), .Z(n31577) );
  XNOR U31317 ( .A(n31576), .B(n31580), .Z(n31578) );
  XNOR U31318 ( .A(n31379), .B(n31493), .Z(n31495) );
  XNOR U31319 ( .A(n31581), .B(n31582), .Z(n31379) );
  AND U31320 ( .A(n306), .B(n31583), .Z(n31582) );
  XNOR U31321 ( .A(n31584), .B(n31585), .Z(n31583) );
  AND U31322 ( .A(n31385), .B(n31388), .Z(n31493) );
  XOR U31323 ( .A(n31586), .B(n31542), .Z(n31388) );
  XNOR U31324 ( .A(p_input[2048]), .B(p_input[288]), .Z(n31542) );
  XOR U31325 ( .A(n31519), .B(n31518), .Z(n31586) );
  XOR U31326 ( .A(n31587), .B(n31530), .Z(n31518) );
  XOR U31327 ( .A(n31504), .B(n31503), .Z(n31530) );
  XNOR U31328 ( .A(n31588), .B(n31509), .Z(n31503) );
  XOR U31329 ( .A(p_input[2072]), .B(p_input[312]), .Z(n31509) );
  XOR U31330 ( .A(n31500), .B(n31508), .Z(n31588) );
  XOR U31331 ( .A(n31589), .B(n31505), .Z(n31508) );
  XOR U31332 ( .A(p_input[2070]), .B(p_input[310]), .Z(n31505) );
  XNOR U31333 ( .A(p_input[2071]), .B(p_input[311]), .Z(n31589) );
  XNOR U31334 ( .A(n28684), .B(p_input[306]), .Z(n31500) );
  XNOR U31335 ( .A(n31514), .B(n31513), .Z(n31504) );
  XOR U31336 ( .A(n31590), .B(n31510), .Z(n31513) );
  XOR U31337 ( .A(p_input[2067]), .B(p_input[307]), .Z(n31510) );
  XNOR U31338 ( .A(p_input[2068]), .B(p_input[308]), .Z(n31590) );
  XOR U31339 ( .A(p_input[2069]), .B(p_input[309]), .Z(n31514) );
  XNOR U31340 ( .A(n31529), .B(n31515), .Z(n31587) );
  XNOR U31341 ( .A(n28686), .B(p_input[289]), .Z(n31515) );
  XNOR U31342 ( .A(n31591), .B(n31536), .Z(n31529) );
  XNOR U31343 ( .A(n31525), .B(n31524), .Z(n31536) );
  XOR U31344 ( .A(n31592), .B(n31521), .Z(n31524) );
  XNOR U31345 ( .A(n28322), .B(p_input[314]), .Z(n31521) );
  XNOR U31346 ( .A(p_input[2075]), .B(p_input[315]), .Z(n31592) );
  XOR U31347 ( .A(p_input[2076]), .B(p_input[316]), .Z(n31525) );
  XNOR U31348 ( .A(n31535), .B(n31526), .Z(n31591) );
  XNOR U31349 ( .A(n28689), .B(p_input[305]), .Z(n31526) );
  XOR U31350 ( .A(n31593), .B(n31541), .Z(n31535) );
  XNOR U31351 ( .A(p_input[2079]), .B(p_input[319]), .Z(n31541) );
  XOR U31352 ( .A(n31532), .B(n31540), .Z(n31593) );
  XOR U31353 ( .A(n31594), .B(n31537), .Z(n31540) );
  XOR U31354 ( .A(p_input[2077]), .B(p_input[317]), .Z(n31537) );
  XNOR U31355 ( .A(p_input[2078]), .B(p_input[318]), .Z(n31594) );
  XNOR U31356 ( .A(n28326), .B(p_input[313]), .Z(n31532) );
  XNOR U31357 ( .A(n31553), .B(n31552), .Z(n31519) );
  XNOR U31358 ( .A(n31595), .B(n31559), .Z(n31552) );
  XNOR U31359 ( .A(n31548), .B(n31547), .Z(n31559) );
  XOR U31360 ( .A(n31596), .B(n31544), .Z(n31547) );
  XNOR U31361 ( .A(n28694), .B(p_input[299]), .Z(n31544) );
  XNOR U31362 ( .A(p_input[2060]), .B(p_input[300]), .Z(n31596) );
  XOR U31363 ( .A(p_input[2061]), .B(p_input[301]), .Z(n31548) );
  XNOR U31364 ( .A(n31558), .B(n31549), .Z(n31595) );
  XNOR U31365 ( .A(n28330), .B(p_input[290]), .Z(n31549) );
  XOR U31366 ( .A(n31597), .B(n31564), .Z(n31558) );
  XNOR U31367 ( .A(p_input[2064]), .B(p_input[304]), .Z(n31564) );
  XOR U31368 ( .A(n31555), .B(n31563), .Z(n31597) );
  XOR U31369 ( .A(n31598), .B(n31560), .Z(n31563) );
  XOR U31370 ( .A(p_input[2062]), .B(p_input[302]), .Z(n31560) );
  XNOR U31371 ( .A(p_input[2063]), .B(p_input[303]), .Z(n31598) );
  XNOR U31372 ( .A(n28697), .B(p_input[298]), .Z(n31555) );
  XNOR U31373 ( .A(n31570), .B(n31569), .Z(n31553) );
  XNOR U31374 ( .A(n31599), .B(n31575), .Z(n31569) );
  XOR U31375 ( .A(p_input[2057]), .B(p_input[297]), .Z(n31575) );
  XOR U31376 ( .A(n31566), .B(n31574), .Z(n31599) );
  XOR U31377 ( .A(n31600), .B(n31571), .Z(n31574) );
  XOR U31378 ( .A(p_input[2055]), .B(p_input[295]), .Z(n31571) );
  XNOR U31379 ( .A(p_input[2056]), .B(p_input[296]), .Z(n31600) );
  XNOR U31380 ( .A(n28337), .B(p_input[291]), .Z(n31566) );
  XNOR U31381 ( .A(n31580), .B(n31579), .Z(n31570) );
  XOR U31382 ( .A(n31601), .B(n31576), .Z(n31579) );
  XOR U31383 ( .A(p_input[2052]), .B(p_input[292]), .Z(n31576) );
  XNOR U31384 ( .A(p_input[2053]), .B(p_input[293]), .Z(n31601) );
  XOR U31385 ( .A(p_input[2054]), .B(p_input[294]), .Z(n31580) );
  XNOR U31386 ( .A(n31602), .B(n31603), .Z(n31385) );
  AND U31387 ( .A(n306), .B(n31604), .Z(n31603) );
  XNOR U31388 ( .A(n31605), .B(n31606), .Z(n306) );
  AND U31389 ( .A(n31607), .B(n31608), .Z(n31606) );
  XOR U31390 ( .A(n31399), .B(n31605), .Z(n31608) );
  XNOR U31391 ( .A(n31609), .B(n31605), .Z(n31607) );
  XOR U31392 ( .A(n31610), .B(n31611), .Z(n31605) );
  AND U31393 ( .A(n31612), .B(n31613), .Z(n31611) );
  XOR U31394 ( .A(n31414), .B(n31610), .Z(n31613) );
  XOR U31395 ( .A(n31610), .B(n31415), .Z(n31612) );
  XOR U31396 ( .A(n31614), .B(n31615), .Z(n31610) );
  AND U31397 ( .A(n31616), .B(n31617), .Z(n31615) );
  XOR U31398 ( .A(n31442), .B(n31614), .Z(n31617) );
  XOR U31399 ( .A(n31614), .B(n31443), .Z(n31616) );
  XOR U31400 ( .A(n31618), .B(n31619), .Z(n31614) );
  AND U31401 ( .A(n31620), .B(n31621), .Z(n31619) );
  XOR U31402 ( .A(n31491), .B(n31618), .Z(n31621) );
  XOR U31403 ( .A(n31618), .B(n31492), .Z(n31620) );
  XOR U31404 ( .A(n31622), .B(n31623), .Z(n31618) );
  AND U31405 ( .A(n31624), .B(n31625), .Z(n31623) );
  XOR U31406 ( .A(n31622), .B(n31584), .Z(n31625) );
  XNOR U31407 ( .A(n31626), .B(n31627), .Z(n31335) );
  AND U31408 ( .A(n310), .B(n31628), .Z(n31627) );
  XNOR U31409 ( .A(n31629), .B(n31630), .Z(n310) );
  AND U31410 ( .A(n31631), .B(n31632), .Z(n31630) );
  XOR U31411 ( .A(n31629), .B(n31345), .Z(n31632) );
  XNOR U31412 ( .A(n31629), .B(n31295), .Z(n31631) );
  XOR U31413 ( .A(n31633), .B(n31634), .Z(n31629) );
  AND U31414 ( .A(n31635), .B(n31636), .Z(n31634) );
  XNOR U31415 ( .A(n31355), .B(n31633), .Z(n31636) );
  XOR U31416 ( .A(n31633), .B(n31305), .Z(n31635) );
  XOR U31417 ( .A(n31637), .B(n31638), .Z(n31633) );
  AND U31418 ( .A(n31639), .B(n31640), .Z(n31638) );
  XNOR U31419 ( .A(n31365), .B(n31637), .Z(n31640) );
  XOR U31420 ( .A(n31637), .B(n31314), .Z(n31639) );
  XOR U31421 ( .A(n31641), .B(n31642), .Z(n31637) );
  AND U31422 ( .A(n31643), .B(n31644), .Z(n31642) );
  XOR U31423 ( .A(n31641), .B(n31322), .Z(n31643) );
  XOR U31424 ( .A(n31645), .B(n31646), .Z(n31286) );
  AND U31425 ( .A(n314), .B(n31628), .Z(n31646) );
  XNOR U31426 ( .A(n31626), .B(n31645), .Z(n31628) );
  XNOR U31427 ( .A(n31647), .B(n31648), .Z(n314) );
  AND U31428 ( .A(n31649), .B(n31650), .Z(n31648) );
  XNOR U31429 ( .A(n31651), .B(n31647), .Z(n31650) );
  IV U31430 ( .A(n31345), .Z(n31651) );
  XOR U31431 ( .A(n31609), .B(n31652), .Z(n31345) );
  AND U31432 ( .A(n317), .B(n31653), .Z(n31652) );
  XOR U31433 ( .A(n31398), .B(n31395), .Z(n31653) );
  IV U31434 ( .A(n31609), .Z(n31398) );
  XNOR U31435 ( .A(n31295), .B(n31647), .Z(n31649) );
  XOR U31436 ( .A(n31654), .B(n31655), .Z(n31295) );
  AND U31437 ( .A(n333), .B(n31656), .Z(n31655) );
  XOR U31438 ( .A(n31657), .B(n31658), .Z(n31647) );
  AND U31439 ( .A(n31659), .B(n31660), .Z(n31658) );
  XNOR U31440 ( .A(n31657), .B(n31355), .Z(n31660) );
  XOR U31441 ( .A(n31415), .B(n31661), .Z(n31355) );
  AND U31442 ( .A(n317), .B(n31662), .Z(n31661) );
  XOR U31443 ( .A(n31411), .B(n31415), .Z(n31662) );
  XNOR U31444 ( .A(n31663), .B(n31657), .Z(n31659) );
  IV U31445 ( .A(n31305), .Z(n31663) );
  XOR U31446 ( .A(n31664), .B(n31665), .Z(n31305) );
  AND U31447 ( .A(n333), .B(n31666), .Z(n31665) );
  XOR U31448 ( .A(n31667), .B(n31668), .Z(n31657) );
  AND U31449 ( .A(n31669), .B(n31670), .Z(n31668) );
  XNOR U31450 ( .A(n31667), .B(n31365), .Z(n31670) );
  XOR U31451 ( .A(n31443), .B(n31671), .Z(n31365) );
  AND U31452 ( .A(n317), .B(n31672), .Z(n31671) );
  XOR U31453 ( .A(n31439), .B(n31443), .Z(n31672) );
  XOR U31454 ( .A(n31314), .B(n31667), .Z(n31669) );
  XOR U31455 ( .A(n31673), .B(n31674), .Z(n31314) );
  AND U31456 ( .A(n333), .B(n31675), .Z(n31674) );
  XOR U31457 ( .A(n31641), .B(n31676), .Z(n31667) );
  AND U31458 ( .A(n31677), .B(n31644), .Z(n31676) );
  XNOR U31459 ( .A(n31375), .B(n31641), .Z(n31644) );
  XOR U31460 ( .A(n31492), .B(n31678), .Z(n31375) );
  AND U31461 ( .A(n317), .B(n31679), .Z(n31678) );
  XOR U31462 ( .A(n31488), .B(n31492), .Z(n31679) );
  XNOR U31463 ( .A(n31680), .B(n31641), .Z(n31677) );
  IV U31464 ( .A(n31322), .Z(n31680) );
  XOR U31465 ( .A(n31681), .B(n31682), .Z(n31322) );
  AND U31466 ( .A(n333), .B(n31683), .Z(n31682) );
  XOR U31467 ( .A(n31684), .B(n31685), .Z(n31641) );
  AND U31468 ( .A(n31686), .B(n31687), .Z(n31685) );
  XNOR U31469 ( .A(n31684), .B(n31383), .Z(n31687) );
  XOR U31470 ( .A(n31585), .B(n31688), .Z(n31383) );
  AND U31471 ( .A(n317), .B(n31689), .Z(n31688) );
  XOR U31472 ( .A(n31581), .B(n31585), .Z(n31689) );
  XNOR U31473 ( .A(n31690), .B(n31684), .Z(n31686) );
  IV U31474 ( .A(n31332), .Z(n31690) );
  XOR U31475 ( .A(n31691), .B(n31692), .Z(n31332) );
  AND U31476 ( .A(n333), .B(n31693), .Z(n31692) );
  AND U31477 ( .A(n31645), .B(n31626), .Z(n31684) );
  XNOR U31478 ( .A(n31694), .B(n31695), .Z(n31626) );
  AND U31479 ( .A(n317), .B(n31604), .Z(n31695) );
  XNOR U31480 ( .A(n31602), .B(n31694), .Z(n31604) );
  XNOR U31481 ( .A(n31696), .B(n31697), .Z(n317) );
  AND U31482 ( .A(n31698), .B(n31699), .Z(n31697) );
  XNOR U31483 ( .A(n31696), .B(n31395), .Z(n31699) );
  IV U31484 ( .A(n31399), .Z(n31395) );
  XOR U31485 ( .A(n31700), .B(n31701), .Z(n31399) );
  AND U31486 ( .A(n321), .B(n31702), .Z(n31701) );
  XOR U31487 ( .A(n31703), .B(n31700), .Z(n31702) );
  XNOR U31488 ( .A(n31696), .B(n31609), .Z(n31698) );
  XOR U31489 ( .A(n31704), .B(n31705), .Z(n31609) );
  AND U31490 ( .A(n329), .B(n31656), .Z(n31705) );
  XOR U31491 ( .A(n31654), .B(n31704), .Z(n31656) );
  XOR U31492 ( .A(n31706), .B(n31707), .Z(n31696) );
  AND U31493 ( .A(n31708), .B(n31709), .Z(n31707) );
  XNOR U31494 ( .A(n31706), .B(n31411), .Z(n31709) );
  IV U31495 ( .A(n31414), .Z(n31411) );
  XOR U31496 ( .A(n31710), .B(n31711), .Z(n31414) );
  AND U31497 ( .A(n321), .B(n31712), .Z(n31711) );
  XOR U31498 ( .A(n31713), .B(n31710), .Z(n31712) );
  XOR U31499 ( .A(n31415), .B(n31706), .Z(n31708) );
  XOR U31500 ( .A(n31714), .B(n31715), .Z(n31415) );
  AND U31501 ( .A(n329), .B(n31666), .Z(n31715) );
  XOR U31502 ( .A(n31714), .B(n31664), .Z(n31666) );
  XOR U31503 ( .A(n31716), .B(n31717), .Z(n31706) );
  AND U31504 ( .A(n31718), .B(n31719), .Z(n31717) );
  XNOR U31505 ( .A(n31716), .B(n31439), .Z(n31719) );
  IV U31506 ( .A(n31442), .Z(n31439) );
  XOR U31507 ( .A(n31720), .B(n31721), .Z(n31442) );
  AND U31508 ( .A(n321), .B(n31722), .Z(n31721) );
  XNOR U31509 ( .A(n31723), .B(n31720), .Z(n31722) );
  XOR U31510 ( .A(n31443), .B(n31716), .Z(n31718) );
  XOR U31511 ( .A(n31724), .B(n31725), .Z(n31443) );
  AND U31512 ( .A(n329), .B(n31675), .Z(n31725) );
  XOR U31513 ( .A(n31724), .B(n31673), .Z(n31675) );
  XOR U31514 ( .A(n31726), .B(n31727), .Z(n31716) );
  AND U31515 ( .A(n31728), .B(n31729), .Z(n31727) );
  XNOR U31516 ( .A(n31726), .B(n31488), .Z(n31729) );
  IV U31517 ( .A(n31491), .Z(n31488) );
  XOR U31518 ( .A(n31730), .B(n31731), .Z(n31491) );
  AND U31519 ( .A(n321), .B(n31732), .Z(n31731) );
  XOR U31520 ( .A(n31733), .B(n31730), .Z(n31732) );
  XOR U31521 ( .A(n31492), .B(n31726), .Z(n31728) );
  XOR U31522 ( .A(n31734), .B(n31735), .Z(n31492) );
  AND U31523 ( .A(n329), .B(n31683), .Z(n31735) );
  XOR U31524 ( .A(n31734), .B(n31681), .Z(n31683) );
  XOR U31525 ( .A(n31622), .B(n31736), .Z(n31726) );
  AND U31526 ( .A(n31624), .B(n31737), .Z(n31736) );
  XNOR U31527 ( .A(n31622), .B(n31581), .Z(n31737) );
  IV U31528 ( .A(n31584), .Z(n31581) );
  XOR U31529 ( .A(n31738), .B(n31739), .Z(n31584) );
  AND U31530 ( .A(n321), .B(n31740), .Z(n31739) );
  XNOR U31531 ( .A(n31741), .B(n31738), .Z(n31740) );
  XOR U31532 ( .A(n31585), .B(n31622), .Z(n31624) );
  XOR U31533 ( .A(n31742), .B(n31743), .Z(n31585) );
  AND U31534 ( .A(n329), .B(n31693), .Z(n31743) );
  XOR U31535 ( .A(n31742), .B(n31691), .Z(n31693) );
  AND U31536 ( .A(n31694), .B(n31602), .Z(n31622) );
  XNOR U31537 ( .A(n31744), .B(n31745), .Z(n31602) );
  AND U31538 ( .A(n321), .B(n31746), .Z(n31745) );
  XNOR U31539 ( .A(n31747), .B(n31744), .Z(n31746) );
  XNOR U31540 ( .A(n31748), .B(n31749), .Z(n321) );
  AND U31541 ( .A(n31750), .B(n31751), .Z(n31749) );
  XOR U31542 ( .A(n31703), .B(n31748), .Z(n31751) );
  AND U31543 ( .A(n31752), .B(n31753), .Z(n31703) );
  XNOR U31544 ( .A(n31700), .B(n31748), .Z(n31750) );
  XNOR U31545 ( .A(n31754), .B(n31755), .Z(n31700) );
  AND U31546 ( .A(n325), .B(n31756), .Z(n31755) );
  XNOR U31547 ( .A(n31757), .B(n31758), .Z(n31756) );
  XOR U31548 ( .A(n31759), .B(n31760), .Z(n31748) );
  AND U31549 ( .A(n31761), .B(n31762), .Z(n31760) );
  XNOR U31550 ( .A(n31759), .B(n31752), .Z(n31762) );
  IV U31551 ( .A(n31713), .Z(n31752) );
  XOR U31552 ( .A(n31763), .B(n31764), .Z(n31713) );
  XOR U31553 ( .A(n31765), .B(n31753), .Z(n31764) );
  AND U31554 ( .A(n31723), .B(n31766), .Z(n31753) );
  AND U31555 ( .A(n31767), .B(n31768), .Z(n31765) );
  XOR U31556 ( .A(n31769), .B(n31763), .Z(n31767) );
  XNOR U31557 ( .A(n31710), .B(n31759), .Z(n31761) );
  XNOR U31558 ( .A(n31770), .B(n31771), .Z(n31710) );
  AND U31559 ( .A(n325), .B(n31772), .Z(n31771) );
  XNOR U31560 ( .A(n31773), .B(n31774), .Z(n31772) );
  XOR U31561 ( .A(n31775), .B(n31776), .Z(n31759) );
  AND U31562 ( .A(n31777), .B(n31778), .Z(n31776) );
  XNOR U31563 ( .A(n31775), .B(n31723), .Z(n31778) );
  XOR U31564 ( .A(n31779), .B(n31768), .Z(n31723) );
  XNOR U31565 ( .A(n31780), .B(n31763), .Z(n31768) );
  XOR U31566 ( .A(n31781), .B(n31782), .Z(n31763) );
  AND U31567 ( .A(n31783), .B(n31784), .Z(n31782) );
  XOR U31568 ( .A(n31785), .B(n31781), .Z(n31783) );
  XNOR U31569 ( .A(n31786), .B(n31787), .Z(n31780) );
  AND U31570 ( .A(n31788), .B(n31789), .Z(n31787) );
  XOR U31571 ( .A(n31786), .B(n31790), .Z(n31788) );
  XNOR U31572 ( .A(n31769), .B(n31766), .Z(n31779) );
  AND U31573 ( .A(n31791), .B(n31792), .Z(n31766) );
  XOR U31574 ( .A(n31793), .B(n31794), .Z(n31769) );
  AND U31575 ( .A(n31795), .B(n31796), .Z(n31794) );
  XOR U31576 ( .A(n31793), .B(n31797), .Z(n31795) );
  XNOR U31577 ( .A(n31720), .B(n31775), .Z(n31777) );
  XNOR U31578 ( .A(n31798), .B(n31799), .Z(n31720) );
  AND U31579 ( .A(n325), .B(n31800), .Z(n31799) );
  XNOR U31580 ( .A(n31801), .B(n31802), .Z(n31800) );
  XOR U31581 ( .A(n31803), .B(n31804), .Z(n31775) );
  AND U31582 ( .A(n31805), .B(n31806), .Z(n31804) );
  XNOR U31583 ( .A(n31803), .B(n31791), .Z(n31806) );
  IV U31584 ( .A(n31733), .Z(n31791) );
  XNOR U31585 ( .A(n31807), .B(n31784), .Z(n31733) );
  XNOR U31586 ( .A(n31808), .B(n31790), .Z(n31784) );
  XOR U31587 ( .A(n31809), .B(n31810), .Z(n31790) );
  AND U31588 ( .A(n31811), .B(n31812), .Z(n31810) );
  XOR U31589 ( .A(n31809), .B(n31813), .Z(n31811) );
  XNOR U31590 ( .A(n31789), .B(n31781), .Z(n31808) );
  XOR U31591 ( .A(n31814), .B(n31815), .Z(n31781) );
  AND U31592 ( .A(n31816), .B(n31817), .Z(n31815) );
  XNOR U31593 ( .A(n31818), .B(n31814), .Z(n31816) );
  XNOR U31594 ( .A(n31819), .B(n31786), .Z(n31789) );
  XOR U31595 ( .A(n31820), .B(n31821), .Z(n31786) );
  AND U31596 ( .A(n31822), .B(n31823), .Z(n31821) );
  XOR U31597 ( .A(n31820), .B(n31824), .Z(n31822) );
  XNOR U31598 ( .A(n31825), .B(n31826), .Z(n31819) );
  AND U31599 ( .A(n31827), .B(n31828), .Z(n31826) );
  XNOR U31600 ( .A(n31825), .B(n31829), .Z(n31827) );
  XNOR U31601 ( .A(n31785), .B(n31792), .Z(n31807) );
  AND U31602 ( .A(n31741), .B(n31830), .Z(n31792) );
  XOR U31603 ( .A(n31797), .B(n31796), .Z(n31785) );
  XNOR U31604 ( .A(n31831), .B(n31793), .Z(n31796) );
  XOR U31605 ( .A(n31832), .B(n31833), .Z(n31793) );
  AND U31606 ( .A(n31834), .B(n31835), .Z(n31833) );
  XOR U31607 ( .A(n31832), .B(n31836), .Z(n31834) );
  XNOR U31608 ( .A(n31837), .B(n31838), .Z(n31831) );
  AND U31609 ( .A(n31839), .B(n31840), .Z(n31838) );
  XOR U31610 ( .A(n31837), .B(n31841), .Z(n31839) );
  XOR U31611 ( .A(n31842), .B(n31843), .Z(n31797) );
  AND U31612 ( .A(n31844), .B(n31845), .Z(n31843) );
  XOR U31613 ( .A(n31842), .B(n31846), .Z(n31844) );
  XNOR U31614 ( .A(n31730), .B(n31803), .Z(n31805) );
  XNOR U31615 ( .A(n31847), .B(n31848), .Z(n31730) );
  AND U31616 ( .A(n325), .B(n31849), .Z(n31848) );
  XNOR U31617 ( .A(n31850), .B(n31851), .Z(n31849) );
  XOR U31618 ( .A(n31852), .B(n31853), .Z(n31803) );
  AND U31619 ( .A(n31854), .B(n31855), .Z(n31853) );
  XNOR U31620 ( .A(n31852), .B(n31741), .Z(n31855) );
  XOR U31621 ( .A(n31856), .B(n31817), .Z(n31741) );
  XNOR U31622 ( .A(n31857), .B(n31824), .Z(n31817) );
  XOR U31623 ( .A(n31813), .B(n31812), .Z(n31824) );
  XNOR U31624 ( .A(n31858), .B(n31809), .Z(n31812) );
  XOR U31625 ( .A(n31859), .B(n31860), .Z(n31809) );
  AND U31626 ( .A(n31861), .B(n31862), .Z(n31860) );
  XOR U31627 ( .A(n31859), .B(n31863), .Z(n31861) );
  XNOR U31628 ( .A(n31864), .B(n31865), .Z(n31858) );
  NOR U31629 ( .A(n31866), .B(n31867), .Z(n31865) );
  XNOR U31630 ( .A(n31864), .B(n31868), .Z(n31866) );
  XOR U31631 ( .A(n31869), .B(n31870), .Z(n31813) );
  NOR U31632 ( .A(n31871), .B(n31872), .Z(n31870) );
  XNOR U31633 ( .A(n31869), .B(n31873), .Z(n31871) );
  XNOR U31634 ( .A(n31823), .B(n31814), .Z(n31857) );
  XOR U31635 ( .A(n31874), .B(n31875), .Z(n31814) );
  NOR U31636 ( .A(n31876), .B(n31877), .Z(n31875) );
  XNOR U31637 ( .A(n31874), .B(n31878), .Z(n31876) );
  XOR U31638 ( .A(n31879), .B(n31829), .Z(n31823) );
  XNOR U31639 ( .A(n31880), .B(n31881), .Z(n31829) );
  NOR U31640 ( .A(n31882), .B(n31883), .Z(n31881) );
  XNOR U31641 ( .A(n31880), .B(n31884), .Z(n31882) );
  XNOR U31642 ( .A(n31828), .B(n31820), .Z(n31879) );
  XOR U31643 ( .A(n31885), .B(n31886), .Z(n31820) );
  AND U31644 ( .A(n31887), .B(n31888), .Z(n31886) );
  XOR U31645 ( .A(n31885), .B(n31889), .Z(n31887) );
  XNOR U31646 ( .A(n31890), .B(n31825), .Z(n31828) );
  XOR U31647 ( .A(n31891), .B(n31892), .Z(n31825) );
  AND U31648 ( .A(n31893), .B(n31894), .Z(n31892) );
  XOR U31649 ( .A(n31891), .B(n31895), .Z(n31893) );
  XNOR U31650 ( .A(n31896), .B(n31897), .Z(n31890) );
  NOR U31651 ( .A(n31898), .B(n31899), .Z(n31897) );
  XOR U31652 ( .A(n31896), .B(n31900), .Z(n31898) );
  XOR U31653 ( .A(n31818), .B(n31830), .Z(n31856) );
  NOR U31654 ( .A(n31747), .B(n31901), .Z(n31830) );
  XNOR U31655 ( .A(n31836), .B(n31835), .Z(n31818) );
  XNOR U31656 ( .A(n31902), .B(n31841), .Z(n31835) );
  XOR U31657 ( .A(n31903), .B(n31904), .Z(n31841) );
  NOR U31658 ( .A(n31905), .B(n31906), .Z(n31904) );
  XNOR U31659 ( .A(n31903), .B(n31907), .Z(n31905) );
  XNOR U31660 ( .A(n31840), .B(n31832), .Z(n31902) );
  XOR U31661 ( .A(n31908), .B(n31909), .Z(n31832) );
  AND U31662 ( .A(n31910), .B(n31911), .Z(n31909) );
  XNOR U31663 ( .A(n31908), .B(n31912), .Z(n31910) );
  XNOR U31664 ( .A(n31913), .B(n31837), .Z(n31840) );
  XOR U31665 ( .A(n31914), .B(n31915), .Z(n31837) );
  AND U31666 ( .A(n31916), .B(n31917), .Z(n31915) );
  XOR U31667 ( .A(n31914), .B(n31918), .Z(n31916) );
  XNOR U31668 ( .A(n31919), .B(n31920), .Z(n31913) );
  NOR U31669 ( .A(n31921), .B(n31922), .Z(n31920) );
  XOR U31670 ( .A(n31919), .B(n31923), .Z(n31921) );
  XOR U31671 ( .A(n31846), .B(n31845), .Z(n31836) );
  XNOR U31672 ( .A(n31924), .B(n31842), .Z(n31845) );
  XOR U31673 ( .A(n31925), .B(n31926), .Z(n31842) );
  AND U31674 ( .A(n31927), .B(n31928), .Z(n31926) );
  XOR U31675 ( .A(n31925), .B(n31929), .Z(n31927) );
  XNOR U31676 ( .A(n31930), .B(n31931), .Z(n31924) );
  NOR U31677 ( .A(n31932), .B(n31933), .Z(n31931) );
  XNOR U31678 ( .A(n31930), .B(n31934), .Z(n31932) );
  XOR U31679 ( .A(n31935), .B(n31936), .Z(n31846) );
  NOR U31680 ( .A(n31937), .B(n31938), .Z(n31936) );
  XNOR U31681 ( .A(n31935), .B(n31939), .Z(n31937) );
  XNOR U31682 ( .A(n31738), .B(n31852), .Z(n31854) );
  XNOR U31683 ( .A(n31940), .B(n31941), .Z(n31738) );
  AND U31684 ( .A(n325), .B(n31942), .Z(n31941) );
  XNOR U31685 ( .A(n31943), .B(n31944), .Z(n31942) );
  AND U31686 ( .A(n31744), .B(n31747), .Z(n31852) );
  XOR U31687 ( .A(n31945), .B(n31901), .Z(n31747) );
  XNOR U31688 ( .A(p_input[2048]), .B(p_input[320]), .Z(n31901) );
  XOR U31689 ( .A(n31878), .B(n31877), .Z(n31945) );
  XOR U31690 ( .A(n31946), .B(n31889), .Z(n31877) );
  XOR U31691 ( .A(n31863), .B(n31862), .Z(n31889) );
  XNOR U31692 ( .A(n31947), .B(n31868), .Z(n31862) );
  XOR U31693 ( .A(p_input[2072]), .B(p_input[344]), .Z(n31868) );
  XOR U31694 ( .A(n31859), .B(n31867), .Z(n31947) );
  XOR U31695 ( .A(n31948), .B(n31864), .Z(n31867) );
  XOR U31696 ( .A(p_input[2070]), .B(p_input[342]), .Z(n31864) );
  XNOR U31697 ( .A(p_input[2071]), .B(p_input[343]), .Z(n31948) );
  XNOR U31698 ( .A(n28684), .B(p_input[338]), .Z(n31859) );
  XNOR U31699 ( .A(n31873), .B(n31872), .Z(n31863) );
  XOR U31700 ( .A(n31949), .B(n31869), .Z(n31872) );
  XOR U31701 ( .A(p_input[2067]), .B(p_input[339]), .Z(n31869) );
  XNOR U31702 ( .A(p_input[2068]), .B(p_input[340]), .Z(n31949) );
  XOR U31703 ( .A(p_input[2069]), .B(p_input[341]), .Z(n31873) );
  XNOR U31704 ( .A(n31888), .B(n31874), .Z(n31946) );
  XNOR U31705 ( .A(n28686), .B(p_input[321]), .Z(n31874) );
  XNOR U31706 ( .A(n31950), .B(n31895), .Z(n31888) );
  XNOR U31707 ( .A(n31884), .B(n31883), .Z(n31895) );
  XOR U31708 ( .A(n31951), .B(n31880), .Z(n31883) );
  XNOR U31709 ( .A(n28322), .B(p_input[346]), .Z(n31880) );
  XNOR U31710 ( .A(p_input[2075]), .B(p_input[347]), .Z(n31951) );
  XOR U31711 ( .A(p_input[2076]), .B(p_input[348]), .Z(n31884) );
  XNOR U31712 ( .A(n31894), .B(n31885), .Z(n31950) );
  XNOR U31713 ( .A(n28689), .B(p_input[337]), .Z(n31885) );
  XOR U31714 ( .A(n31952), .B(n31900), .Z(n31894) );
  XNOR U31715 ( .A(p_input[2079]), .B(p_input[351]), .Z(n31900) );
  XOR U31716 ( .A(n31891), .B(n31899), .Z(n31952) );
  XOR U31717 ( .A(n31953), .B(n31896), .Z(n31899) );
  XOR U31718 ( .A(p_input[2077]), .B(p_input[349]), .Z(n31896) );
  XNOR U31719 ( .A(p_input[2078]), .B(p_input[350]), .Z(n31953) );
  XNOR U31720 ( .A(n28326), .B(p_input[345]), .Z(n31891) );
  XNOR U31721 ( .A(n31912), .B(n31911), .Z(n31878) );
  XNOR U31722 ( .A(n31954), .B(n31918), .Z(n31911) );
  XNOR U31723 ( .A(n31907), .B(n31906), .Z(n31918) );
  XOR U31724 ( .A(n31955), .B(n31903), .Z(n31906) );
  XNOR U31725 ( .A(n28694), .B(p_input[331]), .Z(n31903) );
  XNOR U31726 ( .A(p_input[2060]), .B(p_input[332]), .Z(n31955) );
  XOR U31727 ( .A(p_input[2061]), .B(p_input[333]), .Z(n31907) );
  XNOR U31728 ( .A(n31917), .B(n31908), .Z(n31954) );
  XNOR U31729 ( .A(n28330), .B(p_input[322]), .Z(n31908) );
  XOR U31730 ( .A(n31956), .B(n31923), .Z(n31917) );
  XNOR U31731 ( .A(p_input[2064]), .B(p_input[336]), .Z(n31923) );
  XOR U31732 ( .A(n31914), .B(n31922), .Z(n31956) );
  XOR U31733 ( .A(n31957), .B(n31919), .Z(n31922) );
  XOR U31734 ( .A(p_input[2062]), .B(p_input[334]), .Z(n31919) );
  XNOR U31735 ( .A(p_input[2063]), .B(p_input[335]), .Z(n31957) );
  XNOR U31736 ( .A(n28697), .B(p_input[330]), .Z(n31914) );
  XNOR U31737 ( .A(n31929), .B(n31928), .Z(n31912) );
  XNOR U31738 ( .A(n31958), .B(n31934), .Z(n31928) );
  XOR U31739 ( .A(p_input[2057]), .B(p_input[329]), .Z(n31934) );
  XOR U31740 ( .A(n31925), .B(n31933), .Z(n31958) );
  XOR U31741 ( .A(n31959), .B(n31930), .Z(n31933) );
  XOR U31742 ( .A(p_input[2055]), .B(p_input[327]), .Z(n31930) );
  XNOR U31743 ( .A(p_input[2056]), .B(p_input[328]), .Z(n31959) );
  XNOR U31744 ( .A(n28337), .B(p_input[323]), .Z(n31925) );
  XNOR U31745 ( .A(n31939), .B(n31938), .Z(n31929) );
  XOR U31746 ( .A(n31960), .B(n31935), .Z(n31938) );
  XOR U31747 ( .A(p_input[2052]), .B(p_input[324]), .Z(n31935) );
  XNOR U31748 ( .A(p_input[2053]), .B(p_input[325]), .Z(n31960) );
  XOR U31749 ( .A(p_input[2054]), .B(p_input[326]), .Z(n31939) );
  XNOR U31750 ( .A(n31961), .B(n31962), .Z(n31744) );
  AND U31751 ( .A(n325), .B(n31963), .Z(n31962) );
  XNOR U31752 ( .A(n31964), .B(n31965), .Z(n325) );
  AND U31753 ( .A(n31966), .B(n31967), .Z(n31965) );
  XOR U31754 ( .A(n31758), .B(n31964), .Z(n31967) );
  XNOR U31755 ( .A(n31968), .B(n31964), .Z(n31966) );
  XOR U31756 ( .A(n31969), .B(n31970), .Z(n31964) );
  AND U31757 ( .A(n31971), .B(n31972), .Z(n31970) );
  XOR U31758 ( .A(n31773), .B(n31969), .Z(n31972) );
  XOR U31759 ( .A(n31969), .B(n31774), .Z(n31971) );
  XOR U31760 ( .A(n31973), .B(n31974), .Z(n31969) );
  AND U31761 ( .A(n31975), .B(n31976), .Z(n31974) );
  XOR U31762 ( .A(n31801), .B(n31973), .Z(n31976) );
  XOR U31763 ( .A(n31973), .B(n31802), .Z(n31975) );
  XOR U31764 ( .A(n31977), .B(n31978), .Z(n31973) );
  AND U31765 ( .A(n31979), .B(n31980), .Z(n31978) );
  XOR U31766 ( .A(n31850), .B(n31977), .Z(n31980) );
  XOR U31767 ( .A(n31977), .B(n31851), .Z(n31979) );
  XOR U31768 ( .A(n31981), .B(n31982), .Z(n31977) );
  AND U31769 ( .A(n31983), .B(n31984), .Z(n31982) );
  XOR U31770 ( .A(n31981), .B(n31943), .Z(n31984) );
  XNOR U31771 ( .A(n31985), .B(n31986), .Z(n31694) );
  AND U31772 ( .A(n329), .B(n31987), .Z(n31986) );
  XNOR U31773 ( .A(n31988), .B(n31989), .Z(n329) );
  AND U31774 ( .A(n31990), .B(n31991), .Z(n31989) );
  XOR U31775 ( .A(n31988), .B(n31704), .Z(n31991) );
  XNOR U31776 ( .A(n31988), .B(n31654), .Z(n31990) );
  XOR U31777 ( .A(n31992), .B(n31993), .Z(n31988) );
  AND U31778 ( .A(n31994), .B(n31995), .Z(n31993) );
  XNOR U31779 ( .A(n31714), .B(n31992), .Z(n31995) );
  XOR U31780 ( .A(n31992), .B(n31664), .Z(n31994) );
  XOR U31781 ( .A(n31996), .B(n31997), .Z(n31992) );
  AND U31782 ( .A(n31998), .B(n31999), .Z(n31997) );
  XNOR U31783 ( .A(n31724), .B(n31996), .Z(n31999) );
  XOR U31784 ( .A(n31996), .B(n31673), .Z(n31998) );
  XOR U31785 ( .A(n32000), .B(n32001), .Z(n31996) );
  AND U31786 ( .A(n32002), .B(n32003), .Z(n32001) );
  XOR U31787 ( .A(n32000), .B(n31681), .Z(n32002) );
  XOR U31788 ( .A(n32004), .B(n32005), .Z(n31645) );
  AND U31789 ( .A(n333), .B(n31987), .Z(n32005) );
  XNOR U31790 ( .A(n31985), .B(n32004), .Z(n31987) );
  XNOR U31791 ( .A(n32006), .B(n32007), .Z(n333) );
  AND U31792 ( .A(n32008), .B(n32009), .Z(n32007) );
  XNOR U31793 ( .A(n32010), .B(n32006), .Z(n32009) );
  IV U31794 ( .A(n31704), .Z(n32010) );
  XOR U31795 ( .A(n31968), .B(n32011), .Z(n31704) );
  AND U31796 ( .A(n336), .B(n32012), .Z(n32011) );
  XOR U31797 ( .A(n31757), .B(n31754), .Z(n32012) );
  IV U31798 ( .A(n31968), .Z(n31757) );
  XNOR U31799 ( .A(n31654), .B(n32006), .Z(n32008) );
  XOR U31800 ( .A(n32013), .B(n32014), .Z(n31654) );
  AND U31801 ( .A(n352), .B(n32015), .Z(n32014) );
  XOR U31802 ( .A(n32016), .B(n32017), .Z(n32006) );
  AND U31803 ( .A(n32018), .B(n32019), .Z(n32017) );
  XNOR U31804 ( .A(n32016), .B(n31714), .Z(n32019) );
  XOR U31805 ( .A(n31774), .B(n32020), .Z(n31714) );
  AND U31806 ( .A(n336), .B(n32021), .Z(n32020) );
  XOR U31807 ( .A(n31770), .B(n31774), .Z(n32021) );
  XNOR U31808 ( .A(n32022), .B(n32016), .Z(n32018) );
  IV U31809 ( .A(n31664), .Z(n32022) );
  XOR U31810 ( .A(n32023), .B(n32024), .Z(n31664) );
  AND U31811 ( .A(n352), .B(n32025), .Z(n32024) );
  XOR U31812 ( .A(n32026), .B(n32027), .Z(n32016) );
  AND U31813 ( .A(n32028), .B(n32029), .Z(n32027) );
  XNOR U31814 ( .A(n32026), .B(n31724), .Z(n32029) );
  XOR U31815 ( .A(n31802), .B(n32030), .Z(n31724) );
  AND U31816 ( .A(n336), .B(n32031), .Z(n32030) );
  XOR U31817 ( .A(n31798), .B(n31802), .Z(n32031) );
  XOR U31818 ( .A(n31673), .B(n32026), .Z(n32028) );
  XOR U31819 ( .A(n32032), .B(n32033), .Z(n31673) );
  AND U31820 ( .A(n352), .B(n32034), .Z(n32033) );
  XOR U31821 ( .A(n32000), .B(n32035), .Z(n32026) );
  AND U31822 ( .A(n32036), .B(n32003), .Z(n32035) );
  XNOR U31823 ( .A(n31734), .B(n32000), .Z(n32003) );
  XOR U31824 ( .A(n31851), .B(n32037), .Z(n31734) );
  AND U31825 ( .A(n336), .B(n32038), .Z(n32037) );
  XOR U31826 ( .A(n31847), .B(n31851), .Z(n32038) );
  XNOR U31827 ( .A(n32039), .B(n32000), .Z(n32036) );
  IV U31828 ( .A(n31681), .Z(n32039) );
  XOR U31829 ( .A(n32040), .B(n32041), .Z(n31681) );
  AND U31830 ( .A(n352), .B(n32042), .Z(n32041) );
  XOR U31831 ( .A(n32043), .B(n32044), .Z(n32000) );
  AND U31832 ( .A(n32045), .B(n32046), .Z(n32044) );
  XNOR U31833 ( .A(n32043), .B(n31742), .Z(n32046) );
  XOR U31834 ( .A(n31944), .B(n32047), .Z(n31742) );
  AND U31835 ( .A(n336), .B(n32048), .Z(n32047) );
  XOR U31836 ( .A(n31940), .B(n31944), .Z(n32048) );
  XNOR U31837 ( .A(n32049), .B(n32043), .Z(n32045) );
  IV U31838 ( .A(n31691), .Z(n32049) );
  XOR U31839 ( .A(n32050), .B(n32051), .Z(n31691) );
  AND U31840 ( .A(n352), .B(n32052), .Z(n32051) );
  AND U31841 ( .A(n32004), .B(n31985), .Z(n32043) );
  XNOR U31842 ( .A(n32053), .B(n32054), .Z(n31985) );
  AND U31843 ( .A(n336), .B(n31963), .Z(n32054) );
  XNOR U31844 ( .A(n31961), .B(n32053), .Z(n31963) );
  XNOR U31845 ( .A(n32055), .B(n32056), .Z(n336) );
  AND U31846 ( .A(n32057), .B(n32058), .Z(n32056) );
  XNOR U31847 ( .A(n32055), .B(n31754), .Z(n32058) );
  IV U31848 ( .A(n31758), .Z(n31754) );
  XOR U31849 ( .A(n32059), .B(n32060), .Z(n31758) );
  AND U31850 ( .A(n340), .B(n32061), .Z(n32060) );
  XOR U31851 ( .A(n32062), .B(n32059), .Z(n32061) );
  XNOR U31852 ( .A(n32055), .B(n31968), .Z(n32057) );
  XOR U31853 ( .A(n32063), .B(n32064), .Z(n31968) );
  AND U31854 ( .A(n348), .B(n32015), .Z(n32064) );
  XOR U31855 ( .A(n32013), .B(n32063), .Z(n32015) );
  XOR U31856 ( .A(n32065), .B(n32066), .Z(n32055) );
  AND U31857 ( .A(n32067), .B(n32068), .Z(n32066) );
  XNOR U31858 ( .A(n32065), .B(n31770), .Z(n32068) );
  IV U31859 ( .A(n31773), .Z(n31770) );
  XOR U31860 ( .A(n32069), .B(n32070), .Z(n31773) );
  AND U31861 ( .A(n340), .B(n32071), .Z(n32070) );
  XOR U31862 ( .A(n32072), .B(n32069), .Z(n32071) );
  XOR U31863 ( .A(n31774), .B(n32065), .Z(n32067) );
  XOR U31864 ( .A(n32073), .B(n32074), .Z(n31774) );
  AND U31865 ( .A(n348), .B(n32025), .Z(n32074) );
  XOR U31866 ( .A(n32073), .B(n32023), .Z(n32025) );
  XOR U31867 ( .A(n32075), .B(n32076), .Z(n32065) );
  AND U31868 ( .A(n32077), .B(n32078), .Z(n32076) );
  XNOR U31869 ( .A(n32075), .B(n31798), .Z(n32078) );
  IV U31870 ( .A(n31801), .Z(n31798) );
  XOR U31871 ( .A(n32079), .B(n32080), .Z(n31801) );
  AND U31872 ( .A(n340), .B(n32081), .Z(n32080) );
  XNOR U31873 ( .A(n32082), .B(n32079), .Z(n32081) );
  XOR U31874 ( .A(n31802), .B(n32075), .Z(n32077) );
  XOR U31875 ( .A(n32083), .B(n32084), .Z(n31802) );
  AND U31876 ( .A(n348), .B(n32034), .Z(n32084) );
  XOR U31877 ( .A(n32083), .B(n32032), .Z(n32034) );
  XOR U31878 ( .A(n32085), .B(n32086), .Z(n32075) );
  AND U31879 ( .A(n32087), .B(n32088), .Z(n32086) );
  XNOR U31880 ( .A(n32085), .B(n31847), .Z(n32088) );
  IV U31881 ( .A(n31850), .Z(n31847) );
  XOR U31882 ( .A(n32089), .B(n32090), .Z(n31850) );
  AND U31883 ( .A(n340), .B(n32091), .Z(n32090) );
  XOR U31884 ( .A(n32092), .B(n32089), .Z(n32091) );
  XOR U31885 ( .A(n31851), .B(n32085), .Z(n32087) );
  XOR U31886 ( .A(n32093), .B(n32094), .Z(n31851) );
  AND U31887 ( .A(n348), .B(n32042), .Z(n32094) );
  XOR U31888 ( .A(n32093), .B(n32040), .Z(n32042) );
  XOR U31889 ( .A(n31981), .B(n32095), .Z(n32085) );
  AND U31890 ( .A(n31983), .B(n32096), .Z(n32095) );
  XNOR U31891 ( .A(n31981), .B(n31940), .Z(n32096) );
  IV U31892 ( .A(n31943), .Z(n31940) );
  XOR U31893 ( .A(n32097), .B(n32098), .Z(n31943) );
  AND U31894 ( .A(n340), .B(n32099), .Z(n32098) );
  XNOR U31895 ( .A(n32100), .B(n32097), .Z(n32099) );
  XOR U31896 ( .A(n31944), .B(n31981), .Z(n31983) );
  XOR U31897 ( .A(n32101), .B(n32102), .Z(n31944) );
  AND U31898 ( .A(n348), .B(n32052), .Z(n32102) );
  XOR U31899 ( .A(n32101), .B(n32050), .Z(n32052) );
  AND U31900 ( .A(n32053), .B(n31961), .Z(n31981) );
  XNOR U31901 ( .A(n32103), .B(n32104), .Z(n31961) );
  AND U31902 ( .A(n340), .B(n32105), .Z(n32104) );
  XNOR U31903 ( .A(n32106), .B(n32103), .Z(n32105) );
  XNOR U31904 ( .A(n32107), .B(n32108), .Z(n340) );
  AND U31905 ( .A(n32109), .B(n32110), .Z(n32108) );
  XOR U31906 ( .A(n32062), .B(n32107), .Z(n32110) );
  AND U31907 ( .A(n32111), .B(n32112), .Z(n32062) );
  XNOR U31908 ( .A(n32059), .B(n32107), .Z(n32109) );
  XNOR U31909 ( .A(n32113), .B(n32114), .Z(n32059) );
  AND U31910 ( .A(n344), .B(n32115), .Z(n32114) );
  XNOR U31911 ( .A(n32116), .B(n32117), .Z(n32115) );
  XOR U31912 ( .A(n32118), .B(n32119), .Z(n32107) );
  AND U31913 ( .A(n32120), .B(n32121), .Z(n32119) );
  XNOR U31914 ( .A(n32118), .B(n32111), .Z(n32121) );
  IV U31915 ( .A(n32072), .Z(n32111) );
  XOR U31916 ( .A(n32122), .B(n32123), .Z(n32072) );
  XOR U31917 ( .A(n32124), .B(n32112), .Z(n32123) );
  AND U31918 ( .A(n32082), .B(n32125), .Z(n32112) );
  AND U31919 ( .A(n32126), .B(n32127), .Z(n32124) );
  XOR U31920 ( .A(n32128), .B(n32122), .Z(n32126) );
  XNOR U31921 ( .A(n32069), .B(n32118), .Z(n32120) );
  XNOR U31922 ( .A(n32129), .B(n32130), .Z(n32069) );
  AND U31923 ( .A(n344), .B(n32131), .Z(n32130) );
  XNOR U31924 ( .A(n32132), .B(n32133), .Z(n32131) );
  XOR U31925 ( .A(n32134), .B(n32135), .Z(n32118) );
  AND U31926 ( .A(n32136), .B(n32137), .Z(n32135) );
  XNOR U31927 ( .A(n32134), .B(n32082), .Z(n32137) );
  XOR U31928 ( .A(n32138), .B(n32127), .Z(n32082) );
  XNOR U31929 ( .A(n32139), .B(n32122), .Z(n32127) );
  XOR U31930 ( .A(n32140), .B(n32141), .Z(n32122) );
  AND U31931 ( .A(n32142), .B(n32143), .Z(n32141) );
  XOR U31932 ( .A(n32144), .B(n32140), .Z(n32142) );
  XNOR U31933 ( .A(n32145), .B(n32146), .Z(n32139) );
  AND U31934 ( .A(n32147), .B(n32148), .Z(n32146) );
  XOR U31935 ( .A(n32145), .B(n32149), .Z(n32147) );
  XNOR U31936 ( .A(n32128), .B(n32125), .Z(n32138) );
  AND U31937 ( .A(n32150), .B(n32151), .Z(n32125) );
  XOR U31938 ( .A(n32152), .B(n32153), .Z(n32128) );
  AND U31939 ( .A(n32154), .B(n32155), .Z(n32153) );
  XOR U31940 ( .A(n32152), .B(n32156), .Z(n32154) );
  XNOR U31941 ( .A(n32079), .B(n32134), .Z(n32136) );
  XNOR U31942 ( .A(n32157), .B(n32158), .Z(n32079) );
  AND U31943 ( .A(n344), .B(n32159), .Z(n32158) );
  XNOR U31944 ( .A(n32160), .B(n32161), .Z(n32159) );
  XOR U31945 ( .A(n32162), .B(n32163), .Z(n32134) );
  AND U31946 ( .A(n32164), .B(n32165), .Z(n32163) );
  XNOR U31947 ( .A(n32162), .B(n32150), .Z(n32165) );
  IV U31948 ( .A(n32092), .Z(n32150) );
  XNOR U31949 ( .A(n32166), .B(n32143), .Z(n32092) );
  XNOR U31950 ( .A(n32167), .B(n32149), .Z(n32143) );
  XOR U31951 ( .A(n32168), .B(n32169), .Z(n32149) );
  AND U31952 ( .A(n32170), .B(n32171), .Z(n32169) );
  XOR U31953 ( .A(n32168), .B(n32172), .Z(n32170) );
  XNOR U31954 ( .A(n32148), .B(n32140), .Z(n32167) );
  XOR U31955 ( .A(n32173), .B(n32174), .Z(n32140) );
  AND U31956 ( .A(n32175), .B(n32176), .Z(n32174) );
  XNOR U31957 ( .A(n32177), .B(n32173), .Z(n32175) );
  XNOR U31958 ( .A(n32178), .B(n32145), .Z(n32148) );
  XOR U31959 ( .A(n32179), .B(n32180), .Z(n32145) );
  AND U31960 ( .A(n32181), .B(n32182), .Z(n32180) );
  XOR U31961 ( .A(n32179), .B(n32183), .Z(n32181) );
  XNOR U31962 ( .A(n32184), .B(n32185), .Z(n32178) );
  AND U31963 ( .A(n32186), .B(n32187), .Z(n32185) );
  XNOR U31964 ( .A(n32184), .B(n32188), .Z(n32186) );
  XNOR U31965 ( .A(n32144), .B(n32151), .Z(n32166) );
  AND U31966 ( .A(n32100), .B(n32189), .Z(n32151) );
  XOR U31967 ( .A(n32156), .B(n32155), .Z(n32144) );
  XNOR U31968 ( .A(n32190), .B(n32152), .Z(n32155) );
  XOR U31969 ( .A(n32191), .B(n32192), .Z(n32152) );
  AND U31970 ( .A(n32193), .B(n32194), .Z(n32192) );
  XOR U31971 ( .A(n32191), .B(n32195), .Z(n32193) );
  XNOR U31972 ( .A(n32196), .B(n32197), .Z(n32190) );
  AND U31973 ( .A(n32198), .B(n32199), .Z(n32197) );
  XOR U31974 ( .A(n32196), .B(n32200), .Z(n32198) );
  XOR U31975 ( .A(n32201), .B(n32202), .Z(n32156) );
  AND U31976 ( .A(n32203), .B(n32204), .Z(n32202) );
  XOR U31977 ( .A(n32201), .B(n32205), .Z(n32203) );
  XNOR U31978 ( .A(n32089), .B(n32162), .Z(n32164) );
  XNOR U31979 ( .A(n32206), .B(n32207), .Z(n32089) );
  AND U31980 ( .A(n344), .B(n32208), .Z(n32207) );
  XNOR U31981 ( .A(n32209), .B(n32210), .Z(n32208) );
  XOR U31982 ( .A(n32211), .B(n32212), .Z(n32162) );
  AND U31983 ( .A(n32213), .B(n32214), .Z(n32212) );
  XNOR U31984 ( .A(n32211), .B(n32100), .Z(n32214) );
  XOR U31985 ( .A(n32215), .B(n32176), .Z(n32100) );
  XNOR U31986 ( .A(n32216), .B(n32183), .Z(n32176) );
  XOR U31987 ( .A(n32172), .B(n32171), .Z(n32183) );
  XNOR U31988 ( .A(n32217), .B(n32168), .Z(n32171) );
  XOR U31989 ( .A(n32218), .B(n32219), .Z(n32168) );
  AND U31990 ( .A(n32220), .B(n32221), .Z(n32219) );
  XOR U31991 ( .A(n32218), .B(n32222), .Z(n32220) );
  XNOR U31992 ( .A(n32223), .B(n32224), .Z(n32217) );
  NOR U31993 ( .A(n32225), .B(n32226), .Z(n32224) );
  XNOR U31994 ( .A(n32223), .B(n32227), .Z(n32225) );
  XOR U31995 ( .A(n32228), .B(n32229), .Z(n32172) );
  NOR U31996 ( .A(n32230), .B(n32231), .Z(n32229) );
  XNOR U31997 ( .A(n32228), .B(n32232), .Z(n32230) );
  XNOR U31998 ( .A(n32182), .B(n32173), .Z(n32216) );
  XOR U31999 ( .A(n32233), .B(n32234), .Z(n32173) );
  NOR U32000 ( .A(n32235), .B(n32236), .Z(n32234) );
  XNOR U32001 ( .A(n32233), .B(n32237), .Z(n32235) );
  XOR U32002 ( .A(n32238), .B(n32188), .Z(n32182) );
  XNOR U32003 ( .A(n32239), .B(n32240), .Z(n32188) );
  NOR U32004 ( .A(n32241), .B(n32242), .Z(n32240) );
  XNOR U32005 ( .A(n32239), .B(n32243), .Z(n32241) );
  XNOR U32006 ( .A(n32187), .B(n32179), .Z(n32238) );
  XOR U32007 ( .A(n32244), .B(n32245), .Z(n32179) );
  AND U32008 ( .A(n32246), .B(n32247), .Z(n32245) );
  XOR U32009 ( .A(n32244), .B(n32248), .Z(n32246) );
  XNOR U32010 ( .A(n32249), .B(n32184), .Z(n32187) );
  XOR U32011 ( .A(n32250), .B(n32251), .Z(n32184) );
  AND U32012 ( .A(n32252), .B(n32253), .Z(n32251) );
  XOR U32013 ( .A(n32250), .B(n32254), .Z(n32252) );
  XNOR U32014 ( .A(n32255), .B(n32256), .Z(n32249) );
  NOR U32015 ( .A(n32257), .B(n32258), .Z(n32256) );
  XOR U32016 ( .A(n32255), .B(n32259), .Z(n32257) );
  XOR U32017 ( .A(n32177), .B(n32189), .Z(n32215) );
  NOR U32018 ( .A(n32106), .B(n32260), .Z(n32189) );
  XNOR U32019 ( .A(n32195), .B(n32194), .Z(n32177) );
  XNOR U32020 ( .A(n32261), .B(n32200), .Z(n32194) );
  XOR U32021 ( .A(n32262), .B(n32263), .Z(n32200) );
  NOR U32022 ( .A(n32264), .B(n32265), .Z(n32263) );
  XNOR U32023 ( .A(n32262), .B(n32266), .Z(n32264) );
  XNOR U32024 ( .A(n32199), .B(n32191), .Z(n32261) );
  XOR U32025 ( .A(n32267), .B(n32268), .Z(n32191) );
  AND U32026 ( .A(n32269), .B(n32270), .Z(n32268) );
  XNOR U32027 ( .A(n32267), .B(n32271), .Z(n32269) );
  XNOR U32028 ( .A(n32272), .B(n32196), .Z(n32199) );
  XOR U32029 ( .A(n32273), .B(n32274), .Z(n32196) );
  AND U32030 ( .A(n32275), .B(n32276), .Z(n32274) );
  XOR U32031 ( .A(n32273), .B(n32277), .Z(n32275) );
  XNOR U32032 ( .A(n32278), .B(n32279), .Z(n32272) );
  NOR U32033 ( .A(n32280), .B(n32281), .Z(n32279) );
  XOR U32034 ( .A(n32278), .B(n32282), .Z(n32280) );
  XOR U32035 ( .A(n32205), .B(n32204), .Z(n32195) );
  XNOR U32036 ( .A(n32283), .B(n32201), .Z(n32204) );
  XOR U32037 ( .A(n32284), .B(n32285), .Z(n32201) );
  AND U32038 ( .A(n32286), .B(n32287), .Z(n32285) );
  XOR U32039 ( .A(n32284), .B(n32288), .Z(n32286) );
  XNOR U32040 ( .A(n32289), .B(n32290), .Z(n32283) );
  NOR U32041 ( .A(n32291), .B(n32292), .Z(n32290) );
  XNOR U32042 ( .A(n32289), .B(n32293), .Z(n32291) );
  XOR U32043 ( .A(n32294), .B(n32295), .Z(n32205) );
  NOR U32044 ( .A(n32296), .B(n32297), .Z(n32295) );
  XNOR U32045 ( .A(n32294), .B(n32298), .Z(n32296) );
  XNOR U32046 ( .A(n32097), .B(n32211), .Z(n32213) );
  XNOR U32047 ( .A(n32299), .B(n32300), .Z(n32097) );
  AND U32048 ( .A(n344), .B(n32301), .Z(n32300) );
  XNOR U32049 ( .A(n32302), .B(n32303), .Z(n32301) );
  AND U32050 ( .A(n32103), .B(n32106), .Z(n32211) );
  XOR U32051 ( .A(n32304), .B(n32260), .Z(n32106) );
  XNOR U32052 ( .A(p_input[2048]), .B(p_input[352]), .Z(n32260) );
  XOR U32053 ( .A(n32237), .B(n32236), .Z(n32304) );
  XOR U32054 ( .A(n32305), .B(n32248), .Z(n32236) );
  XOR U32055 ( .A(n32222), .B(n32221), .Z(n32248) );
  XNOR U32056 ( .A(n32306), .B(n32227), .Z(n32221) );
  XOR U32057 ( .A(p_input[2072]), .B(p_input[376]), .Z(n32227) );
  XOR U32058 ( .A(n32218), .B(n32226), .Z(n32306) );
  XOR U32059 ( .A(n32307), .B(n32223), .Z(n32226) );
  XOR U32060 ( .A(p_input[2070]), .B(p_input[374]), .Z(n32223) );
  XNOR U32061 ( .A(p_input[2071]), .B(p_input[375]), .Z(n32307) );
  XNOR U32062 ( .A(n28684), .B(p_input[370]), .Z(n32218) );
  XNOR U32063 ( .A(n32232), .B(n32231), .Z(n32222) );
  XOR U32064 ( .A(n32308), .B(n32228), .Z(n32231) );
  XOR U32065 ( .A(p_input[2067]), .B(p_input[371]), .Z(n32228) );
  XNOR U32066 ( .A(p_input[2068]), .B(p_input[372]), .Z(n32308) );
  XOR U32067 ( .A(p_input[2069]), .B(p_input[373]), .Z(n32232) );
  XNOR U32068 ( .A(n32247), .B(n32233), .Z(n32305) );
  XNOR U32069 ( .A(n28686), .B(p_input[353]), .Z(n32233) );
  XNOR U32070 ( .A(n32309), .B(n32254), .Z(n32247) );
  XNOR U32071 ( .A(n32243), .B(n32242), .Z(n32254) );
  XOR U32072 ( .A(n32310), .B(n32239), .Z(n32242) );
  XNOR U32073 ( .A(n28322), .B(p_input[378]), .Z(n32239) );
  XNOR U32074 ( .A(p_input[2075]), .B(p_input[379]), .Z(n32310) );
  XOR U32075 ( .A(p_input[2076]), .B(p_input[380]), .Z(n32243) );
  XNOR U32076 ( .A(n32253), .B(n32244), .Z(n32309) );
  XNOR U32077 ( .A(n28689), .B(p_input[369]), .Z(n32244) );
  XOR U32078 ( .A(n32311), .B(n32259), .Z(n32253) );
  XNOR U32079 ( .A(p_input[2079]), .B(p_input[383]), .Z(n32259) );
  XOR U32080 ( .A(n32250), .B(n32258), .Z(n32311) );
  XOR U32081 ( .A(n32312), .B(n32255), .Z(n32258) );
  XOR U32082 ( .A(p_input[2077]), .B(p_input[381]), .Z(n32255) );
  XNOR U32083 ( .A(p_input[2078]), .B(p_input[382]), .Z(n32312) );
  XNOR U32084 ( .A(n28326), .B(p_input[377]), .Z(n32250) );
  XNOR U32085 ( .A(n32271), .B(n32270), .Z(n32237) );
  XNOR U32086 ( .A(n32313), .B(n32277), .Z(n32270) );
  XNOR U32087 ( .A(n32266), .B(n32265), .Z(n32277) );
  XOR U32088 ( .A(n32314), .B(n32262), .Z(n32265) );
  XNOR U32089 ( .A(n28694), .B(p_input[363]), .Z(n32262) );
  XNOR U32090 ( .A(p_input[2060]), .B(p_input[364]), .Z(n32314) );
  XOR U32091 ( .A(p_input[2061]), .B(p_input[365]), .Z(n32266) );
  XNOR U32092 ( .A(n32276), .B(n32267), .Z(n32313) );
  XNOR U32093 ( .A(n28330), .B(p_input[354]), .Z(n32267) );
  XOR U32094 ( .A(n32315), .B(n32282), .Z(n32276) );
  XNOR U32095 ( .A(p_input[2064]), .B(p_input[368]), .Z(n32282) );
  XOR U32096 ( .A(n32273), .B(n32281), .Z(n32315) );
  XOR U32097 ( .A(n32316), .B(n32278), .Z(n32281) );
  XOR U32098 ( .A(p_input[2062]), .B(p_input[366]), .Z(n32278) );
  XNOR U32099 ( .A(p_input[2063]), .B(p_input[367]), .Z(n32316) );
  XNOR U32100 ( .A(n28697), .B(p_input[362]), .Z(n32273) );
  XNOR U32101 ( .A(n32288), .B(n32287), .Z(n32271) );
  XNOR U32102 ( .A(n32317), .B(n32293), .Z(n32287) );
  XOR U32103 ( .A(p_input[2057]), .B(p_input[361]), .Z(n32293) );
  XOR U32104 ( .A(n32284), .B(n32292), .Z(n32317) );
  XOR U32105 ( .A(n32318), .B(n32289), .Z(n32292) );
  XOR U32106 ( .A(p_input[2055]), .B(p_input[359]), .Z(n32289) );
  XNOR U32107 ( .A(p_input[2056]), .B(p_input[360]), .Z(n32318) );
  XNOR U32108 ( .A(n28337), .B(p_input[355]), .Z(n32284) );
  XNOR U32109 ( .A(n32298), .B(n32297), .Z(n32288) );
  XOR U32110 ( .A(n32319), .B(n32294), .Z(n32297) );
  XOR U32111 ( .A(p_input[2052]), .B(p_input[356]), .Z(n32294) );
  XNOR U32112 ( .A(p_input[2053]), .B(p_input[357]), .Z(n32319) );
  XOR U32113 ( .A(p_input[2054]), .B(p_input[358]), .Z(n32298) );
  XNOR U32114 ( .A(n32320), .B(n32321), .Z(n32103) );
  AND U32115 ( .A(n344), .B(n32322), .Z(n32321) );
  XNOR U32116 ( .A(n32323), .B(n32324), .Z(n344) );
  AND U32117 ( .A(n32325), .B(n32326), .Z(n32324) );
  XOR U32118 ( .A(n32117), .B(n32323), .Z(n32326) );
  XNOR U32119 ( .A(n32327), .B(n32323), .Z(n32325) );
  XOR U32120 ( .A(n32328), .B(n32329), .Z(n32323) );
  AND U32121 ( .A(n32330), .B(n32331), .Z(n32329) );
  XOR U32122 ( .A(n32132), .B(n32328), .Z(n32331) );
  XOR U32123 ( .A(n32328), .B(n32133), .Z(n32330) );
  XOR U32124 ( .A(n32332), .B(n32333), .Z(n32328) );
  AND U32125 ( .A(n32334), .B(n32335), .Z(n32333) );
  XOR U32126 ( .A(n32160), .B(n32332), .Z(n32335) );
  XOR U32127 ( .A(n32332), .B(n32161), .Z(n32334) );
  XOR U32128 ( .A(n32336), .B(n32337), .Z(n32332) );
  AND U32129 ( .A(n32338), .B(n32339), .Z(n32337) );
  XOR U32130 ( .A(n32209), .B(n32336), .Z(n32339) );
  XOR U32131 ( .A(n32336), .B(n32210), .Z(n32338) );
  XOR U32132 ( .A(n32340), .B(n32341), .Z(n32336) );
  AND U32133 ( .A(n32342), .B(n32343), .Z(n32341) );
  XOR U32134 ( .A(n32340), .B(n32302), .Z(n32343) );
  XNOR U32135 ( .A(n32344), .B(n32345), .Z(n32053) );
  AND U32136 ( .A(n348), .B(n32346), .Z(n32345) );
  XNOR U32137 ( .A(n32347), .B(n32348), .Z(n348) );
  AND U32138 ( .A(n32349), .B(n32350), .Z(n32348) );
  XOR U32139 ( .A(n32347), .B(n32063), .Z(n32350) );
  XNOR U32140 ( .A(n32347), .B(n32013), .Z(n32349) );
  XOR U32141 ( .A(n32351), .B(n32352), .Z(n32347) );
  AND U32142 ( .A(n32353), .B(n32354), .Z(n32352) );
  XNOR U32143 ( .A(n32073), .B(n32351), .Z(n32354) );
  XOR U32144 ( .A(n32351), .B(n32023), .Z(n32353) );
  XOR U32145 ( .A(n32355), .B(n32356), .Z(n32351) );
  AND U32146 ( .A(n32357), .B(n32358), .Z(n32356) );
  XNOR U32147 ( .A(n32083), .B(n32355), .Z(n32358) );
  XOR U32148 ( .A(n32355), .B(n32032), .Z(n32357) );
  XOR U32149 ( .A(n32359), .B(n32360), .Z(n32355) );
  AND U32150 ( .A(n32361), .B(n32362), .Z(n32360) );
  XOR U32151 ( .A(n32359), .B(n32040), .Z(n32361) );
  XOR U32152 ( .A(n32363), .B(n32364), .Z(n32004) );
  AND U32153 ( .A(n352), .B(n32346), .Z(n32364) );
  XNOR U32154 ( .A(n32344), .B(n32363), .Z(n32346) );
  XNOR U32155 ( .A(n32365), .B(n32366), .Z(n352) );
  AND U32156 ( .A(n32367), .B(n32368), .Z(n32366) );
  XNOR U32157 ( .A(n32369), .B(n32365), .Z(n32368) );
  IV U32158 ( .A(n32063), .Z(n32369) );
  XOR U32159 ( .A(n32327), .B(n32370), .Z(n32063) );
  AND U32160 ( .A(n355), .B(n32371), .Z(n32370) );
  XOR U32161 ( .A(n32116), .B(n32113), .Z(n32371) );
  IV U32162 ( .A(n32327), .Z(n32116) );
  XNOR U32163 ( .A(n32013), .B(n32365), .Z(n32367) );
  XOR U32164 ( .A(n32372), .B(n32373), .Z(n32013) );
  AND U32165 ( .A(n371), .B(n32374), .Z(n32373) );
  XOR U32166 ( .A(n32375), .B(n32376), .Z(n32365) );
  AND U32167 ( .A(n32377), .B(n32378), .Z(n32376) );
  XNOR U32168 ( .A(n32375), .B(n32073), .Z(n32378) );
  XOR U32169 ( .A(n32133), .B(n32379), .Z(n32073) );
  AND U32170 ( .A(n355), .B(n32380), .Z(n32379) );
  XOR U32171 ( .A(n32129), .B(n32133), .Z(n32380) );
  XNOR U32172 ( .A(n32381), .B(n32375), .Z(n32377) );
  IV U32173 ( .A(n32023), .Z(n32381) );
  XOR U32174 ( .A(n32382), .B(n32383), .Z(n32023) );
  AND U32175 ( .A(n371), .B(n32384), .Z(n32383) );
  XOR U32176 ( .A(n32385), .B(n32386), .Z(n32375) );
  AND U32177 ( .A(n32387), .B(n32388), .Z(n32386) );
  XNOR U32178 ( .A(n32385), .B(n32083), .Z(n32388) );
  XOR U32179 ( .A(n32161), .B(n32389), .Z(n32083) );
  AND U32180 ( .A(n355), .B(n32390), .Z(n32389) );
  XOR U32181 ( .A(n32157), .B(n32161), .Z(n32390) );
  XOR U32182 ( .A(n32032), .B(n32385), .Z(n32387) );
  XOR U32183 ( .A(n32391), .B(n32392), .Z(n32032) );
  AND U32184 ( .A(n371), .B(n32393), .Z(n32392) );
  XOR U32185 ( .A(n32359), .B(n32394), .Z(n32385) );
  AND U32186 ( .A(n32395), .B(n32362), .Z(n32394) );
  XNOR U32187 ( .A(n32093), .B(n32359), .Z(n32362) );
  XOR U32188 ( .A(n32210), .B(n32396), .Z(n32093) );
  AND U32189 ( .A(n355), .B(n32397), .Z(n32396) );
  XOR U32190 ( .A(n32206), .B(n32210), .Z(n32397) );
  XNOR U32191 ( .A(n32398), .B(n32359), .Z(n32395) );
  IV U32192 ( .A(n32040), .Z(n32398) );
  XOR U32193 ( .A(n32399), .B(n32400), .Z(n32040) );
  AND U32194 ( .A(n371), .B(n32401), .Z(n32400) );
  XOR U32195 ( .A(n32402), .B(n32403), .Z(n32359) );
  AND U32196 ( .A(n32404), .B(n32405), .Z(n32403) );
  XNOR U32197 ( .A(n32402), .B(n32101), .Z(n32405) );
  XOR U32198 ( .A(n32303), .B(n32406), .Z(n32101) );
  AND U32199 ( .A(n355), .B(n32407), .Z(n32406) );
  XOR U32200 ( .A(n32299), .B(n32303), .Z(n32407) );
  XNOR U32201 ( .A(n32408), .B(n32402), .Z(n32404) );
  IV U32202 ( .A(n32050), .Z(n32408) );
  XOR U32203 ( .A(n32409), .B(n32410), .Z(n32050) );
  AND U32204 ( .A(n371), .B(n32411), .Z(n32410) );
  AND U32205 ( .A(n32363), .B(n32344), .Z(n32402) );
  XNOR U32206 ( .A(n32412), .B(n32413), .Z(n32344) );
  AND U32207 ( .A(n355), .B(n32322), .Z(n32413) );
  XNOR U32208 ( .A(n32320), .B(n32412), .Z(n32322) );
  XNOR U32209 ( .A(n32414), .B(n32415), .Z(n355) );
  AND U32210 ( .A(n32416), .B(n32417), .Z(n32415) );
  XNOR U32211 ( .A(n32414), .B(n32113), .Z(n32417) );
  IV U32212 ( .A(n32117), .Z(n32113) );
  XOR U32213 ( .A(n32418), .B(n32419), .Z(n32117) );
  AND U32214 ( .A(n359), .B(n32420), .Z(n32419) );
  XOR U32215 ( .A(n32421), .B(n32418), .Z(n32420) );
  XNOR U32216 ( .A(n32414), .B(n32327), .Z(n32416) );
  XOR U32217 ( .A(n32422), .B(n32423), .Z(n32327) );
  AND U32218 ( .A(n367), .B(n32374), .Z(n32423) );
  XOR U32219 ( .A(n32372), .B(n32422), .Z(n32374) );
  XOR U32220 ( .A(n32424), .B(n32425), .Z(n32414) );
  AND U32221 ( .A(n32426), .B(n32427), .Z(n32425) );
  XNOR U32222 ( .A(n32424), .B(n32129), .Z(n32427) );
  IV U32223 ( .A(n32132), .Z(n32129) );
  XOR U32224 ( .A(n32428), .B(n32429), .Z(n32132) );
  AND U32225 ( .A(n359), .B(n32430), .Z(n32429) );
  XOR U32226 ( .A(n32431), .B(n32428), .Z(n32430) );
  XOR U32227 ( .A(n32133), .B(n32424), .Z(n32426) );
  XOR U32228 ( .A(n32432), .B(n32433), .Z(n32133) );
  AND U32229 ( .A(n367), .B(n32384), .Z(n32433) );
  XOR U32230 ( .A(n32432), .B(n32382), .Z(n32384) );
  XOR U32231 ( .A(n32434), .B(n32435), .Z(n32424) );
  AND U32232 ( .A(n32436), .B(n32437), .Z(n32435) );
  XNOR U32233 ( .A(n32434), .B(n32157), .Z(n32437) );
  IV U32234 ( .A(n32160), .Z(n32157) );
  XOR U32235 ( .A(n32438), .B(n32439), .Z(n32160) );
  AND U32236 ( .A(n359), .B(n32440), .Z(n32439) );
  XNOR U32237 ( .A(n32441), .B(n32438), .Z(n32440) );
  XOR U32238 ( .A(n32161), .B(n32434), .Z(n32436) );
  XOR U32239 ( .A(n32442), .B(n32443), .Z(n32161) );
  AND U32240 ( .A(n367), .B(n32393), .Z(n32443) );
  XOR U32241 ( .A(n32442), .B(n32391), .Z(n32393) );
  XOR U32242 ( .A(n32444), .B(n32445), .Z(n32434) );
  AND U32243 ( .A(n32446), .B(n32447), .Z(n32445) );
  XNOR U32244 ( .A(n32444), .B(n32206), .Z(n32447) );
  IV U32245 ( .A(n32209), .Z(n32206) );
  XOR U32246 ( .A(n32448), .B(n32449), .Z(n32209) );
  AND U32247 ( .A(n359), .B(n32450), .Z(n32449) );
  XOR U32248 ( .A(n32451), .B(n32448), .Z(n32450) );
  XOR U32249 ( .A(n32210), .B(n32444), .Z(n32446) );
  XOR U32250 ( .A(n32452), .B(n32453), .Z(n32210) );
  AND U32251 ( .A(n367), .B(n32401), .Z(n32453) );
  XOR U32252 ( .A(n32452), .B(n32399), .Z(n32401) );
  XOR U32253 ( .A(n32340), .B(n32454), .Z(n32444) );
  AND U32254 ( .A(n32342), .B(n32455), .Z(n32454) );
  XNOR U32255 ( .A(n32340), .B(n32299), .Z(n32455) );
  IV U32256 ( .A(n32302), .Z(n32299) );
  XOR U32257 ( .A(n32456), .B(n32457), .Z(n32302) );
  AND U32258 ( .A(n359), .B(n32458), .Z(n32457) );
  XNOR U32259 ( .A(n32459), .B(n32456), .Z(n32458) );
  XOR U32260 ( .A(n32303), .B(n32340), .Z(n32342) );
  XOR U32261 ( .A(n32460), .B(n32461), .Z(n32303) );
  AND U32262 ( .A(n367), .B(n32411), .Z(n32461) );
  XOR U32263 ( .A(n32460), .B(n32409), .Z(n32411) );
  AND U32264 ( .A(n32412), .B(n32320), .Z(n32340) );
  XNOR U32265 ( .A(n32462), .B(n32463), .Z(n32320) );
  AND U32266 ( .A(n359), .B(n32464), .Z(n32463) );
  XNOR U32267 ( .A(n32465), .B(n32462), .Z(n32464) );
  XNOR U32268 ( .A(n32466), .B(n32467), .Z(n359) );
  AND U32269 ( .A(n32468), .B(n32469), .Z(n32467) );
  XOR U32270 ( .A(n32421), .B(n32466), .Z(n32469) );
  AND U32271 ( .A(n32470), .B(n32471), .Z(n32421) );
  XNOR U32272 ( .A(n32418), .B(n32466), .Z(n32468) );
  XNOR U32273 ( .A(n32472), .B(n32473), .Z(n32418) );
  AND U32274 ( .A(n363), .B(n32474), .Z(n32473) );
  XNOR U32275 ( .A(n32475), .B(n32476), .Z(n32474) );
  XOR U32276 ( .A(n32477), .B(n32478), .Z(n32466) );
  AND U32277 ( .A(n32479), .B(n32480), .Z(n32478) );
  XNOR U32278 ( .A(n32477), .B(n32470), .Z(n32480) );
  IV U32279 ( .A(n32431), .Z(n32470) );
  XOR U32280 ( .A(n32481), .B(n32482), .Z(n32431) );
  XOR U32281 ( .A(n32483), .B(n32471), .Z(n32482) );
  AND U32282 ( .A(n32441), .B(n32484), .Z(n32471) );
  AND U32283 ( .A(n32485), .B(n32486), .Z(n32483) );
  XOR U32284 ( .A(n32487), .B(n32481), .Z(n32485) );
  XNOR U32285 ( .A(n32428), .B(n32477), .Z(n32479) );
  XNOR U32286 ( .A(n32488), .B(n32489), .Z(n32428) );
  AND U32287 ( .A(n363), .B(n32490), .Z(n32489) );
  XNOR U32288 ( .A(n32491), .B(n32492), .Z(n32490) );
  XOR U32289 ( .A(n32493), .B(n32494), .Z(n32477) );
  AND U32290 ( .A(n32495), .B(n32496), .Z(n32494) );
  XNOR U32291 ( .A(n32493), .B(n32441), .Z(n32496) );
  XOR U32292 ( .A(n32497), .B(n32486), .Z(n32441) );
  XNOR U32293 ( .A(n32498), .B(n32481), .Z(n32486) );
  XOR U32294 ( .A(n32499), .B(n32500), .Z(n32481) );
  AND U32295 ( .A(n32501), .B(n32502), .Z(n32500) );
  XOR U32296 ( .A(n32503), .B(n32499), .Z(n32501) );
  XNOR U32297 ( .A(n32504), .B(n32505), .Z(n32498) );
  AND U32298 ( .A(n32506), .B(n32507), .Z(n32505) );
  XOR U32299 ( .A(n32504), .B(n32508), .Z(n32506) );
  XNOR U32300 ( .A(n32487), .B(n32484), .Z(n32497) );
  AND U32301 ( .A(n32509), .B(n32510), .Z(n32484) );
  XOR U32302 ( .A(n32511), .B(n32512), .Z(n32487) );
  AND U32303 ( .A(n32513), .B(n32514), .Z(n32512) );
  XOR U32304 ( .A(n32511), .B(n32515), .Z(n32513) );
  XNOR U32305 ( .A(n32438), .B(n32493), .Z(n32495) );
  XNOR U32306 ( .A(n32516), .B(n32517), .Z(n32438) );
  AND U32307 ( .A(n363), .B(n32518), .Z(n32517) );
  XNOR U32308 ( .A(n32519), .B(n32520), .Z(n32518) );
  XOR U32309 ( .A(n32521), .B(n32522), .Z(n32493) );
  AND U32310 ( .A(n32523), .B(n32524), .Z(n32522) );
  XNOR U32311 ( .A(n32521), .B(n32509), .Z(n32524) );
  IV U32312 ( .A(n32451), .Z(n32509) );
  XNOR U32313 ( .A(n32525), .B(n32502), .Z(n32451) );
  XNOR U32314 ( .A(n32526), .B(n32508), .Z(n32502) );
  XOR U32315 ( .A(n32527), .B(n32528), .Z(n32508) );
  AND U32316 ( .A(n32529), .B(n32530), .Z(n32528) );
  XOR U32317 ( .A(n32527), .B(n32531), .Z(n32529) );
  XNOR U32318 ( .A(n32507), .B(n32499), .Z(n32526) );
  XOR U32319 ( .A(n32532), .B(n32533), .Z(n32499) );
  AND U32320 ( .A(n32534), .B(n32535), .Z(n32533) );
  XNOR U32321 ( .A(n32536), .B(n32532), .Z(n32534) );
  XNOR U32322 ( .A(n32537), .B(n32504), .Z(n32507) );
  XOR U32323 ( .A(n32538), .B(n32539), .Z(n32504) );
  AND U32324 ( .A(n32540), .B(n32541), .Z(n32539) );
  XOR U32325 ( .A(n32538), .B(n32542), .Z(n32540) );
  XNOR U32326 ( .A(n32543), .B(n32544), .Z(n32537) );
  AND U32327 ( .A(n32545), .B(n32546), .Z(n32544) );
  XNOR U32328 ( .A(n32543), .B(n32547), .Z(n32545) );
  XNOR U32329 ( .A(n32503), .B(n32510), .Z(n32525) );
  AND U32330 ( .A(n32459), .B(n32548), .Z(n32510) );
  XOR U32331 ( .A(n32515), .B(n32514), .Z(n32503) );
  XNOR U32332 ( .A(n32549), .B(n32511), .Z(n32514) );
  XOR U32333 ( .A(n32550), .B(n32551), .Z(n32511) );
  AND U32334 ( .A(n32552), .B(n32553), .Z(n32551) );
  XOR U32335 ( .A(n32550), .B(n32554), .Z(n32552) );
  XNOR U32336 ( .A(n32555), .B(n32556), .Z(n32549) );
  AND U32337 ( .A(n32557), .B(n32558), .Z(n32556) );
  XOR U32338 ( .A(n32555), .B(n32559), .Z(n32557) );
  XOR U32339 ( .A(n32560), .B(n32561), .Z(n32515) );
  AND U32340 ( .A(n32562), .B(n32563), .Z(n32561) );
  XOR U32341 ( .A(n32560), .B(n32564), .Z(n32562) );
  XNOR U32342 ( .A(n32448), .B(n32521), .Z(n32523) );
  XNOR U32343 ( .A(n32565), .B(n32566), .Z(n32448) );
  AND U32344 ( .A(n363), .B(n32567), .Z(n32566) );
  XNOR U32345 ( .A(n32568), .B(n32569), .Z(n32567) );
  XOR U32346 ( .A(n32570), .B(n32571), .Z(n32521) );
  AND U32347 ( .A(n32572), .B(n32573), .Z(n32571) );
  XNOR U32348 ( .A(n32570), .B(n32459), .Z(n32573) );
  XOR U32349 ( .A(n32574), .B(n32535), .Z(n32459) );
  XNOR U32350 ( .A(n32575), .B(n32542), .Z(n32535) );
  XOR U32351 ( .A(n32531), .B(n32530), .Z(n32542) );
  XNOR U32352 ( .A(n32576), .B(n32527), .Z(n32530) );
  XOR U32353 ( .A(n32577), .B(n32578), .Z(n32527) );
  AND U32354 ( .A(n32579), .B(n32580), .Z(n32578) );
  XOR U32355 ( .A(n32577), .B(n32581), .Z(n32579) );
  XNOR U32356 ( .A(n32582), .B(n32583), .Z(n32576) );
  NOR U32357 ( .A(n32584), .B(n32585), .Z(n32583) );
  XNOR U32358 ( .A(n32582), .B(n32586), .Z(n32584) );
  XOR U32359 ( .A(n32587), .B(n32588), .Z(n32531) );
  NOR U32360 ( .A(n32589), .B(n32590), .Z(n32588) );
  XNOR U32361 ( .A(n32587), .B(n32591), .Z(n32589) );
  XNOR U32362 ( .A(n32541), .B(n32532), .Z(n32575) );
  XOR U32363 ( .A(n32592), .B(n32593), .Z(n32532) );
  NOR U32364 ( .A(n32594), .B(n32595), .Z(n32593) );
  XNOR U32365 ( .A(n32592), .B(n32596), .Z(n32594) );
  XOR U32366 ( .A(n32597), .B(n32547), .Z(n32541) );
  XNOR U32367 ( .A(n32598), .B(n32599), .Z(n32547) );
  NOR U32368 ( .A(n32600), .B(n32601), .Z(n32599) );
  XNOR U32369 ( .A(n32598), .B(n32602), .Z(n32600) );
  XNOR U32370 ( .A(n32546), .B(n32538), .Z(n32597) );
  XOR U32371 ( .A(n32603), .B(n32604), .Z(n32538) );
  AND U32372 ( .A(n32605), .B(n32606), .Z(n32604) );
  XOR U32373 ( .A(n32603), .B(n32607), .Z(n32605) );
  XNOR U32374 ( .A(n32608), .B(n32543), .Z(n32546) );
  XOR U32375 ( .A(n32609), .B(n32610), .Z(n32543) );
  AND U32376 ( .A(n32611), .B(n32612), .Z(n32610) );
  XOR U32377 ( .A(n32609), .B(n32613), .Z(n32611) );
  XNOR U32378 ( .A(n32614), .B(n32615), .Z(n32608) );
  NOR U32379 ( .A(n32616), .B(n32617), .Z(n32615) );
  XOR U32380 ( .A(n32614), .B(n32618), .Z(n32616) );
  XOR U32381 ( .A(n32536), .B(n32548), .Z(n32574) );
  NOR U32382 ( .A(n32465), .B(n32619), .Z(n32548) );
  XNOR U32383 ( .A(n32554), .B(n32553), .Z(n32536) );
  XNOR U32384 ( .A(n32620), .B(n32559), .Z(n32553) );
  XOR U32385 ( .A(n32621), .B(n32622), .Z(n32559) );
  NOR U32386 ( .A(n32623), .B(n32624), .Z(n32622) );
  XNOR U32387 ( .A(n32621), .B(n32625), .Z(n32623) );
  XNOR U32388 ( .A(n32558), .B(n32550), .Z(n32620) );
  XOR U32389 ( .A(n32626), .B(n32627), .Z(n32550) );
  AND U32390 ( .A(n32628), .B(n32629), .Z(n32627) );
  XNOR U32391 ( .A(n32626), .B(n32630), .Z(n32628) );
  XNOR U32392 ( .A(n32631), .B(n32555), .Z(n32558) );
  XOR U32393 ( .A(n32632), .B(n32633), .Z(n32555) );
  AND U32394 ( .A(n32634), .B(n32635), .Z(n32633) );
  XOR U32395 ( .A(n32632), .B(n32636), .Z(n32634) );
  XNOR U32396 ( .A(n32637), .B(n32638), .Z(n32631) );
  NOR U32397 ( .A(n32639), .B(n32640), .Z(n32638) );
  XOR U32398 ( .A(n32637), .B(n32641), .Z(n32639) );
  XOR U32399 ( .A(n32564), .B(n32563), .Z(n32554) );
  XNOR U32400 ( .A(n32642), .B(n32560), .Z(n32563) );
  XOR U32401 ( .A(n32643), .B(n32644), .Z(n32560) );
  AND U32402 ( .A(n32645), .B(n32646), .Z(n32644) );
  XOR U32403 ( .A(n32643), .B(n32647), .Z(n32645) );
  XNOR U32404 ( .A(n32648), .B(n32649), .Z(n32642) );
  NOR U32405 ( .A(n32650), .B(n32651), .Z(n32649) );
  XNOR U32406 ( .A(n32648), .B(n32652), .Z(n32650) );
  XOR U32407 ( .A(n32653), .B(n32654), .Z(n32564) );
  NOR U32408 ( .A(n32655), .B(n32656), .Z(n32654) );
  XNOR U32409 ( .A(n32653), .B(n32657), .Z(n32655) );
  XNOR U32410 ( .A(n32456), .B(n32570), .Z(n32572) );
  XNOR U32411 ( .A(n32658), .B(n32659), .Z(n32456) );
  AND U32412 ( .A(n363), .B(n32660), .Z(n32659) );
  XNOR U32413 ( .A(n32661), .B(n32662), .Z(n32660) );
  AND U32414 ( .A(n32462), .B(n32465), .Z(n32570) );
  XOR U32415 ( .A(n32663), .B(n32619), .Z(n32465) );
  XNOR U32416 ( .A(p_input[2048]), .B(p_input[384]), .Z(n32619) );
  XOR U32417 ( .A(n32596), .B(n32595), .Z(n32663) );
  XOR U32418 ( .A(n32664), .B(n32607), .Z(n32595) );
  XOR U32419 ( .A(n32581), .B(n32580), .Z(n32607) );
  XNOR U32420 ( .A(n32665), .B(n32586), .Z(n32580) );
  XOR U32421 ( .A(p_input[2072]), .B(p_input[408]), .Z(n32586) );
  XOR U32422 ( .A(n32577), .B(n32585), .Z(n32665) );
  XOR U32423 ( .A(n32666), .B(n32582), .Z(n32585) );
  XOR U32424 ( .A(p_input[2070]), .B(p_input[406]), .Z(n32582) );
  XNOR U32425 ( .A(p_input[2071]), .B(p_input[407]), .Z(n32666) );
  XNOR U32426 ( .A(n28684), .B(p_input[402]), .Z(n32577) );
  XNOR U32427 ( .A(n32591), .B(n32590), .Z(n32581) );
  XOR U32428 ( .A(n32667), .B(n32587), .Z(n32590) );
  XOR U32429 ( .A(p_input[2067]), .B(p_input[403]), .Z(n32587) );
  XNOR U32430 ( .A(p_input[2068]), .B(p_input[404]), .Z(n32667) );
  XOR U32431 ( .A(p_input[2069]), .B(p_input[405]), .Z(n32591) );
  XNOR U32432 ( .A(n32606), .B(n32592), .Z(n32664) );
  XNOR U32433 ( .A(n28686), .B(p_input[385]), .Z(n32592) );
  XNOR U32434 ( .A(n32668), .B(n32613), .Z(n32606) );
  XNOR U32435 ( .A(n32602), .B(n32601), .Z(n32613) );
  XOR U32436 ( .A(n32669), .B(n32598), .Z(n32601) );
  XNOR U32437 ( .A(n28322), .B(p_input[410]), .Z(n32598) );
  XNOR U32438 ( .A(p_input[2075]), .B(p_input[411]), .Z(n32669) );
  XOR U32439 ( .A(p_input[2076]), .B(p_input[412]), .Z(n32602) );
  XNOR U32440 ( .A(n32612), .B(n32603), .Z(n32668) );
  XNOR U32441 ( .A(n28689), .B(p_input[401]), .Z(n32603) );
  XOR U32442 ( .A(n32670), .B(n32618), .Z(n32612) );
  XNOR U32443 ( .A(p_input[2079]), .B(p_input[415]), .Z(n32618) );
  XOR U32444 ( .A(n32609), .B(n32617), .Z(n32670) );
  XOR U32445 ( .A(n32671), .B(n32614), .Z(n32617) );
  XOR U32446 ( .A(p_input[2077]), .B(p_input[413]), .Z(n32614) );
  XNOR U32447 ( .A(p_input[2078]), .B(p_input[414]), .Z(n32671) );
  XNOR U32448 ( .A(n28326), .B(p_input[409]), .Z(n32609) );
  XNOR U32449 ( .A(n32630), .B(n32629), .Z(n32596) );
  XNOR U32450 ( .A(n32672), .B(n32636), .Z(n32629) );
  XNOR U32451 ( .A(n32625), .B(n32624), .Z(n32636) );
  XOR U32452 ( .A(n32673), .B(n32621), .Z(n32624) );
  XNOR U32453 ( .A(n28694), .B(p_input[395]), .Z(n32621) );
  XNOR U32454 ( .A(p_input[2060]), .B(p_input[396]), .Z(n32673) );
  XOR U32455 ( .A(p_input[2061]), .B(p_input[397]), .Z(n32625) );
  XNOR U32456 ( .A(n32635), .B(n32626), .Z(n32672) );
  XNOR U32457 ( .A(n28330), .B(p_input[386]), .Z(n32626) );
  XOR U32458 ( .A(n32674), .B(n32641), .Z(n32635) );
  XNOR U32459 ( .A(p_input[2064]), .B(p_input[400]), .Z(n32641) );
  XOR U32460 ( .A(n32632), .B(n32640), .Z(n32674) );
  XOR U32461 ( .A(n32675), .B(n32637), .Z(n32640) );
  XOR U32462 ( .A(p_input[2062]), .B(p_input[398]), .Z(n32637) );
  XNOR U32463 ( .A(p_input[2063]), .B(p_input[399]), .Z(n32675) );
  XNOR U32464 ( .A(n28697), .B(p_input[394]), .Z(n32632) );
  XNOR U32465 ( .A(n32647), .B(n32646), .Z(n32630) );
  XNOR U32466 ( .A(n32676), .B(n32652), .Z(n32646) );
  XOR U32467 ( .A(p_input[2057]), .B(p_input[393]), .Z(n32652) );
  XOR U32468 ( .A(n32643), .B(n32651), .Z(n32676) );
  XOR U32469 ( .A(n32677), .B(n32648), .Z(n32651) );
  XOR U32470 ( .A(p_input[2055]), .B(p_input[391]), .Z(n32648) );
  XNOR U32471 ( .A(p_input[2056]), .B(p_input[392]), .Z(n32677) );
  XNOR U32472 ( .A(n28337), .B(p_input[387]), .Z(n32643) );
  XNOR U32473 ( .A(n32657), .B(n32656), .Z(n32647) );
  XOR U32474 ( .A(n32678), .B(n32653), .Z(n32656) );
  XOR U32475 ( .A(p_input[2052]), .B(p_input[388]), .Z(n32653) );
  XNOR U32476 ( .A(p_input[2053]), .B(p_input[389]), .Z(n32678) );
  XOR U32477 ( .A(p_input[2054]), .B(p_input[390]), .Z(n32657) );
  XNOR U32478 ( .A(n32679), .B(n32680), .Z(n32462) );
  AND U32479 ( .A(n363), .B(n32681), .Z(n32680) );
  XNOR U32480 ( .A(n32682), .B(n32683), .Z(n363) );
  AND U32481 ( .A(n32684), .B(n32685), .Z(n32683) );
  XOR U32482 ( .A(n32476), .B(n32682), .Z(n32685) );
  XNOR U32483 ( .A(n32686), .B(n32682), .Z(n32684) );
  XOR U32484 ( .A(n32687), .B(n32688), .Z(n32682) );
  AND U32485 ( .A(n32689), .B(n32690), .Z(n32688) );
  XOR U32486 ( .A(n32491), .B(n32687), .Z(n32690) );
  XOR U32487 ( .A(n32687), .B(n32492), .Z(n32689) );
  XOR U32488 ( .A(n32691), .B(n32692), .Z(n32687) );
  AND U32489 ( .A(n32693), .B(n32694), .Z(n32692) );
  XOR U32490 ( .A(n32519), .B(n32691), .Z(n32694) );
  XOR U32491 ( .A(n32691), .B(n32520), .Z(n32693) );
  XOR U32492 ( .A(n32695), .B(n32696), .Z(n32691) );
  AND U32493 ( .A(n32697), .B(n32698), .Z(n32696) );
  XOR U32494 ( .A(n32568), .B(n32695), .Z(n32698) );
  XOR U32495 ( .A(n32695), .B(n32569), .Z(n32697) );
  XOR U32496 ( .A(n32699), .B(n32700), .Z(n32695) );
  AND U32497 ( .A(n32701), .B(n32702), .Z(n32700) );
  XOR U32498 ( .A(n32699), .B(n32661), .Z(n32702) );
  XNOR U32499 ( .A(n32703), .B(n32704), .Z(n32412) );
  AND U32500 ( .A(n367), .B(n32705), .Z(n32704) );
  XNOR U32501 ( .A(n32706), .B(n32707), .Z(n367) );
  AND U32502 ( .A(n32708), .B(n32709), .Z(n32707) );
  XOR U32503 ( .A(n32706), .B(n32422), .Z(n32709) );
  XNOR U32504 ( .A(n32706), .B(n32372), .Z(n32708) );
  XOR U32505 ( .A(n32710), .B(n32711), .Z(n32706) );
  AND U32506 ( .A(n32712), .B(n32713), .Z(n32711) );
  XNOR U32507 ( .A(n32432), .B(n32710), .Z(n32713) );
  XOR U32508 ( .A(n32710), .B(n32382), .Z(n32712) );
  XOR U32509 ( .A(n32714), .B(n32715), .Z(n32710) );
  AND U32510 ( .A(n32716), .B(n32717), .Z(n32715) );
  XNOR U32511 ( .A(n32442), .B(n32714), .Z(n32717) );
  XOR U32512 ( .A(n32714), .B(n32391), .Z(n32716) );
  XOR U32513 ( .A(n32718), .B(n32719), .Z(n32714) );
  AND U32514 ( .A(n32720), .B(n32721), .Z(n32719) );
  XOR U32515 ( .A(n32718), .B(n32399), .Z(n32720) );
  XOR U32516 ( .A(n32722), .B(n32723), .Z(n32363) );
  AND U32517 ( .A(n371), .B(n32705), .Z(n32723) );
  XNOR U32518 ( .A(n32703), .B(n32722), .Z(n32705) );
  XNOR U32519 ( .A(n32724), .B(n32725), .Z(n371) );
  AND U32520 ( .A(n32726), .B(n32727), .Z(n32725) );
  XNOR U32521 ( .A(n32728), .B(n32724), .Z(n32727) );
  IV U32522 ( .A(n32422), .Z(n32728) );
  XOR U32523 ( .A(n32686), .B(n32729), .Z(n32422) );
  AND U32524 ( .A(n374), .B(n32730), .Z(n32729) );
  XOR U32525 ( .A(n32475), .B(n32472), .Z(n32730) );
  IV U32526 ( .A(n32686), .Z(n32475) );
  XNOR U32527 ( .A(n32372), .B(n32724), .Z(n32726) );
  XOR U32528 ( .A(n32731), .B(n32732), .Z(n32372) );
  AND U32529 ( .A(n390), .B(n32733), .Z(n32732) );
  XOR U32530 ( .A(n32734), .B(n32735), .Z(n32724) );
  AND U32531 ( .A(n32736), .B(n32737), .Z(n32735) );
  XNOR U32532 ( .A(n32734), .B(n32432), .Z(n32737) );
  XOR U32533 ( .A(n32492), .B(n32738), .Z(n32432) );
  AND U32534 ( .A(n374), .B(n32739), .Z(n32738) );
  XOR U32535 ( .A(n32488), .B(n32492), .Z(n32739) );
  XNOR U32536 ( .A(n32740), .B(n32734), .Z(n32736) );
  IV U32537 ( .A(n32382), .Z(n32740) );
  XOR U32538 ( .A(n32741), .B(n32742), .Z(n32382) );
  AND U32539 ( .A(n390), .B(n32743), .Z(n32742) );
  XOR U32540 ( .A(n32744), .B(n32745), .Z(n32734) );
  AND U32541 ( .A(n32746), .B(n32747), .Z(n32745) );
  XNOR U32542 ( .A(n32744), .B(n32442), .Z(n32747) );
  XOR U32543 ( .A(n32520), .B(n32748), .Z(n32442) );
  AND U32544 ( .A(n374), .B(n32749), .Z(n32748) );
  XOR U32545 ( .A(n32516), .B(n32520), .Z(n32749) );
  XOR U32546 ( .A(n32391), .B(n32744), .Z(n32746) );
  XOR U32547 ( .A(n32750), .B(n32751), .Z(n32391) );
  AND U32548 ( .A(n390), .B(n32752), .Z(n32751) );
  XOR U32549 ( .A(n32718), .B(n32753), .Z(n32744) );
  AND U32550 ( .A(n32754), .B(n32721), .Z(n32753) );
  XNOR U32551 ( .A(n32452), .B(n32718), .Z(n32721) );
  XOR U32552 ( .A(n32569), .B(n32755), .Z(n32452) );
  AND U32553 ( .A(n374), .B(n32756), .Z(n32755) );
  XOR U32554 ( .A(n32565), .B(n32569), .Z(n32756) );
  XNOR U32555 ( .A(n32757), .B(n32718), .Z(n32754) );
  IV U32556 ( .A(n32399), .Z(n32757) );
  XOR U32557 ( .A(n32758), .B(n32759), .Z(n32399) );
  AND U32558 ( .A(n390), .B(n32760), .Z(n32759) );
  XOR U32559 ( .A(n32761), .B(n32762), .Z(n32718) );
  AND U32560 ( .A(n32763), .B(n32764), .Z(n32762) );
  XNOR U32561 ( .A(n32761), .B(n32460), .Z(n32764) );
  XOR U32562 ( .A(n32662), .B(n32765), .Z(n32460) );
  AND U32563 ( .A(n374), .B(n32766), .Z(n32765) );
  XOR U32564 ( .A(n32658), .B(n32662), .Z(n32766) );
  XNOR U32565 ( .A(n32767), .B(n32761), .Z(n32763) );
  IV U32566 ( .A(n32409), .Z(n32767) );
  XOR U32567 ( .A(n32768), .B(n32769), .Z(n32409) );
  AND U32568 ( .A(n390), .B(n32770), .Z(n32769) );
  AND U32569 ( .A(n32722), .B(n32703), .Z(n32761) );
  XNOR U32570 ( .A(n32771), .B(n32772), .Z(n32703) );
  AND U32571 ( .A(n374), .B(n32681), .Z(n32772) );
  XNOR U32572 ( .A(n32679), .B(n32771), .Z(n32681) );
  XNOR U32573 ( .A(n32773), .B(n32774), .Z(n374) );
  AND U32574 ( .A(n32775), .B(n32776), .Z(n32774) );
  XNOR U32575 ( .A(n32773), .B(n32472), .Z(n32776) );
  IV U32576 ( .A(n32476), .Z(n32472) );
  XOR U32577 ( .A(n32777), .B(n32778), .Z(n32476) );
  AND U32578 ( .A(n378), .B(n32779), .Z(n32778) );
  XOR U32579 ( .A(n32780), .B(n32777), .Z(n32779) );
  XNOR U32580 ( .A(n32773), .B(n32686), .Z(n32775) );
  XOR U32581 ( .A(n32781), .B(n32782), .Z(n32686) );
  AND U32582 ( .A(n386), .B(n32733), .Z(n32782) );
  XOR U32583 ( .A(n32731), .B(n32781), .Z(n32733) );
  XOR U32584 ( .A(n32783), .B(n32784), .Z(n32773) );
  AND U32585 ( .A(n32785), .B(n32786), .Z(n32784) );
  XNOR U32586 ( .A(n32783), .B(n32488), .Z(n32786) );
  IV U32587 ( .A(n32491), .Z(n32488) );
  XOR U32588 ( .A(n32787), .B(n32788), .Z(n32491) );
  AND U32589 ( .A(n378), .B(n32789), .Z(n32788) );
  XOR U32590 ( .A(n32790), .B(n32787), .Z(n32789) );
  XOR U32591 ( .A(n32492), .B(n32783), .Z(n32785) );
  XOR U32592 ( .A(n32791), .B(n32792), .Z(n32492) );
  AND U32593 ( .A(n386), .B(n32743), .Z(n32792) );
  XOR U32594 ( .A(n32791), .B(n32741), .Z(n32743) );
  XOR U32595 ( .A(n32793), .B(n32794), .Z(n32783) );
  AND U32596 ( .A(n32795), .B(n32796), .Z(n32794) );
  XNOR U32597 ( .A(n32793), .B(n32516), .Z(n32796) );
  IV U32598 ( .A(n32519), .Z(n32516) );
  XOR U32599 ( .A(n32797), .B(n32798), .Z(n32519) );
  AND U32600 ( .A(n378), .B(n32799), .Z(n32798) );
  XNOR U32601 ( .A(n32800), .B(n32797), .Z(n32799) );
  XOR U32602 ( .A(n32520), .B(n32793), .Z(n32795) );
  XOR U32603 ( .A(n32801), .B(n32802), .Z(n32520) );
  AND U32604 ( .A(n386), .B(n32752), .Z(n32802) );
  XOR U32605 ( .A(n32801), .B(n32750), .Z(n32752) );
  XOR U32606 ( .A(n32803), .B(n32804), .Z(n32793) );
  AND U32607 ( .A(n32805), .B(n32806), .Z(n32804) );
  XNOR U32608 ( .A(n32803), .B(n32565), .Z(n32806) );
  IV U32609 ( .A(n32568), .Z(n32565) );
  XOR U32610 ( .A(n32807), .B(n32808), .Z(n32568) );
  AND U32611 ( .A(n378), .B(n32809), .Z(n32808) );
  XOR U32612 ( .A(n32810), .B(n32807), .Z(n32809) );
  XOR U32613 ( .A(n32569), .B(n32803), .Z(n32805) );
  XOR U32614 ( .A(n32811), .B(n32812), .Z(n32569) );
  AND U32615 ( .A(n386), .B(n32760), .Z(n32812) );
  XOR U32616 ( .A(n32811), .B(n32758), .Z(n32760) );
  XOR U32617 ( .A(n32699), .B(n32813), .Z(n32803) );
  AND U32618 ( .A(n32701), .B(n32814), .Z(n32813) );
  XNOR U32619 ( .A(n32699), .B(n32658), .Z(n32814) );
  IV U32620 ( .A(n32661), .Z(n32658) );
  XOR U32621 ( .A(n32815), .B(n32816), .Z(n32661) );
  AND U32622 ( .A(n378), .B(n32817), .Z(n32816) );
  XNOR U32623 ( .A(n32818), .B(n32815), .Z(n32817) );
  XOR U32624 ( .A(n32662), .B(n32699), .Z(n32701) );
  XOR U32625 ( .A(n32819), .B(n32820), .Z(n32662) );
  AND U32626 ( .A(n386), .B(n32770), .Z(n32820) );
  XOR U32627 ( .A(n32819), .B(n32768), .Z(n32770) );
  AND U32628 ( .A(n32771), .B(n32679), .Z(n32699) );
  XNOR U32629 ( .A(n32821), .B(n32822), .Z(n32679) );
  AND U32630 ( .A(n378), .B(n32823), .Z(n32822) );
  XNOR U32631 ( .A(n32824), .B(n32821), .Z(n32823) );
  XNOR U32632 ( .A(n32825), .B(n32826), .Z(n378) );
  AND U32633 ( .A(n32827), .B(n32828), .Z(n32826) );
  XOR U32634 ( .A(n32780), .B(n32825), .Z(n32828) );
  AND U32635 ( .A(n32829), .B(n32830), .Z(n32780) );
  XNOR U32636 ( .A(n32777), .B(n32825), .Z(n32827) );
  XNOR U32637 ( .A(n32831), .B(n32832), .Z(n32777) );
  AND U32638 ( .A(n382), .B(n32833), .Z(n32832) );
  XNOR U32639 ( .A(n32834), .B(n32835), .Z(n32833) );
  XOR U32640 ( .A(n32836), .B(n32837), .Z(n32825) );
  AND U32641 ( .A(n32838), .B(n32839), .Z(n32837) );
  XNOR U32642 ( .A(n32836), .B(n32829), .Z(n32839) );
  IV U32643 ( .A(n32790), .Z(n32829) );
  XOR U32644 ( .A(n32840), .B(n32841), .Z(n32790) );
  XOR U32645 ( .A(n32842), .B(n32830), .Z(n32841) );
  AND U32646 ( .A(n32800), .B(n32843), .Z(n32830) );
  AND U32647 ( .A(n32844), .B(n32845), .Z(n32842) );
  XOR U32648 ( .A(n32846), .B(n32840), .Z(n32844) );
  XNOR U32649 ( .A(n32787), .B(n32836), .Z(n32838) );
  XNOR U32650 ( .A(n32847), .B(n32848), .Z(n32787) );
  AND U32651 ( .A(n382), .B(n32849), .Z(n32848) );
  XNOR U32652 ( .A(n32850), .B(n32851), .Z(n32849) );
  XOR U32653 ( .A(n32852), .B(n32853), .Z(n32836) );
  AND U32654 ( .A(n32854), .B(n32855), .Z(n32853) );
  XNOR U32655 ( .A(n32852), .B(n32800), .Z(n32855) );
  XOR U32656 ( .A(n32856), .B(n32845), .Z(n32800) );
  XNOR U32657 ( .A(n32857), .B(n32840), .Z(n32845) );
  XOR U32658 ( .A(n32858), .B(n32859), .Z(n32840) );
  AND U32659 ( .A(n32860), .B(n32861), .Z(n32859) );
  XOR U32660 ( .A(n32862), .B(n32858), .Z(n32860) );
  XNOR U32661 ( .A(n32863), .B(n32864), .Z(n32857) );
  AND U32662 ( .A(n32865), .B(n32866), .Z(n32864) );
  XOR U32663 ( .A(n32863), .B(n32867), .Z(n32865) );
  XNOR U32664 ( .A(n32846), .B(n32843), .Z(n32856) );
  AND U32665 ( .A(n32868), .B(n32869), .Z(n32843) );
  XOR U32666 ( .A(n32870), .B(n32871), .Z(n32846) );
  AND U32667 ( .A(n32872), .B(n32873), .Z(n32871) );
  XOR U32668 ( .A(n32870), .B(n32874), .Z(n32872) );
  XNOR U32669 ( .A(n32797), .B(n32852), .Z(n32854) );
  XNOR U32670 ( .A(n32875), .B(n32876), .Z(n32797) );
  AND U32671 ( .A(n382), .B(n32877), .Z(n32876) );
  XNOR U32672 ( .A(n32878), .B(n32879), .Z(n32877) );
  XOR U32673 ( .A(n32880), .B(n32881), .Z(n32852) );
  AND U32674 ( .A(n32882), .B(n32883), .Z(n32881) );
  XNOR U32675 ( .A(n32880), .B(n32868), .Z(n32883) );
  IV U32676 ( .A(n32810), .Z(n32868) );
  XNOR U32677 ( .A(n32884), .B(n32861), .Z(n32810) );
  XNOR U32678 ( .A(n32885), .B(n32867), .Z(n32861) );
  XOR U32679 ( .A(n32886), .B(n32887), .Z(n32867) );
  AND U32680 ( .A(n32888), .B(n32889), .Z(n32887) );
  XOR U32681 ( .A(n32886), .B(n32890), .Z(n32888) );
  XNOR U32682 ( .A(n32866), .B(n32858), .Z(n32885) );
  XOR U32683 ( .A(n32891), .B(n32892), .Z(n32858) );
  AND U32684 ( .A(n32893), .B(n32894), .Z(n32892) );
  XNOR U32685 ( .A(n32895), .B(n32891), .Z(n32893) );
  XNOR U32686 ( .A(n32896), .B(n32863), .Z(n32866) );
  XOR U32687 ( .A(n32897), .B(n32898), .Z(n32863) );
  AND U32688 ( .A(n32899), .B(n32900), .Z(n32898) );
  XOR U32689 ( .A(n32897), .B(n32901), .Z(n32899) );
  XNOR U32690 ( .A(n32902), .B(n32903), .Z(n32896) );
  AND U32691 ( .A(n32904), .B(n32905), .Z(n32903) );
  XNOR U32692 ( .A(n32902), .B(n32906), .Z(n32904) );
  XNOR U32693 ( .A(n32862), .B(n32869), .Z(n32884) );
  AND U32694 ( .A(n32818), .B(n32907), .Z(n32869) );
  XOR U32695 ( .A(n32874), .B(n32873), .Z(n32862) );
  XNOR U32696 ( .A(n32908), .B(n32870), .Z(n32873) );
  XOR U32697 ( .A(n32909), .B(n32910), .Z(n32870) );
  AND U32698 ( .A(n32911), .B(n32912), .Z(n32910) );
  XOR U32699 ( .A(n32909), .B(n32913), .Z(n32911) );
  XNOR U32700 ( .A(n32914), .B(n32915), .Z(n32908) );
  AND U32701 ( .A(n32916), .B(n32917), .Z(n32915) );
  XOR U32702 ( .A(n32914), .B(n32918), .Z(n32916) );
  XOR U32703 ( .A(n32919), .B(n32920), .Z(n32874) );
  AND U32704 ( .A(n32921), .B(n32922), .Z(n32920) );
  XOR U32705 ( .A(n32919), .B(n32923), .Z(n32921) );
  XNOR U32706 ( .A(n32807), .B(n32880), .Z(n32882) );
  XNOR U32707 ( .A(n32924), .B(n32925), .Z(n32807) );
  AND U32708 ( .A(n382), .B(n32926), .Z(n32925) );
  XNOR U32709 ( .A(n32927), .B(n32928), .Z(n32926) );
  XOR U32710 ( .A(n32929), .B(n32930), .Z(n32880) );
  AND U32711 ( .A(n32931), .B(n32932), .Z(n32930) );
  XNOR U32712 ( .A(n32929), .B(n32818), .Z(n32932) );
  XOR U32713 ( .A(n32933), .B(n32894), .Z(n32818) );
  XNOR U32714 ( .A(n32934), .B(n32901), .Z(n32894) );
  XOR U32715 ( .A(n32890), .B(n32889), .Z(n32901) );
  XNOR U32716 ( .A(n32935), .B(n32886), .Z(n32889) );
  XOR U32717 ( .A(n32936), .B(n32937), .Z(n32886) );
  AND U32718 ( .A(n32938), .B(n32939), .Z(n32937) );
  XOR U32719 ( .A(n32936), .B(n32940), .Z(n32938) );
  XNOR U32720 ( .A(n32941), .B(n32942), .Z(n32935) );
  NOR U32721 ( .A(n32943), .B(n32944), .Z(n32942) );
  XNOR U32722 ( .A(n32941), .B(n32945), .Z(n32943) );
  XOR U32723 ( .A(n32946), .B(n32947), .Z(n32890) );
  NOR U32724 ( .A(n32948), .B(n32949), .Z(n32947) );
  XNOR U32725 ( .A(n32946), .B(n32950), .Z(n32948) );
  XNOR U32726 ( .A(n32900), .B(n32891), .Z(n32934) );
  XOR U32727 ( .A(n32951), .B(n32952), .Z(n32891) );
  NOR U32728 ( .A(n32953), .B(n32954), .Z(n32952) );
  XNOR U32729 ( .A(n32951), .B(n32955), .Z(n32953) );
  XOR U32730 ( .A(n32956), .B(n32906), .Z(n32900) );
  XNOR U32731 ( .A(n32957), .B(n32958), .Z(n32906) );
  NOR U32732 ( .A(n32959), .B(n32960), .Z(n32958) );
  XNOR U32733 ( .A(n32957), .B(n32961), .Z(n32959) );
  XNOR U32734 ( .A(n32905), .B(n32897), .Z(n32956) );
  XOR U32735 ( .A(n32962), .B(n32963), .Z(n32897) );
  AND U32736 ( .A(n32964), .B(n32965), .Z(n32963) );
  XOR U32737 ( .A(n32962), .B(n32966), .Z(n32964) );
  XNOR U32738 ( .A(n32967), .B(n32902), .Z(n32905) );
  XOR U32739 ( .A(n32968), .B(n32969), .Z(n32902) );
  AND U32740 ( .A(n32970), .B(n32971), .Z(n32969) );
  XOR U32741 ( .A(n32968), .B(n32972), .Z(n32970) );
  XNOR U32742 ( .A(n32973), .B(n32974), .Z(n32967) );
  NOR U32743 ( .A(n32975), .B(n32976), .Z(n32974) );
  XOR U32744 ( .A(n32973), .B(n32977), .Z(n32975) );
  XOR U32745 ( .A(n32895), .B(n32907), .Z(n32933) );
  NOR U32746 ( .A(n32824), .B(n32978), .Z(n32907) );
  XNOR U32747 ( .A(n32913), .B(n32912), .Z(n32895) );
  XNOR U32748 ( .A(n32979), .B(n32918), .Z(n32912) );
  XOR U32749 ( .A(n32980), .B(n32981), .Z(n32918) );
  NOR U32750 ( .A(n32982), .B(n32983), .Z(n32981) );
  XNOR U32751 ( .A(n32980), .B(n32984), .Z(n32982) );
  XNOR U32752 ( .A(n32917), .B(n32909), .Z(n32979) );
  XOR U32753 ( .A(n32985), .B(n32986), .Z(n32909) );
  AND U32754 ( .A(n32987), .B(n32988), .Z(n32986) );
  XNOR U32755 ( .A(n32985), .B(n32989), .Z(n32987) );
  XNOR U32756 ( .A(n32990), .B(n32914), .Z(n32917) );
  XOR U32757 ( .A(n32991), .B(n32992), .Z(n32914) );
  AND U32758 ( .A(n32993), .B(n32994), .Z(n32992) );
  XOR U32759 ( .A(n32991), .B(n32995), .Z(n32993) );
  XNOR U32760 ( .A(n32996), .B(n32997), .Z(n32990) );
  NOR U32761 ( .A(n32998), .B(n32999), .Z(n32997) );
  XOR U32762 ( .A(n32996), .B(n33000), .Z(n32998) );
  XOR U32763 ( .A(n32923), .B(n32922), .Z(n32913) );
  XNOR U32764 ( .A(n33001), .B(n32919), .Z(n32922) );
  XOR U32765 ( .A(n33002), .B(n33003), .Z(n32919) );
  AND U32766 ( .A(n33004), .B(n33005), .Z(n33003) );
  XOR U32767 ( .A(n33002), .B(n33006), .Z(n33004) );
  XNOR U32768 ( .A(n33007), .B(n33008), .Z(n33001) );
  NOR U32769 ( .A(n33009), .B(n33010), .Z(n33008) );
  XNOR U32770 ( .A(n33007), .B(n33011), .Z(n33009) );
  XOR U32771 ( .A(n33012), .B(n33013), .Z(n32923) );
  NOR U32772 ( .A(n33014), .B(n33015), .Z(n33013) );
  XNOR U32773 ( .A(n33012), .B(n33016), .Z(n33014) );
  XNOR U32774 ( .A(n32815), .B(n32929), .Z(n32931) );
  XNOR U32775 ( .A(n33017), .B(n33018), .Z(n32815) );
  AND U32776 ( .A(n382), .B(n33019), .Z(n33018) );
  XNOR U32777 ( .A(n33020), .B(n33021), .Z(n33019) );
  AND U32778 ( .A(n32821), .B(n32824), .Z(n32929) );
  XOR U32779 ( .A(n33022), .B(n32978), .Z(n32824) );
  XNOR U32780 ( .A(p_input[2048]), .B(p_input[416]), .Z(n32978) );
  XOR U32781 ( .A(n32955), .B(n32954), .Z(n33022) );
  XOR U32782 ( .A(n33023), .B(n32966), .Z(n32954) );
  XOR U32783 ( .A(n32940), .B(n32939), .Z(n32966) );
  XNOR U32784 ( .A(n33024), .B(n32945), .Z(n32939) );
  XOR U32785 ( .A(p_input[2072]), .B(p_input[440]), .Z(n32945) );
  XOR U32786 ( .A(n32936), .B(n32944), .Z(n33024) );
  XOR U32787 ( .A(n33025), .B(n32941), .Z(n32944) );
  XOR U32788 ( .A(p_input[2070]), .B(p_input[438]), .Z(n32941) );
  XNOR U32789 ( .A(p_input[2071]), .B(p_input[439]), .Z(n33025) );
  XNOR U32790 ( .A(n28684), .B(p_input[434]), .Z(n32936) );
  XNOR U32791 ( .A(n32950), .B(n32949), .Z(n32940) );
  XOR U32792 ( .A(n33026), .B(n32946), .Z(n32949) );
  XOR U32793 ( .A(p_input[2067]), .B(p_input[435]), .Z(n32946) );
  XNOR U32794 ( .A(p_input[2068]), .B(p_input[436]), .Z(n33026) );
  XOR U32795 ( .A(p_input[2069]), .B(p_input[437]), .Z(n32950) );
  XNOR U32796 ( .A(n32965), .B(n32951), .Z(n33023) );
  XNOR U32797 ( .A(n28686), .B(p_input[417]), .Z(n32951) );
  XNOR U32798 ( .A(n33027), .B(n32972), .Z(n32965) );
  XNOR U32799 ( .A(n32961), .B(n32960), .Z(n32972) );
  XOR U32800 ( .A(n33028), .B(n32957), .Z(n32960) );
  XNOR U32801 ( .A(n28322), .B(p_input[442]), .Z(n32957) );
  XNOR U32802 ( .A(p_input[2075]), .B(p_input[443]), .Z(n33028) );
  XOR U32803 ( .A(p_input[2076]), .B(p_input[444]), .Z(n32961) );
  XNOR U32804 ( .A(n32971), .B(n32962), .Z(n33027) );
  XNOR U32805 ( .A(n28689), .B(p_input[433]), .Z(n32962) );
  XOR U32806 ( .A(n33029), .B(n32977), .Z(n32971) );
  XNOR U32807 ( .A(p_input[2079]), .B(p_input[447]), .Z(n32977) );
  XOR U32808 ( .A(n32968), .B(n32976), .Z(n33029) );
  XOR U32809 ( .A(n33030), .B(n32973), .Z(n32976) );
  XOR U32810 ( .A(p_input[2077]), .B(p_input[445]), .Z(n32973) );
  XNOR U32811 ( .A(p_input[2078]), .B(p_input[446]), .Z(n33030) );
  XNOR U32812 ( .A(n28326), .B(p_input[441]), .Z(n32968) );
  XNOR U32813 ( .A(n32989), .B(n32988), .Z(n32955) );
  XNOR U32814 ( .A(n33031), .B(n32995), .Z(n32988) );
  XNOR U32815 ( .A(n32984), .B(n32983), .Z(n32995) );
  XOR U32816 ( .A(n33032), .B(n32980), .Z(n32983) );
  XNOR U32817 ( .A(n28694), .B(p_input[427]), .Z(n32980) );
  XNOR U32818 ( .A(p_input[2060]), .B(p_input[428]), .Z(n33032) );
  XOR U32819 ( .A(p_input[2061]), .B(p_input[429]), .Z(n32984) );
  XNOR U32820 ( .A(n32994), .B(n32985), .Z(n33031) );
  XNOR U32821 ( .A(n28330), .B(p_input[418]), .Z(n32985) );
  XOR U32822 ( .A(n33033), .B(n33000), .Z(n32994) );
  XNOR U32823 ( .A(p_input[2064]), .B(p_input[432]), .Z(n33000) );
  XOR U32824 ( .A(n32991), .B(n32999), .Z(n33033) );
  XOR U32825 ( .A(n33034), .B(n32996), .Z(n32999) );
  XOR U32826 ( .A(p_input[2062]), .B(p_input[430]), .Z(n32996) );
  XNOR U32827 ( .A(p_input[2063]), .B(p_input[431]), .Z(n33034) );
  XNOR U32828 ( .A(n28697), .B(p_input[426]), .Z(n32991) );
  XNOR U32829 ( .A(n33006), .B(n33005), .Z(n32989) );
  XNOR U32830 ( .A(n33035), .B(n33011), .Z(n33005) );
  XOR U32831 ( .A(p_input[2057]), .B(p_input[425]), .Z(n33011) );
  XOR U32832 ( .A(n33002), .B(n33010), .Z(n33035) );
  XOR U32833 ( .A(n33036), .B(n33007), .Z(n33010) );
  XOR U32834 ( .A(p_input[2055]), .B(p_input[423]), .Z(n33007) );
  XNOR U32835 ( .A(p_input[2056]), .B(p_input[424]), .Z(n33036) );
  XNOR U32836 ( .A(n28337), .B(p_input[419]), .Z(n33002) );
  XNOR U32837 ( .A(n33016), .B(n33015), .Z(n33006) );
  XOR U32838 ( .A(n33037), .B(n33012), .Z(n33015) );
  XOR U32839 ( .A(p_input[2052]), .B(p_input[420]), .Z(n33012) );
  XNOR U32840 ( .A(p_input[2053]), .B(p_input[421]), .Z(n33037) );
  XOR U32841 ( .A(p_input[2054]), .B(p_input[422]), .Z(n33016) );
  XNOR U32842 ( .A(n33038), .B(n33039), .Z(n32821) );
  AND U32843 ( .A(n382), .B(n33040), .Z(n33039) );
  XNOR U32844 ( .A(n33041), .B(n33042), .Z(n382) );
  AND U32845 ( .A(n33043), .B(n33044), .Z(n33042) );
  XOR U32846 ( .A(n32835), .B(n33041), .Z(n33044) );
  XNOR U32847 ( .A(n33045), .B(n33041), .Z(n33043) );
  XOR U32848 ( .A(n33046), .B(n33047), .Z(n33041) );
  AND U32849 ( .A(n33048), .B(n33049), .Z(n33047) );
  XOR U32850 ( .A(n32850), .B(n33046), .Z(n33049) );
  XOR U32851 ( .A(n33046), .B(n32851), .Z(n33048) );
  XOR U32852 ( .A(n33050), .B(n33051), .Z(n33046) );
  AND U32853 ( .A(n33052), .B(n33053), .Z(n33051) );
  XOR U32854 ( .A(n32878), .B(n33050), .Z(n33053) );
  XOR U32855 ( .A(n33050), .B(n32879), .Z(n33052) );
  XOR U32856 ( .A(n33054), .B(n33055), .Z(n33050) );
  AND U32857 ( .A(n33056), .B(n33057), .Z(n33055) );
  XOR U32858 ( .A(n32927), .B(n33054), .Z(n33057) );
  XOR U32859 ( .A(n33054), .B(n32928), .Z(n33056) );
  XOR U32860 ( .A(n33058), .B(n33059), .Z(n33054) );
  AND U32861 ( .A(n33060), .B(n33061), .Z(n33059) );
  XOR U32862 ( .A(n33058), .B(n33020), .Z(n33061) );
  XNOR U32863 ( .A(n33062), .B(n33063), .Z(n32771) );
  AND U32864 ( .A(n386), .B(n33064), .Z(n33063) );
  XNOR U32865 ( .A(n33065), .B(n33066), .Z(n386) );
  AND U32866 ( .A(n33067), .B(n33068), .Z(n33066) );
  XOR U32867 ( .A(n33065), .B(n32781), .Z(n33068) );
  XNOR U32868 ( .A(n33065), .B(n32731), .Z(n33067) );
  XOR U32869 ( .A(n33069), .B(n33070), .Z(n33065) );
  AND U32870 ( .A(n33071), .B(n33072), .Z(n33070) );
  XNOR U32871 ( .A(n32791), .B(n33069), .Z(n33072) );
  XOR U32872 ( .A(n33069), .B(n32741), .Z(n33071) );
  XOR U32873 ( .A(n33073), .B(n33074), .Z(n33069) );
  AND U32874 ( .A(n33075), .B(n33076), .Z(n33074) );
  XNOR U32875 ( .A(n32801), .B(n33073), .Z(n33076) );
  XOR U32876 ( .A(n33073), .B(n32750), .Z(n33075) );
  XOR U32877 ( .A(n33077), .B(n33078), .Z(n33073) );
  AND U32878 ( .A(n33079), .B(n33080), .Z(n33078) );
  XOR U32879 ( .A(n33077), .B(n32758), .Z(n33079) );
  XOR U32880 ( .A(n33081), .B(n33082), .Z(n32722) );
  AND U32881 ( .A(n390), .B(n33064), .Z(n33082) );
  XNOR U32882 ( .A(n33062), .B(n33081), .Z(n33064) );
  XNOR U32883 ( .A(n33083), .B(n33084), .Z(n390) );
  AND U32884 ( .A(n33085), .B(n33086), .Z(n33084) );
  XNOR U32885 ( .A(n33087), .B(n33083), .Z(n33086) );
  IV U32886 ( .A(n32781), .Z(n33087) );
  XOR U32887 ( .A(n33045), .B(n33088), .Z(n32781) );
  AND U32888 ( .A(n393), .B(n33089), .Z(n33088) );
  XOR U32889 ( .A(n32834), .B(n32831), .Z(n33089) );
  IV U32890 ( .A(n33045), .Z(n32834) );
  XNOR U32891 ( .A(n32731), .B(n33083), .Z(n33085) );
  XOR U32892 ( .A(n33090), .B(n33091), .Z(n32731) );
  AND U32893 ( .A(n409), .B(n33092), .Z(n33091) );
  XOR U32894 ( .A(n33093), .B(n33094), .Z(n33083) );
  AND U32895 ( .A(n33095), .B(n33096), .Z(n33094) );
  XNOR U32896 ( .A(n33093), .B(n32791), .Z(n33096) );
  XOR U32897 ( .A(n32851), .B(n33097), .Z(n32791) );
  AND U32898 ( .A(n393), .B(n33098), .Z(n33097) );
  XOR U32899 ( .A(n32847), .B(n32851), .Z(n33098) );
  XNOR U32900 ( .A(n33099), .B(n33093), .Z(n33095) );
  IV U32901 ( .A(n32741), .Z(n33099) );
  XOR U32902 ( .A(n33100), .B(n33101), .Z(n32741) );
  AND U32903 ( .A(n409), .B(n33102), .Z(n33101) );
  XOR U32904 ( .A(n33103), .B(n33104), .Z(n33093) );
  AND U32905 ( .A(n33105), .B(n33106), .Z(n33104) );
  XNOR U32906 ( .A(n33103), .B(n32801), .Z(n33106) );
  XOR U32907 ( .A(n32879), .B(n33107), .Z(n32801) );
  AND U32908 ( .A(n393), .B(n33108), .Z(n33107) );
  XOR U32909 ( .A(n32875), .B(n32879), .Z(n33108) );
  XOR U32910 ( .A(n32750), .B(n33103), .Z(n33105) );
  XOR U32911 ( .A(n33109), .B(n33110), .Z(n32750) );
  AND U32912 ( .A(n409), .B(n33111), .Z(n33110) );
  XOR U32913 ( .A(n33077), .B(n33112), .Z(n33103) );
  AND U32914 ( .A(n33113), .B(n33080), .Z(n33112) );
  XNOR U32915 ( .A(n32811), .B(n33077), .Z(n33080) );
  XOR U32916 ( .A(n32928), .B(n33114), .Z(n32811) );
  AND U32917 ( .A(n393), .B(n33115), .Z(n33114) );
  XOR U32918 ( .A(n32924), .B(n32928), .Z(n33115) );
  XNOR U32919 ( .A(n33116), .B(n33077), .Z(n33113) );
  IV U32920 ( .A(n32758), .Z(n33116) );
  XOR U32921 ( .A(n33117), .B(n33118), .Z(n32758) );
  AND U32922 ( .A(n409), .B(n33119), .Z(n33118) );
  XOR U32923 ( .A(n33120), .B(n33121), .Z(n33077) );
  AND U32924 ( .A(n33122), .B(n33123), .Z(n33121) );
  XNOR U32925 ( .A(n33120), .B(n32819), .Z(n33123) );
  XOR U32926 ( .A(n33021), .B(n33124), .Z(n32819) );
  AND U32927 ( .A(n393), .B(n33125), .Z(n33124) );
  XOR U32928 ( .A(n33017), .B(n33021), .Z(n33125) );
  XNOR U32929 ( .A(n33126), .B(n33120), .Z(n33122) );
  IV U32930 ( .A(n32768), .Z(n33126) );
  XOR U32931 ( .A(n33127), .B(n33128), .Z(n32768) );
  AND U32932 ( .A(n409), .B(n33129), .Z(n33128) );
  AND U32933 ( .A(n33081), .B(n33062), .Z(n33120) );
  XNOR U32934 ( .A(n33130), .B(n33131), .Z(n33062) );
  AND U32935 ( .A(n393), .B(n33040), .Z(n33131) );
  XNOR U32936 ( .A(n33038), .B(n33130), .Z(n33040) );
  XNOR U32937 ( .A(n33132), .B(n33133), .Z(n393) );
  AND U32938 ( .A(n33134), .B(n33135), .Z(n33133) );
  XNOR U32939 ( .A(n33132), .B(n32831), .Z(n33135) );
  IV U32940 ( .A(n32835), .Z(n32831) );
  XOR U32941 ( .A(n33136), .B(n33137), .Z(n32835) );
  AND U32942 ( .A(n397), .B(n33138), .Z(n33137) );
  XOR U32943 ( .A(n33139), .B(n33136), .Z(n33138) );
  XNOR U32944 ( .A(n33132), .B(n33045), .Z(n33134) );
  XOR U32945 ( .A(n33140), .B(n33141), .Z(n33045) );
  AND U32946 ( .A(n405), .B(n33092), .Z(n33141) );
  XOR U32947 ( .A(n33090), .B(n33140), .Z(n33092) );
  XOR U32948 ( .A(n33142), .B(n33143), .Z(n33132) );
  AND U32949 ( .A(n33144), .B(n33145), .Z(n33143) );
  XNOR U32950 ( .A(n33142), .B(n32847), .Z(n33145) );
  IV U32951 ( .A(n32850), .Z(n32847) );
  XOR U32952 ( .A(n33146), .B(n33147), .Z(n32850) );
  AND U32953 ( .A(n397), .B(n33148), .Z(n33147) );
  XOR U32954 ( .A(n33149), .B(n33146), .Z(n33148) );
  XOR U32955 ( .A(n32851), .B(n33142), .Z(n33144) );
  XOR U32956 ( .A(n33150), .B(n33151), .Z(n32851) );
  AND U32957 ( .A(n405), .B(n33102), .Z(n33151) );
  XOR U32958 ( .A(n33150), .B(n33100), .Z(n33102) );
  XOR U32959 ( .A(n33152), .B(n33153), .Z(n33142) );
  AND U32960 ( .A(n33154), .B(n33155), .Z(n33153) );
  XNOR U32961 ( .A(n33152), .B(n32875), .Z(n33155) );
  IV U32962 ( .A(n32878), .Z(n32875) );
  XOR U32963 ( .A(n33156), .B(n33157), .Z(n32878) );
  AND U32964 ( .A(n397), .B(n33158), .Z(n33157) );
  XNOR U32965 ( .A(n33159), .B(n33156), .Z(n33158) );
  XOR U32966 ( .A(n32879), .B(n33152), .Z(n33154) );
  XOR U32967 ( .A(n33160), .B(n33161), .Z(n32879) );
  AND U32968 ( .A(n405), .B(n33111), .Z(n33161) );
  XOR U32969 ( .A(n33160), .B(n33109), .Z(n33111) );
  XOR U32970 ( .A(n33162), .B(n33163), .Z(n33152) );
  AND U32971 ( .A(n33164), .B(n33165), .Z(n33163) );
  XNOR U32972 ( .A(n33162), .B(n32924), .Z(n33165) );
  IV U32973 ( .A(n32927), .Z(n32924) );
  XOR U32974 ( .A(n33166), .B(n33167), .Z(n32927) );
  AND U32975 ( .A(n397), .B(n33168), .Z(n33167) );
  XOR U32976 ( .A(n33169), .B(n33166), .Z(n33168) );
  XOR U32977 ( .A(n32928), .B(n33162), .Z(n33164) );
  XOR U32978 ( .A(n33170), .B(n33171), .Z(n32928) );
  AND U32979 ( .A(n405), .B(n33119), .Z(n33171) );
  XOR U32980 ( .A(n33170), .B(n33117), .Z(n33119) );
  XOR U32981 ( .A(n33058), .B(n33172), .Z(n33162) );
  AND U32982 ( .A(n33060), .B(n33173), .Z(n33172) );
  XNOR U32983 ( .A(n33058), .B(n33017), .Z(n33173) );
  IV U32984 ( .A(n33020), .Z(n33017) );
  XOR U32985 ( .A(n33174), .B(n33175), .Z(n33020) );
  AND U32986 ( .A(n397), .B(n33176), .Z(n33175) );
  XNOR U32987 ( .A(n33177), .B(n33174), .Z(n33176) );
  XOR U32988 ( .A(n33021), .B(n33058), .Z(n33060) );
  XOR U32989 ( .A(n33178), .B(n33179), .Z(n33021) );
  AND U32990 ( .A(n405), .B(n33129), .Z(n33179) );
  XOR U32991 ( .A(n33178), .B(n33127), .Z(n33129) );
  AND U32992 ( .A(n33130), .B(n33038), .Z(n33058) );
  XNOR U32993 ( .A(n33180), .B(n33181), .Z(n33038) );
  AND U32994 ( .A(n397), .B(n33182), .Z(n33181) );
  XNOR U32995 ( .A(n33183), .B(n33180), .Z(n33182) );
  XNOR U32996 ( .A(n33184), .B(n33185), .Z(n397) );
  AND U32997 ( .A(n33186), .B(n33187), .Z(n33185) );
  XOR U32998 ( .A(n33139), .B(n33184), .Z(n33187) );
  AND U32999 ( .A(n33188), .B(n33189), .Z(n33139) );
  XNOR U33000 ( .A(n33136), .B(n33184), .Z(n33186) );
  XNOR U33001 ( .A(n33190), .B(n33191), .Z(n33136) );
  AND U33002 ( .A(n401), .B(n33192), .Z(n33191) );
  XNOR U33003 ( .A(n33193), .B(n33194), .Z(n33192) );
  XOR U33004 ( .A(n33195), .B(n33196), .Z(n33184) );
  AND U33005 ( .A(n33197), .B(n33198), .Z(n33196) );
  XNOR U33006 ( .A(n33195), .B(n33188), .Z(n33198) );
  IV U33007 ( .A(n33149), .Z(n33188) );
  XOR U33008 ( .A(n33199), .B(n33200), .Z(n33149) );
  XOR U33009 ( .A(n33201), .B(n33189), .Z(n33200) );
  AND U33010 ( .A(n33159), .B(n33202), .Z(n33189) );
  AND U33011 ( .A(n33203), .B(n33204), .Z(n33201) );
  XOR U33012 ( .A(n33205), .B(n33199), .Z(n33203) );
  XNOR U33013 ( .A(n33146), .B(n33195), .Z(n33197) );
  XNOR U33014 ( .A(n33206), .B(n33207), .Z(n33146) );
  AND U33015 ( .A(n401), .B(n33208), .Z(n33207) );
  XNOR U33016 ( .A(n33209), .B(n33210), .Z(n33208) );
  XOR U33017 ( .A(n33211), .B(n33212), .Z(n33195) );
  AND U33018 ( .A(n33213), .B(n33214), .Z(n33212) );
  XNOR U33019 ( .A(n33211), .B(n33159), .Z(n33214) );
  XOR U33020 ( .A(n33215), .B(n33204), .Z(n33159) );
  XNOR U33021 ( .A(n33216), .B(n33199), .Z(n33204) );
  XOR U33022 ( .A(n33217), .B(n33218), .Z(n33199) );
  AND U33023 ( .A(n33219), .B(n33220), .Z(n33218) );
  XOR U33024 ( .A(n33221), .B(n33217), .Z(n33219) );
  XNOR U33025 ( .A(n33222), .B(n33223), .Z(n33216) );
  AND U33026 ( .A(n33224), .B(n33225), .Z(n33223) );
  XOR U33027 ( .A(n33222), .B(n33226), .Z(n33224) );
  XNOR U33028 ( .A(n33205), .B(n33202), .Z(n33215) );
  AND U33029 ( .A(n33227), .B(n33228), .Z(n33202) );
  XOR U33030 ( .A(n33229), .B(n33230), .Z(n33205) );
  AND U33031 ( .A(n33231), .B(n33232), .Z(n33230) );
  XOR U33032 ( .A(n33229), .B(n33233), .Z(n33231) );
  XNOR U33033 ( .A(n33156), .B(n33211), .Z(n33213) );
  XNOR U33034 ( .A(n33234), .B(n33235), .Z(n33156) );
  AND U33035 ( .A(n401), .B(n33236), .Z(n33235) );
  XNOR U33036 ( .A(n33237), .B(n33238), .Z(n33236) );
  XOR U33037 ( .A(n33239), .B(n33240), .Z(n33211) );
  AND U33038 ( .A(n33241), .B(n33242), .Z(n33240) );
  XNOR U33039 ( .A(n33239), .B(n33227), .Z(n33242) );
  IV U33040 ( .A(n33169), .Z(n33227) );
  XNOR U33041 ( .A(n33243), .B(n33220), .Z(n33169) );
  XNOR U33042 ( .A(n33244), .B(n33226), .Z(n33220) );
  XOR U33043 ( .A(n33245), .B(n33246), .Z(n33226) );
  AND U33044 ( .A(n33247), .B(n33248), .Z(n33246) );
  XOR U33045 ( .A(n33245), .B(n33249), .Z(n33247) );
  XNOR U33046 ( .A(n33225), .B(n33217), .Z(n33244) );
  XOR U33047 ( .A(n33250), .B(n33251), .Z(n33217) );
  AND U33048 ( .A(n33252), .B(n33253), .Z(n33251) );
  XNOR U33049 ( .A(n33254), .B(n33250), .Z(n33252) );
  XNOR U33050 ( .A(n33255), .B(n33222), .Z(n33225) );
  XOR U33051 ( .A(n33256), .B(n33257), .Z(n33222) );
  AND U33052 ( .A(n33258), .B(n33259), .Z(n33257) );
  XOR U33053 ( .A(n33256), .B(n33260), .Z(n33258) );
  XNOR U33054 ( .A(n33261), .B(n33262), .Z(n33255) );
  AND U33055 ( .A(n33263), .B(n33264), .Z(n33262) );
  XNOR U33056 ( .A(n33261), .B(n33265), .Z(n33263) );
  XNOR U33057 ( .A(n33221), .B(n33228), .Z(n33243) );
  AND U33058 ( .A(n33177), .B(n33266), .Z(n33228) );
  XOR U33059 ( .A(n33233), .B(n33232), .Z(n33221) );
  XNOR U33060 ( .A(n33267), .B(n33229), .Z(n33232) );
  XOR U33061 ( .A(n33268), .B(n33269), .Z(n33229) );
  AND U33062 ( .A(n33270), .B(n33271), .Z(n33269) );
  XOR U33063 ( .A(n33268), .B(n33272), .Z(n33270) );
  XNOR U33064 ( .A(n33273), .B(n33274), .Z(n33267) );
  AND U33065 ( .A(n33275), .B(n33276), .Z(n33274) );
  XOR U33066 ( .A(n33273), .B(n33277), .Z(n33275) );
  XOR U33067 ( .A(n33278), .B(n33279), .Z(n33233) );
  AND U33068 ( .A(n33280), .B(n33281), .Z(n33279) );
  XOR U33069 ( .A(n33278), .B(n33282), .Z(n33280) );
  XNOR U33070 ( .A(n33166), .B(n33239), .Z(n33241) );
  XNOR U33071 ( .A(n33283), .B(n33284), .Z(n33166) );
  AND U33072 ( .A(n401), .B(n33285), .Z(n33284) );
  XNOR U33073 ( .A(n33286), .B(n33287), .Z(n33285) );
  XOR U33074 ( .A(n33288), .B(n33289), .Z(n33239) );
  AND U33075 ( .A(n33290), .B(n33291), .Z(n33289) );
  XNOR U33076 ( .A(n33288), .B(n33177), .Z(n33291) );
  XOR U33077 ( .A(n33292), .B(n33253), .Z(n33177) );
  XNOR U33078 ( .A(n33293), .B(n33260), .Z(n33253) );
  XOR U33079 ( .A(n33249), .B(n33248), .Z(n33260) );
  XNOR U33080 ( .A(n33294), .B(n33245), .Z(n33248) );
  XOR U33081 ( .A(n33295), .B(n33296), .Z(n33245) );
  AND U33082 ( .A(n33297), .B(n33298), .Z(n33296) );
  XOR U33083 ( .A(n33295), .B(n33299), .Z(n33297) );
  XNOR U33084 ( .A(n33300), .B(n33301), .Z(n33294) );
  NOR U33085 ( .A(n33302), .B(n33303), .Z(n33301) );
  XNOR U33086 ( .A(n33300), .B(n33304), .Z(n33302) );
  XOR U33087 ( .A(n33305), .B(n33306), .Z(n33249) );
  NOR U33088 ( .A(n33307), .B(n33308), .Z(n33306) );
  XNOR U33089 ( .A(n33305), .B(n33309), .Z(n33307) );
  XNOR U33090 ( .A(n33259), .B(n33250), .Z(n33293) );
  XOR U33091 ( .A(n33310), .B(n33311), .Z(n33250) );
  NOR U33092 ( .A(n33312), .B(n33313), .Z(n33311) );
  XNOR U33093 ( .A(n33310), .B(n33314), .Z(n33312) );
  XOR U33094 ( .A(n33315), .B(n33265), .Z(n33259) );
  XNOR U33095 ( .A(n33316), .B(n33317), .Z(n33265) );
  NOR U33096 ( .A(n33318), .B(n33319), .Z(n33317) );
  XNOR U33097 ( .A(n33316), .B(n33320), .Z(n33318) );
  XNOR U33098 ( .A(n33264), .B(n33256), .Z(n33315) );
  XOR U33099 ( .A(n33321), .B(n33322), .Z(n33256) );
  AND U33100 ( .A(n33323), .B(n33324), .Z(n33322) );
  XOR U33101 ( .A(n33321), .B(n33325), .Z(n33323) );
  XNOR U33102 ( .A(n33326), .B(n33261), .Z(n33264) );
  XOR U33103 ( .A(n33327), .B(n33328), .Z(n33261) );
  AND U33104 ( .A(n33329), .B(n33330), .Z(n33328) );
  XOR U33105 ( .A(n33327), .B(n33331), .Z(n33329) );
  XNOR U33106 ( .A(n33332), .B(n33333), .Z(n33326) );
  NOR U33107 ( .A(n33334), .B(n33335), .Z(n33333) );
  XOR U33108 ( .A(n33332), .B(n33336), .Z(n33334) );
  XOR U33109 ( .A(n33254), .B(n33266), .Z(n33292) );
  NOR U33110 ( .A(n33183), .B(n33337), .Z(n33266) );
  XNOR U33111 ( .A(n33272), .B(n33271), .Z(n33254) );
  XNOR U33112 ( .A(n33338), .B(n33277), .Z(n33271) );
  XOR U33113 ( .A(n33339), .B(n33340), .Z(n33277) );
  NOR U33114 ( .A(n33341), .B(n33342), .Z(n33340) );
  XNOR U33115 ( .A(n33339), .B(n33343), .Z(n33341) );
  XNOR U33116 ( .A(n33276), .B(n33268), .Z(n33338) );
  XOR U33117 ( .A(n33344), .B(n33345), .Z(n33268) );
  AND U33118 ( .A(n33346), .B(n33347), .Z(n33345) );
  XNOR U33119 ( .A(n33344), .B(n33348), .Z(n33346) );
  XNOR U33120 ( .A(n33349), .B(n33273), .Z(n33276) );
  XOR U33121 ( .A(n33350), .B(n33351), .Z(n33273) );
  AND U33122 ( .A(n33352), .B(n33353), .Z(n33351) );
  XOR U33123 ( .A(n33350), .B(n33354), .Z(n33352) );
  XNOR U33124 ( .A(n33355), .B(n33356), .Z(n33349) );
  NOR U33125 ( .A(n33357), .B(n33358), .Z(n33356) );
  XOR U33126 ( .A(n33355), .B(n33359), .Z(n33357) );
  XOR U33127 ( .A(n33282), .B(n33281), .Z(n33272) );
  XNOR U33128 ( .A(n33360), .B(n33278), .Z(n33281) );
  XOR U33129 ( .A(n33361), .B(n33362), .Z(n33278) );
  AND U33130 ( .A(n33363), .B(n33364), .Z(n33362) );
  XOR U33131 ( .A(n33361), .B(n33365), .Z(n33363) );
  XNOR U33132 ( .A(n33366), .B(n33367), .Z(n33360) );
  NOR U33133 ( .A(n33368), .B(n33369), .Z(n33367) );
  XNOR U33134 ( .A(n33366), .B(n33370), .Z(n33368) );
  XOR U33135 ( .A(n33371), .B(n33372), .Z(n33282) );
  NOR U33136 ( .A(n33373), .B(n33374), .Z(n33372) );
  XNOR U33137 ( .A(n33371), .B(n33375), .Z(n33373) );
  XNOR U33138 ( .A(n33174), .B(n33288), .Z(n33290) );
  XNOR U33139 ( .A(n33376), .B(n33377), .Z(n33174) );
  AND U33140 ( .A(n401), .B(n33378), .Z(n33377) );
  XNOR U33141 ( .A(n33379), .B(n33380), .Z(n33378) );
  AND U33142 ( .A(n33180), .B(n33183), .Z(n33288) );
  XOR U33143 ( .A(n33381), .B(n33337), .Z(n33183) );
  XNOR U33144 ( .A(p_input[2048]), .B(p_input[448]), .Z(n33337) );
  XOR U33145 ( .A(n33314), .B(n33313), .Z(n33381) );
  XOR U33146 ( .A(n33382), .B(n33325), .Z(n33313) );
  XOR U33147 ( .A(n33299), .B(n33298), .Z(n33325) );
  XNOR U33148 ( .A(n33383), .B(n33304), .Z(n33298) );
  XOR U33149 ( .A(p_input[2072]), .B(p_input[472]), .Z(n33304) );
  XOR U33150 ( .A(n33295), .B(n33303), .Z(n33383) );
  XOR U33151 ( .A(n33384), .B(n33300), .Z(n33303) );
  XOR U33152 ( .A(p_input[2070]), .B(p_input[470]), .Z(n33300) );
  XNOR U33153 ( .A(p_input[2071]), .B(p_input[471]), .Z(n33384) );
  XNOR U33154 ( .A(n28684), .B(p_input[466]), .Z(n33295) );
  XNOR U33155 ( .A(n33309), .B(n33308), .Z(n33299) );
  XOR U33156 ( .A(n33385), .B(n33305), .Z(n33308) );
  XOR U33157 ( .A(p_input[2067]), .B(p_input[467]), .Z(n33305) );
  XNOR U33158 ( .A(p_input[2068]), .B(p_input[468]), .Z(n33385) );
  XOR U33159 ( .A(p_input[2069]), .B(p_input[469]), .Z(n33309) );
  XNOR U33160 ( .A(n33324), .B(n33310), .Z(n33382) );
  XNOR U33161 ( .A(n28686), .B(p_input[449]), .Z(n33310) );
  XNOR U33162 ( .A(n33386), .B(n33331), .Z(n33324) );
  XNOR U33163 ( .A(n33320), .B(n33319), .Z(n33331) );
  XOR U33164 ( .A(n33387), .B(n33316), .Z(n33319) );
  XNOR U33165 ( .A(n28322), .B(p_input[474]), .Z(n33316) );
  XNOR U33166 ( .A(p_input[2075]), .B(p_input[475]), .Z(n33387) );
  XOR U33167 ( .A(p_input[2076]), .B(p_input[476]), .Z(n33320) );
  XNOR U33168 ( .A(n33330), .B(n33321), .Z(n33386) );
  XNOR U33169 ( .A(n28689), .B(p_input[465]), .Z(n33321) );
  XOR U33170 ( .A(n33388), .B(n33336), .Z(n33330) );
  XNOR U33171 ( .A(p_input[2079]), .B(p_input[479]), .Z(n33336) );
  XOR U33172 ( .A(n33327), .B(n33335), .Z(n33388) );
  XOR U33173 ( .A(n33389), .B(n33332), .Z(n33335) );
  XOR U33174 ( .A(p_input[2077]), .B(p_input[477]), .Z(n33332) );
  XNOR U33175 ( .A(p_input[2078]), .B(p_input[478]), .Z(n33389) );
  XNOR U33176 ( .A(n28326), .B(p_input[473]), .Z(n33327) );
  XNOR U33177 ( .A(n33348), .B(n33347), .Z(n33314) );
  XNOR U33178 ( .A(n33390), .B(n33354), .Z(n33347) );
  XNOR U33179 ( .A(n33343), .B(n33342), .Z(n33354) );
  XOR U33180 ( .A(n33391), .B(n33339), .Z(n33342) );
  XNOR U33181 ( .A(n28694), .B(p_input[459]), .Z(n33339) );
  XNOR U33182 ( .A(p_input[2060]), .B(p_input[460]), .Z(n33391) );
  XOR U33183 ( .A(p_input[2061]), .B(p_input[461]), .Z(n33343) );
  XNOR U33184 ( .A(n33353), .B(n33344), .Z(n33390) );
  XNOR U33185 ( .A(n28330), .B(p_input[450]), .Z(n33344) );
  XOR U33186 ( .A(n33392), .B(n33359), .Z(n33353) );
  XNOR U33187 ( .A(p_input[2064]), .B(p_input[464]), .Z(n33359) );
  XOR U33188 ( .A(n33350), .B(n33358), .Z(n33392) );
  XOR U33189 ( .A(n33393), .B(n33355), .Z(n33358) );
  XOR U33190 ( .A(p_input[2062]), .B(p_input[462]), .Z(n33355) );
  XNOR U33191 ( .A(p_input[2063]), .B(p_input[463]), .Z(n33393) );
  XNOR U33192 ( .A(n28697), .B(p_input[458]), .Z(n33350) );
  XNOR U33193 ( .A(n33365), .B(n33364), .Z(n33348) );
  XNOR U33194 ( .A(n33394), .B(n33370), .Z(n33364) );
  XOR U33195 ( .A(p_input[2057]), .B(p_input[457]), .Z(n33370) );
  XOR U33196 ( .A(n33361), .B(n33369), .Z(n33394) );
  XOR U33197 ( .A(n33395), .B(n33366), .Z(n33369) );
  XOR U33198 ( .A(p_input[2055]), .B(p_input[455]), .Z(n33366) );
  XNOR U33199 ( .A(p_input[2056]), .B(p_input[456]), .Z(n33395) );
  XNOR U33200 ( .A(n28337), .B(p_input[451]), .Z(n33361) );
  XNOR U33201 ( .A(n33375), .B(n33374), .Z(n33365) );
  XOR U33202 ( .A(n33396), .B(n33371), .Z(n33374) );
  XOR U33203 ( .A(p_input[2052]), .B(p_input[452]), .Z(n33371) );
  XNOR U33204 ( .A(p_input[2053]), .B(p_input[453]), .Z(n33396) );
  XOR U33205 ( .A(p_input[2054]), .B(p_input[454]), .Z(n33375) );
  XNOR U33206 ( .A(n33397), .B(n33398), .Z(n33180) );
  AND U33207 ( .A(n401), .B(n33399), .Z(n33398) );
  XNOR U33208 ( .A(n33400), .B(n33401), .Z(n401) );
  AND U33209 ( .A(n33402), .B(n33403), .Z(n33401) );
  XOR U33210 ( .A(n33194), .B(n33400), .Z(n33403) );
  XNOR U33211 ( .A(n33404), .B(n33400), .Z(n33402) );
  XOR U33212 ( .A(n33405), .B(n33406), .Z(n33400) );
  AND U33213 ( .A(n33407), .B(n33408), .Z(n33406) );
  XOR U33214 ( .A(n33209), .B(n33405), .Z(n33408) );
  XOR U33215 ( .A(n33405), .B(n33210), .Z(n33407) );
  XOR U33216 ( .A(n33409), .B(n33410), .Z(n33405) );
  AND U33217 ( .A(n33411), .B(n33412), .Z(n33410) );
  XOR U33218 ( .A(n33237), .B(n33409), .Z(n33412) );
  XOR U33219 ( .A(n33409), .B(n33238), .Z(n33411) );
  XOR U33220 ( .A(n33413), .B(n33414), .Z(n33409) );
  AND U33221 ( .A(n33415), .B(n33416), .Z(n33414) );
  XOR U33222 ( .A(n33286), .B(n33413), .Z(n33416) );
  XOR U33223 ( .A(n33413), .B(n33287), .Z(n33415) );
  XOR U33224 ( .A(n33417), .B(n33418), .Z(n33413) );
  AND U33225 ( .A(n33419), .B(n33420), .Z(n33418) );
  XOR U33226 ( .A(n33417), .B(n33379), .Z(n33420) );
  XNOR U33227 ( .A(n33421), .B(n33422), .Z(n33130) );
  AND U33228 ( .A(n405), .B(n33423), .Z(n33422) );
  XNOR U33229 ( .A(n33424), .B(n33425), .Z(n405) );
  AND U33230 ( .A(n33426), .B(n33427), .Z(n33425) );
  XOR U33231 ( .A(n33424), .B(n33140), .Z(n33427) );
  XNOR U33232 ( .A(n33424), .B(n33090), .Z(n33426) );
  XOR U33233 ( .A(n33428), .B(n33429), .Z(n33424) );
  AND U33234 ( .A(n33430), .B(n33431), .Z(n33429) );
  XNOR U33235 ( .A(n33150), .B(n33428), .Z(n33431) );
  XOR U33236 ( .A(n33428), .B(n33100), .Z(n33430) );
  XOR U33237 ( .A(n33432), .B(n33433), .Z(n33428) );
  AND U33238 ( .A(n33434), .B(n33435), .Z(n33433) );
  XNOR U33239 ( .A(n33160), .B(n33432), .Z(n33435) );
  XOR U33240 ( .A(n33432), .B(n33109), .Z(n33434) );
  XOR U33241 ( .A(n33436), .B(n33437), .Z(n33432) );
  AND U33242 ( .A(n33438), .B(n33439), .Z(n33437) );
  XOR U33243 ( .A(n33436), .B(n33117), .Z(n33438) );
  XOR U33244 ( .A(n33440), .B(n33441), .Z(n33081) );
  AND U33245 ( .A(n409), .B(n33423), .Z(n33441) );
  XNOR U33246 ( .A(n33421), .B(n33440), .Z(n33423) );
  XNOR U33247 ( .A(n33442), .B(n33443), .Z(n409) );
  AND U33248 ( .A(n33444), .B(n33445), .Z(n33443) );
  XNOR U33249 ( .A(n33446), .B(n33442), .Z(n33445) );
  IV U33250 ( .A(n33140), .Z(n33446) );
  XOR U33251 ( .A(n33404), .B(n33447), .Z(n33140) );
  AND U33252 ( .A(n412), .B(n33448), .Z(n33447) );
  XOR U33253 ( .A(n33193), .B(n33190), .Z(n33448) );
  IV U33254 ( .A(n33404), .Z(n33193) );
  XNOR U33255 ( .A(n33090), .B(n33442), .Z(n33444) );
  XOR U33256 ( .A(n33449), .B(n33450), .Z(n33090) );
  AND U33257 ( .A(n428), .B(n33451), .Z(n33450) );
  XOR U33258 ( .A(n33452), .B(n33453), .Z(n33442) );
  AND U33259 ( .A(n33454), .B(n33455), .Z(n33453) );
  XNOR U33260 ( .A(n33452), .B(n33150), .Z(n33455) );
  XOR U33261 ( .A(n33210), .B(n33456), .Z(n33150) );
  AND U33262 ( .A(n412), .B(n33457), .Z(n33456) );
  XOR U33263 ( .A(n33206), .B(n33210), .Z(n33457) );
  XNOR U33264 ( .A(n33458), .B(n33452), .Z(n33454) );
  IV U33265 ( .A(n33100), .Z(n33458) );
  XOR U33266 ( .A(n33459), .B(n33460), .Z(n33100) );
  AND U33267 ( .A(n428), .B(n33461), .Z(n33460) );
  XOR U33268 ( .A(n33462), .B(n33463), .Z(n33452) );
  AND U33269 ( .A(n33464), .B(n33465), .Z(n33463) );
  XNOR U33270 ( .A(n33462), .B(n33160), .Z(n33465) );
  XOR U33271 ( .A(n33238), .B(n33466), .Z(n33160) );
  AND U33272 ( .A(n412), .B(n33467), .Z(n33466) );
  XOR U33273 ( .A(n33234), .B(n33238), .Z(n33467) );
  XOR U33274 ( .A(n33109), .B(n33462), .Z(n33464) );
  XOR U33275 ( .A(n33468), .B(n33469), .Z(n33109) );
  AND U33276 ( .A(n428), .B(n33470), .Z(n33469) );
  XOR U33277 ( .A(n33436), .B(n33471), .Z(n33462) );
  AND U33278 ( .A(n33472), .B(n33439), .Z(n33471) );
  XNOR U33279 ( .A(n33170), .B(n33436), .Z(n33439) );
  XOR U33280 ( .A(n33287), .B(n33473), .Z(n33170) );
  AND U33281 ( .A(n412), .B(n33474), .Z(n33473) );
  XOR U33282 ( .A(n33283), .B(n33287), .Z(n33474) );
  XNOR U33283 ( .A(n33475), .B(n33436), .Z(n33472) );
  IV U33284 ( .A(n33117), .Z(n33475) );
  XOR U33285 ( .A(n33476), .B(n33477), .Z(n33117) );
  AND U33286 ( .A(n428), .B(n33478), .Z(n33477) );
  XOR U33287 ( .A(n33479), .B(n33480), .Z(n33436) );
  AND U33288 ( .A(n33481), .B(n33482), .Z(n33480) );
  XNOR U33289 ( .A(n33479), .B(n33178), .Z(n33482) );
  XOR U33290 ( .A(n33380), .B(n33483), .Z(n33178) );
  AND U33291 ( .A(n412), .B(n33484), .Z(n33483) );
  XOR U33292 ( .A(n33376), .B(n33380), .Z(n33484) );
  XNOR U33293 ( .A(n33485), .B(n33479), .Z(n33481) );
  IV U33294 ( .A(n33127), .Z(n33485) );
  XOR U33295 ( .A(n33486), .B(n33487), .Z(n33127) );
  AND U33296 ( .A(n428), .B(n33488), .Z(n33487) );
  AND U33297 ( .A(n33440), .B(n33421), .Z(n33479) );
  XNOR U33298 ( .A(n33489), .B(n33490), .Z(n33421) );
  AND U33299 ( .A(n412), .B(n33399), .Z(n33490) );
  XNOR U33300 ( .A(n33397), .B(n33489), .Z(n33399) );
  XNOR U33301 ( .A(n33491), .B(n33492), .Z(n412) );
  AND U33302 ( .A(n33493), .B(n33494), .Z(n33492) );
  XNOR U33303 ( .A(n33491), .B(n33190), .Z(n33494) );
  IV U33304 ( .A(n33194), .Z(n33190) );
  XOR U33305 ( .A(n33495), .B(n33496), .Z(n33194) );
  AND U33306 ( .A(n416), .B(n33497), .Z(n33496) );
  XOR U33307 ( .A(n33498), .B(n33495), .Z(n33497) );
  XNOR U33308 ( .A(n33491), .B(n33404), .Z(n33493) );
  XOR U33309 ( .A(n33499), .B(n33500), .Z(n33404) );
  AND U33310 ( .A(n424), .B(n33451), .Z(n33500) );
  XOR U33311 ( .A(n33449), .B(n33499), .Z(n33451) );
  XOR U33312 ( .A(n33501), .B(n33502), .Z(n33491) );
  AND U33313 ( .A(n33503), .B(n33504), .Z(n33502) );
  XNOR U33314 ( .A(n33501), .B(n33206), .Z(n33504) );
  IV U33315 ( .A(n33209), .Z(n33206) );
  XOR U33316 ( .A(n33505), .B(n33506), .Z(n33209) );
  AND U33317 ( .A(n416), .B(n33507), .Z(n33506) );
  XOR U33318 ( .A(n33508), .B(n33505), .Z(n33507) );
  XOR U33319 ( .A(n33210), .B(n33501), .Z(n33503) );
  XOR U33320 ( .A(n33509), .B(n33510), .Z(n33210) );
  AND U33321 ( .A(n424), .B(n33461), .Z(n33510) );
  XOR U33322 ( .A(n33509), .B(n33459), .Z(n33461) );
  XOR U33323 ( .A(n33511), .B(n33512), .Z(n33501) );
  AND U33324 ( .A(n33513), .B(n33514), .Z(n33512) );
  XNOR U33325 ( .A(n33511), .B(n33234), .Z(n33514) );
  IV U33326 ( .A(n33237), .Z(n33234) );
  XOR U33327 ( .A(n33515), .B(n33516), .Z(n33237) );
  AND U33328 ( .A(n416), .B(n33517), .Z(n33516) );
  XNOR U33329 ( .A(n33518), .B(n33515), .Z(n33517) );
  XOR U33330 ( .A(n33238), .B(n33511), .Z(n33513) );
  XOR U33331 ( .A(n33519), .B(n33520), .Z(n33238) );
  AND U33332 ( .A(n424), .B(n33470), .Z(n33520) );
  XOR U33333 ( .A(n33519), .B(n33468), .Z(n33470) );
  XOR U33334 ( .A(n33521), .B(n33522), .Z(n33511) );
  AND U33335 ( .A(n33523), .B(n33524), .Z(n33522) );
  XNOR U33336 ( .A(n33521), .B(n33283), .Z(n33524) );
  IV U33337 ( .A(n33286), .Z(n33283) );
  XOR U33338 ( .A(n33525), .B(n33526), .Z(n33286) );
  AND U33339 ( .A(n416), .B(n33527), .Z(n33526) );
  XOR U33340 ( .A(n33528), .B(n33525), .Z(n33527) );
  XOR U33341 ( .A(n33287), .B(n33521), .Z(n33523) );
  XOR U33342 ( .A(n33529), .B(n33530), .Z(n33287) );
  AND U33343 ( .A(n424), .B(n33478), .Z(n33530) );
  XOR U33344 ( .A(n33529), .B(n33476), .Z(n33478) );
  XOR U33345 ( .A(n33417), .B(n33531), .Z(n33521) );
  AND U33346 ( .A(n33419), .B(n33532), .Z(n33531) );
  XNOR U33347 ( .A(n33417), .B(n33376), .Z(n33532) );
  IV U33348 ( .A(n33379), .Z(n33376) );
  XOR U33349 ( .A(n33533), .B(n33534), .Z(n33379) );
  AND U33350 ( .A(n416), .B(n33535), .Z(n33534) );
  XNOR U33351 ( .A(n33536), .B(n33533), .Z(n33535) );
  XOR U33352 ( .A(n33380), .B(n33417), .Z(n33419) );
  XOR U33353 ( .A(n33537), .B(n33538), .Z(n33380) );
  AND U33354 ( .A(n424), .B(n33488), .Z(n33538) );
  XOR U33355 ( .A(n33537), .B(n33486), .Z(n33488) );
  AND U33356 ( .A(n33489), .B(n33397), .Z(n33417) );
  XNOR U33357 ( .A(n33539), .B(n33540), .Z(n33397) );
  AND U33358 ( .A(n416), .B(n33541), .Z(n33540) );
  XNOR U33359 ( .A(n33542), .B(n33539), .Z(n33541) );
  XNOR U33360 ( .A(n33543), .B(n33544), .Z(n416) );
  AND U33361 ( .A(n33545), .B(n33546), .Z(n33544) );
  XOR U33362 ( .A(n33498), .B(n33543), .Z(n33546) );
  AND U33363 ( .A(n33547), .B(n33548), .Z(n33498) );
  XNOR U33364 ( .A(n33495), .B(n33543), .Z(n33545) );
  XNOR U33365 ( .A(n33549), .B(n33550), .Z(n33495) );
  AND U33366 ( .A(n420), .B(n33551), .Z(n33550) );
  XNOR U33367 ( .A(n33552), .B(n33553), .Z(n33551) );
  XOR U33368 ( .A(n33554), .B(n33555), .Z(n33543) );
  AND U33369 ( .A(n33556), .B(n33557), .Z(n33555) );
  XNOR U33370 ( .A(n33554), .B(n33547), .Z(n33557) );
  IV U33371 ( .A(n33508), .Z(n33547) );
  XOR U33372 ( .A(n33558), .B(n33559), .Z(n33508) );
  XOR U33373 ( .A(n33560), .B(n33548), .Z(n33559) );
  AND U33374 ( .A(n33518), .B(n33561), .Z(n33548) );
  AND U33375 ( .A(n33562), .B(n33563), .Z(n33560) );
  XOR U33376 ( .A(n33564), .B(n33558), .Z(n33562) );
  XNOR U33377 ( .A(n33505), .B(n33554), .Z(n33556) );
  XNOR U33378 ( .A(n33565), .B(n33566), .Z(n33505) );
  AND U33379 ( .A(n420), .B(n33567), .Z(n33566) );
  XNOR U33380 ( .A(n33568), .B(n33569), .Z(n33567) );
  XOR U33381 ( .A(n33570), .B(n33571), .Z(n33554) );
  AND U33382 ( .A(n33572), .B(n33573), .Z(n33571) );
  XNOR U33383 ( .A(n33570), .B(n33518), .Z(n33573) );
  XOR U33384 ( .A(n33574), .B(n33563), .Z(n33518) );
  XNOR U33385 ( .A(n33575), .B(n33558), .Z(n33563) );
  XOR U33386 ( .A(n33576), .B(n33577), .Z(n33558) );
  AND U33387 ( .A(n33578), .B(n33579), .Z(n33577) );
  XOR U33388 ( .A(n33580), .B(n33576), .Z(n33578) );
  XNOR U33389 ( .A(n33581), .B(n33582), .Z(n33575) );
  AND U33390 ( .A(n33583), .B(n33584), .Z(n33582) );
  XOR U33391 ( .A(n33581), .B(n33585), .Z(n33583) );
  XNOR U33392 ( .A(n33564), .B(n33561), .Z(n33574) );
  AND U33393 ( .A(n33586), .B(n33587), .Z(n33561) );
  XOR U33394 ( .A(n33588), .B(n33589), .Z(n33564) );
  AND U33395 ( .A(n33590), .B(n33591), .Z(n33589) );
  XOR U33396 ( .A(n33588), .B(n33592), .Z(n33590) );
  XNOR U33397 ( .A(n33515), .B(n33570), .Z(n33572) );
  XNOR U33398 ( .A(n33593), .B(n33594), .Z(n33515) );
  AND U33399 ( .A(n420), .B(n33595), .Z(n33594) );
  XNOR U33400 ( .A(n33596), .B(n33597), .Z(n33595) );
  XOR U33401 ( .A(n33598), .B(n33599), .Z(n33570) );
  AND U33402 ( .A(n33600), .B(n33601), .Z(n33599) );
  XNOR U33403 ( .A(n33598), .B(n33586), .Z(n33601) );
  IV U33404 ( .A(n33528), .Z(n33586) );
  XNOR U33405 ( .A(n33602), .B(n33579), .Z(n33528) );
  XNOR U33406 ( .A(n33603), .B(n33585), .Z(n33579) );
  XOR U33407 ( .A(n33604), .B(n33605), .Z(n33585) );
  AND U33408 ( .A(n33606), .B(n33607), .Z(n33605) );
  XOR U33409 ( .A(n33604), .B(n33608), .Z(n33606) );
  XNOR U33410 ( .A(n33584), .B(n33576), .Z(n33603) );
  XOR U33411 ( .A(n33609), .B(n33610), .Z(n33576) );
  AND U33412 ( .A(n33611), .B(n33612), .Z(n33610) );
  XNOR U33413 ( .A(n33613), .B(n33609), .Z(n33611) );
  XNOR U33414 ( .A(n33614), .B(n33581), .Z(n33584) );
  XOR U33415 ( .A(n33615), .B(n33616), .Z(n33581) );
  AND U33416 ( .A(n33617), .B(n33618), .Z(n33616) );
  XOR U33417 ( .A(n33615), .B(n33619), .Z(n33617) );
  XNOR U33418 ( .A(n33620), .B(n33621), .Z(n33614) );
  AND U33419 ( .A(n33622), .B(n33623), .Z(n33621) );
  XNOR U33420 ( .A(n33620), .B(n33624), .Z(n33622) );
  XNOR U33421 ( .A(n33580), .B(n33587), .Z(n33602) );
  AND U33422 ( .A(n33536), .B(n33625), .Z(n33587) );
  XOR U33423 ( .A(n33592), .B(n33591), .Z(n33580) );
  XNOR U33424 ( .A(n33626), .B(n33588), .Z(n33591) );
  XOR U33425 ( .A(n33627), .B(n33628), .Z(n33588) );
  AND U33426 ( .A(n33629), .B(n33630), .Z(n33628) );
  XOR U33427 ( .A(n33627), .B(n33631), .Z(n33629) );
  XNOR U33428 ( .A(n33632), .B(n33633), .Z(n33626) );
  AND U33429 ( .A(n33634), .B(n33635), .Z(n33633) );
  XOR U33430 ( .A(n33632), .B(n33636), .Z(n33634) );
  XOR U33431 ( .A(n33637), .B(n33638), .Z(n33592) );
  AND U33432 ( .A(n33639), .B(n33640), .Z(n33638) );
  XOR U33433 ( .A(n33637), .B(n33641), .Z(n33639) );
  XNOR U33434 ( .A(n33525), .B(n33598), .Z(n33600) );
  XNOR U33435 ( .A(n33642), .B(n33643), .Z(n33525) );
  AND U33436 ( .A(n420), .B(n33644), .Z(n33643) );
  XNOR U33437 ( .A(n33645), .B(n33646), .Z(n33644) );
  XOR U33438 ( .A(n33647), .B(n33648), .Z(n33598) );
  AND U33439 ( .A(n33649), .B(n33650), .Z(n33648) );
  XNOR U33440 ( .A(n33647), .B(n33536), .Z(n33650) );
  XOR U33441 ( .A(n33651), .B(n33612), .Z(n33536) );
  XNOR U33442 ( .A(n33652), .B(n33619), .Z(n33612) );
  XOR U33443 ( .A(n33608), .B(n33607), .Z(n33619) );
  XNOR U33444 ( .A(n33653), .B(n33604), .Z(n33607) );
  XOR U33445 ( .A(n33654), .B(n33655), .Z(n33604) );
  AND U33446 ( .A(n33656), .B(n33657), .Z(n33655) );
  XOR U33447 ( .A(n33654), .B(n33658), .Z(n33656) );
  XNOR U33448 ( .A(n33659), .B(n33660), .Z(n33653) );
  NOR U33449 ( .A(n33661), .B(n33662), .Z(n33660) );
  XNOR U33450 ( .A(n33659), .B(n33663), .Z(n33661) );
  XOR U33451 ( .A(n33664), .B(n33665), .Z(n33608) );
  NOR U33452 ( .A(n33666), .B(n33667), .Z(n33665) );
  XNOR U33453 ( .A(n33664), .B(n33668), .Z(n33666) );
  XNOR U33454 ( .A(n33618), .B(n33609), .Z(n33652) );
  XOR U33455 ( .A(n33669), .B(n33670), .Z(n33609) );
  NOR U33456 ( .A(n33671), .B(n33672), .Z(n33670) );
  XNOR U33457 ( .A(n33669), .B(n33673), .Z(n33671) );
  XOR U33458 ( .A(n33674), .B(n33624), .Z(n33618) );
  XNOR U33459 ( .A(n33675), .B(n33676), .Z(n33624) );
  NOR U33460 ( .A(n33677), .B(n33678), .Z(n33676) );
  XNOR U33461 ( .A(n33675), .B(n33679), .Z(n33677) );
  XNOR U33462 ( .A(n33623), .B(n33615), .Z(n33674) );
  XOR U33463 ( .A(n33680), .B(n33681), .Z(n33615) );
  AND U33464 ( .A(n33682), .B(n33683), .Z(n33681) );
  XOR U33465 ( .A(n33680), .B(n33684), .Z(n33682) );
  XNOR U33466 ( .A(n33685), .B(n33620), .Z(n33623) );
  XOR U33467 ( .A(n33686), .B(n33687), .Z(n33620) );
  AND U33468 ( .A(n33688), .B(n33689), .Z(n33687) );
  XOR U33469 ( .A(n33686), .B(n33690), .Z(n33688) );
  XNOR U33470 ( .A(n33691), .B(n33692), .Z(n33685) );
  NOR U33471 ( .A(n33693), .B(n33694), .Z(n33692) );
  XOR U33472 ( .A(n33691), .B(n33695), .Z(n33693) );
  XOR U33473 ( .A(n33613), .B(n33625), .Z(n33651) );
  NOR U33474 ( .A(n33542), .B(n33696), .Z(n33625) );
  XNOR U33475 ( .A(n33631), .B(n33630), .Z(n33613) );
  XNOR U33476 ( .A(n33697), .B(n33636), .Z(n33630) );
  XOR U33477 ( .A(n33698), .B(n33699), .Z(n33636) );
  NOR U33478 ( .A(n33700), .B(n33701), .Z(n33699) );
  XNOR U33479 ( .A(n33698), .B(n33702), .Z(n33700) );
  XNOR U33480 ( .A(n33635), .B(n33627), .Z(n33697) );
  XOR U33481 ( .A(n33703), .B(n33704), .Z(n33627) );
  AND U33482 ( .A(n33705), .B(n33706), .Z(n33704) );
  XNOR U33483 ( .A(n33703), .B(n33707), .Z(n33705) );
  XNOR U33484 ( .A(n33708), .B(n33632), .Z(n33635) );
  XOR U33485 ( .A(n33709), .B(n33710), .Z(n33632) );
  AND U33486 ( .A(n33711), .B(n33712), .Z(n33710) );
  XOR U33487 ( .A(n33709), .B(n33713), .Z(n33711) );
  XNOR U33488 ( .A(n33714), .B(n33715), .Z(n33708) );
  NOR U33489 ( .A(n33716), .B(n33717), .Z(n33715) );
  XOR U33490 ( .A(n33714), .B(n33718), .Z(n33716) );
  XOR U33491 ( .A(n33641), .B(n33640), .Z(n33631) );
  XNOR U33492 ( .A(n33719), .B(n33637), .Z(n33640) );
  XOR U33493 ( .A(n33720), .B(n33721), .Z(n33637) );
  AND U33494 ( .A(n33722), .B(n33723), .Z(n33721) );
  XOR U33495 ( .A(n33720), .B(n33724), .Z(n33722) );
  XNOR U33496 ( .A(n33725), .B(n33726), .Z(n33719) );
  NOR U33497 ( .A(n33727), .B(n33728), .Z(n33726) );
  XNOR U33498 ( .A(n33725), .B(n33729), .Z(n33727) );
  XOR U33499 ( .A(n33730), .B(n33731), .Z(n33641) );
  NOR U33500 ( .A(n33732), .B(n33733), .Z(n33731) );
  XNOR U33501 ( .A(n33730), .B(n33734), .Z(n33732) );
  XNOR U33502 ( .A(n33533), .B(n33647), .Z(n33649) );
  XNOR U33503 ( .A(n33735), .B(n33736), .Z(n33533) );
  AND U33504 ( .A(n420), .B(n33737), .Z(n33736) );
  XNOR U33505 ( .A(n33738), .B(n33739), .Z(n33737) );
  AND U33506 ( .A(n33539), .B(n33542), .Z(n33647) );
  XOR U33507 ( .A(n33740), .B(n33696), .Z(n33542) );
  XNOR U33508 ( .A(p_input[2048]), .B(p_input[480]), .Z(n33696) );
  XOR U33509 ( .A(n33673), .B(n33672), .Z(n33740) );
  XOR U33510 ( .A(n33741), .B(n33684), .Z(n33672) );
  XOR U33511 ( .A(n33658), .B(n33657), .Z(n33684) );
  XNOR U33512 ( .A(n33742), .B(n33663), .Z(n33657) );
  XOR U33513 ( .A(p_input[2072]), .B(p_input[504]), .Z(n33663) );
  XOR U33514 ( .A(n33654), .B(n33662), .Z(n33742) );
  XOR U33515 ( .A(n33743), .B(n33659), .Z(n33662) );
  XOR U33516 ( .A(p_input[2070]), .B(p_input[502]), .Z(n33659) );
  XNOR U33517 ( .A(p_input[2071]), .B(p_input[503]), .Z(n33743) );
  XNOR U33518 ( .A(n28684), .B(p_input[498]), .Z(n33654) );
  XNOR U33519 ( .A(n33668), .B(n33667), .Z(n33658) );
  XOR U33520 ( .A(n33744), .B(n33664), .Z(n33667) );
  XOR U33521 ( .A(p_input[2067]), .B(p_input[499]), .Z(n33664) );
  XNOR U33522 ( .A(p_input[2068]), .B(p_input[500]), .Z(n33744) );
  XOR U33523 ( .A(p_input[2069]), .B(p_input[501]), .Z(n33668) );
  XNOR U33524 ( .A(n33683), .B(n33669), .Z(n33741) );
  XNOR U33525 ( .A(n28686), .B(p_input[481]), .Z(n33669) );
  XNOR U33526 ( .A(n33745), .B(n33690), .Z(n33683) );
  XNOR U33527 ( .A(n33679), .B(n33678), .Z(n33690) );
  XOR U33528 ( .A(n33746), .B(n33675), .Z(n33678) );
  XNOR U33529 ( .A(n28322), .B(p_input[506]), .Z(n33675) );
  XNOR U33530 ( .A(p_input[2075]), .B(p_input[507]), .Z(n33746) );
  XOR U33531 ( .A(p_input[2076]), .B(p_input[508]), .Z(n33679) );
  XNOR U33532 ( .A(n33689), .B(n33680), .Z(n33745) );
  XNOR U33533 ( .A(n28689), .B(p_input[497]), .Z(n33680) );
  XOR U33534 ( .A(n33747), .B(n33695), .Z(n33689) );
  XNOR U33535 ( .A(p_input[2079]), .B(p_input[511]), .Z(n33695) );
  XOR U33536 ( .A(n33686), .B(n33694), .Z(n33747) );
  XOR U33537 ( .A(n33748), .B(n33691), .Z(n33694) );
  XOR U33538 ( .A(p_input[2077]), .B(p_input[509]), .Z(n33691) );
  XNOR U33539 ( .A(p_input[2078]), .B(p_input[510]), .Z(n33748) );
  XNOR U33540 ( .A(n28326), .B(p_input[505]), .Z(n33686) );
  XNOR U33541 ( .A(n33707), .B(n33706), .Z(n33673) );
  XNOR U33542 ( .A(n33749), .B(n33713), .Z(n33706) );
  XNOR U33543 ( .A(n33702), .B(n33701), .Z(n33713) );
  XOR U33544 ( .A(n33750), .B(n33698), .Z(n33701) );
  XNOR U33545 ( .A(n28694), .B(p_input[491]), .Z(n33698) );
  XNOR U33546 ( .A(p_input[2060]), .B(p_input[492]), .Z(n33750) );
  XOR U33547 ( .A(p_input[2061]), .B(p_input[493]), .Z(n33702) );
  XNOR U33548 ( .A(n33712), .B(n33703), .Z(n33749) );
  XNOR U33549 ( .A(n28330), .B(p_input[482]), .Z(n33703) );
  XOR U33550 ( .A(n33751), .B(n33718), .Z(n33712) );
  XNOR U33551 ( .A(p_input[2064]), .B(p_input[496]), .Z(n33718) );
  XOR U33552 ( .A(n33709), .B(n33717), .Z(n33751) );
  XOR U33553 ( .A(n33752), .B(n33714), .Z(n33717) );
  XOR U33554 ( .A(p_input[2062]), .B(p_input[494]), .Z(n33714) );
  XNOR U33555 ( .A(p_input[2063]), .B(p_input[495]), .Z(n33752) );
  XNOR U33556 ( .A(n28697), .B(p_input[490]), .Z(n33709) );
  XNOR U33557 ( .A(n33724), .B(n33723), .Z(n33707) );
  XNOR U33558 ( .A(n33753), .B(n33729), .Z(n33723) );
  XOR U33559 ( .A(p_input[2057]), .B(p_input[489]), .Z(n33729) );
  XOR U33560 ( .A(n33720), .B(n33728), .Z(n33753) );
  XOR U33561 ( .A(n33754), .B(n33725), .Z(n33728) );
  XOR U33562 ( .A(p_input[2055]), .B(p_input[487]), .Z(n33725) );
  XNOR U33563 ( .A(p_input[2056]), .B(p_input[488]), .Z(n33754) );
  XNOR U33564 ( .A(n28337), .B(p_input[483]), .Z(n33720) );
  XNOR U33565 ( .A(n33734), .B(n33733), .Z(n33724) );
  XOR U33566 ( .A(n33755), .B(n33730), .Z(n33733) );
  XOR U33567 ( .A(p_input[2052]), .B(p_input[484]), .Z(n33730) );
  XNOR U33568 ( .A(p_input[2053]), .B(p_input[485]), .Z(n33755) );
  XOR U33569 ( .A(p_input[2054]), .B(p_input[486]), .Z(n33734) );
  XNOR U33570 ( .A(n33756), .B(n33757), .Z(n33539) );
  AND U33571 ( .A(n420), .B(n33758), .Z(n33757) );
  XNOR U33572 ( .A(n33759), .B(n33760), .Z(n420) );
  AND U33573 ( .A(n33761), .B(n33762), .Z(n33760) );
  XOR U33574 ( .A(n33553), .B(n33759), .Z(n33762) );
  XNOR U33575 ( .A(n33763), .B(n33759), .Z(n33761) );
  XOR U33576 ( .A(n33764), .B(n33765), .Z(n33759) );
  AND U33577 ( .A(n33766), .B(n33767), .Z(n33765) );
  XOR U33578 ( .A(n33568), .B(n33764), .Z(n33767) );
  XOR U33579 ( .A(n33764), .B(n33569), .Z(n33766) );
  XOR U33580 ( .A(n33768), .B(n33769), .Z(n33764) );
  AND U33581 ( .A(n33770), .B(n33771), .Z(n33769) );
  XOR U33582 ( .A(n33596), .B(n33768), .Z(n33771) );
  XOR U33583 ( .A(n33768), .B(n33597), .Z(n33770) );
  XOR U33584 ( .A(n33772), .B(n33773), .Z(n33768) );
  AND U33585 ( .A(n33774), .B(n33775), .Z(n33773) );
  XOR U33586 ( .A(n33645), .B(n33772), .Z(n33775) );
  XOR U33587 ( .A(n33772), .B(n33646), .Z(n33774) );
  XOR U33588 ( .A(n33776), .B(n33777), .Z(n33772) );
  AND U33589 ( .A(n33778), .B(n33779), .Z(n33777) );
  XOR U33590 ( .A(n33776), .B(n33738), .Z(n33779) );
  XNOR U33591 ( .A(n33780), .B(n33781), .Z(n33489) );
  AND U33592 ( .A(n424), .B(n33782), .Z(n33781) );
  XNOR U33593 ( .A(n33783), .B(n33784), .Z(n424) );
  AND U33594 ( .A(n33785), .B(n33786), .Z(n33784) );
  XOR U33595 ( .A(n33783), .B(n33499), .Z(n33786) );
  XNOR U33596 ( .A(n33783), .B(n33449), .Z(n33785) );
  XOR U33597 ( .A(n33787), .B(n33788), .Z(n33783) );
  AND U33598 ( .A(n33789), .B(n33790), .Z(n33788) );
  XNOR U33599 ( .A(n33509), .B(n33787), .Z(n33790) );
  XOR U33600 ( .A(n33787), .B(n33459), .Z(n33789) );
  XOR U33601 ( .A(n33791), .B(n33792), .Z(n33787) );
  AND U33602 ( .A(n33793), .B(n33794), .Z(n33792) );
  XNOR U33603 ( .A(n33519), .B(n33791), .Z(n33794) );
  XOR U33604 ( .A(n33791), .B(n33468), .Z(n33793) );
  XOR U33605 ( .A(n33795), .B(n33796), .Z(n33791) );
  AND U33606 ( .A(n33797), .B(n33798), .Z(n33796) );
  XOR U33607 ( .A(n33795), .B(n33476), .Z(n33797) );
  XOR U33608 ( .A(n33799), .B(n33800), .Z(n33440) );
  AND U33609 ( .A(n428), .B(n33782), .Z(n33800) );
  XNOR U33610 ( .A(n33780), .B(n33799), .Z(n33782) );
  XNOR U33611 ( .A(n33801), .B(n33802), .Z(n428) );
  AND U33612 ( .A(n33803), .B(n33804), .Z(n33802) );
  XNOR U33613 ( .A(n33805), .B(n33801), .Z(n33804) );
  IV U33614 ( .A(n33499), .Z(n33805) );
  XOR U33615 ( .A(n33763), .B(n33806), .Z(n33499) );
  AND U33616 ( .A(n431), .B(n33807), .Z(n33806) );
  XOR U33617 ( .A(n33552), .B(n33549), .Z(n33807) );
  IV U33618 ( .A(n33763), .Z(n33552) );
  XNOR U33619 ( .A(n33449), .B(n33801), .Z(n33803) );
  XOR U33620 ( .A(n33808), .B(n33809), .Z(n33449) );
  AND U33621 ( .A(n447), .B(n33810), .Z(n33809) );
  XOR U33622 ( .A(n33811), .B(n33812), .Z(n33801) );
  AND U33623 ( .A(n33813), .B(n33814), .Z(n33812) );
  XNOR U33624 ( .A(n33811), .B(n33509), .Z(n33814) );
  XOR U33625 ( .A(n33569), .B(n33815), .Z(n33509) );
  AND U33626 ( .A(n431), .B(n33816), .Z(n33815) );
  XOR U33627 ( .A(n33565), .B(n33569), .Z(n33816) );
  XNOR U33628 ( .A(n33817), .B(n33811), .Z(n33813) );
  IV U33629 ( .A(n33459), .Z(n33817) );
  XOR U33630 ( .A(n33818), .B(n33819), .Z(n33459) );
  AND U33631 ( .A(n447), .B(n33820), .Z(n33819) );
  XOR U33632 ( .A(n33821), .B(n33822), .Z(n33811) );
  AND U33633 ( .A(n33823), .B(n33824), .Z(n33822) );
  XNOR U33634 ( .A(n33821), .B(n33519), .Z(n33824) );
  XOR U33635 ( .A(n33597), .B(n33825), .Z(n33519) );
  AND U33636 ( .A(n431), .B(n33826), .Z(n33825) );
  XOR U33637 ( .A(n33593), .B(n33597), .Z(n33826) );
  XOR U33638 ( .A(n33468), .B(n33821), .Z(n33823) );
  XOR U33639 ( .A(n33827), .B(n33828), .Z(n33468) );
  AND U33640 ( .A(n447), .B(n33829), .Z(n33828) );
  XOR U33641 ( .A(n33795), .B(n33830), .Z(n33821) );
  AND U33642 ( .A(n33831), .B(n33798), .Z(n33830) );
  XNOR U33643 ( .A(n33529), .B(n33795), .Z(n33798) );
  XOR U33644 ( .A(n33646), .B(n33832), .Z(n33529) );
  AND U33645 ( .A(n431), .B(n33833), .Z(n33832) );
  XOR U33646 ( .A(n33642), .B(n33646), .Z(n33833) );
  XNOR U33647 ( .A(n33834), .B(n33795), .Z(n33831) );
  IV U33648 ( .A(n33476), .Z(n33834) );
  XOR U33649 ( .A(n33835), .B(n33836), .Z(n33476) );
  AND U33650 ( .A(n447), .B(n33837), .Z(n33836) );
  XOR U33651 ( .A(n33838), .B(n33839), .Z(n33795) );
  AND U33652 ( .A(n33840), .B(n33841), .Z(n33839) );
  XNOR U33653 ( .A(n33838), .B(n33537), .Z(n33841) );
  XOR U33654 ( .A(n33739), .B(n33842), .Z(n33537) );
  AND U33655 ( .A(n431), .B(n33843), .Z(n33842) );
  XOR U33656 ( .A(n33735), .B(n33739), .Z(n33843) );
  XNOR U33657 ( .A(n33844), .B(n33838), .Z(n33840) );
  IV U33658 ( .A(n33486), .Z(n33844) );
  XOR U33659 ( .A(n33845), .B(n33846), .Z(n33486) );
  AND U33660 ( .A(n447), .B(n33847), .Z(n33846) );
  AND U33661 ( .A(n33799), .B(n33780), .Z(n33838) );
  XNOR U33662 ( .A(n33848), .B(n33849), .Z(n33780) );
  AND U33663 ( .A(n431), .B(n33758), .Z(n33849) );
  XNOR U33664 ( .A(n33756), .B(n33848), .Z(n33758) );
  XNOR U33665 ( .A(n33850), .B(n33851), .Z(n431) );
  AND U33666 ( .A(n33852), .B(n33853), .Z(n33851) );
  XNOR U33667 ( .A(n33850), .B(n33549), .Z(n33853) );
  IV U33668 ( .A(n33553), .Z(n33549) );
  XOR U33669 ( .A(n33854), .B(n33855), .Z(n33553) );
  AND U33670 ( .A(n435), .B(n33856), .Z(n33855) );
  XOR U33671 ( .A(n33857), .B(n33854), .Z(n33856) );
  XNOR U33672 ( .A(n33850), .B(n33763), .Z(n33852) );
  XOR U33673 ( .A(n33858), .B(n33859), .Z(n33763) );
  AND U33674 ( .A(n443), .B(n33810), .Z(n33859) );
  XOR U33675 ( .A(n33808), .B(n33858), .Z(n33810) );
  XOR U33676 ( .A(n33860), .B(n33861), .Z(n33850) );
  AND U33677 ( .A(n33862), .B(n33863), .Z(n33861) );
  XNOR U33678 ( .A(n33860), .B(n33565), .Z(n33863) );
  IV U33679 ( .A(n33568), .Z(n33565) );
  XOR U33680 ( .A(n33864), .B(n33865), .Z(n33568) );
  AND U33681 ( .A(n435), .B(n33866), .Z(n33865) );
  XOR U33682 ( .A(n33867), .B(n33864), .Z(n33866) );
  XOR U33683 ( .A(n33569), .B(n33860), .Z(n33862) );
  XOR U33684 ( .A(n33868), .B(n33869), .Z(n33569) );
  AND U33685 ( .A(n443), .B(n33820), .Z(n33869) );
  XOR U33686 ( .A(n33868), .B(n33818), .Z(n33820) );
  XOR U33687 ( .A(n33870), .B(n33871), .Z(n33860) );
  AND U33688 ( .A(n33872), .B(n33873), .Z(n33871) );
  XNOR U33689 ( .A(n33870), .B(n33593), .Z(n33873) );
  IV U33690 ( .A(n33596), .Z(n33593) );
  XOR U33691 ( .A(n33874), .B(n33875), .Z(n33596) );
  AND U33692 ( .A(n435), .B(n33876), .Z(n33875) );
  XNOR U33693 ( .A(n33877), .B(n33874), .Z(n33876) );
  XOR U33694 ( .A(n33597), .B(n33870), .Z(n33872) );
  XOR U33695 ( .A(n33878), .B(n33879), .Z(n33597) );
  AND U33696 ( .A(n443), .B(n33829), .Z(n33879) );
  XOR U33697 ( .A(n33878), .B(n33827), .Z(n33829) );
  XOR U33698 ( .A(n33880), .B(n33881), .Z(n33870) );
  AND U33699 ( .A(n33882), .B(n33883), .Z(n33881) );
  XNOR U33700 ( .A(n33880), .B(n33642), .Z(n33883) );
  IV U33701 ( .A(n33645), .Z(n33642) );
  XOR U33702 ( .A(n33884), .B(n33885), .Z(n33645) );
  AND U33703 ( .A(n435), .B(n33886), .Z(n33885) );
  XOR U33704 ( .A(n33887), .B(n33884), .Z(n33886) );
  XOR U33705 ( .A(n33646), .B(n33880), .Z(n33882) );
  XOR U33706 ( .A(n33888), .B(n33889), .Z(n33646) );
  AND U33707 ( .A(n443), .B(n33837), .Z(n33889) );
  XOR U33708 ( .A(n33888), .B(n33835), .Z(n33837) );
  XOR U33709 ( .A(n33776), .B(n33890), .Z(n33880) );
  AND U33710 ( .A(n33778), .B(n33891), .Z(n33890) );
  XNOR U33711 ( .A(n33776), .B(n33735), .Z(n33891) );
  IV U33712 ( .A(n33738), .Z(n33735) );
  XOR U33713 ( .A(n33892), .B(n33893), .Z(n33738) );
  AND U33714 ( .A(n435), .B(n33894), .Z(n33893) );
  XNOR U33715 ( .A(n33895), .B(n33892), .Z(n33894) );
  XOR U33716 ( .A(n33739), .B(n33776), .Z(n33778) );
  XOR U33717 ( .A(n33896), .B(n33897), .Z(n33739) );
  AND U33718 ( .A(n443), .B(n33847), .Z(n33897) );
  XOR U33719 ( .A(n33896), .B(n33845), .Z(n33847) );
  AND U33720 ( .A(n33848), .B(n33756), .Z(n33776) );
  XNOR U33721 ( .A(n33898), .B(n33899), .Z(n33756) );
  AND U33722 ( .A(n435), .B(n33900), .Z(n33899) );
  XNOR U33723 ( .A(n33901), .B(n33898), .Z(n33900) );
  XNOR U33724 ( .A(n33902), .B(n33903), .Z(n435) );
  AND U33725 ( .A(n33904), .B(n33905), .Z(n33903) );
  XOR U33726 ( .A(n33857), .B(n33902), .Z(n33905) );
  AND U33727 ( .A(n33906), .B(n33907), .Z(n33857) );
  XNOR U33728 ( .A(n33854), .B(n33902), .Z(n33904) );
  XNOR U33729 ( .A(n33908), .B(n33909), .Z(n33854) );
  AND U33730 ( .A(n439), .B(n33910), .Z(n33909) );
  XNOR U33731 ( .A(n33911), .B(n33912), .Z(n33910) );
  XOR U33732 ( .A(n33913), .B(n33914), .Z(n33902) );
  AND U33733 ( .A(n33915), .B(n33916), .Z(n33914) );
  XNOR U33734 ( .A(n33913), .B(n33906), .Z(n33916) );
  IV U33735 ( .A(n33867), .Z(n33906) );
  XOR U33736 ( .A(n33917), .B(n33918), .Z(n33867) );
  XOR U33737 ( .A(n33919), .B(n33907), .Z(n33918) );
  AND U33738 ( .A(n33877), .B(n33920), .Z(n33907) );
  AND U33739 ( .A(n33921), .B(n33922), .Z(n33919) );
  XOR U33740 ( .A(n33923), .B(n33917), .Z(n33921) );
  XNOR U33741 ( .A(n33864), .B(n33913), .Z(n33915) );
  XNOR U33742 ( .A(n33924), .B(n33925), .Z(n33864) );
  AND U33743 ( .A(n439), .B(n33926), .Z(n33925) );
  XNOR U33744 ( .A(n33927), .B(n33928), .Z(n33926) );
  XOR U33745 ( .A(n33929), .B(n33930), .Z(n33913) );
  AND U33746 ( .A(n33931), .B(n33932), .Z(n33930) );
  XNOR U33747 ( .A(n33929), .B(n33877), .Z(n33932) );
  XOR U33748 ( .A(n33933), .B(n33922), .Z(n33877) );
  XNOR U33749 ( .A(n33934), .B(n33917), .Z(n33922) );
  XOR U33750 ( .A(n33935), .B(n33936), .Z(n33917) );
  AND U33751 ( .A(n33937), .B(n33938), .Z(n33936) );
  XOR U33752 ( .A(n33939), .B(n33935), .Z(n33937) );
  XNOR U33753 ( .A(n33940), .B(n33941), .Z(n33934) );
  AND U33754 ( .A(n33942), .B(n33943), .Z(n33941) );
  XOR U33755 ( .A(n33940), .B(n33944), .Z(n33942) );
  XNOR U33756 ( .A(n33923), .B(n33920), .Z(n33933) );
  AND U33757 ( .A(n33945), .B(n33946), .Z(n33920) );
  XOR U33758 ( .A(n33947), .B(n33948), .Z(n33923) );
  AND U33759 ( .A(n33949), .B(n33950), .Z(n33948) );
  XOR U33760 ( .A(n33947), .B(n33951), .Z(n33949) );
  XNOR U33761 ( .A(n33874), .B(n33929), .Z(n33931) );
  XNOR U33762 ( .A(n33952), .B(n33953), .Z(n33874) );
  AND U33763 ( .A(n439), .B(n33954), .Z(n33953) );
  XNOR U33764 ( .A(n33955), .B(n33956), .Z(n33954) );
  XOR U33765 ( .A(n33957), .B(n33958), .Z(n33929) );
  AND U33766 ( .A(n33959), .B(n33960), .Z(n33958) );
  XNOR U33767 ( .A(n33957), .B(n33945), .Z(n33960) );
  IV U33768 ( .A(n33887), .Z(n33945) );
  XNOR U33769 ( .A(n33961), .B(n33938), .Z(n33887) );
  XNOR U33770 ( .A(n33962), .B(n33944), .Z(n33938) );
  XOR U33771 ( .A(n33963), .B(n33964), .Z(n33944) );
  AND U33772 ( .A(n33965), .B(n33966), .Z(n33964) );
  XOR U33773 ( .A(n33963), .B(n33967), .Z(n33965) );
  XNOR U33774 ( .A(n33943), .B(n33935), .Z(n33962) );
  XOR U33775 ( .A(n33968), .B(n33969), .Z(n33935) );
  AND U33776 ( .A(n33970), .B(n33971), .Z(n33969) );
  XNOR U33777 ( .A(n33972), .B(n33968), .Z(n33970) );
  XNOR U33778 ( .A(n33973), .B(n33940), .Z(n33943) );
  XOR U33779 ( .A(n33974), .B(n33975), .Z(n33940) );
  AND U33780 ( .A(n33976), .B(n33977), .Z(n33975) );
  XOR U33781 ( .A(n33974), .B(n33978), .Z(n33976) );
  XNOR U33782 ( .A(n33979), .B(n33980), .Z(n33973) );
  AND U33783 ( .A(n33981), .B(n33982), .Z(n33980) );
  XNOR U33784 ( .A(n33979), .B(n33983), .Z(n33981) );
  XNOR U33785 ( .A(n33939), .B(n33946), .Z(n33961) );
  AND U33786 ( .A(n33895), .B(n33984), .Z(n33946) );
  XOR U33787 ( .A(n33951), .B(n33950), .Z(n33939) );
  XNOR U33788 ( .A(n33985), .B(n33947), .Z(n33950) );
  XOR U33789 ( .A(n33986), .B(n33987), .Z(n33947) );
  AND U33790 ( .A(n33988), .B(n33989), .Z(n33987) );
  XOR U33791 ( .A(n33986), .B(n33990), .Z(n33988) );
  XNOR U33792 ( .A(n33991), .B(n33992), .Z(n33985) );
  AND U33793 ( .A(n33993), .B(n33994), .Z(n33992) );
  XOR U33794 ( .A(n33991), .B(n33995), .Z(n33993) );
  XOR U33795 ( .A(n33996), .B(n33997), .Z(n33951) );
  AND U33796 ( .A(n33998), .B(n33999), .Z(n33997) );
  XOR U33797 ( .A(n33996), .B(n34000), .Z(n33998) );
  XNOR U33798 ( .A(n33884), .B(n33957), .Z(n33959) );
  XNOR U33799 ( .A(n34001), .B(n34002), .Z(n33884) );
  AND U33800 ( .A(n439), .B(n34003), .Z(n34002) );
  XNOR U33801 ( .A(n34004), .B(n34005), .Z(n34003) );
  XOR U33802 ( .A(n34006), .B(n34007), .Z(n33957) );
  AND U33803 ( .A(n34008), .B(n34009), .Z(n34007) );
  XNOR U33804 ( .A(n34006), .B(n33895), .Z(n34009) );
  XOR U33805 ( .A(n34010), .B(n33971), .Z(n33895) );
  XNOR U33806 ( .A(n34011), .B(n33978), .Z(n33971) );
  XOR U33807 ( .A(n33967), .B(n33966), .Z(n33978) );
  XNOR U33808 ( .A(n34012), .B(n33963), .Z(n33966) );
  XOR U33809 ( .A(n34013), .B(n34014), .Z(n33963) );
  AND U33810 ( .A(n34015), .B(n34016), .Z(n34014) );
  XOR U33811 ( .A(n34013), .B(n34017), .Z(n34015) );
  XNOR U33812 ( .A(n34018), .B(n34019), .Z(n34012) );
  NOR U33813 ( .A(n34020), .B(n34021), .Z(n34019) );
  XNOR U33814 ( .A(n34018), .B(n34022), .Z(n34020) );
  XOR U33815 ( .A(n34023), .B(n34024), .Z(n33967) );
  NOR U33816 ( .A(n34025), .B(n34026), .Z(n34024) );
  XNOR U33817 ( .A(n34023), .B(n34027), .Z(n34025) );
  XNOR U33818 ( .A(n33977), .B(n33968), .Z(n34011) );
  XOR U33819 ( .A(n34028), .B(n34029), .Z(n33968) );
  NOR U33820 ( .A(n34030), .B(n34031), .Z(n34029) );
  XNOR U33821 ( .A(n34028), .B(n34032), .Z(n34030) );
  XOR U33822 ( .A(n34033), .B(n33983), .Z(n33977) );
  XNOR U33823 ( .A(n34034), .B(n34035), .Z(n33983) );
  NOR U33824 ( .A(n34036), .B(n34037), .Z(n34035) );
  XNOR U33825 ( .A(n34034), .B(n34038), .Z(n34036) );
  XNOR U33826 ( .A(n33982), .B(n33974), .Z(n34033) );
  XOR U33827 ( .A(n34039), .B(n34040), .Z(n33974) );
  AND U33828 ( .A(n34041), .B(n34042), .Z(n34040) );
  XOR U33829 ( .A(n34039), .B(n34043), .Z(n34041) );
  XNOR U33830 ( .A(n34044), .B(n33979), .Z(n33982) );
  XOR U33831 ( .A(n34045), .B(n34046), .Z(n33979) );
  AND U33832 ( .A(n34047), .B(n34048), .Z(n34046) );
  XOR U33833 ( .A(n34045), .B(n34049), .Z(n34047) );
  XNOR U33834 ( .A(n34050), .B(n34051), .Z(n34044) );
  NOR U33835 ( .A(n34052), .B(n34053), .Z(n34051) );
  XOR U33836 ( .A(n34050), .B(n34054), .Z(n34052) );
  XOR U33837 ( .A(n33972), .B(n33984), .Z(n34010) );
  NOR U33838 ( .A(n33901), .B(n34055), .Z(n33984) );
  XNOR U33839 ( .A(n33990), .B(n33989), .Z(n33972) );
  XNOR U33840 ( .A(n34056), .B(n33995), .Z(n33989) );
  XOR U33841 ( .A(n34057), .B(n34058), .Z(n33995) );
  NOR U33842 ( .A(n34059), .B(n34060), .Z(n34058) );
  XNOR U33843 ( .A(n34057), .B(n34061), .Z(n34059) );
  XNOR U33844 ( .A(n33994), .B(n33986), .Z(n34056) );
  XOR U33845 ( .A(n34062), .B(n34063), .Z(n33986) );
  AND U33846 ( .A(n34064), .B(n34065), .Z(n34063) );
  XNOR U33847 ( .A(n34062), .B(n34066), .Z(n34064) );
  XNOR U33848 ( .A(n34067), .B(n33991), .Z(n33994) );
  XOR U33849 ( .A(n34068), .B(n34069), .Z(n33991) );
  AND U33850 ( .A(n34070), .B(n34071), .Z(n34069) );
  XOR U33851 ( .A(n34068), .B(n34072), .Z(n34070) );
  XNOR U33852 ( .A(n34073), .B(n34074), .Z(n34067) );
  NOR U33853 ( .A(n34075), .B(n34076), .Z(n34074) );
  XOR U33854 ( .A(n34073), .B(n34077), .Z(n34075) );
  XOR U33855 ( .A(n34000), .B(n33999), .Z(n33990) );
  XNOR U33856 ( .A(n34078), .B(n33996), .Z(n33999) );
  XOR U33857 ( .A(n34079), .B(n34080), .Z(n33996) );
  AND U33858 ( .A(n34081), .B(n34082), .Z(n34080) );
  XOR U33859 ( .A(n34079), .B(n34083), .Z(n34081) );
  XNOR U33860 ( .A(n34084), .B(n34085), .Z(n34078) );
  NOR U33861 ( .A(n34086), .B(n34087), .Z(n34085) );
  XNOR U33862 ( .A(n34084), .B(n34088), .Z(n34086) );
  XOR U33863 ( .A(n34089), .B(n34090), .Z(n34000) );
  NOR U33864 ( .A(n34091), .B(n34092), .Z(n34090) );
  XNOR U33865 ( .A(n34089), .B(n34093), .Z(n34091) );
  XNOR U33866 ( .A(n33892), .B(n34006), .Z(n34008) );
  XNOR U33867 ( .A(n34094), .B(n34095), .Z(n33892) );
  AND U33868 ( .A(n439), .B(n34096), .Z(n34095) );
  XNOR U33869 ( .A(n34097), .B(n34098), .Z(n34096) );
  AND U33870 ( .A(n33898), .B(n33901), .Z(n34006) );
  XOR U33871 ( .A(n34099), .B(n34055), .Z(n33901) );
  XNOR U33872 ( .A(p_input[2048]), .B(p_input[512]), .Z(n34055) );
  XOR U33873 ( .A(n34032), .B(n34031), .Z(n34099) );
  XOR U33874 ( .A(n34100), .B(n34043), .Z(n34031) );
  XOR U33875 ( .A(n34017), .B(n34016), .Z(n34043) );
  XNOR U33876 ( .A(n34101), .B(n34022), .Z(n34016) );
  XOR U33877 ( .A(p_input[2072]), .B(p_input[536]), .Z(n34022) );
  XOR U33878 ( .A(n34013), .B(n34021), .Z(n34101) );
  XOR U33879 ( .A(n34102), .B(n34018), .Z(n34021) );
  XOR U33880 ( .A(p_input[2070]), .B(p_input[534]), .Z(n34018) );
  XNOR U33881 ( .A(p_input[2071]), .B(p_input[535]), .Z(n34102) );
  XNOR U33882 ( .A(n28684), .B(p_input[530]), .Z(n34013) );
  XNOR U33883 ( .A(n34027), .B(n34026), .Z(n34017) );
  XOR U33884 ( .A(n34103), .B(n34023), .Z(n34026) );
  XOR U33885 ( .A(p_input[2067]), .B(p_input[531]), .Z(n34023) );
  XNOR U33886 ( .A(p_input[2068]), .B(p_input[532]), .Z(n34103) );
  XOR U33887 ( .A(p_input[2069]), .B(p_input[533]), .Z(n34027) );
  XNOR U33888 ( .A(n34042), .B(n34028), .Z(n34100) );
  XNOR U33889 ( .A(n28686), .B(p_input[513]), .Z(n34028) );
  XNOR U33890 ( .A(n34104), .B(n34049), .Z(n34042) );
  XNOR U33891 ( .A(n34038), .B(n34037), .Z(n34049) );
  XOR U33892 ( .A(n34105), .B(n34034), .Z(n34037) );
  XNOR U33893 ( .A(n28322), .B(p_input[538]), .Z(n34034) );
  XNOR U33894 ( .A(p_input[2075]), .B(p_input[539]), .Z(n34105) );
  XOR U33895 ( .A(p_input[2076]), .B(p_input[540]), .Z(n34038) );
  XNOR U33896 ( .A(n34048), .B(n34039), .Z(n34104) );
  XNOR U33897 ( .A(n28689), .B(p_input[529]), .Z(n34039) );
  XOR U33898 ( .A(n34106), .B(n34054), .Z(n34048) );
  XNOR U33899 ( .A(p_input[2079]), .B(p_input[543]), .Z(n34054) );
  XOR U33900 ( .A(n34045), .B(n34053), .Z(n34106) );
  XOR U33901 ( .A(n34107), .B(n34050), .Z(n34053) );
  XOR U33902 ( .A(p_input[2077]), .B(p_input[541]), .Z(n34050) );
  XNOR U33903 ( .A(p_input[2078]), .B(p_input[542]), .Z(n34107) );
  XNOR U33904 ( .A(n28326), .B(p_input[537]), .Z(n34045) );
  XNOR U33905 ( .A(n34066), .B(n34065), .Z(n34032) );
  XNOR U33906 ( .A(n34108), .B(n34072), .Z(n34065) );
  XNOR U33907 ( .A(n34061), .B(n34060), .Z(n34072) );
  XOR U33908 ( .A(n34109), .B(n34057), .Z(n34060) );
  XNOR U33909 ( .A(n28694), .B(p_input[523]), .Z(n34057) );
  XNOR U33910 ( .A(p_input[2060]), .B(p_input[524]), .Z(n34109) );
  XOR U33911 ( .A(p_input[2061]), .B(p_input[525]), .Z(n34061) );
  XNOR U33912 ( .A(n34071), .B(n34062), .Z(n34108) );
  XNOR U33913 ( .A(n28330), .B(p_input[514]), .Z(n34062) );
  XOR U33914 ( .A(n34110), .B(n34077), .Z(n34071) );
  XNOR U33915 ( .A(p_input[2064]), .B(p_input[528]), .Z(n34077) );
  XOR U33916 ( .A(n34068), .B(n34076), .Z(n34110) );
  XOR U33917 ( .A(n34111), .B(n34073), .Z(n34076) );
  XOR U33918 ( .A(p_input[2062]), .B(p_input[526]), .Z(n34073) );
  XNOR U33919 ( .A(p_input[2063]), .B(p_input[527]), .Z(n34111) );
  XNOR U33920 ( .A(n28697), .B(p_input[522]), .Z(n34068) );
  XNOR U33921 ( .A(n34083), .B(n34082), .Z(n34066) );
  XNOR U33922 ( .A(n34112), .B(n34088), .Z(n34082) );
  XOR U33923 ( .A(p_input[2057]), .B(p_input[521]), .Z(n34088) );
  XOR U33924 ( .A(n34079), .B(n34087), .Z(n34112) );
  XOR U33925 ( .A(n34113), .B(n34084), .Z(n34087) );
  XOR U33926 ( .A(p_input[2055]), .B(p_input[519]), .Z(n34084) );
  XNOR U33927 ( .A(p_input[2056]), .B(p_input[520]), .Z(n34113) );
  XNOR U33928 ( .A(n28337), .B(p_input[515]), .Z(n34079) );
  XNOR U33929 ( .A(n34093), .B(n34092), .Z(n34083) );
  XOR U33930 ( .A(n34114), .B(n34089), .Z(n34092) );
  XOR U33931 ( .A(p_input[2052]), .B(p_input[516]), .Z(n34089) );
  XNOR U33932 ( .A(p_input[2053]), .B(p_input[517]), .Z(n34114) );
  XOR U33933 ( .A(p_input[2054]), .B(p_input[518]), .Z(n34093) );
  XNOR U33934 ( .A(n34115), .B(n34116), .Z(n33898) );
  AND U33935 ( .A(n439), .B(n34117), .Z(n34116) );
  XNOR U33936 ( .A(n34118), .B(n34119), .Z(n439) );
  AND U33937 ( .A(n34120), .B(n34121), .Z(n34119) );
  XOR U33938 ( .A(n33912), .B(n34118), .Z(n34121) );
  XNOR U33939 ( .A(n34122), .B(n34118), .Z(n34120) );
  XOR U33940 ( .A(n34123), .B(n34124), .Z(n34118) );
  AND U33941 ( .A(n34125), .B(n34126), .Z(n34124) );
  XOR U33942 ( .A(n33927), .B(n34123), .Z(n34126) );
  XOR U33943 ( .A(n34123), .B(n33928), .Z(n34125) );
  XOR U33944 ( .A(n34127), .B(n34128), .Z(n34123) );
  AND U33945 ( .A(n34129), .B(n34130), .Z(n34128) );
  XOR U33946 ( .A(n33955), .B(n34127), .Z(n34130) );
  XOR U33947 ( .A(n34127), .B(n33956), .Z(n34129) );
  XOR U33948 ( .A(n34131), .B(n34132), .Z(n34127) );
  AND U33949 ( .A(n34133), .B(n34134), .Z(n34132) );
  XOR U33950 ( .A(n34004), .B(n34131), .Z(n34134) );
  XOR U33951 ( .A(n34131), .B(n34005), .Z(n34133) );
  XOR U33952 ( .A(n34135), .B(n34136), .Z(n34131) );
  AND U33953 ( .A(n34137), .B(n34138), .Z(n34136) );
  XOR U33954 ( .A(n34135), .B(n34097), .Z(n34138) );
  XNOR U33955 ( .A(n34139), .B(n34140), .Z(n33848) );
  AND U33956 ( .A(n443), .B(n34141), .Z(n34140) );
  XNOR U33957 ( .A(n34142), .B(n34143), .Z(n443) );
  AND U33958 ( .A(n34144), .B(n34145), .Z(n34143) );
  XOR U33959 ( .A(n34142), .B(n33858), .Z(n34145) );
  XNOR U33960 ( .A(n34142), .B(n33808), .Z(n34144) );
  XOR U33961 ( .A(n34146), .B(n34147), .Z(n34142) );
  AND U33962 ( .A(n34148), .B(n34149), .Z(n34147) );
  XNOR U33963 ( .A(n33868), .B(n34146), .Z(n34149) );
  XOR U33964 ( .A(n34146), .B(n33818), .Z(n34148) );
  XOR U33965 ( .A(n34150), .B(n34151), .Z(n34146) );
  AND U33966 ( .A(n34152), .B(n34153), .Z(n34151) );
  XNOR U33967 ( .A(n33878), .B(n34150), .Z(n34153) );
  XOR U33968 ( .A(n34150), .B(n33827), .Z(n34152) );
  XOR U33969 ( .A(n34154), .B(n34155), .Z(n34150) );
  AND U33970 ( .A(n34156), .B(n34157), .Z(n34155) );
  XOR U33971 ( .A(n34154), .B(n33835), .Z(n34156) );
  XOR U33972 ( .A(n34158), .B(n34159), .Z(n33799) );
  AND U33973 ( .A(n447), .B(n34141), .Z(n34159) );
  XNOR U33974 ( .A(n34139), .B(n34158), .Z(n34141) );
  XNOR U33975 ( .A(n34160), .B(n34161), .Z(n447) );
  AND U33976 ( .A(n34162), .B(n34163), .Z(n34161) );
  XNOR U33977 ( .A(n34164), .B(n34160), .Z(n34163) );
  IV U33978 ( .A(n33858), .Z(n34164) );
  XOR U33979 ( .A(n34122), .B(n34165), .Z(n33858) );
  AND U33980 ( .A(n450), .B(n34166), .Z(n34165) );
  XOR U33981 ( .A(n33911), .B(n33908), .Z(n34166) );
  IV U33982 ( .A(n34122), .Z(n33911) );
  XNOR U33983 ( .A(n33808), .B(n34160), .Z(n34162) );
  XOR U33984 ( .A(n34167), .B(n34168), .Z(n33808) );
  AND U33985 ( .A(n466), .B(n34169), .Z(n34168) );
  XOR U33986 ( .A(n34170), .B(n34171), .Z(n34160) );
  AND U33987 ( .A(n34172), .B(n34173), .Z(n34171) );
  XNOR U33988 ( .A(n34170), .B(n33868), .Z(n34173) );
  XOR U33989 ( .A(n33928), .B(n34174), .Z(n33868) );
  AND U33990 ( .A(n450), .B(n34175), .Z(n34174) );
  XOR U33991 ( .A(n33924), .B(n33928), .Z(n34175) );
  XNOR U33992 ( .A(n34176), .B(n34170), .Z(n34172) );
  IV U33993 ( .A(n33818), .Z(n34176) );
  XOR U33994 ( .A(n34177), .B(n34178), .Z(n33818) );
  AND U33995 ( .A(n466), .B(n34179), .Z(n34178) );
  XOR U33996 ( .A(n34180), .B(n34181), .Z(n34170) );
  AND U33997 ( .A(n34182), .B(n34183), .Z(n34181) );
  XNOR U33998 ( .A(n34180), .B(n33878), .Z(n34183) );
  XOR U33999 ( .A(n33956), .B(n34184), .Z(n33878) );
  AND U34000 ( .A(n450), .B(n34185), .Z(n34184) );
  XOR U34001 ( .A(n33952), .B(n33956), .Z(n34185) );
  XOR U34002 ( .A(n33827), .B(n34180), .Z(n34182) );
  XOR U34003 ( .A(n34186), .B(n34187), .Z(n33827) );
  AND U34004 ( .A(n466), .B(n34188), .Z(n34187) );
  XOR U34005 ( .A(n34154), .B(n34189), .Z(n34180) );
  AND U34006 ( .A(n34190), .B(n34157), .Z(n34189) );
  XNOR U34007 ( .A(n33888), .B(n34154), .Z(n34157) );
  XOR U34008 ( .A(n34005), .B(n34191), .Z(n33888) );
  AND U34009 ( .A(n450), .B(n34192), .Z(n34191) );
  XOR U34010 ( .A(n34001), .B(n34005), .Z(n34192) );
  XNOR U34011 ( .A(n34193), .B(n34154), .Z(n34190) );
  IV U34012 ( .A(n33835), .Z(n34193) );
  XOR U34013 ( .A(n34194), .B(n34195), .Z(n33835) );
  AND U34014 ( .A(n466), .B(n34196), .Z(n34195) );
  XOR U34015 ( .A(n34197), .B(n34198), .Z(n34154) );
  AND U34016 ( .A(n34199), .B(n34200), .Z(n34198) );
  XNOR U34017 ( .A(n34197), .B(n33896), .Z(n34200) );
  XOR U34018 ( .A(n34098), .B(n34201), .Z(n33896) );
  AND U34019 ( .A(n450), .B(n34202), .Z(n34201) );
  XOR U34020 ( .A(n34094), .B(n34098), .Z(n34202) );
  XNOR U34021 ( .A(n34203), .B(n34197), .Z(n34199) );
  IV U34022 ( .A(n33845), .Z(n34203) );
  XOR U34023 ( .A(n34204), .B(n34205), .Z(n33845) );
  AND U34024 ( .A(n466), .B(n34206), .Z(n34205) );
  AND U34025 ( .A(n34158), .B(n34139), .Z(n34197) );
  XNOR U34026 ( .A(n34207), .B(n34208), .Z(n34139) );
  AND U34027 ( .A(n450), .B(n34117), .Z(n34208) );
  XNOR U34028 ( .A(n34115), .B(n34207), .Z(n34117) );
  XNOR U34029 ( .A(n34209), .B(n34210), .Z(n450) );
  AND U34030 ( .A(n34211), .B(n34212), .Z(n34210) );
  XNOR U34031 ( .A(n34209), .B(n33908), .Z(n34212) );
  IV U34032 ( .A(n33912), .Z(n33908) );
  XOR U34033 ( .A(n34213), .B(n34214), .Z(n33912) );
  AND U34034 ( .A(n454), .B(n34215), .Z(n34214) );
  XOR U34035 ( .A(n34216), .B(n34213), .Z(n34215) );
  XNOR U34036 ( .A(n34209), .B(n34122), .Z(n34211) );
  XOR U34037 ( .A(n34217), .B(n34218), .Z(n34122) );
  AND U34038 ( .A(n462), .B(n34169), .Z(n34218) );
  XOR U34039 ( .A(n34167), .B(n34217), .Z(n34169) );
  XOR U34040 ( .A(n34219), .B(n34220), .Z(n34209) );
  AND U34041 ( .A(n34221), .B(n34222), .Z(n34220) );
  XNOR U34042 ( .A(n34219), .B(n33924), .Z(n34222) );
  IV U34043 ( .A(n33927), .Z(n33924) );
  XOR U34044 ( .A(n34223), .B(n34224), .Z(n33927) );
  AND U34045 ( .A(n454), .B(n34225), .Z(n34224) );
  XOR U34046 ( .A(n34226), .B(n34223), .Z(n34225) );
  XOR U34047 ( .A(n33928), .B(n34219), .Z(n34221) );
  XOR U34048 ( .A(n34227), .B(n34228), .Z(n33928) );
  AND U34049 ( .A(n462), .B(n34179), .Z(n34228) );
  XOR U34050 ( .A(n34227), .B(n34177), .Z(n34179) );
  XOR U34051 ( .A(n34229), .B(n34230), .Z(n34219) );
  AND U34052 ( .A(n34231), .B(n34232), .Z(n34230) );
  XNOR U34053 ( .A(n34229), .B(n33952), .Z(n34232) );
  IV U34054 ( .A(n33955), .Z(n33952) );
  XOR U34055 ( .A(n34233), .B(n34234), .Z(n33955) );
  AND U34056 ( .A(n454), .B(n34235), .Z(n34234) );
  XNOR U34057 ( .A(n34236), .B(n34233), .Z(n34235) );
  XOR U34058 ( .A(n33956), .B(n34229), .Z(n34231) );
  XOR U34059 ( .A(n34237), .B(n34238), .Z(n33956) );
  AND U34060 ( .A(n462), .B(n34188), .Z(n34238) );
  XOR U34061 ( .A(n34237), .B(n34186), .Z(n34188) );
  XOR U34062 ( .A(n34239), .B(n34240), .Z(n34229) );
  AND U34063 ( .A(n34241), .B(n34242), .Z(n34240) );
  XNOR U34064 ( .A(n34239), .B(n34001), .Z(n34242) );
  IV U34065 ( .A(n34004), .Z(n34001) );
  XOR U34066 ( .A(n34243), .B(n34244), .Z(n34004) );
  AND U34067 ( .A(n454), .B(n34245), .Z(n34244) );
  XOR U34068 ( .A(n34246), .B(n34243), .Z(n34245) );
  XOR U34069 ( .A(n34005), .B(n34239), .Z(n34241) );
  XOR U34070 ( .A(n34247), .B(n34248), .Z(n34005) );
  AND U34071 ( .A(n462), .B(n34196), .Z(n34248) );
  XOR U34072 ( .A(n34247), .B(n34194), .Z(n34196) );
  XOR U34073 ( .A(n34135), .B(n34249), .Z(n34239) );
  AND U34074 ( .A(n34137), .B(n34250), .Z(n34249) );
  XNOR U34075 ( .A(n34135), .B(n34094), .Z(n34250) );
  IV U34076 ( .A(n34097), .Z(n34094) );
  XOR U34077 ( .A(n34251), .B(n34252), .Z(n34097) );
  AND U34078 ( .A(n454), .B(n34253), .Z(n34252) );
  XNOR U34079 ( .A(n34254), .B(n34251), .Z(n34253) );
  XOR U34080 ( .A(n34098), .B(n34135), .Z(n34137) );
  XOR U34081 ( .A(n34255), .B(n34256), .Z(n34098) );
  AND U34082 ( .A(n462), .B(n34206), .Z(n34256) );
  XOR U34083 ( .A(n34255), .B(n34204), .Z(n34206) );
  AND U34084 ( .A(n34207), .B(n34115), .Z(n34135) );
  XNOR U34085 ( .A(n34257), .B(n34258), .Z(n34115) );
  AND U34086 ( .A(n454), .B(n34259), .Z(n34258) );
  XNOR U34087 ( .A(n34260), .B(n34257), .Z(n34259) );
  XNOR U34088 ( .A(n34261), .B(n34262), .Z(n454) );
  AND U34089 ( .A(n34263), .B(n34264), .Z(n34262) );
  XOR U34090 ( .A(n34216), .B(n34261), .Z(n34264) );
  AND U34091 ( .A(n34265), .B(n34266), .Z(n34216) );
  XNOR U34092 ( .A(n34213), .B(n34261), .Z(n34263) );
  XNOR U34093 ( .A(n34267), .B(n34268), .Z(n34213) );
  AND U34094 ( .A(n458), .B(n34269), .Z(n34268) );
  XNOR U34095 ( .A(n34270), .B(n34271), .Z(n34269) );
  XOR U34096 ( .A(n34272), .B(n34273), .Z(n34261) );
  AND U34097 ( .A(n34274), .B(n34275), .Z(n34273) );
  XNOR U34098 ( .A(n34272), .B(n34265), .Z(n34275) );
  IV U34099 ( .A(n34226), .Z(n34265) );
  XOR U34100 ( .A(n34276), .B(n34277), .Z(n34226) );
  XOR U34101 ( .A(n34278), .B(n34266), .Z(n34277) );
  AND U34102 ( .A(n34236), .B(n34279), .Z(n34266) );
  AND U34103 ( .A(n34280), .B(n34281), .Z(n34278) );
  XOR U34104 ( .A(n34282), .B(n34276), .Z(n34280) );
  XNOR U34105 ( .A(n34223), .B(n34272), .Z(n34274) );
  XNOR U34106 ( .A(n34283), .B(n34284), .Z(n34223) );
  AND U34107 ( .A(n458), .B(n34285), .Z(n34284) );
  XNOR U34108 ( .A(n34286), .B(n34287), .Z(n34285) );
  XOR U34109 ( .A(n34288), .B(n34289), .Z(n34272) );
  AND U34110 ( .A(n34290), .B(n34291), .Z(n34289) );
  XNOR U34111 ( .A(n34288), .B(n34236), .Z(n34291) );
  XOR U34112 ( .A(n34292), .B(n34281), .Z(n34236) );
  XNOR U34113 ( .A(n34293), .B(n34276), .Z(n34281) );
  XOR U34114 ( .A(n34294), .B(n34295), .Z(n34276) );
  AND U34115 ( .A(n34296), .B(n34297), .Z(n34295) );
  XOR U34116 ( .A(n34298), .B(n34294), .Z(n34296) );
  XNOR U34117 ( .A(n34299), .B(n34300), .Z(n34293) );
  AND U34118 ( .A(n34301), .B(n34302), .Z(n34300) );
  XOR U34119 ( .A(n34299), .B(n34303), .Z(n34301) );
  XNOR U34120 ( .A(n34282), .B(n34279), .Z(n34292) );
  AND U34121 ( .A(n34304), .B(n34305), .Z(n34279) );
  XOR U34122 ( .A(n34306), .B(n34307), .Z(n34282) );
  AND U34123 ( .A(n34308), .B(n34309), .Z(n34307) );
  XOR U34124 ( .A(n34306), .B(n34310), .Z(n34308) );
  XNOR U34125 ( .A(n34233), .B(n34288), .Z(n34290) );
  XNOR U34126 ( .A(n34311), .B(n34312), .Z(n34233) );
  AND U34127 ( .A(n458), .B(n34313), .Z(n34312) );
  XNOR U34128 ( .A(n34314), .B(n34315), .Z(n34313) );
  XOR U34129 ( .A(n34316), .B(n34317), .Z(n34288) );
  AND U34130 ( .A(n34318), .B(n34319), .Z(n34317) );
  XNOR U34131 ( .A(n34316), .B(n34304), .Z(n34319) );
  IV U34132 ( .A(n34246), .Z(n34304) );
  XNOR U34133 ( .A(n34320), .B(n34297), .Z(n34246) );
  XNOR U34134 ( .A(n34321), .B(n34303), .Z(n34297) );
  XOR U34135 ( .A(n34322), .B(n34323), .Z(n34303) );
  AND U34136 ( .A(n34324), .B(n34325), .Z(n34323) );
  XOR U34137 ( .A(n34322), .B(n34326), .Z(n34324) );
  XNOR U34138 ( .A(n34302), .B(n34294), .Z(n34321) );
  XOR U34139 ( .A(n34327), .B(n34328), .Z(n34294) );
  AND U34140 ( .A(n34329), .B(n34330), .Z(n34328) );
  XNOR U34141 ( .A(n34331), .B(n34327), .Z(n34329) );
  XNOR U34142 ( .A(n34332), .B(n34299), .Z(n34302) );
  XOR U34143 ( .A(n34333), .B(n34334), .Z(n34299) );
  AND U34144 ( .A(n34335), .B(n34336), .Z(n34334) );
  XOR U34145 ( .A(n34333), .B(n34337), .Z(n34335) );
  XNOR U34146 ( .A(n34338), .B(n34339), .Z(n34332) );
  AND U34147 ( .A(n34340), .B(n34341), .Z(n34339) );
  XNOR U34148 ( .A(n34338), .B(n34342), .Z(n34340) );
  XNOR U34149 ( .A(n34298), .B(n34305), .Z(n34320) );
  AND U34150 ( .A(n34254), .B(n34343), .Z(n34305) );
  XOR U34151 ( .A(n34310), .B(n34309), .Z(n34298) );
  XNOR U34152 ( .A(n34344), .B(n34306), .Z(n34309) );
  XOR U34153 ( .A(n34345), .B(n34346), .Z(n34306) );
  AND U34154 ( .A(n34347), .B(n34348), .Z(n34346) );
  XOR U34155 ( .A(n34345), .B(n34349), .Z(n34347) );
  XNOR U34156 ( .A(n34350), .B(n34351), .Z(n34344) );
  AND U34157 ( .A(n34352), .B(n34353), .Z(n34351) );
  XOR U34158 ( .A(n34350), .B(n34354), .Z(n34352) );
  XOR U34159 ( .A(n34355), .B(n34356), .Z(n34310) );
  AND U34160 ( .A(n34357), .B(n34358), .Z(n34356) );
  XOR U34161 ( .A(n34355), .B(n34359), .Z(n34357) );
  XNOR U34162 ( .A(n34243), .B(n34316), .Z(n34318) );
  XNOR U34163 ( .A(n34360), .B(n34361), .Z(n34243) );
  AND U34164 ( .A(n458), .B(n34362), .Z(n34361) );
  XNOR U34165 ( .A(n34363), .B(n34364), .Z(n34362) );
  XOR U34166 ( .A(n34365), .B(n34366), .Z(n34316) );
  AND U34167 ( .A(n34367), .B(n34368), .Z(n34366) );
  XNOR U34168 ( .A(n34365), .B(n34254), .Z(n34368) );
  XOR U34169 ( .A(n34369), .B(n34330), .Z(n34254) );
  XNOR U34170 ( .A(n34370), .B(n34337), .Z(n34330) );
  XOR U34171 ( .A(n34326), .B(n34325), .Z(n34337) );
  XNOR U34172 ( .A(n34371), .B(n34322), .Z(n34325) );
  XOR U34173 ( .A(n34372), .B(n34373), .Z(n34322) );
  AND U34174 ( .A(n34374), .B(n34375), .Z(n34373) );
  XOR U34175 ( .A(n34372), .B(n34376), .Z(n34374) );
  XNOR U34176 ( .A(n34377), .B(n34378), .Z(n34371) );
  NOR U34177 ( .A(n34379), .B(n34380), .Z(n34378) );
  XNOR U34178 ( .A(n34377), .B(n34381), .Z(n34379) );
  XOR U34179 ( .A(n34382), .B(n34383), .Z(n34326) );
  NOR U34180 ( .A(n34384), .B(n34385), .Z(n34383) );
  XNOR U34181 ( .A(n34382), .B(n34386), .Z(n34384) );
  XNOR U34182 ( .A(n34336), .B(n34327), .Z(n34370) );
  XOR U34183 ( .A(n34387), .B(n34388), .Z(n34327) );
  NOR U34184 ( .A(n34389), .B(n34390), .Z(n34388) );
  XNOR U34185 ( .A(n34387), .B(n34391), .Z(n34389) );
  XOR U34186 ( .A(n34392), .B(n34342), .Z(n34336) );
  XNOR U34187 ( .A(n34393), .B(n34394), .Z(n34342) );
  NOR U34188 ( .A(n34395), .B(n34396), .Z(n34394) );
  XNOR U34189 ( .A(n34393), .B(n34397), .Z(n34395) );
  XNOR U34190 ( .A(n34341), .B(n34333), .Z(n34392) );
  XOR U34191 ( .A(n34398), .B(n34399), .Z(n34333) );
  AND U34192 ( .A(n34400), .B(n34401), .Z(n34399) );
  XOR U34193 ( .A(n34398), .B(n34402), .Z(n34400) );
  XNOR U34194 ( .A(n34403), .B(n34338), .Z(n34341) );
  XOR U34195 ( .A(n34404), .B(n34405), .Z(n34338) );
  AND U34196 ( .A(n34406), .B(n34407), .Z(n34405) );
  XOR U34197 ( .A(n34404), .B(n34408), .Z(n34406) );
  XNOR U34198 ( .A(n34409), .B(n34410), .Z(n34403) );
  NOR U34199 ( .A(n34411), .B(n34412), .Z(n34410) );
  XOR U34200 ( .A(n34409), .B(n34413), .Z(n34411) );
  XOR U34201 ( .A(n34331), .B(n34343), .Z(n34369) );
  NOR U34202 ( .A(n34260), .B(n34414), .Z(n34343) );
  XNOR U34203 ( .A(n34349), .B(n34348), .Z(n34331) );
  XNOR U34204 ( .A(n34415), .B(n34354), .Z(n34348) );
  XOR U34205 ( .A(n34416), .B(n34417), .Z(n34354) );
  NOR U34206 ( .A(n34418), .B(n34419), .Z(n34417) );
  XNOR U34207 ( .A(n34416), .B(n34420), .Z(n34418) );
  XNOR U34208 ( .A(n34353), .B(n34345), .Z(n34415) );
  XOR U34209 ( .A(n34421), .B(n34422), .Z(n34345) );
  AND U34210 ( .A(n34423), .B(n34424), .Z(n34422) );
  XNOR U34211 ( .A(n34421), .B(n34425), .Z(n34423) );
  XNOR U34212 ( .A(n34426), .B(n34350), .Z(n34353) );
  XOR U34213 ( .A(n34427), .B(n34428), .Z(n34350) );
  AND U34214 ( .A(n34429), .B(n34430), .Z(n34428) );
  XOR U34215 ( .A(n34427), .B(n34431), .Z(n34429) );
  XNOR U34216 ( .A(n34432), .B(n34433), .Z(n34426) );
  NOR U34217 ( .A(n34434), .B(n34435), .Z(n34433) );
  XOR U34218 ( .A(n34432), .B(n34436), .Z(n34434) );
  XOR U34219 ( .A(n34359), .B(n34358), .Z(n34349) );
  XNOR U34220 ( .A(n34437), .B(n34355), .Z(n34358) );
  XOR U34221 ( .A(n34438), .B(n34439), .Z(n34355) );
  AND U34222 ( .A(n34440), .B(n34441), .Z(n34439) );
  XOR U34223 ( .A(n34438), .B(n34442), .Z(n34440) );
  XNOR U34224 ( .A(n34443), .B(n34444), .Z(n34437) );
  NOR U34225 ( .A(n34445), .B(n34446), .Z(n34444) );
  XNOR U34226 ( .A(n34443), .B(n34447), .Z(n34445) );
  XOR U34227 ( .A(n34448), .B(n34449), .Z(n34359) );
  NOR U34228 ( .A(n34450), .B(n34451), .Z(n34449) );
  XNOR U34229 ( .A(n34448), .B(n34452), .Z(n34450) );
  XNOR U34230 ( .A(n34251), .B(n34365), .Z(n34367) );
  XNOR U34231 ( .A(n34453), .B(n34454), .Z(n34251) );
  AND U34232 ( .A(n458), .B(n34455), .Z(n34454) );
  XNOR U34233 ( .A(n34456), .B(n34457), .Z(n34455) );
  AND U34234 ( .A(n34257), .B(n34260), .Z(n34365) );
  XOR U34235 ( .A(n34458), .B(n34414), .Z(n34260) );
  XNOR U34236 ( .A(p_input[2048]), .B(p_input[544]), .Z(n34414) );
  XOR U34237 ( .A(n34391), .B(n34390), .Z(n34458) );
  XOR U34238 ( .A(n34459), .B(n34402), .Z(n34390) );
  XOR U34239 ( .A(n34376), .B(n34375), .Z(n34402) );
  XNOR U34240 ( .A(n34460), .B(n34381), .Z(n34375) );
  XOR U34241 ( .A(p_input[2072]), .B(p_input[568]), .Z(n34381) );
  XOR U34242 ( .A(n34372), .B(n34380), .Z(n34460) );
  XOR U34243 ( .A(n34461), .B(n34377), .Z(n34380) );
  XOR U34244 ( .A(p_input[2070]), .B(p_input[566]), .Z(n34377) );
  XNOR U34245 ( .A(p_input[2071]), .B(p_input[567]), .Z(n34461) );
  XNOR U34246 ( .A(n28684), .B(p_input[562]), .Z(n34372) );
  XNOR U34247 ( .A(n34386), .B(n34385), .Z(n34376) );
  XOR U34248 ( .A(n34462), .B(n34382), .Z(n34385) );
  XOR U34249 ( .A(p_input[2067]), .B(p_input[563]), .Z(n34382) );
  XNOR U34250 ( .A(p_input[2068]), .B(p_input[564]), .Z(n34462) );
  XOR U34251 ( .A(p_input[2069]), .B(p_input[565]), .Z(n34386) );
  XNOR U34252 ( .A(n34401), .B(n34387), .Z(n34459) );
  XNOR U34253 ( .A(n28686), .B(p_input[545]), .Z(n34387) );
  XNOR U34254 ( .A(n34463), .B(n34408), .Z(n34401) );
  XNOR U34255 ( .A(n34397), .B(n34396), .Z(n34408) );
  XOR U34256 ( .A(n34464), .B(n34393), .Z(n34396) );
  XNOR U34257 ( .A(n28322), .B(p_input[570]), .Z(n34393) );
  XNOR U34258 ( .A(p_input[2075]), .B(p_input[571]), .Z(n34464) );
  XOR U34259 ( .A(p_input[2076]), .B(p_input[572]), .Z(n34397) );
  XNOR U34260 ( .A(n34407), .B(n34398), .Z(n34463) );
  XNOR U34261 ( .A(n28689), .B(p_input[561]), .Z(n34398) );
  XOR U34262 ( .A(n34465), .B(n34413), .Z(n34407) );
  XNOR U34263 ( .A(p_input[2079]), .B(p_input[575]), .Z(n34413) );
  XOR U34264 ( .A(n34404), .B(n34412), .Z(n34465) );
  XOR U34265 ( .A(n34466), .B(n34409), .Z(n34412) );
  XOR U34266 ( .A(p_input[2077]), .B(p_input[573]), .Z(n34409) );
  XNOR U34267 ( .A(p_input[2078]), .B(p_input[574]), .Z(n34466) );
  XNOR U34268 ( .A(n28326), .B(p_input[569]), .Z(n34404) );
  XNOR U34269 ( .A(n34425), .B(n34424), .Z(n34391) );
  XNOR U34270 ( .A(n34467), .B(n34431), .Z(n34424) );
  XNOR U34271 ( .A(n34420), .B(n34419), .Z(n34431) );
  XOR U34272 ( .A(n34468), .B(n34416), .Z(n34419) );
  XNOR U34273 ( .A(n28694), .B(p_input[555]), .Z(n34416) );
  XNOR U34274 ( .A(p_input[2060]), .B(p_input[556]), .Z(n34468) );
  XOR U34275 ( .A(p_input[2061]), .B(p_input[557]), .Z(n34420) );
  XNOR U34276 ( .A(n34430), .B(n34421), .Z(n34467) );
  XNOR U34277 ( .A(n28330), .B(p_input[546]), .Z(n34421) );
  XOR U34278 ( .A(n34469), .B(n34436), .Z(n34430) );
  XNOR U34279 ( .A(p_input[2064]), .B(p_input[560]), .Z(n34436) );
  XOR U34280 ( .A(n34427), .B(n34435), .Z(n34469) );
  XOR U34281 ( .A(n34470), .B(n34432), .Z(n34435) );
  XOR U34282 ( .A(p_input[2062]), .B(p_input[558]), .Z(n34432) );
  XNOR U34283 ( .A(p_input[2063]), .B(p_input[559]), .Z(n34470) );
  XNOR U34284 ( .A(n28697), .B(p_input[554]), .Z(n34427) );
  XNOR U34285 ( .A(n34442), .B(n34441), .Z(n34425) );
  XNOR U34286 ( .A(n34471), .B(n34447), .Z(n34441) );
  XOR U34287 ( .A(p_input[2057]), .B(p_input[553]), .Z(n34447) );
  XOR U34288 ( .A(n34438), .B(n34446), .Z(n34471) );
  XOR U34289 ( .A(n34472), .B(n34443), .Z(n34446) );
  XOR U34290 ( .A(p_input[2055]), .B(p_input[551]), .Z(n34443) );
  XNOR U34291 ( .A(p_input[2056]), .B(p_input[552]), .Z(n34472) );
  XNOR U34292 ( .A(n28337), .B(p_input[547]), .Z(n34438) );
  XNOR U34293 ( .A(n34452), .B(n34451), .Z(n34442) );
  XOR U34294 ( .A(n34473), .B(n34448), .Z(n34451) );
  XOR U34295 ( .A(p_input[2052]), .B(p_input[548]), .Z(n34448) );
  XNOR U34296 ( .A(p_input[2053]), .B(p_input[549]), .Z(n34473) );
  XOR U34297 ( .A(p_input[2054]), .B(p_input[550]), .Z(n34452) );
  XNOR U34298 ( .A(n34474), .B(n34475), .Z(n34257) );
  AND U34299 ( .A(n458), .B(n34476), .Z(n34475) );
  XNOR U34300 ( .A(n34477), .B(n34478), .Z(n458) );
  AND U34301 ( .A(n34479), .B(n34480), .Z(n34478) );
  XOR U34302 ( .A(n34271), .B(n34477), .Z(n34480) );
  XNOR U34303 ( .A(n34481), .B(n34477), .Z(n34479) );
  XOR U34304 ( .A(n34482), .B(n34483), .Z(n34477) );
  AND U34305 ( .A(n34484), .B(n34485), .Z(n34483) );
  XOR U34306 ( .A(n34286), .B(n34482), .Z(n34485) );
  XOR U34307 ( .A(n34482), .B(n34287), .Z(n34484) );
  XOR U34308 ( .A(n34486), .B(n34487), .Z(n34482) );
  AND U34309 ( .A(n34488), .B(n34489), .Z(n34487) );
  XOR U34310 ( .A(n34314), .B(n34486), .Z(n34489) );
  XOR U34311 ( .A(n34486), .B(n34315), .Z(n34488) );
  XOR U34312 ( .A(n34490), .B(n34491), .Z(n34486) );
  AND U34313 ( .A(n34492), .B(n34493), .Z(n34491) );
  XOR U34314 ( .A(n34363), .B(n34490), .Z(n34493) );
  XOR U34315 ( .A(n34490), .B(n34364), .Z(n34492) );
  XOR U34316 ( .A(n34494), .B(n34495), .Z(n34490) );
  AND U34317 ( .A(n34496), .B(n34497), .Z(n34495) );
  XOR U34318 ( .A(n34494), .B(n34456), .Z(n34497) );
  XNOR U34319 ( .A(n34498), .B(n34499), .Z(n34207) );
  AND U34320 ( .A(n462), .B(n34500), .Z(n34499) );
  XNOR U34321 ( .A(n34501), .B(n34502), .Z(n462) );
  AND U34322 ( .A(n34503), .B(n34504), .Z(n34502) );
  XOR U34323 ( .A(n34501), .B(n34217), .Z(n34504) );
  XNOR U34324 ( .A(n34501), .B(n34167), .Z(n34503) );
  XOR U34325 ( .A(n34505), .B(n34506), .Z(n34501) );
  AND U34326 ( .A(n34507), .B(n34508), .Z(n34506) );
  XNOR U34327 ( .A(n34227), .B(n34505), .Z(n34508) );
  XOR U34328 ( .A(n34505), .B(n34177), .Z(n34507) );
  XOR U34329 ( .A(n34509), .B(n34510), .Z(n34505) );
  AND U34330 ( .A(n34511), .B(n34512), .Z(n34510) );
  XNOR U34331 ( .A(n34237), .B(n34509), .Z(n34512) );
  XOR U34332 ( .A(n34509), .B(n34186), .Z(n34511) );
  XOR U34333 ( .A(n34513), .B(n34514), .Z(n34509) );
  AND U34334 ( .A(n34515), .B(n34516), .Z(n34514) );
  XOR U34335 ( .A(n34513), .B(n34194), .Z(n34515) );
  XOR U34336 ( .A(n34517), .B(n34518), .Z(n34158) );
  AND U34337 ( .A(n466), .B(n34500), .Z(n34518) );
  XNOR U34338 ( .A(n34498), .B(n34517), .Z(n34500) );
  XNOR U34339 ( .A(n34519), .B(n34520), .Z(n466) );
  AND U34340 ( .A(n34521), .B(n34522), .Z(n34520) );
  XNOR U34341 ( .A(n34523), .B(n34519), .Z(n34522) );
  IV U34342 ( .A(n34217), .Z(n34523) );
  XOR U34343 ( .A(n34481), .B(n34524), .Z(n34217) );
  AND U34344 ( .A(n469), .B(n34525), .Z(n34524) );
  XOR U34345 ( .A(n34270), .B(n34267), .Z(n34525) );
  IV U34346 ( .A(n34481), .Z(n34270) );
  XNOR U34347 ( .A(n34167), .B(n34519), .Z(n34521) );
  XOR U34348 ( .A(n34526), .B(n34527), .Z(n34167) );
  AND U34349 ( .A(n485), .B(n34528), .Z(n34527) );
  XOR U34350 ( .A(n34529), .B(n34530), .Z(n34519) );
  AND U34351 ( .A(n34531), .B(n34532), .Z(n34530) );
  XNOR U34352 ( .A(n34529), .B(n34227), .Z(n34532) );
  XOR U34353 ( .A(n34287), .B(n34533), .Z(n34227) );
  AND U34354 ( .A(n469), .B(n34534), .Z(n34533) );
  XOR U34355 ( .A(n34283), .B(n34287), .Z(n34534) );
  XNOR U34356 ( .A(n34535), .B(n34529), .Z(n34531) );
  IV U34357 ( .A(n34177), .Z(n34535) );
  XOR U34358 ( .A(n34536), .B(n34537), .Z(n34177) );
  AND U34359 ( .A(n485), .B(n34538), .Z(n34537) );
  XOR U34360 ( .A(n34539), .B(n34540), .Z(n34529) );
  AND U34361 ( .A(n34541), .B(n34542), .Z(n34540) );
  XNOR U34362 ( .A(n34539), .B(n34237), .Z(n34542) );
  XOR U34363 ( .A(n34315), .B(n34543), .Z(n34237) );
  AND U34364 ( .A(n469), .B(n34544), .Z(n34543) );
  XOR U34365 ( .A(n34311), .B(n34315), .Z(n34544) );
  XOR U34366 ( .A(n34186), .B(n34539), .Z(n34541) );
  XOR U34367 ( .A(n34545), .B(n34546), .Z(n34186) );
  AND U34368 ( .A(n485), .B(n34547), .Z(n34546) );
  XOR U34369 ( .A(n34513), .B(n34548), .Z(n34539) );
  AND U34370 ( .A(n34549), .B(n34516), .Z(n34548) );
  XNOR U34371 ( .A(n34247), .B(n34513), .Z(n34516) );
  XOR U34372 ( .A(n34364), .B(n34550), .Z(n34247) );
  AND U34373 ( .A(n469), .B(n34551), .Z(n34550) );
  XOR U34374 ( .A(n34360), .B(n34364), .Z(n34551) );
  XNOR U34375 ( .A(n34552), .B(n34513), .Z(n34549) );
  IV U34376 ( .A(n34194), .Z(n34552) );
  XOR U34377 ( .A(n34553), .B(n34554), .Z(n34194) );
  AND U34378 ( .A(n485), .B(n34555), .Z(n34554) );
  XOR U34379 ( .A(n34556), .B(n34557), .Z(n34513) );
  AND U34380 ( .A(n34558), .B(n34559), .Z(n34557) );
  XNOR U34381 ( .A(n34556), .B(n34255), .Z(n34559) );
  XOR U34382 ( .A(n34457), .B(n34560), .Z(n34255) );
  AND U34383 ( .A(n469), .B(n34561), .Z(n34560) );
  XOR U34384 ( .A(n34453), .B(n34457), .Z(n34561) );
  XNOR U34385 ( .A(n34562), .B(n34556), .Z(n34558) );
  IV U34386 ( .A(n34204), .Z(n34562) );
  XOR U34387 ( .A(n34563), .B(n34564), .Z(n34204) );
  AND U34388 ( .A(n485), .B(n34565), .Z(n34564) );
  AND U34389 ( .A(n34517), .B(n34498), .Z(n34556) );
  XNOR U34390 ( .A(n34566), .B(n34567), .Z(n34498) );
  AND U34391 ( .A(n469), .B(n34476), .Z(n34567) );
  XNOR U34392 ( .A(n34474), .B(n34566), .Z(n34476) );
  XNOR U34393 ( .A(n34568), .B(n34569), .Z(n469) );
  AND U34394 ( .A(n34570), .B(n34571), .Z(n34569) );
  XNOR U34395 ( .A(n34568), .B(n34267), .Z(n34571) );
  IV U34396 ( .A(n34271), .Z(n34267) );
  XOR U34397 ( .A(n34572), .B(n34573), .Z(n34271) );
  AND U34398 ( .A(n473), .B(n34574), .Z(n34573) );
  XOR U34399 ( .A(n34575), .B(n34572), .Z(n34574) );
  XNOR U34400 ( .A(n34568), .B(n34481), .Z(n34570) );
  XOR U34401 ( .A(n34576), .B(n34577), .Z(n34481) );
  AND U34402 ( .A(n481), .B(n34528), .Z(n34577) );
  XOR U34403 ( .A(n34526), .B(n34576), .Z(n34528) );
  XOR U34404 ( .A(n34578), .B(n34579), .Z(n34568) );
  AND U34405 ( .A(n34580), .B(n34581), .Z(n34579) );
  XNOR U34406 ( .A(n34578), .B(n34283), .Z(n34581) );
  IV U34407 ( .A(n34286), .Z(n34283) );
  XOR U34408 ( .A(n34582), .B(n34583), .Z(n34286) );
  AND U34409 ( .A(n473), .B(n34584), .Z(n34583) );
  XOR U34410 ( .A(n34585), .B(n34582), .Z(n34584) );
  XOR U34411 ( .A(n34287), .B(n34578), .Z(n34580) );
  XOR U34412 ( .A(n34586), .B(n34587), .Z(n34287) );
  AND U34413 ( .A(n481), .B(n34538), .Z(n34587) );
  XOR U34414 ( .A(n34586), .B(n34536), .Z(n34538) );
  XOR U34415 ( .A(n34588), .B(n34589), .Z(n34578) );
  AND U34416 ( .A(n34590), .B(n34591), .Z(n34589) );
  XNOR U34417 ( .A(n34588), .B(n34311), .Z(n34591) );
  IV U34418 ( .A(n34314), .Z(n34311) );
  XOR U34419 ( .A(n34592), .B(n34593), .Z(n34314) );
  AND U34420 ( .A(n473), .B(n34594), .Z(n34593) );
  XNOR U34421 ( .A(n34595), .B(n34592), .Z(n34594) );
  XOR U34422 ( .A(n34315), .B(n34588), .Z(n34590) );
  XOR U34423 ( .A(n34596), .B(n34597), .Z(n34315) );
  AND U34424 ( .A(n481), .B(n34547), .Z(n34597) );
  XOR U34425 ( .A(n34596), .B(n34545), .Z(n34547) );
  XOR U34426 ( .A(n34598), .B(n34599), .Z(n34588) );
  AND U34427 ( .A(n34600), .B(n34601), .Z(n34599) );
  XNOR U34428 ( .A(n34598), .B(n34360), .Z(n34601) );
  IV U34429 ( .A(n34363), .Z(n34360) );
  XOR U34430 ( .A(n34602), .B(n34603), .Z(n34363) );
  AND U34431 ( .A(n473), .B(n34604), .Z(n34603) );
  XOR U34432 ( .A(n34605), .B(n34602), .Z(n34604) );
  XOR U34433 ( .A(n34364), .B(n34598), .Z(n34600) );
  XOR U34434 ( .A(n34606), .B(n34607), .Z(n34364) );
  AND U34435 ( .A(n481), .B(n34555), .Z(n34607) );
  XOR U34436 ( .A(n34606), .B(n34553), .Z(n34555) );
  XOR U34437 ( .A(n34494), .B(n34608), .Z(n34598) );
  AND U34438 ( .A(n34496), .B(n34609), .Z(n34608) );
  XNOR U34439 ( .A(n34494), .B(n34453), .Z(n34609) );
  IV U34440 ( .A(n34456), .Z(n34453) );
  XOR U34441 ( .A(n34610), .B(n34611), .Z(n34456) );
  AND U34442 ( .A(n473), .B(n34612), .Z(n34611) );
  XNOR U34443 ( .A(n34613), .B(n34610), .Z(n34612) );
  XOR U34444 ( .A(n34457), .B(n34494), .Z(n34496) );
  XOR U34445 ( .A(n34614), .B(n34615), .Z(n34457) );
  AND U34446 ( .A(n481), .B(n34565), .Z(n34615) );
  XOR U34447 ( .A(n34614), .B(n34563), .Z(n34565) );
  AND U34448 ( .A(n34566), .B(n34474), .Z(n34494) );
  XNOR U34449 ( .A(n34616), .B(n34617), .Z(n34474) );
  AND U34450 ( .A(n473), .B(n34618), .Z(n34617) );
  XNOR U34451 ( .A(n34619), .B(n34616), .Z(n34618) );
  XNOR U34452 ( .A(n34620), .B(n34621), .Z(n473) );
  AND U34453 ( .A(n34622), .B(n34623), .Z(n34621) );
  XOR U34454 ( .A(n34575), .B(n34620), .Z(n34623) );
  AND U34455 ( .A(n34624), .B(n34625), .Z(n34575) );
  XNOR U34456 ( .A(n34572), .B(n34620), .Z(n34622) );
  XNOR U34457 ( .A(n34626), .B(n34627), .Z(n34572) );
  AND U34458 ( .A(n477), .B(n34628), .Z(n34627) );
  XNOR U34459 ( .A(n34629), .B(n34630), .Z(n34628) );
  XOR U34460 ( .A(n34631), .B(n34632), .Z(n34620) );
  AND U34461 ( .A(n34633), .B(n34634), .Z(n34632) );
  XNOR U34462 ( .A(n34631), .B(n34624), .Z(n34634) );
  IV U34463 ( .A(n34585), .Z(n34624) );
  XOR U34464 ( .A(n34635), .B(n34636), .Z(n34585) );
  XOR U34465 ( .A(n34637), .B(n34625), .Z(n34636) );
  AND U34466 ( .A(n34595), .B(n34638), .Z(n34625) );
  AND U34467 ( .A(n34639), .B(n34640), .Z(n34637) );
  XOR U34468 ( .A(n34641), .B(n34635), .Z(n34639) );
  XNOR U34469 ( .A(n34582), .B(n34631), .Z(n34633) );
  XNOR U34470 ( .A(n34642), .B(n34643), .Z(n34582) );
  AND U34471 ( .A(n477), .B(n34644), .Z(n34643) );
  XNOR U34472 ( .A(n34645), .B(n34646), .Z(n34644) );
  XOR U34473 ( .A(n34647), .B(n34648), .Z(n34631) );
  AND U34474 ( .A(n34649), .B(n34650), .Z(n34648) );
  XNOR U34475 ( .A(n34647), .B(n34595), .Z(n34650) );
  XOR U34476 ( .A(n34651), .B(n34640), .Z(n34595) );
  XNOR U34477 ( .A(n34652), .B(n34635), .Z(n34640) );
  XOR U34478 ( .A(n34653), .B(n34654), .Z(n34635) );
  AND U34479 ( .A(n34655), .B(n34656), .Z(n34654) );
  XOR U34480 ( .A(n34657), .B(n34653), .Z(n34655) );
  XNOR U34481 ( .A(n34658), .B(n34659), .Z(n34652) );
  AND U34482 ( .A(n34660), .B(n34661), .Z(n34659) );
  XOR U34483 ( .A(n34658), .B(n34662), .Z(n34660) );
  XNOR U34484 ( .A(n34641), .B(n34638), .Z(n34651) );
  AND U34485 ( .A(n34663), .B(n34664), .Z(n34638) );
  XOR U34486 ( .A(n34665), .B(n34666), .Z(n34641) );
  AND U34487 ( .A(n34667), .B(n34668), .Z(n34666) );
  XOR U34488 ( .A(n34665), .B(n34669), .Z(n34667) );
  XNOR U34489 ( .A(n34592), .B(n34647), .Z(n34649) );
  XNOR U34490 ( .A(n34670), .B(n34671), .Z(n34592) );
  AND U34491 ( .A(n477), .B(n34672), .Z(n34671) );
  XNOR U34492 ( .A(n34673), .B(n34674), .Z(n34672) );
  XOR U34493 ( .A(n34675), .B(n34676), .Z(n34647) );
  AND U34494 ( .A(n34677), .B(n34678), .Z(n34676) );
  XNOR U34495 ( .A(n34675), .B(n34663), .Z(n34678) );
  IV U34496 ( .A(n34605), .Z(n34663) );
  XNOR U34497 ( .A(n34679), .B(n34656), .Z(n34605) );
  XNOR U34498 ( .A(n34680), .B(n34662), .Z(n34656) );
  XOR U34499 ( .A(n34681), .B(n34682), .Z(n34662) );
  AND U34500 ( .A(n34683), .B(n34684), .Z(n34682) );
  XOR U34501 ( .A(n34681), .B(n34685), .Z(n34683) );
  XNOR U34502 ( .A(n34661), .B(n34653), .Z(n34680) );
  XOR U34503 ( .A(n34686), .B(n34687), .Z(n34653) );
  AND U34504 ( .A(n34688), .B(n34689), .Z(n34687) );
  XNOR U34505 ( .A(n34690), .B(n34686), .Z(n34688) );
  XNOR U34506 ( .A(n34691), .B(n34658), .Z(n34661) );
  XOR U34507 ( .A(n34692), .B(n34693), .Z(n34658) );
  AND U34508 ( .A(n34694), .B(n34695), .Z(n34693) );
  XOR U34509 ( .A(n34692), .B(n34696), .Z(n34694) );
  XNOR U34510 ( .A(n34697), .B(n34698), .Z(n34691) );
  AND U34511 ( .A(n34699), .B(n34700), .Z(n34698) );
  XNOR U34512 ( .A(n34697), .B(n34701), .Z(n34699) );
  XNOR U34513 ( .A(n34657), .B(n34664), .Z(n34679) );
  AND U34514 ( .A(n34613), .B(n34702), .Z(n34664) );
  XOR U34515 ( .A(n34669), .B(n34668), .Z(n34657) );
  XNOR U34516 ( .A(n34703), .B(n34665), .Z(n34668) );
  XOR U34517 ( .A(n34704), .B(n34705), .Z(n34665) );
  AND U34518 ( .A(n34706), .B(n34707), .Z(n34705) );
  XOR U34519 ( .A(n34704), .B(n34708), .Z(n34706) );
  XNOR U34520 ( .A(n34709), .B(n34710), .Z(n34703) );
  AND U34521 ( .A(n34711), .B(n34712), .Z(n34710) );
  XOR U34522 ( .A(n34709), .B(n34713), .Z(n34711) );
  XOR U34523 ( .A(n34714), .B(n34715), .Z(n34669) );
  AND U34524 ( .A(n34716), .B(n34717), .Z(n34715) );
  XOR U34525 ( .A(n34714), .B(n34718), .Z(n34716) );
  XNOR U34526 ( .A(n34602), .B(n34675), .Z(n34677) );
  XNOR U34527 ( .A(n34719), .B(n34720), .Z(n34602) );
  AND U34528 ( .A(n477), .B(n34721), .Z(n34720) );
  XNOR U34529 ( .A(n34722), .B(n34723), .Z(n34721) );
  XOR U34530 ( .A(n34724), .B(n34725), .Z(n34675) );
  AND U34531 ( .A(n34726), .B(n34727), .Z(n34725) );
  XNOR U34532 ( .A(n34724), .B(n34613), .Z(n34727) );
  XOR U34533 ( .A(n34728), .B(n34689), .Z(n34613) );
  XNOR U34534 ( .A(n34729), .B(n34696), .Z(n34689) );
  XOR U34535 ( .A(n34685), .B(n34684), .Z(n34696) );
  XNOR U34536 ( .A(n34730), .B(n34681), .Z(n34684) );
  XOR U34537 ( .A(n34731), .B(n34732), .Z(n34681) );
  AND U34538 ( .A(n34733), .B(n34734), .Z(n34732) );
  XOR U34539 ( .A(n34731), .B(n34735), .Z(n34733) );
  XNOR U34540 ( .A(n34736), .B(n34737), .Z(n34730) );
  NOR U34541 ( .A(n34738), .B(n34739), .Z(n34737) );
  XNOR U34542 ( .A(n34736), .B(n34740), .Z(n34738) );
  XOR U34543 ( .A(n34741), .B(n34742), .Z(n34685) );
  NOR U34544 ( .A(n34743), .B(n34744), .Z(n34742) );
  XNOR U34545 ( .A(n34741), .B(n34745), .Z(n34743) );
  XNOR U34546 ( .A(n34695), .B(n34686), .Z(n34729) );
  XOR U34547 ( .A(n34746), .B(n34747), .Z(n34686) );
  NOR U34548 ( .A(n34748), .B(n34749), .Z(n34747) );
  XNOR U34549 ( .A(n34746), .B(n34750), .Z(n34748) );
  XOR U34550 ( .A(n34751), .B(n34701), .Z(n34695) );
  XNOR U34551 ( .A(n34752), .B(n34753), .Z(n34701) );
  NOR U34552 ( .A(n34754), .B(n34755), .Z(n34753) );
  XNOR U34553 ( .A(n34752), .B(n34756), .Z(n34754) );
  XNOR U34554 ( .A(n34700), .B(n34692), .Z(n34751) );
  XOR U34555 ( .A(n34757), .B(n34758), .Z(n34692) );
  AND U34556 ( .A(n34759), .B(n34760), .Z(n34758) );
  XOR U34557 ( .A(n34757), .B(n34761), .Z(n34759) );
  XNOR U34558 ( .A(n34762), .B(n34697), .Z(n34700) );
  XOR U34559 ( .A(n34763), .B(n34764), .Z(n34697) );
  AND U34560 ( .A(n34765), .B(n34766), .Z(n34764) );
  XOR U34561 ( .A(n34763), .B(n34767), .Z(n34765) );
  XNOR U34562 ( .A(n34768), .B(n34769), .Z(n34762) );
  NOR U34563 ( .A(n34770), .B(n34771), .Z(n34769) );
  XOR U34564 ( .A(n34768), .B(n34772), .Z(n34770) );
  XOR U34565 ( .A(n34690), .B(n34702), .Z(n34728) );
  NOR U34566 ( .A(n34619), .B(n34773), .Z(n34702) );
  XNOR U34567 ( .A(n34708), .B(n34707), .Z(n34690) );
  XNOR U34568 ( .A(n34774), .B(n34713), .Z(n34707) );
  XOR U34569 ( .A(n34775), .B(n34776), .Z(n34713) );
  NOR U34570 ( .A(n34777), .B(n34778), .Z(n34776) );
  XNOR U34571 ( .A(n34775), .B(n34779), .Z(n34777) );
  XNOR U34572 ( .A(n34712), .B(n34704), .Z(n34774) );
  XOR U34573 ( .A(n34780), .B(n34781), .Z(n34704) );
  AND U34574 ( .A(n34782), .B(n34783), .Z(n34781) );
  XNOR U34575 ( .A(n34780), .B(n34784), .Z(n34782) );
  XNOR U34576 ( .A(n34785), .B(n34709), .Z(n34712) );
  XOR U34577 ( .A(n34786), .B(n34787), .Z(n34709) );
  AND U34578 ( .A(n34788), .B(n34789), .Z(n34787) );
  XOR U34579 ( .A(n34786), .B(n34790), .Z(n34788) );
  XNOR U34580 ( .A(n34791), .B(n34792), .Z(n34785) );
  NOR U34581 ( .A(n34793), .B(n34794), .Z(n34792) );
  XOR U34582 ( .A(n34791), .B(n34795), .Z(n34793) );
  XOR U34583 ( .A(n34718), .B(n34717), .Z(n34708) );
  XNOR U34584 ( .A(n34796), .B(n34714), .Z(n34717) );
  XOR U34585 ( .A(n34797), .B(n34798), .Z(n34714) );
  AND U34586 ( .A(n34799), .B(n34800), .Z(n34798) );
  XOR U34587 ( .A(n34797), .B(n34801), .Z(n34799) );
  XNOR U34588 ( .A(n34802), .B(n34803), .Z(n34796) );
  NOR U34589 ( .A(n34804), .B(n34805), .Z(n34803) );
  XNOR U34590 ( .A(n34802), .B(n34806), .Z(n34804) );
  XOR U34591 ( .A(n34807), .B(n34808), .Z(n34718) );
  NOR U34592 ( .A(n34809), .B(n34810), .Z(n34808) );
  XNOR U34593 ( .A(n34807), .B(n34811), .Z(n34809) );
  XNOR U34594 ( .A(n34610), .B(n34724), .Z(n34726) );
  XNOR U34595 ( .A(n34812), .B(n34813), .Z(n34610) );
  AND U34596 ( .A(n477), .B(n34814), .Z(n34813) );
  XNOR U34597 ( .A(n34815), .B(n34816), .Z(n34814) );
  AND U34598 ( .A(n34616), .B(n34619), .Z(n34724) );
  XOR U34599 ( .A(n34817), .B(n34773), .Z(n34619) );
  XNOR U34600 ( .A(p_input[2048]), .B(p_input[576]), .Z(n34773) );
  XOR U34601 ( .A(n34750), .B(n34749), .Z(n34817) );
  XOR U34602 ( .A(n34818), .B(n34761), .Z(n34749) );
  XOR U34603 ( .A(n34735), .B(n34734), .Z(n34761) );
  XNOR U34604 ( .A(n34819), .B(n34740), .Z(n34734) );
  XOR U34605 ( .A(p_input[2072]), .B(p_input[600]), .Z(n34740) );
  XOR U34606 ( .A(n34731), .B(n34739), .Z(n34819) );
  XOR U34607 ( .A(n34820), .B(n34736), .Z(n34739) );
  XOR U34608 ( .A(p_input[2070]), .B(p_input[598]), .Z(n34736) );
  XNOR U34609 ( .A(p_input[2071]), .B(p_input[599]), .Z(n34820) );
  XNOR U34610 ( .A(n28684), .B(p_input[594]), .Z(n34731) );
  XNOR U34611 ( .A(n34745), .B(n34744), .Z(n34735) );
  XOR U34612 ( .A(n34821), .B(n34741), .Z(n34744) );
  XOR U34613 ( .A(p_input[2067]), .B(p_input[595]), .Z(n34741) );
  XNOR U34614 ( .A(p_input[2068]), .B(p_input[596]), .Z(n34821) );
  XOR U34615 ( .A(p_input[2069]), .B(p_input[597]), .Z(n34745) );
  XNOR U34616 ( .A(n34760), .B(n34746), .Z(n34818) );
  XNOR U34617 ( .A(n28686), .B(p_input[577]), .Z(n34746) );
  XNOR U34618 ( .A(n34822), .B(n34767), .Z(n34760) );
  XNOR U34619 ( .A(n34756), .B(n34755), .Z(n34767) );
  XOR U34620 ( .A(n34823), .B(n34752), .Z(n34755) );
  XNOR U34621 ( .A(n28322), .B(p_input[602]), .Z(n34752) );
  XNOR U34622 ( .A(p_input[2075]), .B(p_input[603]), .Z(n34823) );
  XOR U34623 ( .A(p_input[2076]), .B(p_input[604]), .Z(n34756) );
  XNOR U34624 ( .A(n34766), .B(n34757), .Z(n34822) );
  XNOR U34625 ( .A(n28689), .B(p_input[593]), .Z(n34757) );
  XOR U34626 ( .A(n34824), .B(n34772), .Z(n34766) );
  XNOR U34627 ( .A(p_input[2079]), .B(p_input[607]), .Z(n34772) );
  XOR U34628 ( .A(n34763), .B(n34771), .Z(n34824) );
  XOR U34629 ( .A(n34825), .B(n34768), .Z(n34771) );
  XOR U34630 ( .A(p_input[2077]), .B(p_input[605]), .Z(n34768) );
  XNOR U34631 ( .A(p_input[2078]), .B(p_input[606]), .Z(n34825) );
  XNOR U34632 ( .A(n28326), .B(p_input[601]), .Z(n34763) );
  XNOR U34633 ( .A(n34784), .B(n34783), .Z(n34750) );
  XNOR U34634 ( .A(n34826), .B(n34790), .Z(n34783) );
  XNOR U34635 ( .A(n34779), .B(n34778), .Z(n34790) );
  XOR U34636 ( .A(n34827), .B(n34775), .Z(n34778) );
  XNOR U34637 ( .A(n28694), .B(p_input[587]), .Z(n34775) );
  XNOR U34638 ( .A(p_input[2060]), .B(p_input[588]), .Z(n34827) );
  XOR U34639 ( .A(p_input[2061]), .B(p_input[589]), .Z(n34779) );
  XNOR U34640 ( .A(n34789), .B(n34780), .Z(n34826) );
  XNOR U34641 ( .A(n28330), .B(p_input[578]), .Z(n34780) );
  XOR U34642 ( .A(n34828), .B(n34795), .Z(n34789) );
  XNOR U34643 ( .A(p_input[2064]), .B(p_input[592]), .Z(n34795) );
  XOR U34644 ( .A(n34786), .B(n34794), .Z(n34828) );
  XOR U34645 ( .A(n34829), .B(n34791), .Z(n34794) );
  XOR U34646 ( .A(p_input[2062]), .B(p_input[590]), .Z(n34791) );
  XNOR U34647 ( .A(p_input[2063]), .B(p_input[591]), .Z(n34829) );
  XNOR U34648 ( .A(n28697), .B(p_input[586]), .Z(n34786) );
  XNOR U34649 ( .A(n34801), .B(n34800), .Z(n34784) );
  XNOR U34650 ( .A(n34830), .B(n34806), .Z(n34800) );
  XOR U34651 ( .A(p_input[2057]), .B(p_input[585]), .Z(n34806) );
  XOR U34652 ( .A(n34797), .B(n34805), .Z(n34830) );
  XOR U34653 ( .A(n34831), .B(n34802), .Z(n34805) );
  XOR U34654 ( .A(p_input[2055]), .B(p_input[583]), .Z(n34802) );
  XNOR U34655 ( .A(p_input[2056]), .B(p_input[584]), .Z(n34831) );
  XNOR U34656 ( .A(n28337), .B(p_input[579]), .Z(n34797) );
  XNOR U34657 ( .A(n34811), .B(n34810), .Z(n34801) );
  XOR U34658 ( .A(n34832), .B(n34807), .Z(n34810) );
  XOR U34659 ( .A(p_input[2052]), .B(p_input[580]), .Z(n34807) );
  XNOR U34660 ( .A(p_input[2053]), .B(p_input[581]), .Z(n34832) );
  XOR U34661 ( .A(p_input[2054]), .B(p_input[582]), .Z(n34811) );
  XNOR U34662 ( .A(n34833), .B(n34834), .Z(n34616) );
  AND U34663 ( .A(n477), .B(n34835), .Z(n34834) );
  XNOR U34664 ( .A(n34836), .B(n34837), .Z(n477) );
  AND U34665 ( .A(n34838), .B(n34839), .Z(n34837) );
  XOR U34666 ( .A(n34630), .B(n34836), .Z(n34839) );
  XNOR U34667 ( .A(n34840), .B(n34836), .Z(n34838) );
  XOR U34668 ( .A(n34841), .B(n34842), .Z(n34836) );
  AND U34669 ( .A(n34843), .B(n34844), .Z(n34842) );
  XOR U34670 ( .A(n34645), .B(n34841), .Z(n34844) );
  XOR U34671 ( .A(n34841), .B(n34646), .Z(n34843) );
  XOR U34672 ( .A(n34845), .B(n34846), .Z(n34841) );
  AND U34673 ( .A(n34847), .B(n34848), .Z(n34846) );
  XOR U34674 ( .A(n34673), .B(n34845), .Z(n34848) );
  XOR U34675 ( .A(n34845), .B(n34674), .Z(n34847) );
  XOR U34676 ( .A(n34849), .B(n34850), .Z(n34845) );
  AND U34677 ( .A(n34851), .B(n34852), .Z(n34850) );
  XOR U34678 ( .A(n34722), .B(n34849), .Z(n34852) );
  XOR U34679 ( .A(n34849), .B(n34723), .Z(n34851) );
  XOR U34680 ( .A(n34853), .B(n34854), .Z(n34849) );
  AND U34681 ( .A(n34855), .B(n34856), .Z(n34854) );
  XOR U34682 ( .A(n34853), .B(n34815), .Z(n34856) );
  XNOR U34683 ( .A(n34857), .B(n34858), .Z(n34566) );
  AND U34684 ( .A(n481), .B(n34859), .Z(n34858) );
  XNOR U34685 ( .A(n34860), .B(n34861), .Z(n481) );
  AND U34686 ( .A(n34862), .B(n34863), .Z(n34861) );
  XOR U34687 ( .A(n34860), .B(n34576), .Z(n34863) );
  XNOR U34688 ( .A(n34860), .B(n34526), .Z(n34862) );
  XOR U34689 ( .A(n34864), .B(n34865), .Z(n34860) );
  AND U34690 ( .A(n34866), .B(n34867), .Z(n34865) );
  XNOR U34691 ( .A(n34586), .B(n34864), .Z(n34867) );
  XOR U34692 ( .A(n34864), .B(n34536), .Z(n34866) );
  XOR U34693 ( .A(n34868), .B(n34869), .Z(n34864) );
  AND U34694 ( .A(n34870), .B(n34871), .Z(n34869) );
  XNOR U34695 ( .A(n34596), .B(n34868), .Z(n34871) );
  XOR U34696 ( .A(n34868), .B(n34545), .Z(n34870) );
  XOR U34697 ( .A(n34872), .B(n34873), .Z(n34868) );
  AND U34698 ( .A(n34874), .B(n34875), .Z(n34873) );
  XOR U34699 ( .A(n34872), .B(n34553), .Z(n34874) );
  XOR U34700 ( .A(n34876), .B(n34877), .Z(n34517) );
  AND U34701 ( .A(n485), .B(n34859), .Z(n34877) );
  XNOR U34702 ( .A(n34857), .B(n34876), .Z(n34859) );
  XNOR U34703 ( .A(n34878), .B(n34879), .Z(n485) );
  AND U34704 ( .A(n34880), .B(n34881), .Z(n34879) );
  XNOR U34705 ( .A(n34882), .B(n34878), .Z(n34881) );
  IV U34706 ( .A(n34576), .Z(n34882) );
  XOR U34707 ( .A(n34840), .B(n34883), .Z(n34576) );
  AND U34708 ( .A(n488), .B(n34884), .Z(n34883) );
  XOR U34709 ( .A(n34629), .B(n34626), .Z(n34884) );
  IV U34710 ( .A(n34840), .Z(n34629) );
  XNOR U34711 ( .A(n34526), .B(n34878), .Z(n34880) );
  XOR U34712 ( .A(n34885), .B(n34886), .Z(n34526) );
  AND U34713 ( .A(n504), .B(n34887), .Z(n34886) );
  XOR U34714 ( .A(n34888), .B(n34889), .Z(n34878) );
  AND U34715 ( .A(n34890), .B(n34891), .Z(n34889) );
  XNOR U34716 ( .A(n34888), .B(n34586), .Z(n34891) );
  XOR U34717 ( .A(n34646), .B(n34892), .Z(n34586) );
  AND U34718 ( .A(n488), .B(n34893), .Z(n34892) );
  XOR U34719 ( .A(n34642), .B(n34646), .Z(n34893) );
  XNOR U34720 ( .A(n34894), .B(n34888), .Z(n34890) );
  IV U34721 ( .A(n34536), .Z(n34894) );
  XOR U34722 ( .A(n34895), .B(n34896), .Z(n34536) );
  AND U34723 ( .A(n504), .B(n34897), .Z(n34896) );
  XOR U34724 ( .A(n34898), .B(n34899), .Z(n34888) );
  AND U34725 ( .A(n34900), .B(n34901), .Z(n34899) );
  XNOR U34726 ( .A(n34898), .B(n34596), .Z(n34901) );
  XOR U34727 ( .A(n34674), .B(n34902), .Z(n34596) );
  AND U34728 ( .A(n488), .B(n34903), .Z(n34902) );
  XOR U34729 ( .A(n34670), .B(n34674), .Z(n34903) );
  XOR U34730 ( .A(n34545), .B(n34898), .Z(n34900) );
  XOR U34731 ( .A(n34904), .B(n34905), .Z(n34545) );
  AND U34732 ( .A(n504), .B(n34906), .Z(n34905) );
  XOR U34733 ( .A(n34872), .B(n34907), .Z(n34898) );
  AND U34734 ( .A(n34908), .B(n34875), .Z(n34907) );
  XNOR U34735 ( .A(n34606), .B(n34872), .Z(n34875) );
  XOR U34736 ( .A(n34723), .B(n34909), .Z(n34606) );
  AND U34737 ( .A(n488), .B(n34910), .Z(n34909) );
  XOR U34738 ( .A(n34719), .B(n34723), .Z(n34910) );
  XNOR U34739 ( .A(n34911), .B(n34872), .Z(n34908) );
  IV U34740 ( .A(n34553), .Z(n34911) );
  XOR U34741 ( .A(n34912), .B(n34913), .Z(n34553) );
  AND U34742 ( .A(n504), .B(n34914), .Z(n34913) );
  XOR U34743 ( .A(n34915), .B(n34916), .Z(n34872) );
  AND U34744 ( .A(n34917), .B(n34918), .Z(n34916) );
  XNOR U34745 ( .A(n34915), .B(n34614), .Z(n34918) );
  XOR U34746 ( .A(n34816), .B(n34919), .Z(n34614) );
  AND U34747 ( .A(n488), .B(n34920), .Z(n34919) );
  XOR U34748 ( .A(n34812), .B(n34816), .Z(n34920) );
  XNOR U34749 ( .A(n34921), .B(n34915), .Z(n34917) );
  IV U34750 ( .A(n34563), .Z(n34921) );
  XOR U34751 ( .A(n34922), .B(n34923), .Z(n34563) );
  AND U34752 ( .A(n504), .B(n34924), .Z(n34923) );
  AND U34753 ( .A(n34876), .B(n34857), .Z(n34915) );
  XNOR U34754 ( .A(n34925), .B(n34926), .Z(n34857) );
  AND U34755 ( .A(n488), .B(n34835), .Z(n34926) );
  XNOR U34756 ( .A(n34833), .B(n34925), .Z(n34835) );
  XNOR U34757 ( .A(n34927), .B(n34928), .Z(n488) );
  AND U34758 ( .A(n34929), .B(n34930), .Z(n34928) );
  XNOR U34759 ( .A(n34927), .B(n34626), .Z(n34930) );
  IV U34760 ( .A(n34630), .Z(n34626) );
  XOR U34761 ( .A(n34931), .B(n34932), .Z(n34630) );
  AND U34762 ( .A(n492), .B(n34933), .Z(n34932) );
  XOR U34763 ( .A(n34934), .B(n34931), .Z(n34933) );
  XNOR U34764 ( .A(n34927), .B(n34840), .Z(n34929) );
  XOR U34765 ( .A(n34935), .B(n34936), .Z(n34840) );
  AND U34766 ( .A(n500), .B(n34887), .Z(n34936) );
  XOR U34767 ( .A(n34885), .B(n34935), .Z(n34887) );
  XOR U34768 ( .A(n34937), .B(n34938), .Z(n34927) );
  AND U34769 ( .A(n34939), .B(n34940), .Z(n34938) );
  XNOR U34770 ( .A(n34937), .B(n34642), .Z(n34940) );
  IV U34771 ( .A(n34645), .Z(n34642) );
  XOR U34772 ( .A(n34941), .B(n34942), .Z(n34645) );
  AND U34773 ( .A(n492), .B(n34943), .Z(n34942) );
  XOR U34774 ( .A(n34944), .B(n34941), .Z(n34943) );
  XOR U34775 ( .A(n34646), .B(n34937), .Z(n34939) );
  XOR U34776 ( .A(n34945), .B(n34946), .Z(n34646) );
  AND U34777 ( .A(n500), .B(n34897), .Z(n34946) );
  XOR U34778 ( .A(n34945), .B(n34895), .Z(n34897) );
  XOR U34779 ( .A(n34947), .B(n34948), .Z(n34937) );
  AND U34780 ( .A(n34949), .B(n34950), .Z(n34948) );
  XNOR U34781 ( .A(n34947), .B(n34670), .Z(n34950) );
  IV U34782 ( .A(n34673), .Z(n34670) );
  XOR U34783 ( .A(n34951), .B(n34952), .Z(n34673) );
  AND U34784 ( .A(n492), .B(n34953), .Z(n34952) );
  XNOR U34785 ( .A(n34954), .B(n34951), .Z(n34953) );
  XOR U34786 ( .A(n34674), .B(n34947), .Z(n34949) );
  XOR U34787 ( .A(n34955), .B(n34956), .Z(n34674) );
  AND U34788 ( .A(n500), .B(n34906), .Z(n34956) );
  XOR U34789 ( .A(n34955), .B(n34904), .Z(n34906) );
  XOR U34790 ( .A(n34957), .B(n34958), .Z(n34947) );
  AND U34791 ( .A(n34959), .B(n34960), .Z(n34958) );
  XNOR U34792 ( .A(n34957), .B(n34719), .Z(n34960) );
  IV U34793 ( .A(n34722), .Z(n34719) );
  XOR U34794 ( .A(n34961), .B(n34962), .Z(n34722) );
  AND U34795 ( .A(n492), .B(n34963), .Z(n34962) );
  XOR U34796 ( .A(n34964), .B(n34961), .Z(n34963) );
  XOR U34797 ( .A(n34723), .B(n34957), .Z(n34959) );
  XOR U34798 ( .A(n34965), .B(n34966), .Z(n34723) );
  AND U34799 ( .A(n500), .B(n34914), .Z(n34966) );
  XOR U34800 ( .A(n34965), .B(n34912), .Z(n34914) );
  XOR U34801 ( .A(n34853), .B(n34967), .Z(n34957) );
  AND U34802 ( .A(n34855), .B(n34968), .Z(n34967) );
  XNOR U34803 ( .A(n34853), .B(n34812), .Z(n34968) );
  IV U34804 ( .A(n34815), .Z(n34812) );
  XOR U34805 ( .A(n34969), .B(n34970), .Z(n34815) );
  AND U34806 ( .A(n492), .B(n34971), .Z(n34970) );
  XNOR U34807 ( .A(n34972), .B(n34969), .Z(n34971) );
  XOR U34808 ( .A(n34816), .B(n34853), .Z(n34855) );
  XOR U34809 ( .A(n34973), .B(n34974), .Z(n34816) );
  AND U34810 ( .A(n500), .B(n34924), .Z(n34974) );
  XOR U34811 ( .A(n34973), .B(n34922), .Z(n34924) );
  AND U34812 ( .A(n34925), .B(n34833), .Z(n34853) );
  XNOR U34813 ( .A(n34975), .B(n34976), .Z(n34833) );
  AND U34814 ( .A(n492), .B(n34977), .Z(n34976) );
  XNOR U34815 ( .A(n34978), .B(n34975), .Z(n34977) );
  XNOR U34816 ( .A(n34979), .B(n34980), .Z(n492) );
  AND U34817 ( .A(n34981), .B(n34982), .Z(n34980) );
  XOR U34818 ( .A(n34934), .B(n34979), .Z(n34982) );
  AND U34819 ( .A(n34983), .B(n34984), .Z(n34934) );
  XNOR U34820 ( .A(n34931), .B(n34979), .Z(n34981) );
  XNOR U34821 ( .A(n34985), .B(n34986), .Z(n34931) );
  AND U34822 ( .A(n496), .B(n34987), .Z(n34986) );
  XNOR U34823 ( .A(n34988), .B(n34989), .Z(n34987) );
  XOR U34824 ( .A(n34990), .B(n34991), .Z(n34979) );
  AND U34825 ( .A(n34992), .B(n34993), .Z(n34991) );
  XNOR U34826 ( .A(n34990), .B(n34983), .Z(n34993) );
  IV U34827 ( .A(n34944), .Z(n34983) );
  XOR U34828 ( .A(n34994), .B(n34995), .Z(n34944) );
  XOR U34829 ( .A(n34996), .B(n34984), .Z(n34995) );
  AND U34830 ( .A(n34954), .B(n34997), .Z(n34984) );
  AND U34831 ( .A(n34998), .B(n34999), .Z(n34996) );
  XOR U34832 ( .A(n35000), .B(n34994), .Z(n34998) );
  XNOR U34833 ( .A(n34941), .B(n34990), .Z(n34992) );
  XNOR U34834 ( .A(n35001), .B(n35002), .Z(n34941) );
  AND U34835 ( .A(n496), .B(n35003), .Z(n35002) );
  XNOR U34836 ( .A(n35004), .B(n35005), .Z(n35003) );
  XOR U34837 ( .A(n35006), .B(n35007), .Z(n34990) );
  AND U34838 ( .A(n35008), .B(n35009), .Z(n35007) );
  XNOR U34839 ( .A(n35006), .B(n34954), .Z(n35009) );
  XOR U34840 ( .A(n35010), .B(n34999), .Z(n34954) );
  XNOR U34841 ( .A(n35011), .B(n34994), .Z(n34999) );
  XOR U34842 ( .A(n35012), .B(n35013), .Z(n34994) );
  AND U34843 ( .A(n35014), .B(n35015), .Z(n35013) );
  XOR U34844 ( .A(n35016), .B(n35012), .Z(n35014) );
  XNOR U34845 ( .A(n35017), .B(n35018), .Z(n35011) );
  AND U34846 ( .A(n35019), .B(n35020), .Z(n35018) );
  XOR U34847 ( .A(n35017), .B(n35021), .Z(n35019) );
  XNOR U34848 ( .A(n35000), .B(n34997), .Z(n35010) );
  AND U34849 ( .A(n35022), .B(n35023), .Z(n34997) );
  XOR U34850 ( .A(n35024), .B(n35025), .Z(n35000) );
  AND U34851 ( .A(n35026), .B(n35027), .Z(n35025) );
  XOR U34852 ( .A(n35024), .B(n35028), .Z(n35026) );
  XNOR U34853 ( .A(n34951), .B(n35006), .Z(n35008) );
  XNOR U34854 ( .A(n35029), .B(n35030), .Z(n34951) );
  AND U34855 ( .A(n496), .B(n35031), .Z(n35030) );
  XNOR U34856 ( .A(n35032), .B(n35033), .Z(n35031) );
  XOR U34857 ( .A(n35034), .B(n35035), .Z(n35006) );
  AND U34858 ( .A(n35036), .B(n35037), .Z(n35035) );
  XNOR U34859 ( .A(n35034), .B(n35022), .Z(n35037) );
  IV U34860 ( .A(n34964), .Z(n35022) );
  XNOR U34861 ( .A(n35038), .B(n35015), .Z(n34964) );
  XNOR U34862 ( .A(n35039), .B(n35021), .Z(n35015) );
  XOR U34863 ( .A(n35040), .B(n35041), .Z(n35021) );
  AND U34864 ( .A(n35042), .B(n35043), .Z(n35041) );
  XOR U34865 ( .A(n35040), .B(n35044), .Z(n35042) );
  XNOR U34866 ( .A(n35020), .B(n35012), .Z(n35039) );
  XOR U34867 ( .A(n35045), .B(n35046), .Z(n35012) );
  AND U34868 ( .A(n35047), .B(n35048), .Z(n35046) );
  XNOR U34869 ( .A(n35049), .B(n35045), .Z(n35047) );
  XNOR U34870 ( .A(n35050), .B(n35017), .Z(n35020) );
  XOR U34871 ( .A(n35051), .B(n35052), .Z(n35017) );
  AND U34872 ( .A(n35053), .B(n35054), .Z(n35052) );
  XOR U34873 ( .A(n35051), .B(n35055), .Z(n35053) );
  XNOR U34874 ( .A(n35056), .B(n35057), .Z(n35050) );
  AND U34875 ( .A(n35058), .B(n35059), .Z(n35057) );
  XNOR U34876 ( .A(n35056), .B(n35060), .Z(n35058) );
  XNOR U34877 ( .A(n35016), .B(n35023), .Z(n35038) );
  AND U34878 ( .A(n34972), .B(n35061), .Z(n35023) );
  XOR U34879 ( .A(n35028), .B(n35027), .Z(n35016) );
  XNOR U34880 ( .A(n35062), .B(n35024), .Z(n35027) );
  XOR U34881 ( .A(n35063), .B(n35064), .Z(n35024) );
  AND U34882 ( .A(n35065), .B(n35066), .Z(n35064) );
  XOR U34883 ( .A(n35063), .B(n35067), .Z(n35065) );
  XNOR U34884 ( .A(n35068), .B(n35069), .Z(n35062) );
  AND U34885 ( .A(n35070), .B(n35071), .Z(n35069) );
  XOR U34886 ( .A(n35068), .B(n35072), .Z(n35070) );
  XOR U34887 ( .A(n35073), .B(n35074), .Z(n35028) );
  AND U34888 ( .A(n35075), .B(n35076), .Z(n35074) );
  XOR U34889 ( .A(n35073), .B(n35077), .Z(n35075) );
  XNOR U34890 ( .A(n34961), .B(n35034), .Z(n35036) );
  XNOR U34891 ( .A(n35078), .B(n35079), .Z(n34961) );
  AND U34892 ( .A(n496), .B(n35080), .Z(n35079) );
  XNOR U34893 ( .A(n35081), .B(n35082), .Z(n35080) );
  XOR U34894 ( .A(n35083), .B(n35084), .Z(n35034) );
  AND U34895 ( .A(n35085), .B(n35086), .Z(n35084) );
  XNOR U34896 ( .A(n35083), .B(n34972), .Z(n35086) );
  XOR U34897 ( .A(n35087), .B(n35048), .Z(n34972) );
  XNOR U34898 ( .A(n35088), .B(n35055), .Z(n35048) );
  XOR U34899 ( .A(n35044), .B(n35043), .Z(n35055) );
  XNOR U34900 ( .A(n35089), .B(n35040), .Z(n35043) );
  XOR U34901 ( .A(n35090), .B(n35091), .Z(n35040) );
  AND U34902 ( .A(n35092), .B(n35093), .Z(n35091) );
  XOR U34903 ( .A(n35090), .B(n35094), .Z(n35092) );
  XNOR U34904 ( .A(n35095), .B(n35096), .Z(n35089) );
  NOR U34905 ( .A(n35097), .B(n35098), .Z(n35096) );
  XNOR U34906 ( .A(n35095), .B(n35099), .Z(n35097) );
  XOR U34907 ( .A(n35100), .B(n35101), .Z(n35044) );
  NOR U34908 ( .A(n35102), .B(n35103), .Z(n35101) );
  XNOR U34909 ( .A(n35100), .B(n35104), .Z(n35102) );
  XNOR U34910 ( .A(n35054), .B(n35045), .Z(n35088) );
  XOR U34911 ( .A(n35105), .B(n35106), .Z(n35045) );
  NOR U34912 ( .A(n35107), .B(n35108), .Z(n35106) );
  XNOR U34913 ( .A(n35105), .B(n35109), .Z(n35107) );
  XOR U34914 ( .A(n35110), .B(n35060), .Z(n35054) );
  XNOR U34915 ( .A(n35111), .B(n35112), .Z(n35060) );
  NOR U34916 ( .A(n35113), .B(n35114), .Z(n35112) );
  XNOR U34917 ( .A(n35111), .B(n35115), .Z(n35113) );
  XNOR U34918 ( .A(n35059), .B(n35051), .Z(n35110) );
  XOR U34919 ( .A(n35116), .B(n35117), .Z(n35051) );
  AND U34920 ( .A(n35118), .B(n35119), .Z(n35117) );
  XOR U34921 ( .A(n35116), .B(n35120), .Z(n35118) );
  XNOR U34922 ( .A(n35121), .B(n35056), .Z(n35059) );
  XOR U34923 ( .A(n35122), .B(n35123), .Z(n35056) );
  AND U34924 ( .A(n35124), .B(n35125), .Z(n35123) );
  XOR U34925 ( .A(n35122), .B(n35126), .Z(n35124) );
  XNOR U34926 ( .A(n35127), .B(n35128), .Z(n35121) );
  NOR U34927 ( .A(n35129), .B(n35130), .Z(n35128) );
  XOR U34928 ( .A(n35127), .B(n35131), .Z(n35129) );
  XOR U34929 ( .A(n35049), .B(n35061), .Z(n35087) );
  NOR U34930 ( .A(n34978), .B(n35132), .Z(n35061) );
  XNOR U34931 ( .A(n35067), .B(n35066), .Z(n35049) );
  XNOR U34932 ( .A(n35133), .B(n35072), .Z(n35066) );
  XOR U34933 ( .A(n35134), .B(n35135), .Z(n35072) );
  NOR U34934 ( .A(n35136), .B(n35137), .Z(n35135) );
  XNOR U34935 ( .A(n35134), .B(n35138), .Z(n35136) );
  XNOR U34936 ( .A(n35071), .B(n35063), .Z(n35133) );
  XOR U34937 ( .A(n35139), .B(n35140), .Z(n35063) );
  AND U34938 ( .A(n35141), .B(n35142), .Z(n35140) );
  XNOR U34939 ( .A(n35139), .B(n35143), .Z(n35141) );
  XNOR U34940 ( .A(n35144), .B(n35068), .Z(n35071) );
  XOR U34941 ( .A(n35145), .B(n35146), .Z(n35068) );
  AND U34942 ( .A(n35147), .B(n35148), .Z(n35146) );
  XOR U34943 ( .A(n35145), .B(n35149), .Z(n35147) );
  XNOR U34944 ( .A(n35150), .B(n35151), .Z(n35144) );
  NOR U34945 ( .A(n35152), .B(n35153), .Z(n35151) );
  XOR U34946 ( .A(n35150), .B(n35154), .Z(n35152) );
  XOR U34947 ( .A(n35077), .B(n35076), .Z(n35067) );
  XNOR U34948 ( .A(n35155), .B(n35073), .Z(n35076) );
  XOR U34949 ( .A(n35156), .B(n35157), .Z(n35073) );
  AND U34950 ( .A(n35158), .B(n35159), .Z(n35157) );
  XOR U34951 ( .A(n35156), .B(n35160), .Z(n35158) );
  XNOR U34952 ( .A(n35161), .B(n35162), .Z(n35155) );
  NOR U34953 ( .A(n35163), .B(n35164), .Z(n35162) );
  XNOR U34954 ( .A(n35161), .B(n35165), .Z(n35163) );
  XOR U34955 ( .A(n35166), .B(n35167), .Z(n35077) );
  NOR U34956 ( .A(n35168), .B(n35169), .Z(n35167) );
  XNOR U34957 ( .A(n35166), .B(n35170), .Z(n35168) );
  XNOR U34958 ( .A(n34969), .B(n35083), .Z(n35085) );
  XNOR U34959 ( .A(n35171), .B(n35172), .Z(n34969) );
  AND U34960 ( .A(n496), .B(n35173), .Z(n35172) );
  XNOR U34961 ( .A(n35174), .B(n35175), .Z(n35173) );
  AND U34962 ( .A(n34975), .B(n34978), .Z(n35083) );
  XOR U34963 ( .A(n35176), .B(n35132), .Z(n34978) );
  XNOR U34964 ( .A(p_input[2048]), .B(p_input[608]), .Z(n35132) );
  XOR U34965 ( .A(n35109), .B(n35108), .Z(n35176) );
  XOR U34966 ( .A(n35177), .B(n35120), .Z(n35108) );
  XOR U34967 ( .A(n35094), .B(n35093), .Z(n35120) );
  XNOR U34968 ( .A(n35178), .B(n35099), .Z(n35093) );
  XOR U34969 ( .A(p_input[2072]), .B(p_input[632]), .Z(n35099) );
  XOR U34970 ( .A(n35090), .B(n35098), .Z(n35178) );
  XOR U34971 ( .A(n35179), .B(n35095), .Z(n35098) );
  XOR U34972 ( .A(p_input[2070]), .B(p_input[630]), .Z(n35095) );
  XNOR U34973 ( .A(p_input[2071]), .B(p_input[631]), .Z(n35179) );
  XNOR U34974 ( .A(n28684), .B(p_input[626]), .Z(n35090) );
  XNOR U34975 ( .A(n35104), .B(n35103), .Z(n35094) );
  XOR U34976 ( .A(n35180), .B(n35100), .Z(n35103) );
  XOR U34977 ( .A(p_input[2067]), .B(p_input[627]), .Z(n35100) );
  XNOR U34978 ( .A(p_input[2068]), .B(p_input[628]), .Z(n35180) );
  XOR U34979 ( .A(p_input[2069]), .B(p_input[629]), .Z(n35104) );
  XNOR U34980 ( .A(n35119), .B(n35105), .Z(n35177) );
  XNOR U34981 ( .A(n28686), .B(p_input[609]), .Z(n35105) );
  XNOR U34982 ( .A(n35181), .B(n35126), .Z(n35119) );
  XNOR U34983 ( .A(n35115), .B(n35114), .Z(n35126) );
  XOR U34984 ( .A(n35182), .B(n35111), .Z(n35114) );
  XNOR U34985 ( .A(n28322), .B(p_input[634]), .Z(n35111) );
  XNOR U34986 ( .A(p_input[2075]), .B(p_input[635]), .Z(n35182) );
  XOR U34987 ( .A(p_input[2076]), .B(p_input[636]), .Z(n35115) );
  XNOR U34988 ( .A(n35125), .B(n35116), .Z(n35181) );
  XNOR U34989 ( .A(n28689), .B(p_input[625]), .Z(n35116) );
  XOR U34990 ( .A(n35183), .B(n35131), .Z(n35125) );
  XNOR U34991 ( .A(p_input[2079]), .B(p_input[639]), .Z(n35131) );
  XOR U34992 ( .A(n35122), .B(n35130), .Z(n35183) );
  XOR U34993 ( .A(n35184), .B(n35127), .Z(n35130) );
  XOR U34994 ( .A(p_input[2077]), .B(p_input[637]), .Z(n35127) );
  XNOR U34995 ( .A(p_input[2078]), .B(p_input[638]), .Z(n35184) );
  XNOR U34996 ( .A(n28326), .B(p_input[633]), .Z(n35122) );
  XNOR U34997 ( .A(n35143), .B(n35142), .Z(n35109) );
  XNOR U34998 ( .A(n35185), .B(n35149), .Z(n35142) );
  XNOR U34999 ( .A(n35138), .B(n35137), .Z(n35149) );
  XOR U35000 ( .A(n35186), .B(n35134), .Z(n35137) );
  XNOR U35001 ( .A(n28694), .B(p_input[619]), .Z(n35134) );
  XNOR U35002 ( .A(p_input[2060]), .B(p_input[620]), .Z(n35186) );
  XOR U35003 ( .A(p_input[2061]), .B(p_input[621]), .Z(n35138) );
  XNOR U35004 ( .A(n35148), .B(n35139), .Z(n35185) );
  XNOR U35005 ( .A(n28330), .B(p_input[610]), .Z(n35139) );
  XOR U35006 ( .A(n35187), .B(n35154), .Z(n35148) );
  XNOR U35007 ( .A(p_input[2064]), .B(p_input[624]), .Z(n35154) );
  XOR U35008 ( .A(n35145), .B(n35153), .Z(n35187) );
  XOR U35009 ( .A(n35188), .B(n35150), .Z(n35153) );
  XOR U35010 ( .A(p_input[2062]), .B(p_input[622]), .Z(n35150) );
  XNOR U35011 ( .A(p_input[2063]), .B(p_input[623]), .Z(n35188) );
  XNOR U35012 ( .A(n28697), .B(p_input[618]), .Z(n35145) );
  XNOR U35013 ( .A(n35160), .B(n35159), .Z(n35143) );
  XNOR U35014 ( .A(n35189), .B(n35165), .Z(n35159) );
  XOR U35015 ( .A(p_input[2057]), .B(p_input[617]), .Z(n35165) );
  XOR U35016 ( .A(n35156), .B(n35164), .Z(n35189) );
  XOR U35017 ( .A(n35190), .B(n35161), .Z(n35164) );
  XOR U35018 ( .A(p_input[2055]), .B(p_input[615]), .Z(n35161) );
  XNOR U35019 ( .A(p_input[2056]), .B(p_input[616]), .Z(n35190) );
  XNOR U35020 ( .A(n28337), .B(p_input[611]), .Z(n35156) );
  XNOR U35021 ( .A(n35170), .B(n35169), .Z(n35160) );
  XOR U35022 ( .A(n35191), .B(n35166), .Z(n35169) );
  XOR U35023 ( .A(p_input[2052]), .B(p_input[612]), .Z(n35166) );
  XNOR U35024 ( .A(p_input[2053]), .B(p_input[613]), .Z(n35191) );
  XOR U35025 ( .A(p_input[2054]), .B(p_input[614]), .Z(n35170) );
  XNOR U35026 ( .A(n35192), .B(n35193), .Z(n34975) );
  AND U35027 ( .A(n496), .B(n35194), .Z(n35193) );
  XNOR U35028 ( .A(n35195), .B(n35196), .Z(n496) );
  AND U35029 ( .A(n35197), .B(n35198), .Z(n35196) );
  XOR U35030 ( .A(n34989), .B(n35195), .Z(n35198) );
  XNOR U35031 ( .A(n35199), .B(n35195), .Z(n35197) );
  XOR U35032 ( .A(n35200), .B(n35201), .Z(n35195) );
  AND U35033 ( .A(n35202), .B(n35203), .Z(n35201) );
  XOR U35034 ( .A(n35004), .B(n35200), .Z(n35203) );
  XOR U35035 ( .A(n35200), .B(n35005), .Z(n35202) );
  XOR U35036 ( .A(n35204), .B(n35205), .Z(n35200) );
  AND U35037 ( .A(n35206), .B(n35207), .Z(n35205) );
  XOR U35038 ( .A(n35032), .B(n35204), .Z(n35207) );
  XOR U35039 ( .A(n35204), .B(n35033), .Z(n35206) );
  XOR U35040 ( .A(n35208), .B(n35209), .Z(n35204) );
  AND U35041 ( .A(n35210), .B(n35211), .Z(n35209) );
  XOR U35042 ( .A(n35081), .B(n35208), .Z(n35211) );
  XOR U35043 ( .A(n35208), .B(n35082), .Z(n35210) );
  XOR U35044 ( .A(n35212), .B(n35213), .Z(n35208) );
  AND U35045 ( .A(n35214), .B(n35215), .Z(n35213) );
  XOR U35046 ( .A(n35212), .B(n35174), .Z(n35215) );
  XNOR U35047 ( .A(n35216), .B(n35217), .Z(n34925) );
  AND U35048 ( .A(n500), .B(n35218), .Z(n35217) );
  XNOR U35049 ( .A(n35219), .B(n35220), .Z(n500) );
  AND U35050 ( .A(n35221), .B(n35222), .Z(n35220) );
  XOR U35051 ( .A(n35219), .B(n34935), .Z(n35222) );
  XNOR U35052 ( .A(n35219), .B(n34885), .Z(n35221) );
  XOR U35053 ( .A(n35223), .B(n35224), .Z(n35219) );
  AND U35054 ( .A(n35225), .B(n35226), .Z(n35224) );
  XNOR U35055 ( .A(n34945), .B(n35223), .Z(n35226) );
  XOR U35056 ( .A(n35223), .B(n34895), .Z(n35225) );
  XOR U35057 ( .A(n35227), .B(n35228), .Z(n35223) );
  AND U35058 ( .A(n35229), .B(n35230), .Z(n35228) );
  XNOR U35059 ( .A(n34955), .B(n35227), .Z(n35230) );
  XOR U35060 ( .A(n35227), .B(n34904), .Z(n35229) );
  XOR U35061 ( .A(n35231), .B(n35232), .Z(n35227) );
  AND U35062 ( .A(n35233), .B(n35234), .Z(n35232) );
  XOR U35063 ( .A(n35231), .B(n34912), .Z(n35233) );
  XOR U35064 ( .A(n35235), .B(n35236), .Z(n34876) );
  AND U35065 ( .A(n504), .B(n35218), .Z(n35236) );
  XNOR U35066 ( .A(n35216), .B(n35235), .Z(n35218) );
  XNOR U35067 ( .A(n35237), .B(n35238), .Z(n504) );
  AND U35068 ( .A(n35239), .B(n35240), .Z(n35238) );
  XNOR U35069 ( .A(n35241), .B(n35237), .Z(n35240) );
  IV U35070 ( .A(n34935), .Z(n35241) );
  XOR U35071 ( .A(n35199), .B(n35242), .Z(n34935) );
  AND U35072 ( .A(n507), .B(n35243), .Z(n35242) );
  XOR U35073 ( .A(n34988), .B(n34985), .Z(n35243) );
  IV U35074 ( .A(n35199), .Z(n34988) );
  XNOR U35075 ( .A(n34885), .B(n35237), .Z(n35239) );
  XOR U35076 ( .A(n35244), .B(n35245), .Z(n34885) );
  AND U35077 ( .A(n523), .B(n35246), .Z(n35245) );
  XOR U35078 ( .A(n35247), .B(n35248), .Z(n35237) );
  AND U35079 ( .A(n35249), .B(n35250), .Z(n35248) );
  XNOR U35080 ( .A(n35247), .B(n34945), .Z(n35250) );
  XOR U35081 ( .A(n35005), .B(n35251), .Z(n34945) );
  AND U35082 ( .A(n507), .B(n35252), .Z(n35251) );
  XOR U35083 ( .A(n35001), .B(n35005), .Z(n35252) );
  XNOR U35084 ( .A(n35253), .B(n35247), .Z(n35249) );
  IV U35085 ( .A(n34895), .Z(n35253) );
  XOR U35086 ( .A(n35254), .B(n35255), .Z(n34895) );
  AND U35087 ( .A(n523), .B(n35256), .Z(n35255) );
  XOR U35088 ( .A(n35257), .B(n35258), .Z(n35247) );
  AND U35089 ( .A(n35259), .B(n35260), .Z(n35258) );
  XNOR U35090 ( .A(n35257), .B(n34955), .Z(n35260) );
  XOR U35091 ( .A(n35033), .B(n35261), .Z(n34955) );
  AND U35092 ( .A(n507), .B(n35262), .Z(n35261) );
  XOR U35093 ( .A(n35029), .B(n35033), .Z(n35262) );
  XOR U35094 ( .A(n34904), .B(n35257), .Z(n35259) );
  XOR U35095 ( .A(n35263), .B(n35264), .Z(n34904) );
  AND U35096 ( .A(n523), .B(n35265), .Z(n35264) );
  XOR U35097 ( .A(n35231), .B(n35266), .Z(n35257) );
  AND U35098 ( .A(n35267), .B(n35234), .Z(n35266) );
  XNOR U35099 ( .A(n34965), .B(n35231), .Z(n35234) );
  XOR U35100 ( .A(n35082), .B(n35268), .Z(n34965) );
  AND U35101 ( .A(n507), .B(n35269), .Z(n35268) );
  XOR U35102 ( .A(n35078), .B(n35082), .Z(n35269) );
  XNOR U35103 ( .A(n35270), .B(n35231), .Z(n35267) );
  IV U35104 ( .A(n34912), .Z(n35270) );
  XOR U35105 ( .A(n35271), .B(n35272), .Z(n34912) );
  AND U35106 ( .A(n523), .B(n35273), .Z(n35272) );
  XOR U35107 ( .A(n35274), .B(n35275), .Z(n35231) );
  AND U35108 ( .A(n35276), .B(n35277), .Z(n35275) );
  XNOR U35109 ( .A(n35274), .B(n34973), .Z(n35277) );
  XOR U35110 ( .A(n35175), .B(n35278), .Z(n34973) );
  AND U35111 ( .A(n507), .B(n35279), .Z(n35278) );
  XOR U35112 ( .A(n35171), .B(n35175), .Z(n35279) );
  XNOR U35113 ( .A(n35280), .B(n35274), .Z(n35276) );
  IV U35114 ( .A(n34922), .Z(n35280) );
  XOR U35115 ( .A(n35281), .B(n35282), .Z(n34922) );
  AND U35116 ( .A(n523), .B(n35283), .Z(n35282) );
  AND U35117 ( .A(n35235), .B(n35216), .Z(n35274) );
  XNOR U35118 ( .A(n35284), .B(n35285), .Z(n35216) );
  AND U35119 ( .A(n507), .B(n35194), .Z(n35285) );
  XNOR U35120 ( .A(n35192), .B(n35284), .Z(n35194) );
  XNOR U35121 ( .A(n35286), .B(n35287), .Z(n507) );
  AND U35122 ( .A(n35288), .B(n35289), .Z(n35287) );
  XNOR U35123 ( .A(n35286), .B(n34985), .Z(n35289) );
  IV U35124 ( .A(n34989), .Z(n34985) );
  XOR U35125 ( .A(n35290), .B(n35291), .Z(n34989) );
  AND U35126 ( .A(n511), .B(n35292), .Z(n35291) );
  XOR U35127 ( .A(n35293), .B(n35290), .Z(n35292) );
  XNOR U35128 ( .A(n35286), .B(n35199), .Z(n35288) );
  XOR U35129 ( .A(n35294), .B(n35295), .Z(n35199) );
  AND U35130 ( .A(n519), .B(n35246), .Z(n35295) );
  XOR U35131 ( .A(n35244), .B(n35294), .Z(n35246) );
  XOR U35132 ( .A(n35296), .B(n35297), .Z(n35286) );
  AND U35133 ( .A(n35298), .B(n35299), .Z(n35297) );
  XNOR U35134 ( .A(n35296), .B(n35001), .Z(n35299) );
  IV U35135 ( .A(n35004), .Z(n35001) );
  XOR U35136 ( .A(n35300), .B(n35301), .Z(n35004) );
  AND U35137 ( .A(n511), .B(n35302), .Z(n35301) );
  XOR U35138 ( .A(n35303), .B(n35300), .Z(n35302) );
  XOR U35139 ( .A(n35005), .B(n35296), .Z(n35298) );
  XOR U35140 ( .A(n35304), .B(n35305), .Z(n35005) );
  AND U35141 ( .A(n519), .B(n35256), .Z(n35305) );
  XOR U35142 ( .A(n35304), .B(n35254), .Z(n35256) );
  XOR U35143 ( .A(n35306), .B(n35307), .Z(n35296) );
  AND U35144 ( .A(n35308), .B(n35309), .Z(n35307) );
  XNOR U35145 ( .A(n35306), .B(n35029), .Z(n35309) );
  IV U35146 ( .A(n35032), .Z(n35029) );
  XOR U35147 ( .A(n35310), .B(n35311), .Z(n35032) );
  AND U35148 ( .A(n511), .B(n35312), .Z(n35311) );
  XNOR U35149 ( .A(n35313), .B(n35310), .Z(n35312) );
  XOR U35150 ( .A(n35033), .B(n35306), .Z(n35308) );
  XOR U35151 ( .A(n35314), .B(n35315), .Z(n35033) );
  AND U35152 ( .A(n519), .B(n35265), .Z(n35315) );
  XOR U35153 ( .A(n35314), .B(n35263), .Z(n35265) );
  XOR U35154 ( .A(n35316), .B(n35317), .Z(n35306) );
  AND U35155 ( .A(n35318), .B(n35319), .Z(n35317) );
  XNOR U35156 ( .A(n35316), .B(n35078), .Z(n35319) );
  IV U35157 ( .A(n35081), .Z(n35078) );
  XOR U35158 ( .A(n35320), .B(n35321), .Z(n35081) );
  AND U35159 ( .A(n511), .B(n35322), .Z(n35321) );
  XOR U35160 ( .A(n35323), .B(n35320), .Z(n35322) );
  XOR U35161 ( .A(n35082), .B(n35316), .Z(n35318) );
  XOR U35162 ( .A(n35324), .B(n35325), .Z(n35082) );
  AND U35163 ( .A(n519), .B(n35273), .Z(n35325) );
  XOR U35164 ( .A(n35324), .B(n35271), .Z(n35273) );
  XOR U35165 ( .A(n35212), .B(n35326), .Z(n35316) );
  AND U35166 ( .A(n35214), .B(n35327), .Z(n35326) );
  XNOR U35167 ( .A(n35212), .B(n35171), .Z(n35327) );
  IV U35168 ( .A(n35174), .Z(n35171) );
  XOR U35169 ( .A(n35328), .B(n35329), .Z(n35174) );
  AND U35170 ( .A(n511), .B(n35330), .Z(n35329) );
  XNOR U35171 ( .A(n35331), .B(n35328), .Z(n35330) );
  XOR U35172 ( .A(n35175), .B(n35212), .Z(n35214) );
  XOR U35173 ( .A(n35332), .B(n35333), .Z(n35175) );
  AND U35174 ( .A(n519), .B(n35283), .Z(n35333) );
  XOR U35175 ( .A(n35332), .B(n35281), .Z(n35283) );
  AND U35176 ( .A(n35284), .B(n35192), .Z(n35212) );
  XNOR U35177 ( .A(n35334), .B(n35335), .Z(n35192) );
  AND U35178 ( .A(n511), .B(n35336), .Z(n35335) );
  XNOR U35179 ( .A(n35337), .B(n35334), .Z(n35336) );
  XNOR U35180 ( .A(n35338), .B(n35339), .Z(n511) );
  AND U35181 ( .A(n35340), .B(n35341), .Z(n35339) );
  XOR U35182 ( .A(n35293), .B(n35338), .Z(n35341) );
  AND U35183 ( .A(n35342), .B(n35343), .Z(n35293) );
  XNOR U35184 ( .A(n35290), .B(n35338), .Z(n35340) );
  XNOR U35185 ( .A(n35344), .B(n35345), .Z(n35290) );
  AND U35186 ( .A(n515), .B(n35346), .Z(n35345) );
  XNOR U35187 ( .A(n35347), .B(n35348), .Z(n35346) );
  XOR U35188 ( .A(n35349), .B(n35350), .Z(n35338) );
  AND U35189 ( .A(n35351), .B(n35352), .Z(n35350) );
  XNOR U35190 ( .A(n35349), .B(n35342), .Z(n35352) );
  IV U35191 ( .A(n35303), .Z(n35342) );
  XOR U35192 ( .A(n35353), .B(n35354), .Z(n35303) );
  XOR U35193 ( .A(n35355), .B(n35343), .Z(n35354) );
  AND U35194 ( .A(n35313), .B(n35356), .Z(n35343) );
  AND U35195 ( .A(n35357), .B(n35358), .Z(n35355) );
  XOR U35196 ( .A(n35359), .B(n35353), .Z(n35357) );
  XNOR U35197 ( .A(n35300), .B(n35349), .Z(n35351) );
  XNOR U35198 ( .A(n35360), .B(n35361), .Z(n35300) );
  AND U35199 ( .A(n515), .B(n35362), .Z(n35361) );
  XNOR U35200 ( .A(n35363), .B(n35364), .Z(n35362) );
  XOR U35201 ( .A(n35365), .B(n35366), .Z(n35349) );
  AND U35202 ( .A(n35367), .B(n35368), .Z(n35366) );
  XNOR U35203 ( .A(n35365), .B(n35313), .Z(n35368) );
  XOR U35204 ( .A(n35369), .B(n35358), .Z(n35313) );
  XNOR U35205 ( .A(n35370), .B(n35353), .Z(n35358) );
  XOR U35206 ( .A(n35371), .B(n35372), .Z(n35353) );
  AND U35207 ( .A(n35373), .B(n35374), .Z(n35372) );
  XOR U35208 ( .A(n35375), .B(n35371), .Z(n35373) );
  XNOR U35209 ( .A(n35376), .B(n35377), .Z(n35370) );
  AND U35210 ( .A(n35378), .B(n35379), .Z(n35377) );
  XOR U35211 ( .A(n35376), .B(n35380), .Z(n35378) );
  XNOR U35212 ( .A(n35359), .B(n35356), .Z(n35369) );
  AND U35213 ( .A(n35381), .B(n35382), .Z(n35356) );
  XOR U35214 ( .A(n35383), .B(n35384), .Z(n35359) );
  AND U35215 ( .A(n35385), .B(n35386), .Z(n35384) );
  XOR U35216 ( .A(n35383), .B(n35387), .Z(n35385) );
  XNOR U35217 ( .A(n35310), .B(n35365), .Z(n35367) );
  XNOR U35218 ( .A(n35388), .B(n35389), .Z(n35310) );
  AND U35219 ( .A(n515), .B(n35390), .Z(n35389) );
  XNOR U35220 ( .A(n35391), .B(n35392), .Z(n35390) );
  XOR U35221 ( .A(n35393), .B(n35394), .Z(n35365) );
  AND U35222 ( .A(n35395), .B(n35396), .Z(n35394) );
  XNOR U35223 ( .A(n35393), .B(n35381), .Z(n35396) );
  IV U35224 ( .A(n35323), .Z(n35381) );
  XNOR U35225 ( .A(n35397), .B(n35374), .Z(n35323) );
  XNOR U35226 ( .A(n35398), .B(n35380), .Z(n35374) );
  XOR U35227 ( .A(n35399), .B(n35400), .Z(n35380) );
  AND U35228 ( .A(n35401), .B(n35402), .Z(n35400) );
  XOR U35229 ( .A(n35399), .B(n35403), .Z(n35401) );
  XNOR U35230 ( .A(n35379), .B(n35371), .Z(n35398) );
  XOR U35231 ( .A(n35404), .B(n35405), .Z(n35371) );
  AND U35232 ( .A(n35406), .B(n35407), .Z(n35405) );
  XNOR U35233 ( .A(n35408), .B(n35404), .Z(n35406) );
  XNOR U35234 ( .A(n35409), .B(n35376), .Z(n35379) );
  XOR U35235 ( .A(n35410), .B(n35411), .Z(n35376) );
  AND U35236 ( .A(n35412), .B(n35413), .Z(n35411) );
  XOR U35237 ( .A(n35410), .B(n35414), .Z(n35412) );
  XNOR U35238 ( .A(n35415), .B(n35416), .Z(n35409) );
  AND U35239 ( .A(n35417), .B(n35418), .Z(n35416) );
  XNOR U35240 ( .A(n35415), .B(n35419), .Z(n35417) );
  XNOR U35241 ( .A(n35375), .B(n35382), .Z(n35397) );
  AND U35242 ( .A(n35331), .B(n35420), .Z(n35382) );
  XOR U35243 ( .A(n35387), .B(n35386), .Z(n35375) );
  XNOR U35244 ( .A(n35421), .B(n35383), .Z(n35386) );
  XOR U35245 ( .A(n35422), .B(n35423), .Z(n35383) );
  AND U35246 ( .A(n35424), .B(n35425), .Z(n35423) );
  XOR U35247 ( .A(n35422), .B(n35426), .Z(n35424) );
  XNOR U35248 ( .A(n35427), .B(n35428), .Z(n35421) );
  AND U35249 ( .A(n35429), .B(n35430), .Z(n35428) );
  XOR U35250 ( .A(n35427), .B(n35431), .Z(n35429) );
  XOR U35251 ( .A(n35432), .B(n35433), .Z(n35387) );
  AND U35252 ( .A(n35434), .B(n35435), .Z(n35433) );
  XOR U35253 ( .A(n35432), .B(n35436), .Z(n35434) );
  XNOR U35254 ( .A(n35320), .B(n35393), .Z(n35395) );
  XNOR U35255 ( .A(n35437), .B(n35438), .Z(n35320) );
  AND U35256 ( .A(n515), .B(n35439), .Z(n35438) );
  XNOR U35257 ( .A(n35440), .B(n35441), .Z(n35439) );
  XOR U35258 ( .A(n35442), .B(n35443), .Z(n35393) );
  AND U35259 ( .A(n35444), .B(n35445), .Z(n35443) );
  XNOR U35260 ( .A(n35442), .B(n35331), .Z(n35445) );
  XOR U35261 ( .A(n35446), .B(n35407), .Z(n35331) );
  XNOR U35262 ( .A(n35447), .B(n35414), .Z(n35407) );
  XOR U35263 ( .A(n35403), .B(n35402), .Z(n35414) );
  XNOR U35264 ( .A(n35448), .B(n35399), .Z(n35402) );
  XOR U35265 ( .A(n35449), .B(n35450), .Z(n35399) );
  AND U35266 ( .A(n35451), .B(n35452), .Z(n35450) );
  XOR U35267 ( .A(n35449), .B(n35453), .Z(n35451) );
  XNOR U35268 ( .A(n35454), .B(n35455), .Z(n35448) );
  NOR U35269 ( .A(n35456), .B(n35457), .Z(n35455) );
  XNOR U35270 ( .A(n35454), .B(n35458), .Z(n35456) );
  XOR U35271 ( .A(n35459), .B(n35460), .Z(n35403) );
  NOR U35272 ( .A(n35461), .B(n35462), .Z(n35460) );
  XNOR U35273 ( .A(n35459), .B(n35463), .Z(n35461) );
  XNOR U35274 ( .A(n35413), .B(n35404), .Z(n35447) );
  XOR U35275 ( .A(n35464), .B(n35465), .Z(n35404) );
  NOR U35276 ( .A(n35466), .B(n35467), .Z(n35465) );
  XNOR U35277 ( .A(n35464), .B(n35468), .Z(n35466) );
  XOR U35278 ( .A(n35469), .B(n35419), .Z(n35413) );
  XNOR U35279 ( .A(n35470), .B(n35471), .Z(n35419) );
  NOR U35280 ( .A(n35472), .B(n35473), .Z(n35471) );
  XNOR U35281 ( .A(n35470), .B(n35474), .Z(n35472) );
  XNOR U35282 ( .A(n35418), .B(n35410), .Z(n35469) );
  XOR U35283 ( .A(n35475), .B(n35476), .Z(n35410) );
  AND U35284 ( .A(n35477), .B(n35478), .Z(n35476) );
  XOR U35285 ( .A(n35475), .B(n35479), .Z(n35477) );
  XNOR U35286 ( .A(n35480), .B(n35415), .Z(n35418) );
  XOR U35287 ( .A(n35481), .B(n35482), .Z(n35415) );
  AND U35288 ( .A(n35483), .B(n35484), .Z(n35482) );
  XOR U35289 ( .A(n35481), .B(n35485), .Z(n35483) );
  XNOR U35290 ( .A(n35486), .B(n35487), .Z(n35480) );
  NOR U35291 ( .A(n35488), .B(n35489), .Z(n35487) );
  XOR U35292 ( .A(n35486), .B(n35490), .Z(n35488) );
  XOR U35293 ( .A(n35408), .B(n35420), .Z(n35446) );
  NOR U35294 ( .A(n35337), .B(n35491), .Z(n35420) );
  XNOR U35295 ( .A(n35426), .B(n35425), .Z(n35408) );
  XNOR U35296 ( .A(n35492), .B(n35431), .Z(n35425) );
  XOR U35297 ( .A(n35493), .B(n35494), .Z(n35431) );
  NOR U35298 ( .A(n35495), .B(n35496), .Z(n35494) );
  XNOR U35299 ( .A(n35493), .B(n35497), .Z(n35495) );
  XNOR U35300 ( .A(n35430), .B(n35422), .Z(n35492) );
  XOR U35301 ( .A(n35498), .B(n35499), .Z(n35422) );
  AND U35302 ( .A(n35500), .B(n35501), .Z(n35499) );
  XNOR U35303 ( .A(n35498), .B(n35502), .Z(n35500) );
  XNOR U35304 ( .A(n35503), .B(n35427), .Z(n35430) );
  XOR U35305 ( .A(n35504), .B(n35505), .Z(n35427) );
  AND U35306 ( .A(n35506), .B(n35507), .Z(n35505) );
  XOR U35307 ( .A(n35504), .B(n35508), .Z(n35506) );
  XNOR U35308 ( .A(n35509), .B(n35510), .Z(n35503) );
  NOR U35309 ( .A(n35511), .B(n35512), .Z(n35510) );
  XOR U35310 ( .A(n35509), .B(n35513), .Z(n35511) );
  XOR U35311 ( .A(n35436), .B(n35435), .Z(n35426) );
  XNOR U35312 ( .A(n35514), .B(n35432), .Z(n35435) );
  XOR U35313 ( .A(n35515), .B(n35516), .Z(n35432) );
  AND U35314 ( .A(n35517), .B(n35518), .Z(n35516) );
  XOR U35315 ( .A(n35515), .B(n35519), .Z(n35517) );
  XNOR U35316 ( .A(n35520), .B(n35521), .Z(n35514) );
  NOR U35317 ( .A(n35522), .B(n35523), .Z(n35521) );
  XNOR U35318 ( .A(n35520), .B(n35524), .Z(n35522) );
  XOR U35319 ( .A(n35525), .B(n35526), .Z(n35436) );
  NOR U35320 ( .A(n35527), .B(n35528), .Z(n35526) );
  XNOR U35321 ( .A(n35525), .B(n35529), .Z(n35527) );
  XNOR U35322 ( .A(n35328), .B(n35442), .Z(n35444) );
  XNOR U35323 ( .A(n35530), .B(n35531), .Z(n35328) );
  AND U35324 ( .A(n515), .B(n35532), .Z(n35531) );
  XNOR U35325 ( .A(n35533), .B(n35534), .Z(n35532) );
  AND U35326 ( .A(n35334), .B(n35337), .Z(n35442) );
  XOR U35327 ( .A(n35535), .B(n35491), .Z(n35337) );
  XNOR U35328 ( .A(p_input[2048]), .B(p_input[640]), .Z(n35491) );
  XOR U35329 ( .A(n35468), .B(n35467), .Z(n35535) );
  XOR U35330 ( .A(n35536), .B(n35479), .Z(n35467) );
  XOR U35331 ( .A(n35453), .B(n35452), .Z(n35479) );
  XNOR U35332 ( .A(n35537), .B(n35458), .Z(n35452) );
  XOR U35333 ( .A(p_input[2072]), .B(p_input[664]), .Z(n35458) );
  XOR U35334 ( .A(n35449), .B(n35457), .Z(n35537) );
  XOR U35335 ( .A(n35538), .B(n35454), .Z(n35457) );
  XOR U35336 ( .A(p_input[2070]), .B(p_input[662]), .Z(n35454) );
  XNOR U35337 ( .A(p_input[2071]), .B(p_input[663]), .Z(n35538) );
  XNOR U35338 ( .A(n28684), .B(p_input[658]), .Z(n35449) );
  XNOR U35339 ( .A(n35463), .B(n35462), .Z(n35453) );
  XOR U35340 ( .A(n35539), .B(n35459), .Z(n35462) );
  XOR U35341 ( .A(p_input[2067]), .B(p_input[659]), .Z(n35459) );
  XNOR U35342 ( .A(p_input[2068]), .B(p_input[660]), .Z(n35539) );
  XOR U35343 ( .A(p_input[2069]), .B(p_input[661]), .Z(n35463) );
  XNOR U35344 ( .A(n35478), .B(n35464), .Z(n35536) );
  XNOR U35345 ( .A(n28686), .B(p_input[641]), .Z(n35464) );
  XNOR U35346 ( .A(n35540), .B(n35485), .Z(n35478) );
  XNOR U35347 ( .A(n35474), .B(n35473), .Z(n35485) );
  XOR U35348 ( .A(n35541), .B(n35470), .Z(n35473) );
  XNOR U35349 ( .A(n28322), .B(p_input[666]), .Z(n35470) );
  XNOR U35350 ( .A(p_input[2075]), .B(p_input[667]), .Z(n35541) );
  XOR U35351 ( .A(p_input[2076]), .B(p_input[668]), .Z(n35474) );
  XNOR U35352 ( .A(n35484), .B(n35475), .Z(n35540) );
  XNOR U35353 ( .A(n28689), .B(p_input[657]), .Z(n35475) );
  XOR U35354 ( .A(n35542), .B(n35490), .Z(n35484) );
  XNOR U35355 ( .A(p_input[2079]), .B(p_input[671]), .Z(n35490) );
  XOR U35356 ( .A(n35481), .B(n35489), .Z(n35542) );
  XOR U35357 ( .A(n35543), .B(n35486), .Z(n35489) );
  XOR U35358 ( .A(p_input[2077]), .B(p_input[669]), .Z(n35486) );
  XNOR U35359 ( .A(p_input[2078]), .B(p_input[670]), .Z(n35543) );
  XNOR U35360 ( .A(n28326), .B(p_input[665]), .Z(n35481) );
  XNOR U35361 ( .A(n35502), .B(n35501), .Z(n35468) );
  XNOR U35362 ( .A(n35544), .B(n35508), .Z(n35501) );
  XNOR U35363 ( .A(n35497), .B(n35496), .Z(n35508) );
  XOR U35364 ( .A(n35545), .B(n35493), .Z(n35496) );
  XNOR U35365 ( .A(n28694), .B(p_input[651]), .Z(n35493) );
  XNOR U35366 ( .A(p_input[2060]), .B(p_input[652]), .Z(n35545) );
  XOR U35367 ( .A(p_input[2061]), .B(p_input[653]), .Z(n35497) );
  XNOR U35368 ( .A(n35507), .B(n35498), .Z(n35544) );
  XNOR U35369 ( .A(n28330), .B(p_input[642]), .Z(n35498) );
  XOR U35370 ( .A(n35546), .B(n35513), .Z(n35507) );
  XNOR U35371 ( .A(p_input[2064]), .B(p_input[656]), .Z(n35513) );
  XOR U35372 ( .A(n35504), .B(n35512), .Z(n35546) );
  XOR U35373 ( .A(n35547), .B(n35509), .Z(n35512) );
  XOR U35374 ( .A(p_input[2062]), .B(p_input[654]), .Z(n35509) );
  XNOR U35375 ( .A(p_input[2063]), .B(p_input[655]), .Z(n35547) );
  XNOR U35376 ( .A(n28697), .B(p_input[650]), .Z(n35504) );
  XNOR U35377 ( .A(n35519), .B(n35518), .Z(n35502) );
  XNOR U35378 ( .A(n35548), .B(n35524), .Z(n35518) );
  XOR U35379 ( .A(p_input[2057]), .B(p_input[649]), .Z(n35524) );
  XOR U35380 ( .A(n35515), .B(n35523), .Z(n35548) );
  XOR U35381 ( .A(n35549), .B(n35520), .Z(n35523) );
  XOR U35382 ( .A(p_input[2055]), .B(p_input[647]), .Z(n35520) );
  XNOR U35383 ( .A(p_input[2056]), .B(p_input[648]), .Z(n35549) );
  XNOR U35384 ( .A(n28337), .B(p_input[643]), .Z(n35515) );
  XNOR U35385 ( .A(n35529), .B(n35528), .Z(n35519) );
  XOR U35386 ( .A(n35550), .B(n35525), .Z(n35528) );
  XOR U35387 ( .A(p_input[2052]), .B(p_input[644]), .Z(n35525) );
  XNOR U35388 ( .A(p_input[2053]), .B(p_input[645]), .Z(n35550) );
  XOR U35389 ( .A(p_input[2054]), .B(p_input[646]), .Z(n35529) );
  XNOR U35390 ( .A(n35551), .B(n35552), .Z(n35334) );
  AND U35391 ( .A(n515), .B(n35553), .Z(n35552) );
  XNOR U35392 ( .A(n35554), .B(n35555), .Z(n515) );
  AND U35393 ( .A(n35556), .B(n35557), .Z(n35555) );
  XOR U35394 ( .A(n35348), .B(n35554), .Z(n35557) );
  XNOR U35395 ( .A(n35558), .B(n35554), .Z(n35556) );
  XOR U35396 ( .A(n35559), .B(n35560), .Z(n35554) );
  AND U35397 ( .A(n35561), .B(n35562), .Z(n35560) );
  XOR U35398 ( .A(n35363), .B(n35559), .Z(n35562) );
  XOR U35399 ( .A(n35559), .B(n35364), .Z(n35561) );
  XOR U35400 ( .A(n35563), .B(n35564), .Z(n35559) );
  AND U35401 ( .A(n35565), .B(n35566), .Z(n35564) );
  XOR U35402 ( .A(n35391), .B(n35563), .Z(n35566) );
  XOR U35403 ( .A(n35563), .B(n35392), .Z(n35565) );
  XOR U35404 ( .A(n35567), .B(n35568), .Z(n35563) );
  AND U35405 ( .A(n35569), .B(n35570), .Z(n35568) );
  XOR U35406 ( .A(n35440), .B(n35567), .Z(n35570) );
  XOR U35407 ( .A(n35567), .B(n35441), .Z(n35569) );
  XOR U35408 ( .A(n35571), .B(n35572), .Z(n35567) );
  AND U35409 ( .A(n35573), .B(n35574), .Z(n35572) );
  XOR U35410 ( .A(n35571), .B(n35533), .Z(n35574) );
  XNOR U35411 ( .A(n35575), .B(n35576), .Z(n35284) );
  AND U35412 ( .A(n519), .B(n35577), .Z(n35576) );
  XNOR U35413 ( .A(n35578), .B(n35579), .Z(n519) );
  AND U35414 ( .A(n35580), .B(n35581), .Z(n35579) );
  XOR U35415 ( .A(n35578), .B(n35294), .Z(n35581) );
  XNOR U35416 ( .A(n35578), .B(n35244), .Z(n35580) );
  XOR U35417 ( .A(n35582), .B(n35583), .Z(n35578) );
  AND U35418 ( .A(n35584), .B(n35585), .Z(n35583) );
  XNOR U35419 ( .A(n35304), .B(n35582), .Z(n35585) );
  XOR U35420 ( .A(n35582), .B(n35254), .Z(n35584) );
  XOR U35421 ( .A(n35586), .B(n35587), .Z(n35582) );
  AND U35422 ( .A(n35588), .B(n35589), .Z(n35587) );
  XNOR U35423 ( .A(n35314), .B(n35586), .Z(n35589) );
  XOR U35424 ( .A(n35586), .B(n35263), .Z(n35588) );
  XOR U35425 ( .A(n35590), .B(n35591), .Z(n35586) );
  AND U35426 ( .A(n35592), .B(n35593), .Z(n35591) );
  XOR U35427 ( .A(n35590), .B(n35271), .Z(n35592) );
  XOR U35428 ( .A(n35594), .B(n35595), .Z(n35235) );
  AND U35429 ( .A(n523), .B(n35577), .Z(n35595) );
  XNOR U35430 ( .A(n35575), .B(n35594), .Z(n35577) );
  XNOR U35431 ( .A(n35596), .B(n35597), .Z(n523) );
  AND U35432 ( .A(n35598), .B(n35599), .Z(n35597) );
  XNOR U35433 ( .A(n35600), .B(n35596), .Z(n35599) );
  IV U35434 ( .A(n35294), .Z(n35600) );
  XOR U35435 ( .A(n35558), .B(n35601), .Z(n35294) );
  AND U35436 ( .A(n526), .B(n35602), .Z(n35601) );
  XOR U35437 ( .A(n35347), .B(n35344), .Z(n35602) );
  IV U35438 ( .A(n35558), .Z(n35347) );
  XNOR U35439 ( .A(n35244), .B(n35596), .Z(n35598) );
  XOR U35440 ( .A(n35603), .B(n35604), .Z(n35244) );
  AND U35441 ( .A(n542), .B(n35605), .Z(n35604) );
  XOR U35442 ( .A(n35606), .B(n35607), .Z(n35596) );
  AND U35443 ( .A(n35608), .B(n35609), .Z(n35607) );
  XNOR U35444 ( .A(n35606), .B(n35304), .Z(n35609) );
  XOR U35445 ( .A(n35364), .B(n35610), .Z(n35304) );
  AND U35446 ( .A(n526), .B(n35611), .Z(n35610) );
  XOR U35447 ( .A(n35360), .B(n35364), .Z(n35611) );
  XNOR U35448 ( .A(n35612), .B(n35606), .Z(n35608) );
  IV U35449 ( .A(n35254), .Z(n35612) );
  XOR U35450 ( .A(n35613), .B(n35614), .Z(n35254) );
  AND U35451 ( .A(n542), .B(n35615), .Z(n35614) );
  XOR U35452 ( .A(n35616), .B(n35617), .Z(n35606) );
  AND U35453 ( .A(n35618), .B(n35619), .Z(n35617) );
  XNOR U35454 ( .A(n35616), .B(n35314), .Z(n35619) );
  XOR U35455 ( .A(n35392), .B(n35620), .Z(n35314) );
  AND U35456 ( .A(n526), .B(n35621), .Z(n35620) );
  XOR U35457 ( .A(n35388), .B(n35392), .Z(n35621) );
  XOR U35458 ( .A(n35263), .B(n35616), .Z(n35618) );
  XOR U35459 ( .A(n35622), .B(n35623), .Z(n35263) );
  AND U35460 ( .A(n542), .B(n35624), .Z(n35623) );
  XOR U35461 ( .A(n35590), .B(n35625), .Z(n35616) );
  AND U35462 ( .A(n35626), .B(n35593), .Z(n35625) );
  XNOR U35463 ( .A(n35324), .B(n35590), .Z(n35593) );
  XOR U35464 ( .A(n35441), .B(n35627), .Z(n35324) );
  AND U35465 ( .A(n526), .B(n35628), .Z(n35627) );
  XOR U35466 ( .A(n35437), .B(n35441), .Z(n35628) );
  XNOR U35467 ( .A(n35629), .B(n35590), .Z(n35626) );
  IV U35468 ( .A(n35271), .Z(n35629) );
  XOR U35469 ( .A(n35630), .B(n35631), .Z(n35271) );
  AND U35470 ( .A(n542), .B(n35632), .Z(n35631) );
  XOR U35471 ( .A(n35633), .B(n35634), .Z(n35590) );
  AND U35472 ( .A(n35635), .B(n35636), .Z(n35634) );
  XNOR U35473 ( .A(n35633), .B(n35332), .Z(n35636) );
  XOR U35474 ( .A(n35534), .B(n35637), .Z(n35332) );
  AND U35475 ( .A(n526), .B(n35638), .Z(n35637) );
  XOR U35476 ( .A(n35530), .B(n35534), .Z(n35638) );
  XNOR U35477 ( .A(n35639), .B(n35633), .Z(n35635) );
  IV U35478 ( .A(n35281), .Z(n35639) );
  XOR U35479 ( .A(n35640), .B(n35641), .Z(n35281) );
  AND U35480 ( .A(n542), .B(n35642), .Z(n35641) );
  AND U35481 ( .A(n35594), .B(n35575), .Z(n35633) );
  XNOR U35482 ( .A(n35643), .B(n35644), .Z(n35575) );
  AND U35483 ( .A(n526), .B(n35553), .Z(n35644) );
  XNOR U35484 ( .A(n35551), .B(n35643), .Z(n35553) );
  XNOR U35485 ( .A(n35645), .B(n35646), .Z(n526) );
  AND U35486 ( .A(n35647), .B(n35648), .Z(n35646) );
  XNOR U35487 ( .A(n35645), .B(n35344), .Z(n35648) );
  IV U35488 ( .A(n35348), .Z(n35344) );
  XOR U35489 ( .A(n35649), .B(n35650), .Z(n35348) );
  AND U35490 ( .A(n530), .B(n35651), .Z(n35650) );
  XOR U35491 ( .A(n35652), .B(n35649), .Z(n35651) );
  XNOR U35492 ( .A(n35645), .B(n35558), .Z(n35647) );
  XOR U35493 ( .A(n35653), .B(n35654), .Z(n35558) );
  AND U35494 ( .A(n538), .B(n35605), .Z(n35654) );
  XOR U35495 ( .A(n35603), .B(n35653), .Z(n35605) );
  XOR U35496 ( .A(n35655), .B(n35656), .Z(n35645) );
  AND U35497 ( .A(n35657), .B(n35658), .Z(n35656) );
  XNOR U35498 ( .A(n35655), .B(n35360), .Z(n35658) );
  IV U35499 ( .A(n35363), .Z(n35360) );
  XOR U35500 ( .A(n35659), .B(n35660), .Z(n35363) );
  AND U35501 ( .A(n530), .B(n35661), .Z(n35660) );
  XOR U35502 ( .A(n35662), .B(n35659), .Z(n35661) );
  XOR U35503 ( .A(n35364), .B(n35655), .Z(n35657) );
  XOR U35504 ( .A(n35663), .B(n35664), .Z(n35364) );
  AND U35505 ( .A(n538), .B(n35615), .Z(n35664) );
  XOR U35506 ( .A(n35663), .B(n35613), .Z(n35615) );
  XOR U35507 ( .A(n35665), .B(n35666), .Z(n35655) );
  AND U35508 ( .A(n35667), .B(n35668), .Z(n35666) );
  XNOR U35509 ( .A(n35665), .B(n35388), .Z(n35668) );
  IV U35510 ( .A(n35391), .Z(n35388) );
  XOR U35511 ( .A(n35669), .B(n35670), .Z(n35391) );
  AND U35512 ( .A(n530), .B(n35671), .Z(n35670) );
  XNOR U35513 ( .A(n35672), .B(n35669), .Z(n35671) );
  XOR U35514 ( .A(n35392), .B(n35665), .Z(n35667) );
  XOR U35515 ( .A(n35673), .B(n35674), .Z(n35392) );
  AND U35516 ( .A(n538), .B(n35624), .Z(n35674) );
  XOR U35517 ( .A(n35673), .B(n35622), .Z(n35624) );
  XOR U35518 ( .A(n35675), .B(n35676), .Z(n35665) );
  AND U35519 ( .A(n35677), .B(n35678), .Z(n35676) );
  XNOR U35520 ( .A(n35675), .B(n35437), .Z(n35678) );
  IV U35521 ( .A(n35440), .Z(n35437) );
  XOR U35522 ( .A(n35679), .B(n35680), .Z(n35440) );
  AND U35523 ( .A(n530), .B(n35681), .Z(n35680) );
  XOR U35524 ( .A(n35682), .B(n35679), .Z(n35681) );
  XOR U35525 ( .A(n35441), .B(n35675), .Z(n35677) );
  XOR U35526 ( .A(n35683), .B(n35684), .Z(n35441) );
  AND U35527 ( .A(n538), .B(n35632), .Z(n35684) );
  XOR U35528 ( .A(n35683), .B(n35630), .Z(n35632) );
  XOR U35529 ( .A(n35571), .B(n35685), .Z(n35675) );
  AND U35530 ( .A(n35573), .B(n35686), .Z(n35685) );
  XNOR U35531 ( .A(n35571), .B(n35530), .Z(n35686) );
  IV U35532 ( .A(n35533), .Z(n35530) );
  XOR U35533 ( .A(n35687), .B(n35688), .Z(n35533) );
  AND U35534 ( .A(n530), .B(n35689), .Z(n35688) );
  XNOR U35535 ( .A(n35690), .B(n35687), .Z(n35689) );
  XOR U35536 ( .A(n35534), .B(n35571), .Z(n35573) );
  XOR U35537 ( .A(n35691), .B(n35692), .Z(n35534) );
  AND U35538 ( .A(n538), .B(n35642), .Z(n35692) );
  XOR U35539 ( .A(n35691), .B(n35640), .Z(n35642) );
  AND U35540 ( .A(n35643), .B(n35551), .Z(n35571) );
  XNOR U35541 ( .A(n35693), .B(n35694), .Z(n35551) );
  AND U35542 ( .A(n530), .B(n35695), .Z(n35694) );
  XNOR U35543 ( .A(n35696), .B(n35693), .Z(n35695) );
  XNOR U35544 ( .A(n35697), .B(n35698), .Z(n530) );
  AND U35545 ( .A(n35699), .B(n35700), .Z(n35698) );
  XOR U35546 ( .A(n35652), .B(n35697), .Z(n35700) );
  AND U35547 ( .A(n35701), .B(n35702), .Z(n35652) );
  XNOR U35548 ( .A(n35649), .B(n35697), .Z(n35699) );
  XNOR U35549 ( .A(n35703), .B(n35704), .Z(n35649) );
  AND U35550 ( .A(n534), .B(n35705), .Z(n35704) );
  XNOR U35551 ( .A(n35706), .B(n35707), .Z(n35705) );
  XOR U35552 ( .A(n35708), .B(n35709), .Z(n35697) );
  AND U35553 ( .A(n35710), .B(n35711), .Z(n35709) );
  XNOR U35554 ( .A(n35708), .B(n35701), .Z(n35711) );
  IV U35555 ( .A(n35662), .Z(n35701) );
  XOR U35556 ( .A(n35712), .B(n35713), .Z(n35662) );
  XOR U35557 ( .A(n35714), .B(n35702), .Z(n35713) );
  AND U35558 ( .A(n35672), .B(n35715), .Z(n35702) );
  AND U35559 ( .A(n35716), .B(n35717), .Z(n35714) );
  XOR U35560 ( .A(n35718), .B(n35712), .Z(n35716) );
  XNOR U35561 ( .A(n35659), .B(n35708), .Z(n35710) );
  XNOR U35562 ( .A(n35719), .B(n35720), .Z(n35659) );
  AND U35563 ( .A(n534), .B(n35721), .Z(n35720) );
  XNOR U35564 ( .A(n35722), .B(n35723), .Z(n35721) );
  XOR U35565 ( .A(n35724), .B(n35725), .Z(n35708) );
  AND U35566 ( .A(n35726), .B(n35727), .Z(n35725) );
  XNOR U35567 ( .A(n35724), .B(n35672), .Z(n35727) );
  XOR U35568 ( .A(n35728), .B(n35717), .Z(n35672) );
  XNOR U35569 ( .A(n35729), .B(n35712), .Z(n35717) );
  XOR U35570 ( .A(n35730), .B(n35731), .Z(n35712) );
  AND U35571 ( .A(n35732), .B(n35733), .Z(n35731) );
  XOR U35572 ( .A(n35734), .B(n35730), .Z(n35732) );
  XNOR U35573 ( .A(n35735), .B(n35736), .Z(n35729) );
  AND U35574 ( .A(n35737), .B(n35738), .Z(n35736) );
  XOR U35575 ( .A(n35735), .B(n35739), .Z(n35737) );
  XNOR U35576 ( .A(n35718), .B(n35715), .Z(n35728) );
  AND U35577 ( .A(n35740), .B(n35741), .Z(n35715) );
  XOR U35578 ( .A(n35742), .B(n35743), .Z(n35718) );
  AND U35579 ( .A(n35744), .B(n35745), .Z(n35743) );
  XOR U35580 ( .A(n35742), .B(n35746), .Z(n35744) );
  XNOR U35581 ( .A(n35669), .B(n35724), .Z(n35726) );
  XNOR U35582 ( .A(n35747), .B(n35748), .Z(n35669) );
  AND U35583 ( .A(n534), .B(n35749), .Z(n35748) );
  XNOR U35584 ( .A(n35750), .B(n35751), .Z(n35749) );
  XOR U35585 ( .A(n35752), .B(n35753), .Z(n35724) );
  AND U35586 ( .A(n35754), .B(n35755), .Z(n35753) );
  XNOR U35587 ( .A(n35752), .B(n35740), .Z(n35755) );
  IV U35588 ( .A(n35682), .Z(n35740) );
  XNOR U35589 ( .A(n35756), .B(n35733), .Z(n35682) );
  XNOR U35590 ( .A(n35757), .B(n35739), .Z(n35733) );
  XOR U35591 ( .A(n35758), .B(n35759), .Z(n35739) );
  AND U35592 ( .A(n35760), .B(n35761), .Z(n35759) );
  XOR U35593 ( .A(n35758), .B(n35762), .Z(n35760) );
  XNOR U35594 ( .A(n35738), .B(n35730), .Z(n35757) );
  XOR U35595 ( .A(n35763), .B(n35764), .Z(n35730) );
  AND U35596 ( .A(n35765), .B(n35766), .Z(n35764) );
  XNOR U35597 ( .A(n35767), .B(n35763), .Z(n35765) );
  XNOR U35598 ( .A(n35768), .B(n35735), .Z(n35738) );
  XOR U35599 ( .A(n35769), .B(n35770), .Z(n35735) );
  AND U35600 ( .A(n35771), .B(n35772), .Z(n35770) );
  XOR U35601 ( .A(n35769), .B(n35773), .Z(n35771) );
  XNOR U35602 ( .A(n35774), .B(n35775), .Z(n35768) );
  AND U35603 ( .A(n35776), .B(n35777), .Z(n35775) );
  XNOR U35604 ( .A(n35774), .B(n35778), .Z(n35776) );
  XNOR U35605 ( .A(n35734), .B(n35741), .Z(n35756) );
  AND U35606 ( .A(n35690), .B(n35779), .Z(n35741) );
  XOR U35607 ( .A(n35746), .B(n35745), .Z(n35734) );
  XNOR U35608 ( .A(n35780), .B(n35742), .Z(n35745) );
  XOR U35609 ( .A(n35781), .B(n35782), .Z(n35742) );
  AND U35610 ( .A(n35783), .B(n35784), .Z(n35782) );
  XOR U35611 ( .A(n35781), .B(n35785), .Z(n35783) );
  XNOR U35612 ( .A(n35786), .B(n35787), .Z(n35780) );
  AND U35613 ( .A(n35788), .B(n35789), .Z(n35787) );
  XOR U35614 ( .A(n35786), .B(n35790), .Z(n35788) );
  XOR U35615 ( .A(n35791), .B(n35792), .Z(n35746) );
  AND U35616 ( .A(n35793), .B(n35794), .Z(n35792) );
  XOR U35617 ( .A(n35791), .B(n35795), .Z(n35793) );
  XNOR U35618 ( .A(n35679), .B(n35752), .Z(n35754) );
  XNOR U35619 ( .A(n35796), .B(n35797), .Z(n35679) );
  AND U35620 ( .A(n534), .B(n35798), .Z(n35797) );
  XNOR U35621 ( .A(n35799), .B(n35800), .Z(n35798) );
  XOR U35622 ( .A(n35801), .B(n35802), .Z(n35752) );
  AND U35623 ( .A(n35803), .B(n35804), .Z(n35802) );
  XNOR U35624 ( .A(n35801), .B(n35690), .Z(n35804) );
  XOR U35625 ( .A(n35805), .B(n35766), .Z(n35690) );
  XNOR U35626 ( .A(n35806), .B(n35773), .Z(n35766) );
  XOR U35627 ( .A(n35762), .B(n35761), .Z(n35773) );
  XNOR U35628 ( .A(n35807), .B(n35758), .Z(n35761) );
  XOR U35629 ( .A(n35808), .B(n35809), .Z(n35758) );
  AND U35630 ( .A(n35810), .B(n35811), .Z(n35809) );
  XOR U35631 ( .A(n35808), .B(n35812), .Z(n35810) );
  XNOR U35632 ( .A(n35813), .B(n35814), .Z(n35807) );
  NOR U35633 ( .A(n35815), .B(n35816), .Z(n35814) );
  XNOR U35634 ( .A(n35813), .B(n35817), .Z(n35815) );
  XOR U35635 ( .A(n35818), .B(n35819), .Z(n35762) );
  NOR U35636 ( .A(n35820), .B(n35821), .Z(n35819) );
  XNOR U35637 ( .A(n35818), .B(n35822), .Z(n35820) );
  XNOR U35638 ( .A(n35772), .B(n35763), .Z(n35806) );
  XOR U35639 ( .A(n35823), .B(n35824), .Z(n35763) );
  NOR U35640 ( .A(n35825), .B(n35826), .Z(n35824) );
  XNOR U35641 ( .A(n35823), .B(n35827), .Z(n35825) );
  XOR U35642 ( .A(n35828), .B(n35778), .Z(n35772) );
  XNOR U35643 ( .A(n35829), .B(n35830), .Z(n35778) );
  NOR U35644 ( .A(n35831), .B(n35832), .Z(n35830) );
  XNOR U35645 ( .A(n35829), .B(n35833), .Z(n35831) );
  XNOR U35646 ( .A(n35777), .B(n35769), .Z(n35828) );
  XOR U35647 ( .A(n35834), .B(n35835), .Z(n35769) );
  AND U35648 ( .A(n35836), .B(n35837), .Z(n35835) );
  XOR U35649 ( .A(n35834), .B(n35838), .Z(n35836) );
  XNOR U35650 ( .A(n35839), .B(n35774), .Z(n35777) );
  XOR U35651 ( .A(n35840), .B(n35841), .Z(n35774) );
  AND U35652 ( .A(n35842), .B(n35843), .Z(n35841) );
  XOR U35653 ( .A(n35840), .B(n35844), .Z(n35842) );
  XNOR U35654 ( .A(n35845), .B(n35846), .Z(n35839) );
  NOR U35655 ( .A(n35847), .B(n35848), .Z(n35846) );
  XOR U35656 ( .A(n35845), .B(n35849), .Z(n35847) );
  XOR U35657 ( .A(n35767), .B(n35779), .Z(n35805) );
  NOR U35658 ( .A(n35696), .B(n35850), .Z(n35779) );
  XNOR U35659 ( .A(n35785), .B(n35784), .Z(n35767) );
  XNOR U35660 ( .A(n35851), .B(n35790), .Z(n35784) );
  XOR U35661 ( .A(n35852), .B(n35853), .Z(n35790) );
  NOR U35662 ( .A(n35854), .B(n35855), .Z(n35853) );
  XNOR U35663 ( .A(n35852), .B(n35856), .Z(n35854) );
  XNOR U35664 ( .A(n35789), .B(n35781), .Z(n35851) );
  XOR U35665 ( .A(n35857), .B(n35858), .Z(n35781) );
  AND U35666 ( .A(n35859), .B(n35860), .Z(n35858) );
  XNOR U35667 ( .A(n35857), .B(n35861), .Z(n35859) );
  XNOR U35668 ( .A(n35862), .B(n35786), .Z(n35789) );
  XOR U35669 ( .A(n35863), .B(n35864), .Z(n35786) );
  AND U35670 ( .A(n35865), .B(n35866), .Z(n35864) );
  XOR U35671 ( .A(n35863), .B(n35867), .Z(n35865) );
  XNOR U35672 ( .A(n35868), .B(n35869), .Z(n35862) );
  NOR U35673 ( .A(n35870), .B(n35871), .Z(n35869) );
  XOR U35674 ( .A(n35868), .B(n35872), .Z(n35870) );
  XOR U35675 ( .A(n35795), .B(n35794), .Z(n35785) );
  XNOR U35676 ( .A(n35873), .B(n35791), .Z(n35794) );
  XOR U35677 ( .A(n35874), .B(n35875), .Z(n35791) );
  AND U35678 ( .A(n35876), .B(n35877), .Z(n35875) );
  XOR U35679 ( .A(n35874), .B(n35878), .Z(n35876) );
  XNOR U35680 ( .A(n35879), .B(n35880), .Z(n35873) );
  NOR U35681 ( .A(n35881), .B(n35882), .Z(n35880) );
  XNOR U35682 ( .A(n35879), .B(n35883), .Z(n35881) );
  XOR U35683 ( .A(n35884), .B(n35885), .Z(n35795) );
  NOR U35684 ( .A(n35886), .B(n35887), .Z(n35885) );
  XNOR U35685 ( .A(n35884), .B(n35888), .Z(n35886) );
  XNOR U35686 ( .A(n35687), .B(n35801), .Z(n35803) );
  XNOR U35687 ( .A(n35889), .B(n35890), .Z(n35687) );
  AND U35688 ( .A(n534), .B(n35891), .Z(n35890) );
  XNOR U35689 ( .A(n35892), .B(n35893), .Z(n35891) );
  AND U35690 ( .A(n35693), .B(n35696), .Z(n35801) );
  XOR U35691 ( .A(n35894), .B(n35850), .Z(n35696) );
  XNOR U35692 ( .A(p_input[2048]), .B(p_input[672]), .Z(n35850) );
  XOR U35693 ( .A(n35827), .B(n35826), .Z(n35894) );
  XOR U35694 ( .A(n35895), .B(n35838), .Z(n35826) );
  XOR U35695 ( .A(n35812), .B(n35811), .Z(n35838) );
  XNOR U35696 ( .A(n35896), .B(n35817), .Z(n35811) );
  XOR U35697 ( .A(p_input[2072]), .B(p_input[696]), .Z(n35817) );
  XOR U35698 ( .A(n35808), .B(n35816), .Z(n35896) );
  XOR U35699 ( .A(n35897), .B(n35813), .Z(n35816) );
  XOR U35700 ( .A(p_input[2070]), .B(p_input[694]), .Z(n35813) );
  XNOR U35701 ( .A(p_input[2071]), .B(p_input[695]), .Z(n35897) );
  XNOR U35702 ( .A(n28684), .B(p_input[690]), .Z(n35808) );
  XNOR U35703 ( .A(n35822), .B(n35821), .Z(n35812) );
  XOR U35704 ( .A(n35898), .B(n35818), .Z(n35821) );
  XOR U35705 ( .A(p_input[2067]), .B(p_input[691]), .Z(n35818) );
  XNOR U35706 ( .A(p_input[2068]), .B(p_input[692]), .Z(n35898) );
  XOR U35707 ( .A(p_input[2069]), .B(p_input[693]), .Z(n35822) );
  XNOR U35708 ( .A(n35837), .B(n35823), .Z(n35895) );
  XNOR U35709 ( .A(n28686), .B(p_input[673]), .Z(n35823) );
  XNOR U35710 ( .A(n35899), .B(n35844), .Z(n35837) );
  XNOR U35711 ( .A(n35833), .B(n35832), .Z(n35844) );
  XOR U35712 ( .A(n35900), .B(n35829), .Z(n35832) );
  XNOR U35713 ( .A(n28322), .B(p_input[698]), .Z(n35829) );
  XNOR U35714 ( .A(p_input[2075]), .B(p_input[699]), .Z(n35900) );
  XOR U35715 ( .A(p_input[2076]), .B(p_input[700]), .Z(n35833) );
  XNOR U35716 ( .A(n35843), .B(n35834), .Z(n35899) );
  XNOR U35717 ( .A(n28689), .B(p_input[689]), .Z(n35834) );
  XOR U35718 ( .A(n35901), .B(n35849), .Z(n35843) );
  XNOR U35719 ( .A(p_input[2079]), .B(p_input[703]), .Z(n35849) );
  XOR U35720 ( .A(n35840), .B(n35848), .Z(n35901) );
  XOR U35721 ( .A(n35902), .B(n35845), .Z(n35848) );
  XOR U35722 ( .A(p_input[2077]), .B(p_input[701]), .Z(n35845) );
  XNOR U35723 ( .A(p_input[2078]), .B(p_input[702]), .Z(n35902) );
  XNOR U35724 ( .A(n28326), .B(p_input[697]), .Z(n35840) );
  XNOR U35725 ( .A(n35861), .B(n35860), .Z(n35827) );
  XNOR U35726 ( .A(n35903), .B(n35867), .Z(n35860) );
  XNOR U35727 ( .A(n35856), .B(n35855), .Z(n35867) );
  XOR U35728 ( .A(n35904), .B(n35852), .Z(n35855) );
  XNOR U35729 ( .A(n28694), .B(p_input[683]), .Z(n35852) );
  XNOR U35730 ( .A(p_input[2060]), .B(p_input[684]), .Z(n35904) );
  XOR U35731 ( .A(p_input[2061]), .B(p_input[685]), .Z(n35856) );
  XNOR U35732 ( .A(n35866), .B(n35857), .Z(n35903) );
  XNOR U35733 ( .A(n28330), .B(p_input[674]), .Z(n35857) );
  XOR U35734 ( .A(n35905), .B(n35872), .Z(n35866) );
  XNOR U35735 ( .A(p_input[2064]), .B(p_input[688]), .Z(n35872) );
  XOR U35736 ( .A(n35863), .B(n35871), .Z(n35905) );
  XOR U35737 ( .A(n35906), .B(n35868), .Z(n35871) );
  XOR U35738 ( .A(p_input[2062]), .B(p_input[686]), .Z(n35868) );
  XNOR U35739 ( .A(p_input[2063]), .B(p_input[687]), .Z(n35906) );
  XNOR U35740 ( .A(n28697), .B(p_input[682]), .Z(n35863) );
  XNOR U35741 ( .A(n35878), .B(n35877), .Z(n35861) );
  XNOR U35742 ( .A(n35907), .B(n35883), .Z(n35877) );
  XOR U35743 ( .A(p_input[2057]), .B(p_input[681]), .Z(n35883) );
  XOR U35744 ( .A(n35874), .B(n35882), .Z(n35907) );
  XOR U35745 ( .A(n35908), .B(n35879), .Z(n35882) );
  XOR U35746 ( .A(p_input[2055]), .B(p_input[679]), .Z(n35879) );
  XNOR U35747 ( .A(p_input[2056]), .B(p_input[680]), .Z(n35908) );
  XNOR U35748 ( .A(n28337), .B(p_input[675]), .Z(n35874) );
  XNOR U35749 ( .A(n35888), .B(n35887), .Z(n35878) );
  XOR U35750 ( .A(n35909), .B(n35884), .Z(n35887) );
  XOR U35751 ( .A(p_input[2052]), .B(p_input[676]), .Z(n35884) );
  XNOR U35752 ( .A(p_input[2053]), .B(p_input[677]), .Z(n35909) );
  XOR U35753 ( .A(p_input[2054]), .B(p_input[678]), .Z(n35888) );
  XNOR U35754 ( .A(n35910), .B(n35911), .Z(n35693) );
  AND U35755 ( .A(n534), .B(n35912), .Z(n35911) );
  XNOR U35756 ( .A(n35913), .B(n35914), .Z(n534) );
  AND U35757 ( .A(n35915), .B(n35916), .Z(n35914) );
  XOR U35758 ( .A(n35707), .B(n35913), .Z(n35916) );
  XNOR U35759 ( .A(n35917), .B(n35913), .Z(n35915) );
  XOR U35760 ( .A(n35918), .B(n35919), .Z(n35913) );
  AND U35761 ( .A(n35920), .B(n35921), .Z(n35919) );
  XOR U35762 ( .A(n35722), .B(n35918), .Z(n35921) );
  XOR U35763 ( .A(n35918), .B(n35723), .Z(n35920) );
  XOR U35764 ( .A(n35922), .B(n35923), .Z(n35918) );
  AND U35765 ( .A(n35924), .B(n35925), .Z(n35923) );
  XOR U35766 ( .A(n35750), .B(n35922), .Z(n35925) );
  XOR U35767 ( .A(n35922), .B(n35751), .Z(n35924) );
  XOR U35768 ( .A(n35926), .B(n35927), .Z(n35922) );
  AND U35769 ( .A(n35928), .B(n35929), .Z(n35927) );
  XOR U35770 ( .A(n35799), .B(n35926), .Z(n35929) );
  XOR U35771 ( .A(n35926), .B(n35800), .Z(n35928) );
  XOR U35772 ( .A(n35930), .B(n35931), .Z(n35926) );
  AND U35773 ( .A(n35932), .B(n35933), .Z(n35931) );
  XOR U35774 ( .A(n35930), .B(n35892), .Z(n35933) );
  XNOR U35775 ( .A(n35934), .B(n35935), .Z(n35643) );
  AND U35776 ( .A(n538), .B(n35936), .Z(n35935) );
  XNOR U35777 ( .A(n35937), .B(n35938), .Z(n538) );
  AND U35778 ( .A(n35939), .B(n35940), .Z(n35938) );
  XOR U35779 ( .A(n35937), .B(n35653), .Z(n35940) );
  XNOR U35780 ( .A(n35937), .B(n35603), .Z(n35939) );
  XOR U35781 ( .A(n35941), .B(n35942), .Z(n35937) );
  AND U35782 ( .A(n35943), .B(n35944), .Z(n35942) );
  XNOR U35783 ( .A(n35663), .B(n35941), .Z(n35944) );
  XOR U35784 ( .A(n35941), .B(n35613), .Z(n35943) );
  XOR U35785 ( .A(n35945), .B(n35946), .Z(n35941) );
  AND U35786 ( .A(n35947), .B(n35948), .Z(n35946) );
  XNOR U35787 ( .A(n35673), .B(n35945), .Z(n35948) );
  XOR U35788 ( .A(n35945), .B(n35622), .Z(n35947) );
  XOR U35789 ( .A(n35949), .B(n35950), .Z(n35945) );
  AND U35790 ( .A(n35951), .B(n35952), .Z(n35950) );
  XOR U35791 ( .A(n35949), .B(n35630), .Z(n35951) );
  XOR U35792 ( .A(n35953), .B(n35954), .Z(n35594) );
  AND U35793 ( .A(n542), .B(n35936), .Z(n35954) );
  XNOR U35794 ( .A(n35934), .B(n35953), .Z(n35936) );
  XNOR U35795 ( .A(n35955), .B(n35956), .Z(n542) );
  AND U35796 ( .A(n35957), .B(n35958), .Z(n35956) );
  XNOR U35797 ( .A(n35959), .B(n35955), .Z(n35958) );
  IV U35798 ( .A(n35653), .Z(n35959) );
  XOR U35799 ( .A(n35917), .B(n35960), .Z(n35653) );
  AND U35800 ( .A(n545), .B(n35961), .Z(n35960) );
  XOR U35801 ( .A(n35706), .B(n35703), .Z(n35961) );
  IV U35802 ( .A(n35917), .Z(n35706) );
  XNOR U35803 ( .A(n35603), .B(n35955), .Z(n35957) );
  XOR U35804 ( .A(n35962), .B(n35963), .Z(n35603) );
  AND U35805 ( .A(n561), .B(n35964), .Z(n35963) );
  XOR U35806 ( .A(n35965), .B(n35966), .Z(n35955) );
  AND U35807 ( .A(n35967), .B(n35968), .Z(n35966) );
  XNOR U35808 ( .A(n35965), .B(n35663), .Z(n35968) );
  XOR U35809 ( .A(n35723), .B(n35969), .Z(n35663) );
  AND U35810 ( .A(n545), .B(n35970), .Z(n35969) );
  XOR U35811 ( .A(n35719), .B(n35723), .Z(n35970) );
  XNOR U35812 ( .A(n35971), .B(n35965), .Z(n35967) );
  IV U35813 ( .A(n35613), .Z(n35971) );
  XOR U35814 ( .A(n35972), .B(n35973), .Z(n35613) );
  AND U35815 ( .A(n561), .B(n35974), .Z(n35973) );
  XOR U35816 ( .A(n35975), .B(n35976), .Z(n35965) );
  AND U35817 ( .A(n35977), .B(n35978), .Z(n35976) );
  XNOR U35818 ( .A(n35975), .B(n35673), .Z(n35978) );
  XOR U35819 ( .A(n35751), .B(n35979), .Z(n35673) );
  AND U35820 ( .A(n545), .B(n35980), .Z(n35979) );
  XOR U35821 ( .A(n35747), .B(n35751), .Z(n35980) );
  XOR U35822 ( .A(n35622), .B(n35975), .Z(n35977) );
  XOR U35823 ( .A(n35981), .B(n35982), .Z(n35622) );
  AND U35824 ( .A(n561), .B(n35983), .Z(n35982) );
  XOR U35825 ( .A(n35949), .B(n35984), .Z(n35975) );
  AND U35826 ( .A(n35985), .B(n35952), .Z(n35984) );
  XNOR U35827 ( .A(n35683), .B(n35949), .Z(n35952) );
  XOR U35828 ( .A(n35800), .B(n35986), .Z(n35683) );
  AND U35829 ( .A(n545), .B(n35987), .Z(n35986) );
  XOR U35830 ( .A(n35796), .B(n35800), .Z(n35987) );
  XNOR U35831 ( .A(n35988), .B(n35949), .Z(n35985) );
  IV U35832 ( .A(n35630), .Z(n35988) );
  XOR U35833 ( .A(n35989), .B(n35990), .Z(n35630) );
  AND U35834 ( .A(n561), .B(n35991), .Z(n35990) );
  XOR U35835 ( .A(n35992), .B(n35993), .Z(n35949) );
  AND U35836 ( .A(n35994), .B(n35995), .Z(n35993) );
  XNOR U35837 ( .A(n35992), .B(n35691), .Z(n35995) );
  XOR U35838 ( .A(n35893), .B(n35996), .Z(n35691) );
  AND U35839 ( .A(n545), .B(n35997), .Z(n35996) );
  XOR U35840 ( .A(n35889), .B(n35893), .Z(n35997) );
  XNOR U35841 ( .A(n35998), .B(n35992), .Z(n35994) );
  IV U35842 ( .A(n35640), .Z(n35998) );
  XOR U35843 ( .A(n35999), .B(n36000), .Z(n35640) );
  AND U35844 ( .A(n561), .B(n36001), .Z(n36000) );
  AND U35845 ( .A(n35953), .B(n35934), .Z(n35992) );
  XNOR U35846 ( .A(n36002), .B(n36003), .Z(n35934) );
  AND U35847 ( .A(n545), .B(n35912), .Z(n36003) );
  XNOR U35848 ( .A(n35910), .B(n36002), .Z(n35912) );
  XNOR U35849 ( .A(n36004), .B(n36005), .Z(n545) );
  AND U35850 ( .A(n36006), .B(n36007), .Z(n36005) );
  XNOR U35851 ( .A(n36004), .B(n35703), .Z(n36007) );
  IV U35852 ( .A(n35707), .Z(n35703) );
  XOR U35853 ( .A(n36008), .B(n36009), .Z(n35707) );
  AND U35854 ( .A(n549), .B(n36010), .Z(n36009) );
  XOR U35855 ( .A(n36011), .B(n36008), .Z(n36010) );
  XNOR U35856 ( .A(n36004), .B(n35917), .Z(n36006) );
  XOR U35857 ( .A(n36012), .B(n36013), .Z(n35917) );
  AND U35858 ( .A(n557), .B(n35964), .Z(n36013) );
  XOR U35859 ( .A(n35962), .B(n36012), .Z(n35964) );
  XOR U35860 ( .A(n36014), .B(n36015), .Z(n36004) );
  AND U35861 ( .A(n36016), .B(n36017), .Z(n36015) );
  XNOR U35862 ( .A(n36014), .B(n35719), .Z(n36017) );
  IV U35863 ( .A(n35722), .Z(n35719) );
  XOR U35864 ( .A(n36018), .B(n36019), .Z(n35722) );
  AND U35865 ( .A(n549), .B(n36020), .Z(n36019) );
  XOR U35866 ( .A(n36021), .B(n36018), .Z(n36020) );
  XOR U35867 ( .A(n35723), .B(n36014), .Z(n36016) );
  XOR U35868 ( .A(n36022), .B(n36023), .Z(n35723) );
  AND U35869 ( .A(n557), .B(n35974), .Z(n36023) );
  XOR U35870 ( .A(n36022), .B(n35972), .Z(n35974) );
  XOR U35871 ( .A(n36024), .B(n36025), .Z(n36014) );
  AND U35872 ( .A(n36026), .B(n36027), .Z(n36025) );
  XNOR U35873 ( .A(n36024), .B(n35747), .Z(n36027) );
  IV U35874 ( .A(n35750), .Z(n35747) );
  XOR U35875 ( .A(n36028), .B(n36029), .Z(n35750) );
  AND U35876 ( .A(n549), .B(n36030), .Z(n36029) );
  XNOR U35877 ( .A(n36031), .B(n36028), .Z(n36030) );
  XOR U35878 ( .A(n35751), .B(n36024), .Z(n36026) );
  XOR U35879 ( .A(n36032), .B(n36033), .Z(n35751) );
  AND U35880 ( .A(n557), .B(n35983), .Z(n36033) );
  XOR U35881 ( .A(n36032), .B(n35981), .Z(n35983) );
  XOR U35882 ( .A(n36034), .B(n36035), .Z(n36024) );
  AND U35883 ( .A(n36036), .B(n36037), .Z(n36035) );
  XNOR U35884 ( .A(n36034), .B(n35796), .Z(n36037) );
  IV U35885 ( .A(n35799), .Z(n35796) );
  XOR U35886 ( .A(n36038), .B(n36039), .Z(n35799) );
  AND U35887 ( .A(n549), .B(n36040), .Z(n36039) );
  XOR U35888 ( .A(n36041), .B(n36038), .Z(n36040) );
  XOR U35889 ( .A(n35800), .B(n36034), .Z(n36036) );
  XOR U35890 ( .A(n36042), .B(n36043), .Z(n35800) );
  AND U35891 ( .A(n557), .B(n35991), .Z(n36043) );
  XOR U35892 ( .A(n36042), .B(n35989), .Z(n35991) );
  XOR U35893 ( .A(n35930), .B(n36044), .Z(n36034) );
  AND U35894 ( .A(n35932), .B(n36045), .Z(n36044) );
  XNOR U35895 ( .A(n35930), .B(n35889), .Z(n36045) );
  IV U35896 ( .A(n35892), .Z(n35889) );
  XOR U35897 ( .A(n36046), .B(n36047), .Z(n35892) );
  AND U35898 ( .A(n549), .B(n36048), .Z(n36047) );
  XNOR U35899 ( .A(n36049), .B(n36046), .Z(n36048) );
  XOR U35900 ( .A(n35893), .B(n35930), .Z(n35932) );
  XOR U35901 ( .A(n36050), .B(n36051), .Z(n35893) );
  AND U35902 ( .A(n557), .B(n36001), .Z(n36051) );
  XOR U35903 ( .A(n36050), .B(n35999), .Z(n36001) );
  AND U35904 ( .A(n36002), .B(n35910), .Z(n35930) );
  XNOR U35905 ( .A(n36052), .B(n36053), .Z(n35910) );
  AND U35906 ( .A(n549), .B(n36054), .Z(n36053) );
  XNOR U35907 ( .A(n36055), .B(n36052), .Z(n36054) );
  XNOR U35908 ( .A(n36056), .B(n36057), .Z(n549) );
  AND U35909 ( .A(n36058), .B(n36059), .Z(n36057) );
  XOR U35910 ( .A(n36011), .B(n36056), .Z(n36059) );
  AND U35911 ( .A(n36060), .B(n36061), .Z(n36011) );
  XNOR U35912 ( .A(n36008), .B(n36056), .Z(n36058) );
  XNOR U35913 ( .A(n36062), .B(n36063), .Z(n36008) );
  AND U35914 ( .A(n553), .B(n36064), .Z(n36063) );
  XNOR U35915 ( .A(n36065), .B(n36066), .Z(n36064) );
  XOR U35916 ( .A(n36067), .B(n36068), .Z(n36056) );
  AND U35917 ( .A(n36069), .B(n36070), .Z(n36068) );
  XNOR U35918 ( .A(n36067), .B(n36060), .Z(n36070) );
  IV U35919 ( .A(n36021), .Z(n36060) );
  XOR U35920 ( .A(n36071), .B(n36072), .Z(n36021) );
  XOR U35921 ( .A(n36073), .B(n36061), .Z(n36072) );
  AND U35922 ( .A(n36031), .B(n36074), .Z(n36061) );
  AND U35923 ( .A(n36075), .B(n36076), .Z(n36073) );
  XOR U35924 ( .A(n36077), .B(n36071), .Z(n36075) );
  XNOR U35925 ( .A(n36018), .B(n36067), .Z(n36069) );
  XNOR U35926 ( .A(n36078), .B(n36079), .Z(n36018) );
  AND U35927 ( .A(n553), .B(n36080), .Z(n36079) );
  XNOR U35928 ( .A(n36081), .B(n36082), .Z(n36080) );
  XOR U35929 ( .A(n36083), .B(n36084), .Z(n36067) );
  AND U35930 ( .A(n36085), .B(n36086), .Z(n36084) );
  XNOR U35931 ( .A(n36083), .B(n36031), .Z(n36086) );
  XOR U35932 ( .A(n36087), .B(n36076), .Z(n36031) );
  XNOR U35933 ( .A(n36088), .B(n36071), .Z(n36076) );
  XOR U35934 ( .A(n36089), .B(n36090), .Z(n36071) );
  AND U35935 ( .A(n36091), .B(n36092), .Z(n36090) );
  XOR U35936 ( .A(n36093), .B(n36089), .Z(n36091) );
  XNOR U35937 ( .A(n36094), .B(n36095), .Z(n36088) );
  AND U35938 ( .A(n36096), .B(n36097), .Z(n36095) );
  XOR U35939 ( .A(n36094), .B(n36098), .Z(n36096) );
  XNOR U35940 ( .A(n36077), .B(n36074), .Z(n36087) );
  AND U35941 ( .A(n36099), .B(n36100), .Z(n36074) );
  XOR U35942 ( .A(n36101), .B(n36102), .Z(n36077) );
  AND U35943 ( .A(n36103), .B(n36104), .Z(n36102) );
  XOR U35944 ( .A(n36101), .B(n36105), .Z(n36103) );
  XNOR U35945 ( .A(n36028), .B(n36083), .Z(n36085) );
  XNOR U35946 ( .A(n36106), .B(n36107), .Z(n36028) );
  AND U35947 ( .A(n553), .B(n36108), .Z(n36107) );
  XNOR U35948 ( .A(n36109), .B(n36110), .Z(n36108) );
  XOR U35949 ( .A(n36111), .B(n36112), .Z(n36083) );
  AND U35950 ( .A(n36113), .B(n36114), .Z(n36112) );
  XNOR U35951 ( .A(n36111), .B(n36099), .Z(n36114) );
  IV U35952 ( .A(n36041), .Z(n36099) );
  XNOR U35953 ( .A(n36115), .B(n36092), .Z(n36041) );
  XNOR U35954 ( .A(n36116), .B(n36098), .Z(n36092) );
  XOR U35955 ( .A(n36117), .B(n36118), .Z(n36098) );
  AND U35956 ( .A(n36119), .B(n36120), .Z(n36118) );
  XOR U35957 ( .A(n36117), .B(n36121), .Z(n36119) );
  XNOR U35958 ( .A(n36097), .B(n36089), .Z(n36116) );
  XOR U35959 ( .A(n36122), .B(n36123), .Z(n36089) );
  AND U35960 ( .A(n36124), .B(n36125), .Z(n36123) );
  XNOR U35961 ( .A(n36126), .B(n36122), .Z(n36124) );
  XNOR U35962 ( .A(n36127), .B(n36094), .Z(n36097) );
  XOR U35963 ( .A(n36128), .B(n36129), .Z(n36094) );
  AND U35964 ( .A(n36130), .B(n36131), .Z(n36129) );
  XOR U35965 ( .A(n36128), .B(n36132), .Z(n36130) );
  XNOR U35966 ( .A(n36133), .B(n36134), .Z(n36127) );
  AND U35967 ( .A(n36135), .B(n36136), .Z(n36134) );
  XNOR U35968 ( .A(n36133), .B(n36137), .Z(n36135) );
  XNOR U35969 ( .A(n36093), .B(n36100), .Z(n36115) );
  AND U35970 ( .A(n36049), .B(n36138), .Z(n36100) );
  XOR U35971 ( .A(n36105), .B(n36104), .Z(n36093) );
  XNOR U35972 ( .A(n36139), .B(n36101), .Z(n36104) );
  XOR U35973 ( .A(n36140), .B(n36141), .Z(n36101) );
  AND U35974 ( .A(n36142), .B(n36143), .Z(n36141) );
  XOR U35975 ( .A(n36140), .B(n36144), .Z(n36142) );
  XNOR U35976 ( .A(n36145), .B(n36146), .Z(n36139) );
  AND U35977 ( .A(n36147), .B(n36148), .Z(n36146) );
  XOR U35978 ( .A(n36145), .B(n36149), .Z(n36147) );
  XOR U35979 ( .A(n36150), .B(n36151), .Z(n36105) );
  AND U35980 ( .A(n36152), .B(n36153), .Z(n36151) );
  XOR U35981 ( .A(n36150), .B(n36154), .Z(n36152) );
  XNOR U35982 ( .A(n36038), .B(n36111), .Z(n36113) );
  XNOR U35983 ( .A(n36155), .B(n36156), .Z(n36038) );
  AND U35984 ( .A(n553), .B(n36157), .Z(n36156) );
  XNOR U35985 ( .A(n36158), .B(n36159), .Z(n36157) );
  XOR U35986 ( .A(n36160), .B(n36161), .Z(n36111) );
  AND U35987 ( .A(n36162), .B(n36163), .Z(n36161) );
  XNOR U35988 ( .A(n36160), .B(n36049), .Z(n36163) );
  XOR U35989 ( .A(n36164), .B(n36125), .Z(n36049) );
  XNOR U35990 ( .A(n36165), .B(n36132), .Z(n36125) );
  XOR U35991 ( .A(n36121), .B(n36120), .Z(n36132) );
  XNOR U35992 ( .A(n36166), .B(n36117), .Z(n36120) );
  XOR U35993 ( .A(n36167), .B(n36168), .Z(n36117) );
  AND U35994 ( .A(n36169), .B(n36170), .Z(n36168) );
  XOR U35995 ( .A(n36167), .B(n36171), .Z(n36169) );
  XNOR U35996 ( .A(n36172), .B(n36173), .Z(n36166) );
  NOR U35997 ( .A(n36174), .B(n36175), .Z(n36173) );
  XNOR U35998 ( .A(n36172), .B(n36176), .Z(n36174) );
  XOR U35999 ( .A(n36177), .B(n36178), .Z(n36121) );
  NOR U36000 ( .A(n36179), .B(n36180), .Z(n36178) );
  XNOR U36001 ( .A(n36177), .B(n36181), .Z(n36179) );
  XNOR U36002 ( .A(n36131), .B(n36122), .Z(n36165) );
  XOR U36003 ( .A(n36182), .B(n36183), .Z(n36122) );
  NOR U36004 ( .A(n36184), .B(n36185), .Z(n36183) );
  XNOR U36005 ( .A(n36182), .B(n36186), .Z(n36184) );
  XOR U36006 ( .A(n36187), .B(n36137), .Z(n36131) );
  XNOR U36007 ( .A(n36188), .B(n36189), .Z(n36137) );
  NOR U36008 ( .A(n36190), .B(n36191), .Z(n36189) );
  XNOR U36009 ( .A(n36188), .B(n36192), .Z(n36190) );
  XNOR U36010 ( .A(n36136), .B(n36128), .Z(n36187) );
  XOR U36011 ( .A(n36193), .B(n36194), .Z(n36128) );
  AND U36012 ( .A(n36195), .B(n36196), .Z(n36194) );
  XOR U36013 ( .A(n36193), .B(n36197), .Z(n36195) );
  XNOR U36014 ( .A(n36198), .B(n36133), .Z(n36136) );
  XOR U36015 ( .A(n36199), .B(n36200), .Z(n36133) );
  AND U36016 ( .A(n36201), .B(n36202), .Z(n36200) );
  XOR U36017 ( .A(n36199), .B(n36203), .Z(n36201) );
  XNOR U36018 ( .A(n36204), .B(n36205), .Z(n36198) );
  NOR U36019 ( .A(n36206), .B(n36207), .Z(n36205) );
  XOR U36020 ( .A(n36204), .B(n36208), .Z(n36206) );
  XOR U36021 ( .A(n36126), .B(n36138), .Z(n36164) );
  NOR U36022 ( .A(n36055), .B(n36209), .Z(n36138) );
  XNOR U36023 ( .A(n36144), .B(n36143), .Z(n36126) );
  XNOR U36024 ( .A(n36210), .B(n36149), .Z(n36143) );
  XOR U36025 ( .A(n36211), .B(n36212), .Z(n36149) );
  NOR U36026 ( .A(n36213), .B(n36214), .Z(n36212) );
  XNOR U36027 ( .A(n36211), .B(n36215), .Z(n36213) );
  XNOR U36028 ( .A(n36148), .B(n36140), .Z(n36210) );
  XOR U36029 ( .A(n36216), .B(n36217), .Z(n36140) );
  AND U36030 ( .A(n36218), .B(n36219), .Z(n36217) );
  XNOR U36031 ( .A(n36216), .B(n36220), .Z(n36218) );
  XNOR U36032 ( .A(n36221), .B(n36145), .Z(n36148) );
  XOR U36033 ( .A(n36222), .B(n36223), .Z(n36145) );
  AND U36034 ( .A(n36224), .B(n36225), .Z(n36223) );
  XOR U36035 ( .A(n36222), .B(n36226), .Z(n36224) );
  XNOR U36036 ( .A(n36227), .B(n36228), .Z(n36221) );
  NOR U36037 ( .A(n36229), .B(n36230), .Z(n36228) );
  XOR U36038 ( .A(n36227), .B(n36231), .Z(n36229) );
  XOR U36039 ( .A(n36154), .B(n36153), .Z(n36144) );
  XNOR U36040 ( .A(n36232), .B(n36150), .Z(n36153) );
  XOR U36041 ( .A(n36233), .B(n36234), .Z(n36150) );
  AND U36042 ( .A(n36235), .B(n36236), .Z(n36234) );
  XOR U36043 ( .A(n36233), .B(n36237), .Z(n36235) );
  XNOR U36044 ( .A(n36238), .B(n36239), .Z(n36232) );
  NOR U36045 ( .A(n36240), .B(n36241), .Z(n36239) );
  XNOR U36046 ( .A(n36238), .B(n36242), .Z(n36240) );
  XOR U36047 ( .A(n36243), .B(n36244), .Z(n36154) );
  NOR U36048 ( .A(n36245), .B(n36246), .Z(n36244) );
  XNOR U36049 ( .A(n36243), .B(n36247), .Z(n36245) );
  XNOR U36050 ( .A(n36046), .B(n36160), .Z(n36162) );
  XNOR U36051 ( .A(n36248), .B(n36249), .Z(n36046) );
  AND U36052 ( .A(n553), .B(n36250), .Z(n36249) );
  XNOR U36053 ( .A(n36251), .B(n36252), .Z(n36250) );
  AND U36054 ( .A(n36052), .B(n36055), .Z(n36160) );
  XOR U36055 ( .A(n36253), .B(n36209), .Z(n36055) );
  XNOR U36056 ( .A(p_input[2048]), .B(p_input[704]), .Z(n36209) );
  XOR U36057 ( .A(n36186), .B(n36185), .Z(n36253) );
  XOR U36058 ( .A(n36254), .B(n36197), .Z(n36185) );
  XOR U36059 ( .A(n36171), .B(n36170), .Z(n36197) );
  XNOR U36060 ( .A(n36255), .B(n36176), .Z(n36170) );
  XOR U36061 ( .A(p_input[2072]), .B(p_input[728]), .Z(n36176) );
  XOR U36062 ( .A(n36167), .B(n36175), .Z(n36255) );
  XOR U36063 ( .A(n36256), .B(n36172), .Z(n36175) );
  XOR U36064 ( .A(p_input[2070]), .B(p_input[726]), .Z(n36172) );
  XNOR U36065 ( .A(p_input[2071]), .B(p_input[727]), .Z(n36256) );
  XNOR U36066 ( .A(n28684), .B(p_input[722]), .Z(n36167) );
  XNOR U36067 ( .A(n36181), .B(n36180), .Z(n36171) );
  XOR U36068 ( .A(n36257), .B(n36177), .Z(n36180) );
  XOR U36069 ( .A(p_input[2067]), .B(p_input[723]), .Z(n36177) );
  XNOR U36070 ( .A(p_input[2068]), .B(p_input[724]), .Z(n36257) );
  XOR U36071 ( .A(p_input[2069]), .B(p_input[725]), .Z(n36181) );
  XNOR U36072 ( .A(n36196), .B(n36182), .Z(n36254) );
  XNOR U36073 ( .A(n28686), .B(p_input[705]), .Z(n36182) );
  XNOR U36074 ( .A(n36258), .B(n36203), .Z(n36196) );
  XNOR U36075 ( .A(n36192), .B(n36191), .Z(n36203) );
  XOR U36076 ( .A(n36259), .B(n36188), .Z(n36191) );
  XNOR U36077 ( .A(n28322), .B(p_input[730]), .Z(n36188) );
  XNOR U36078 ( .A(p_input[2075]), .B(p_input[731]), .Z(n36259) );
  XOR U36079 ( .A(p_input[2076]), .B(p_input[732]), .Z(n36192) );
  XNOR U36080 ( .A(n36202), .B(n36193), .Z(n36258) );
  XNOR U36081 ( .A(n28689), .B(p_input[721]), .Z(n36193) );
  XOR U36082 ( .A(n36260), .B(n36208), .Z(n36202) );
  XNOR U36083 ( .A(p_input[2079]), .B(p_input[735]), .Z(n36208) );
  XOR U36084 ( .A(n36199), .B(n36207), .Z(n36260) );
  XOR U36085 ( .A(n36261), .B(n36204), .Z(n36207) );
  XOR U36086 ( .A(p_input[2077]), .B(p_input[733]), .Z(n36204) );
  XNOR U36087 ( .A(p_input[2078]), .B(p_input[734]), .Z(n36261) );
  XNOR U36088 ( .A(n28326), .B(p_input[729]), .Z(n36199) );
  XNOR U36089 ( .A(n36220), .B(n36219), .Z(n36186) );
  XNOR U36090 ( .A(n36262), .B(n36226), .Z(n36219) );
  XNOR U36091 ( .A(n36215), .B(n36214), .Z(n36226) );
  XOR U36092 ( .A(n36263), .B(n36211), .Z(n36214) );
  XNOR U36093 ( .A(n28694), .B(p_input[715]), .Z(n36211) );
  XNOR U36094 ( .A(p_input[2060]), .B(p_input[716]), .Z(n36263) );
  XOR U36095 ( .A(p_input[2061]), .B(p_input[717]), .Z(n36215) );
  XNOR U36096 ( .A(n36225), .B(n36216), .Z(n36262) );
  XNOR U36097 ( .A(n28330), .B(p_input[706]), .Z(n36216) );
  XOR U36098 ( .A(n36264), .B(n36231), .Z(n36225) );
  XNOR U36099 ( .A(p_input[2064]), .B(p_input[720]), .Z(n36231) );
  XOR U36100 ( .A(n36222), .B(n36230), .Z(n36264) );
  XOR U36101 ( .A(n36265), .B(n36227), .Z(n36230) );
  XOR U36102 ( .A(p_input[2062]), .B(p_input[718]), .Z(n36227) );
  XNOR U36103 ( .A(p_input[2063]), .B(p_input[719]), .Z(n36265) );
  XNOR U36104 ( .A(n28697), .B(p_input[714]), .Z(n36222) );
  XNOR U36105 ( .A(n36237), .B(n36236), .Z(n36220) );
  XNOR U36106 ( .A(n36266), .B(n36242), .Z(n36236) );
  XOR U36107 ( .A(p_input[2057]), .B(p_input[713]), .Z(n36242) );
  XOR U36108 ( .A(n36233), .B(n36241), .Z(n36266) );
  XOR U36109 ( .A(n36267), .B(n36238), .Z(n36241) );
  XOR U36110 ( .A(p_input[2055]), .B(p_input[711]), .Z(n36238) );
  XNOR U36111 ( .A(p_input[2056]), .B(p_input[712]), .Z(n36267) );
  XNOR U36112 ( .A(n28337), .B(p_input[707]), .Z(n36233) );
  XNOR U36113 ( .A(n36247), .B(n36246), .Z(n36237) );
  XOR U36114 ( .A(n36268), .B(n36243), .Z(n36246) );
  XOR U36115 ( .A(p_input[2052]), .B(p_input[708]), .Z(n36243) );
  XNOR U36116 ( .A(p_input[2053]), .B(p_input[709]), .Z(n36268) );
  XOR U36117 ( .A(p_input[2054]), .B(p_input[710]), .Z(n36247) );
  XNOR U36118 ( .A(n36269), .B(n36270), .Z(n36052) );
  AND U36119 ( .A(n553), .B(n36271), .Z(n36270) );
  XNOR U36120 ( .A(n36272), .B(n36273), .Z(n553) );
  AND U36121 ( .A(n36274), .B(n36275), .Z(n36273) );
  XOR U36122 ( .A(n36066), .B(n36272), .Z(n36275) );
  XNOR U36123 ( .A(n36276), .B(n36272), .Z(n36274) );
  XOR U36124 ( .A(n36277), .B(n36278), .Z(n36272) );
  AND U36125 ( .A(n36279), .B(n36280), .Z(n36278) );
  XOR U36126 ( .A(n36081), .B(n36277), .Z(n36280) );
  XOR U36127 ( .A(n36277), .B(n36082), .Z(n36279) );
  XOR U36128 ( .A(n36281), .B(n36282), .Z(n36277) );
  AND U36129 ( .A(n36283), .B(n36284), .Z(n36282) );
  XOR U36130 ( .A(n36109), .B(n36281), .Z(n36284) );
  XOR U36131 ( .A(n36281), .B(n36110), .Z(n36283) );
  XOR U36132 ( .A(n36285), .B(n36286), .Z(n36281) );
  AND U36133 ( .A(n36287), .B(n36288), .Z(n36286) );
  XOR U36134 ( .A(n36158), .B(n36285), .Z(n36288) );
  XOR U36135 ( .A(n36285), .B(n36159), .Z(n36287) );
  XOR U36136 ( .A(n36289), .B(n36290), .Z(n36285) );
  AND U36137 ( .A(n36291), .B(n36292), .Z(n36290) );
  XOR U36138 ( .A(n36289), .B(n36251), .Z(n36292) );
  XNOR U36139 ( .A(n36293), .B(n36294), .Z(n36002) );
  AND U36140 ( .A(n557), .B(n36295), .Z(n36294) );
  XNOR U36141 ( .A(n36296), .B(n36297), .Z(n557) );
  AND U36142 ( .A(n36298), .B(n36299), .Z(n36297) );
  XOR U36143 ( .A(n36296), .B(n36012), .Z(n36299) );
  XNOR U36144 ( .A(n36296), .B(n35962), .Z(n36298) );
  XOR U36145 ( .A(n36300), .B(n36301), .Z(n36296) );
  AND U36146 ( .A(n36302), .B(n36303), .Z(n36301) );
  XNOR U36147 ( .A(n36022), .B(n36300), .Z(n36303) );
  XOR U36148 ( .A(n36300), .B(n35972), .Z(n36302) );
  XOR U36149 ( .A(n36304), .B(n36305), .Z(n36300) );
  AND U36150 ( .A(n36306), .B(n36307), .Z(n36305) );
  XNOR U36151 ( .A(n36032), .B(n36304), .Z(n36307) );
  XOR U36152 ( .A(n36304), .B(n35981), .Z(n36306) );
  XOR U36153 ( .A(n36308), .B(n36309), .Z(n36304) );
  AND U36154 ( .A(n36310), .B(n36311), .Z(n36309) );
  XOR U36155 ( .A(n36308), .B(n35989), .Z(n36310) );
  XOR U36156 ( .A(n36312), .B(n36313), .Z(n35953) );
  AND U36157 ( .A(n561), .B(n36295), .Z(n36313) );
  XNOR U36158 ( .A(n36293), .B(n36312), .Z(n36295) );
  XNOR U36159 ( .A(n36314), .B(n36315), .Z(n561) );
  AND U36160 ( .A(n36316), .B(n36317), .Z(n36315) );
  XNOR U36161 ( .A(n36318), .B(n36314), .Z(n36317) );
  IV U36162 ( .A(n36012), .Z(n36318) );
  XOR U36163 ( .A(n36276), .B(n36319), .Z(n36012) );
  AND U36164 ( .A(n564), .B(n36320), .Z(n36319) );
  XOR U36165 ( .A(n36065), .B(n36062), .Z(n36320) );
  IV U36166 ( .A(n36276), .Z(n36065) );
  XNOR U36167 ( .A(n35962), .B(n36314), .Z(n36316) );
  XOR U36168 ( .A(n36321), .B(n36322), .Z(n35962) );
  AND U36169 ( .A(n580), .B(n36323), .Z(n36322) );
  XOR U36170 ( .A(n36324), .B(n36325), .Z(n36314) );
  AND U36171 ( .A(n36326), .B(n36327), .Z(n36325) );
  XNOR U36172 ( .A(n36324), .B(n36022), .Z(n36327) );
  XOR U36173 ( .A(n36082), .B(n36328), .Z(n36022) );
  AND U36174 ( .A(n564), .B(n36329), .Z(n36328) );
  XOR U36175 ( .A(n36078), .B(n36082), .Z(n36329) );
  XNOR U36176 ( .A(n36330), .B(n36324), .Z(n36326) );
  IV U36177 ( .A(n35972), .Z(n36330) );
  XOR U36178 ( .A(n36331), .B(n36332), .Z(n35972) );
  AND U36179 ( .A(n580), .B(n36333), .Z(n36332) );
  XOR U36180 ( .A(n36334), .B(n36335), .Z(n36324) );
  AND U36181 ( .A(n36336), .B(n36337), .Z(n36335) );
  XNOR U36182 ( .A(n36334), .B(n36032), .Z(n36337) );
  XOR U36183 ( .A(n36110), .B(n36338), .Z(n36032) );
  AND U36184 ( .A(n564), .B(n36339), .Z(n36338) );
  XOR U36185 ( .A(n36106), .B(n36110), .Z(n36339) );
  XOR U36186 ( .A(n35981), .B(n36334), .Z(n36336) );
  XOR U36187 ( .A(n36340), .B(n36341), .Z(n35981) );
  AND U36188 ( .A(n580), .B(n36342), .Z(n36341) );
  XOR U36189 ( .A(n36308), .B(n36343), .Z(n36334) );
  AND U36190 ( .A(n36344), .B(n36311), .Z(n36343) );
  XNOR U36191 ( .A(n36042), .B(n36308), .Z(n36311) );
  XOR U36192 ( .A(n36159), .B(n36345), .Z(n36042) );
  AND U36193 ( .A(n564), .B(n36346), .Z(n36345) );
  XOR U36194 ( .A(n36155), .B(n36159), .Z(n36346) );
  XNOR U36195 ( .A(n36347), .B(n36308), .Z(n36344) );
  IV U36196 ( .A(n35989), .Z(n36347) );
  XOR U36197 ( .A(n36348), .B(n36349), .Z(n35989) );
  AND U36198 ( .A(n580), .B(n36350), .Z(n36349) );
  XOR U36199 ( .A(n36351), .B(n36352), .Z(n36308) );
  AND U36200 ( .A(n36353), .B(n36354), .Z(n36352) );
  XNOR U36201 ( .A(n36351), .B(n36050), .Z(n36354) );
  XOR U36202 ( .A(n36252), .B(n36355), .Z(n36050) );
  AND U36203 ( .A(n564), .B(n36356), .Z(n36355) );
  XOR U36204 ( .A(n36248), .B(n36252), .Z(n36356) );
  XNOR U36205 ( .A(n36357), .B(n36351), .Z(n36353) );
  IV U36206 ( .A(n35999), .Z(n36357) );
  XOR U36207 ( .A(n36358), .B(n36359), .Z(n35999) );
  AND U36208 ( .A(n580), .B(n36360), .Z(n36359) );
  AND U36209 ( .A(n36312), .B(n36293), .Z(n36351) );
  XNOR U36210 ( .A(n36361), .B(n36362), .Z(n36293) );
  AND U36211 ( .A(n564), .B(n36271), .Z(n36362) );
  XNOR U36212 ( .A(n36269), .B(n36361), .Z(n36271) );
  XNOR U36213 ( .A(n36363), .B(n36364), .Z(n564) );
  AND U36214 ( .A(n36365), .B(n36366), .Z(n36364) );
  XNOR U36215 ( .A(n36363), .B(n36062), .Z(n36366) );
  IV U36216 ( .A(n36066), .Z(n36062) );
  XOR U36217 ( .A(n36367), .B(n36368), .Z(n36066) );
  AND U36218 ( .A(n568), .B(n36369), .Z(n36368) );
  XOR U36219 ( .A(n36370), .B(n36367), .Z(n36369) );
  XNOR U36220 ( .A(n36363), .B(n36276), .Z(n36365) );
  XOR U36221 ( .A(n36371), .B(n36372), .Z(n36276) );
  AND U36222 ( .A(n576), .B(n36323), .Z(n36372) );
  XOR U36223 ( .A(n36321), .B(n36371), .Z(n36323) );
  XOR U36224 ( .A(n36373), .B(n36374), .Z(n36363) );
  AND U36225 ( .A(n36375), .B(n36376), .Z(n36374) );
  XNOR U36226 ( .A(n36373), .B(n36078), .Z(n36376) );
  IV U36227 ( .A(n36081), .Z(n36078) );
  XOR U36228 ( .A(n36377), .B(n36378), .Z(n36081) );
  AND U36229 ( .A(n568), .B(n36379), .Z(n36378) );
  XOR U36230 ( .A(n36380), .B(n36377), .Z(n36379) );
  XOR U36231 ( .A(n36082), .B(n36373), .Z(n36375) );
  XOR U36232 ( .A(n36381), .B(n36382), .Z(n36082) );
  AND U36233 ( .A(n576), .B(n36333), .Z(n36382) );
  XOR U36234 ( .A(n36381), .B(n36331), .Z(n36333) );
  XOR U36235 ( .A(n36383), .B(n36384), .Z(n36373) );
  AND U36236 ( .A(n36385), .B(n36386), .Z(n36384) );
  XNOR U36237 ( .A(n36383), .B(n36106), .Z(n36386) );
  IV U36238 ( .A(n36109), .Z(n36106) );
  XOR U36239 ( .A(n36387), .B(n36388), .Z(n36109) );
  AND U36240 ( .A(n568), .B(n36389), .Z(n36388) );
  XNOR U36241 ( .A(n36390), .B(n36387), .Z(n36389) );
  XOR U36242 ( .A(n36110), .B(n36383), .Z(n36385) );
  XOR U36243 ( .A(n36391), .B(n36392), .Z(n36110) );
  AND U36244 ( .A(n576), .B(n36342), .Z(n36392) );
  XOR U36245 ( .A(n36391), .B(n36340), .Z(n36342) );
  XOR U36246 ( .A(n36393), .B(n36394), .Z(n36383) );
  AND U36247 ( .A(n36395), .B(n36396), .Z(n36394) );
  XNOR U36248 ( .A(n36393), .B(n36155), .Z(n36396) );
  IV U36249 ( .A(n36158), .Z(n36155) );
  XOR U36250 ( .A(n36397), .B(n36398), .Z(n36158) );
  AND U36251 ( .A(n568), .B(n36399), .Z(n36398) );
  XOR U36252 ( .A(n36400), .B(n36397), .Z(n36399) );
  XOR U36253 ( .A(n36159), .B(n36393), .Z(n36395) );
  XOR U36254 ( .A(n36401), .B(n36402), .Z(n36159) );
  AND U36255 ( .A(n576), .B(n36350), .Z(n36402) );
  XOR U36256 ( .A(n36401), .B(n36348), .Z(n36350) );
  XOR U36257 ( .A(n36289), .B(n36403), .Z(n36393) );
  AND U36258 ( .A(n36291), .B(n36404), .Z(n36403) );
  XNOR U36259 ( .A(n36289), .B(n36248), .Z(n36404) );
  IV U36260 ( .A(n36251), .Z(n36248) );
  XOR U36261 ( .A(n36405), .B(n36406), .Z(n36251) );
  AND U36262 ( .A(n568), .B(n36407), .Z(n36406) );
  XNOR U36263 ( .A(n36408), .B(n36405), .Z(n36407) );
  XOR U36264 ( .A(n36252), .B(n36289), .Z(n36291) );
  XOR U36265 ( .A(n36409), .B(n36410), .Z(n36252) );
  AND U36266 ( .A(n576), .B(n36360), .Z(n36410) );
  XOR U36267 ( .A(n36409), .B(n36358), .Z(n36360) );
  AND U36268 ( .A(n36361), .B(n36269), .Z(n36289) );
  XNOR U36269 ( .A(n36411), .B(n36412), .Z(n36269) );
  AND U36270 ( .A(n568), .B(n36413), .Z(n36412) );
  XNOR U36271 ( .A(n36414), .B(n36411), .Z(n36413) );
  XNOR U36272 ( .A(n36415), .B(n36416), .Z(n568) );
  AND U36273 ( .A(n36417), .B(n36418), .Z(n36416) );
  XOR U36274 ( .A(n36370), .B(n36415), .Z(n36418) );
  AND U36275 ( .A(n36419), .B(n36420), .Z(n36370) );
  XNOR U36276 ( .A(n36367), .B(n36415), .Z(n36417) );
  XNOR U36277 ( .A(n36421), .B(n36422), .Z(n36367) );
  AND U36278 ( .A(n572), .B(n36423), .Z(n36422) );
  XNOR U36279 ( .A(n36424), .B(n36425), .Z(n36423) );
  XOR U36280 ( .A(n36426), .B(n36427), .Z(n36415) );
  AND U36281 ( .A(n36428), .B(n36429), .Z(n36427) );
  XNOR U36282 ( .A(n36426), .B(n36419), .Z(n36429) );
  IV U36283 ( .A(n36380), .Z(n36419) );
  XOR U36284 ( .A(n36430), .B(n36431), .Z(n36380) );
  XOR U36285 ( .A(n36432), .B(n36420), .Z(n36431) );
  AND U36286 ( .A(n36390), .B(n36433), .Z(n36420) );
  AND U36287 ( .A(n36434), .B(n36435), .Z(n36432) );
  XOR U36288 ( .A(n36436), .B(n36430), .Z(n36434) );
  XNOR U36289 ( .A(n36377), .B(n36426), .Z(n36428) );
  XNOR U36290 ( .A(n36437), .B(n36438), .Z(n36377) );
  AND U36291 ( .A(n572), .B(n36439), .Z(n36438) );
  XNOR U36292 ( .A(n36440), .B(n36441), .Z(n36439) );
  XOR U36293 ( .A(n36442), .B(n36443), .Z(n36426) );
  AND U36294 ( .A(n36444), .B(n36445), .Z(n36443) );
  XNOR U36295 ( .A(n36442), .B(n36390), .Z(n36445) );
  XOR U36296 ( .A(n36446), .B(n36435), .Z(n36390) );
  XNOR U36297 ( .A(n36447), .B(n36430), .Z(n36435) );
  XOR U36298 ( .A(n36448), .B(n36449), .Z(n36430) );
  AND U36299 ( .A(n36450), .B(n36451), .Z(n36449) );
  XOR U36300 ( .A(n36452), .B(n36448), .Z(n36450) );
  XNOR U36301 ( .A(n36453), .B(n36454), .Z(n36447) );
  AND U36302 ( .A(n36455), .B(n36456), .Z(n36454) );
  XOR U36303 ( .A(n36453), .B(n36457), .Z(n36455) );
  XNOR U36304 ( .A(n36436), .B(n36433), .Z(n36446) );
  AND U36305 ( .A(n36458), .B(n36459), .Z(n36433) );
  XOR U36306 ( .A(n36460), .B(n36461), .Z(n36436) );
  AND U36307 ( .A(n36462), .B(n36463), .Z(n36461) );
  XOR U36308 ( .A(n36460), .B(n36464), .Z(n36462) );
  XNOR U36309 ( .A(n36387), .B(n36442), .Z(n36444) );
  XNOR U36310 ( .A(n36465), .B(n36466), .Z(n36387) );
  AND U36311 ( .A(n572), .B(n36467), .Z(n36466) );
  XNOR U36312 ( .A(n36468), .B(n36469), .Z(n36467) );
  XOR U36313 ( .A(n36470), .B(n36471), .Z(n36442) );
  AND U36314 ( .A(n36472), .B(n36473), .Z(n36471) );
  XNOR U36315 ( .A(n36470), .B(n36458), .Z(n36473) );
  IV U36316 ( .A(n36400), .Z(n36458) );
  XNOR U36317 ( .A(n36474), .B(n36451), .Z(n36400) );
  XNOR U36318 ( .A(n36475), .B(n36457), .Z(n36451) );
  XOR U36319 ( .A(n36476), .B(n36477), .Z(n36457) );
  AND U36320 ( .A(n36478), .B(n36479), .Z(n36477) );
  XOR U36321 ( .A(n36476), .B(n36480), .Z(n36478) );
  XNOR U36322 ( .A(n36456), .B(n36448), .Z(n36475) );
  XOR U36323 ( .A(n36481), .B(n36482), .Z(n36448) );
  AND U36324 ( .A(n36483), .B(n36484), .Z(n36482) );
  XNOR U36325 ( .A(n36485), .B(n36481), .Z(n36483) );
  XNOR U36326 ( .A(n36486), .B(n36453), .Z(n36456) );
  XOR U36327 ( .A(n36487), .B(n36488), .Z(n36453) );
  AND U36328 ( .A(n36489), .B(n36490), .Z(n36488) );
  XOR U36329 ( .A(n36487), .B(n36491), .Z(n36489) );
  XNOR U36330 ( .A(n36492), .B(n36493), .Z(n36486) );
  AND U36331 ( .A(n36494), .B(n36495), .Z(n36493) );
  XNOR U36332 ( .A(n36492), .B(n36496), .Z(n36494) );
  XNOR U36333 ( .A(n36452), .B(n36459), .Z(n36474) );
  AND U36334 ( .A(n36408), .B(n36497), .Z(n36459) );
  XOR U36335 ( .A(n36464), .B(n36463), .Z(n36452) );
  XNOR U36336 ( .A(n36498), .B(n36460), .Z(n36463) );
  XOR U36337 ( .A(n36499), .B(n36500), .Z(n36460) );
  AND U36338 ( .A(n36501), .B(n36502), .Z(n36500) );
  XOR U36339 ( .A(n36499), .B(n36503), .Z(n36501) );
  XNOR U36340 ( .A(n36504), .B(n36505), .Z(n36498) );
  AND U36341 ( .A(n36506), .B(n36507), .Z(n36505) );
  XOR U36342 ( .A(n36504), .B(n36508), .Z(n36506) );
  XOR U36343 ( .A(n36509), .B(n36510), .Z(n36464) );
  AND U36344 ( .A(n36511), .B(n36512), .Z(n36510) );
  XOR U36345 ( .A(n36509), .B(n36513), .Z(n36511) );
  XNOR U36346 ( .A(n36397), .B(n36470), .Z(n36472) );
  XNOR U36347 ( .A(n36514), .B(n36515), .Z(n36397) );
  AND U36348 ( .A(n572), .B(n36516), .Z(n36515) );
  XNOR U36349 ( .A(n36517), .B(n36518), .Z(n36516) );
  XOR U36350 ( .A(n36519), .B(n36520), .Z(n36470) );
  AND U36351 ( .A(n36521), .B(n36522), .Z(n36520) );
  XNOR U36352 ( .A(n36519), .B(n36408), .Z(n36522) );
  XOR U36353 ( .A(n36523), .B(n36484), .Z(n36408) );
  XNOR U36354 ( .A(n36524), .B(n36491), .Z(n36484) );
  XOR U36355 ( .A(n36480), .B(n36479), .Z(n36491) );
  XNOR U36356 ( .A(n36525), .B(n36476), .Z(n36479) );
  XOR U36357 ( .A(n36526), .B(n36527), .Z(n36476) );
  AND U36358 ( .A(n36528), .B(n36529), .Z(n36527) );
  XOR U36359 ( .A(n36526), .B(n36530), .Z(n36528) );
  XNOR U36360 ( .A(n36531), .B(n36532), .Z(n36525) );
  NOR U36361 ( .A(n36533), .B(n36534), .Z(n36532) );
  XNOR U36362 ( .A(n36531), .B(n36535), .Z(n36533) );
  XOR U36363 ( .A(n36536), .B(n36537), .Z(n36480) );
  NOR U36364 ( .A(n36538), .B(n36539), .Z(n36537) );
  XNOR U36365 ( .A(n36536), .B(n36540), .Z(n36538) );
  XNOR U36366 ( .A(n36490), .B(n36481), .Z(n36524) );
  XOR U36367 ( .A(n36541), .B(n36542), .Z(n36481) );
  NOR U36368 ( .A(n36543), .B(n36544), .Z(n36542) );
  XNOR U36369 ( .A(n36541), .B(n36545), .Z(n36543) );
  XOR U36370 ( .A(n36546), .B(n36496), .Z(n36490) );
  XNOR U36371 ( .A(n36547), .B(n36548), .Z(n36496) );
  NOR U36372 ( .A(n36549), .B(n36550), .Z(n36548) );
  XNOR U36373 ( .A(n36547), .B(n36551), .Z(n36549) );
  XNOR U36374 ( .A(n36495), .B(n36487), .Z(n36546) );
  XOR U36375 ( .A(n36552), .B(n36553), .Z(n36487) );
  AND U36376 ( .A(n36554), .B(n36555), .Z(n36553) );
  XOR U36377 ( .A(n36552), .B(n36556), .Z(n36554) );
  XNOR U36378 ( .A(n36557), .B(n36492), .Z(n36495) );
  XOR U36379 ( .A(n36558), .B(n36559), .Z(n36492) );
  AND U36380 ( .A(n36560), .B(n36561), .Z(n36559) );
  XOR U36381 ( .A(n36558), .B(n36562), .Z(n36560) );
  XNOR U36382 ( .A(n36563), .B(n36564), .Z(n36557) );
  NOR U36383 ( .A(n36565), .B(n36566), .Z(n36564) );
  XOR U36384 ( .A(n36563), .B(n36567), .Z(n36565) );
  XOR U36385 ( .A(n36485), .B(n36497), .Z(n36523) );
  NOR U36386 ( .A(n36414), .B(n36568), .Z(n36497) );
  XNOR U36387 ( .A(n36503), .B(n36502), .Z(n36485) );
  XNOR U36388 ( .A(n36569), .B(n36508), .Z(n36502) );
  XOR U36389 ( .A(n36570), .B(n36571), .Z(n36508) );
  NOR U36390 ( .A(n36572), .B(n36573), .Z(n36571) );
  XNOR U36391 ( .A(n36570), .B(n36574), .Z(n36572) );
  XNOR U36392 ( .A(n36507), .B(n36499), .Z(n36569) );
  XOR U36393 ( .A(n36575), .B(n36576), .Z(n36499) );
  AND U36394 ( .A(n36577), .B(n36578), .Z(n36576) );
  XNOR U36395 ( .A(n36575), .B(n36579), .Z(n36577) );
  XNOR U36396 ( .A(n36580), .B(n36504), .Z(n36507) );
  XOR U36397 ( .A(n36581), .B(n36582), .Z(n36504) );
  AND U36398 ( .A(n36583), .B(n36584), .Z(n36582) );
  XOR U36399 ( .A(n36581), .B(n36585), .Z(n36583) );
  XNOR U36400 ( .A(n36586), .B(n36587), .Z(n36580) );
  NOR U36401 ( .A(n36588), .B(n36589), .Z(n36587) );
  XOR U36402 ( .A(n36586), .B(n36590), .Z(n36588) );
  XOR U36403 ( .A(n36513), .B(n36512), .Z(n36503) );
  XNOR U36404 ( .A(n36591), .B(n36509), .Z(n36512) );
  XOR U36405 ( .A(n36592), .B(n36593), .Z(n36509) );
  AND U36406 ( .A(n36594), .B(n36595), .Z(n36593) );
  XOR U36407 ( .A(n36592), .B(n36596), .Z(n36594) );
  XNOR U36408 ( .A(n36597), .B(n36598), .Z(n36591) );
  NOR U36409 ( .A(n36599), .B(n36600), .Z(n36598) );
  XNOR U36410 ( .A(n36597), .B(n36601), .Z(n36599) );
  XOR U36411 ( .A(n36602), .B(n36603), .Z(n36513) );
  NOR U36412 ( .A(n36604), .B(n36605), .Z(n36603) );
  XNOR U36413 ( .A(n36602), .B(n36606), .Z(n36604) );
  XNOR U36414 ( .A(n36405), .B(n36519), .Z(n36521) );
  XNOR U36415 ( .A(n36607), .B(n36608), .Z(n36405) );
  AND U36416 ( .A(n572), .B(n36609), .Z(n36608) );
  XNOR U36417 ( .A(n36610), .B(n36611), .Z(n36609) );
  AND U36418 ( .A(n36411), .B(n36414), .Z(n36519) );
  XOR U36419 ( .A(n36612), .B(n36568), .Z(n36414) );
  XNOR U36420 ( .A(p_input[2048]), .B(p_input[736]), .Z(n36568) );
  XOR U36421 ( .A(n36545), .B(n36544), .Z(n36612) );
  XOR U36422 ( .A(n36613), .B(n36556), .Z(n36544) );
  XOR U36423 ( .A(n36530), .B(n36529), .Z(n36556) );
  XNOR U36424 ( .A(n36614), .B(n36535), .Z(n36529) );
  XOR U36425 ( .A(p_input[2072]), .B(p_input[760]), .Z(n36535) );
  XOR U36426 ( .A(n36526), .B(n36534), .Z(n36614) );
  XOR U36427 ( .A(n36615), .B(n36531), .Z(n36534) );
  XOR U36428 ( .A(p_input[2070]), .B(p_input[758]), .Z(n36531) );
  XNOR U36429 ( .A(p_input[2071]), .B(p_input[759]), .Z(n36615) );
  XNOR U36430 ( .A(n28684), .B(p_input[754]), .Z(n36526) );
  XNOR U36431 ( .A(n36540), .B(n36539), .Z(n36530) );
  XOR U36432 ( .A(n36616), .B(n36536), .Z(n36539) );
  XOR U36433 ( .A(p_input[2067]), .B(p_input[755]), .Z(n36536) );
  XNOR U36434 ( .A(p_input[2068]), .B(p_input[756]), .Z(n36616) );
  XOR U36435 ( .A(p_input[2069]), .B(p_input[757]), .Z(n36540) );
  XNOR U36436 ( .A(n36555), .B(n36541), .Z(n36613) );
  XNOR U36437 ( .A(n28686), .B(p_input[737]), .Z(n36541) );
  XNOR U36438 ( .A(n36617), .B(n36562), .Z(n36555) );
  XNOR U36439 ( .A(n36551), .B(n36550), .Z(n36562) );
  XOR U36440 ( .A(n36618), .B(n36547), .Z(n36550) );
  XNOR U36441 ( .A(n28322), .B(p_input[762]), .Z(n36547) );
  XNOR U36442 ( .A(p_input[2075]), .B(p_input[763]), .Z(n36618) );
  XOR U36443 ( .A(p_input[2076]), .B(p_input[764]), .Z(n36551) );
  XNOR U36444 ( .A(n36561), .B(n36552), .Z(n36617) );
  XNOR U36445 ( .A(n28689), .B(p_input[753]), .Z(n36552) );
  XOR U36446 ( .A(n36619), .B(n36567), .Z(n36561) );
  XNOR U36447 ( .A(p_input[2079]), .B(p_input[767]), .Z(n36567) );
  XOR U36448 ( .A(n36558), .B(n36566), .Z(n36619) );
  XOR U36449 ( .A(n36620), .B(n36563), .Z(n36566) );
  XOR U36450 ( .A(p_input[2077]), .B(p_input[765]), .Z(n36563) );
  XNOR U36451 ( .A(p_input[2078]), .B(p_input[766]), .Z(n36620) );
  XNOR U36452 ( .A(n28326), .B(p_input[761]), .Z(n36558) );
  XNOR U36453 ( .A(n36579), .B(n36578), .Z(n36545) );
  XNOR U36454 ( .A(n36621), .B(n36585), .Z(n36578) );
  XNOR U36455 ( .A(n36574), .B(n36573), .Z(n36585) );
  XOR U36456 ( .A(n36622), .B(n36570), .Z(n36573) );
  XNOR U36457 ( .A(n28694), .B(p_input[747]), .Z(n36570) );
  XNOR U36458 ( .A(p_input[2060]), .B(p_input[748]), .Z(n36622) );
  XOR U36459 ( .A(p_input[2061]), .B(p_input[749]), .Z(n36574) );
  XNOR U36460 ( .A(n36584), .B(n36575), .Z(n36621) );
  XNOR U36461 ( .A(n28330), .B(p_input[738]), .Z(n36575) );
  XOR U36462 ( .A(n36623), .B(n36590), .Z(n36584) );
  XNOR U36463 ( .A(p_input[2064]), .B(p_input[752]), .Z(n36590) );
  XOR U36464 ( .A(n36581), .B(n36589), .Z(n36623) );
  XOR U36465 ( .A(n36624), .B(n36586), .Z(n36589) );
  XOR U36466 ( .A(p_input[2062]), .B(p_input[750]), .Z(n36586) );
  XNOR U36467 ( .A(p_input[2063]), .B(p_input[751]), .Z(n36624) );
  XNOR U36468 ( .A(n28697), .B(p_input[746]), .Z(n36581) );
  XNOR U36469 ( .A(n36596), .B(n36595), .Z(n36579) );
  XNOR U36470 ( .A(n36625), .B(n36601), .Z(n36595) );
  XOR U36471 ( .A(p_input[2057]), .B(p_input[745]), .Z(n36601) );
  XOR U36472 ( .A(n36592), .B(n36600), .Z(n36625) );
  XOR U36473 ( .A(n36626), .B(n36597), .Z(n36600) );
  XOR U36474 ( .A(p_input[2055]), .B(p_input[743]), .Z(n36597) );
  XNOR U36475 ( .A(p_input[2056]), .B(p_input[744]), .Z(n36626) );
  XNOR U36476 ( .A(n28337), .B(p_input[739]), .Z(n36592) );
  XNOR U36477 ( .A(n36606), .B(n36605), .Z(n36596) );
  XOR U36478 ( .A(n36627), .B(n36602), .Z(n36605) );
  XOR U36479 ( .A(p_input[2052]), .B(p_input[740]), .Z(n36602) );
  XNOR U36480 ( .A(p_input[2053]), .B(p_input[741]), .Z(n36627) );
  XOR U36481 ( .A(p_input[2054]), .B(p_input[742]), .Z(n36606) );
  XNOR U36482 ( .A(n36628), .B(n36629), .Z(n36411) );
  AND U36483 ( .A(n572), .B(n36630), .Z(n36629) );
  XNOR U36484 ( .A(n36631), .B(n36632), .Z(n572) );
  AND U36485 ( .A(n36633), .B(n36634), .Z(n36632) );
  XOR U36486 ( .A(n36425), .B(n36631), .Z(n36634) );
  XNOR U36487 ( .A(n36635), .B(n36631), .Z(n36633) );
  XOR U36488 ( .A(n36636), .B(n36637), .Z(n36631) );
  AND U36489 ( .A(n36638), .B(n36639), .Z(n36637) );
  XOR U36490 ( .A(n36440), .B(n36636), .Z(n36639) );
  XOR U36491 ( .A(n36636), .B(n36441), .Z(n36638) );
  XOR U36492 ( .A(n36640), .B(n36641), .Z(n36636) );
  AND U36493 ( .A(n36642), .B(n36643), .Z(n36641) );
  XOR U36494 ( .A(n36468), .B(n36640), .Z(n36643) );
  XOR U36495 ( .A(n36640), .B(n36469), .Z(n36642) );
  XOR U36496 ( .A(n36644), .B(n36645), .Z(n36640) );
  AND U36497 ( .A(n36646), .B(n36647), .Z(n36645) );
  XOR U36498 ( .A(n36517), .B(n36644), .Z(n36647) );
  XOR U36499 ( .A(n36644), .B(n36518), .Z(n36646) );
  XOR U36500 ( .A(n36648), .B(n36649), .Z(n36644) );
  AND U36501 ( .A(n36650), .B(n36651), .Z(n36649) );
  XOR U36502 ( .A(n36648), .B(n36610), .Z(n36651) );
  XNOR U36503 ( .A(n36652), .B(n36653), .Z(n36361) );
  AND U36504 ( .A(n576), .B(n36654), .Z(n36653) );
  XNOR U36505 ( .A(n36655), .B(n36656), .Z(n576) );
  AND U36506 ( .A(n36657), .B(n36658), .Z(n36656) );
  XOR U36507 ( .A(n36655), .B(n36371), .Z(n36658) );
  XNOR U36508 ( .A(n36655), .B(n36321), .Z(n36657) );
  XOR U36509 ( .A(n36659), .B(n36660), .Z(n36655) );
  AND U36510 ( .A(n36661), .B(n36662), .Z(n36660) );
  XNOR U36511 ( .A(n36381), .B(n36659), .Z(n36662) );
  XOR U36512 ( .A(n36659), .B(n36331), .Z(n36661) );
  XOR U36513 ( .A(n36663), .B(n36664), .Z(n36659) );
  AND U36514 ( .A(n36665), .B(n36666), .Z(n36664) );
  XNOR U36515 ( .A(n36391), .B(n36663), .Z(n36666) );
  XOR U36516 ( .A(n36663), .B(n36340), .Z(n36665) );
  XOR U36517 ( .A(n36667), .B(n36668), .Z(n36663) );
  AND U36518 ( .A(n36669), .B(n36670), .Z(n36668) );
  XOR U36519 ( .A(n36667), .B(n36348), .Z(n36669) );
  XOR U36520 ( .A(n36671), .B(n36672), .Z(n36312) );
  AND U36521 ( .A(n580), .B(n36654), .Z(n36672) );
  XNOR U36522 ( .A(n36652), .B(n36671), .Z(n36654) );
  XNOR U36523 ( .A(n36673), .B(n36674), .Z(n580) );
  AND U36524 ( .A(n36675), .B(n36676), .Z(n36674) );
  XNOR U36525 ( .A(n36677), .B(n36673), .Z(n36676) );
  IV U36526 ( .A(n36371), .Z(n36677) );
  XOR U36527 ( .A(n36635), .B(n36678), .Z(n36371) );
  AND U36528 ( .A(n583), .B(n36679), .Z(n36678) );
  XOR U36529 ( .A(n36424), .B(n36421), .Z(n36679) );
  IV U36530 ( .A(n36635), .Z(n36424) );
  XNOR U36531 ( .A(n36321), .B(n36673), .Z(n36675) );
  XOR U36532 ( .A(n36680), .B(n36681), .Z(n36321) );
  AND U36533 ( .A(n599), .B(n36682), .Z(n36681) );
  XOR U36534 ( .A(n36683), .B(n36684), .Z(n36673) );
  AND U36535 ( .A(n36685), .B(n36686), .Z(n36684) );
  XNOR U36536 ( .A(n36683), .B(n36381), .Z(n36686) );
  XOR U36537 ( .A(n36441), .B(n36687), .Z(n36381) );
  AND U36538 ( .A(n583), .B(n36688), .Z(n36687) );
  XOR U36539 ( .A(n36437), .B(n36441), .Z(n36688) );
  XNOR U36540 ( .A(n36689), .B(n36683), .Z(n36685) );
  IV U36541 ( .A(n36331), .Z(n36689) );
  XOR U36542 ( .A(n36690), .B(n36691), .Z(n36331) );
  AND U36543 ( .A(n599), .B(n36692), .Z(n36691) );
  XOR U36544 ( .A(n36693), .B(n36694), .Z(n36683) );
  AND U36545 ( .A(n36695), .B(n36696), .Z(n36694) );
  XNOR U36546 ( .A(n36693), .B(n36391), .Z(n36696) );
  XOR U36547 ( .A(n36469), .B(n36697), .Z(n36391) );
  AND U36548 ( .A(n583), .B(n36698), .Z(n36697) );
  XOR U36549 ( .A(n36465), .B(n36469), .Z(n36698) );
  XOR U36550 ( .A(n36340), .B(n36693), .Z(n36695) );
  XOR U36551 ( .A(n36699), .B(n36700), .Z(n36340) );
  AND U36552 ( .A(n599), .B(n36701), .Z(n36700) );
  XOR U36553 ( .A(n36667), .B(n36702), .Z(n36693) );
  AND U36554 ( .A(n36703), .B(n36670), .Z(n36702) );
  XNOR U36555 ( .A(n36401), .B(n36667), .Z(n36670) );
  XOR U36556 ( .A(n36518), .B(n36704), .Z(n36401) );
  AND U36557 ( .A(n583), .B(n36705), .Z(n36704) );
  XOR U36558 ( .A(n36514), .B(n36518), .Z(n36705) );
  XNOR U36559 ( .A(n36706), .B(n36667), .Z(n36703) );
  IV U36560 ( .A(n36348), .Z(n36706) );
  XOR U36561 ( .A(n36707), .B(n36708), .Z(n36348) );
  AND U36562 ( .A(n599), .B(n36709), .Z(n36708) );
  XOR U36563 ( .A(n36710), .B(n36711), .Z(n36667) );
  AND U36564 ( .A(n36712), .B(n36713), .Z(n36711) );
  XNOR U36565 ( .A(n36710), .B(n36409), .Z(n36713) );
  XOR U36566 ( .A(n36611), .B(n36714), .Z(n36409) );
  AND U36567 ( .A(n583), .B(n36715), .Z(n36714) );
  XOR U36568 ( .A(n36607), .B(n36611), .Z(n36715) );
  XNOR U36569 ( .A(n36716), .B(n36710), .Z(n36712) );
  IV U36570 ( .A(n36358), .Z(n36716) );
  XOR U36571 ( .A(n36717), .B(n36718), .Z(n36358) );
  AND U36572 ( .A(n599), .B(n36719), .Z(n36718) );
  AND U36573 ( .A(n36671), .B(n36652), .Z(n36710) );
  XNOR U36574 ( .A(n36720), .B(n36721), .Z(n36652) );
  AND U36575 ( .A(n583), .B(n36630), .Z(n36721) );
  XNOR U36576 ( .A(n36628), .B(n36720), .Z(n36630) );
  XNOR U36577 ( .A(n36722), .B(n36723), .Z(n583) );
  AND U36578 ( .A(n36724), .B(n36725), .Z(n36723) );
  XNOR U36579 ( .A(n36722), .B(n36421), .Z(n36725) );
  IV U36580 ( .A(n36425), .Z(n36421) );
  XOR U36581 ( .A(n36726), .B(n36727), .Z(n36425) );
  AND U36582 ( .A(n587), .B(n36728), .Z(n36727) );
  XOR U36583 ( .A(n36729), .B(n36726), .Z(n36728) );
  XNOR U36584 ( .A(n36722), .B(n36635), .Z(n36724) );
  XOR U36585 ( .A(n36730), .B(n36731), .Z(n36635) );
  AND U36586 ( .A(n595), .B(n36682), .Z(n36731) );
  XOR U36587 ( .A(n36680), .B(n36730), .Z(n36682) );
  XOR U36588 ( .A(n36732), .B(n36733), .Z(n36722) );
  AND U36589 ( .A(n36734), .B(n36735), .Z(n36733) );
  XNOR U36590 ( .A(n36732), .B(n36437), .Z(n36735) );
  IV U36591 ( .A(n36440), .Z(n36437) );
  XOR U36592 ( .A(n36736), .B(n36737), .Z(n36440) );
  AND U36593 ( .A(n587), .B(n36738), .Z(n36737) );
  XOR U36594 ( .A(n36739), .B(n36736), .Z(n36738) );
  XOR U36595 ( .A(n36441), .B(n36732), .Z(n36734) );
  XOR U36596 ( .A(n36740), .B(n36741), .Z(n36441) );
  AND U36597 ( .A(n595), .B(n36692), .Z(n36741) );
  XOR U36598 ( .A(n36740), .B(n36690), .Z(n36692) );
  XOR U36599 ( .A(n36742), .B(n36743), .Z(n36732) );
  AND U36600 ( .A(n36744), .B(n36745), .Z(n36743) );
  XNOR U36601 ( .A(n36742), .B(n36465), .Z(n36745) );
  IV U36602 ( .A(n36468), .Z(n36465) );
  XOR U36603 ( .A(n36746), .B(n36747), .Z(n36468) );
  AND U36604 ( .A(n587), .B(n36748), .Z(n36747) );
  XNOR U36605 ( .A(n36749), .B(n36746), .Z(n36748) );
  XOR U36606 ( .A(n36469), .B(n36742), .Z(n36744) );
  XOR U36607 ( .A(n36750), .B(n36751), .Z(n36469) );
  AND U36608 ( .A(n595), .B(n36701), .Z(n36751) );
  XOR U36609 ( .A(n36750), .B(n36699), .Z(n36701) );
  XOR U36610 ( .A(n36752), .B(n36753), .Z(n36742) );
  AND U36611 ( .A(n36754), .B(n36755), .Z(n36753) );
  XNOR U36612 ( .A(n36752), .B(n36514), .Z(n36755) );
  IV U36613 ( .A(n36517), .Z(n36514) );
  XOR U36614 ( .A(n36756), .B(n36757), .Z(n36517) );
  AND U36615 ( .A(n587), .B(n36758), .Z(n36757) );
  XOR U36616 ( .A(n36759), .B(n36756), .Z(n36758) );
  XOR U36617 ( .A(n36518), .B(n36752), .Z(n36754) );
  XOR U36618 ( .A(n36760), .B(n36761), .Z(n36518) );
  AND U36619 ( .A(n595), .B(n36709), .Z(n36761) );
  XOR U36620 ( .A(n36760), .B(n36707), .Z(n36709) );
  XOR U36621 ( .A(n36648), .B(n36762), .Z(n36752) );
  AND U36622 ( .A(n36650), .B(n36763), .Z(n36762) );
  XNOR U36623 ( .A(n36648), .B(n36607), .Z(n36763) );
  IV U36624 ( .A(n36610), .Z(n36607) );
  XOR U36625 ( .A(n36764), .B(n36765), .Z(n36610) );
  AND U36626 ( .A(n587), .B(n36766), .Z(n36765) );
  XNOR U36627 ( .A(n36767), .B(n36764), .Z(n36766) );
  XOR U36628 ( .A(n36611), .B(n36648), .Z(n36650) );
  XOR U36629 ( .A(n36768), .B(n36769), .Z(n36611) );
  AND U36630 ( .A(n595), .B(n36719), .Z(n36769) );
  XOR U36631 ( .A(n36768), .B(n36717), .Z(n36719) );
  AND U36632 ( .A(n36720), .B(n36628), .Z(n36648) );
  XNOR U36633 ( .A(n36770), .B(n36771), .Z(n36628) );
  AND U36634 ( .A(n587), .B(n36772), .Z(n36771) );
  XNOR U36635 ( .A(n36773), .B(n36770), .Z(n36772) );
  XNOR U36636 ( .A(n36774), .B(n36775), .Z(n587) );
  AND U36637 ( .A(n36776), .B(n36777), .Z(n36775) );
  XOR U36638 ( .A(n36729), .B(n36774), .Z(n36777) );
  AND U36639 ( .A(n36778), .B(n36779), .Z(n36729) );
  XNOR U36640 ( .A(n36726), .B(n36774), .Z(n36776) );
  XNOR U36641 ( .A(n36780), .B(n36781), .Z(n36726) );
  AND U36642 ( .A(n591), .B(n36782), .Z(n36781) );
  XNOR U36643 ( .A(n36783), .B(n36784), .Z(n36782) );
  XOR U36644 ( .A(n36785), .B(n36786), .Z(n36774) );
  AND U36645 ( .A(n36787), .B(n36788), .Z(n36786) );
  XNOR U36646 ( .A(n36785), .B(n36778), .Z(n36788) );
  IV U36647 ( .A(n36739), .Z(n36778) );
  XOR U36648 ( .A(n36789), .B(n36790), .Z(n36739) );
  XOR U36649 ( .A(n36791), .B(n36779), .Z(n36790) );
  AND U36650 ( .A(n36749), .B(n36792), .Z(n36779) );
  AND U36651 ( .A(n36793), .B(n36794), .Z(n36791) );
  XOR U36652 ( .A(n36795), .B(n36789), .Z(n36793) );
  XNOR U36653 ( .A(n36736), .B(n36785), .Z(n36787) );
  XNOR U36654 ( .A(n36796), .B(n36797), .Z(n36736) );
  AND U36655 ( .A(n591), .B(n36798), .Z(n36797) );
  XNOR U36656 ( .A(n36799), .B(n36800), .Z(n36798) );
  XOR U36657 ( .A(n36801), .B(n36802), .Z(n36785) );
  AND U36658 ( .A(n36803), .B(n36804), .Z(n36802) );
  XNOR U36659 ( .A(n36801), .B(n36749), .Z(n36804) );
  XOR U36660 ( .A(n36805), .B(n36794), .Z(n36749) );
  XNOR U36661 ( .A(n36806), .B(n36789), .Z(n36794) );
  XOR U36662 ( .A(n36807), .B(n36808), .Z(n36789) );
  AND U36663 ( .A(n36809), .B(n36810), .Z(n36808) );
  XOR U36664 ( .A(n36811), .B(n36807), .Z(n36809) );
  XNOR U36665 ( .A(n36812), .B(n36813), .Z(n36806) );
  AND U36666 ( .A(n36814), .B(n36815), .Z(n36813) );
  XOR U36667 ( .A(n36812), .B(n36816), .Z(n36814) );
  XNOR U36668 ( .A(n36795), .B(n36792), .Z(n36805) );
  AND U36669 ( .A(n36817), .B(n36818), .Z(n36792) );
  XOR U36670 ( .A(n36819), .B(n36820), .Z(n36795) );
  AND U36671 ( .A(n36821), .B(n36822), .Z(n36820) );
  XOR U36672 ( .A(n36819), .B(n36823), .Z(n36821) );
  XNOR U36673 ( .A(n36746), .B(n36801), .Z(n36803) );
  XNOR U36674 ( .A(n36824), .B(n36825), .Z(n36746) );
  AND U36675 ( .A(n591), .B(n36826), .Z(n36825) );
  XNOR U36676 ( .A(n36827), .B(n36828), .Z(n36826) );
  XOR U36677 ( .A(n36829), .B(n36830), .Z(n36801) );
  AND U36678 ( .A(n36831), .B(n36832), .Z(n36830) );
  XNOR U36679 ( .A(n36829), .B(n36817), .Z(n36832) );
  IV U36680 ( .A(n36759), .Z(n36817) );
  XNOR U36681 ( .A(n36833), .B(n36810), .Z(n36759) );
  XNOR U36682 ( .A(n36834), .B(n36816), .Z(n36810) );
  XOR U36683 ( .A(n36835), .B(n36836), .Z(n36816) );
  AND U36684 ( .A(n36837), .B(n36838), .Z(n36836) );
  XOR U36685 ( .A(n36835), .B(n36839), .Z(n36837) );
  XNOR U36686 ( .A(n36815), .B(n36807), .Z(n36834) );
  XOR U36687 ( .A(n36840), .B(n36841), .Z(n36807) );
  AND U36688 ( .A(n36842), .B(n36843), .Z(n36841) );
  XNOR U36689 ( .A(n36844), .B(n36840), .Z(n36842) );
  XNOR U36690 ( .A(n36845), .B(n36812), .Z(n36815) );
  XOR U36691 ( .A(n36846), .B(n36847), .Z(n36812) );
  AND U36692 ( .A(n36848), .B(n36849), .Z(n36847) );
  XOR U36693 ( .A(n36846), .B(n36850), .Z(n36848) );
  XNOR U36694 ( .A(n36851), .B(n36852), .Z(n36845) );
  AND U36695 ( .A(n36853), .B(n36854), .Z(n36852) );
  XNOR U36696 ( .A(n36851), .B(n36855), .Z(n36853) );
  XNOR U36697 ( .A(n36811), .B(n36818), .Z(n36833) );
  AND U36698 ( .A(n36767), .B(n36856), .Z(n36818) );
  XOR U36699 ( .A(n36823), .B(n36822), .Z(n36811) );
  XNOR U36700 ( .A(n36857), .B(n36819), .Z(n36822) );
  XOR U36701 ( .A(n36858), .B(n36859), .Z(n36819) );
  AND U36702 ( .A(n36860), .B(n36861), .Z(n36859) );
  XOR U36703 ( .A(n36858), .B(n36862), .Z(n36860) );
  XNOR U36704 ( .A(n36863), .B(n36864), .Z(n36857) );
  AND U36705 ( .A(n36865), .B(n36866), .Z(n36864) );
  XOR U36706 ( .A(n36863), .B(n36867), .Z(n36865) );
  XOR U36707 ( .A(n36868), .B(n36869), .Z(n36823) );
  AND U36708 ( .A(n36870), .B(n36871), .Z(n36869) );
  XOR U36709 ( .A(n36868), .B(n36872), .Z(n36870) );
  XNOR U36710 ( .A(n36756), .B(n36829), .Z(n36831) );
  XNOR U36711 ( .A(n36873), .B(n36874), .Z(n36756) );
  AND U36712 ( .A(n591), .B(n36875), .Z(n36874) );
  XNOR U36713 ( .A(n36876), .B(n36877), .Z(n36875) );
  XOR U36714 ( .A(n36878), .B(n36879), .Z(n36829) );
  AND U36715 ( .A(n36880), .B(n36881), .Z(n36879) );
  XNOR U36716 ( .A(n36878), .B(n36767), .Z(n36881) );
  XOR U36717 ( .A(n36882), .B(n36843), .Z(n36767) );
  XNOR U36718 ( .A(n36883), .B(n36850), .Z(n36843) );
  XOR U36719 ( .A(n36839), .B(n36838), .Z(n36850) );
  XNOR U36720 ( .A(n36884), .B(n36835), .Z(n36838) );
  XOR U36721 ( .A(n36885), .B(n36886), .Z(n36835) );
  AND U36722 ( .A(n36887), .B(n36888), .Z(n36886) );
  XOR U36723 ( .A(n36885), .B(n36889), .Z(n36887) );
  XNOR U36724 ( .A(n36890), .B(n36891), .Z(n36884) );
  NOR U36725 ( .A(n36892), .B(n36893), .Z(n36891) );
  XNOR U36726 ( .A(n36890), .B(n36894), .Z(n36892) );
  XOR U36727 ( .A(n36895), .B(n36896), .Z(n36839) );
  NOR U36728 ( .A(n36897), .B(n36898), .Z(n36896) );
  XNOR U36729 ( .A(n36895), .B(n36899), .Z(n36897) );
  XNOR U36730 ( .A(n36849), .B(n36840), .Z(n36883) );
  XOR U36731 ( .A(n36900), .B(n36901), .Z(n36840) );
  NOR U36732 ( .A(n36902), .B(n36903), .Z(n36901) );
  XNOR U36733 ( .A(n36900), .B(n36904), .Z(n36902) );
  XOR U36734 ( .A(n36905), .B(n36855), .Z(n36849) );
  XNOR U36735 ( .A(n36906), .B(n36907), .Z(n36855) );
  NOR U36736 ( .A(n36908), .B(n36909), .Z(n36907) );
  XNOR U36737 ( .A(n36906), .B(n36910), .Z(n36908) );
  XNOR U36738 ( .A(n36854), .B(n36846), .Z(n36905) );
  XOR U36739 ( .A(n36911), .B(n36912), .Z(n36846) );
  AND U36740 ( .A(n36913), .B(n36914), .Z(n36912) );
  XOR U36741 ( .A(n36911), .B(n36915), .Z(n36913) );
  XNOR U36742 ( .A(n36916), .B(n36851), .Z(n36854) );
  XOR U36743 ( .A(n36917), .B(n36918), .Z(n36851) );
  AND U36744 ( .A(n36919), .B(n36920), .Z(n36918) );
  XOR U36745 ( .A(n36917), .B(n36921), .Z(n36919) );
  XNOR U36746 ( .A(n36922), .B(n36923), .Z(n36916) );
  NOR U36747 ( .A(n36924), .B(n36925), .Z(n36923) );
  XOR U36748 ( .A(n36922), .B(n36926), .Z(n36924) );
  XOR U36749 ( .A(n36844), .B(n36856), .Z(n36882) );
  NOR U36750 ( .A(n36773), .B(n36927), .Z(n36856) );
  XNOR U36751 ( .A(n36862), .B(n36861), .Z(n36844) );
  XNOR U36752 ( .A(n36928), .B(n36867), .Z(n36861) );
  XOR U36753 ( .A(n36929), .B(n36930), .Z(n36867) );
  NOR U36754 ( .A(n36931), .B(n36932), .Z(n36930) );
  XNOR U36755 ( .A(n36929), .B(n36933), .Z(n36931) );
  XNOR U36756 ( .A(n36866), .B(n36858), .Z(n36928) );
  XOR U36757 ( .A(n36934), .B(n36935), .Z(n36858) );
  AND U36758 ( .A(n36936), .B(n36937), .Z(n36935) );
  XNOR U36759 ( .A(n36934), .B(n36938), .Z(n36936) );
  XNOR U36760 ( .A(n36939), .B(n36863), .Z(n36866) );
  XOR U36761 ( .A(n36940), .B(n36941), .Z(n36863) );
  AND U36762 ( .A(n36942), .B(n36943), .Z(n36941) );
  XOR U36763 ( .A(n36940), .B(n36944), .Z(n36942) );
  XNOR U36764 ( .A(n36945), .B(n36946), .Z(n36939) );
  NOR U36765 ( .A(n36947), .B(n36948), .Z(n36946) );
  XOR U36766 ( .A(n36945), .B(n36949), .Z(n36947) );
  XOR U36767 ( .A(n36872), .B(n36871), .Z(n36862) );
  XNOR U36768 ( .A(n36950), .B(n36868), .Z(n36871) );
  XOR U36769 ( .A(n36951), .B(n36952), .Z(n36868) );
  AND U36770 ( .A(n36953), .B(n36954), .Z(n36952) );
  XOR U36771 ( .A(n36951), .B(n36955), .Z(n36953) );
  XNOR U36772 ( .A(n36956), .B(n36957), .Z(n36950) );
  NOR U36773 ( .A(n36958), .B(n36959), .Z(n36957) );
  XNOR U36774 ( .A(n36956), .B(n36960), .Z(n36958) );
  XOR U36775 ( .A(n36961), .B(n36962), .Z(n36872) );
  NOR U36776 ( .A(n36963), .B(n36964), .Z(n36962) );
  XNOR U36777 ( .A(n36961), .B(n36965), .Z(n36963) );
  XNOR U36778 ( .A(n36764), .B(n36878), .Z(n36880) );
  XNOR U36779 ( .A(n36966), .B(n36967), .Z(n36764) );
  AND U36780 ( .A(n591), .B(n36968), .Z(n36967) );
  XNOR U36781 ( .A(n36969), .B(n36970), .Z(n36968) );
  AND U36782 ( .A(n36770), .B(n36773), .Z(n36878) );
  XOR U36783 ( .A(n36971), .B(n36927), .Z(n36773) );
  XNOR U36784 ( .A(p_input[2048]), .B(p_input[768]), .Z(n36927) );
  XOR U36785 ( .A(n36904), .B(n36903), .Z(n36971) );
  XOR U36786 ( .A(n36972), .B(n36915), .Z(n36903) );
  XOR U36787 ( .A(n36889), .B(n36888), .Z(n36915) );
  XNOR U36788 ( .A(n36973), .B(n36894), .Z(n36888) );
  XOR U36789 ( .A(p_input[2072]), .B(p_input[792]), .Z(n36894) );
  XOR U36790 ( .A(n36885), .B(n36893), .Z(n36973) );
  XOR U36791 ( .A(n36974), .B(n36890), .Z(n36893) );
  XOR U36792 ( .A(p_input[2070]), .B(p_input[790]), .Z(n36890) );
  XNOR U36793 ( .A(p_input[2071]), .B(p_input[791]), .Z(n36974) );
  XNOR U36794 ( .A(n28684), .B(p_input[786]), .Z(n36885) );
  XNOR U36795 ( .A(n36899), .B(n36898), .Z(n36889) );
  XOR U36796 ( .A(n36975), .B(n36895), .Z(n36898) );
  XOR U36797 ( .A(p_input[2067]), .B(p_input[787]), .Z(n36895) );
  XNOR U36798 ( .A(p_input[2068]), .B(p_input[788]), .Z(n36975) );
  XOR U36799 ( .A(p_input[2069]), .B(p_input[789]), .Z(n36899) );
  XNOR U36800 ( .A(n36914), .B(n36900), .Z(n36972) );
  XNOR U36801 ( .A(n28686), .B(p_input[769]), .Z(n36900) );
  XNOR U36802 ( .A(n36976), .B(n36921), .Z(n36914) );
  XNOR U36803 ( .A(n36910), .B(n36909), .Z(n36921) );
  XOR U36804 ( .A(n36977), .B(n36906), .Z(n36909) );
  XNOR U36805 ( .A(n28322), .B(p_input[794]), .Z(n36906) );
  XNOR U36806 ( .A(p_input[2075]), .B(p_input[795]), .Z(n36977) );
  XOR U36807 ( .A(p_input[2076]), .B(p_input[796]), .Z(n36910) );
  XNOR U36808 ( .A(n36920), .B(n36911), .Z(n36976) );
  XNOR U36809 ( .A(n28689), .B(p_input[785]), .Z(n36911) );
  XOR U36810 ( .A(n36978), .B(n36926), .Z(n36920) );
  XNOR U36811 ( .A(p_input[2079]), .B(p_input[799]), .Z(n36926) );
  XOR U36812 ( .A(n36917), .B(n36925), .Z(n36978) );
  XOR U36813 ( .A(n36979), .B(n36922), .Z(n36925) );
  XOR U36814 ( .A(p_input[2077]), .B(p_input[797]), .Z(n36922) );
  XNOR U36815 ( .A(p_input[2078]), .B(p_input[798]), .Z(n36979) );
  XNOR U36816 ( .A(n28326), .B(p_input[793]), .Z(n36917) );
  XNOR U36817 ( .A(n36938), .B(n36937), .Z(n36904) );
  XNOR U36818 ( .A(n36980), .B(n36944), .Z(n36937) );
  XNOR U36819 ( .A(n36933), .B(n36932), .Z(n36944) );
  XOR U36820 ( .A(n36981), .B(n36929), .Z(n36932) );
  XNOR U36821 ( .A(n28694), .B(p_input[779]), .Z(n36929) );
  XNOR U36822 ( .A(p_input[2060]), .B(p_input[780]), .Z(n36981) );
  XOR U36823 ( .A(p_input[2061]), .B(p_input[781]), .Z(n36933) );
  XNOR U36824 ( .A(n36943), .B(n36934), .Z(n36980) );
  XNOR U36825 ( .A(n28330), .B(p_input[770]), .Z(n36934) );
  XOR U36826 ( .A(n36982), .B(n36949), .Z(n36943) );
  XNOR U36827 ( .A(p_input[2064]), .B(p_input[784]), .Z(n36949) );
  XOR U36828 ( .A(n36940), .B(n36948), .Z(n36982) );
  XOR U36829 ( .A(n36983), .B(n36945), .Z(n36948) );
  XOR U36830 ( .A(p_input[2062]), .B(p_input[782]), .Z(n36945) );
  XNOR U36831 ( .A(p_input[2063]), .B(p_input[783]), .Z(n36983) );
  XNOR U36832 ( .A(n28697), .B(p_input[778]), .Z(n36940) );
  XNOR U36833 ( .A(n36955), .B(n36954), .Z(n36938) );
  XNOR U36834 ( .A(n36984), .B(n36960), .Z(n36954) );
  XOR U36835 ( .A(p_input[2057]), .B(p_input[777]), .Z(n36960) );
  XOR U36836 ( .A(n36951), .B(n36959), .Z(n36984) );
  XOR U36837 ( .A(n36985), .B(n36956), .Z(n36959) );
  XOR U36838 ( .A(p_input[2055]), .B(p_input[775]), .Z(n36956) );
  XNOR U36839 ( .A(p_input[2056]), .B(p_input[776]), .Z(n36985) );
  XNOR U36840 ( .A(n28337), .B(p_input[771]), .Z(n36951) );
  XNOR U36841 ( .A(n36965), .B(n36964), .Z(n36955) );
  XOR U36842 ( .A(n36986), .B(n36961), .Z(n36964) );
  XOR U36843 ( .A(p_input[2052]), .B(p_input[772]), .Z(n36961) );
  XNOR U36844 ( .A(p_input[2053]), .B(p_input[773]), .Z(n36986) );
  XOR U36845 ( .A(p_input[2054]), .B(p_input[774]), .Z(n36965) );
  XNOR U36846 ( .A(n36987), .B(n36988), .Z(n36770) );
  AND U36847 ( .A(n591), .B(n36989), .Z(n36988) );
  XNOR U36848 ( .A(n36990), .B(n36991), .Z(n591) );
  AND U36849 ( .A(n36992), .B(n36993), .Z(n36991) );
  XOR U36850 ( .A(n36784), .B(n36990), .Z(n36993) );
  XNOR U36851 ( .A(n36994), .B(n36990), .Z(n36992) );
  XOR U36852 ( .A(n36995), .B(n36996), .Z(n36990) );
  AND U36853 ( .A(n36997), .B(n36998), .Z(n36996) );
  XOR U36854 ( .A(n36799), .B(n36995), .Z(n36998) );
  XOR U36855 ( .A(n36995), .B(n36800), .Z(n36997) );
  XOR U36856 ( .A(n36999), .B(n37000), .Z(n36995) );
  AND U36857 ( .A(n37001), .B(n37002), .Z(n37000) );
  XOR U36858 ( .A(n36827), .B(n36999), .Z(n37002) );
  XOR U36859 ( .A(n36999), .B(n36828), .Z(n37001) );
  XOR U36860 ( .A(n37003), .B(n37004), .Z(n36999) );
  AND U36861 ( .A(n37005), .B(n37006), .Z(n37004) );
  XOR U36862 ( .A(n36876), .B(n37003), .Z(n37006) );
  XOR U36863 ( .A(n37003), .B(n36877), .Z(n37005) );
  XOR U36864 ( .A(n37007), .B(n37008), .Z(n37003) );
  AND U36865 ( .A(n37009), .B(n37010), .Z(n37008) );
  XOR U36866 ( .A(n37007), .B(n36969), .Z(n37010) );
  XNOR U36867 ( .A(n37011), .B(n37012), .Z(n36720) );
  AND U36868 ( .A(n595), .B(n37013), .Z(n37012) );
  XNOR U36869 ( .A(n37014), .B(n37015), .Z(n595) );
  AND U36870 ( .A(n37016), .B(n37017), .Z(n37015) );
  XOR U36871 ( .A(n37014), .B(n36730), .Z(n37017) );
  XNOR U36872 ( .A(n37014), .B(n36680), .Z(n37016) );
  XOR U36873 ( .A(n37018), .B(n37019), .Z(n37014) );
  AND U36874 ( .A(n37020), .B(n37021), .Z(n37019) );
  XNOR U36875 ( .A(n36740), .B(n37018), .Z(n37021) );
  XOR U36876 ( .A(n37018), .B(n36690), .Z(n37020) );
  XOR U36877 ( .A(n37022), .B(n37023), .Z(n37018) );
  AND U36878 ( .A(n37024), .B(n37025), .Z(n37023) );
  XNOR U36879 ( .A(n36750), .B(n37022), .Z(n37025) );
  XOR U36880 ( .A(n37022), .B(n36699), .Z(n37024) );
  XOR U36881 ( .A(n37026), .B(n37027), .Z(n37022) );
  AND U36882 ( .A(n37028), .B(n37029), .Z(n37027) );
  XOR U36883 ( .A(n37026), .B(n36707), .Z(n37028) );
  XOR U36884 ( .A(n37030), .B(n37031), .Z(n36671) );
  AND U36885 ( .A(n599), .B(n37013), .Z(n37031) );
  XNOR U36886 ( .A(n37011), .B(n37030), .Z(n37013) );
  XNOR U36887 ( .A(n37032), .B(n37033), .Z(n599) );
  AND U36888 ( .A(n37034), .B(n37035), .Z(n37033) );
  XNOR U36889 ( .A(n37036), .B(n37032), .Z(n37035) );
  IV U36890 ( .A(n36730), .Z(n37036) );
  XOR U36891 ( .A(n36994), .B(n37037), .Z(n36730) );
  AND U36892 ( .A(n602), .B(n37038), .Z(n37037) );
  XOR U36893 ( .A(n36783), .B(n36780), .Z(n37038) );
  IV U36894 ( .A(n36994), .Z(n36783) );
  XNOR U36895 ( .A(n36680), .B(n37032), .Z(n37034) );
  XOR U36896 ( .A(n37039), .B(n37040), .Z(n36680) );
  AND U36897 ( .A(n618), .B(n37041), .Z(n37040) );
  XOR U36898 ( .A(n37042), .B(n37043), .Z(n37032) );
  AND U36899 ( .A(n37044), .B(n37045), .Z(n37043) );
  XNOR U36900 ( .A(n37042), .B(n36740), .Z(n37045) );
  XOR U36901 ( .A(n36800), .B(n37046), .Z(n36740) );
  AND U36902 ( .A(n602), .B(n37047), .Z(n37046) );
  XOR U36903 ( .A(n36796), .B(n36800), .Z(n37047) );
  XNOR U36904 ( .A(n37048), .B(n37042), .Z(n37044) );
  IV U36905 ( .A(n36690), .Z(n37048) );
  XOR U36906 ( .A(n37049), .B(n37050), .Z(n36690) );
  AND U36907 ( .A(n618), .B(n37051), .Z(n37050) );
  XOR U36908 ( .A(n37052), .B(n37053), .Z(n37042) );
  AND U36909 ( .A(n37054), .B(n37055), .Z(n37053) );
  XNOR U36910 ( .A(n37052), .B(n36750), .Z(n37055) );
  XOR U36911 ( .A(n36828), .B(n37056), .Z(n36750) );
  AND U36912 ( .A(n602), .B(n37057), .Z(n37056) );
  XOR U36913 ( .A(n36824), .B(n36828), .Z(n37057) );
  XOR U36914 ( .A(n36699), .B(n37052), .Z(n37054) );
  XOR U36915 ( .A(n37058), .B(n37059), .Z(n36699) );
  AND U36916 ( .A(n618), .B(n37060), .Z(n37059) );
  XOR U36917 ( .A(n37026), .B(n37061), .Z(n37052) );
  AND U36918 ( .A(n37062), .B(n37029), .Z(n37061) );
  XNOR U36919 ( .A(n36760), .B(n37026), .Z(n37029) );
  XOR U36920 ( .A(n36877), .B(n37063), .Z(n36760) );
  AND U36921 ( .A(n602), .B(n37064), .Z(n37063) );
  XOR U36922 ( .A(n36873), .B(n36877), .Z(n37064) );
  XNOR U36923 ( .A(n37065), .B(n37026), .Z(n37062) );
  IV U36924 ( .A(n36707), .Z(n37065) );
  XOR U36925 ( .A(n37066), .B(n37067), .Z(n36707) );
  AND U36926 ( .A(n618), .B(n37068), .Z(n37067) );
  XOR U36927 ( .A(n37069), .B(n37070), .Z(n37026) );
  AND U36928 ( .A(n37071), .B(n37072), .Z(n37070) );
  XNOR U36929 ( .A(n37069), .B(n36768), .Z(n37072) );
  XOR U36930 ( .A(n36970), .B(n37073), .Z(n36768) );
  AND U36931 ( .A(n602), .B(n37074), .Z(n37073) );
  XOR U36932 ( .A(n36966), .B(n36970), .Z(n37074) );
  XNOR U36933 ( .A(n37075), .B(n37069), .Z(n37071) );
  IV U36934 ( .A(n36717), .Z(n37075) );
  XOR U36935 ( .A(n37076), .B(n37077), .Z(n36717) );
  AND U36936 ( .A(n618), .B(n37078), .Z(n37077) );
  AND U36937 ( .A(n37030), .B(n37011), .Z(n37069) );
  XNOR U36938 ( .A(n37079), .B(n37080), .Z(n37011) );
  AND U36939 ( .A(n602), .B(n36989), .Z(n37080) );
  XNOR U36940 ( .A(n36987), .B(n37079), .Z(n36989) );
  XNOR U36941 ( .A(n37081), .B(n37082), .Z(n602) );
  AND U36942 ( .A(n37083), .B(n37084), .Z(n37082) );
  XNOR U36943 ( .A(n37081), .B(n36780), .Z(n37084) );
  IV U36944 ( .A(n36784), .Z(n36780) );
  XOR U36945 ( .A(n37085), .B(n37086), .Z(n36784) );
  AND U36946 ( .A(n606), .B(n37087), .Z(n37086) );
  XOR U36947 ( .A(n37088), .B(n37085), .Z(n37087) );
  XNOR U36948 ( .A(n37081), .B(n36994), .Z(n37083) );
  XOR U36949 ( .A(n37089), .B(n37090), .Z(n36994) );
  AND U36950 ( .A(n614), .B(n37041), .Z(n37090) );
  XOR U36951 ( .A(n37039), .B(n37089), .Z(n37041) );
  XOR U36952 ( .A(n37091), .B(n37092), .Z(n37081) );
  AND U36953 ( .A(n37093), .B(n37094), .Z(n37092) );
  XNOR U36954 ( .A(n37091), .B(n36796), .Z(n37094) );
  IV U36955 ( .A(n36799), .Z(n36796) );
  XOR U36956 ( .A(n37095), .B(n37096), .Z(n36799) );
  AND U36957 ( .A(n606), .B(n37097), .Z(n37096) );
  XOR U36958 ( .A(n37098), .B(n37095), .Z(n37097) );
  XOR U36959 ( .A(n36800), .B(n37091), .Z(n37093) );
  XOR U36960 ( .A(n37099), .B(n37100), .Z(n36800) );
  AND U36961 ( .A(n614), .B(n37051), .Z(n37100) );
  XOR U36962 ( .A(n37099), .B(n37049), .Z(n37051) );
  XOR U36963 ( .A(n37101), .B(n37102), .Z(n37091) );
  AND U36964 ( .A(n37103), .B(n37104), .Z(n37102) );
  XNOR U36965 ( .A(n37101), .B(n36824), .Z(n37104) );
  IV U36966 ( .A(n36827), .Z(n36824) );
  XOR U36967 ( .A(n37105), .B(n37106), .Z(n36827) );
  AND U36968 ( .A(n606), .B(n37107), .Z(n37106) );
  XNOR U36969 ( .A(n37108), .B(n37105), .Z(n37107) );
  XOR U36970 ( .A(n36828), .B(n37101), .Z(n37103) );
  XOR U36971 ( .A(n37109), .B(n37110), .Z(n36828) );
  AND U36972 ( .A(n614), .B(n37060), .Z(n37110) );
  XOR U36973 ( .A(n37109), .B(n37058), .Z(n37060) );
  XOR U36974 ( .A(n37111), .B(n37112), .Z(n37101) );
  AND U36975 ( .A(n37113), .B(n37114), .Z(n37112) );
  XNOR U36976 ( .A(n37111), .B(n36873), .Z(n37114) );
  IV U36977 ( .A(n36876), .Z(n36873) );
  XOR U36978 ( .A(n37115), .B(n37116), .Z(n36876) );
  AND U36979 ( .A(n606), .B(n37117), .Z(n37116) );
  XOR U36980 ( .A(n37118), .B(n37115), .Z(n37117) );
  XOR U36981 ( .A(n36877), .B(n37111), .Z(n37113) );
  XOR U36982 ( .A(n37119), .B(n37120), .Z(n36877) );
  AND U36983 ( .A(n614), .B(n37068), .Z(n37120) );
  XOR U36984 ( .A(n37119), .B(n37066), .Z(n37068) );
  XOR U36985 ( .A(n37007), .B(n37121), .Z(n37111) );
  AND U36986 ( .A(n37009), .B(n37122), .Z(n37121) );
  XNOR U36987 ( .A(n37007), .B(n36966), .Z(n37122) );
  IV U36988 ( .A(n36969), .Z(n36966) );
  XOR U36989 ( .A(n37123), .B(n37124), .Z(n36969) );
  AND U36990 ( .A(n606), .B(n37125), .Z(n37124) );
  XNOR U36991 ( .A(n37126), .B(n37123), .Z(n37125) );
  XOR U36992 ( .A(n36970), .B(n37007), .Z(n37009) );
  XOR U36993 ( .A(n37127), .B(n37128), .Z(n36970) );
  AND U36994 ( .A(n614), .B(n37078), .Z(n37128) );
  XOR U36995 ( .A(n37127), .B(n37076), .Z(n37078) );
  AND U36996 ( .A(n37079), .B(n36987), .Z(n37007) );
  XNOR U36997 ( .A(n37129), .B(n37130), .Z(n36987) );
  AND U36998 ( .A(n606), .B(n37131), .Z(n37130) );
  XNOR U36999 ( .A(n37132), .B(n37129), .Z(n37131) );
  XNOR U37000 ( .A(n37133), .B(n37134), .Z(n606) );
  AND U37001 ( .A(n37135), .B(n37136), .Z(n37134) );
  XOR U37002 ( .A(n37088), .B(n37133), .Z(n37136) );
  AND U37003 ( .A(n37137), .B(n37138), .Z(n37088) );
  XNOR U37004 ( .A(n37085), .B(n37133), .Z(n37135) );
  XNOR U37005 ( .A(n37139), .B(n37140), .Z(n37085) );
  AND U37006 ( .A(n610), .B(n37141), .Z(n37140) );
  XNOR U37007 ( .A(n37142), .B(n37143), .Z(n37141) );
  XOR U37008 ( .A(n37144), .B(n37145), .Z(n37133) );
  AND U37009 ( .A(n37146), .B(n37147), .Z(n37145) );
  XNOR U37010 ( .A(n37144), .B(n37137), .Z(n37147) );
  IV U37011 ( .A(n37098), .Z(n37137) );
  XOR U37012 ( .A(n37148), .B(n37149), .Z(n37098) );
  XOR U37013 ( .A(n37150), .B(n37138), .Z(n37149) );
  AND U37014 ( .A(n37108), .B(n37151), .Z(n37138) );
  AND U37015 ( .A(n37152), .B(n37153), .Z(n37150) );
  XOR U37016 ( .A(n37154), .B(n37148), .Z(n37152) );
  XNOR U37017 ( .A(n37095), .B(n37144), .Z(n37146) );
  XNOR U37018 ( .A(n37155), .B(n37156), .Z(n37095) );
  AND U37019 ( .A(n610), .B(n37157), .Z(n37156) );
  XNOR U37020 ( .A(n37158), .B(n37159), .Z(n37157) );
  XOR U37021 ( .A(n37160), .B(n37161), .Z(n37144) );
  AND U37022 ( .A(n37162), .B(n37163), .Z(n37161) );
  XNOR U37023 ( .A(n37160), .B(n37108), .Z(n37163) );
  XOR U37024 ( .A(n37164), .B(n37153), .Z(n37108) );
  XNOR U37025 ( .A(n37165), .B(n37148), .Z(n37153) );
  XOR U37026 ( .A(n37166), .B(n37167), .Z(n37148) );
  AND U37027 ( .A(n37168), .B(n37169), .Z(n37167) );
  XOR U37028 ( .A(n37170), .B(n37166), .Z(n37168) );
  XNOR U37029 ( .A(n37171), .B(n37172), .Z(n37165) );
  AND U37030 ( .A(n37173), .B(n37174), .Z(n37172) );
  XOR U37031 ( .A(n37171), .B(n37175), .Z(n37173) );
  XNOR U37032 ( .A(n37154), .B(n37151), .Z(n37164) );
  AND U37033 ( .A(n37176), .B(n37177), .Z(n37151) );
  XOR U37034 ( .A(n37178), .B(n37179), .Z(n37154) );
  AND U37035 ( .A(n37180), .B(n37181), .Z(n37179) );
  XOR U37036 ( .A(n37178), .B(n37182), .Z(n37180) );
  XNOR U37037 ( .A(n37105), .B(n37160), .Z(n37162) );
  XNOR U37038 ( .A(n37183), .B(n37184), .Z(n37105) );
  AND U37039 ( .A(n610), .B(n37185), .Z(n37184) );
  XNOR U37040 ( .A(n37186), .B(n37187), .Z(n37185) );
  XOR U37041 ( .A(n37188), .B(n37189), .Z(n37160) );
  AND U37042 ( .A(n37190), .B(n37191), .Z(n37189) );
  XNOR U37043 ( .A(n37188), .B(n37176), .Z(n37191) );
  IV U37044 ( .A(n37118), .Z(n37176) );
  XNOR U37045 ( .A(n37192), .B(n37169), .Z(n37118) );
  XNOR U37046 ( .A(n37193), .B(n37175), .Z(n37169) );
  XOR U37047 ( .A(n37194), .B(n37195), .Z(n37175) );
  AND U37048 ( .A(n37196), .B(n37197), .Z(n37195) );
  XOR U37049 ( .A(n37194), .B(n37198), .Z(n37196) );
  XNOR U37050 ( .A(n37174), .B(n37166), .Z(n37193) );
  XOR U37051 ( .A(n37199), .B(n37200), .Z(n37166) );
  AND U37052 ( .A(n37201), .B(n37202), .Z(n37200) );
  XNOR U37053 ( .A(n37203), .B(n37199), .Z(n37201) );
  XNOR U37054 ( .A(n37204), .B(n37171), .Z(n37174) );
  XOR U37055 ( .A(n37205), .B(n37206), .Z(n37171) );
  AND U37056 ( .A(n37207), .B(n37208), .Z(n37206) );
  XOR U37057 ( .A(n37205), .B(n37209), .Z(n37207) );
  XNOR U37058 ( .A(n37210), .B(n37211), .Z(n37204) );
  AND U37059 ( .A(n37212), .B(n37213), .Z(n37211) );
  XNOR U37060 ( .A(n37210), .B(n37214), .Z(n37212) );
  XNOR U37061 ( .A(n37170), .B(n37177), .Z(n37192) );
  AND U37062 ( .A(n37126), .B(n37215), .Z(n37177) );
  XOR U37063 ( .A(n37182), .B(n37181), .Z(n37170) );
  XNOR U37064 ( .A(n37216), .B(n37178), .Z(n37181) );
  XOR U37065 ( .A(n37217), .B(n37218), .Z(n37178) );
  AND U37066 ( .A(n37219), .B(n37220), .Z(n37218) );
  XOR U37067 ( .A(n37217), .B(n37221), .Z(n37219) );
  XNOR U37068 ( .A(n37222), .B(n37223), .Z(n37216) );
  AND U37069 ( .A(n37224), .B(n37225), .Z(n37223) );
  XOR U37070 ( .A(n37222), .B(n37226), .Z(n37224) );
  XOR U37071 ( .A(n37227), .B(n37228), .Z(n37182) );
  AND U37072 ( .A(n37229), .B(n37230), .Z(n37228) );
  XOR U37073 ( .A(n37227), .B(n37231), .Z(n37229) );
  XNOR U37074 ( .A(n37115), .B(n37188), .Z(n37190) );
  XNOR U37075 ( .A(n37232), .B(n37233), .Z(n37115) );
  AND U37076 ( .A(n610), .B(n37234), .Z(n37233) );
  XNOR U37077 ( .A(n37235), .B(n37236), .Z(n37234) );
  XOR U37078 ( .A(n37237), .B(n37238), .Z(n37188) );
  AND U37079 ( .A(n37239), .B(n37240), .Z(n37238) );
  XNOR U37080 ( .A(n37237), .B(n37126), .Z(n37240) );
  XOR U37081 ( .A(n37241), .B(n37202), .Z(n37126) );
  XNOR U37082 ( .A(n37242), .B(n37209), .Z(n37202) );
  XOR U37083 ( .A(n37198), .B(n37197), .Z(n37209) );
  XNOR U37084 ( .A(n37243), .B(n37194), .Z(n37197) );
  XOR U37085 ( .A(n37244), .B(n37245), .Z(n37194) );
  AND U37086 ( .A(n37246), .B(n37247), .Z(n37245) );
  XOR U37087 ( .A(n37244), .B(n37248), .Z(n37246) );
  XNOR U37088 ( .A(n37249), .B(n37250), .Z(n37243) );
  NOR U37089 ( .A(n37251), .B(n37252), .Z(n37250) );
  XNOR U37090 ( .A(n37249), .B(n37253), .Z(n37251) );
  XOR U37091 ( .A(n37254), .B(n37255), .Z(n37198) );
  NOR U37092 ( .A(n37256), .B(n37257), .Z(n37255) );
  XNOR U37093 ( .A(n37254), .B(n37258), .Z(n37256) );
  XNOR U37094 ( .A(n37208), .B(n37199), .Z(n37242) );
  XOR U37095 ( .A(n37259), .B(n37260), .Z(n37199) );
  NOR U37096 ( .A(n37261), .B(n37262), .Z(n37260) );
  XNOR U37097 ( .A(n37259), .B(n37263), .Z(n37261) );
  XOR U37098 ( .A(n37264), .B(n37214), .Z(n37208) );
  XNOR U37099 ( .A(n37265), .B(n37266), .Z(n37214) );
  NOR U37100 ( .A(n37267), .B(n37268), .Z(n37266) );
  XNOR U37101 ( .A(n37265), .B(n37269), .Z(n37267) );
  XNOR U37102 ( .A(n37213), .B(n37205), .Z(n37264) );
  XOR U37103 ( .A(n37270), .B(n37271), .Z(n37205) );
  AND U37104 ( .A(n37272), .B(n37273), .Z(n37271) );
  XOR U37105 ( .A(n37270), .B(n37274), .Z(n37272) );
  XNOR U37106 ( .A(n37275), .B(n37210), .Z(n37213) );
  XOR U37107 ( .A(n37276), .B(n37277), .Z(n37210) );
  AND U37108 ( .A(n37278), .B(n37279), .Z(n37277) );
  XOR U37109 ( .A(n37276), .B(n37280), .Z(n37278) );
  XNOR U37110 ( .A(n37281), .B(n37282), .Z(n37275) );
  NOR U37111 ( .A(n37283), .B(n37284), .Z(n37282) );
  XOR U37112 ( .A(n37281), .B(n37285), .Z(n37283) );
  XOR U37113 ( .A(n37203), .B(n37215), .Z(n37241) );
  NOR U37114 ( .A(n37132), .B(n37286), .Z(n37215) );
  XNOR U37115 ( .A(n37221), .B(n37220), .Z(n37203) );
  XNOR U37116 ( .A(n37287), .B(n37226), .Z(n37220) );
  XOR U37117 ( .A(n37288), .B(n37289), .Z(n37226) );
  NOR U37118 ( .A(n37290), .B(n37291), .Z(n37289) );
  XNOR U37119 ( .A(n37288), .B(n37292), .Z(n37290) );
  XNOR U37120 ( .A(n37225), .B(n37217), .Z(n37287) );
  XOR U37121 ( .A(n37293), .B(n37294), .Z(n37217) );
  AND U37122 ( .A(n37295), .B(n37296), .Z(n37294) );
  XNOR U37123 ( .A(n37293), .B(n37297), .Z(n37295) );
  XNOR U37124 ( .A(n37298), .B(n37222), .Z(n37225) );
  XOR U37125 ( .A(n37299), .B(n37300), .Z(n37222) );
  AND U37126 ( .A(n37301), .B(n37302), .Z(n37300) );
  XOR U37127 ( .A(n37299), .B(n37303), .Z(n37301) );
  XNOR U37128 ( .A(n37304), .B(n37305), .Z(n37298) );
  NOR U37129 ( .A(n37306), .B(n37307), .Z(n37305) );
  XOR U37130 ( .A(n37304), .B(n37308), .Z(n37306) );
  XOR U37131 ( .A(n37231), .B(n37230), .Z(n37221) );
  XNOR U37132 ( .A(n37309), .B(n37227), .Z(n37230) );
  XOR U37133 ( .A(n37310), .B(n37311), .Z(n37227) );
  AND U37134 ( .A(n37312), .B(n37313), .Z(n37311) );
  XOR U37135 ( .A(n37310), .B(n37314), .Z(n37312) );
  XNOR U37136 ( .A(n37315), .B(n37316), .Z(n37309) );
  NOR U37137 ( .A(n37317), .B(n37318), .Z(n37316) );
  XNOR U37138 ( .A(n37315), .B(n37319), .Z(n37317) );
  XOR U37139 ( .A(n37320), .B(n37321), .Z(n37231) );
  NOR U37140 ( .A(n37322), .B(n37323), .Z(n37321) );
  XNOR U37141 ( .A(n37320), .B(n37324), .Z(n37322) );
  XNOR U37142 ( .A(n37123), .B(n37237), .Z(n37239) );
  XNOR U37143 ( .A(n37325), .B(n37326), .Z(n37123) );
  AND U37144 ( .A(n610), .B(n37327), .Z(n37326) );
  XNOR U37145 ( .A(n37328), .B(n37329), .Z(n37327) );
  AND U37146 ( .A(n37129), .B(n37132), .Z(n37237) );
  XOR U37147 ( .A(n37330), .B(n37286), .Z(n37132) );
  XNOR U37148 ( .A(p_input[2048]), .B(p_input[800]), .Z(n37286) );
  XOR U37149 ( .A(n37263), .B(n37262), .Z(n37330) );
  XOR U37150 ( .A(n37331), .B(n37274), .Z(n37262) );
  XOR U37151 ( .A(n37248), .B(n37247), .Z(n37274) );
  XNOR U37152 ( .A(n37332), .B(n37253), .Z(n37247) );
  XOR U37153 ( .A(p_input[2072]), .B(p_input[824]), .Z(n37253) );
  XOR U37154 ( .A(n37244), .B(n37252), .Z(n37332) );
  XOR U37155 ( .A(n37333), .B(n37249), .Z(n37252) );
  XOR U37156 ( .A(p_input[2070]), .B(p_input[822]), .Z(n37249) );
  XNOR U37157 ( .A(p_input[2071]), .B(p_input[823]), .Z(n37333) );
  XNOR U37158 ( .A(n28684), .B(p_input[818]), .Z(n37244) );
  XNOR U37159 ( .A(n37258), .B(n37257), .Z(n37248) );
  XOR U37160 ( .A(n37334), .B(n37254), .Z(n37257) );
  XOR U37161 ( .A(p_input[2067]), .B(p_input[819]), .Z(n37254) );
  XNOR U37162 ( .A(p_input[2068]), .B(p_input[820]), .Z(n37334) );
  XOR U37163 ( .A(p_input[2069]), .B(p_input[821]), .Z(n37258) );
  XNOR U37164 ( .A(n37273), .B(n37259), .Z(n37331) );
  XNOR U37165 ( .A(n28686), .B(p_input[801]), .Z(n37259) );
  XNOR U37166 ( .A(n37335), .B(n37280), .Z(n37273) );
  XNOR U37167 ( .A(n37269), .B(n37268), .Z(n37280) );
  XOR U37168 ( .A(n37336), .B(n37265), .Z(n37268) );
  XNOR U37169 ( .A(n28322), .B(p_input[826]), .Z(n37265) );
  XNOR U37170 ( .A(p_input[2075]), .B(p_input[827]), .Z(n37336) );
  XOR U37171 ( .A(p_input[2076]), .B(p_input[828]), .Z(n37269) );
  XNOR U37172 ( .A(n37279), .B(n37270), .Z(n37335) );
  XNOR U37173 ( .A(n28689), .B(p_input[817]), .Z(n37270) );
  XOR U37174 ( .A(n37337), .B(n37285), .Z(n37279) );
  XNOR U37175 ( .A(p_input[2079]), .B(p_input[831]), .Z(n37285) );
  XOR U37176 ( .A(n37276), .B(n37284), .Z(n37337) );
  XOR U37177 ( .A(n37338), .B(n37281), .Z(n37284) );
  XOR U37178 ( .A(p_input[2077]), .B(p_input[829]), .Z(n37281) );
  XNOR U37179 ( .A(p_input[2078]), .B(p_input[830]), .Z(n37338) );
  XNOR U37180 ( .A(n28326), .B(p_input[825]), .Z(n37276) );
  XNOR U37181 ( .A(n37297), .B(n37296), .Z(n37263) );
  XNOR U37182 ( .A(n37339), .B(n37303), .Z(n37296) );
  XNOR U37183 ( .A(n37292), .B(n37291), .Z(n37303) );
  XOR U37184 ( .A(n37340), .B(n37288), .Z(n37291) );
  XNOR U37185 ( .A(n28694), .B(p_input[811]), .Z(n37288) );
  XNOR U37186 ( .A(p_input[2060]), .B(p_input[812]), .Z(n37340) );
  XOR U37187 ( .A(p_input[2061]), .B(p_input[813]), .Z(n37292) );
  XNOR U37188 ( .A(n37302), .B(n37293), .Z(n37339) );
  XNOR U37189 ( .A(n28330), .B(p_input[802]), .Z(n37293) );
  XOR U37190 ( .A(n37341), .B(n37308), .Z(n37302) );
  XNOR U37191 ( .A(p_input[2064]), .B(p_input[816]), .Z(n37308) );
  XOR U37192 ( .A(n37299), .B(n37307), .Z(n37341) );
  XOR U37193 ( .A(n37342), .B(n37304), .Z(n37307) );
  XOR U37194 ( .A(p_input[2062]), .B(p_input[814]), .Z(n37304) );
  XNOR U37195 ( .A(p_input[2063]), .B(p_input[815]), .Z(n37342) );
  XNOR U37196 ( .A(n28697), .B(p_input[810]), .Z(n37299) );
  XNOR U37197 ( .A(n37314), .B(n37313), .Z(n37297) );
  XNOR U37198 ( .A(n37343), .B(n37319), .Z(n37313) );
  XOR U37199 ( .A(p_input[2057]), .B(p_input[809]), .Z(n37319) );
  XOR U37200 ( .A(n37310), .B(n37318), .Z(n37343) );
  XOR U37201 ( .A(n37344), .B(n37315), .Z(n37318) );
  XOR U37202 ( .A(p_input[2055]), .B(p_input[807]), .Z(n37315) );
  XNOR U37203 ( .A(p_input[2056]), .B(p_input[808]), .Z(n37344) );
  XNOR U37204 ( .A(n28337), .B(p_input[803]), .Z(n37310) );
  XNOR U37205 ( .A(n37324), .B(n37323), .Z(n37314) );
  XOR U37206 ( .A(n37345), .B(n37320), .Z(n37323) );
  XOR U37207 ( .A(p_input[2052]), .B(p_input[804]), .Z(n37320) );
  XNOR U37208 ( .A(p_input[2053]), .B(p_input[805]), .Z(n37345) );
  XOR U37209 ( .A(p_input[2054]), .B(p_input[806]), .Z(n37324) );
  XNOR U37210 ( .A(n37346), .B(n37347), .Z(n37129) );
  AND U37211 ( .A(n610), .B(n37348), .Z(n37347) );
  XNOR U37212 ( .A(n37349), .B(n37350), .Z(n610) );
  AND U37213 ( .A(n37351), .B(n37352), .Z(n37350) );
  XOR U37214 ( .A(n37143), .B(n37349), .Z(n37352) );
  XNOR U37215 ( .A(n37353), .B(n37349), .Z(n37351) );
  XOR U37216 ( .A(n37354), .B(n37355), .Z(n37349) );
  AND U37217 ( .A(n37356), .B(n37357), .Z(n37355) );
  XOR U37218 ( .A(n37158), .B(n37354), .Z(n37357) );
  XOR U37219 ( .A(n37354), .B(n37159), .Z(n37356) );
  XOR U37220 ( .A(n37358), .B(n37359), .Z(n37354) );
  AND U37221 ( .A(n37360), .B(n37361), .Z(n37359) );
  XOR U37222 ( .A(n37186), .B(n37358), .Z(n37361) );
  XOR U37223 ( .A(n37358), .B(n37187), .Z(n37360) );
  XOR U37224 ( .A(n37362), .B(n37363), .Z(n37358) );
  AND U37225 ( .A(n37364), .B(n37365), .Z(n37363) );
  XOR U37226 ( .A(n37235), .B(n37362), .Z(n37365) );
  XOR U37227 ( .A(n37362), .B(n37236), .Z(n37364) );
  XOR U37228 ( .A(n37366), .B(n37367), .Z(n37362) );
  AND U37229 ( .A(n37368), .B(n37369), .Z(n37367) );
  XOR U37230 ( .A(n37366), .B(n37328), .Z(n37369) );
  XNOR U37231 ( .A(n37370), .B(n37371), .Z(n37079) );
  AND U37232 ( .A(n614), .B(n37372), .Z(n37371) );
  XNOR U37233 ( .A(n37373), .B(n37374), .Z(n614) );
  AND U37234 ( .A(n37375), .B(n37376), .Z(n37374) );
  XOR U37235 ( .A(n37373), .B(n37089), .Z(n37376) );
  XNOR U37236 ( .A(n37373), .B(n37039), .Z(n37375) );
  XOR U37237 ( .A(n37377), .B(n37378), .Z(n37373) );
  AND U37238 ( .A(n37379), .B(n37380), .Z(n37378) );
  XNOR U37239 ( .A(n37099), .B(n37377), .Z(n37380) );
  XOR U37240 ( .A(n37377), .B(n37049), .Z(n37379) );
  XOR U37241 ( .A(n37381), .B(n37382), .Z(n37377) );
  AND U37242 ( .A(n37383), .B(n37384), .Z(n37382) );
  XNOR U37243 ( .A(n37109), .B(n37381), .Z(n37384) );
  XOR U37244 ( .A(n37381), .B(n37058), .Z(n37383) );
  XOR U37245 ( .A(n37385), .B(n37386), .Z(n37381) );
  AND U37246 ( .A(n37387), .B(n37388), .Z(n37386) );
  XOR U37247 ( .A(n37385), .B(n37066), .Z(n37387) );
  XOR U37248 ( .A(n37389), .B(n37390), .Z(n37030) );
  AND U37249 ( .A(n618), .B(n37372), .Z(n37390) );
  XNOR U37250 ( .A(n37370), .B(n37389), .Z(n37372) );
  XNOR U37251 ( .A(n37391), .B(n37392), .Z(n618) );
  AND U37252 ( .A(n37393), .B(n37394), .Z(n37392) );
  XNOR U37253 ( .A(n37395), .B(n37391), .Z(n37394) );
  IV U37254 ( .A(n37089), .Z(n37395) );
  XOR U37255 ( .A(n37353), .B(n37396), .Z(n37089) );
  AND U37256 ( .A(n621), .B(n37397), .Z(n37396) );
  XOR U37257 ( .A(n37142), .B(n37139), .Z(n37397) );
  IV U37258 ( .A(n37353), .Z(n37142) );
  XNOR U37259 ( .A(n37039), .B(n37391), .Z(n37393) );
  XOR U37260 ( .A(n37398), .B(n37399), .Z(n37039) );
  AND U37261 ( .A(n637), .B(n37400), .Z(n37399) );
  XOR U37262 ( .A(n37401), .B(n37402), .Z(n37391) );
  AND U37263 ( .A(n37403), .B(n37404), .Z(n37402) );
  XNOR U37264 ( .A(n37401), .B(n37099), .Z(n37404) );
  XOR U37265 ( .A(n37159), .B(n37405), .Z(n37099) );
  AND U37266 ( .A(n621), .B(n37406), .Z(n37405) );
  XOR U37267 ( .A(n37155), .B(n37159), .Z(n37406) );
  XNOR U37268 ( .A(n37407), .B(n37401), .Z(n37403) );
  IV U37269 ( .A(n37049), .Z(n37407) );
  XOR U37270 ( .A(n37408), .B(n37409), .Z(n37049) );
  AND U37271 ( .A(n637), .B(n37410), .Z(n37409) );
  XOR U37272 ( .A(n37411), .B(n37412), .Z(n37401) );
  AND U37273 ( .A(n37413), .B(n37414), .Z(n37412) );
  XNOR U37274 ( .A(n37411), .B(n37109), .Z(n37414) );
  XOR U37275 ( .A(n37187), .B(n37415), .Z(n37109) );
  AND U37276 ( .A(n621), .B(n37416), .Z(n37415) );
  XOR U37277 ( .A(n37183), .B(n37187), .Z(n37416) );
  XOR U37278 ( .A(n37058), .B(n37411), .Z(n37413) );
  XOR U37279 ( .A(n37417), .B(n37418), .Z(n37058) );
  AND U37280 ( .A(n637), .B(n37419), .Z(n37418) );
  XOR U37281 ( .A(n37385), .B(n37420), .Z(n37411) );
  AND U37282 ( .A(n37421), .B(n37388), .Z(n37420) );
  XNOR U37283 ( .A(n37119), .B(n37385), .Z(n37388) );
  XOR U37284 ( .A(n37236), .B(n37422), .Z(n37119) );
  AND U37285 ( .A(n621), .B(n37423), .Z(n37422) );
  XOR U37286 ( .A(n37232), .B(n37236), .Z(n37423) );
  XNOR U37287 ( .A(n37424), .B(n37385), .Z(n37421) );
  IV U37288 ( .A(n37066), .Z(n37424) );
  XOR U37289 ( .A(n37425), .B(n37426), .Z(n37066) );
  AND U37290 ( .A(n637), .B(n37427), .Z(n37426) );
  XOR U37291 ( .A(n37428), .B(n37429), .Z(n37385) );
  AND U37292 ( .A(n37430), .B(n37431), .Z(n37429) );
  XNOR U37293 ( .A(n37428), .B(n37127), .Z(n37431) );
  XOR U37294 ( .A(n37329), .B(n37432), .Z(n37127) );
  AND U37295 ( .A(n621), .B(n37433), .Z(n37432) );
  XOR U37296 ( .A(n37325), .B(n37329), .Z(n37433) );
  XNOR U37297 ( .A(n37434), .B(n37428), .Z(n37430) );
  IV U37298 ( .A(n37076), .Z(n37434) );
  XOR U37299 ( .A(n37435), .B(n37436), .Z(n37076) );
  AND U37300 ( .A(n637), .B(n37437), .Z(n37436) );
  AND U37301 ( .A(n37389), .B(n37370), .Z(n37428) );
  XNOR U37302 ( .A(n37438), .B(n37439), .Z(n37370) );
  AND U37303 ( .A(n621), .B(n37348), .Z(n37439) );
  XNOR U37304 ( .A(n37346), .B(n37438), .Z(n37348) );
  XNOR U37305 ( .A(n37440), .B(n37441), .Z(n621) );
  AND U37306 ( .A(n37442), .B(n37443), .Z(n37441) );
  XNOR U37307 ( .A(n37440), .B(n37139), .Z(n37443) );
  IV U37308 ( .A(n37143), .Z(n37139) );
  XOR U37309 ( .A(n37444), .B(n37445), .Z(n37143) );
  AND U37310 ( .A(n625), .B(n37446), .Z(n37445) );
  XOR U37311 ( .A(n37447), .B(n37444), .Z(n37446) );
  XNOR U37312 ( .A(n37440), .B(n37353), .Z(n37442) );
  XOR U37313 ( .A(n37448), .B(n37449), .Z(n37353) );
  AND U37314 ( .A(n633), .B(n37400), .Z(n37449) );
  XOR U37315 ( .A(n37398), .B(n37448), .Z(n37400) );
  XOR U37316 ( .A(n37450), .B(n37451), .Z(n37440) );
  AND U37317 ( .A(n37452), .B(n37453), .Z(n37451) );
  XNOR U37318 ( .A(n37450), .B(n37155), .Z(n37453) );
  IV U37319 ( .A(n37158), .Z(n37155) );
  XOR U37320 ( .A(n37454), .B(n37455), .Z(n37158) );
  AND U37321 ( .A(n625), .B(n37456), .Z(n37455) );
  XOR U37322 ( .A(n37457), .B(n37454), .Z(n37456) );
  XOR U37323 ( .A(n37159), .B(n37450), .Z(n37452) );
  XOR U37324 ( .A(n37458), .B(n37459), .Z(n37159) );
  AND U37325 ( .A(n633), .B(n37410), .Z(n37459) );
  XOR U37326 ( .A(n37458), .B(n37408), .Z(n37410) );
  XOR U37327 ( .A(n37460), .B(n37461), .Z(n37450) );
  AND U37328 ( .A(n37462), .B(n37463), .Z(n37461) );
  XNOR U37329 ( .A(n37460), .B(n37183), .Z(n37463) );
  IV U37330 ( .A(n37186), .Z(n37183) );
  XOR U37331 ( .A(n37464), .B(n37465), .Z(n37186) );
  AND U37332 ( .A(n625), .B(n37466), .Z(n37465) );
  XNOR U37333 ( .A(n37467), .B(n37464), .Z(n37466) );
  XOR U37334 ( .A(n37187), .B(n37460), .Z(n37462) );
  XOR U37335 ( .A(n37468), .B(n37469), .Z(n37187) );
  AND U37336 ( .A(n633), .B(n37419), .Z(n37469) );
  XOR U37337 ( .A(n37468), .B(n37417), .Z(n37419) );
  XOR U37338 ( .A(n37470), .B(n37471), .Z(n37460) );
  AND U37339 ( .A(n37472), .B(n37473), .Z(n37471) );
  XNOR U37340 ( .A(n37470), .B(n37232), .Z(n37473) );
  IV U37341 ( .A(n37235), .Z(n37232) );
  XOR U37342 ( .A(n37474), .B(n37475), .Z(n37235) );
  AND U37343 ( .A(n625), .B(n37476), .Z(n37475) );
  XOR U37344 ( .A(n37477), .B(n37474), .Z(n37476) );
  XOR U37345 ( .A(n37236), .B(n37470), .Z(n37472) );
  XOR U37346 ( .A(n37478), .B(n37479), .Z(n37236) );
  AND U37347 ( .A(n633), .B(n37427), .Z(n37479) );
  XOR U37348 ( .A(n37478), .B(n37425), .Z(n37427) );
  XOR U37349 ( .A(n37366), .B(n37480), .Z(n37470) );
  AND U37350 ( .A(n37368), .B(n37481), .Z(n37480) );
  XNOR U37351 ( .A(n37366), .B(n37325), .Z(n37481) );
  IV U37352 ( .A(n37328), .Z(n37325) );
  XOR U37353 ( .A(n37482), .B(n37483), .Z(n37328) );
  AND U37354 ( .A(n625), .B(n37484), .Z(n37483) );
  XNOR U37355 ( .A(n37485), .B(n37482), .Z(n37484) );
  XOR U37356 ( .A(n37329), .B(n37366), .Z(n37368) );
  XOR U37357 ( .A(n37486), .B(n37487), .Z(n37329) );
  AND U37358 ( .A(n633), .B(n37437), .Z(n37487) );
  XOR U37359 ( .A(n37486), .B(n37435), .Z(n37437) );
  AND U37360 ( .A(n37438), .B(n37346), .Z(n37366) );
  XNOR U37361 ( .A(n37488), .B(n37489), .Z(n37346) );
  AND U37362 ( .A(n625), .B(n37490), .Z(n37489) );
  XNOR U37363 ( .A(n37491), .B(n37488), .Z(n37490) );
  XNOR U37364 ( .A(n37492), .B(n37493), .Z(n625) );
  AND U37365 ( .A(n37494), .B(n37495), .Z(n37493) );
  XOR U37366 ( .A(n37447), .B(n37492), .Z(n37495) );
  AND U37367 ( .A(n37496), .B(n37497), .Z(n37447) );
  XNOR U37368 ( .A(n37444), .B(n37492), .Z(n37494) );
  XNOR U37369 ( .A(n37498), .B(n37499), .Z(n37444) );
  AND U37370 ( .A(n629), .B(n37500), .Z(n37499) );
  XNOR U37371 ( .A(n37501), .B(n37502), .Z(n37500) );
  XOR U37372 ( .A(n37503), .B(n37504), .Z(n37492) );
  AND U37373 ( .A(n37505), .B(n37506), .Z(n37504) );
  XNOR U37374 ( .A(n37503), .B(n37496), .Z(n37506) );
  IV U37375 ( .A(n37457), .Z(n37496) );
  XOR U37376 ( .A(n37507), .B(n37508), .Z(n37457) );
  XOR U37377 ( .A(n37509), .B(n37497), .Z(n37508) );
  AND U37378 ( .A(n37467), .B(n37510), .Z(n37497) );
  AND U37379 ( .A(n37511), .B(n37512), .Z(n37509) );
  XOR U37380 ( .A(n37513), .B(n37507), .Z(n37511) );
  XNOR U37381 ( .A(n37454), .B(n37503), .Z(n37505) );
  XNOR U37382 ( .A(n37514), .B(n37515), .Z(n37454) );
  AND U37383 ( .A(n629), .B(n37516), .Z(n37515) );
  XNOR U37384 ( .A(n37517), .B(n37518), .Z(n37516) );
  XOR U37385 ( .A(n37519), .B(n37520), .Z(n37503) );
  AND U37386 ( .A(n37521), .B(n37522), .Z(n37520) );
  XNOR U37387 ( .A(n37519), .B(n37467), .Z(n37522) );
  XOR U37388 ( .A(n37523), .B(n37512), .Z(n37467) );
  XNOR U37389 ( .A(n37524), .B(n37507), .Z(n37512) );
  XOR U37390 ( .A(n37525), .B(n37526), .Z(n37507) );
  AND U37391 ( .A(n37527), .B(n37528), .Z(n37526) );
  XOR U37392 ( .A(n37529), .B(n37525), .Z(n37527) );
  XNOR U37393 ( .A(n37530), .B(n37531), .Z(n37524) );
  AND U37394 ( .A(n37532), .B(n37533), .Z(n37531) );
  XOR U37395 ( .A(n37530), .B(n37534), .Z(n37532) );
  XNOR U37396 ( .A(n37513), .B(n37510), .Z(n37523) );
  AND U37397 ( .A(n37535), .B(n37536), .Z(n37510) );
  XOR U37398 ( .A(n37537), .B(n37538), .Z(n37513) );
  AND U37399 ( .A(n37539), .B(n37540), .Z(n37538) );
  XOR U37400 ( .A(n37537), .B(n37541), .Z(n37539) );
  XNOR U37401 ( .A(n37464), .B(n37519), .Z(n37521) );
  XNOR U37402 ( .A(n37542), .B(n37543), .Z(n37464) );
  AND U37403 ( .A(n629), .B(n37544), .Z(n37543) );
  XNOR U37404 ( .A(n37545), .B(n37546), .Z(n37544) );
  XOR U37405 ( .A(n37547), .B(n37548), .Z(n37519) );
  AND U37406 ( .A(n37549), .B(n37550), .Z(n37548) );
  XNOR U37407 ( .A(n37547), .B(n37535), .Z(n37550) );
  IV U37408 ( .A(n37477), .Z(n37535) );
  XNOR U37409 ( .A(n37551), .B(n37528), .Z(n37477) );
  XNOR U37410 ( .A(n37552), .B(n37534), .Z(n37528) );
  XOR U37411 ( .A(n37553), .B(n37554), .Z(n37534) );
  AND U37412 ( .A(n37555), .B(n37556), .Z(n37554) );
  XOR U37413 ( .A(n37553), .B(n37557), .Z(n37555) );
  XNOR U37414 ( .A(n37533), .B(n37525), .Z(n37552) );
  XOR U37415 ( .A(n37558), .B(n37559), .Z(n37525) );
  AND U37416 ( .A(n37560), .B(n37561), .Z(n37559) );
  XNOR U37417 ( .A(n37562), .B(n37558), .Z(n37560) );
  XNOR U37418 ( .A(n37563), .B(n37530), .Z(n37533) );
  XOR U37419 ( .A(n37564), .B(n37565), .Z(n37530) );
  AND U37420 ( .A(n37566), .B(n37567), .Z(n37565) );
  XOR U37421 ( .A(n37564), .B(n37568), .Z(n37566) );
  XNOR U37422 ( .A(n37569), .B(n37570), .Z(n37563) );
  AND U37423 ( .A(n37571), .B(n37572), .Z(n37570) );
  XNOR U37424 ( .A(n37569), .B(n37573), .Z(n37571) );
  XNOR U37425 ( .A(n37529), .B(n37536), .Z(n37551) );
  AND U37426 ( .A(n37485), .B(n37574), .Z(n37536) );
  XOR U37427 ( .A(n37541), .B(n37540), .Z(n37529) );
  XNOR U37428 ( .A(n37575), .B(n37537), .Z(n37540) );
  XOR U37429 ( .A(n37576), .B(n37577), .Z(n37537) );
  AND U37430 ( .A(n37578), .B(n37579), .Z(n37577) );
  XOR U37431 ( .A(n37576), .B(n37580), .Z(n37578) );
  XNOR U37432 ( .A(n37581), .B(n37582), .Z(n37575) );
  AND U37433 ( .A(n37583), .B(n37584), .Z(n37582) );
  XOR U37434 ( .A(n37581), .B(n37585), .Z(n37583) );
  XOR U37435 ( .A(n37586), .B(n37587), .Z(n37541) );
  AND U37436 ( .A(n37588), .B(n37589), .Z(n37587) );
  XOR U37437 ( .A(n37586), .B(n37590), .Z(n37588) );
  XNOR U37438 ( .A(n37474), .B(n37547), .Z(n37549) );
  XNOR U37439 ( .A(n37591), .B(n37592), .Z(n37474) );
  AND U37440 ( .A(n629), .B(n37593), .Z(n37592) );
  XNOR U37441 ( .A(n37594), .B(n37595), .Z(n37593) );
  XOR U37442 ( .A(n37596), .B(n37597), .Z(n37547) );
  AND U37443 ( .A(n37598), .B(n37599), .Z(n37597) );
  XNOR U37444 ( .A(n37596), .B(n37485), .Z(n37599) );
  XOR U37445 ( .A(n37600), .B(n37561), .Z(n37485) );
  XNOR U37446 ( .A(n37601), .B(n37568), .Z(n37561) );
  XOR U37447 ( .A(n37557), .B(n37556), .Z(n37568) );
  XNOR U37448 ( .A(n37602), .B(n37553), .Z(n37556) );
  XOR U37449 ( .A(n37603), .B(n37604), .Z(n37553) );
  AND U37450 ( .A(n37605), .B(n37606), .Z(n37604) );
  XOR U37451 ( .A(n37603), .B(n37607), .Z(n37605) );
  XNOR U37452 ( .A(n37608), .B(n37609), .Z(n37602) );
  NOR U37453 ( .A(n37610), .B(n37611), .Z(n37609) );
  XNOR U37454 ( .A(n37608), .B(n37612), .Z(n37610) );
  XOR U37455 ( .A(n37613), .B(n37614), .Z(n37557) );
  NOR U37456 ( .A(n37615), .B(n37616), .Z(n37614) );
  XNOR U37457 ( .A(n37613), .B(n37617), .Z(n37615) );
  XNOR U37458 ( .A(n37567), .B(n37558), .Z(n37601) );
  XOR U37459 ( .A(n37618), .B(n37619), .Z(n37558) );
  NOR U37460 ( .A(n37620), .B(n37621), .Z(n37619) );
  XNOR U37461 ( .A(n37618), .B(n37622), .Z(n37620) );
  XOR U37462 ( .A(n37623), .B(n37573), .Z(n37567) );
  XNOR U37463 ( .A(n37624), .B(n37625), .Z(n37573) );
  NOR U37464 ( .A(n37626), .B(n37627), .Z(n37625) );
  XNOR U37465 ( .A(n37624), .B(n37628), .Z(n37626) );
  XNOR U37466 ( .A(n37572), .B(n37564), .Z(n37623) );
  XOR U37467 ( .A(n37629), .B(n37630), .Z(n37564) );
  AND U37468 ( .A(n37631), .B(n37632), .Z(n37630) );
  XOR U37469 ( .A(n37629), .B(n37633), .Z(n37631) );
  XNOR U37470 ( .A(n37634), .B(n37569), .Z(n37572) );
  XOR U37471 ( .A(n37635), .B(n37636), .Z(n37569) );
  AND U37472 ( .A(n37637), .B(n37638), .Z(n37636) );
  XOR U37473 ( .A(n37635), .B(n37639), .Z(n37637) );
  XNOR U37474 ( .A(n37640), .B(n37641), .Z(n37634) );
  NOR U37475 ( .A(n37642), .B(n37643), .Z(n37641) );
  XOR U37476 ( .A(n37640), .B(n37644), .Z(n37642) );
  XOR U37477 ( .A(n37562), .B(n37574), .Z(n37600) );
  NOR U37478 ( .A(n37491), .B(n37645), .Z(n37574) );
  XNOR U37479 ( .A(n37580), .B(n37579), .Z(n37562) );
  XNOR U37480 ( .A(n37646), .B(n37585), .Z(n37579) );
  XOR U37481 ( .A(n37647), .B(n37648), .Z(n37585) );
  NOR U37482 ( .A(n37649), .B(n37650), .Z(n37648) );
  XNOR U37483 ( .A(n37647), .B(n37651), .Z(n37649) );
  XNOR U37484 ( .A(n37584), .B(n37576), .Z(n37646) );
  XOR U37485 ( .A(n37652), .B(n37653), .Z(n37576) );
  AND U37486 ( .A(n37654), .B(n37655), .Z(n37653) );
  XNOR U37487 ( .A(n37652), .B(n37656), .Z(n37654) );
  XNOR U37488 ( .A(n37657), .B(n37581), .Z(n37584) );
  XOR U37489 ( .A(n37658), .B(n37659), .Z(n37581) );
  AND U37490 ( .A(n37660), .B(n37661), .Z(n37659) );
  XOR U37491 ( .A(n37658), .B(n37662), .Z(n37660) );
  XNOR U37492 ( .A(n37663), .B(n37664), .Z(n37657) );
  NOR U37493 ( .A(n37665), .B(n37666), .Z(n37664) );
  XOR U37494 ( .A(n37663), .B(n37667), .Z(n37665) );
  XOR U37495 ( .A(n37590), .B(n37589), .Z(n37580) );
  XNOR U37496 ( .A(n37668), .B(n37586), .Z(n37589) );
  XOR U37497 ( .A(n37669), .B(n37670), .Z(n37586) );
  AND U37498 ( .A(n37671), .B(n37672), .Z(n37670) );
  XOR U37499 ( .A(n37669), .B(n37673), .Z(n37671) );
  XNOR U37500 ( .A(n37674), .B(n37675), .Z(n37668) );
  NOR U37501 ( .A(n37676), .B(n37677), .Z(n37675) );
  XNOR U37502 ( .A(n37674), .B(n37678), .Z(n37676) );
  XOR U37503 ( .A(n37679), .B(n37680), .Z(n37590) );
  NOR U37504 ( .A(n37681), .B(n37682), .Z(n37680) );
  XNOR U37505 ( .A(n37679), .B(n37683), .Z(n37681) );
  XNOR U37506 ( .A(n37482), .B(n37596), .Z(n37598) );
  XNOR U37507 ( .A(n37684), .B(n37685), .Z(n37482) );
  AND U37508 ( .A(n629), .B(n37686), .Z(n37685) );
  XNOR U37509 ( .A(n37687), .B(n37688), .Z(n37686) );
  AND U37510 ( .A(n37488), .B(n37491), .Z(n37596) );
  XOR U37511 ( .A(n37689), .B(n37645), .Z(n37491) );
  XNOR U37512 ( .A(p_input[2048]), .B(p_input[832]), .Z(n37645) );
  XOR U37513 ( .A(n37622), .B(n37621), .Z(n37689) );
  XOR U37514 ( .A(n37690), .B(n37633), .Z(n37621) );
  XOR U37515 ( .A(n37607), .B(n37606), .Z(n37633) );
  XNOR U37516 ( .A(n37691), .B(n37612), .Z(n37606) );
  XOR U37517 ( .A(p_input[2072]), .B(p_input[856]), .Z(n37612) );
  XOR U37518 ( .A(n37603), .B(n37611), .Z(n37691) );
  XOR U37519 ( .A(n37692), .B(n37608), .Z(n37611) );
  XOR U37520 ( .A(p_input[2070]), .B(p_input[854]), .Z(n37608) );
  XNOR U37521 ( .A(p_input[2071]), .B(p_input[855]), .Z(n37692) );
  XNOR U37522 ( .A(n28684), .B(p_input[850]), .Z(n37603) );
  XNOR U37523 ( .A(n37617), .B(n37616), .Z(n37607) );
  XOR U37524 ( .A(n37693), .B(n37613), .Z(n37616) );
  XOR U37525 ( .A(p_input[2067]), .B(p_input[851]), .Z(n37613) );
  XNOR U37526 ( .A(p_input[2068]), .B(p_input[852]), .Z(n37693) );
  XOR U37527 ( .A(p_input[2069]), .B(p_input[853]), .Z(n37617) );
  XNOR U37528 ( .A(n37632), .B(n37618), .Z(n37690) );
  XNOR U37529 ( .A(n28686), .B(p_input[833]), .Z(n37618) );
  XNOR U37530 ( .A(n37694), .B(n37639), .Z(n37632) );
  XNOR U37531 ( .A(n37628), .B(n37627), .Z(n37639) );
  XOR U37532 ( .A(n37695), .B(n37624), .Z(n37627) );
  XNOR U37533 ( .A(n28322), .B(p_input[858]), .Z(n37624) );
  XNOR U37534 ( .A(p_input[2075]), .B(p_input[859]), .Z(n37695) );
  XOR U37535 ( .A(p_input[2076]), .B(p_input[860]), .Z(n37628) );
  XNOR U37536 ( .A(n37638), .B(n37629), .Z(n37694) );
  XNOR U37537 ( .A(n28689), .B(p_input[849]), .Z(n37629) );
  XOR U37538 ( .A(n37696), .B(n37644), .Z(n37638) );
  XNOR U37539 ( .A(p_input[2079]), .B(p_input[863]), .Z(n37644) );
  XOR U37540 ( .A(n37635), .B(n37643), .Z(n37696) );
  XOR U37541 ( .A(n37697), .B(n37640), .Z(n37643) );
  XOR U37542 ( .A(p_input[2077]), .B(p_input[861]), .Z(n37640) );
  XNOR U37543 ( .A(p_input[2078]), .B(p_input[862]), .Z(n37697) );
  XNOR U37544 ( .A(n28326), .B(p_input[857]), .Z(n37635) );
  XNOR U37545 ( .A(n37656), .B(n37655), .Z(n37622) );
  XNOR U37546 ( .A(n37698), .B(n37662), .Z(n37655) );
  XNOR U37547 ( .A(n37651), .B(n37650), .Z(n37662) );
  XOR U37548 ( .A(n37699), .B(n37647), .Z(n37650) );
  XNOR U37549 ( .A(n28694), .B(p_input[843]), .Z(n37647) );
  XNOR U37550 ( .A(p_input[2060]), .B(p_input[844]), .Z(n37699) );
  XOR U37551 ( .A(p_input[2061]), .B(p_input[845]), .Z(n37651) );
  XNOR U37552 ( .A(n37661), .B(n37652), .Z(n37698) );
  XNOR U37553 ( .A(n28330), .B(p_input[834]), .Z(n37652) );
  XOR U37554 ( .A(n37700), .B(n37667), .Z(n37661) );
  XNOR U37555 ( .A(p_input[2064]), .B(p_input[848]), .Z(n37667) );
  XOR U37556 ( .A(n37658), .B(n37666), .Z(n37700) );
  XOR U37557 ( .A(n37701), .B(n37663), .Z(n37666) );
  XOR U37558 ( .A(p_input[2062]), .B(p_input[846]), .Z(n37663) );
  XNOR U37559 ( .A(p_input[2063]), .B(p_input[847]), .Z(n37701) );
  XNOR U37560 ( .A(n28697), .B(p_input[842]), .Z(n37658) );
  XNOR U37561 ( .A(n37673), .B(n37672), .Z(n37656) );
  XNOR U37562 ( .A(n37702), .B(n37678), .Z(n37672) );
  XOR U37563 ( .A(p_input[2057]), .B(p_input[841]), .Z(n37678) );
  XOR U37564 ( .A(n37669), .B(n37677), .Z(n37702) );
  XOR U37565 ( .A(n37703), .B(n37674), .Z(n37677) );
  XOR U37566 ( .A(p_input[2055]), .B(p_input[839]), .Z(n37674) );
  XNOR U37567 ( .A(p_input[2056]), .B(p_input[840]), .Z(n37703) );
  XNOR U37568 ( .A(n28337), .B(p_input[835]), .Z(n37669) );
  XNOR U37569 ( .A(n37683), .B(n37682), .Z(n37673) );
  XOR U37570 ( .A(n37704), .B(n37679), .Z(n37682) );
  XOR U37571 ( .A(p_input[2052]), .B(p_input[836]), .Z(n37679) );
  XNOR U37572 ( .A(p_input[2053]), .B(p_input[837]), .Z(n37704) );
  XOR U37573 ( .A(p_input[2054]), .B(p_input[838]), .Z(n37683) );
  XNOR U37574 ( .A(n37705), .B(n37706), .Z(n37488) );
  AND U37575 ( .A(n629), .B(n37707), .Z(n37706) );
  XNOR U37576 ( .A(n37708), .B(n37709), .Z(n629) );
  AND U37577 ( .A(n37710), .B(n37711), .Z(n37709) );
  XOR U37578 ( .A(n37502), .B(n37708), .Z(n37711) );
  XNOR U37579 ( .A(n37712), .B(n37708), .Z(n37710) );
  XOR U37580 ( .A(n37713), .B(n37714), .Z(n37708) );
  AND U37581 ( .A(n37715), .B(n37716), .Z(n37714) );
  XOR U37582 ( .A(n37517), .B(n37713), .Z(n37716) );
  XOR U37583 ( .A(n37713), .B(n37518), .Z(n37715) );
  XOR U37584 ( .A(n37717), .B(n37718), .Z(n37713) );
  AND U37585 ( .A(n37719), .B(n37720), .Z(n37718) );
  XOR U37586 ( .A(n37545), .B(n37717), .Z(n37720) );
  XOR U37587 ( .A(n37717), .B(n37546), .Z(n37719) );
  XOR U37588 ( .A(n37721), .B(n37722), .Z(n37717) );
  AND U37589 ( .A(n37723), .B(n37724), .Z(n37722) );
  XOR U37590 ( .A(n37594), .B(n37721), .Z(n37724) );
  XOR U37591 ( .A(n37721), .B(n37595), .Z(n37723) );
  XOR U37592 ( .A(n37725), .B(n37726), .Z(n37721) );
  AND U37593 ( .A(n37727), .B(n37728), .Z(n37726) );
  XOR U37594 ( .A(n37725), .B(n37687), .Z(n37728) );
  XNOR U37595 ( .A(n37729), .B(n37730), .Z(n37438) );
  AND U37596 ( .A(n633), .B(n37731), .Z(n37730) );
  XNOR U37597 ( .A(n37732), .B(n37733), .Z(n633) );
  AND U37598 ( .A(n37734), .B(n37735), .Z(n37733) );
  XOR U37599 ( .A(n37732), .B(n37448), .Z(n37735) );
  XNOR U37600 ( .A(n37732), .B(n37398), .Z(n37734) );
  XOR U37601 ( .A(n37736), .B(n37737), .Z(n37732) );
  AND U37602 ( .A(n37738), .B(n37739), .Z(n37737) );
  XNOR U37603 ( .A(n37458), .B(n37736), .Z(n37739) );
  XOR U37604 ( .A(n37736), .B(n37408), .Z(n37738) );
  XOR U37605 ( .A(n37740), .B(n37741), .Z(n37736) );
  AND U37606 ( .A(n37742), .B(n37743), .Z(n37741) );
  XNOR U37607 ( .A(n37468), .B(n37740), .Z(n37743) );
  XOR U37608 ( .A(n37740), .B(n37417), .Z(n37742) );
  XOR U37609 ( .A(n37744), .B(n37745), .Z(n37740) );
  AND U37610 ( .A(n37746), .B(n37747), .Z(n37745) );
  XOR U37611 ( .A(n37744), .B(n37425), .Z(n37746) );
  XOR U37612 ( .A(n37748), .B(n37749), .Z(n37389) );
  AND U37613 ( .A(n637), .B(n37731), .Z(n37749) );
  XNOR U37614 ( .A(n37729), .B(n37748), .Z(n37731) );
  XNOR U37615 ( .A(n37750), .B(n37751), .Z(n637) );
  AND U37616 ( .A(n37752), .B(n37753), .Z(n37751) );
  XNOR U37617 ( .A(n37754), .B(n37750), .Z(n37753) );
  IV U37618 ( .A(n37448), .Z(n37754) );
  XOR U37619 ( .A(n37712), .B(n37755), .Z(n37448) );
  AND U37620 ( .A(n640), .B(n37756), .Z(n37755) );
  XOR U37621 ( .A(n37501), .B(n37498), .Z(n37756) );
  IV U37622 ( .A(n37712), .Z(n37501) );
  XNOR U37623 ( .A(n37398), .B(n37750), .Z(n37752) );
  XOR U37624 ( .A(n37757), .B(n37758), .Z(n37398) );
  AND U37625 ( .A(n656), .B(n37759), .Z(n37758) );
  XOR U37626 ( .A(n37760), .B(n37761), .Z(n37750) );
  AND U37627 ( .A(n37762), .B(n37763), .Z(n37761) );
  XNOR U37628 ( .A(n37760), .B(n37458), .Z(n37763) );
  XOR U37629 ( .A(n37518), .B(n37764), .Z(n37458) );
  AND U37630 ( .A(n640), .B(n37765), .Z(n37764) );
  XOR U37631 ( .A(n37514), .B(n37518), .Z(n37765) );
  XNOR U37632 ( .A(n37766), .B(n37760), .Z(n37762) );
  IV U37633 ( .A(n37408), .Z(n37766) );
  XOR U37634 ( .A(n37767), .B(n37768), .Z(n37408) );
  AND U37635 ( .A(n656), .B(n37769), .Z(n37768) );
  XOR U37636 ( .A(n37770), .B(n37771), .Z(n37760) );
  AND U37637 ( .A(n37772), .B(n37773), .Z(n37771) );
  XNOR U37638 ( .A(n37770), .B(n37468), .Z(n37773) );
  XOR U37639 ( .A(n37546), .B(n37774), .Z(n37468) );
  AND U37640 ( .A(n640), .B(n37775), .Z(n37774) );
  XOR U37641 ( .A(n37542), .B(n37546), .Z(n37775) );
  XOR U37642 ( .A(n37417), .B(n37770), .Z(n37772) );
  XOR U37643 ( .A(n37776), .B(n37777), .Z(n37417) );
  AND U37644 ( .A(n656), .B(n37778), .Z(n37777) );
  XOR U37645 ( .A(n37744), .B(n37779), .Z(n37770) );
  AND U37646 ( .A(n37780), .B(n37747), .Z(n37779) );
  XNOR U37647 ( .A(n37478), .B(n37744), .Z(n37747) );
  XOR U37648 ( .A(n37595), .B(n37781), .Z(n37478) );
  AND U37649 ( .A(n640), .B(n37782), .Z(n37781) );
  XOR U37650 ( .A(n37591), .B(n37595), .Z(n37782) );
  XNOR U37651 ( .A(n37783), .B(n37744), .Z(n37780) );
  IV U37652 ( .A(n37425), .Z(n37783) );
  XOR U37653 ( .A(n37784), .B(n37785), .Z(n37425) );
  AND U37654 ( .A(n656), .B(n37786), .Z(n37785) );
  XOR U37655 ( .A(n37787), .B(n37788), .Z(n37744) );
  AND U37656 ( .A(n37789), .B(n37790), .Z(n37788) );
  XNOR U37657 ( .A(n37787), .B(n37486), .Z(n37790) );
  XOR U37658 ( .A(n37688), .B(n37791), .Z(n37486) );
  AND U37659 ( .A(n640), .B(n37792), .Z(n37791) );
  XOR U37660 ( .A(n37684), .B(n37688), .Z(n37792) );
  XNOR U37661 ( .A(n37793), .B(n37787), .Z(n37789) );
  IV U37662 ( .A(n37435), .Z(n37793) );
  XOR U37663 ( .A(n37794), .B(n37795), .Z(n37435) );
  AND U37664 ( .A(n656), .B(n37796), .Z(n37795) );
  AND U37665 ( .A(n37748), .B(n37729), .Z(n37787) );
  XNOR U37666 ( .A(n37797), .B(n37798), .Z(n37729) );
  AND U37667 ( .A(n640), .B(n37707), .Z(n37798) );
  XNOR U37668 ( .A(n37705), .B(n37797), .Z(n37707) );
  XNOR U37669 ( .A(n37799), .B(n37800), .Z(n640) );
  AND U37670 ( .A(n37801), .B(n37802), .Z(n37800) );
  XNOR U37671 ( .A(n37799), .B(n37498), .Z(n37802) );
  IV U37672 ( .A(n37502), .Z(n37498) );
  XOR U37673 ( .A(n37803), .B(n37804), .Z(n37502) );
  AND U37674 ( .A(n644), .B(n37805), .Z(n37804) );
  XOR U37675 ( .A(n37806), .B(n37803), .Z(n37805) );
  XNOR U37676 ( .A(n37799), .B(n37712), .Z(n37801) );
  XOR U37677 ( .A(n37807), .B(n37808), .Z(n37712) );
  AND U37678 ( .A(n652), .B(n37759), .Z(n37808) );
  XOR U37679 ( .A(n37757), .B(n37807), .Z(n37759) );
  XOR U37680 ( .A(n37809), .B(n37810), .Z(n37799) );
  AND U37681 ( .A(n37811), .B(n37812), .Z(n37810) );
  XNOR U37682 ( .A(n37809), .B(n37514), .Z(n37812) );
  IV U37683 ( .A(n37517), .Z(n37514) );
  XOR U37684 ( .A(n37813), .B(n37814), .Z(n37517) );
  AND U37685 ( .A(n644), .B(n37815), .Z(n37814) );
  XOR U37686 ( .A(n37816), .B(n37813), .Z(n37815) );
  XOR U37687 ( .A(n37518), .B(n37809), .Z(n37811) );
  XOR U37688 ( .A(n37817), .B(n37818), .Z(n37518) );
  AND U37689 ( .A(n652), .B(n37769), .Z(n37818) );
  XOR U37690 ( .A(n37817), .B(n37767), .Z(n37769) );
  XOR U37691 ( .A(n37819), .B(n37820), .Z(n37809) );
  AND U37692 ( .A(n37821), .B(n37822), .Z(n37820) );
  XNOR U37693 ( .A(n37819), .B(n37542), .Z(n37822) );
  IV U37694 ( .A(n37545), .Z(n37542) );
  XOR U37695 ( .A(n37823), .B(n37824), .Z(n37545) );
  AND U37696 ( .A(n644), .B(n37825), .Z(n37824) );
  XNOR U37697 ( .A(n37826), .B(n37823), .Z(n37825) );
  XOR U37698 ( .A(n37546), .B(n37819), .Z(n37821) );
  XOR U37699 ( .A(n37827), .B(n37828), .Z(n37546) );
  AND U37700 ( .A(n652), .B(n37778), .Z(n37828) );
  XOR U37701 ( .A(n37827), .B(n37776), .Z(n37778) );
  XOR U37702 ( .A(n37829), .B(n37830), .Z(n37819) );
  AND U37703 ( .A(n37831), .B(n37832), .Z(n37830) );
  XNOR U37704 ( .A(n37829), .B(n37591), .Z(n37832) );
  IV U37705 ( .A(n37594), .Z(n37591) );
  XOR U37706 ( .A(n37833), .B(n37834), .Z(n37594) );
  AND U37707 ( .A(n644), .B(n37835), .Z(n37834) );
  XOR U37708 ( .A(n37836), .B(n37833), .Z(n37835) );
  XOR U37709 ( .A(n37595), .B(n37829), .Z(n37831) );
  XOR U37710 ( .A(n37837), .B(n37838), .Z(n37595) );
  AND U37711 ( .A(n652), .B(n37786), .Z(n37838) );
  XOR U37712 ( .A(n37837), .B(n37784), .Z(n37786) );
  XOR U37713 ( .A(n37725), .B(n37839), .Z(n37829) );
  AND U37714 ( .A(n37727), .B(n37840), .Z(n37839) );
  XNOR U37715 ( .A(n37725), .B(n37684), .Z(n37840) );
  IV U37716 ( .A(n37687), .Z(n37684) );
  XOR U37717 ( .A(n37841), .B(n37842), .Z(n37687) );
  AND U37718 ( .A(n644), .B(n37843), .Z(n37842) );
  XNOR U37719 ( .A(n37844), .B(n37841), .Z(n37843) );
  XOR U37720 ( .A(n37688), .B(n37725), .Z(n37727) );
  XOR U37721 ( .A(n37845), .B(n37846), .Z(n37688) );
  AND U37722 ( .A(n652), .B(n37796), .Z(n37846) );
  XOR U37723 ( .A(n37845), .B(n37794), .Z(n37796) );
  AND U37724 ( .A(n37797), .B(n37705), .Z(n37725) );
  XNOR U37725 ( .A(n37847), .B(n37848), .Z(n37705) );
  AND U37726 ( .A(n644), .B(n37849), .Z(n37848) );
  XNOR U37727 ( .A(n37850), .B(n37847), .Z(n37849) );
  XNOR U37728 ( .A(n37851), .B(n37852), .Z(n644) );
  AND U37729 ( .A(n37853), .B(n37854), .Z(n37852) );
  XOR U37730 ( .A(n37806), .B(n37851), .Z(n37854) );
  AND U37731 ( .A(n37855), .B(n37856), .Z(n37806) );
  XNOR U37732 ( .A(n37803), .B(n37851), .Z(n37853) );
  XNOR U37733 ( .A(n37857), .B(n37858), .Z(n37803) );
  AND U37734 ( .A(n648), .B(n37859), .Z(n37858) );
  XNOR U37735 ( .A(n37860), .B(n37861), .Z(n37859) );
  XOR U37736 ( .A(n37862), .B(n37863), .Z(n37851) );
  AND U37737 ( .A(n37864), .B(n37865), .Z(n37863) );
  XNOR U37738 ( .A(n37862), .B(n37855), .Z(n37865) );
  IV U37739 ( .A(n37816), .Z(n37855) );
  XOR U37740 ( .A(n37866), .B(n37867), .Z(n37816) );
  XOR U37741 ( .A(n37868), .B(n37856), .Z(n37867) );
  AND U37742 ( .A(n37826), .B(n37869), .Z(n37856) );
  AND U37743 ( .A(n37870), .B(n37871), .Z(n37868) );
  XOR U37744 ( .A(n37872), .B(n37866), .Z(n37870) );
  XNOR U37745 ( .A(n37813), .B(n37862), .Z(n37864) );
  XNOR U37746 ( .A(n37873), .B(n37874), .Z(n37813) );
  AND U37747 ( .A(n648), .B(n37875), .Z(n37874) );
  XNOR U37748 ( .A(n37876), .B(n37877), .Z(n37875) );
  XOR U37749 ( .A(n37878), .B(n37879), .Z(n37862) );
  AND U37750 ( .A(n37880), .B(n37881), .Z(n37879) );
  XNOR U37751 ( .A(n37878), .B(n37826), .Z(n37881) );
  XOR U37752 ( .A(n37882), .B(n37871), .Z(n37826) );
  XNOR U37753 ( .A(n37883), .B(n37866), .Z(n37871) );
  XOR U37754 ( .A(n37884), .B(n37885), .Z(n37866) );
  AND U37755 ( .A(n37886), .B(n37887), .Z(n37885) );
  XOR U37756 ( .A(n37888), .B(n37884), .Z(n37886) );
  XNOR U37757 ( .A(n37889), .B(n37890), .Z(n37883) );
  AND U37758 ( .A(n37891), .B(n37892), .Z(n37890) );
  XOR U37759 ( .A(n37889), .B(n37893), .Z(n37891) );
  XNOR U37760 ( .A(n37872), .B(n37869), .Z(n37882) );
  AND U37761 ( .A(n37894), .B(n37895), .Z(n37869) );
  XOR U37762 ( .A(n37896), .B(n37897), .Z(n37872) );
  AND U37763 ( .A(n37898), .B(n37899), .Z(n37897) );
  XOR U37764 ( .A(n37896), .B(n37900), .Z(n37898) );
  XNOR U37765 ( .A(n37823), .B(n37878), .Z(n37880) );
  XNOR U37766 ( .A(n37901), .B(n37902), .Z(n37823) );
  AND U37767 ( .A(n648), .B(n37903), .Z(n37902) );
  XNOR U37768 ( .A(n37904), .B(n37905), .Z(n37903) );
  XOR U37769 ( .A(n37906), .B(n37907), .Z(n37878) );
  AND U37770 ( .A(n37908), .B(n37909), .Z(n37907) );
  XNOR U37771 ( .A(n37906), .B(n37894), .Z(n37909) );
  IV U37772 ( .A(n37836), .Z(n37894) );
  XNOR U37773 ( .A(n37910), .B(n37887), .Z(n37836) );
  XNOR U37774 ( .A(n37911), .B(n37893), .Z(n37887) );
  XOR U37775 ( .A(n37912), .B(n37913), .Z(n37893) );
  AND U37776 ( .A(n37914), .B(n37915), .Z(n37913) );
  XOR U37777 ( .A(n37912), .B(n37916), .Z(n37914) );
  XNOR U37778 ( .A(n37892), .B(n37884), .Z(n37911) );
  XOR U37779 ( .A(n37917), .B(n37918), .Z(n37884) );
  AND U37780 ( .A(n37919), .B(n37920), .Z(n37918) );
  XNOR U37781 ( .A(n37921), .B(n37917), .Z(n37919) );
  XNOR U37782 ( .A(n37922), .B(n37889), .Z(n37892) );
  XOR U37783 ( .A(n37923), .B(n37924), .Z(n37889) );
  AND U37784 ( .A(n37925), .B(n37926), .Z(n37924) );
  XOR U37785 ( .A(n37923), .B(n37927), .Z(n37925) );
  XNOR U37786 ( .A(n37928), .B(n37929), .Z(n37922) );
  AND U37787 ( .A(n37930), .B(n37931), .Z(n37929) );
  XNOR U37788 ( .A(n37928), .B(n37932), .Z(n37930) );
  XNOR U37789 ( .A(n37888), .B(n37895), .Z(n37910) );
  AND U37790 ( .A(n37844), .B(n37933), .Z(n37895) );
  XOR U37791 ( .A(n37900), .B(n37899), .Z(n37888) );
  XNOR U37792 ( .A(n37934), .B(n37896), .Z(n37899) );
  XOR U37793 ( .A(n37935), .B(n37936), .Z(n37896) );
  AND U37794 ( .A(n37937), .B(n37938), .Z(n37936) );
  XOR U37795 ( .A(n37935), .B(n37939), .Z(n37937) );
  XNOR U37796 ( .A(n37940), .B(n37941), .Z(n37934) );
  AND U37797 ( .A(n37942), .B(n37943), .Z(n37941) );
  XOR U37798 ( .A(n37940), .B(n37944), .Z(n37942) );
  XOR U37799 ( .A(n37945), .B(n37946), .Z(n37900) );
  AND U37800 ( .A(n37947), .B(n37948), .Z(n37946) );
  XOR U37801 ( .A(n37945), .B(n37949), .Z(n37947) );
  XNOR U37802 ( .A(n37833), .B(n37906), .Z(n37908) );
  XNOR U37803 ( .A(n37950), .B(n37951), .Z(n37833) );
  AND U37804 ( .A(n648), .B(n37952), .Z(n37951) );
  XNOR U37805 ( .A(n37953), .B(n37954), .Z(n37952) );
  XOR U37806 ( .A(n37955), .B(n37956), .Z(n37906) );
  AND U37807 ( .A(n37957), .B(n37958), .Z(n37956) );
  XNOR U37808 ( .A(n37955), .B(n37844), .Z(n37958) );
  XOR U37809 ( .A(n37959), .B(n37920), .Z(n37844) );
  XNOR U37810 ( .A(n37960), .B(n37927), .Z(n37920) );
  XOR U37811 ( .A(n37916), .B(n37915), .Z(n37927) );
  XNOR U37812 ( .A(n37961), .B(n37912), .Z(n37915) );
  XOR U37813 ( .A(n37962), .B(n37963), .Z(n37912) );
  AND U37814 ( .A(n37964), .B(n37965), .Z(n37963) );
  XOR U37815 ( .A(n37962), .B(n37966), .Z(n37964) );
  XNOR U37816 ( .A(n37967), .B(n37968), .Z(n37961) );
  NOR U37817 ( .A(n37969), .B(n37970), .Z(n37968) );
  XNOR U37818 ( .A(n37967), .B(n37971), .Z(n37969) );
  XOR U37819 ( .A(n37972), .B(n37973), .Z(n37916) );
  NOR U37820 ( .A(n37974), .B(n37975), .Z(n37973) );
  XNOR U37821 ( .A(n37972), .B(n37976), .Z(n37974) );
  XNOR U37822 ( .A(n37926), .B(n37917), .Z(n37960) );
  XOR U37823 ( .A(n37977), .B(n37978), .Z(n37917) );
  NOR U37824 ( .A(n37979), .B(n37980), .Z(n37978) );
  XNOR U37825 ( .A(n37977), .B(n37981), .Z(n37979) );
  XOR U37826 ( .A(n37982), .B(n37932), .Z(n37926) );
  XNOR U37827 ( .A(n37983), .B(n37984), .Z(n37932) );
  NOR U37828 ( .A(n37985), .B(n37986), .Z(n37984) );
  XNOR U37829 ( .A(n37983), .B(n37987), .Z(n37985) );
  XNOR U37830 ( .A(n37931), .B(n37923), .Z(n37982) );
  XOR U37831 ( .A(n37988), .B(n37989), .Z(n37923) );
  AND U37832 ( .A(n37990), .B(n37991), .Z(n37989) );
  XOR U37833 ( .A(n37988), .B(n37992), .Z(n37990) );
  XNOR U37834 ( .A(n37993), .B(n37928), .Z(n37931) );
  XOR U37835 ( .A(n37994), .B(n37995), .Z(n37928) );
  AND U37836 ( .A(n37996), .B(n37997), .Z(n37995) );
  XOR U37837 ( .A(n37994), .B(n37998), .Z(n37996) );
  XNOR U37838 ( .A(n37999), .B(n38000), .Z(n37993) );
  NOR U37839 ( .A(n38001), .B(n38002), .Z(n38000) );
  XOR U37840 ( .A(n37999), .B(n38003), .Z(n38001) );
  XOR U37841 ( .A(n37921), .B(n37933), .Z(n37959) );
  NOR U37842 ( .A(n37850), .B(n38004), .Z(n37933) );
  XNOR U37843 ( .A(n37939), .B(n37938), .Z(n37921) );
  XNOR U37844 ( .A(n38005), .B(n37944), .Z(n37938) );
  XOR U37845 ( .A(n38006), .B(n38007), .Z(n37944) );
  NOR U37846 ( .A(n38008), .B(n38009), .Z(n38007) );
  XNOR U37847 ( .A(n38006), .B(n38010), .Z(n38008) );
  XNOR U37848 ( .A(n37943), .B(n37935), .Z(n38005) );
  XOR U37849 ( .A(n38011), .B(n38012), .Z(n37935) );
  AND U37850 ( .A(n38013), .B(n38014), .Z(n38012) );
  XNOR U37851 ( .A(n38011), .B(n38015), .Z(n38013) );
  XNOR U37852 ( .A(n38016), .B(n37940), .Z(n37943) );
  XOR U37853 ( .A(n38017), .B(n38018), .Z(n37940) );
  AND U37854 ( .A(n38019), .B(n38020), .Z(n38018) );
  XOR U37855 ( .A(n38017), .B(n38021), .Z(n38019) );
  XNOR U37856 ( .A(n38022), .B(n38023), .Z(n38016) );
  NOR U37857 ( .A(n38024), .B(n38025), .Z(n38023) );
  XOR U37858 ( .A(n38022), .B(n38026), .Z(n38024) );
  XOR U37859 ( .A(n37949), .B(n37948), .Z(n37939) );
  XNOR U37860 ( .A(n38027), .B(n37945), .Z(n37948) );
  XOR U37861 ( .A(n38028), .B(n38029), .Z(n37945) );
  AND U37862 ( .A(n38030), .B(n38031), .Z(n38029) );
  XOR U37863 ( .A(n38028), .B(n38032), .Z(n38030) );
  XNOR U37864 ( .A(n38033), .B(n38034), .Z(n38027) );
  NOR U37865 ( .A(n38035), .B(n38036), .Z(n38034) );
  XNOR U37866 ( .A(n38033), .B(n38037), .Z(n38035) );
  XOR U37867 ( .A(n38038), .B(n38039), .Z(n37949) );
  NOR U37868 ( .A(n38040), .B(n38041), .Z(n38039) );
  XNOR U37869 ( .A(n38038), .B(n38042), .Z(n38040) );
  XNOR U37870 ( .A(n37841), .B(n37955), .Z(n37957) );
  XNOR U37871 ( .A(n38043), .B(n38044), .Z(n37841) );
  AND U37872 ( .A(n648), .B(n38045), .Z(n38044) );
  XNOR U37873 ( .A(n38046), .B(n38047), .Z(n38045) );
  AND U37874 ( .A(n37847), .B(n37850), .Z(n37955) );
  XOR U37875 ( .A(n38048), .B(n38004), .Z(n37850) );
  XNOR U37876 ( .A(p_input[2048]), .B(p_input[864]), .Z(n38004) );
  XOR U37877 ( .A(n37981), .B(n37980), .Z(n38048) );
  XOR U37878 ( .A(n38049), .B(n37992), .Z(n37980) );
  XOR U37879 ( .A(n37966), .B(n37965), .Z(n37992) );
  XNOR U37880 ( .A(n38050), .B(n37971), .Z(n37965) );
  XOR U37881 ( .A(p_input[2072]), .B(p_input[888]), .Z(n37971) );
  XOR U37882 ( .A(n37962), .B(n37970), .Z(n38050) );
  XOR U37883 ( .A(n38051), .B(n37967), .Z(n37970) );
  XOR U37884 ( .A(p_input[2070]), .B(p_input[886]), .Z(n37967) );
  XNOR U37885 ( .A(p_input[2071]), .B(p_input[887]), .Z(n38051) );
  XNOR U37886 ( .A(n28684), .B(p_input[882]), .Z(n37962) );
  XNOR U37887 ( .A(n37976), .B(n37975), .Z(n37966) );
  XOR U37888 ( .A(n38052), .B(n37972), .Z(n37975) );
  XOR U37889 ( .A(p_input[2067]), .B(p_input[883]), .Z(n37972) );
  XNOR U37890 ( .A(p_input[2068]), .B(p_input[884]), .Z(n38052) );
  XOR U37891 ( .A(p_input[2069]), .B(p_input[885]), .Z(n37976) );
  XNOR U37892 ( .A(n37991), .B(n37977), .Z(n38049) );
  XNOR U37893 ( .A(n28686), .B(p_input[865]), .Z(n37977) );
  XNOR U37894 ( .A(n38053), .B(n37998), .Z(n37991) );
  XNOR U37895 ( .A(n37987), .B(n37986), .Z(n37998) );
  XOR U37896 ( .A(n38054), .B(n37983), .Z(n37986) );
  XNOR U37897 ( .A(n28322), .B(p_input[890]), .Z(n37983) );
  XNOR U37898 ( .A(p_input[2075]), .B(p_input[891]), .Z(n38054) );
  XOR U37899 ( .A(p_input[2076]), .B(p_input[892]), .Z(n37987) );
  XNOR U37900 ( .A(n37997), .B(n37988), .Z(n38053) );
  XNOR U37901 ( .A(n28689), .B(p_input[881]), .Z(n37988) );
  XOR U37902 ( .A(n38055), .B(n38003), .Z(n37997) );
  XNOR U37903 ( .A(p_input[2079]), .B(p_input[895]), .Z(n38003) );
  XOR U37904 ( .A(n37994), .B(n38002), .Z(n38055) );
  XOR U37905 ( .A(n38056), .B(n37999), .Z(n38002) );
  XOR U37906 ( .A(p_input[2077]), .B(p_input[893]), .Z(n37999) );
  XNOR U37907 ( .A(p_input[2078]), .B(p_input[894]), .Z(n38056) );
  XNOR U37908 ( .A(n28326), .B(p_input[889]), .Z(n37994) );
  XNOR U37909 ( .A(n38015), .B(n38014), .Z(n37981) );
  XNOR U37910 ( .A(n38057), .B(n38021), .Z(n38014) );
  XNOR U37911 ( .A(n38010), .B(n38009), .Z(n38021) );
  XOR U37912 ( .A(n38058), .B(n38006), .Z(n38009) );
  XNOR U37913 ( .A(n28694), .B(p_input[875]), .Z(n38006) );
  XNOR U37914 ( .A(p_input[2060]), .B(p_input[876]), .Z(n38058) );
  XOR U37915 ( .A(p_input[2061]), .B(p_input[877]), .Z(n38010) );
  XNOR U37916 ( .A(n38020), .B(n38011), .Z(n38057) );
  XNOR U37917 ( .A(n28330), .B(p_input[866]), .Z(n38011) );
  XOR U37918 ( .A(n38059), .B(n38026), .Z(n38020) );
  XNOR U37919 ( .A(p_input[2064]), .B(p_input[880]), .Z(n38026) );
  XOR U37920 ( .A(n38017), .B(n38025), .Z(n38059) );
  XOR U37921 ( .A(n38060), .B(n38022), .Z(n38025) );
  XOR U37922 ( .A(p_input[2062]), .B(p_input[878]), .Z(n38022) );
  XNOR U37923 ( .A(p_input[2063]), .B(p_input[879]), .Z(n38060) );
  XNOR U37924 ( .A(n28697), .B(p_input[874]), .Z(n38017) );
  XNOR U37925 ( .A(n38032), .B(n38031), .Z(n38015) );
  XNOR U37926 ( .A(n38061), .B(n38037), .Z(n38031) );
  XOR U37927 ( .A(p_input[2057]), .B(p_input[873]), .Z(n38037) );
  XOR U37928 ( .A(n38028), .B(n38036), .Z(n38061) );
  XOR U37929 ( .A(n38062), .B(n38033), .Z(n38036) );
  XOR U37930 ( .A(p_input[2055]), .B(p_input[871]), .Z(n38033) );
  XNOR U37931 ( .A(p_input[2056]), .B(p_input[872]), .Z(n38062) );
  XNOR U37932 ( .A(n28337), .B(p_input[867]), .Z(n38028) );
  XNOR U37933 ( .A(n38042), .B(n38041), .Z(n38032) );
  XOR U37934 ( .A(n38063), .B(n38038), .Z(n38041) );
  XOR U37935 ( .A(p_input[2052]), .B(p_input[868]), .Z(n38038) );
  XNOR U37936 ( .A(p_input[2053]), .B(p_input[869]), .Z(n38063) );
  XOR U37937 ( .A(p_input[2054]), .B(p_input[870]), .Z(n38042) );
  XNOR U37938 ( .A(n38064), .B(n38065), .Z(n37847) );
  AND U37939 ( .A(n648), .B(n38066), .Z(n38065) );
  XNOR U37940 ( .A(n38067), .B(n38068), .Z(n648) );
  AND U37941 ( .A(n38069), .B(n38070), .Z(n38068) );
  XOR U37942 ( .A(n37861), .B(n38067), .Z(n38070) );
  XNOR U37943 ( .A(n38071), .B(n38067), .Z(n38069) );
  XOR U37944 ( .A(n38072), .B(n38073), .Z(n38067) );
  AND U37945 ( .A(n38074), .B(n38075), .Z(n38073) );
  XOR U37946 ( .A(n37876), .B(n38072), .Z(n38075) );
  XOR U37947 ( .A(n38072), .B(n37877), .Z(n38074) );
  XOR U37948 ( .A(n38076), .B(n38077), .Z(n38072) );
  AND U37949 ( .A(n38078), .B(n38079), .Z(n38077) );
  XOR U37950 ( .A(n37904), .B(n38076), .Z(n38079) );
  XOR U37951 ( .A(n38076), .B(n37905), .Z(n38078) );
  XOR U37952 ( .A(n38080), .B(n38081), .Z(n38076) );
  AND U37953 ( .A(n38082), .B(n38083), .Z(n38081) );
  XOR U37954 ( .A(n37953), .B(n38080), .Z(n38083) );
  XOR U37955 ( .A(n38080), .B(n37954), .Z(n38082) );
  XOR U37956 ( .A(n38084), .B(n38085), .Z(n38080) );
  AND U37957 ( .A(n38086), .B(n38087), .Z(n38085) );
  XOR U37958 ( .A(n38084), .B(n38046), .Z(n38087) );
  XNOR U37959 ( .A(n38088), .B(n38089), .Z(n37797) );
  AND U37960 ( .A(n652), .B(n38090), .Z(n38089) );
  XNOR U37961 ( .A(n38091), .B(n38092), .Z(n652) );
  AND U37962 ( .A(n38093), .B(n38094), .Z(n38092) );
  XOR U37963 ( .A(n38091), .B(n37807), .Z(n38094) );
  XNOR U37964 ( .A(n38091), .B(n37757), .Z(n38093) );
  XOR U37965 ( .A(n38095), .B(n38096), .Z(n38091) );
  AND U37966 ( .A(n38097), .B(n38098), .Z(n38096) );
  XNOR U37967 ( .A(n37817), .B(n38095), .Z(n38098) );
  XOR U37968 ( .A(n38095), .B(n37767), .Z(n38097) );
  XOR U37969 ( .A(n38099), .B(n38100), .Z(n38095) );
  AND U37970 ( .A(n38101), .B(n38102), .Z(n38100) );
  XNOR U37971 ( .A(n37827), .B(n38099), .Z(n38102) );
  XOR U37972 ( .A(n38099), .B(n37776), .Z(n38101) );
  XOR U37973 ( .A(n38103), .B(n38104), .Z(n38099) );
  AND U37974 ( .A(n38105), .B(n38106), .Z(n38104) );
  XOR U37975 ( .A(n38103), .B(n37784), .Z(n38105) );
  XOR U37976 ( .A(n38107), .B(n38108), .Z(n37748) );
  AND U37977 ( .A(n656), .B(n38090), .Z(n38108) );
  XNOR U37978 ( .A(n38088), .B(n38107), .Z(n38090) );
  XNOR U37979 ( .A(n38109), .B(n38110), .Z(n656) );
  AND U37980 ( .A(n38111), .B(n38112), .Z(n38110) );
  XNOR U37981 ( .A(n38113), .B(n38109), .Z(n38112) );
  IV U37982 ( .A(n37807), .Z(n38113) );
  XOR U37983 ( .A(n38071), .B(n38114), .Z(n37807) );
  AND U37984 ( .A(n659), .B(n38115), .Z(n38114) );
  XOR U37985 ( .A(n37860), .B(n37857), .Z(n38115) );
  IV U37986 ( .A(n38071), .Z(n37860) );
  XNOR U37987 ( .A(n37757), .B(n38109), .Z(n38111) );
  XOR U37988 ( .A(n38116), .B(n38117), .Z(n37757) );
  AND U37989 ( .A(n675), .B(n38118), .Z(n38117) );
  XOR U37990 ( .A(n38119), .B(n38120), .Z(n38109) );
  AND U37991 ( .A(n38121), .B(n38122), .Z(n38120) );
  XNOR U37992 ( .A(n38119), .B(n37817), .Z(n38122) );
  XOR U37993 ( .A(n37877), .B(n38123), .Z(n37817) );
  AND U37994 ( .A(n659), .B(n38124), .Z(n38123) );
  XOR U37995 ( .A(n37873), .B(n37877), .Z(n38124) );
  XNOR U37996 ( .A(n38125), .B(n38119), .Z(n38121) );
  IV U37997 ( .A(n37767), .Z(n38125) );
  XOR U37998 ( .A(n38126), .B(n38127), .Z(n37767) );
  AND U37999 ( .A(n675), .B(n38128), .Z(n38127) );
  XOR U38000 ( .A(n38129), .B(n38130), .Z(n38119) );
  AND U38001 ( .A(n38131), .B(n38132), .Z(n38130) );
  XNOR U38002 ( .A(n38129), .B(n37827), .Z(n38132) );
  XOR U38003 ( .A(n37905), .B(n38133), .Z(n37827) );
  AND U38004 ( .A(n659), .B(n38134), .Z(n38133) );
  XOR U38005 ( .A(n37901), .B(n37905), .Z(n38134) );
  XOR U38006 ( .A(n37776), .B(n38129), .Z(n38131) );
  XOR U38007 ( .A(n38135), .B(n38136), .Z(n37776) );
  AND U38008 ( .A(n675), .B(n38137), .Z(n38136) );
  XOR U38009 ( .A(n38103), .B(n38138), .Z(n38129) );
  AND U38010 ( .A(n38139), .B(n38106), .Z(n38138) );
  XNOR U38011 ( .A(n37837), .B(n38103), .Z(n38106) );
  XOR U38012 ( .A(n37954), .B(n38140), .Z(n37837) );
  AND U38013 ( .A(n659), .B(n38141), .Z(n38140) );
  XOR U38014 ( .A(n37950), .B(n37954), .Z(n38141) );
  XNOR U38015 ( .A(n38142), .B(n38103), .Z(n38139) );
  IV U38016 ( .A(n37784), .Z(n38142) );
  XOR U38017 ( .A(n38143), .B(n38144), .Z(n37784) );
  AND U38018 ( .A(n675), .B(n38145), .Z(n38144) );
  XOR U38019 ( .A(n38146), .B(n38147), .Z(n38103) );
  AND U38020 ( .A(n38148), .B(n38149), .Z(n38147) );
  XNOR U38021 ( .A(n38146), .B(n37845), .Z(n38149) );
  XOR U38022 ( .A(n38047), .B(n38150), .Z(n37845) );
  AND U38023 ( .A(n659), .B(n38151), .Z(n38150) );
  XOR U38024 ( .A(n38043), .B(n38047), .Z(n38151) );
  XNOR U38025 ( .A(n38152), .B(n38146), .Z(n38148) );
  IV U38026 ( .A(n37794), .Z(n38152) );
  XOR U38027 ( .A(n38153), .B(n38154), .Z(n37794) );
  AND U38028 ( .A(n675), .B(n38155), .Z(n38154) );
  AND U38029 ( .A(n38107), .B(n38088), .Z(n38146) );
  XNOR U38030 ( .A(n38156), .B(n38157), .Z(n38088) );
  AND U38031 ( .A(n659), .B(n38066), .Z(n38157) );
  XNOR U38032 ( .A(n38064), .B(n38156), .Z(n38066) );
  XNOR U38033 ( .A(n38158), .B(n38159), .Z(n659) );
  AND U38034 ( .A(n38160), .B(n38161), .Z(n38159) );
  XNOR U38035 ( .A(n38158), .B(n37857), .Z(n38161) );
  IV U38036 ( .A(n37861), .Z(n37857) );
  XOR U38037 ( .A(n38162), .B(n38163), .Z(n37861) );
  AND U38038 ( .A(n663), .B(n38164), .Z(n38163) );
  XOR U38039 ( .A(n38165), .B(n38162), .Z(n38164) );
  XNOR U38040 ( .A(n38158), .B(n38071), .Z(n38160) );
  XOR U38041 ( .A(n38166), .B(n38167), .Z(n38071) );
  AND U38042 ( .A(n671), .B(n38118), .Z(n38167) );
  XOR U38043 ( .A(n38116), .B(n38166), .Z(n38118) );
  XOR U38044 ( .A(n38168), .B(n38169), .Z(n38158) );
  AND U38045 ( .A(n38170), .B(n38171), .Z(n38169) );
  XNOR U38046 ( .A(n38168), .B(n37873), .Z(n38171) );
  IV U38047 ( .A(n37876), .Z(n37873) );
  XOR U38048 ( .A(n38172), .B(n38173), .Z(n37876) );
  AND U38049 ( .A(n663), .B(n38174), .Z(n38173) );
  XOR U38050 ( .A(n38175), .B(n38172), .Z(n38174) );
  XOR U38051 ( .A(n37877), .B(n38168), .Z(n38170) );
  XOR U38052 ( .A(n38176), .B(n38177), .Z(n37877) );
  AND U38053 ( .A(n671), .B(n38128), .Z(n38177) );
  XOR U38054 ( .A(n38176), .B(n38126), .Z(n38128) );
  XOR U38055 ( .A(n38178), .B(n38179), .Z(n38168) );
  AND U38056 ( .A(n38180), .B(n38181), .Z(n38179) );
  XNOR U38057 ( .A(n38178), .B(n37901), .Z(n38181) );
  IV U38058 ( .A(n37904), .Z(n37901) );
  XOR U38059 ( .A(n38182), .B(n38183), .Z(n37904) );
  AND U38060 ( .A(n663), .B(n38184), .Z(n38183) );
  XNOR U38061 ( .A(n38185), .B(n38182), .Z(n38184) );
  XOR U38062 ( .A(n37905), .B(n38178), .Z(n38180) );
  XOR U38063 ( .A(n38186), .B(n38187), .Z(n37905) );
  AND U38064 ( .A(n671), .B(n38137), .Z(n38187) );
  XOR U38065 ( .A(n38186), .B(n38135), .Z(n38137) );
  XOR U38066 ( .A(n38188), .B(n38189), .Z(n38178) );
  AND U38067 ( .A(n38190), .B(n38191), .Z(n38189) );
  XNOR U38068 ( .A(n38188), .B(n37950), .Z(n38191) );
  IV U38069 ( .A(n37953), .Z(n37950) );
  XOR U38070 ( .A(n38192), .B(n38193), .Z(n37953) );
  AND U38071 ( .A(n663), .B(n38194), .Z(n38193) );
  XOR U38072 ( .A(n38195), .B(n38192), .Z(n38194) );
  XOR U38073 ( .A(n37954), .B(n38188), .Z(n38190) );
  XOR U38074 ( .A(n38196), .B(n38197), .Z(n37954) );
  AND U38075 ( .A(n671), .B(n38145), .Z(n38197) );
  XOR U38076 ( .A(n38196), .B(n38143), .Z(n38145) );
  XOR U38077 ( .A(n38084), .B(n38198), .Z(n38188) );
  AND U38078 ( .A(n38086), .B(n38199), .Z(n38198) );
  XNOR U38079 ( .A(n38084), .B(n38043), .Z(n38199) );
  IV U38080 ( .A(n38046), .Z(n38043) );
  XOR U38081 ( .A(n38200), .B(n38201), .Z(n38046) );
  AND U38082 ( .A(n663), .B(n38202), .Z(n38201) );
  XNOR U38083 ( .A(n38203), .B(n38200), .Z(n38202) );
  XOR U38084 ( .A(n38047), .B(n38084), .Z(n38086) );
  XOR U38085 ( .A(n38204), .B(n38205), .Z(n38047) );
  AND U38086 ( .A(n671), .B(n38155), .Z(n38205) );
  XOR U38087 ( .A(n38204), .B(n38153), .Z(n38155) );
  AND U38088 ( .A(n38156), .B(n38064), .Z(n38084) );
  XNOR U38089 ( .A(n38206), .B(n38207), .Z(n38064) );
  AND U38090 ( .A(n663), .B(n38208), .Z(n38207) );
  XNOR U38091 ( .A(n38209), .B(n38206), .Z(n38208) );
  XNOR U38092 ( .A(n38210), .B(n38211), .Z(n663) );
  AND U38093 ( .A(n38212), .B(n38213), .Z(n38211) );
  XOR U38094 ( .A(n38165), .B(n38210), .Z(n38213) );
  AND U38095 ( .A(n38214), .B(n38215), .Z(n38165) );
  XNOR U38096 ( .A(n38162), .B(n38210), .Z(n38212) );
  XNOR U38097 ( .A(n38216), .B(n38217), .Z(n38162) );
  AND U38098 ( .A(n667), .B(n38218), .Z(n38217) );
  XNOR U38099 ( .A(n38219), .B(n38220), .Z(n38218) );
  XOR U38100 ( .A(n38221), .B(n38222), .Z(n38210) );
  AND U38101 ( .A(n38223), .B(n38224), .Z(n38222) );
  XNOR U38102 ( .A(n38221), .B(n38214), .Z(n38224) );
  IV U38103 ( .A(n38175), .Z(n38214) );
  XOR U38104 ( .A(n38225), .B(n38226), .Z(n38175) );
  XOR U38105 ( .A(n38227), .B(n38215), .Z(n38226) );
  AND U38106 ( .A(n38185), .B(n38228), .Z(n38215) );
  AND U38107 ( .A(n38229), .B(n38230), .Z(n38227) );
  XOR U38108 ( .A(n38231), .B(n38225), .Z(n38229) );
  XNOR U38109 ( .A(n38172), .B(n38221), .Z(n38223) );
  XNOR U38110 ( .A(n38232), .B(n38233), .Z(n38172) );
  AND U38111 ( .A(n667), .B(n38234), .Z(n38233) );
  XNOR U38112 ( .A(n38235), .B(n38236), .Z(n38234) );
  XOR U38113 ( .A(n38237), .B(n38238), .Z(n38221) );
  AND U38114 ( .A(n38239), .B(n38240), .Z(n38238) );
  XNOR U38115 ( .A(n38237), .B(n38185), .Z(n38240) );
  XOR U38116 ( .A(n38241), .B(n38230), .Z(n38185) );
  XNOR U38117 ( .A(n38242), .B(n38225), .Z(n38230) );
  XOR U38118 ( .A(n38243), .B(n38244), .Z(n38225) );
  AND U38119 ( .A(n38245), .B(n38246), .Z(n38244) );
  XOR U38120 ( .A(n38247), .B(n38243), .Z(n38245) );
  XNOR U38121 ( .A(n38248), .B(n38249), .Z(n38242) );
  AND U38122 ( .A(n38250), .B(n38251), .Z(n38249) );
  XOR U38123 ( .A(n38248), .B(n38252), .Z(n38250) );
  XNOR U38124 ( .A(n38231), .B(n38228), .Z(n38241) );
  AND U38125 ( .A(n38253), .B(n38254), .Z(n38228) );
  XOR U38126 ( .A(n38255), .B(n38256), .Z(n38231) );
  AND U38127 ( .A(n38257), .B(n38258), .Z(n38256) );
  XOR U38128 ( .A(n38255), .B(n38259), .Z(n38257) );
  XNOR U38129 ( .A(n38182), .B(n38237), .Z(n38239) );
  XNOR U38130 ( .A(n38260), .B(n38261), .Z(n38182) );
  AND U38131 ( .A(n667), .B(n38262), .Z(n38261) );
  XNOR U38132 ( .A(n38263), .B(n38264), .Z(n38262) );
  XOR U38133 ( .A(n38265), .B(n38266), .Z(n38237) );
  AND U38134 ( .A(n38267), .B(n38268), .Z(n38266) );
  XNOR U38135 ( .A(n38265), .B(n38253), .Z(n38268) );
  IV U38136 ( .A(n38195), .Z(n38253) );
  XNOR U38137 ( .A(n38269), .B(n38246), .Z(n38195) );
  XNOR U38138 ( .A(n38270), .B(n38252), .Z(n38246) );
  XOR U38139 ( .A(n38271), .B(n38272), .Z(n38252) );
  AND U38140 ( .A(n38273), .B(n38274), .Z(n38272) );
  XOR U38141 ( .A(n38271), .B(n38275), .Z(n38273) );
  XNOR U38142 ( .A(n38251), .B(n38243), .Z(n38270) );
  XOR U38143 ( .A(n38276), .B(n38277), .Z(n38243) );
  AND U38144 ( .A(n38278), .B(n38279), .Z(n38277) );
  XNOR U38145 ( .A(n38280), .B(n38276), .Z(n38278) );
  XNOR U38146 ( .A(n38281), .B(n38248), .Z(n38251) );
  XOR U38147 ( .A(n38282), .B(n38283), .Z(n38248) );
  AND U38148 ( .A(n38284), .B(n38285), .Z(n38283) );
  XOR U38149 ( .A(n38282), .B(n38286), .Z(n38284) );
  XNOR U38150 ( .A(n38287), .B(n38288), .Z(n38281) );
  AND U38151 ( .A(n38289), .B(n38290), .Z(n38288) );
  XNOR U38152 ( .A(n38287), .B(n38291), .Z(n38289) );
  XNOR U38153 ( .A(n38247), .B(n38254), .Z(n38269) );
  AND U38154 ( .A(n38203), .B(n38292), .Z(n38254) );
  XOR U38155 ( .A(n38259), .B(n38258), .Z(n38247) );
  XNOR U38156 ( .A(n38293), .B(n38255), .Z(n38258) );
  XOR U38157 ( .A(n38294), .B(n38295), .Z(n38255) );
  AND U38158 ( .A(n38296), .B(n38297), .Z(n38295) );
  XOR U38159 ( .A(n38294), .B(n38298), .Z(n38296) );
  XNOR U38160 ( .A(n38299), .B(n38300), .Z(n38293) );
  AND U38161 ( .A(n38301), .B(n38302), .Z(n38300) );
  XOR U38162 ( .A(n38299), .B(n38303), .Z(n38301) );
  XOR U38163 ( .A(n38304), .B(n38305), .Z(n38259) );
  AND U38164 ( .A(n38306), .B(n38307), .Z(n38305) );
  XOR U38165 ( .A(n38304), .B(n38308), .Z(n38306) );
  XNOR U38166 ( .A(n38192), .B(n38265), .Z(n38267) );
  XNOR U38167 ( .A(n38309), .B(n38310), .Z(n38192) );
  AND U38168 ( .A(n667), .B(n38311), .Z(n38310) );
  XNOR U38169 ( .A(n38312), .B(n38313), .Z(n38311) );
  XOR U38170 ( .A(n38314), .B(n38315), .Z(n38265) );
  AND U38171 ( .A(n38316), .B(n38317), .Z(n38315) );
  XNOR U38172 ( .A(n38314), .B(n38203), .Z(n38317) );
  XOR U38173 ( .A(n38318), .B(n38279), .Z(n38203) );
  XNOR U38174 ( .A(n38319), .B(n38286), .Z(n38279) );
  XOR U38175 ( .A(n38275), .B(n38274), .Z(n38286) );
  XNOR U38176 ( .A(n38320), .B(n38271), .Z(n38274) );
  XOR U38177 ( .A(n38321), .B(n38322), .Z(n38271) );
  AND U38178 ( .A(n38323), .B(n38324), .Z(n38322) );
  XOR U38179 ( .A(n38321), .B(n38325), .Z(n38323) );
  XNOR U38180 ( .A(n38326), .B(n38327), .Z(n38320) );
  NOR U38181 ( .A(n38328), .B(n38329), .Z(n38327) );
  XNOR U38182 ( .A(n38326), .B(n38330), .Z(n38328) );
  XOR U38183 ( .A(n38331), .B(n38332), .Z(n38275) );
  NOR U38184 ( .A(n38333), .B(n38334), .Z(n38332) );
  XNOR U38185 ( .A(n38331), .B(n38335), .Z(n38333) );
  XNOR U38186 ( .A(n38285), .B(n38276), .Z(n38319) );
  XOR U38187 ( .A(n38336), .B(n38337), .Z(n38276) );
  NOR U38188 ( .A(n38338), .B(n38339), .Z(n38337) );
  XNOR U38189 ( .A(n38336), .B(n38340), .Z(n38338) );
  XOR U38190 ( .A(n38341), .B(n38291), .Z(n38285) );
  XNOR U38191 ( .A(n38342), .B(n38343), .Z(n38291) );
  NOR U38192 ( .A(n38344), .B(n38345), .Z(n38343) );
  XNOR U38193 ( .A(n38342), .B(n38346), .Z(n38344) );
  XNOR U38194 ( .A(n38290), .B(n38282), .Z(n38341) );
  XOR U38195 ( .A(n38347), .B(n38348), .Z(n38282) );
  AND U38196 ( .A(n38349), .B(n38350), .Z(n38348) );
  XOR U38197 ( .A(n38347), .B(n38351), .Z(n38349) );
  XNOR U38198 ( .A(n38352), .B(n38287), .Z(n38290) );
  XOR U38199 ( .A(n38353), .B(n38354), .Z(n38287) );
  AND U38200 ( .A(n38355), .B(n38356), .Z(n38354) );
  XOR U38201 ( .A(n38353), .B(n38357), .Z(n38355) );
  XNOR U38202 ( .A(n38358), .B(n38359), .Z(n38352) );
  NOR U38203 ( .A(n38360), .B(n38361), .Z(n38359) );
  XOR U38204 ( .A(n38358), .B(n38362), .Z(n38360) );
  XOR U38205 ( .A(n38280), .B(n38292), .Z(n38318) );
  NOR U38206 ( .A(n38209), .B(n38363), .Z(n38292) );
  XNOR U38207 ( .A(n38298), .B(n38297), .Z(n38280) );
  XNOR U38208 ( .A(n38364), .B(n38303), .Z(n38297) );
  XOR U38209 ( .A(n38365), .B(n38366), .Z(n38303) );
  NOR U38210 ( .A(n38367), .B(n38368), .Z(n38366) );
  XNOR U38211 ( .A(n38365), .B(n38369), .Z(n38367) );
  XNOR U38212 ( .A(n38302), .B(n38294), .Z(n38364) );
  XOR U38213 ( .A(n38370), .B(n38371), .Z(n38294) );
  AND U38214 ( .A(n38372), .B(n38373), .Z(n38371) );
  XNOR U38215 ( .A(n38370), .B(n38374), .Z(n38372) );
  XNOR U38216 ( .A(n38375), .B(n38299), .Z(n38302) );
  XOR U38217 ( .A(n38376), .B(n38377), .Z(n38299) );
  AND U38218 ( .A(n38378), .B(n38379), .Z(n38377) );
  XOR U38219 ( .A(n38376), .B(n38380), .Z(n38378) );
  XNOR U38220 ( .A(n38381), .B(n38382), .Z(n38375) );
  NOR U38221 ( .A(n38383), .B(n38384), .Z(n38382) );
  XOR U38222 ( .A(n38381), .B(n38385), .Z(n38383) );
  XOR U38223 ( .A(n38308), .B(n38307), .Z(n38298) );
  XNOR U38224 ( .A(n38386), .B(n38304), .Z(n38307) );
  XOR U38225 ( .A(n38387), .B(n38388), .Z(n38304) );
  AND U38226 ( .A(n38389), .B(n38390), .Z(n38388) );
  XOR U38227 ( .A(n38387), .B(n38391), .Z(n38389) );
  XNOR U38228 ( .A(n38392), .B(n38393), .Z(n38386) );
  NOR U38229 ( .A(n38394), .B(n38395), .Z(n38393) );
  XNOR U38230 ( .A(n38392), .B(n38396), .Z(n38394) );
  XOR U38231 ( .A(n38397), .B(n38398), .Z(n38308) );
  NOR U38232 ( .A(n38399), .B(n38400), .Z(n38398) );
  XNOR U38233 ( .A(n38397), .B(n38401), .Z(n38399) );
  XNOR U38234 ( .A(n38200), .B(n38314), .Z(n38316) );
  XNOR U38235 ( .A(n38402), .B(n38403), .Z(n38200) );
  AND U38236 ( .A(n667), .B(n38404), .Z(n38403) );
  XNOR U38237 ( .A(n38405), .B(n38406), .Z(n38404) );
  AND U38238 ( .A(n38206), .B(n38209), .Z(n38314) );
  XOR U38239 ( .A(n38407), .B(n38363), .Z(n38209) );
  XNOR U38240 ( .A(p_input[2048]), .B(p_input[896]), .Z(n38363) );
  XOR U38241 ( .A(n38340), .B(n38339), .Z(n38407) );
  XOR U38242 ( .A(n38408), .B(n38351), .Z(n38339) );
  XOR U38243 ( .A(n38325), .B(n38324), .Z(n38351) );
  XNOR U38244 ( .A(n38409), .B(n38330), .Z(n38324) );
  XOR U38245 ( .A(p_input[2072]), .B(p_input[920]), .Z(n38330) );
  XOR U38246 ( .A(n38321), .B(n38329), .Z(n38409) );
  XOR U38247 ( .A(n38410), .B(n38326), .Z(n38329) );
  XOR U38248 ( .A(p_input[2070]), .B(p_input[918]), .Z(n38326) );
  XNOR U38249 ( .A(p_input[2071]), .B(p_input[919]), .Z(n38410) );
  XNOR U38250 ( .A(n28684), .B(p_input[914]), .Z(n38321) );
  XNOR U38251 ( .A(n38335), .B(n38334), .Z(n38325) );
  XOR U38252 ( .A(n38411), .B(n38331), .Z(n38334) );
  XOR U38253 ( .A(p_input[2067]), .B(p_input[915]), .Z(n38331) );
  XNOR U38254 ( .A(p_input[2068]), .B(p_input[916]), .Z(n38411) );
  XOR U38255 ( .A(p_input[2069]), .B(p_input[917]), .Z(n38335) );
  XNOR U38256 ( .A(n38350), .B(n38336), .Z(n38408) );
  XNOR U38257 ( .A(n28686), .B(p_input[897]), .Z(n38336) );
  XNOR U38258 ( .A(n38412), .B(n38357), .Z(n38350) );
  XNOR U38259 ( .A(n38346), .B(n38345), .Z(n38357) );
  XOR U38260 ( .A(n38413), .B(n38342), .Z(n38345) );
  XNOR U38261 ( .A(n28322), .B(p_input[922]), .Z(n38342) );
  XNOR U38262 ( .A(p_input[2075]), .B(p_input[923]), .Z(n38413) );
  XOR U38263 ( .A(p_input[2076]), .B(p_input[924]), .Z(n38346) );
  XNOR U38264 ( .A(n38356), .B(n38347), .Z(n38412) );
  XNOR U38265 ( .A(n28689), .B(p_input[913]), .Z(n38347) );
  XOR U38266 ( .A(n38414), .B(n38362), .Z(n38356) );
  XNOR U38267 ( .A(p_input[2079]), .B(p_input[927]), .Z(n38362) );
  XOR U38268 ( .A(n38353), .B(n38361), .Z(n38414) );
  XOR U38269 ( .A(n38415), .B(n38358), .Z(n38361) );
  XOR U38270 ( .A(p_input[2077]), .B(p_input[925]), .Z(n38358) );
  XNOR U38271 ( .A(p_input[2078]), .B(p_input[926]), .Z(n38415) );
  XNOR U38272 ( .A(n28326), .B(p_input[921]), .Z(n38353) );
  XNOR U38273 ( .A(n38374), .B(n38373), .Z(n38340) );
  XNOR U38274 ( .A(n38416), .B(n38380), .Z(n38373) );
  XNOR U38275 ( .A(n38369), .B(n38368), .Z(n38380) );
  XOR U38276 ( .A(n38417), .B(n38365), .Z(n38368) );
  XNOR U38277 ( .A(n28694), .B(p_input[907]), .Z(n38365) );
  XNOR U38278 ( .A(p_input[2060]), .B(p_input[908]), .Z(n38417) );
  XOR U38279 ( .A(p_input[2061]), .B(p_input[909]), .Z(n38369) );
  XNOR U38280 ( .A(n38379), .B(n38370), .Z(n38416) );
  XNOR U38281 ( .A(n28330), .B(p_input[898]), .Z(n38370) );
  XOR U38282 ( .A(n38418), .B(n38385), .Z(n38379) );
  XNOR U38283 ( .A(p_input[2064]), .B(p_input[912]), .Z(n38385) );
  XOR U38284 ( .A(n38376), .B(n38384), .Z(n38418) );
  XOR U38285 ( .A(n38419), .B(n38381), .Z(n38384) );
  XOR U38286 ( .A(p_input[2062]), .B(p_input[910]), .Z(n38381) );
  XNOR U38287 ( .A(p_input[2063]), .B(p_input[911]), .Z(n38419) );
  XNOR U38288 ( .A(n28697), .B(p_input[906]), .Z(n38376) );
  XNOR U38289 ( .A(n38391), .B(n38390), .Z(n38374) );
  XNOR U38290 ( .A(n38420), .B(n38396), .Z(n38390) );
  XOR U38291 ( .A(p_input[2057]), .B(p_input[905]), .Z(n38396) );
  XOR U38292 ( .A(n38387), .B(n38395), .Z(n38420) );
  XOR U38293 ( .A(n38421), .B(n38392), .Z(n38395) );
  XOR U38294 ( .A(p_input[2055]), .B(p_input[903]), .Z(n38392) );
  XNOR U38295 ( .A(p_input[2056]), .B(p_input[904]), .Z(n38421) );
  XNOR U38296 ( .A(n28337), .B(p_input[899]), .Z(n38387) );
  XNOR U38297 ( .A(n38401), .B(n38400), .Z(n38391) );
  XOR U38298 ( .A(n38422), .B(n38397), .Z(n38400) );
  XOR U38299 ( .A(p_input[2052]), .B(p_input[900]), .Z(n38397) );
  XNOR U38300 ( .A(p_input[2053]), .B(p_input[901]), .Z(n38422) );
  XOR U38301 ( .A(p_input[2054]), .B(p_input[902]), .Z(n38401) );
  XNOR U38302 ( .A(n38423), .B(n38424), .Z(n38206) );
  AND U38303 ( .A(n667), .B(n38425), .Z(n38424) );
  XNOR U38304 ( .A(n38426), .B(n38427), .Z(n667) );
  AND U38305 ( .A(n38428), .B(n38429), .Z(n38427) );
  XOR U38306 ( .A(n38220), .B(n38426), .Z(n38429) );
  XNOR U38307 ( .A(n38430), .B(n38426), .Z(n38428) );
  XOR U38308 ( .A(n38431), .B(n38432), .Z(n38426) );
  AND U38309 ( .A(n38433), .B(n38434), .Z(n38432) );
  XOR U38310 ( .A(n38235), .B(n38431), .Z(n38434) );
  XOR U38311 ( .A(n38431), .B(n38236), .Z(n38433) );
  XOR U38312 ( .A(n38435), .B(n38436), .Z(n38431) );
  AND U38313 ( .A(n38437), .B(n38438), .Z(n38436) );
  XOR U38314 ( .A(n38263), .B(n38435), .Z(n38438) );
  XOR U38315 ( .A(n38435), .B(n38264), .Z(n38437) );
  XOR U38316 ( .A(n38439), .B(n38440), .Z(n38435) );
  AND U38317 ( .A(n38441), .B(n38442), .Z(n38440) );
  XOR U38318 ( .A(n38312), .B(n38439), .Z(n38442) );
  XOR U38319 ( .A(n38439), .B(n38313), .Z(n38441) );
  XOR U38320 ( .A(n38443), .B(n38444), .Z(n38439) );
  AND U38321 ( .A(n38445), .B(n38446), .Z(n38444) );
  XOR U38322 ( .A(n38443), .B(n38405), .Z(n38446) );
  XNOR U38323 ( .A(n38447), .B(n38448), .Z(n38156) );
  AND U38324 ( .A(n671), .B(n38449), .Z(n38448) );
  XNOR U38325 ( .A(n38450), .B(n38451), .Z(n671) );
  AND U38326 ( .A(n38452), .B(n38453), .Z(n38451) );
  XOR U38327 ( .A(n38450), .B(n38166), .Z(n38453) );
  XNOR U38328 ( .A(n38450), .B(n38116), .Z(n38452) );
  XOR U38329 ( .A(n38454), .B(n38455), .Z(n38450) );
  AND U38330 ( .A(n38456), .B(n38457), .Z(n38455) );
  XNOR U38331 ( .A(n38176), .B(n38454), .Z(n38457) );
  XOR U38332 ( .A(n38454), .B(n38126), .Z(n38456) );
  XOR U38333 ( .A(n38458), .B(n38459), .Z(n38454) );
  AND U38334 ( .A(n38460), .B(n38461), .Z(n38459) );
  XNOR U38335 ( .A(n38186), .B(n38458), .Z(n38461) );
  XOR U38336 ( .A(n38458), .B(n38135), .Z(n38460) );
  XOR U38337 ( .A(n38462), .B(n38463), .Z(n38458) );
  AND U38338 ( .A(n38464), .B(n38465), .Z(n38463) );
  XOR U38339 ( .A(n38462), .B(n38143), .Z(n38464) );
  XOR U38340 ( .A(n38466), .B(n38467), .Z(n38107) );
  AND U38341 ( .A(n675), .B(n38449), .Z(n38467) );
  XNOR U38342 ( .A(n38447), .B(n38466), .Z(n38449) );
  XNOR U38343 ( .A(n38468), .B(n38469), .Z(n675) );
  AND U38344 ( .A(n38470), .B(n38471), .Z(n38469) );
  XNOR U38345 ( .A(n38472), .B(n38468), .Z(n38471) );
  IV U38346 ( .A(n38166), .Z(n38472) );
  XOR U38347 ( .A(n38430), .B(n38473), .Z(n38166) );
  AND U38348 ( .A(n678), .B(n38474), .Z(n38473) );
  XOR U38349 ( .A(n38219), .B(n38216), .Z(n38474) );
  IV U38350 ( .A(n38430), .Z(n38219) );
  XNOR U38351 ( .A(n38116), .B(n38468), .Z(n38470) );
  XOR U38352 ( .A(n38475), .B(n38476), .Z(n38116) );
  AND U38353 ( .A(n694), .B(n38477), .Z(n38476) );
  XOR U38354 ( .A(n38478), .B(n38479), .Z(n38468) );
  AND U38355 ( .A(n38480), .B(n38481), .Z(n38479) );
  XNOR U38356 ( .A(n38478), .B(n38176), .Z(n38481) );
  XOR U38357 ( .A(n38236), .B(n38482), .Z(n38176) );
  AND U38358 ( .A(n678), .B(n38483), .Z(n38482) );
  XOR U38359 ( .A(n38232), .B(n38236), .Z(n38483) );
  XNOR U38360 ( .A(n38484), .B(n38478), .Z(n38480) );
  IV U38361 ( .A(n38126), .Z(n38484) );
  XOR U38362 ( .A(n38485), .B(n38486), .Z(n38126) );
  AND U38363 ( .A(n694), .B(n38487), .Z(n38486) );
  XOR U38364 ( .A(n38488), .B(n38489), .Z(n38478) );
  AND U38365 ( .A(n38490), .B(n38491), .Z(n38489) );
  XNOR U38366 ( .A(n38488), .B(n38186), .Z(n38491) );
  XOR U38367 ( .A(n38264), .B(n38492), .Z(n38186) );
  AND U38368 ( .A(n678), .B(n38493), .Z(n38492) );
  XOR U38369 ( .A(n38260), .B(n38264), .Z(n38493) );
  XOR U38370 ( .A(n38135), .B(n38488), .Z(n38490) );
  XOR U38371 ( .A(n38494), .B(n38495), .Z(n38135) );
  AND U38372 ( .A(n694), .B(n38496), .Z(n38495) );
  XOR U38373 ( .A(n38462), .B(n38497), .Z(n38488) );
  AND U38374 ( .A(n38498), .B(n38465), .Z(n38497) );
  XNOR U38375 ( .A(n38196), .B(n38462), .Z(n38465) );
  XOR U38376 ( .A(n38313), .B(n38499), .Z(n38196) );
  AND U38377 ( .A(n678), .B(n38500), .Z(n38499) );
  XOR U38378 ( .A(n38309), .B(n38313), .Z(n38500) );
  XNOR U38379 ( .A(n38501), .B(n38462), .Z(n38498) );
  IV U38380 ( .A(n38143), .Z(n38501) );
  XOR U38381 ( .A(n38502), .B(n38503), .Z(n38143) );
  AND U38382 ( .A(n694), .B(n38504), .Z(n38503) );
  XOR U38383 ( .A(n38505), .B(n38506), .Z(n38462) );
  AND U38384 ( .A(n38507), .B(n38508), .Z(n38506) );
  XNOR U38385 ( .A(n38505), .B(n38204), .Z(n38508) );
  XOR U38386 ( .A(n38406), .B(n38509), .Z(n38204) );
  AND U38387 ( .A(n678), .B(n38510), .Z(n38509) );
  XOR U38388 ( .A(n38402), .B(n38406), .Z(n38510) );
  XNOR U38389 ( .A(n38511), .B(n38505), .Z(n38507) );
  IV U38390 ( .A(n38153), .Z(n38511) );
  XOR U38391 ( .A(n38512), .B(n38513), .Z(n38153) );
  AND U38392 ( .A(n694), .B(n38514), .Z(n38513) );
  AND U38393 ( .A(n38466), .B(n38447), .Z(n38505) );
  XNOR U38394 ( .A(n38515), .B(n38516), .Z(n38447) );
  AND U38395 ( .A(n678), .B(n38425), .Z(n38516) );
  XNOR U38396 ( .A(n38423), .B(n38515), .Z(n38425) );
  XNOR U38397 ( .A(n38517), .B(n38518), .Z(n678) );
  AND U38398 ( .A(n38519), .B(n38520), .Z(n38518) );
  XNOR U38399 ( .A(n38517), .B(n38216), .Z(n38520) );
  IV U38400 ( .A(n38220), .Z(n38216) );
  XOR U38401 ( .A(n38521), .B(n38522), .Z(n38220) );
  AND U38402 ( .A(n682), .B(n38523), .Z(n38522) );
  XOR U38403 ( .A(n38524), .B(n38521), .Z(n38523) );
  XNOR U38404 ( .A(n38517), .B(n38430), .Z(n38519) );
  XOR U38405 ( .A(n38525), .B(n38526), .Z(n38430) );
  AND U38406 ( .A(n690), .B(n38477), .Z(n38526) );
  XOR U38407 ( .A(n38475), .B(n38525), .Z(n38477) );
  XOR U38408 ( .A(n38527), .B(n38528), .Z(n38517) );
  AND U38409 ( .A(n38529), .B(n38530), .Z(n38528) );
  XNOR U38410 ( .A(n38527), .B(n38232), .Z(n38530) );
  IV U38411 ( .A(n38235), .Z(n38232) );
  XOR U38412 ( .A(n38531), .B(n38532), .Z(n38235) );
  AND U38413 ( .A(n682), .B(n38533), .Z(n38532) );
  XOR U38414 ( .A(n38534), .B(n38531), .Z(n38533) );
  XOR U38415 ( .A(n38236), .B(n38527), .Z(n38529) );
  XOR U38416 ( .A(n38535), .B(n38536), .Z(n38236) );
  AND U38417 ( .A(n690), .B(n38487), .Z(n38536) );
  XOR U38418 ( .A(n38535), .B(n38485), .Z(n38487) );
  XOR U38419 ( .A(n38537), .B(n38538), .Z(n38527) );
  AND U38420 ( .A(n38539), .B(n38540), .Z(n38538) );
  XNOR U38421 ( .A(n38537), .B(n38260), .Z(n38540) );
  IV U38422 ( .A(n38263), .Z(n38260) );
  XOR U38423 ( .A(n38541), .B(n38542), .Z(n38263) );
  AND U38424 ( .A(n682), .B(n38543), .Z(n38542) );
  XNOR U38425 ( .A(n38544), .B(n38541), .Z(n38543) );
  XOR U38426 ( .A(n38264), .B(n38537), .Z(n38539) );
  XOR U38427 ( .A(n38545), .B(n38546), .Z(n38264) );
  AND U38428 ( .A(n690), .B(n38496), .Z(n38546) );
  XOR U38429 ( .A(n38545), .B(n38494), .Z(n38496) );
  XOR U38430 ( .A(n38547), .B(n38548), .Z(n38537) );
  AND U38431 ( .A(n38549), .B(n38550), .Z(n38548) );
  XNOR U38432 ( .A(n38547), .B(n38309), .Z(n38550) );
  IV U38433 ( .A(n38312), .Z(n38309) );
  XOR U38434 ( .A(n38551), .B(n38552), .Z(n38312) );
  AND U38435 ( .A(n682), .B(n38553), .Z(n38552) );
  XOR U38436 ( .A(n38554), .B(n38551), .Z(n38553) );
  XOR U38437 ( .A(n38313), .B(n38547), .Z(n38549) );
  XOR U38438 ( .A(n38555), .B(n38556), .Z(n38313) );
  AND U38439 ( .A(n690), .B(n38504), .Z(n38556) );
  XOR U38440 ( .A(n38555), .B(n38502), .Z(n38504) );
  XOR U38441 ( .A(n38443), .B(n38557), .Z(n38547) );
  AND U38442 ( .A(n38445), .B(n38558), .Z(n38557) );
  XNOR U38443 ( .A(n38443), .B(n38402), .Z(n38558) );
  IV U38444 ( .A(n38405), .Z(n38402) );
  XOR U38445 ( .A(n38559), .B(n38560), .Z(n38405) );
  AND U38446 ( .A(n682), .B(n38561), .Z(n38560) );
  XNOR U38447 ( .A(n38562), .B(n38559), .Z(n38561) );
  XOR U38448 ( .A(n38406), .B(n38443), .Z(n38445) );
  XOR U38449 ( .A(n38563), .B(n38564), .Z(n38406) );
  AND U38450 ( .A(n690), .B(n38514), .Z(n38564) );
  XOR U38451 ( .A(n38563), .B(n38512), .Z(n38514) );
  AND U38452 ( .A(n38515), .B(n38423), .Z(n38443) );
  XNOR U38453 ( .A(n38565), .B(n38566), .Z(n38423) );
  AND U38454 ( .A(n682), .B(n38567), .Z(n38566) );
  XNOR U38455 ( .A(n38568), .B(n38565), .Z(n38567) );
  XNOR U38456 ( .A(n38569), .B(n38570), .Z(n682) );
  AND U38457 ( .A(n38571), .B(n38572), .Z(n38570) );
  XOR U38458 ( .A(n38524), .B(n38569), .Z(n38572) );
  AND U38459 ( .A(n38573), .B(n38574), .Z(n38524) );
  XNOR U38460 ( .A(n38521), .B(n38569), .Z(n38571) );
  XNOR U38461 ( .A(n38575), .B(n38576), .Z(n38521) );
  AND U38462 ( .A(n686), .B(n38577), .Z(n38576) );
  XNOR U38463 ( .A(n38578), .B(n38579), .Z(n38577) );
  XOR U38464 ( .A(n38580), .B(n38581), .Z(n38569) );
  AND U38465 ( .A(n38582), .B(n38583), .Z(n38581) );
  XNOR U38466 ( .A(n38580), .B(n38573), .Z(n38583) );
  IV U38467 ( .A(n38534), .Z(n38573) );
  XOR U38468 ( .A(n38584), .B(n38585), .Z(n38534) );
  XOR U38469 ( .A(n38586), .B(n38574), .Z(n38585) );
  AND U38470 ( .A(n38544), .B(n38587), .Z(n38574) );
  AND U38471 ( .A(n38588), .B(n38589), .Z(n38586) );
  XOR U38472 ( .A(n38590), .B(n38584), .Z(n38588) );
  XNOR U38473 ( .A(n38531), .B(n38580), .Z(n38582) );
  XNOR U38474 ( .A(n38591), .B(n38592), .Z(n38531) );
  AND U38475 ( .A(n686), .B(n38593), .Z(n38592) );
  XNOR U38476 ( .A(n38594), .B(n38595), .Z(n38593) );
  XOR U38477 ( .A(n38596), .B(n38597), .Z(n38580) );
  AND U38478 ( .A(n38598), .B(n38599), .Z(n38597) );
  XNOR U38479 ( .A(n38596), .B(n38544), .Z(n38599) );
  XOR U38480 ( .A(n38600), .B(n38589), .Z(n38544) );
  XNOR U38481 ( .A(n38601), .B(n38584), .Z(n38589) );
  XOR U38482 ( .A(n38602), .B(n38603), .Z(n38584) );
  AND U38483 ( .A(n38604), .B(n38605), .Z(n38603) );
  XOR U38484 ( .A(n38606), .B(n38602), .Z(n38604) );
  XNOR U38485 ( .A(n38607), .B(n38608), .Z(n38601) );
  AND U38486 ( .A(n38609), .B(n38610), .Z(n38608) );
  XOR U38487 ( .A(n38607), .B(n38611), .Z(n38609) );
  XNOR U38488 ( .A(n38590), .B(n38587), .Z(n38600) );
  AND U38489 ( .A(n38612), .B(n38613), .Z(n38587) );
  XOR U38490 ( .A(n38614), .B(n38615), .Z(n38590) );
  AND U38491 ( .A(n38616), .B(n38617), .Z(n38615) );
  XOR U38492 ( .A(n38614), .B(n38618), .Z(n38616) );
  XNOR U38493 ( .A(n38541), .B(n38596), .Z(n38598) );
  XNOR U38494 ( .A(n38619), .B(n38620), .Z(n38541) );
  AND U38495 ( .A(n686), .B(n38621), .Z(n38620) );
  XNOR U38496 ( .A(n38622), .B(n38623), .Z(n38621) );
  XOR U38497 ( .A(n38624), .B(n38625), .Z(n38596) );
  AND U38498 ( .A(n38626), .B(n38627), .Z(n38625) );
  XNOR U38499 ( .A(n38624), .B(n38612), .Z(n38627) );
  IV U38500 ( .A(n38554), .Z(n38612) );
  XNOR U38501 ( .A(n38628), .B(n38605), .Z(n38554) );
  XNOR U38502 ( .A(n38629), .B(n38611), .Z(n38605) );
  XOR U38503 ( .A(n38630), .B(n38631), .Z(n38611) );
  AND U38504 ( .A(n38632), .B(n38633), .Z(n38631) );
  XOR U38505 ( .A(n38630), .B(n38634), .Z(n38632) );
  XNOR U38506 ( .A(n38610), .B(n38602), .Z(n38629) );
  XOR U38507 ( .A(n38635), .B(n38636), .Z(n38602) );
  AND U38508 ( .A(n38637), .B(n38638), .Z(n38636) );
  XNOR U38509 ( .A(n38639), .B(n38635), .Z(n38637) );
  XNOR U38510 ( .A(n38640), .B(n38607), .Z(n38610) );
  XOR U38511 ( .A(n38641), .B(n38642), .Z(n38607) );
  AND U38512 ( .A(n38643), .B(n38644), .Z(n38642) );
  XOR U38513 ( .A(n38641), .B(n38645), .Z(n38643) );
  XNOR U38514 ( .A(n38646), .B(n38647), .Z(n38640) );
  AND U38515 ( .A(n38648), .B(n38649), .Z(n38647) );
  XNOR U38516 ( .A(n38646), .B(n38650), .Z(n38648) );
  XNOR U38517 ( .A(n38606), .B(n38613), .Z(n38628) );
  AND U38518 ( .A(n38562), .B(n38651), .Z(n38613) );
  XOR U38519 ( .A(n38618), .B(n38617), .Z(n38606) );
  XNOR U38520 ( .A(n38652), .B(n38614), .Z(n38617) );
  XOR U38521 ( .A(n38653), .B(n38654), .Z(n38614) );
  AND U38522 ( .A(n38655), .B(n38656), .Z(n38654) );
  XOR U38523 ( .A(n38653), .B(n38657), .Z(n38655) );
  XNOR U38524 ( .A(n38658), .B(n38659), .Z(n38652) );
  AND U38525 ( .A(n38660), .B(n38661), .Z(n38659) );
  XOR U38526 ( .A(n38658), .B(n38662), .Z(n38660) );
  XOR U38527 ( .A(n38663), .B(n38664), .Z(n38618) );
  AND U38528 ( .A(n38665), .B(n38666), .Z(n38664) );
  XOR U38529 ( .A(n38663), .B(n38667), .Z(n38665) );
  XNOR U38530 ( .A(n38551), .B(n38624), .Z(n38626) );
  XNOR U38531 ( .A(n38668), .B(n38669), .Z(n38551) );
  AND U38532 ( .A(n686), .B(n38670), .Z(n38669) );
  XNOR U38533 ( .A(n38671), .B(n38672), .Z(n38670) );
  XOR U38534 ( .A(n38673), .B(n38674), .Z(n38624) );
  AND U38535 ( .A(n38675), .B(n38676), .Z(n38674) );
  XNOR U38536 ( .A(n38673), .B(n38562), .Z(n38676) );
  XOR U38537 ( .A(n38677), .B(n38638), .Z(n38562) );
  XNOR U38538 ( .A(n38678), .B(n38645), .Z(n38638) );
  XOR U38539 ( .A(n38634), .B(n38633), .Z(n38645) );
  XNOR U38540 ( .A(n38679), .B(n38630), .Z(n38633) );
  XOR U38541 ( .A(n38680), .B(n38681), .Z(n38630) );
  AND U38542 ( .A(n38682), .B(n38683), .Z(n38681) );
  XOR U38543 ( .A(n38680), .B(n38684), .Z(n38682) );
  XNOR U38544 ( .A(n38685), .B(n38686), .Z(n38679) );
  NOR U38545 ( .A(n38687), .B(n38688), .Z(n38686) );
  XNOR U38546 ( .A(n38685), .B(n38689), .Z(n38687) );
  XOR U38547 ( .A(n38690), .B(n38691), .Z(n38634) );
  NOR U38548 ( .A(n38692), .B(n38693), .Z(n38691) );
  XNOR U38549 ( .A(n38690), .B(n38694), .Z(n38692) );
  XNOR U38550 ( .A(n38644), .B(n38635), .Z(n38678) );
  XOR U38551 ( .A(n38695), .B(n38696), .Z(n38635) );
  NOR U38552 ( .A(n38697), .B(n38698), .Z(n38696) );
  XNOR U38553 ( .A(n38695), .B(n38699), .Z(n38697) );
  XOR U38554 ( .A(n38700), .B(n38650), .Z(n38644) );
  XNOR U38555 ( .A(n38701), .B(n38702), .Z(n38650) );
  NOR U38556 ( .A(n38703), .B(n38704), .Z(n38702) );
  XNOR U38557 ( .A(n38701), .B(n38705), .Z(n38703) );
  XNOR U38558 ( .A(n38649), .B(n38641), .Z(n38700) );
  XOR U38559 ( .A(n38706), .B(n38707), .Z(n38641) );
  AND U38560 ( .A(n38708), .B(n38709), .Z(n38707) );
  XOR U38561 ( .A(n38706), .B(n38710), .Z(n38708) );
  XNOR U38562 ( .A(n38711), .B(n38646), .Z(n38649) );
  XOR U38563 ( .A(n38712), .B(n38713), .Z(n38646) );
  AND U38564 ( .A(n38714), .B(n38715), .Z(n38713) );
  XOR U38565 ( .A(n38712), .B(n38716), .Z(n38714) );
  XNOR U38566 ( .A(n38717), .B(n38718), .Z(n38711) );
  NOR U38567 ( .A(n38719), .B(n38720), .Z(n38718) );
  XOR U38568 ( .A(n38717), .B(n38721), .Z(n38719) );
  XOR U38569 ( .A(n38639), .B(n38651), .Z(n38677) );
  NOR U38570 ( .A(n38568), .B(n38722), .Z(n38651) );
  XNOR U38571 ( .A(n38657), .B(n38656), .Z(n38639) );
  XNOR U38572 ( .A(n38723), .B(n38662), .Z(n38656) );
  XOR U38573 ( .A(n38724), .B(n38725), .Z(n38662) );
  NOR U38574 ( .A(n38726), .B(n38727), .Z(n38725) );
  XNOR U38575 ( .A(n38724), .B(n38728), .Z(n38726) );
  XNOR U38576 ( .A(n38661), .B(n38653), .Z(n38723) );
  XOR U38577 ( .A(n38729), .B(n38730), .Z(n38653) );
  AND U38578 ( .A(n38731), .B(n38732), .Z(n38730) );
  XNOR U38579 ( .A(n38729), .B(n38733), .Z(n38731) );
  XNOR U38580 ( .A(n38734), .B(n38658), .Z(n38661) );
  XOR U38581 ( .A(n38735), .B(n38736), .Z(n38658) );
  AND U38582 ( .A(n38737), .B(n38738), .Z(n38736) );
  XOR U38583 ( .A(n38735), .B(n38739), .Z(n38737) );
  XNOR U38584 ( .A(n38740), .B(n38741), .Z(n38734) );
  NOR U38585 ( .A(n38742), .B(n38743), .Z(n38741) );
  XOR U38586 ( .A(n38740), .B(n38744), .Z(n38742) );
  XOR U38587 ( .A(n38667), .B(n38666), .Z(n38657) );
  XNOR U38588 ( .A(n38745), .B(n38663), .Z(n38666) );
  XOR U38589 ( .A(n38746), .B(n38747), .Z(n38663) );
  AND U38590 ( .A(n38748), .B(n38749), .Z(n38747) );
  XOR U38591 ( .A(n38746), .B(n38750), .Z(n38748) );
  XNOR U38592 ( .A(n38751), .B(n38752), .Z(n38745) );
  NOR U38593 ( .A(n38753), .B(n38754), .Z(n38752) );
  XNOR U38594 ( .A(n38751), .B(n38755), .Z(n38753) );
  XOR U38595 ( .A(n38756), .B(n38757), .Z(n38667) );
  NOR U38596 ( .A(n38758), .B(n38759), .Z(n38757) );
  XNOR U38597 ( .A(n38756), .B(n38760), .Z(n38758) );
  XNOR U38598 ( .A(n38559), .B(n38673), .Z(n38675) );
  XNOR U38599 ( .A(n38761), .B(n38762), .Z(n38559) );
  AND U38600 ( .A(n686), .B(n38763), .Z(n38762) );
  XNOR U38601 ( .A(n38764), .B(n38765), .Z(n38763) );
  AND U38602 ( .A(n38565), .B(n38568), .Z(n38673) );
  XOR U38603 ( .A(n38766), .B(n38722), .Z(n38568) );
  XNOR U38604 ( .A(p_input[2048]), .B(p_input[928]), .Z(n38722) );
  XOR U38605 ( .A(n38699), .B(n38698), .Z(n38766) );
  XOR U38606 ( .A(n38767), .B(n38710), .Z(n38698) );
  XOR U38607 ( .A(n38684), .B(n38683), .Z(n38710) );
  XNOR U38608 ( .A(n38768), .B(n38689), .Z(n38683) );
  XOR U38609 ( .A(p_input[2072]), .B(p_input[952]), .Z(n38689) );
  XOR U38610 ( .A(n38680), .B(n38688), .Z(n38768) );
  XOR U38611 ( .A(n38769), .B(n38685), .Z(n38688) );
  XOR U38612 ( .A(p_input[2070]), .B(p_input[950]), .Z(n38685) );
  XNOR U38613 ( .A(p_input[2071]), .B(p_input[951]), .Z(n38769) );
  XNOR U38614 ( .A(n28684), .B(p_input[946]), .Z(n38680) );
  XNOR U38615 ( .A(n38694), .B(n38693), .Z(n38684) );
  XOR U38616 ( .A(n38770), .B(n38690), .Z(n38693) );
  XOR U38617 ( .A(p_input[2067]), .B(p_input[947]), .Z(n38690) );
  XNOR U38618 ( .A(p_input[2068]), .B(p_input[948]), .Z(n38770) );
  XOR U38619 ( .A(p_input[2069]), .B(p_input[949]), .Z(n38694) );
  XNOR U38620 ( .A(n38709), .B(n38695), .Z(n38767) );
  XNOR U38621 ( .A(n28686), .B(p_input[929]), .Z(n38695) );
  XNOR U38622 ( .A(n38771), .B(n38716), .Z(n38709) );
  XNOR U38623 ( .A(n38705), .B(n38704), .Z(n38716) );
  XOR U38624 ( .A(n38772), .B(n38701), .Z(n38704) );
  XNOR U38625 ( .A(n28322), .B(p_input[954]), .Z(n38701) );
  XNOR U38626 ( .A(p_input[2075]), .B(p_input[955]), .Z(n38772) );
  XOR U38627 ( .A(p_input[2076]), .B(p_input[956]), .Z(n38705) );
  XNOR U38628 ( .A(n38715), .B(n38706), .Z(n38771) );
  XNOR U38629 ( .A(n28689), .B(p_input[945]), .Z(n38706) );
  XOR U38630 ( .A(n38773), .B(n38721), .Z(n38715) );
  XNOR U38631 ( .A(p_input[2079]), .B(p_input[959]), .Z(n38721) );
  XOR U38632 ( .A(n38712), .B(n38720), .Z(n38773) );
  XOR U38633 ( .A(n38774), .B(n38717), .Z(n38720) );
  XOR U38634 ( .A(p_input[2077]), .B(p_input[957]), .Z(n38717) );
  XNOR U38635 ( .A(p_input[2078]), .B(p_input[958]), .Z(n38774) );
  XNOR U38636 ( .A(n28326), .B(p_input[953]), .Z(n38712) );
  XNOR U38637 ( .A(n38733), .B(n38732), .Z(n38699) );
  XNOR U38638 ( .A(n38775), .B(n38739), .Z(n38732) );
  XNOR U38639 ( .A(n38728), .B(n38727), .Z(n38739) );
  XOR U38640 ( .A(n38776), .B(n38724), .Z(n38727) );
  XNOR U38641 ( .A(n28694), .B(p_input[939]), .Z(n38724) );
  XNOR U38642 ( .A(p_input[2060]), .B(p_input[940]), .Z(n38776) );
  XOR U38643 ( .A(p_input[2061]), .B(p_input[941]), .Z(n38728) );
  XNOR U38644 ( .A(n38738), .B(n38729), .Z(n38775) );
  XNOR U38645 ( .A(n28330), .B(p_input[930]), .Z(n38729) );
  XOR U38646 ( .A(n38777), .B(n38744), .Z(n38738) );
  XNOR U38647 ( .A(p_input[2064]), .B(p_input[944]), .Z(n38744) );
  XOR U38648 ( .A(n38735), .B(n38743), .Z(n38777) );
  XOR U38649 ( .A(n38778), .B(n38740), .Z(n38743) );
  XOR U38650 ( .A(p_input[2062]), .B(p_input[942]), .Z(n38740) );
  XNOR U38651 ( .A(p_input[2063]), .B(p_input[943]), .Z(n38778) );
  XNOR U38652 ( .A(n28697), .B(p_input[938]), .Z(n38735) );
  XNOR U38653 ( .A(n38750), .B(n38749), .Z(n38733) );
  XNOR U38654 ( .A(n38779), .B(n38755), .Z(n38749) );
  XOR U38655 ( .A(p_input[2057]), .B(p_input[937]), .Z(n38755) );
  XOR U38656 ( .A(n38746), .B(n38754), .Z(n38779) );
  XOR U38657 ( .A(n38780), .B(n38751), .Z(n38754) );
  XOR U38658 ( .A(p_input[2055]), .B(p_input[935]), .Z(n38751) );
  XNOR U38659 ( .A(p_input[2056]), .B(p_input[936]), .Z(n38780) );
  XNOR U38660 ( .A(n28337), .B(p_input[931]), .Z(n38746) );
  XNOR U38661 ( .A(n38760), .B(n38759), .Z(n38750) );
  XOR U38662 ( .A(n38781), .B(n38756), .Z(n38759) );
  XOR U38663 ( .A(p_input[2052]), .B(p_input[932]), .Z(n38756) );
  XNOR U38664 ( .A(p_input[2053]), .B(p_input[933]), .Z(n38781) );
  XOR U38665 ( .A(p_input[2054]), .B(p_input[934]), .Z(n38760) );
  XNOR U38666 ( .A(n38782), .B(n38783), .Z(n38565) );
  AND U38667 ( .A(n686), .B(n38784), .Z(n38783) );
  XNOR U38668 ( .A(n38785), .B(n38786), .Z(n686) );
  AND U38669 ( .A(n38787), .B(n38788), .Z(n38786) );
  XOR U38670 ( .A(n38579), .B(n38785), .Z(n38788) );
  XNOR U38671 ( .A(n38789), .B(n38785), .Z(n38787) );
  XOR U38672 ( .A(n38790), .B(n38791), .Z(n38785) );
  AND U38673 ( .A(n38792), .B(n38793), .Z(n38791) );
  XOR U38674 ( .A(n38594), .B(n38790), .Z(n38793) );
  XOR U38675 ( .A(n38790), .B(n38595), .Z(n38792) );
  XOR U38676 ( .A(n38794), .B(n38795), .Z(n38790) );
  AND U38677 ( .A(n38796), .B(n38797), .Z(n38795) );
  XOR U38678 ( .A(n38622), .B(n38794), .Z(n38797) );
  XOR U38679 ( .A(n38794), .B(n38623), .Z(n38796) );
  XOR U38680 ( .A(n38798), .B(n38799), .Z(n38794) );
  AND U38681 ( .A(n38800), .B(n38801), .Z(n38799) );
  XOR U38682 ( .A(n38671), .B(n38798), .Z(n38801) );
  XOR U38683 ( .A(n38798), .B(n38672), .Z(n38800) );
  XOR U38684 ( .A(n38802), .B(n38803), .Z(n38798) );
  AND U38685 ( .A(n38804), .B(n38805), .Z(n38803) );
  XOR U38686 ( .A(n38802), .B(n38764), .Z(n38805) );
  XNOR U38687 ( .A(n38806), .B(n38807), .Z(n38515) );
  AND U38688 ( .A(n690), .B(n38808), .Z(n38807) );
  XNOR U38689 ( .A(n38809), .B(n38810), .Z(n690) );
  AND U38690 ( .A(n38811), .B(n38812), .Z(n38810) );
  XOR U38691 ( .A(n38809), .B(n38525), .Z(n38812) );
  XNOR U38692 ( .A(n38809), .B(n38475), .Z(n38811) );
  XOR U38693 ( .A(n38813), .B(n38814), .Z(n38809) );
  AND U38694 ( .A(n38815), .B(n38816), .Z(n38814) );
  XNOR U38695 ( .A(n38535), .B(n38813), .Z(n38816) );
  XOR U38696 ( .A(n38813), .B(n38485), .Z(n38815) );
  XOR U38697 ( .A(n38817), .B(n38818), .Z(n38813) );
  AND U38698 ( .A(n38819), .B(n38820), .Z(n38818) );
  XNOR U38699 ( .A(n38545), .B(n38817), .Z(n38820) );
  XOR U38700 ( .A(n38817), .B(n38494), .Z(n38819) );
  XOR U38701 ( .A(n38821), .B(n38822), .Z(n38817) );
  AND U38702 ( .A(n38823), .B(n38824), .Z(n38822) );
  XOR U38703 ( .A(n38821), .B(n38502), .Z(n38823) );
  XOR U38704 ( .A(n38825), .B(n38826), .Z(n38466) );
  AND U38705 ( .A(n694), .B(n38808), .Z(n38826) );
  XNOR U38706 ( .A(n38806), .B(n38825), .Z(n38808) );
  XNOR U38707 ( .A(n38827), .B(n38828), .Z(n694) );
  AND U38708 ( .A(n38829), .B(n38830), .Z(n38828) );
  XNOR U38709 ( .A(n38831), .B(n38827), .Z(n38830) );
  IV U38710 ( .A(n38525), .Z(n38831) );
  XOR U38711 ( .A(n38789), .B(n38832), .Z(n38525) );
  AND U38712 ( .A(n697), .B(n38833), .Z(n38832) );
  XOR U38713 ( .A(n38578), .B(n38575), .Z(n38833) );
  IV U38714 ( .A(n38789), .Z(n38578) );
  XNOR U38715 ( .A(n38475), .B(n38827), .Z(n38829) );
  XOR U38716 ( .A(n38834), .B(n38835), .Z(n38475) );
  AND U38717 ( .A(n713), .B(n38836), .Z(n38835) );
  XOR U38718 ( .A(n38837), .B(n38838), .Z(n38827) );
  AND U38719 ( .A(n38839), .B(n38840), .Z(n38838) );
  XNOR U38720 ( .A(n38837), .B(n38535), .Z(n38840) );
  XOR U38721 ( .A(n38595), .B(n38841), .Z(n38535) );
  AND U38722 ( .A(n697), .B(n38842), .Z(n38841) );
  XOR U38723 ( .A(n38591), .B(n38595), .Z(n38842) );
  XNOR U38724 ( .A(n38843), .B(n38837), .Z(n38839) );
  IV U38725 ( .A(n38485), .Z(n38843) );
  XOR U38726 ( .A(n38844), .B(n38845), .Z(n38485) );
  AND U38727 ( .A(n713), .B(n38846), .Z(n38845) );
  XOR U38728 ( .A(n38847), .B(n38848), .Z(n38837) );
  AND U38729 ( .A(n38849), .B(n38850), .Z(n38848) );
  XNOR U38730 ( .A(n38847), .B(n38545), .Z(n38850) );
  XOR U38731 ( .A(n38623), .B(n38851), .Z(n38545) );
  AND U38732 ( .A(n697), .B(n38852), .Z(n38851) );
  XOR U38733 ( .A(n38619), .B(n38623), .Z(n38852) );
  XOR U38734 ( .A(n38494), .B(n38847), .Z(n38849) );
  XOR U38735 ( .A(n38853), .B(n38854), .Z(n38494) );
  AND U38736 ( .A(n713), .B(n38855), .Z(n38854) );
  XOR U38737 ( .A(n38821), .B(n38856), .Z(n38847) );
  AND U38738 ( .A(n38857), .B(n38824), .Z(n38856) );
  XNOR U38739 ( .A(n38555), .B(n38821), .Z(n38824) );
  XOR U38740 ( .A(n38672), .B(n38858), .Z(n38555) );
  AND U38741 ( .A(n697), .B(n38859), .Z(n38858) );
  XOR U38742 ( .A(n38668), .B(n38672), .Z(n38859) );
  XNOR U38743 ( .A(n38860), .B(n38821), .Z(n38857) );
  IV U38744 ( .A(n38502), .Z(n38860) );
  XOR U38745 ( .A(n38861), .B(n38862), .Z(n38502) );
  AND U38746 ( .A(n713), .B(n38863), .Z(n38862) );
  XOR U38747 ( .A(n38864), .B(n38865), .Z(n38821) );
  AND U38748 ( .A(n38866), .B(n38867), .Z(n38865) );
  XNOR U38749 ( .A(n38864), .B(n38563), .Z(n38867) );
  XOR U38750 ( .A(n38765), .B(n38868), .Z(n38563) );
  AND U38751 ( .A(n697), .B(n38869), .Z(n38868) );
  XOR U38752 ( .A(n38761), .B(n38765), .Z(n38869) );
  XNOR U38753 ( .A(n38870), .B(n38864), .Z(n38866) );
  IV U38754 ( .A(n38512), .Z(n38870) );
  XOR U38755 ( .A(n38871), .B(n38872), .Z(n38512) );
  AND U38756 ( .A(n713), .B(n38873), .Z(n38872) );
  AND U38757 ( .A(n38825), .B(n38806), .Z(n38864) );
  XNOR U38758 ( .A(n38874), .B(n38875), .Z(n38806) );
  AND U38759 ( .A(n697), .B(n38784), .Z(n38875) );
  XNOR U38760 ( .A(n38782), .B(n38874), .Z(n38784) );
  XNOR U38761 ( .A(n38876), .B(n38877), .Z(n697) );
  AND U38762 ( .A(n38878), .B(n38879), .Z(n38877) );
  XNOR U38763 ( .A(n38876), .B(n38575), .Z(n38879) );
  IV U38764 ( .A(n38579), .Z(n38575) );
  XOR U38765 ( .A(n38880), .B(n38881), .Z(n38579) );
  AND U38766 ( .A(n701), .B(n38882), .Z(n38881) );
  XOR U38767 ( .A(n38883), .B(n38880), .Z(n38882) );
  XNOR U38768 ( .A(n38876), .B(n38789), .Z(n38878) );
  XOR U38769 ( .A(n38884), .B(n38885), .Z(n38789) );
  AND U38770 ( .A(n709), .B(n38836), .Z(n38885) );
  XOR U38771 ( .A(n38834), .B(n38884), .Z(n38836) );
  XOR U38772 ( .A(n38886), .B(n38887), .Z(n38876) );
  AND U38773 ( .A(n38888), .B(n38889), .Z(n38887) );
  XNOR U38774 ( .A(n38886), .B(n38591), .Z(n38889) );
  IV U38775 ( .A(n38594), .Z(n38591) );
  XOR U38776 ( .A(n38890), .B(n38891), .Z(n38594) );
  AND U38777 ( .A(n701), .B(n38892), .Z(n38891) );
  XOR U38778 ( .A(n38893), .B(n38890), .Z(n38892) );
  XOR U38779 ( .A(n38595), .B(n38886), .Z(n38888) );
  XOR U38780 ( .A(n38894), .B(n38895), .Z(n38595) );
  AND U38781 ( .A(n709), .B(n38846), .Z(n38895) );
  XOR U38782 ( .A(n38894), .B(n38844), .Z(n38846) );
  XOR U38783 ( .A(n38896), .B(n38897), .Z(n38886) );
  AND U38784 ( .A(n38898), .B(n38899), .Z(n38897) );
  XNOR U38785 ( .A(n38896), .B(n38619), .Z(n38899) );
  IV U38786 ( .A(n38622), .Z(n38619) );
  XOR U38787 ( .A(n38900), .B(n38901), .Z(n38622) );
  AND U38788 ( .A(n701), .B(n38902), .Z(n38901) );
  XNOR U38789 ( .A(n38903), .B(n38900), .Z(n38902) );
  XOR U38790 ( .A(n38623), .B(n38896), .Z(n38898) );
  XOR U38791 ( .A(n38904), .B(n38905), .Z(n38623) );
  AND U38792 ( .A(n709), .B(n38855), .Z(n38905) );
  XOR U38793 ( .A(n38904), .B(n38853), .Z(n38855) );
  XOR U38794 ( .A(n38906), .B(n38907), .Z(n38896) );
  AND U38795 ( .A(n38908), .B(n38909), .Z(n38907) );
  XNOR U38796 ( .A(n38906), .B(n38668), .Z(n38909) );
  IV U38797 ( .A(n38671), .Z(n38668) );
  XOR U38798 ( .A(n38910), .B(n38911), .Z(n38671) );
  AND U38799 ( .A(n701), .B(n38912), .Z(n38911) );
  XOR U38800 ( .A(n38913), .B(n38910), .Z(n38912) );
  XOR U38801 ( .A(n38672), .B(n38906), .Z(n38908) );
  XOR U38802 ( .A(n38914), .B(n38915), .Z(n38672) );
  AND U38803 ( .A(n709), .B(n38863), .Z(n38915) );
  XOR U38804 ( .A(n38914), .B(n38861), .Z(n38863) );
  XOR U38805 ( .A(n38802), .B(n38916), .Z(n38906) );
  AND U38806 ( .A(n38804), .B(n38917), .Z(n38916) );
  XNOR U38807 ( .A(n38802), .B(n38761), .Z(n38917) );
  IV U38808 ( .A(n38764), .Z(n38761) );
  XOR U38809 ( .A(n38918), .B(n38919), .Z(n38764) );
  AND U38810 ( .A(n701), .B(n38920), .Z(n38919) );
  XNOR U38811 ( .A(n38921), .B(n38918), .Z(n38920) );
  XOR U38812 ( .A(n38765), .B(n38802), .Z(n38804) );
  XOR U38813 ( .A(n38922), .B(n38923), .Z(n38765) );
  AND U38814 ( .A(n709), .B(n38873), .Z(n38923) );
  XOR U38815 ( .A(n38922), .B(n38871), .Z(n38873) );
  AND U38816 ( .A(n38874), .B(n38782), .Z(n38802) );
  XNOR U38817 ( .A(n38924), .B(n38925), .Z(n38782) );
  AND U38818 ( .A(n701), .B(n38926), .Z(n38925) );
  XNOR U38819 ( .A(n38927), .B(n38924), .Z(n38926) );
  XNOR U38820 ( .A(n38928), .B(n38929), .Z(n701) );
  AND U38821 ( .A(n38930), .B(n38931), .Z(n38929) );
  XOR U38822 ( .A(n38883), .B(n38928), .Z(n38931) );
  AND U38823 ( .A(n38932), .B(n38933), .Z(n38883) );
  XNOR U38824 ( .A(n38880), .B(n38928), .Z(n38930) );
  XNOR U38825 ( .A(n38934), .B(n38935), .Z(n38880) );
  AND U38826 ( .A(n705), .B(n38936), .Z(n38935) );
  XNOR U38827 ( .A(n38937), .B(n38938), .Z(n38936) );
  XOR U38828 ( .A(n38939), .B(n38940), .Z(n38928) );
  AND U38829 ( .A(n38941), .B(n38942), .Z(n38940) );
  XNOR U38830 ( .A(n38939), .B(n38932), .Z(n38942) );
  IV U38831 ( .A(n38893), .Z(n38932) );
  XOR U38832 ( .A(n38943), .B(n38944), .Z(n38893) );
  XOR U38833 ( .A(n38945), .B(n38933), .Z(n38944) );
  AND U38834 ( .A(n38903), .B(n38946), .Z(n38933) );
  AND U38835 ( .A(n38947), .B(n38948), .Z(n38945) );
  XOR U38836 ( .A(n38949), .B(n38943), .Z(n38947) );
  XNOR U38837 ( .A(n38890), .B(n38939), .Z(n38941) );
  XNOR U38838 ( .A(n38950), .B(n38951), .Z(n38890) );
  AND U38839 ( .A(n705), .B(n38952), .Z(n38951) );
  XNOR U38840 ( .A(n38953), .B(n38954), .Z(n38952) );
  XOR U38841 ( .A(n38955), .B(n38956), .Z(n38939) );
  AND U38842 ( .A(n38957), .B(n38958), .Z(n38956) );
  XNOR U38843 ( .A(n38955), .B(n38903), .Z(n38958) );
  XOR U38844 ( .A(n38959), .B(n38948), .Z(n38903) );
  XNOR U38845 ( .A(n38960), .B(n38943), .Z(n38948) );
  XOR U38846 ( .A(n38961), .B(n38962), .Z(n38943) );
  AND U38847 ( .A(n38963), .B(n38964), .Z(n38962) );
  XOR U38848 ( .A(n38965), .B(n38961), .Z(n38963) );
  XNOR U38849 ( .A(n38966), .B(n38967), .Z(n38960) );
  AND U38850 ( .A(n38968), .B(n38969), .Z(n38967) );
  XOR U38851 ( .A(n38966), .B(n38970), .Z(n38968) );
  XNOR U38852 ( .A(n38949), .B(n38946), .Z(n38959) );
  AND U38853 ( .A(n38971), .B(n38972), .Z(n38946) );
  XOR U38854 ( .A(n38973), .B(n38974), .Z(n38949) );
  AND U38855 ( .A(n38975), .B(n38976), .Z(n38974) );
  XOR U38856 ( .A(n38973), .B(n38977), .Z(n38975) );
  XNOR U38857 ( .A(n38900), .B(n38955), .Z(n38957) );
  XNOR U38858 ( .A(n38978), .B(n38979), .Z(n38900) );
  AND U38859 ( .A(n705), .B(n38980), .Z(n38979) );
  XNOR U38860 ( .A(n38981), .B(n38982), .Z(n38980) );
  XOR U38861 ( .A(n38983), .B(n38984), .Z(n38955) );
  AND U38862 ( .A(n38985), .B(n38986), .Z(n38984) );
  XNOR U38863 ( .A(n38983), .B(n38971), .Z(n38986) );
  IV U38864 ( .A(n38913), .Z(n38971) );
  XNOR U38865 ( .A(n38987), .B(n38964), .Z(n38913) );
  XNOR U38866 ( .A(n38988), .B(n38970), .Z(n38964) );
  XOR U38867 ( .A(n38989), .B(n38990), .Z(n38970) );
  AND U38868 ( .A(n38991), .B(n38992), .Z(n38990) );
  XOR U38869 ( .A(n38989), .B(n38993), .Z(n38991) );
  XNOR U38870 ( .A(n38969), .B(n38961), .Z(n38988) );
  XOR U38871 ( .A(n38994), .B(n38995), .Z(n38961) );
  AND U38872 ( .A(n38996), .B(n38997), .Z(n38995) );
  XNOR U38873 ( .A(n38998), .B(n38994), .Z(n38996) );
  XNOR U38874 ( .A(n38999), .B(n38966), .Z(n38969) );
  XOR U38875 ( .A(n39000), .B(n39001), .Z(n38966) );
  AND U38876 ( .A(n39002), .B(n39003), .Z(n39001) );
  XOR U38877 ( .A(n39000), .B(n39004), .Z(n39002) );
  XNOR U38878 ( .A(n39005), .B(n39006), .Z(n38999) );
  AND U38879 ( .A(n39007), .B(n39008), .Z(n39006) );
  XNOR U38880 ( .A(n39005), .B(n39009), .Z(n39007) );
  XNOR U38881 ( .A(n38965), .B(n38972), .Z(n38987) );
  AND U38882 ( .A(n38921), .B(n39010), .Z(n38972) );
  XOR U38883 ( .A(n38977), .B(n38976), .Z(n38965) );
  XNOR U38884 ( .A(n39011), .B(n38973), .Z(n38976) );
  XOR U38885 ( .A(n39012), .B(n39013), .Z(n38973) );
  AND U38886 ( .A(n39014), .B(n39015), .Z(n39013) );
  XOR U38887 ( .A(n39012), .B(n39016), .Z(n39014) );
  XNOR U38888 ( .A(n39017), .B(n39018), .Z(n39011) );
  AND U38889 ( .A(n39019), .B(n39020), .Z(n39018) );
  XOR U38890 ( .A(n39017), .B(n39021), .Z(n39019) );
  XOR U38891 ( .A(n39022), .B(n39023), .Z(n38977) );
  AND U38892 ( .A(n39024), .B(n39025), .Z(n39023) );
  XOR U38893 ( .A(n39022), .B(n39026), .Z(n39024) );
  XNOR U38894 ( .A(n38910), .B(n38983), .Z(n38985) );
  XNOR U38895 ( .A(n39027), .B(n39028), .Z(n38910) );
  AND U38896 ( .A(n705), .B(n39029), .Z(n39028) );
  XNOR U38897 ( .A(n39030), .B(n39031), .Z(n39029) );
  XOR U38898 ( .A(n39032), .B(n39033), .Z(n38983) );
  AND U38899 ( .A(n39034), .B(n39035), .Z(n39033) );
  XNOR U38900 ( .A(n39032), .B(n38921), .Z(n39035) );
  XOR U38901 ( .A(n39036), .B(n38997), .Z(n38921) );
  XNOR U38902 ( .A(n39037), .B(n39004), .Z(n38997) );
  XOR U38903 ( .A(n38993), .B(n38992), .Z(n39004) );
  XNOR U38904 ( .A(n39038), .B(n38989), .Z(n38992) );
  XOR U38905 ( .A(n39039), .B(n39040), .Z(n38989) );
  AND U38906 ( .A(n39041), .B(n39042), .Z(n39040) );
  XOR U38907 ( .A(n39039), .B(n39043), .Z(n39041) );
  XNOR U38908 ( .A(n39044), .B(n39045), .Z(n39038) );
  NOR U38909 ( .A(n39046), .B(n39047), .Z(n39045) );
  XNOR U38910 ( .A(n39044), .B(n39048), .Z(n39046) );
  XOR U38911 ( .A(n39049), .B(n39050), .Z(n38993) );
  NOR U38912 ( .A(n39051), .B(n39052), .Z(n39050) );
  XNOR U38913 ( .A(n39049), .B(n39053), .Z(n39051) );
  XNOR U38914 ( .A(n39003), .B(n38994), .Z(n39037) );
  XOR U38915 ( .A(n39054), .B(n39055), .Z(n38994) );
  NOR U38916 ( .A(n39056), .B(n39057), .Z(n39055) );
  XNOR U38917 ( .A(n39054), .B(n39058), .Z(n39056) );
  XOR U38918 ( .A(n39059), .B(n39009), .Z(n39003) );
  XNOR U38919 ( .A(n39060), .B(n39061), .Z(n39009) );
  NOR U38920 ( .A(n39062), .B(n39063), .Z(n39061) );
  XNOR U38921 ( .A(n39060), .B(n39064), .Z(n39062) );
  XNOR U38922 ( .A(n39008), .B(n39000), .Z(n39059) );
  XOR U38923 ( .A(n39065), .B(n39066), .Z(n39000) );
  AND U38924 ( .A(n39067), .B(n39068), .Z(n39066) );
  XOR U38925 ( .A(n39065), .B(n39069), .Z(n39067) );
  XNOR U38926 ( .A(n39070), .B(n39005), .Z(n39008) );
  XOR U38927 ( .A(n39071), .B(n39072), .Z(n39005) );
  AND U38928 ( .A(n39073), .B(n39074), .Z(n39072) );
  XOR U38929 ( .A(n39071), .B(n39075), .Z(n39073) );
  XNOR U38930 ( .A(n39076), .B(n39077), .Z(n39070) );
  NOR U38931 ( .A(n39078), .B(n39079), .Z(n39077) );
  XOR U38932 ( .A(n39076), .B(n39080), .Z(n39078) );
  XOR U38933 ( .A(n38998), .B(n39010), .Z(n39036) );
  NOR U38934 ( .A(n38927), .B(n39081), .Z(n39010) );
  XNOR U38935 ( .A(n39016), .B(n39015), .Z(n38998) );
  XNOR U38936 ( .A(n39082), .B(n39021), .Z(n39015) );
  XOR U38937 ( .A(n39083), .B(n39084), .Z(n39021) );
  NOR U38938 ( .A(n39085), .B(n39086), .Z(n39084) );
  XNOR U38939 ( .A(n39083), .B(n39087), .Z(n39085) );
  XNOR U38940 ( .A(n39020), .B(n39012), .Z(n39082) );
  XOR U38941 ( .A(n39088), .B(n39089), .Z(n39012) );
  AND U38942 ( .A(n39090), .B(n39091), .Z(n39089) );
  XNOR U38943 ( .A(n39088), .B(n39092), .Z(n39090) );
  XNOR U38944 ( .A(n39093), .B(n39017), .Z(n39020) );
  XOR U38945 ( .A(n39094), .B(n39095), .Z(n39017) );
  AND U38946 ( .A(n39096), .B(n39097), .Z(n39095) );
  XOR U38947 ( .A(n39094), .B(n39098), .Z(n39096) );
  XNOR U38948 ( .A(n39099), .B(n39100), .Z(n39093) );
  NOR U38949 ( .A(n39101), .B(n39102), .Z(n39100) );
  XOR U38950 ( .A(n39099), .B(n39103), .Z(n39101) );
  XOR U38951 ( .A(n39026), .B(n39025), .Z(n39016) );
  XNOR U38952 ( .A(n39104), .B(n39022), .Z(n39025) );
  XOR U38953 ( .A(n39105), .B(n39106), .Z(n39022) );
  AND U38954 ( .A(n39107), .B(n39108), .Z(n39106) );
  XOR U38955 ( .A(n39105), .B(n39109), .Z(n39107) );
  XNOR U38956 ( .A(n39110), .B(n39111), .Z(n39104) );
  NOR U38957 ( .A(n39112), .B(n39113), .Z(n39111) );
  XNOR U38958 ( .A(n39110), .B(n39114), .Z(n39112) );
  XOR U38959 ( .A(n39115), .B(n39116), .Z(n39026) );
  NOR U38960 ( .A(n39117), .B(n39118), .Z(n39116) );
  XNOR U38961 ( .A(n39115), .B(n39119), .Z(n39117) );
  XNOR U38962 ( .A(n38918), .B(n39032), .Z(n39034) );
  XNOR U38963 ( .A(n39120), .B(n39121), .Z(n38918) );
  AND U38964 ( .A(n705), .B(n39122), .Z(n39121) );
  XNOR U38965 ( .A(n39123), .B(n39124), .Z(n39122) );
  AND U38966 ( .A(n38924), .B(n38927), .Z(n39032) );
  XOR U38967 ( .A(n39125), .B(n39081), .Z(n38927) );
  XNOR U38968 ( .A(p_input[2048]), .B(p_input[960]), .Z(n39081) );
  XOR U38969 ( .A(n39058), .B(n39057), .Z(n39125) );
  XOR U38970 ( .A(n39126), .B(n39069), .Z(n39057) );
  XOR U38971 ( .A(n39043), .B(n39042), .Z(n39069) );
  XNOR U38972 ( .A(n39127), .B(n39048), .Z(n39042) );
  XOR U38973 ( .A(p_input[2072]), .B(p_input[984]), .Z(n39048) );
  XOR U38974 ( .A(n39039), .B(n39047), .Z(n39127) );
  XOR U38975 ( .A(n39128), .B(n39044), .Z(n39047) );
  XOR U38976 ( .A(p_input[2070]), .B(p_input[982]), .Z(n39044) );
  XNOR U38977 ( .A(p_input[2071]), .B(p_input[983]), .Z(n39128) );
  XNOR U38978 ( .A(n28684), .B(p_input[978]), .Z(n39039) );
  XNOR U38979 ( .A(n39053), .B(n39052), .Z(n39043) );
  XOR U38980 ( .A(n39129), .B(n39049), .Z(n39052) );
  XOR U38981 ( .A(p_input[2067]), .B(p_input[979]), .Z(n39049) );
  XNOR U38982 ( .A(p_input[2068]), .B(p_input[980]), .Z(n39129) );
  XOR U38983 ( .A(p_input[2069]), .B(p_input[981]), .Z(n39053) );
  XNOR U38984 ( .A(n39068), .B(n39054), .Z(n39126) );
  XNOR U38985 ( .A(n28686), .B(p_input[961]), .Z(n39054) );
  XNOR U38986 ( .A(n39130), .B(n39075), .Z(n39068) );
  XNOR U38987 ( .A(n39064), .B(n39063), .Z(n39075) );
  XOR U38988 ( .A(n39131), .B(n39060), .Z(n39063) );
  XNOR U38989 ( .A(n28322), .B(p_input[986]), .Z(n39060) );
  XNOR U38990 ( .A(p_input[2075]), .B(p_input[987]), .Z(n39131) );
  XOR U38991 ( .A(p_input[2076]), .B(p_input[988]), .Z(n39064) );
  XNOR U38992 ( .A(n39074), .B(n39065), .Z(n39130) );
  XNOR U38993 ( .A(n28689), .B(p_input[977]), .Z(n39065) );
  XOR U38994 ( .A(n39132), .B(n39080), .Z(n39074) );
  XNOR U38995 ( .A(p_input[2079]), .B(p_input[991]), .Z(n39080) );
  XOR U38996 ( .A(n39071), .B(n39079), .Z(n39132) );
  XOR U38997 ( .A(n39133), .B(n39076), .Z(n39079) );
  XOR U38998 ( .A(p_input[2077]), .B(p_input[989]), .Z(n39076) );
  XNOR U38999 ( .A(p_input[2078]), .B(p_input[990]), .Z(n39133) );
  XNOR U39000 ( .A(n28326), .B(p_input[985]), .Z(n39071) );
  XNOR U39001 ( .A(n39092), .B(n39091), .Z(n39058) );
  XNOR U39002 ( .A(n39134), .B(n39098), .Z(n39091) );
  XNOR U39003 ( .A(n39087), .B(n39086), .Z(n39098) );
  XOR U39004 ( .A(n39135), .B(n39083), .Z(n39086) );
  XNOR U39005 ( .A(n28694), .B(p_input[971]), .Z(n39083) );
  XNOR U39006 ( .A(p_input[2060]), .B(p_input[972]), .Z(n39135) );
  XOR U39007 ( .A(p_input[2061]), .B(p_input[973]), .Z(n39087) );
  XNOR U39008 ( .A(n39097), .B(n39088), .Z(n39134) );
  XNOR U39009 ( .A(n28330), .B(p_input[962]), .Z(n39088) );
  XOR U39010 ( .A(n39136), .B(n39103), .Z(n39097) );
  XNOR U39011 ( .A(p_input[2064]), .B(p_input[976]), .Z(n39103) );
  XOR U39012 ( .A(n39094), .B(n39102), .Z(n39136) );
  XOR U39013 ( .A(n39137), .B(n39099), .Z(n39102) );
  XOR U39014 ( .A(p_input[2062]), .B(p_input[974]), .Z(n39099) );
  XNOR U39015 ( .A(p_input[2063]), .B(p_input[975]), .Z(n39137) );
  XNOR U39016 ( .A(n28697), .B(p_input[970]), .Z(n39094) );
  XNOR U39017 ( .A(n39109), .B(n39108), .Z(n39092) );
  XNOR U39018 ( .A(n39138), .B(n39114), .Z(n39108) );
  XOR U39019 ( .A(p_input[2057]), .B(p_input[969]), .Z(n39114) );
  XOR U39020 ( .A(n39105), .B(n39113), .Z(n39138) );
  XOR U39021 ( .A(n39139), .B(n39110), .Z(n39113) );
  XOR U39022 ( .A(p_input[2055]), .B(p_input[967]), .Z(n39110) );
  XNOR U39023 ( .A(p_input[2056]), .B(p_input[968]), .Z(n39139) );
  XNOR U39024 ( .A(n28337), .B(p_input[963]), .Z(n39105) );
  XNOR U39025 ( .A(n39119), .B(n39118), .Z(n39109) );
  XOR U39026 ( .A(n39140), .B(n39115), .Z(n39118) );
  XOR U39027 ( .A(p_input[2052]), .B(p_input[964]), .Z(n39115) );
  XNOR U39028 ( .A(p_input[2053]), .B(p_input[965]), .Z(n39140) );
  XOR U39029 ( .A(p_input[2054]), .B(p_input[966]), .Z(n39119) );
  XNOR U39030 ( .A(n39141), .B(n39142), .Z(n38924) );
  AND U39031 ( .A(n705), .B(n39143), .Z(n39142) );
  XNOR U39032 ( .A(n39144), .B(n39145), .Z(n705) );
  AND U39033 ( .A(n39146), .B(n39147), .Z(n39145) );
  XOR U39034 ( .A(n38938), .B(n39144), .Z(n39147) );
  XNOR U39035 ( .A(n39148), .B(n39144), .Z(n39146) );
  XOR U39036 ( .A(n39149), .B(n39150), .Z(n39144) );
  AND U39037 ( .A(n39151), .B(n39152), .Z(n39150) );
  XOR U39038 ( .A(n38953), .B(n39149), .Z(n39152) );
  XOR U39039 ( .A(n39149), .B(n38954), .Z(n39151) );
  XOR U39040 ( .A(n39153), .B(n39154), .Z(n39149) );
  AND U39041 ( .A(n39155), .B(n39156), .Z(n39154) );
  XOR U39042 ( .A(n38981), .B(n39153), .Z(n39156) );
  XOR U39043 ( .A(n39153), .B(n38982), .Z(n39155) );
  XOR U39044 ( .A(n39157), .B(n39158), .Z(n39153) );
  AND U39045 ( .A(n39159), .B(n39160), .Z(n39158) );
  XOR U39046 ( .A(n39030), .B(n39157), .Z(n39160) );
  XOR U39047 ( .A(n39157), .B(n39031), .Z(n39159) );
  XOR U39048 ( .A(n39161), .B(n39162), .Z(n39157) );
  AND U39049 ( .A(n39163), .B(n39164), .Z(n39162) );
  XOR U39050 ( .A(n39161), .B(n39123), .Z(n39164) );
  XNOR U39051 ( .A(n39165), .B(n39166), .Z(n38874) );
  AND U39052 ( .A(n709), .B(n39167), .Z(n39166) );
  XNOR U39053 ( .A(n39168), .B(n39169), .Z(n709) );
  AND U39054 ( .A(n39170), .B(n39171), .Z(n39169) );
  XOR U39055 ( .A(n39168), .B(n38884), .Z(n39171) );
  XNOR U39056 ( .A(n39168), .B(n38834), .Z(n39170) );
  XOR U39057 ( .A(n39172), .B(n39173), .Z(n39168) );
  AND U39058 ( .A(n39174), .B(n39175), .Z(n39173) );
  XNOR U39059 ( .A(n38894), .B(n39172), .Z(n39175) );
  XOR U39060 ( .A(n39172), .B(n38844), .Z(n39174) );
  XOR U39061 ( .A(n39176), .B(n39177), .Z(n39172) );
  AND U39062 ( .A(n39178), .B(n39179), .Z(n39177) );
  XNOR U39063 ( .A(n38904), .B(n39176), .Z(n39179) );
  XOR U39064 ( .A(n39176), .B(n38853), .Z(n39178) );
  XOR U39065 ( .A(n39180), .B(n39181), .Z(n39176) );
  AND U39066 ( .A(n39182), .B(n39183), .Z(n39181) );
  XOR U39067 ( .A(n39180), .B(n38861), .Z(n39182) );
  XOR U39068 ( .A(n39184), .B(n39185), .Z(n38825) );
  AND U39069 ( .A(n713), .B(n39167), .Z(n39185) );
  XNOR U39070 ( .A(n39165), .B(n39184), .Z(n39167) );
  XNOR U39071 ( .A(n39186), .B(n39187), .Z(n713) );
  AND U39072 ( .A(n39188), .B(n39189), .Z(n39187) );
  XNOR U39073 ( .A(n39190), .B(n39186), .Z(n39189) );
  IV U39074 ( .A(n38884), .Z(n39190) );
  XOR U39075 ( .A(n39148), .B(n39191), .Z(n38884) );
  AND U39076 ( .A(n716), .B(n39192), .Z(n39191) );
  XOR U39077 ( .A(n38937), .B(n38934), .Z(n39192) );
  IV U39078 ( .A(n39148), .Z(n38937) );
  XNOR U39079 ( .A(n38834), .B(n39186), .Z(n39188) );
  XOR U39080 ( .A(n39193), .B(n39194), .Z(n38834) );
  AND U39081 ( .A(n732), .B(n39195), .Z(n39194) );
  XOR U39082 ( .A(n39196), .B(n39197), .Z(n39186) );
  AND U39083 ( .A(n39198), .B(n39199), .Z(n39197) );
  XNOR U39084 ( .A(n39196), .B(n38894), .Z(n39199) );
  XOR U39085 ( .A(n38954), .B(n39200), .Z(n38894) );
  AND U39086 ( .A(n716), .B(n39201), .Z(n39200) );
  XOR U39087 ( .A(n38950), .B(n38954), .Z(n39201) );
  XNOR U39088 ( .A(n39202), .B(n39196), .Z(n39198) );
  IV U39089 ( .A(n38844), .Z(n39202) );
  XOR U39090 ( .A(n39203), .B(n39204), .Z(n38844) );
  AND U39091 ( .A(n732), .B(n39205), .Z(n39204) );
  XOR U39092 ( .A(n39206), .B(n39207), .Z(n39196) );
  AND U39093 ( .A(n39208), .B(n39209), .Z(n39207) );
  XNOR U39094 ( .A(n39206), .B(n38904), .Z(n39209) );
  XOR U39095 ( .A(n38982), .B(n39210), .Z(n38904) );
  AND U39096 ( .A(n716), .B(n39211), .Z(n39210) );
  XOR U39097 ( .A(n38978), .B(n38982), .Z(n39211) );
  XOR U39098 ( .A(n38853), .B(n39206), .Z(n39208) );
  XOR U39099 ( .A(n39212), .B(n39213), .Z(n38853) );
  AND U39100 ( .A(n732), .B(n39214), .Z(n39213) );
  XOR U39101 ( .A(n39180), .B(n39215), .Z(n39206) );
  AND U39102 ( .A(n39216), .B(n39183), .Z(n39215) );
  XNOR U39103 ( .A(n38914), .B(n39180), .Z(n39183) );
  XOR U39104 ( .A(n39031), .B(n39217), .Z(n38914) );
  AND U39105 ( .A(n716), .B(n39218), .Z(n39217) );
  XOR U39106 ( .A(n39027), .B(n39031), .Z(n39218) );
  XNOR U39107 ( .A(n39219), .B(n39180), .Z(n39216) );
  IV U39108 ( .A(n38861), .Z(n39219) );
  XOR U39109 ( .A(n39220), .B(n39221), .Z(n38861) );
  AND U39110 ( .A(n732), .B(n39222), .Z(n39221) );
  XOR U39111 ( .A(n39223), .B(n39224), .Z(n39180) );
  AND U39112 ( .A(n39225), .B(n39226), .Z(n39224) );
  XNOR U39113 ( .A(n39223), .B(n38922), .Z(n39226) );
  XOR U39114 ( .A(n39124), .B(n39227), .Z(n38922) );
  AND U39115 ( .A(n716), .B(n39228), .Z(n39227) );
  XOR U39116 ( .A(n39120), .B(n39124), .Z(n39228) );
  XNOR U39117 ( .A(n39229), .B(n39223), .Z(n39225) );
  IV U39118 ( .A(n38871), .Z(n39229) );
  XOR U39119 ( .A(n39230), .B(n39231), .Z(n38871) );
  AND U39120 ( .A(n732), .B(n39232), .Z(n39231) );
  AND U39121 ( .A(n39184), .B(n39165), .Z(n39223) );
  XNOR U39122 ( .A(n39233), .B(n39234), .Z(n39165) );
  AND U39123 ( .A(n716), .B(n39143), .Z(n39234) );
  XNOR U39124 ( .A(n39141), .B(n39233), .Z(n39143) );
  XNOR U39125 ( .A(n39235), .B(n39236), .Z(n716) );
  AND U39126 ( .A(n39237), .B(n39238), .Z(n39236) );
  XNOR U39127 ( .A(n39235), .B(n38934), .Z(n39238) );
  IV U39128 ( .A(n38938), .Z(n38934) );
  XOR U39129 ( .A(n39239), .B(n39240), .Z(n38938) );
  AND U39130 ( .A(n720), .B(n39241), .Z(n39240) );
  XOR U39131 ( .A(n39242), .B(n39239), .Z(n39241) );
  XNOR U39132 ( .A(n39235), .B(n39148), .Z(n39237) );
  XOR U39133 ( .A(n39243), .B(n39244), .Z(n39148) );
  AND U39134 ( .A(n728), .B(n39195), .Z(n39244) );
  XOR U39135 ( .A(n39193), .B(n39243), .Z(n39195) );
  XOR U39136 ( .A(n39245), .B(n39246), .Z(n39235) );
  AND U39137 ( .A(n39247), .B(n39248), .Z(n39246) );
  XNOR U39138 ( .A(n39245), .B(n38950), .Z(n39248) );
  IV U39139 ( .A(n38953), .Z(n38950) );
  XOR U39140 ( .A(n39249), .B(n39250), .Z(n38953) );
  AND U39141 ( .A(n720), .B(n39251), .Z(n39250) );
  XOR U39142 ( .A(n39252), .B(n39249), .Z(n39251) );
  XOR U39143 ( .A(n38954), .B(n39245), .Z(n39247) );
  XOR U39144 ( .A(n39253), .B(n39254), .Z(n38954) );
  AND U39145 ( .A(n728), .B(n39205), .Z(n39254) );
  XOR U39146 ( .A(n39253), .B(n39203), .Z(n39205) );
  XOR U39147 ( .A(n39255), .B(n39256), .Z(n39245) );
  AND U39148 ( .A(n39257), .B(n39258), .Z(n39256) );
  XNOR U39149 ( .A(n39255), .B(n38978), .Z(n39258) );
  IV U39150 ( .A(n38981), .Z(n38978) );
  XOR U39151 ( .A(n39259), .B(n39260), .Z(n38981) );
  AND U39152 ( .A(n720), .B(n39261), .Z(n39260) );
  XNOR U39153 ( .A(n39262), .B(n39259), .Z(n39261) );
  XOR U39154 ( .A(n38982), .B(n39255), .Z(n39257) );
  XOR U39155 ( .A(n39263), .B(n39264), .Z(n38982) );
  AND U39156 ( .A(n728), .B(n39214), .Z(n39264) );
  XOR U39157 ( .A(n39263), .B(n39212), .Z(n39214) );
  XOR U39158 ( .A(n39265), .B(n39266), .Z(n39255) );
  AND U39159 ( .A(n39267), .B(n39268), .Z(n39266) );
  XNOR U39160 ( .A(n39265), .B(n39027), .Z(n39268) );
  IV U39161 ( .A(n39030), .Z(n39027) );
  XOR U39162 ( .A(n39269), .B(n39270), .Z(n39030) );
  AND U39163 ( .A(n720), .B(n39271), .Z(n39270) );
  XOR U39164 ( .A(n39272), .B(n39269), .Z(n39271) );
  XOR U39165 ( .A(n39031), .B(n39265), .Z(n39267) );
  XOR U39166 ( .A(n39273), .B(n39274), .Z(n39031) );
  AND U39167 ( .A(n728), .B(n39222), .Z(n39274) );
  XOR U39168 ( .A(n39273), .B(n39220), .Z(n39222) );
  XOR U39169 ( .A(n39161), .B(n39275), .Z(n39265) );
  AND U39170 ( .A(n39163), .B(n39276), .Z(n39275) );
  XNOR U39171 ( .A(n39161), .B(n39120), .Z(n39276) );
  IV U39172 ( .A(n39123), .Z(n39120) );
  XOR U39173 ( .A(n39277), .B(n39278), .Z(n39123) );
  AND U39174 ( .A(n720), .B(n39279), .Z(n39278) );
  XNOR U39175 ( .A(n39280), .B(n39277), .Z(n39279) );
  XOR U39176 ( .A(n39124), .B(n39161), .Z(n39163) );
  XOR U39177 ( .A(n39281), .B(n39282), .Z(n39124) );
  AND U39178 ( .A(n728), .B(n39232), .Z(n39282) );
  XOR U39179 ( .A(n39281), .B(n39230), .Z(n39232) );
  AND U39180 ( .A(n39233), .B(n39141), .Z(n39161) );
  XNOR U39181 ( .A(n39283), .B(n39284), .Z(n39141) );
  AND U39182 ( .A(n720), .B(n39285), .Z(n39284) );
  XNOR U39183 ( .A(n39286), .B(n39283), .Z(n39285) );
  XNOR U39184 ( .A(n39287), .B(n39288), .Z(n720) );
  AND U39185 ( .A(n39289), .B(n39290), .Z(n39288) );
  XOR U39186 ( .A(n39242), .B(n39287), .Z(n39290) );
  AND U39187 ( .A(n39291), .B(n39292), .Z(n39242) );
  XNOR U39188 ( .A(n39239), .B(n39287), .Z(n39289) );
  XNOR U39189 ( .A(n39293), .B(n39294), .Z(n39239) );
  AND U39190 ( .A(n724), .B(n39295), .Z(n39294) );
  XNOR U39191 ( .A(n39296), .B(n39297), .Z(n39295) );
  XOR U39192 ( .A(n39298), .B(n39299), .Z(n39287) );
  AND U39193 ( .A(n39300), .B(n39301), .Z(n39299) );
  XNOR U39194 ( .A(n39298), .B(n39291), .Z(n39301) );
  IV U39195 ( .A(n39252), .Z(n39291) );
  XOR U39196 ( .A(n39302), .B(n39303), .Z(n39252) );
  XOR U39197 ( .A(n39304), .B(n39292), .Z(n39303) );
  AND U39198 ( .A(n39262), .B(n39305), .Z(n39292) );
  AND U39199 ( .A(n39306), .B(n39307), .Z(n39304) );
  XOR U39200 ( .A(n39308), .B(n39302), .Z(n39306) );
  XNOR U39201 ( .A(n39249), .B(n39298), .Z(n39300) );
  XNOR U39202 ( .A(n39309), .B(n39310), .Z(n39249) );
  AND U39203 ( .A(n724), .B(n39311), .Z(n39310) );
  XNOR U39204 ( .A(n39312), .B(n39313), .Z(n39311) );
  XOR U39205 ( .A(n39314), .B(n39315), .Z(n39298) );
  AND U39206 ( .A(n39316), .B(n39317), .Z(n39315) );
  XNOR U39207 ( .A(n39314), .B(n39262), .Z(n39317) );
  XOR U39208 ( .A(n39318), .B(n39307), .Z(n39262) );
  XNOR U39209 ( .A(n39319), .B(n39302), .Z(n39307) );
  XOR U39210 ( .A(n39320), .B(n39321), .Z(n39302) );
  AND U39211 ( .A(n39322), .B(n39323), .Z(n39321) );
  XOR U39212 ( .A(n39324), .B(n39320), .Z(n39322) );
  XNOR U39213 ( .A(n39325), .B(n39326), .Z(n39319) );
  AND U39214 ( .A(n39327), .B(n39328), .Z(n39326) );
  XOR U39215 ( .A(n39325), .B(n39329), .Z(n39327) );
  XNOR U39216 ( .A(n39308), .B(n39305), .Z(n39318) );
  AND U39217 ( .A(n39330), .B(n39331), .Z(n39305) );
  XOR U39218 ( .A(n39332), .B(n39333), .Z(n39308) );
  AND U39219 ( .A(n39334), .B(n39335), .Z(n39333) );
  XOR U39220 ( .A(n39332), .B(n39336), .Z(n39334) );
  XNOR U39221 ( .A(n39259), .B(n39314), .Z(n39316) );
  XNOR U39222 ( .A(n39337), .B(n39338), .Z(n39259) );
  AND U39223 ( .A(n724), .B(n39339), .Z(n39338) );
  XNOR U39224 ( .A(n39340), .B(n39341), .Z(n39339) );
  XOR U39225 ( .A(n39342), .B(n39343), .Z(n39314) );
  AND U39226 ( .A(n39344), .B(n39345), .Z(n39343) );
  XNOR U39227 ( .A(n39342), .B(n39330), .Z(n39345) );
  IV U39228 ( .A(n39272), .Z(n39330) );
  XNOR U39229 ( .A(n39346), .B(n39323), .Z(n39272) );
  XNOR U39230 ( .A(n39347), .B(n39329), .Z(n39323) );
  XOR U39231 ( .A(n39348), .B(n39349), .Z(n39329) );
  AND U39232 ( .A(n39350), .B(n39351), .Z(n39349) );
  XOR U39233 ( .A(n39348), .B(n39352), .Z(n39350) );
  XNOR U39234 ( .A(n39328), .B(n39320), .Z(n39347) );
  XOR U39235 ( .A(n39353), .B(n39354), .Z(n39320) );
  AND U39236 ( .A(n39355), .B(n39356), .Z(n39354) );
  XNOR U39237 ( .A(n39357), .B(n39353), .Z(n39355) );
  XNOR U39238 ( .A(n39358), .B(n39325), .Z(n39328) );
  XOR U39239 ( .A(n39359), .B(n39360), .Z(n39325) );
  AND U39240 ( .A(n39361), .B(n39362), .Z(n39360) );
  XOR U39241 ( .A(n39359), .B(n39363), .Z(n39361) );
  XNOR U39242 ( .A(n39364), .B(n39365), .Z(n39358) );
  AND U39243 ( .A(n39366), .B(n39367), .Z(n39365) );
  XNOR U39244 ( .A(n39364), .B(n39368), .Z(n39366) );
  XNOR U39245 ( .A(n39324), .B(n39331), .Z(n39346) );
  AND U39246 ( .A(n39280), .B(n39369), .Z(n39331) );
  XOR U39247 ( .A(n39336), .B(n39335), .Z(n39324) );
  XNOR U39248 ( .A(n39370), .B(n39332), .Z(n39335) );
  XOR U39249 ( .A(n39371), .B(n39372), .Z(n39332) );
  AND U39250 ( .A(n39373), .B(n39374), .Z(n39372) );
  XOR U39251 ( .A(n39371), .B(n39375), .Z(n39373) );
  XNOR U39252 ( .A(n39376), .B(n39377), .Z(n39370) );
  AND U39253 ( .A(n39378), .B(n39379), .Z(n39377) );
  XOR U39254 ( .A(n39376), .B(n39380), .Z(n39378) );
  XOR U39255 ( .A(n39381), .B(n39382), .Z(n39336) );
  AND U39256 ( .A(n39383), .B(n39384), .Z(n39382) );
  XOR U39257 ( .A(n39381), .B(n39385), .Z(n39383) );
  XNOR U39258 ( .A(n39269), .B(n39342), .Z(n39344) );
  XNOR U39259 ( .A(n39386), .B(n39387), .Z(n39269) );
  AND U39260 ( .A(n724), .B(n39388), .Z(n39387) );
  XNOR U39261 ( .A(n39389), .B(n39390), .Z(n39388) );
  XOR U39262 ( .A(n39391), .B(n39392), .Z(n39342) );
  AND U39263 ( .A(n39393), .B(n39394), .Z(n39392) );
  XNOR U39264 ( .A(n39391), .B(n39280), .Z(n39394) );
  XOR U39265 ( .A(n39395), .B(n39356), .Z(n39280) );
  XNOR U39266 ( .A(n39396), .B(n39363), .Z(n39356) );
  XOR U39267 ( .A(n39352), .B(n39351), .Z(n39363) );
  XNOR U39268 ( .A(n39397), .B(n39348), .Z(n39351) );
  XOR U39269 ( .A(n39398), .B(n39399), .Z(n39348) );
  AND U39270 ( .A(n39400), .B(n39401), .Z(n39399) );
  XNOR U39271 ( .A(n39402), .B(n39403), .Z(n39400) );
  IV U39272 ( .A(n39398), .Z(n39402) );
  XNOR U39273 ( .A(n39404), .B(n39405), .Z(n39397) );
  NOR U39274 ( .A(n39406), .B(n39407), .Z(n39405) );
  XNOR U39275 ( .A(n39404), .B(n39408), .Z(n39406) );
  XOR U39276 ( .A(n39409), .B(n39410), .Z(n39352) );
  NOR U39277 ( .A(n39411), .B(n39412), .Z(n39410) );
  XNOR U39278 ( .A(n39409), .B(n39413), .Z(n39411) );
  XNOR U39279 ( .A(n39362), .B(n39353), .Z(n39396) );
  XOR U39280 ( .A(n39414), .B(n39415), .Z(n39353) );
  AND U39281 ( .A(n39416), .B(n39417), .Z(n39415) );
  XOR U39282 ( .A(n39414), .B(n39418), .Z(n39416) );
  XOR U39283 ( .A(n39419), .B(n39368), .Z(n39362) );
  XOR U39284 ( .A(n39420), .B(n39421), .Z(n39368) );
  NOR U39285 ( .A(n39422), .B(n39423), .Z(n39421) );
  XOR U39286 ( .A(n39420), .B(n39424), .Z(n39422) );
  XNOR U39287 ( .A(n39367), .B(n39359), .Z(n39419) );
  XOR U39288 ( .A(n39425), .B(n39426), .Z(n39359) );
  AND U39289 ( .A(n39427), .B(n39428), .Z(n39426) );
  XOR U39290 ( .A(n39425), .B(n39429), .Z(n39427) );
  XNOR U39291 ( .A(n39430), .B(n39364), .Z(n39367) );
  XOR U39292 ( .A(n39431), .B(n39432), .Z(n39364) );
  AND U39293 ( .A(n39433), .B(n39434), .Z(n39432) );
  XNOR U39294 ( .A(n39435), .B(n39436), .Z(n39433) );
  IV U39295 ( .A(n39431), .Z(n39435) );
  XNOR U39296 ( .A(n39437), .B(n39438), .Z(n39430) );
  NOR U39297 ( .A(n39439), .B(n39440), .Z(n39438) );
  XNOR U39298 ( .A(n39437), .B(n39441), .Z(n39439) );
  XOR U39299 ( .A(n39357), .B(n39369), .Z(n39395) );
  NOR U39300 ( .A(n39286), .B(n39442), .Z(n39369) );
  XNOR U39301 ( .A(n39375), .B(n39374), .Z(n39357) );
  XNOR U39302 ( .A(n39443), .B(n39380), .Z(n39374) );
  XNOR U39303 ( .A(n39444), .B(n39445), .Z(n39380) );
  NOR U39304 ( .A(n39446), .B(n39447), .Z(n39445) );
  XOR U39305 ( .A(n39444), .B(n39448), .Z(n39446) );
  XNOR U39306 ( .A(n39379), .B(n39371), .Z(n39443) );
  XOR U39307 ( .A(n39449), .B(n39450), .Z(n39371) );
  AND U39308 ( .A(n39451), .B(n39452), .Z(n39450) );
  XOR U39309 ( .A(n39449), .B(n39453), .Z(n39451) );
  XNOR U39310 ( .A(n39454), .B(n39376), .Z(n39379) );
  XOR U39311 ( .A(n39455), .B(n39456), .Z(n39376) );
  AND U39312 ( .A(n39457), .B(n39458), .Z(n39456) );
  XNOR U39313 ( .A(n39459), .B(n39460), .Z(n39457) );
  IV U39314 ( .A(n39455), .Z(n39459) );
  XNOR U39315 ( .A(n39461), .B(n39462), .Z(n39454) );
  NOR U39316 ( .A(n39463), .B(n39464), .Z(n39462) );
  XNOR U39317 ( .A(n39461), .B(n39465), .Z(n39463) );
  XOR U39318 ( .A(n39385), .B(n39384), .Z(n39375) );
  XNOR U39319 ( .A(n39466), .B(n39381), .Z(n39384) );
  XOR U39320 ( .A(n39467), .B(n39468), .Z(n39381) );
  AND U39321 ( .A(n39469), .B(n39470), .Z(n39468) );
  XOR U39322 ( .A(n39467), .B(n39471), .Z(n39469) );
  XNOR U39323 ( .A(n39472), .B(n39473), .Z(n39466) );
  NOR U39324 ( .A(n39474), .B(n39475), .Z(n39473) );
  XNOR U39325 ( .A(n39472), .B(n39476), .Z(n39474) );
  XOR U39326 ( .A(n39477), .B(n39478), .Z(n39385) );
  NOR U39327 ( .A(n39479), .B(n39480), .Z(n39478) );
  XNOR U39328 ( .A(n39477), .B(n39481), .Z(n39479) );
  XNOR U39329 ( .A(n39277), .B(n39391), .Z(n39393) );
  XNOR U39330 ( .A(n39482), .B(n39483), .Z(n39277) );
  AND U39331 ( .A(n724), .B(n39484), .Z(n39483) );
  XNOR U39332 ( .A(n39485), .B(n39486), .Z(n39484) );
  AND U39333 ( .A(n39283), .B(n39286), .Z(n39391) );
  XOR U39334 ( .A(n39487), .B(n39442), .Z(n39286) );
  XNOR U39335 ( .A(p_input[2048]), .B(p_input[992]), .Z(n39442) );
  XNOR U39336 ( .A(n39418), .B(n39417), .Z(n39487) );
  XNOR U39337 ( .A(n39488), .B(n39429), .Z(n39417) );
  XOR U39338 ( .A(n39403), .B(n39401), .Z(n39429) );
  XNOR U39339 ( .A(n39489), .B(n39408), .Z(n39401) );
  XOR U39340 ( .A(p_input[1016]), .B(p_input[2072]), .Z(n39408) );
  XOR U39341 ( .A(n39398), .B(n39407), .Z(n39489) );
  XOR U39342 ( .A(n39490), .B(n39404), .Z(n39407) );
  XOR U39343 ( .A(p_input[1014]), .B(p_input[2070]), .Z(n39404) );
  XOR U39344 ( .A(p_input[1015]), .B(n29410), .Z(n39490) );
  XOR U39345 ( .A(p_input[1010]), .B(p_input[2066]), .Z(n39398) );
  XNOR U39346 ( .A(n39413), .B(n39412), .Z(n39403) );
  XOR U39347 ( .A(n39491), .B(n39409), .Z(n39412) );
  XOR U39348 ( .A(p_input[1011]), .B(p_input[2067]), .Z(n39409) );
  XOR U39349 ( .A(p_input[1012]), .B(n29412), .Z(n39491) );
  XOR U39350 ( .A(p_input[1013]), .B(p_input[2069]), .Z(n39413) );
  XNOR U39351 ( .A(n39428), .B(n39414), .Z(n39488) );
  XNOR U39352 ( .A(n28686), .B(p_input[993]), .Z(n39414) );
  XNOR U39353 ( .A(n39492), .B(n39436), .Z(n39428) );
  XNOR U39354 ( .A(n39424), .B(n39423), .Z(n39436) );
  XNOR U39355 ( .A(n39493), .B(n39420), .Z(n39423) );
  XNOR U39356 ( .A(p_input[1018]), .B(p_input[2074]), .Z(n39420) );
  XOR U39357 ( .A(p_input[1019]), .B(n29415), .Z(n39493) );
  XOR U39358 ( .A(p_input[1020]), .B(p_input[2076]), .Z(n39424) );
  XOR U39359 ( .A(n39434), .B(n39494), .Z(n39492) );
  IV U39360 ( .A(n39425), .Z(n39494) );
  XOR U39361 ( .A(p_input[1009]), .B(p_input[2065]), .Z(n39425) );
  XNOR U39362 ( .A(n39495), .B(n39441), .Z(n39434) );
  XNOR U39363 ( .A(p_input[1023]), .B(n29418), .Z(n39441) );
  XOR U39364 ( .A(n39431), .B(n39440), .Z(n39495) );
  XOR U39365 ( .A(n39496), .B(n39437), .Z(n39440) );
  XOR U39366 ( .A(p_input[1021]), .B(p_input[2077]), .Z(n39437) );
  XOR U39367 ( .A(p_input[1022]), .B(n29420), .Z(n39496) );
  XOR U39368 ( .A(p_input[1017]), .B(p_input[2073]), .Z(n39431) );
  XOR U39369 ( .A(n39453), .B(n39452), .Z(n39418) );
  XNOR U39370 ( .A(n39497), .B(n39460), .Z(n39452) );
  XNOR U39371 ( .A(n39448), .B(n39447), .Z(n39460) );
  XNOR U39372 ( .A(n39498), .B(n39444), .Z(n39447) );
  XNOR U39373 ( .A(p_input[1003]), .B(p_input[2059]), .Z(n39444) );
  XOR U39374 ( .A(p_input[1004]), .B(n28329), .Z(n39498) );
  XOR U39375 ( .A(p_input[1005]), .B(p_input[2061]), .Z(n39448) );
  XNOR U39376 ( .A(n39458), .B(n39449), .Z(n39497) );
  XNOR U39377 ( .A(n28330), .B(p_input[994]), .Z(n39449) );
  XNOR U39378 ( .A(n39499), .B(n39465), .Z(n39458) );
  XNOR U39379 ( .A(p_input[1008]), .B(n28332), .Z(n39465) );
  XOR U39380 ( .A(n39455), .B(n39464), .Z(n39499) );
  XOR U39381 ( .A(n39500), .B(n39461), .Z(n39464) );
  XOR U39382 ( .A(p_input[1006]), .B(p_input[2062]), .Z(n39461) );
  XOR U39383 ( .A(p_input[1007]), .B(n28334), .Z(n39500) );
  XOR U39384 ( .A(p_input[1002]), .B(p_input[2058]), .Z(n39455) );
  XOR U39385 ( .A(n39471), .B(n39470), .Z(n39453) );
  XNOR U39386 ( .A(n39501), .B(n39476), .Z(n39470) );
  XOR U39387 ( .A(p_input[1001]), .B(p_input[2057]), .Z(n39476) );
  XOR U39388 ( .A(n39467), .B(n39475), .Z(n39501) );
  XOR U39389 ( .A(n39502), .B(n39472), .Z(n39475) );
  XOR U39390 ( .A(p_input[2055]), .B(p_input[999]), .Z(n39472) );
  XOR U39391 ( .A(p_input[1000]), .B(n29427), .Z(n39502) );
  XNOR U39392 ( .A(n28337), .B(p_input[995]), .Z(n39467) );
  XNOR U39393 ( .A(n39481), .B(n39480), .Z(n39471) );
  XOR U39394 ( .A(n39503), .B(n39477), .Z(n39480) );
  XOR U39395 ( .A(p_input[2052]), .B(p_input[996]), .Z(n39477) );
  XNOR U39396 ( .A(p_input[2053]), .B(p_input[997]), .Z(n39503) );
  XOR U39397 ( .A(p_input[2054]), .B(p_input[998]), .Z(n39481) );
  XNOR U39398 ( .A(n39504), .B(n39505), .Z(n39283) );
  AND U39399 ( .A(n724), .B(n39506), .Z(n39505) );
  XNOR U39400 ( .A(n39507), .B(n39508), .Z(n724) );
  AND U39401 ( .A(n39509), .B(n39510), .Z(n39508) );
  XOR U39402 ( .A(n39297), .B(n39507), .Z(n39510) );
  XNOR U39403 ( .A(n39511), .B(n39507), .Z(n39509) );
  XOR U39404 ( .A(n39512), .B(n39513), .Z(n39507) );
  AND U39405 ( .A(n39514), .B(n39515), .Z(n39513) );
  XOR U39406 ( .A(n39312), .B(n39512), .Z(n39515) );
  XOR U39407 ( .A(n39512), .B(n39313), .Z(n39514) );
  XOR U39408 ( .A(n39516), .B(n39517), .Z(n39512) );
  AND U39409 ( .A(n39518), .B(n39519), .Z(n39517) );
  XOR U39410 ( .A(n39340), .B(n39516), .Z(n39519) );
  XOR U39411 ( .A(n39516), .B(n39341), .Z(n39518) );
  XOR U39412 ( .A(n39520), .B(n39521), .Z(n39516) );
  AND U39413 ( .A(n39522), .B(n39523), .Z(n39521) );
  XOR U39414 ( .A(n39389), .B(n39520), .Z(n39523) );
  XOR U39415 ( .A(n39520), .B(n39390), .Z(n39522) );
  XOR U39416 ( .A(n39524), .B(n39525), .Z(n39520) );
  AND U39417 ( .A(n39526), .B(n39527), .Z(n39525) );
  XOR U39418 ( .A(n39524), .B(n39485), .Z(n39527) );
  XNOR U39419 ( .A(n39528), .B(n39529), .Z(n39233) );
  AND U39420 ( .A(n728), .B(n39530), .Z(n39529) );
  XNOR U39421 ( .A(n39531), .B(n39532), .Z(n728) );
  AND U39422 ( .A(n39533), .B(n39534), .Z(n39532) );
  XOR U39423 ( .A(n39531), .B(n39243), .Z(n39534) );
  XNOR U39424 ( .A(n39531), .B(n39193), .Z(n39533) );
  XOR U39425 ( .A(n39535), .B(n39536), .Z(n39531) );
  AND U39426 ( .A(n39537), .B(n39538), .Z(n39536) );
  XNOR U39427 ( .A(n39253), .B(n39535), .Z(n39538) );
  XOR U39428 ( .A(n39535), .B(n39203), .Z(n39537) );
  XOR U39429 ( .A(n39539), .B(n39540), .Z(n39535) );
  AND U39430 ( .A(n39541), .B(n39542), .Z(n39540) );
  XNOR U39431 ( .A(n39263), .B(n39539), .Z(n39542) );
  XOR U39432 ( .A(n39539), .B(n39212), .Z(n39541) );
  XOR U39433 ( .A(n39543), .B(n39544), .Z(n39539) );
  AND U39434 ( .A(n39545), .B(n39546), .Z(n39544) );
  XOR U39435 ( .A(n39543), .B(n39220), .Z(n39545) );
  XOR U39436 ( .A(n39547), .B(n39548), .Z(n39184) );
  AND U39437 ( .A(n732), .B(n39530), .Z(n39548) );
  XNOR U39438 ( .A(n39528), .B(n39547), .Z(n39530) );
  XNOR U39439 ( .A(n39549), .B(n39550), .Z(n732) );
  AND U39440 ( .A(n39551), .B(n39552), .Z(n39550) );
  XNOR U39441 ( .A(n39553), .B(n39549), .Z(n39552) );
  IV U39442 ( .A(n39243), .Z(n39553) );
  XOR U39443 ( .A(n39511), .B(n39554), .Z(n39243) );
  AND U39444 ( .A(n735), .B(n39555), .Z(n39554) );
  XOR U39445 ( .A(n39296), .B(n39293), .Z(n39555) );
  IV U39446 ( .A(n39511), .Z(n39296) );
  XNOR U39447 ( .A(n39193), .B(n39549), .Z(n39551) );
  XOR U39448 ( .A(n39556), .B(n39557), .Z(n39193) );
  AND U39449 ( .A(n751), .B(n39558), .Z(n39557) );
  XOR U39450 ( .A(n39559), .B(n39560), .Z(n39549) );
  AND U39451 ( .A(n39561), .B(n39562), .Z(n39560) );
  XNOR U39452 ( .A(n39559), .B(n39253), .Z(n39562) );
  XOR U39453 ( .A(n39313), .B(n39563), .Z(n39253) );
  AND U39454 ( .A(n735), .B(n39564), .Z(n39563) );
  XOR U39455 ( .A(n39309), .B(n39313), .Z(n39564) );
  XNOR U39456 ( .A(n39565), .B(n39559), .Z(n39561) );
  IV U39457 ( .A(n39203), .Z(n39565) );
  XOR U39458 ( .A(n39566), .B(n39567), .Z(n39203) );
  AND U39459 ( .A(n751), .B(n39568), .Z(n39567) );
  XOR U39460 ( .A(n39569), .B(n39570), .Z(n39559) );
  AND U39461 ( .A(n39571), .B(n39572), .Z(n39570) );
  XNOR U39462 ( .A(n39569), .B(n39263), .Z(n39572) );
  XOR U39463 ( .A(n39341), .B(n39573), .Z(n39263) );
  AND U39464 ( .A(n735), .B(n39574), .Z(n39573) );
  XOR U39465 ( .A(n39337), .B(n39341), .Z(n39574) );
  XOR U39466 ( .A(n39212), .B(n39569), .Z(n39571) );
  XOR U39467 ( .A(n39575), .B(n39576), .Z(n39212) );
  AND U39468 ( .A(n751), .B(n39577), .Z(n39576) );
  XOR U39469 ( .A(n39543), .B(n39578), .Z(n39569) );
  AND U39470 ( .A(n39579), .B(n39546), .Z(n39578) );
  XNOR U39471 ( .A(n39273), .B(n39543), .Z(n39546) );
  XOR U39472 ( .A(n39390), .B(n39580), .Z(n39273) );
  AND U39473 ( .A(n735), .B(n39581), .Z(n39580) );
  XOR U39474 ( .A(n39386), .B(n39390), .Z(n39581) );
  XNOR U39475 ( .A(n39582), .B(n39543), .Z(n39579) );
  IV U39476 ( .A(n39220), .Z(n39582) );
  XOR U39477 ( .A(n39583), .B(n39584), .Z(n39220) );
  AND U39478 ( .A(n751), .B(n39585), .Z(n39584) );
  XOR U39479 ( .A(n39586), .B(n39587), .Z(n39543) );
  AND U39480 ( .A(n39588), .B(n39589), .Z(n39587) );
  XNOR U39481 ( .A(n39586), .B(n39281), .Z(n39589) );
  XOR U39482 ( .A(n39486), .B(n39590), .Z(n39281) );
  AND U39483 ( .A(n735), .B(n39591), .Z(n39590) );
  XOR U39484 ( .A(n39482), .B(n39486), .Z(n39591) );
  XNOR U39485 ( .A(n39592), .B(n39586), .Z(n39588) );
  IV U39486 ( .A(n39230), .Z(n39592) );
  XOR U39487 ( .A(n39593), .B(n39594), .Z(n39230) );
  AND U39488 ( .A(n751), .B(n39595), .Z(n39594) );
  AND U39489 ( .A(n39547), .B(n39528), .Z(n39586) );
  XNOR U39490 ( .A(n39596), .B(n39597), .Z(n39528) );
  AND U39491 ( .A(n735), .B(n39506), .Z(n39597) );
  XNOR U39492 ( .A(n39504), .B(n39596), .Z(n39506) );
  XNOR U39493 ( .A(n39598), .B(n39599), .Z(n735) );
  AND U39494 ( .A(n39600), .B(n39601), .Z(n39599) );
  XNOR U39495 ( .A(n39598), .B(n39293), .Z(n39601) );
  IV U39496 ( .A(n39297), .Z(n39293) );
  XOR U39497 ( .A(n39602), .B(n39603), .Z(n39297) );
  AND U39498 ( .A(n739), .B(n39604), .Z(n39603) );
  XOR U39499 ( .A(n39605), .B(n39602), .Z(n39604) );
  XNOR U39500 ( .A(n39598), .B(n39511), .Z(n39600) );
  XOR U39501 ( .A(n39606), .B(n39607), .Z(n39511) );
  AND U39502 ( .A(n747), .B(n39558), .Z(n39607) );
  XOR U39503 ( .A(n39556), .B(n39606), .Z(n39558) );
  XOR U39504 ( .A(n39608), .B(n39609), .Z(n39598) );
  AND U39505 ( .A(n39610), .B(n39611), .Z(n39609) );
  XNOR U39506 ( .A(n39608), .B(n39309), .Z(n39611) );
  IV U39507 ( .A(n39312), .Z(n39309) );
  XOR U39508 ( .A(n39612), .B(n39613), .Z(n39312) );
  AND U39509 ( .A(n739), .B(n39614), .Z(n39613) );
  XOR U39510 ( .A(n39615), .B(n39612), .Z(n39614) );
  XOR U39511 ( .A(n39313), .B(n39608), .Z(n39610) );
  XOR U39512 ( .A(n39616), .B(n39617), .Z(n39313) );
  AND U39513 ( .A(n747), .B(n39568), .Z(n39617) );
  XOR U39514 ( .A(n39616), .B(n39566), .Z(n39568) );
  XOR U39515 ( .A(n39618), .B(n39619), .Z(n39608) );
  AND U39516 ( .A(n39620), .B(n39621), .Z(n39619) );
  XNOR U39517 ( .A(n39618), .B(n39337), .Z(n39621) );
  IV U39518 ( .A(n39340), .Z(n39337) );
  XOR U39519 ( .A(n39622), .B(n39623), .Z(n39340) );
  AND U39520 ( .A(n739), .B(n39624), .Z(n39623) );
  XNOR U39521 ( .A(n39625), .B(n39622), .Z(n39624) );
  XOR U39522 ( .A(n39341), .B(n39618), .Z(n39620) );
  XOR U39523 ( .A(n39626), .B(n39627), .Z(n39341) );
  AND U39524 ( .A(n747), .B(n39577), .Z(n39627) );
  XOR U39525 ( .A(n39626), .B(n39575), .Z(n39577) );
  XOR U39526 ( .A(n39628), .B(n39629), .Z(n39618) );
  AND U39527 ( .A(n39630), .B(n39631), .Z(n39629) );
  XNOR U39528 ( .A(n39628), .B(n39386), .Z(n39631) );
  IV U39529 ( .A(n39389), .Z(n39386) );
  XOR U39530 ( .A(n39632), .B(n39633), .Z(n39389) );
  AND U39531 ( .A(n739), .B(n39634), .Z(n39633) );
  XOR U39532 ( .A(n39635), .B(n39632), .Z(n39634) );
  XOR U39533 ( .A(n39390), .B(n39628), .Z(n39630) );
  XOR U39534 ( .A(n39636), .B(n39637), .Z(n39390) );
  AND U39535 ( .A(n747), .B(n39585), .Z(n39637) );
  XOR U39536 ( .A(n39636), .B(n39583), .Z(n39585) );
  XOR U39537 ( .A(n39524), .B(n39638), .Z(n39628) );
  AND U39538 ( .A(n39526), .B(n39639), .Z(n39638) );
  XNOR U39539 ( .A(n39524), .B(n39482), .Z(n39639) );
  IV U39540 ( .A(n39485), .Z(n39482) );
  XOR U39541 ( .A(n39640), .B(n39641), .Z(n39485) );
  AND U39542 ( .A(n739), .B(n39642), .Z(n39641) );
  XNOR U39543 ( .A(n39643), .B(n39640), .Z(n39642) );
  XOR U39544 ( .A(n39486), .B(n39524), .Z(n39526) );
  XOR U39545 ( .A(n39644), .B(n39645), .Z(n39486) );
  AND U39546 ( .A(n747), .B(n39595), .Z(n39645) );
  XOR U39547 ( .A(n39644), .B(n39593), .Z(n39595) );
  AND U39548 ( .A(n39596), .B(n39504), .Z(n39524) );
  XNOR U39549 ( .A(n39646), .B(n39647), .Z(n39504) );
  AND U39550 ( .A(n739), .B(n39648), .Z(n39647) );
  XNOR U39551 ( .A(n39649), .B(n39646), .Z(n39648) );
  XNOR U39552 ( .A(n39650), .B(n39651), .Z(n739) );
  AND U39553 ( .A(n39652), .B(n39653), .Z(n39651) );
  XOR U39554 ( .A(n39605), .B(n39650), .Z(n39653) );
  AND U39555 ( .A(n39654), .B(n39655), .Z(n39605) );
  XNOR U39556 ( .A(n39602), .B(n39650), .Z(n39652) );
  XNOR U39557 ( .A(n39656), .B(n39657), .Z(n39602) );
  AND U39558 ( .A(n743), .B(n39658), .Z(n39657) );
  XNOR U39559 ( .A(n39659), .B(n39660), .Z(n39658) );
  XOR U39560 ( .A(n39661), .B(n39662), .Z(n39650) );
  AND U39561 ( .A(n39663), .B(n39664), .Z(n39662) );
  XNOR U39562 ( .A(n39661), .B(n39654), .Z(n39664) );
  IV U39563 ( .A(n39615), .Z(n39654) );
  XOR U39564 ( .A(n39665), .B(n39666), .Z(n39615) );
  XOR U39565 ( .A(n39667), .B(n39655), .Z(n39666) );
  AND U39566 ( .A(n39625), .B(n39668), .Z(n39655) );
  AND U39567 ( .A(n39669), .B(n39670), .Z(n39667) );
  XOR U39568 ( .A(n39671), .B(n39665), .Z(n39669) );
  XNOR U39569 ( .A(n39612), .B(n39661), .Z(n39663) );
  XNOR U39570 ( .A(n39672), .B(n39673), .Z(n39612) );
  AND U39571 ( .A(n743), .B(n39674), .Z(n39673) );
  XNOR U39572 ( .A(n39675), .B(n39676), .Z(n39674) );
  XOR U39573 ( .A(n39677), .B(n39678), .Z(n39661) );
  AND U39574 ( .A(n39679), .B(n39680), .Z(n39678) );
  XNOR U39575 ( .A(n39677), .B(n39625), .Z(n39680) );
  XOR U39576 ( .A(n39681), .B(n39670), .Z(n39625) );
  XNOR U39577 ( .A(n39682), .B(n39665), .Z(n39670) );
  XOR U39578 ( .A(n39683), .B(n39684), .Z(n39665) );
  AND U39579 ( .A(n39685), .B(n39686), .Z(n39684) );
  XOR U39580 ( .A(n39687), .B(n39683), .Z(n39685) );
  XNOR U39581 ( .A(n39688), .B(n39689), .Z(n39682) );
  AND U39582 ( .A(n39690), .B(n39691), .Z(n39689) );
  XOR U39583 ( .A(n39688), .B(n39692), .Z(n39690) );
  XNOR U39584 ( .A(n39671), .B(n39668), .Z(n39681) );
  AND U39585 ( .A(n39693), .B(n39694), .Z(n39668) );
  XOR U39586 ( .A(n39695), .B(n39696), .Z(n39671) );
  AND U39587 ( .A(n39697), .B(n39698), .Z(n39696) );
  XOR U39588 ( .A(n39695), .B(n39699), .Z(n39697) );
  XNOR U39589 ( .A(n39622), .B(n39677), .Z(n39679) );
  XNOR U39590 ( .A(n39700), .B(n39701), .Z(n39622) );
  AND U39591 ( .A(n743), .B(n39702), .Z(n39701) );
  XNOR U39592 ( .A(n39703), .B(n39704), .Z(n39702) );
  XOR U39593 ( .A(n39705), .B(n39706), .Z(n39677) );
  AND U39594 ( .A(n39707), .B(n39708), .Z(n39706) );
  XNOR U39595 ( .A(n39705), .B(n39693), .Z(n39708) );
  IV U39596 ( .A(n39635), .Z(n39693) );
  XNOR U39597 ( .A(n39709), .B(n39686), .Z(n39635) );
  XNOR U39598 ( .A(n39710), .B(n39692), .Z(n39686) );
  XOR U39599 ( .A(n39711), .B(n39712), .Z(n39692) );
  AND U39600 ( .A(n39713), .B(n39714), .Z(n39712) );
  XOR U39601 ( .A(n39711), .B(n39715), .Z(n39713) );
  XNOR U39602 ( .A(n39691), .B(n39683), .Z(n39710) );
  XOR U39603 ( .A(n39716), .B(n39717), .Z(n39683) );
  AND U39604 ( .A(n39718), .B(n39719), .Z(n39717) );
  XNOR U39605 ( .A(n39720), .B(n39716), .Z(n39718) );
  XNOR U39606 ( .A(n39721), .B(n39688), .Z(n39691) );
  XOR U39607 ( .A(n39722), .B(n39723), .Z(n39688) );
  AND U39608 ( .A(n39724), .B(n39725), .Z(n39723) );
  XOR U39609 ( .A(n39722), .B(n39726), .Z(n39724) );
  XNOR U39610 ( .A(n39727), .B(n39728), .Z(n39721) );
  AND U39611 ( .A(n39729), .B(n39730), .Z(n39728) );
  XNOR U39612 ( .A(n39727), .B(n39731), .Z(n39729) );
  XNOR U39613 ( .A(n39687), .B(n39694), .Z(n39709) );
  AND U39614 ( .A(n39643), .B(n39732), .Z(n39694) );
  XOR U39615 ( .A(n39699), .B(n39698), .Z(n39687) );
  XNOR U39616 ( .A(n39733), .B(n39695), .Z(n39698) );
  XOR U39617 ( .A(n39734), .B(n39735), .Z(n39695) );
  AND U39618 ( .A(n39736), .B(n39737), .Z(n39735) );
  XOR U39619 ( .A(n39734), .B(n39738), .Z(n39736) );
  XNOR U39620 ( .A(n39739), .B(n39740), .Z(n39733) );
  AND U39621 ( .A(n39741), .B(n39742), .Z(n39740) );
  XOR U39622 ( .A(n39739), .B(n39743), .Z(n39741) );
  XOR U39623 ( .A(n39744), .B(n39745), .Z(n39699) );
  AND U39624 ( .A(n39746), .B(n39747), .Z(n39745) );
  XOR U39625 ( .A(n39744), .B(n39748), .Z(n39746) );
  XNOR U39626 ( .A(n39632), .B(n39705), .Z(n39707) );
  XNOR U39627 ( .A(n39749), .B(n39750), .Z(n39632) );
  AND U39628 ( .A(n743), .B(n39751), .Z(n39750) );
  XNOR U39629 ( .A(n39752), .B(n39753), .Z(n39751) );
  XOR U39630 ( .A(n39754), .B(n39755), .Z(n39705) );
  AND U39631 ( .A(n39756), .B(n39757), .Z(n39755) );
  XNOR U39632 ( .A(n39754), .B(n39643), .Z(n39757) );
  XOR U39633 ( .A(n39758), .B(n39719), .Z(n39643) );
  XNOR U39634 ( .A(n39759), .B(n39726), .Z(n39719) );
  XOR U39635 ( .A(n39715), .B(n39714), .Z(n39726) );
  XNOR U39636 ( .A(n39760), .B(n39711), .Z(n39714) );
  XOR U39637 ( .A(n39761), .B(n39762), .Z(n39711) );
  AND U39638 ( .A(n39763), .B(n39764), .Z(n39762) );
  XNOR U39639 ( .A(n39765), .B(n39766), .Z(n39763) );
  IV U39640 ( .A(n39761), .Z(n39765) );
  XNOR U39641 ( .A(n39767), .B(n39768), .Z(n39760) );
  NOR U39642 ( .A(n39769), .B(n39770), .Z(n39768) );
  XNOR U39643 ( .A(n39767), .B(n39771), .Z(n39769) );
  XOR U39644 ( .A(n39772), .B(n39773), .Z(n39715) );
  NOR U39645 ( .A(n39774), .B(n39775), .Z(n39773) );
  XNOR U39646 ( .A(n39772), .B(n39776), .Z(n39774) );
  XNOR U39647 ( .A(n39725), .B(n39716), .Z(n39759) );
  XOR U39648 ( .A(n39777), .B(n39778), .Z(n39716) );
  AND U39649 ( .A(n39779), .B(n39780), .Z(n39778) );
  XOR U39650 ( .A(n39777), .B(n39781), .Z(n39779) );
  XOR U39651 ( .A(n39782), .B(n39731), .Z(n39725) );
  XOR U39652 ( .A(n39783), .B(n39784), .Z(n39731) );
  NOR U39653 ( .A(n39785), .B(n39786), .Z(n39784) );
  XOR U39654 ( .A(n39783), .B(n39787), .Z(n39785) );
  XNOR U39655 ( .A(n39730), .B(n39722), .Z(n39782) );
  XOR U39656 ( .A(n39788), .B(n39789), .Z(n39722) );
  AND U39657 ( .A(n39790), .B(n39791), .Z(n39789) );
  XOR U39658 ( .A(n39788), .B(n39792), .Z(n39790) );
  XNOR U39659 ( .A(n39793), .B(n39727), .Z(n39730) );
  XOR U39660 ( .A(n39794), .B(n39795), .Z(n39727) );
  AND U39661 ( .A(n39796), .B(n39797), .Z(n39795) );
  XNOR U39662 ( .A(n39798), .B(n39799), .Z(n39796) );
  IV U39663 ( .A(n39794), .Z(n39798) );
  XNOR U39664 ( .A(n39800), .B(n39801), .Z(n39793) );
  NOR U39665 ( .A(n39802), .B(n39803), .Z(n39801) );
  XNOR U39666 ( .A(n39800), .B(n39804), .Z(n39802) );
  XOR U39667 ( .A(n39720), .B(n39732), .Z(n39758) );
  NOR U39668 ( .A(n39649), .B(n39805), .Z(n39732) );
  XNOR U39669 ( .A(n39738), .B(n39737), .Z(n39720) );
  XNOR U39670 ( .A(n39806), .B(n39743), .Z(n39737) );
  XNOR U39671 ( .A(n39807), .B(n39808), .Z(n39743) );
  NOR U39672 ( .A(n39809), .B(n39810), .Z(n39808) );
  XOR U39673 ( .A(n39807), .B(n39811), .Z(n39809) );
  XNOR U39674 ( .A(n39742), .B(n39734), .Z(n39806) );
  XOR U39675 ( .A(n39812), .B(n39813), .Z(n39734) );
  AND U39676 ( .A(n39814), .B(n39815), .Z(n39813) );
  XOR U39677 ( .A(n39812), .B(n39816), .Z(n39814) );
  XNOR U39678 ( .A(n39817), .B(n39739), .Z(n39742) );
  XOR U39679 ( .A(n39818), .B(n39819), .Z(n39739) );
  AND U39680 ( .A(n39820), .B(n39821), .Z(n39819) );
  XNOR U39681 ( .A(n39822), .B(n39823), .Z(n39820) );
  IV U39682 ( .A(n39818), .Z(n39822) );
  XNOR U39683 ( .A(n39824), .B(n39825), .Z(n39817) );
  NOR U39684 ( .A(n39826), .B(n39827), .Z(n39825) );
  XNOR U39685 ( .A(n39824), .B(n39828), .Z(n39826) );
  XOR U39686 ( .A(n39748), .B(n39747), .Z(n39738) );
  XNOR U39687 ( .A(n39829), .B(n39744), .Z(n39747) );
  XOR U39688 ( .A(n39830), .B(n39831), .Z(n39744) );
  AND U39689 ( .A(n39832), .B(n39833), .Z(n39831) );
  XNOR U39690 ( .A(n39834), .B(n39835), .Z(n39832) );
  IV U39691 ( .A(n39830), .Z(n39834) );
  XNOR U39692 ( .A(n39836), .B(n39837), .Z(n39829) );
  NOR U39693 ( .A(n39838), .B(n39839), .Z(n39837) );
  XNOR U39694 ( .A(n39836), .B(n39840), .Z(n39838) );
  XOR U39695 ( .A(n39841), .B(n39842), .Z(n39748) );
  NOR U39696 ( .A(n39843), .B(n39844), .Z(n39842) );
  XNOR U39697 ( .A(n39841), .B(n39845), .Z(n39843) );
  XNOR U39698 ( .A(n39640), .B(n39754), .Z(n39756) );
  XNOR U39699 ( .A(n39846), .B(n39847), .Z(n39640) );
  AND U39700 ( .A(n743), .B(n39848), .Z(n39847) );
  XNOR U39701 ( .A(n39849), .B(n39850), .Z(n39848) );
  AND U39702 ( .A(n39646), .B(n39649), .Z(n39754) );
  XOR U39703 ( .A(n39851), .B(n39805), .Z(n39649) );
  XNOR U39704 ( .A(p_input[1024]), .B(p_input[2048]), .Z(n39805) );
  XNOR U39705 ( .A(n39781), .B(n39780), .Z(n39851) );
  XNOR U39706 ( .A(n39852), .B(n39792), .Z(n39780) );
  XOR U39707 ( .A(n39766), .B(n39764), .Z(n39792) );
  XNOR U39708 ( .A(n39853), .B(n39771), .Z(n39764) );
  XOR U39709 ( .A(p_input[1048]), .B(p_input[2072]), .Z(n39771) );
  XOR U39710 ( .A(n39761), .B(n39770), .Z(n39853) );
  XOR U39711 ( .A(n39854), .B(n39767), .Z(n39770) );
  XOR U39712 ( .A(p_input[1046]), .B(p_input[2070]), .Z(n39767) );
  XOR U39713 ( .A(p_input[1047]), .B(n29410), .Z(n39854) );
  XOR U39714 ( .A(p_input[1042]), .B(p_input[2066]), .Z(n39761) );
  XNOR U39715 ( .A(n39776), .B(n39775), .Z(n39766) );
  XOR U39716 ( .A(n39855), .B(n39772), .Z(n39775) );
  XOR U39717 ( .A(p_input[1043]), .B(p_input[2067]), .Z(n39772) );
  XOR U39718 ( .A(p_input[1044]), .B(n29412), .Z(n39855) );
  XOR U39719 ( .A(p_input[1045]), .B(p_input[2069]), .Z(n39776) );
  XOR U39720 ( .A(n39791), .B(n39856), .Z(n39852) );
  IV U39721 ( .A(n39777), .Z(n39856) );
  XOR U39722 ( .A(p_input[1025]), .B(p_input[2049]), .Z(n39777) );
  XNOR U39723 ( .A(n39857), .B(n39799), .Z(n39791) );
  XNOR U39724 ( .A(n39787), .B(n39786), .Z(n39799) );
  XNOR U39725 ( .A(n39858), .B(n39783), .Z(n39786) );
  XNOR U39726 ( .A(p_input[1050]), .B(p_input[2074]), .Z(n39783) );
  XOR U39727 ( .A(p_input[1051]), .B(n29415), .Z(n39858) );
  XOR U39728 ( .A(p_input[1052]), .B(p_input[2076]), .Z(n39787) );
  XOR U39729 ( .A(n39797), .B(n39859), .Z(n39857) );
  IV U39730 ( .A(n39788), .Z(n39859) );
  XOR U39731 ( .A(p_input[1041]), .B(p_input[2065]), .Z(n39788) );
  XNOR U39732 ( .A(n39860), .B(n39804), .Z(n39797) );
  XNOR U39733 ( .A(p_input[1055]), .B(n29418), .Z(n39804) );
  XOR U39734 ( .A(n39794), .B(n39803), .Z(n39860) );
  XOR U39735 ( .A(n39861), .B(n39800), .Z(n39803) );
  XOR U39736 ( .A(p_input[1053]), .B(p_input[2077]), .Z(n39800) );
  XOR U39737 ( .A(p_input[1054]), .B(n29420), .Z(n39861) );
  XOR U39738 ( .A(p_input[1049]), .B(p_input[2073]), .Z(n39794) );
  XOR U39739 ( .A(n39816), .B(n39815), .Z(n39781) );
  XNOR U39740 ( .A(n39862), .B(n39823), .Z(n39815) );
  XNOR U39741 ( .A(n39811), .B(n39810), .Z(n39823) );
  XNOR U39742 ( .A(n39863), .B(n39807), .Z(n39810) );
  XNOR U39743 ( .A(p_input[1035]), .B(p_input[2059]), .Z(n39807) );
  XOR U39744 ( .A(p_input[1036]), .B(n28329), .Z(n39863) );
  XOR U39745 ( .A(p_input[1037]), .B(p_input[2061]), .Z(n39811) );
  XOR U39746 ( .A(n39821), .B(n39864), .Z(n39862) );
  IV U39747 ( .A(n39812), .Z(n39864) );
  XOR U39748 ( .A(p_input[1026]), .B(p_input[2050]), .Z(n39812) );
  XNOR U39749 ( .A(n39865), .B(n39828), .Z(n39821) );
  XNOR U39750 ( .A(p_input[1040]), .B(n28332), .Z(n39828) );
  XOR U39751 ( .A(n39818), .B(n39827), .Z(n39865) );
  XOR U39752 ( .A(n39866), .B(n39824), .Z(n39827) );
  XOR U39753 ( .A(p_input[1038]), .B(p_input[2062]), .Z(n39824) );
  XOR U39754 ( .A(p_input[1039]), .B(n28334), .Z(n39866) );
  XOR U39755 ( .A(p_input[1034]), .B(p_input[2058]), .Z(n39818) );
  XOR U39756 ( .A(n39835), .B(n39833), .Z(n39816) );
  XNOR U39757 ( .A(n39867), .B(n39840), .Z(n39833) );
  XOR U39758 ( .A(p_input[1033]), .B(p_input[2057]), .Z(n39840) );
  XOR U39759 ( .A(n39830), .B(n39839), .Z(n39867) );
  XOR U39760 ( .A(n39868), .B(n39836), .Z(n39839) );
  XOR U39761 ( .A(p_input[1031]), .B(p_input[2055]), .Z(n39836) );
  XOR U39762 ( .A(p_input[1032]), .B(n29427), .Z(n39868) );
  XOR U39763 ( .A(p_input[1027]), .B(p_input[2051]), .Z(n39830) );
  XNOR U39764 ( .A(n39845), .B(n39844), .Z(n39835) );
  XOR U39765 ( .A(n39869), .B(n39841), .Z(n39844) );
  XOR U39766 ( .A(p_input[1028]), .B(p_input[2052]), .Z(n39841) );
  XOR U39767 ( .A(p_input[1029]), .B(n29429), .Z(n39869) );
  XOR U39768 ( .A(p_input[1030]), .B(p_input[2054]), .Z(n39845) );
  XNOR U39769 ( .A(n39870), .B(n39871), .Z(n39646) );
  AND U39770 ( .A(n743), .B(n39872), .Z(n39871) );
  XNOR U39771 ( .A(n39873), .B(n39874), .Z(n743) );
  AND U39772 ( .A(n39875), .B(n39876), .Z(n39874) );
  XOR U39773 ( .A(n39660), .B(n39873), .Z(n39876) );
  XNOR U39774 ( .A(n39877), .B(n39873), .Z(n39875) );
  XOR U39775 ( .A(n39878), .B(n39879), .Z(n39873) );
  AND U39776 ( .A(n39880), .B(n39881), .Z(n39879) );
  XOR U39777 ( .A(n39675), .B(n39878), .Z(n39881) );
  XOR U39778 ( .A(n39878), .B(n39676), .Z(n39880) );
  XOR U39779 ( .A(n39882), .B(n39883), .Z(n39878) );
  AND U39780 ( .A(n39884), .B(n39885), .Z(n39883) );
  XOR U39781 ( .A(n39703), .B(n39882), .Z(n39885) );
  XOR U39782 ( .A(n39882), .B(n39704), .Z(n39884) );
  XOR U39783 ( .A(n39886), .B(n39887), .Z(n39882) );
  AND U39784 ( .A(n39888), .B(n39889), .Z(n39887) );
  XOR U39785 ( .A(n39752), .B(n39886), .Z(n39889) );
  XOR U39786 ( .A(n39886), .B(n39753), .Z(n39888) );
  XOR U39787 ( .A(n39890), .B(n39891), .Z(n39886) );
  AND U39788 ( .A(n39892), .B(n39893), .Z(n39891) );
  XOR U39789 ( .A(n39890), .B(n39849), .Z(n39893) );
  XNOR U39790 ( .A(n39894), .B(n39895), .Z(n39596) );
  AND U39791 ( .A(n747), .B(n39896), .Z(n39895) );
  XNOR U39792 ( .A(n39897), .B(n39898), .Z(n747) );
  AND U39793 ( .A(n39899), .B(n39900), .Z(n39898) );
  XOR U39794 ( .A(n39897), .B(n39606), .Z(n39900) );
  XNOR U39795 ( .A(n39897), .B(n39556), .Z(n39899) );
  XOR U39796 ( .A(n39901), .B(n39902), .Z(n39897) );
  AND U39797 ( .A(n39903), .B(n39904), .Z(n39902) );
  XNOR U39798 ( .A(n39616), .B(n39901), .Z(n39904) );
  XOR U39799 ( .A(n39901), .B(n39566), .Z(n39903) );
  XOR U39800 ( .A(n39905), .B(n39906), .Z(n39901) );
  AND U39801 ( .A(n39907), .B(n39908), .Z(n39906) );
  XNOR U39802 ( .A(n39626), .B(n39905), .Z(n39908) );
  XOR U39803 ( .A(n39905), .B(n39575), .Z(n39907) );
  XOR U39804 ( .A(n39909), .B(n39910), .Z(n39905) );
  AND U39805 ( .A(n39911), .B(n39912), .Z(n39910) );
  XOR U39806 ( .A(n39909), .B(n39583), .Z(n39911) );
  XOR U39807 ( .A(n39913), .B(n39914), .Z(n39547) );
  AND U39808 ( .A(n751), .B(n39896), .Z(n39914) );
  XNOR U39809 ( .A(n39894), .B(n39913), .Z(n39896) );
  XNOR U39810 ( .A(n39915), .B(n39916), .Z(n751) );
  AND U39811 ( .A(n39917), .B(n39918), .Z(n39916) );
  XNOR U39812 ( .A(n39919), .B(n39915), .Z(n39918) );
  IV U39813 ( .A(n39606), .Z(n39919) );
  XOR U39814 ( .A(n39877), .B(n39920), .Z(n39606) );
  AND U39815 ( .A(n754), .B(n39921), .Z(n39920) );
  XOR U39816 ( .A(n39659), .B(n39656), .Z(n39921) );
  IV U39817 ( .A(n39877), .Z(n39659) );
  XNOR U39818 ( .A(n39556), .B(n39915), .Z(n39917) );
  XOR U39819 ( .A(n39922), .B(n39923), .Z(n39556) );
  AND U39820 ( .A(n770), .B(n39924), .Z(n39923) );
  XOR U39821 ( .A(n39925), .B(n39926), .Z(n39915) );
  AND U39822 ( .A(n39927), .B(n39928), .Z(n39926) );
  XNOR U39823 ( .A(n39925), .B(n39616), .Z(n39928) );
  XOR U39824 ( .A(n39676), .B(n39929), .Z(n39616) );
  AND U39825 ( .A(n754), .B(n39930), .Z(n39929) );
  XOR U39826 ( .A(n39672), .B(n39676), .Z(n39930) );
  XNOR U39827 ( .A(n39931), .B(n39925), .Z(n39927) );
  IV U39828 ( .A(n39566), .Z(n39931) );
  XOR U39829 ( .A(n39932), .B(n39933), .Z(n39566) );
  AND U39830 ( .A(n770), .B(n39934), .Z(n39933) );
  XOR U39831 ( .A(n39935), .B(n39936), .Z(n39925) );
  AND U39832 ( .A(n39937), .B(n39938), .Z(n39936) );
  XNOR U39833 ( .A(n39935), .B(n39626), .Z(n39938) );
  XOR U39834 ( .A(n39704), .B(n39939), .Z(n39626) );
  AND U39835 ( .A(n754), .B(n39940), .Z(n39939) );
  XOR U39836 ( .A(n39700), .B(n39704), .Z(n39940) );
  XOR U39837 ( .A(n39575), .B(n39935), .Z(n39937) );
  XOR U39838 ( .A(n39941), .B(n39942), .Z(n39575) );
  AND U39839 ( .A(n770), .B(n39943), .Z(n39942) );
  XOR U39840 ( .A(n39909), .B(n39944), .Z(n39935) );
  AND U39841 ( .A(n39945), .B(n39912), .Z(n39944) );
  XNOR U39842 ( .A(n39636), .B(n39909), .Z(n39912) );
  XOR U39843 ( .A(n39753), .B(n39946), .Z(n39636) );
  AND U39844 ( .A(n754), .B(n39947), .Z(n39946) );
  XOR U39845 ( .A(n39749), .B(n39753), .Z(n39947) );
  XNOR U39846 ( .A(n39948), .B(n39909), .Z(n39945) );
  IV U39847 ( .A(n39583), .Z(n39948) );
  XOR U39848 ( .A(n39949), .B(n39950), .Z(n39583) );
  AND U39849 ( .A(n770), .B(n39951), .Z(n39950) );
  XOR U39850 ( .A(n39952), .B(n39953), .Z(n39909) );
  AND U39851 ( .A(n39954), .B(n39955), .Z(n39953) );
  XNOR U39852 ( .A(n39952), .B(n39644), .Z(n39955) );
  XOR U39853 ( .A(n39850), .B(n39956), .Z(n39644) );
  AND U39854 ( .A(n754), .B(n39957), .Z(n39956) );
  XOR U39855 ( .A(n39846), .B(n39850), .Z(n39957) );
  XNOR U39856 ( .A(n39958), .B(n39952), .Z(n39954) );
  IV U39857 ( .A(n39593), .Z(n39958) );
  XOR U39858 ( .A(n39959), .B(n39960), .Z(n39593) );
  AND U39859 ( .A(n770), .B(n39961), .Z(n39960) );
  AND U39860 ( .A(n39913), .B(n39894), .Z(n39952) );
  XNOR U39861 ( .A(n39962), .B(n39963), .Z(n39894) );
  AND U39862 ( .A(n754), .B(n39872), .Z(n39963) );
  XNOR U39863 ( .A(n39870), .B(n39962), .Z(n39872) );
  XNOR U39864 ( .A(n39964), .B(n39965), .Z(n754) );
  AND U39865 ( .A(n39966), .B(n39967), .Z(n39965) );
  XNOR U39866 ( .A(n39964), .B(n39656), .Z(n39967) );
  IV U39867 ( .A(n39660), .Z(n39656) );
  XOR U39868 ( .A(n39968), .B(n39969), .Z(n39660) );
  AND U39869 ( .A(n758), .B(n39970), .Z(n39969) );
  XOR U39870 ( .A(n39971), .B(n39968), .Z(n39970) );
  XNOR U39871 ( .A(n39964), .B(n39877), .Z(n39966) );
  XOR U39872 ( .A(n39972), .B(n39973), .Z(n39877) );
  AND U39873 ( .A(n766), .B(n39924), .Z(n39973) );
  XOR U39874 ( .A(n39922), .B(n39972), .Z(n39924) );
  XOR U39875 ( .A(n39974), .B(n39975), .Z(n39964) );
  AND U39876 ( .A(n39976), .B(n39977), .Z(n39975) );
  XNOR U39877 ( .A(n39974), .B(n39672), .Z(n39977) );
  IV U39878 ( .A(n39675), .Z(n39672) );
  XOR U39879 ( .A(n39978), .B(n39979), .Z(n39675) );
  AND U39880 ( .A(n758), .B(n39980), .Z(n39979) );
  XOR U39881 ( .A(n39981), .B(n39978), .Z(n39980) );
  XOR U39882 ( .A(n39676), .B(n39974), .Z(n39976) );
  XOR U39883 ( .A(n39982), .B(n39983), .Z(n39676) );
  AND U39884 ( .A(n766), .B(n39934), .Z(n39983) );
  XOR U39885 ( .A(n39982), .B(n39932), .Z(n39934) );
  XOR U39886 ( .A(n39984), .B(n39985), .Z(n39974) );
  AND U39887 ( .A(n39986), .B(n39987), .Z(n39985) );
  XNOR U39888 ( .A(n39984), .B(n39700), .Z(n39987) );
  IV U39889 ( .A(n39703), .Z(n39700) );
  XOR U39890 ( .A(n39988), .B(n39989), .Z(n39703) );
  AND U39891 ( .A(n758), .B(n39990), .Z(n39989) );
  XNOR U39892 ( .A(n39991), .B(n39988), .Z(n39990) );
  XOR U39893 ( .A(n39704), .B(n39984), .Z(n39986) );
  XOR U39894 ( .A(n39992), .B(n39993), .Z(n39704) );
  AND U39895 ( .A(n766), .B(n39943), .Z(n39993) );
  XOR U39896 ( .A(n39992), .B(n39941), .Z(n39943) );
  XOR U39897 ( .A(n39994), .B(n39995), .Z(n39984) );
  AND U39898 ( .A(n39996), .B(n39997), .Z(n39995) );
  XNOR U39899 ( .A(n39994), .B(n39749), .Z(n39997) );
  IV U39900 ( .A(n39752), .Z(n39749) );
  XOR U39901 ( .A(n39998), .B(n39999), .Z(n39752) );
  AND U39902 ( .A(n758), .B(n40000), .Z(n39999) );
  XOR U39903 ( .A(n40001), .B(n39998), .Z(n40000) );
  XOR U39904 ( .A(n39753), .B(n39994), .Z(n39996) );
  XOR U39905 ( .A(n40002), .B(n40003), .Z(n39753) );
  AND U39906 ( .A(n766), .B(n39951), .Z(n40003) );
  XOR U39907 ( .A(n40002), .B(n39949), .Z(n39951) );
  XOR U39908 ( .A(n39890), .B(n40004), .Z(n39994) );
  AND U39909 ( .A(n39892), .B(n40005), .Z(n40004) );
  XNOR U39910 ( .A(n39890), .B(n39846), .Z(n40005) );
  IV U39911 ( .A(n39849), .Z(n39846) );
  XOR U39912 ( .A(n40006), .B(n40007), .Z(n39849) );
  AND U39913 ( .A(n758), .B(n40008), .Z(n40007) );
  XNOR U39914 ( .A(n40009), .B(n40006), .Z(n40008) );
  XOR U39915 ( .A(n39850), .B(n39890), .Z(n39892) );
  XOR U39916 ( .A(n40010), .B(n40011), .Z(n39850) );
  AND U39917 ( .A(n766), .B(n39961), .Z(n40011) );
  XOR U39918 ( .A(n40010), .B(n39959), .Z(n39961) );
  AND U39919 ( .A(n39962), .B(n39870), .Z(n39890) );
  XNOR U39920 ( .A(n40012), .B(n40013), .Z(n39870) );
  AND U39921 ( .A(n758), .B(n40014), .Z(n40013) );
  XNOR U39922 ( .A(n40015), .B(n40012), .Z(n40014) );
  XNOR U39923 ( .A(n40016), .B(n40017), .Z(n758) );
  AND U39924 ( .A(n40018), .B(n40019), .Z(n40017) );
  XOR U39925 ( .A(n39971), .B(n40016), .Z(n40019) );
  AND U39926 ( .A(n40020), .B(n40021), .Z(n39971) );
  XNOR U39927 ( .A(n39968), .B(n40016), .Z(n40018) );
  XNOR U39928 ( .A(n40022), .B(n40023), .Z(n39968) );
  AND U39929 ( .A(n762), .B(n40024), .Z(n40023) );
  XNOR U39930 ( .A(n40025), .B(n40026), .Z(n40024) );
  XOR U39931 ( .A(n40027), .B(n40028), .Z(n40016) );
  AND U39932 ( .A(n40029), .B(n40030), .Z(n40028) );
  XNOR U39933 ( .A(n40027), .B(n40020), .Z(n40030) );
  IV U39934 ( .A(n39981), .Z(n40020) );
  XOR U39935 ( .A(n40031), .B(n40032), .Z(n39981) );
  XOR U39936 ( .A(n40033), .B(n40021), .Z(n40032) );
  AND U39937 ( .A(n39991), .B(n40034), .Z(n40021) );
  AND U39938 ( .A(n40035), .B(n40036), .Z(n40033) );
  XOR U39939 ( .A(n40037), .B(n40031), .Z(n40035) );
  XNOR U39940 ( .A(n39978), .B(n40027), .Z(n40029) );
  XNOR U39941 ( .A(n40038), .B(n40039), .Z(n39978) );
  AND U39942 ( .A(n762), .B(n40040), .Z(n40039) );
  XNOR U39943 ( .A(n40041), .B(n40042), .Z(n40040) );
  XOR U39944 ( .A(n40043), .B(n40044), .Z(n40027) );
  AND U39945 ( .A(n40045), .B(n40046), .Z(n40044) );
  XNOR U39946 ( .A(n40043), .B(n39991), .Z(n40046) );
  XOR U39947 ( .A(n40047), .B(n40036), .Z(n39991) );
  XNOR U39948 ( .A(n40048), .B(n40031), .Z(n40036) );
  XOR U39949 ( .A(n40049), .B(n40050), .Z(n40031) );
  AND U39950 ( .A(n40051), .B(n40052), .Z(n40050) );
  XOR U39951 ( .A(n40053), .B(n40049), .Z(n40051) );
  XNOR U39952 ( .A(n40054), .B(n40055), .Z(n40048) );
  AND U39953 ( .A(n40056), .B(n40057), .Z(n40055) );
  XOR U39954 ( .A(n40054), .B(n40058), .Z(n40056) );
  XNOR U39955 ( .A(n40037), .B(n40034), .Z(n40047) );
  AND U39956 ( .A(n40059), .B(n40060), .Z(n40034) );
  XOR U39957 ( .A(n40061), .B(n40062), .Z(n40037) );
  AND U39958 ( .A(n40063), .B(n40064), .Z(n40062) );
  XOR U39959 ( .A(n40061), .B(n40065), .Z(n40063) );
  XNOR U39960 ( .A(n39988), .B(n40043), .Z(n40045) );
  XNOR U39961 ( .A(n40066), .B(n40067), .Z(n39988) );
  AND U39962 ( .A(n762), .B(n40068), .Z(n40067) );
  XNOR U39963 ( .A(n40069), .B(n40070), .Z(n40068) );
  XOR U39964 ( .A(n40071), .B(n40072), .Z(n40043) );
  AND U39965 ( .A(n40073), .B(n40074), .Z(n40072) );
  XNOR U39966 ( .A(n40071), .B(n40059), .Z(n40074) );
  IV U39967 ( .A(n40001), .Z(n40059) );
  XNOR U39968 ( .A(n40075), .B(n40052), .Z(n40001) );
  XNOR U39969 ( .A(n40076), .B(n40058), .Z(n40052) );
  XOR U39970 ( .A(n40077), .B(n40078), .Z(n40058) );
  AND U39971 ( .A(n40079), .B(n40080), .Z(n40078) );
  XOR U39972 ( .A(n40077), .B(n40081), .Z(n40079) );
  XNOR U39973 ( .A(n40057), .B(n40049), .Z(n40076) );
  XOR U39974 ( .A(n40082), .B(n40083), .Z(n40049) );
  AND U39975 ( .A(n40084), .B(n40085), .Z(n40083) );
  XNOR U39976 ( .A(n40086), .B(n40082), .Z(n40084) );
  XNOR U39977 ( .A(n40087), .B(n40054), .Z(n40057) );
  XOR U39978 ( .A(n40088), .B(n40089), .Z(n40054) );
  AND U39979 ( .A(n40090), .B(n40091), .Z(n40089) );
  XOR U39980 ( .A(n40088), .B(n40092), .Z(n40090) );
  XNOR U39981 ( .A(n40093), .B(n40094), .Z(n40087) );
  AND U39982 ( .A(n40095), .B(n40096), .Z(n40094) );
  XNOR U39983 ( .A(n40093), .B(n40097), .Z(n40095) );
  XNOR U39984 ( .A(n40053), .B(n40060), .Z(n40075) );
  AND U39985 ( .A(n40009), .B(n40098), .Z(n40060) );
  XOR U39986 ( .A(n40065), .B(n40064), .Z(n40053) );
  XNOR U39987 ( .A(n40099), .B(n40061), .Z(n40064) );
  XOR U39988 ( .A(n40100), .B(n40101), .Z(n40061) );
  AND U39989 ( .A(n40102), .B(n40103), .Z(n40101) );
  XOR U39990 ( .A(n40100), .B(n40104), .Z(n40102) );
  XNOR U39991 ( .A(n40105), .B(n40106), .Z(n40099) );
  AND U39992 ( .A(n40107), .B(n40108), .Z(n40106) );
  XOR U39993 ( .A(n40105), .B(n40109), .Z(n40107) );
  XOR U39994 ( .A(n40110), .B(n40111), .Z(n40065) );
  AND U39995 ( .A(n40112), .B(n40113), .Z(n40111) );
  XOR U39996 ( .A(n40110), .B(n40114), .Z(n40112) );
  XNOR U39997 ( .A(n39998), .B(n40071), .Z(n40073) );
  XNOR U39998 ( .A(n40115), .B(n40116), .Z(n39998) );
  AND U39999 ( .A(n762), .B(n40117), .Z(n40116) );
  XNOR U40000 ( .A(n40118), .B(n40119), .Z(n40117) );
  XOR U40001 ( .A(n40120), .B(n40121), .Z(n40071) );
  AND U40002 ( .A(n40122), .B(n40123), .Z(n40121) );
  XNOR U40003 ( .A(n40120), .B(n40009), .Z(n40123) );
  XOR U40004 ( .A(n40124), .B(n40085), .Z(n40009) );
  XNOR U40005 ( .A(n40125), .B(n40092), .Z(n40085) );
  XOR U40006 ( .A(n40081), .B(n40080), .Z(n40092) );
  XNOR U40007 ( .A(n40126), .B(n40077), .Z(n40080) );
  XOR U40008 ( .A(n40127), .B(n40128), .Z(n40077) );
  AND U40009 ( .A(n40129), .B(n40130), .Z(n40128) );
  XNOR U40010 ( .A(n40131), .B(n40132), .Z(n40129) );
  IV U40011 ( .A(n40127), .Z(n40131) );
  XNOR U40012 ( .A(n40133), .B(n40134), .Z(n40126) );
  NOR U40013 ( .A(n40135), .B(n40136), .Z(n40134) );
  XNOR U40014 ( .A(n40133), .B(n40137), .Z(n40135) );
  XOR U40015 ( .A(n40138), .B(n40139), .Z(n40081) );
  NOR U40016 ( .A(n40140), .B(n40141), .Z(n40139) );
  XNOR U40017 ( .A(n40138), .B(n40142), .Z(n40140) );
  XNOR U40018 ( .A(n40091), .B(n40082), .Z(n40125) );
  XOR U40019 ( .A(n40143), .B(n40144), .Z(n40082) );
  AND U40020 ( .A(n40145), .B(n40146), .Z(n40144) );
  XOR U40021 ( .A(n40143), .B(n40147), .Z(n40145) );
  XOR U40022 ( .A(n40148), .B(n40097), .Z(n40091) );
  XOR U40023 ( .A(n40149), .B(n40150), .Z(n40097) );
  NOR U40024 ( .A(n40151), .B(n40152), .Z(n40150) );
  XOR U40025 ( .A(n40149), .B(n40153), .Z(n40151) );
  XNOR U40026 ( .A(n40096), .B(n40088), .Z(n40148) );
  XOR U40027 ( .A(n40154), .B(n40155), .Z(n40088) );
  AND U40028 ( .A(n40156), .B(n40157), .Z(n40155) );
  XOR U40029 ( .A(n40154), .B(n40158), .Z(n40156) );
  XNOR U40030 ( .A(n40159), .B(n40093), .Z(n40096) );
  XOR U40031 ( .A(n40160), .B(n40161), .Z(n40093) );
  AND U40032 ( .A(n40162), .B(n40163), .Z(n40161) );
  XNOR U40033 ( .A(n40164), .B(n40165), .Z(n40162) );
  IV U40034 ( .A(n40160), .Z(n40164) );
  XNOR U40035 ( .A(n40166), .B(n40167), .Z(n40159) );
  NOR U40036 ( .A(n40168), .B(n40169), .Z(n40167) );
  XNOR U40037 ( .A(n40166), .B(n40170), .Z(n40168) );
  XOR U40038 ( .A(n40086), .B(n40098), .Z(n40124) );
  NOR U40039 ( .A(n40015), .B(n40171), .Z(n40098) );
  XNOR U40040 ( .A(n40104), .B(n40103), .Z(n40086) );
  XNOR U40041 ( .A(n40172), .B(n40109), .Z(n40103) );
  XNOR U40042 ( .A(n40173), .B(n40174), .Z(n40109) );
  NOR U40043 ( .A(n40175), .B(n40176), .Z(n40174) );
  XOR U40044 ( .A(n40173), .B(n40177), .Z(n40175) );
  XNOR U40045 ( .A(n40108), .B(n40100), .Z(n40172) );
  XOR U40046 ( .A(n40178), .B(n40179), .Z(n40100) );
  AND U40047 ( .A(n40180), .B(n40181), .Z(n40179) );
  XOR U40048 ( .A(n40178), .B(n40182), .Z(n40180) );
  XNOR U40049 ( .A(n40183), .B(n40105), .Z(n40108) );
  XOR U40050 ( .A(n40184), .B(n40185), .Z(n40105) );
  AND U40051 ( .A(n40186), .B(n40187), .Z(n40185) );
  XNOR U40052 ( .A(n40188), .B(n40189), .Z(n40186) );
  IV U40053 ( .A(n40184), .Z(n40188) );
  XNOR U40054 ( .A(n40190), .B(n40191), .Z(n40183) );
  NOR U40055 ( .A(n40192), .B(n40193), .Z(n40191) );
  XNOR U40056 ( .A(n40190), .B(n40194), .Z(n40192) );
  XOR U40057 ( .A(n40114), .B(n40113), .Z(n40104) );
  XNOR U40058 ( .A(n40195), .B(n40110), .Z(n40113) );
  XOR U40059 ( .A(n40196), .B(n40197), .Z(n40110) );
  AND U40060 ( .A(n40198), .B(n40199), .Z(n40197) );
  XNOR U40061 ( .A(n40200), .B(n40201), .Z(n40198) );
  IV U40062 ( .A(n40196), .Z(n40200) );
  XNOR U40063 ( .A(n40202), .B(n40203), .Z(n40195) );
  NOR U40064 ( .A(n40204), .B(n40205), .Z(n40203) );
  XNOR U40065 ( .A(n40202), .B(n40206), .Z(n40204) );
  XOR U40066 ( .A(n40207), .B(n40208), .Z(n40114) );
  NOR U40067 ( .A(n40209), .B(n40210), .Z(n40208) );
  XNOR U40068 ( .A(n40207), .B(n40211), .Z(n40209) );
  XNOR U40069 ( .A(n40006), .B(n40120), .Z(n40122) );
  XNOR U40070 ( .A(n40212), .B(n40213), .Z(n40006) );
  AND U40071 ( .A(n762), .B(n40214), .Z(n40213) );
  XNOR U40072 ( .A(n40215), .B(n40216), .Z(n40214) );
  AND U40073 ( .A(n40012), .B(n40015), .Z(n40120) );
  XOR U40074 ( .A(n40217), .B(n40171), .Z(n40015) );
  XNOR U40075 ( .A(p_input[1056]), .B(p_input[2048]), .Z(n40171) );
  XNOR U40076 ( .A(n40147), .B(n40146), .Z(n40217) );
  XNOR U40077 ( .A(n40218), .B(n40158), .Z(n40146) );
  XOR U40078 ( .A(n40132), .B(n40130), .Z(n40158) );
  XNOR U40079 ( .A(n40219), .B(n40137), .Z(n40130) );
  XOR U40080 ( .A(p_input[1080]), .B(p_input[2072]), .Z(n40137) );
  XOR U40081 ( .A(n40127), .B(n40136), .Z(n40219) );
  XOR U40082 ( .A(n40220), .B(n40133), .Z(n40136) );
  XOR U40083 ( .A(p_input[1078]), .B(p_input[2070]), .Z(n40133) );
  XOR U40084 ( .A(p_input[1079]), .B(n29410), .Z(n40220) );
  XOR U40085 ( .A(p_input[1074]), .B(p_input[2066]), .Z(n40127) );
  XNOR U40086 ( .A(n40142), .B(n40141), .Z(n40132) );
  XOR U40087 ( .A(n40221), .B(n40138), .Z(n40141) );
  XOR U40088 ( .A(p_input[1075]), .B(p_input[2067]), .Z(n40138) );
  XOR U40089 ( .A(p_input[1076]), .B(n29412), .Z(n40221) );
  XOR U40090 ( .A(p_input[1077]), .B(p_input[2069]), .Z(n40142) );
  XOR U40091 ( .A(n40157), .B(n40222), .Z(n40218) );
  IV U40092 ( .A(n40143), .Z(n40222) );
  XOR U40093 ( .A(p_input[1057]), .B(p_input[2049]), .Z(n40143) );
  XNOR U40094 ( .A(n40223), .B(n40165), .Z(n40157) );
  XNOR U40095 ( .A(n40153), .B(n40152), .Z(n40165) );
  XNOR U40096 ( .A(n40224), .B(n40149), .Z(n40152) );
  XNOR U40097 ( .A(p_input[1082]), .B(p_input[2074]), .Z(n40149) );
  XOR U40098 ( .A(p_input[1083]), .B(n29415), .Z(n40224) );
  XOR U40099 ( .A(p_input[1084]), .B(p_input[2076]), .Z(n40153) );
  XOR U40100 ( .A(n40163), .B(n40225), .Z(n40223) );
  IV U40101 ( .A(n40154), .Z(n40225) );
  XOR U40102 ( .A(p_input[1073]), .B(p_input[2065]), .Z(n40154) );
  XNOR U40103 ( .A(n40226), .B(n40170), .Z(n40163) );
  XNOR U40104 ( .A(p_input[1087]), .B(n29418), .Z(n40170) );
  XOR U40105 ( .A(n40160), .B(n40169), .Z(n40226) );
  XOR U40106 ( .A(n40227), .B(n40166), .Z(n40169) );
  XOR U40107 ( .A(p_input[1085]), .B(p_input[2077]), .Z(n40166) );
  XOR U40108 ( .A(p_input[1086]), .B(n29420), .Z(n40227) );
  XOR U40109 ( .A(p_input[1081]), .B(p_input[2073]), .Z(n40160) );
  XOR U40110 ( .A(n40182), .B(n40181), .Z(n40147) );
  XNOR U40111 ( .A(n40228), .B(n40189), .Z(n40181) );
  XNOR U40112 ( .A(n40177), .B(n40176), .Z(n40189) );
  XNOR U40113 ( .A(n40229), .B(n40173), .Z(n40176) );
  XNOR U40114 ( .A(p_input[1067]), .B(p_input[2059]), .Z(n40173) );
  XOR U40115 ( .A(p_input[1068]), .B(n28329), .Z(n40229) );
  XOR U40116 ( .A(p_input[1069]), .B(p_input[2061]), .Z(n40177) );
  XOR U40117 ( .A(n40187), .B(n40230), .Z(n40228) );
  IV U40118 ( .A(n40178), .Z(n40230) );
  XOR U40119 ( .A(p_input[1058]), .B(p_input[2050]), .Z(n40178) );
  XNOR U40120 ( .A(n40231), .B(n40194), .Z(n40187) );
  XNOR U40121 ( .A(p_input[1072]), .B(n28332), .Z(n40194) );
  XOR U40122 ( .A(n40184), .B(n40193), .Z(n40231) );
  XOR U40123 ( .A(n40232), .B(n40190), .Z(n40193) );
  XOR U40124 ( .A(p_input[1070]), .B(p_input[2062]), .Z(n40190) );
  XOR U40125 ( .A(p_input[1071]), .B(n28334), .Z(n40232) );
  XOR U40126 ( .A(p_input[1066]), .B(p_input[2058]), .Z(n40184) );
  XOR U40127 ( .A(n40201), .B(n40199), .Z(n40182) );
  XNOR U40128 ( .A(n40233), .B(n40206), .Z(n40199) );
  XOR U40129 ( .A(p_input[1065]), .B(p_input[2057]), .Z(n40206) );
  XOR U40130 ( .A(n40196), .B(n40205), .Z(n40233) );
  XOR U40131 ( .A(n40234), .B(n40202), .Z(n40205) );
  XOR U40132 ( .A(p_input[1063]), .B(p_input[2055]), .Z(n40202) );
  XOR U40133 ( .A(p_input[1064]), .B(n29427), .Z(n40234) );
  XOR U40134 ( .A(p_input[1059]), .B(p_input[2051]), .Z(n40196) );
  XNOR U40135 ( .A(n40211), .B(n40210), .Z(n40201) );
  XOR U40136 ( .A(n40235), .B(n40207), .Z(n40210) );
  XOR U40137 ( .A(p_input[1060]), .B(p_input[2052]), .Z(n40207) );
  XOR U40138 ( .A(p_input[1061]), .B(n29429), .Z(n40235) );
  XOR U40139 ( .A(p_input[1062]), .B(p_input[2054]), .Z(n40211) );
  XNOR U40140 ( .A(n40236), .B(n40237), .Z(n40012) );
  AND U40141 ( .A(n762), .B(n40238), .Z(n40237) );
  XNOR U40142 ( .A(n40239), .B(n40240), .Z(n762) );
  AND U40143 ( .A(n40241), .B(n40242), .Z(n40240) );
  XOR U40144 ( .A(n40026), .B(n40239), .Z(n40242) );
  XNOR U40145 ( .A(n40243), .B(n40239), .Z(n40241) );
  XOR U40146 ( .A(n40244), .B(n40245), .Z(n40239) );
  AND U40147 ( .A(n40246), .B(n40247), .Z(n40245) );
  XOR U40148 ( .A(n40041), .B(n40244), .Z(n40247) );
  XOR U40149 ( .A(n40244), .B(n40042), .Z(n40246) );
  XOR U40150 ( .A(n40248), .B(n40249), .Z(n40244) );
  AND U40151 ( .A(n40250), .B(n40251), .Z(n40249) );
  XOR U40152 ( .A(n40069), .B(n40248), .Z(n40251) );
  XOR U40153 ( .A(n40248), .B(n40070), .Z(n40250) );
  XOR U40154 ( .A(n40252), .B(n40253), .Z(n40248) );
  AND U40155 ( .A(n40254), .B(n40255), .Z(n40253) );
  XOR U40156 ( .A(n40118), .B(n40252), .Z(n40255) );
  XOR U40157 ( .A(n40252), .B(n40119), .Z(n40254) );
  XOR U40158 ( .A(n40256), .B(n40257), .Z(n40252) );
  AND U40159 ( .A(n40258), .B(n40259), .Z(n40257) );
  XOR U40160 ( .A(n40256), .B(n40215), .Z(n40259) );
  XNOR U40161 ( .A(n40260), .B(n40261), .Z(n39962) );
  AND U40162 ( .A(n766), .B(n40262), .Z(n40261) );
  XNOR U40163 ( .A(n40263), .B(n40264), .Z(n766) );
  AND U40164 ( .A(n40265), .B(n40266), .Z(n40264) );
  XOR U40165 ( .A(n40263), .B(n39972), .Z(n40266) );
  XNOR U40166 ( .A(n40263), .B(n39922), .Z(n40265) );
  XOR U40167 ( .A(n40267), .B(n40268), .Z(n40263) );
  AND U40168 ( .A(n40269), .B(n40270), .Z(n40268) );
  XNOR U40169 ( .A(n39982), .B(n40267), .Z(n40270) );
  XOR U40170 ( .A(n40267), .B(n39932), .Z(n40269) );
  XOR U40171 ( .A(n40271), .B(n40272), .Z(n40267) );
  AND U40172 ( .A(n40273), .B(n40274), .Z(n40272) );
  XNOR U40173 ( .A(n39992), .B(n40271), .Z(n40274) );
  XOR U40174 ( .A(n40271), .B(n39941), .Z(n40273) );
  XOR U40175 ( .A(n40275), .B(n40276), .Z(n40271) );
  AND U40176 ( .A(n40277), .B(n40278), .Z(n40276) );
  XOR U40177 ( .A(n40275), .B(n39949), .Z(n40277) );
  XOR U40178 ( .A(n40279), .B(n40280), .Z(n39913) );
  AND U40179 ( .A(n770), .B(n40262), .Z(n40280) );
  XNOR U40180 ( .A(n40260), .B(n40279), .Z(n40262) );
  XNOR U40181 ( .A(n40281), .B(n40282), .Z(n770) );
  AND U40182 ( .A(n40283), .B(n40284), .Z(n40282) );
  XNOR U40183 ( .A(n40285), .B(n40281), .Z(n40284) );
  IV U40184 ( .A(n39972), .Z(n40285) );
  XOR U40185 ( .A(n40243), .B(n40286), .Z(n39972) );
  AND U40186 ( .A(n773), .B(n40287), .Z(n40286) );
  XOR U40187 ( .A(n40025), .B(n40022), .Z(n40287) );
  IV U40188 ( .A(n40243), .Z(n40025) );
  XNOR U40189 ( .A(n39922), .B(n40281), .Z(n40283) );
  XOR U40190 ( .A(n40288), .B(n40289), .Z(n39922) );
  AND U40191 ( .A(n789), .B(n40290), .Z(n40289) );
  XOR U40192 ( .A(n40291), .B(n40292), .Z(n40281) );
  AND U40193 ( .A(n40293), .B(n40294), .Z(n40292) );
  XNOR U40194 ( .A(n40291), .B(n39982), .Z(n40294) );
  XOR U40195 ( .A(n40042), .B(n40295), .Z(n39982) );
  AND U40196 ( .A(n773), .B(n40296), .Z(n40295) );
  XOR U40197 ( .A(n40038), .B(n40042), .Z(n40296) );
  XNOR U40198 ( .A(n40297), .B(n40291), .Z(n40293) );
  IV U40199 ( .A(n39932), .Z(n40297) );
  XOR U40200 ( .A(n40298), .B(n40299), .Z(n39932) );
  AND U40201 ( .A(n789), .B(n40300), .Z(n40299) );
  XOR U40202 ( .A(n40301), .B(n40302), .Z(n40291) );
  AND U40203 ( .A(n40303), .B(n40304), .Z(n40302) );
  XNOR U40204 ( .A(n40301), .B(n39992), .Z(n40304) );
  XOR U40205 ( .A(n40070), .B(n40305), .Z(n39992) );
  AND U40206 ( .A(n773), .B(n40306), .Z(n40305) );
  XOR U40207 ( .A(n40066), .B(n40070), .Z(n40306) );
  XOR U40208 ( .A(n39941), .B(n40301), .Z(n40303) );
  XOR U40209 ( .A(n40307), .B(n40308), .Z(n39941) );
  AND U40210 ( .A(n789), .B(n40309), .Z(n40308) );
  XOR U40211 ( .A(n40275), .B(n40310), .Z(n40301) );
  AND U40212 ( .A(n40311), .B(n40278), .Z(n40310) );
  XNOR U40213 ( .A(n40002), .B(n40275), .Z(n40278) );
  XOR U40214 ( .A(n40119), .B(n40312), .Z(n40002) );
  AND U40215 ( .A(n773), .B(n40313), .Z(n40312) );
  XOR U40216 ( .A(n40115), .B(n40119), .Z(n40313) );
  XNOR U40217 ( .A(n40314), .B(n40275), .Z(n40311) );
  IV U40218 ( .A(n39949), .Z(n40314) );
  XOR U40219 ( .A(n40315), .B(n40316), .Z(n39949) );
  AND U40220 ( .A(n789), .B(n40317), .Z(n40316) );
  XOR U40221 ( .A(n40318), .B(n40319), .Z(n40275) );
  AND U40222 ( .A(n40320), .B(n40321), .Z(n40319) );
  XNOR U40223 ( .A(n40318), .B(n40010), .Z(n40321) );
  XOR U40224 ( .A(n40216), .B(n40322), .Z(n40010) );
  AND U40225 ( .A(n773), .B(n40323), .Z(n40322) );
  XOR U40226 ( .A(n40212), .B(n40216), .Z(n40323) );
  XNOR U40227 ( .A(n40324), .B(n40318), .Z(n40320) );
  IV U40228 ( .A(n39959), .Z(n40324) );
  XOR U40229 ( .A(n40325), .B(n40326), .Z(n39959) );
  AND U40230 ( .A(n789), .B(n40327), .Z(n40326) );
  AND U40231 ( .A(n40279), .B(n40260), .Z(n40318) );
  XNOR U40232 ( .A(n40328), .B(n40329), .Z(n40260) );
  AND U40233 ( .A(n773), .B(n40238), .Z(n40329) );
  XNOR U40234 ( .A(n40236), .B(n40328), .Z(n40238) );
  XNOR U40235 ( .A(n40330), .B(n40331), .Z(n773) );
  AND U40236 ( .A(n40332), .B(n40333), .Z(n40331) );
  XNOR U40237 ( .A(n40330), .B(n40022), .Z(n40333) );
  IV U40238 ( .A(n40026), .Z(n40022) );
  XOR U40239 ( .A(n40334), .B(n40335), .Z(n40026) );
  AND U40240 ( .A(n777), .B(n40336), .Z(n40335) );
  XOR U40241 ( .A(n40337), .B(n40334), .Z(n40336) );
  XNOR U40242 ( .A(n40330), .B(n40243), .Z(n40332) );
  XOR U40243 ( .A(n40338), .B(n40339), .Z(n40243) );
  AND U40244 ( .A(n785), .B(n40290), .Z(n40339) );
  XOR U40245 ( .A(n40288), .B(n40338), .Z(n40290) );
  XOR U40246 ( .A(n40340), .B(n40341), .Z(n40330) );
  AND U40247 ( .A(n40342), .B(n40343), .Z(n40341) );
  XNOR U40248 ( .A(n40340), .B(n40038), .Z(n40343) );
  IV U40249 ( .A(n40041), .Z(n40038) );
  XOR U40250 ( .A(n40344), .B(n40345), .Z(n40041) );
  AND U40251 ( .A(n777), .B(n40346), .Z(n40345) );
  XOR U40252 ( .A(n40347), .B(n40344), .Z(n40346) );
  XOR U40253 ( .A(n40042), .B(n40340), .Z(n40342) );
  XOR U40254 ( .A(n40348), .B(n40349), .Z(n40042) );
  AND U40255 ( .A(n785), .B(n40300), .Z(n40349) );
  XOR U40256 ( .A(n40348), .B(n40298), .Z(n40300) );
  XOR U40257 ( .A(n40350), .B(n40351), .Z(n40340) );
  AND U40258 ( .A(n40352), .B(n40353), .Z(n40351) );
  XNOR U40259 ( .A(n40350), .B(n40066), .Z(n40353) );
  IV U40260 ( .A(n40069), .Z(n40066) );
  XOR U40261 ( .A(n40354), .B(n40355), .Z(n40069) );
  AND U40262 ( .A(n777), .B(n40356), .Z(n40355) );
  XNOR U40263 ( .A(n40357), .B(n40354), .Z(n40356) );
  XOR U40264 ( .A(n40070), .B(n40350), .Z(n40352) );
  XOR U40265 ( .A(n40358), .B(n40359), .Z(n40070) );
  AND U40266 ( .A(n785), .B(n40309), .Z(n40359) );
  XOR U40267 ( .A(n40358), .B(n40307), .Z(n40309) );
  XOR U40268 ( .A(n40360), .B(n40361), .Z(n40350) );
  AND U40269 ( .A(n40362), .B(n40363), .Z(n40361) );
  XNOR U40270 ( .A(n40360), .B(n40115), .Z(n40363) );
  IV U40271 ( .A(n40118), .Z(n40115) );
  XOR U40272 ( .A(n40364), .B(n40365), .Z(n40118) );
  AND U40273 ( .A(n777), .B(n40366), .Z(n40365) );
  XOR U40274 ( .A(n40367), .B(n40364), .Z(n40366) );
  XOR U40275 ( .A(n40119), .B(n40360), .Z(n40362) );
  XOR U40276 ( .A(n40368), .B(n40369), .Z(n40119) );
  AND U40277 ( .A(n785), .B(n40317), .Z(n40369) );
  XOR U40278 ( .A(n40368), .B(n40315), .Z(n40317) );
  XOR U40279 ( .A(n40256), .B(n40370), .Z(n40360) );
  AND U40280 ( .A(n40258), .B(n40371), .Z(n40370) );
  XNOR U40281 ( .A(n40256), .B(n40212), .Z(n40371) );
  IV U40282 ( .A(n40215), .Z(n40212) );
  XOR U40283 ( .A(n40372), .B(n40373), .Z(n40215) );
  AND U40284 ( .A(n777), .B(n40374), .Z(n40373) );
  XNOR U40285 ( .A(n40375), .B(n40372), .Z(n40374) );
  XOR U40286 ( .A(n40216), .B(n40256), .Z(n40258) );
  XOR U40287 ( .A(n40376), .B(n40377), .Z(n40216) );
  AND U40288 ( .A(n785), .B(n40327), .Z(n40377) );
  XOR U40289 ( .A(n40376), .B(n40325), .Z(n40327) );
  AND U40290 ( .A(n40328), .B(n40236), .Z(n40256) );
  XNOR U40291 ( .A(n40378), .B(n40379), .Z(n40236) );
  AND U40292 ( .A(n777), .B(n40380), .Z(n40379) );
  XNOR U40293 ( .A(n40381), .B(n40378), .Z(n40380) );
  XNOR U40294 ( .A(n40382), .B(n40383), .Z(n777) );
  AND U40295 ( .A(n40384), .B(n40385), .Z(n40383) );
  XOR U40296 ( .A(n40337), .B(n40382), .Z(n40385) );
  AND U40297 ( .A(n40386), .B(n40387), .Z(n40337) );
  XNOR U40298 ( .A(n40334), .B(n40382), .Z(n40384) );
  XNOR U40299 ( .A(n40388), .B(n40389), .Z(n40334) );
  AND U40300 ( .A(n781), .B(n40390), .Z(n40389) );
  XNOR U40301 ( .A(n40391), .B(n40392), .Z(n40390) );
  XOR U40302 ( .A(n40393), .B(n40394), .Z(n40382) );
  AND U40303 ( .A(n40395), .B(n40396), .Z(n40394) );
  XNOR U40304 ( .A(n40393), .B(n40386), .Z(n40396) );
  IV U40305 ( .A(n40347), .Z(n40386) );
  XOR U40306 ( .A(n40397), .B(n40398), .Z(n40347) );
  XOR U40307 ( .A(n40399), .B(n40387), .Z(n40398) );
  AND U40308 ( .A(n40357), .B(n40400), .Z(n40387) );
  AND U40309 ( .A(n40401), .B(n40402), .Z(n40399) );
  XOR U40310 ( .A(n40403), .B(n40397), .Z(n40401) );
  XNOR U40311 ( .A(n40344), .B(n40393), .Z(n40395) );
  XNOR U40312 ( .A(n40404), .B(n40405), .Z(n40344) );
  AND U40313 ( .A(n781), .B(n40406), .Z(n40405) );
  XNOR U40314 ( .A(n40407), .B(n40408), .Z(n40406) );
  XOR U40315 ( .A(n40409), .B(n40410), .Z(n40393) );
  AND U40316 ( .A(n40411), .B(n40412), .Z(n40410) );
  XNOR U40317 ( .A(n40409), .B(n40357), .Z(n40412) );
  XOR U40318 ( .A(n40413), .B(n40402), .Z(n40357) );
  XNOR U40319 ( .A(n40414), .B(n40397), .Z(n40402) );
  XOR U40320 ( .A(n40415), .B(n40416), .Z(n40397) );
  AND U40321 ( .A(n40417), .B(n40418), .Z(n40416) );
  XOR U40322 ( .A(n40419), .B(n40415), .Z(n40417) );
  XNOR U40323 ( .A(n40420), .B(n40421), .Z(n40414) );
  AND U40324 ( .A(n40422), .B(n40423), .Z(n40421) );
  XOR U40325 ( .A(n40420), .B(n40424), .Z(n40422) );
  XNOR U40326 ( .A(n40403), .B(n40400), .Z(n40413) );
  AND U40327 ( .A(n40425), .B(n40426), .Z(n40400) );
  XOR U40328 ( .A(n40427), .B(n40428), .Z(n40403) );
  AND U40329 ( .A(n40429), .B(n40430), .Z(n40428) );
  XOR U40330 ( .A(n40427), .B(n40431), .Z(n40429) );
  XNOR U40331 ( .A(n40354), .B(n40409), .Z(n40411) );
  XNOR U40332 ( .A(n40432), .B(n40433), .Z(n40354) );
  AND U40333 ( .A(n781), .B(n40434), .Z(n40433) );
  XNOR U40334 ( .A(n40435), .B(n40436), .Z(n40434) );
  XOR U40335 ( .A(n40437), .B(n40438), .Z(n40409) );
  AND U40336 ( .A(n40439), .B(n40440), .Z(n40438) );
  XNOR U40337 ( .A(n40437), .B(n40425), .Z(n40440) );
  IV U40338 ( .A(n40367), .Z(n40425) );
  XNOR U40339 ( .A(n40441), .B(n40418), .Z(n40367) );
  XNOR U40340 ( .A(n40442), .B(n40424), .Z(n40418) );
  XOR U40341 ( .A(n40443), .B(n40444), .Z(n40424) );
  AND U40342 ( .A(n40445), .B(n40446), .Z(n40444) );
  XOR U40343 ( .A(n40443), .B(n40447), .Z(n40445) );
  XNOR U40344 ( .A(n40423), .B(n40415), .Z(n40442) );
  XOR U40345 ( .A(n40448), .B(n40449), .Z(n40415) );
  AND U40346 ( .A(n40450), .B(n40451), .Z(n40449) );
  XNOR U40347 ( .A(n40452), .B(n40448), .Z(n40450) );
  XNOR U40348 ( .A(n40453), .B(n40420), .Z(n40423) );
  XOR U40349 ( .A(n40454), .B(n40455), .Z(n40420) );
  AND U40350 ( .A(n40456), .B(n40457), .Z(n40455) );
  XOR U40351 ( .A(n40454), .B(n40458), .Z(n40456) );
  XNOR U40352 ( .A(n40459), .B(n40460), .Z(n40453) );
  AND U40353 ( .A(n40461), .B(n40462), .Z(n40460) );
  XNOR U40354 ( .A(n40459), .B(n40463), .Z(n40461) );
  XNOR U40355 ( .A(n40419), .B(n40426), .Z(n40441) );
  AND U40356 ( .A(n40375), .B(n40464), .Z(n40426) );
  XOR U40357 ( .A(n40431), .B(n40430), .Z(n40419) );
  XNOR U40358 ( .A(n40465), .B(n40427), .Z(n40430) );
  XOR U40359 ( .A(n40466), .B(n40467), .Z(n40427) );
  AND U40360 ( .A(n40468), .B(n40469), .Z(n40467) );
  XOR U40361 ( .A(n40466), .B(n40470), .Z(n40468) );
  XNOR U40362 ( .A(n40471), .B(n40472), .Z(n40465) );
  AND U40363 ( .A(n40473), .B(n40474), .Z(n40472) );
  XOR U40364 ( .A(n40471), .B(n40475), .Z(n40473) );
  XOR U40365 ( .A(n40476), .B(n40477), .Z(n40431) );
  AND U40366 ( .A(n40478), .B(n40479), .Z(n40477) );
  XOR U40367 ( .A(n40476), .B(n40480), .Z(n40478) );
  XNOR U40368 ( .A(n40364), .B(n40437), .Z(n40439) );
  XNOR U40369 ( .A(n40481), .B(n40482), .Z(n40364) );
  AND U40370 ( .A(n781), .B(n40483), .Z(n40482) );
  XNOR U40371 ( .A(n40484), .B(n40485), .Z(n40483) );
  XOR U40372 ( .A(n40486), .B(n40487), .Z(n40437) );
  AND U40373 ( .A(n40488), .B(n40489), .Z(n40487) );
  XNOR U40374 ( .A(n40486), .B(n40375), .Z(n40489) );
  XOR U40375 ( .A(n40490), .B(n40451), .Z(n40375) );
  XNOR U40376 ( .A(n40491), .B(n40458), .Z(n40451) );
  XOR U40377 ( .A(n40447), .B(n40446), .Z(n40458) );
  XNOR U40378 ( .A(n40492), .B(n40443), .Z(n40446) );
  XOR U40379 ( .A(n40493), .B(n40494), .Z(n40443) );
  AND U40380 ( .A(n40495), .B(n40496), .Z(n40494) );
  XNOR U40381 ( .A(n40497), .B(n40498), .Z(n40495) );
  IV U40382 ( .A(n40493), .Z(n40497) );
  XNOR U40383 ( .A(n40499), .B(n40500), .Z(n40492) );
  NOR U40384 ( .A(n40501), .B(n40502), .Z(n40500) );
  XNOR U40385 ( .A(n40499), .B(n40503), .Z(n40501) );
  XOR U40386 ( .A(n40504), .B(n40505), .Z(n40447) );
  NOR U40387 ( .A(n40506), .B(n40507), .Z(n40505) );
  XNOR U40388 ( .A(n40504), .B(n40508), .Z(n40506) );
  XNOR U40389 ( .A(n40457), .B(n40448), .Z(n40491) );
  XOR U40390 ( .A(n40509), .B(n40510), .Z(n40448) );
  AND U40391 ( .A(n40511), .B(n40512), .Z(n40510) );
  XOR U40392 ( .A(n40509), .B(n40513), .Z(n40511) );
  XOR U40393 ( .A(n40514), .B(n40463), .Z(n40457) );
  XOR U40394 ( .A(n40515), .B(n40516), .Z(n40463) );
  NOR U40395 ( .A(n40517), .B(n40518), .Z(n40516) );
  XOR U40396 ( .A(n40515), .B(n40519), .Z(n40517) );
  XNOR U40397 ( .A(n40462), .B(n40454), .Z(n40514) );
  XOR U40398 ( .A(n40520), .B(n40521), .Z(n40454) );
  AND U40399 ( .A(n40522), .B(n40523), .Z(n40521) );
  XOR U40400 ( .A(n40520), .B(n40524), .Z(n40522) );
  XNOR U40401 ( .A(n40525), .B(n40459), .Z(n40462) );
  XOR U40402 ( .A(n40526), .B(n40527), .Z(n40459) );
  AND U40403 ( .A(n40528), .B(n40529), .Z(n40527) );
  XNOR U40404 ( .A(n40530), .B(n40531), .Z(n40528) );
  IV U40405 ( .A(n40526), .Z(n40530) );
  XNOR U40406 ( .A(n40532), .B(n40533), .Z(n40525) );
  NOR U40407 ( .A(n40534), .B(n40535), .Z(n40533) );
  XNOR U40408 ( .A(n40532), .B(n40536), .Z(n40534) );
  XOR U40409 ( .A(n40452), .B(n40464), .Z(n40490) );
  NOR U40410 ( .A(n40381), .B(n40537), .Z(n40464) );
  XNOR U40411 ( .A(n40470), .B(n40469), .Z(n40452) );
  XNOR U40412 ( .A(n40538), .B(n40475), .Z(n40469) );
  XNOR U40413 ( .A(n40539), .B(n40540), .Z(n40475) );
  NOR U40414 ( .A(n40541), .B(n40542), .Z(n40540) );
  XOR U40415 ( .A(n40539), .B(n40543), .Z(n40541) );
  XNOR U40416 ( .A(n40474), .B(n40466), .Z(n40538) );
  XOR U40417 ( .A(n40544), .B(n40545), .Z(n40466) );
  AND U40418 ( .A(n40546), .B(n40547), .Z(n40545) );
  XOR U40419 ( .A(n40544), .B(n40548), .Z(n40546) );
  XNOR U40420 ( .A(n40549), .B(n40471), .Z(n40474) );
  XOR U40421 ( .A(n40550), .B(n40551), .Z(n40471) );
  AND U40422 ( .A(n40552), .B(n40553), .Z(n40551) );
  XNOR U40423 ( .A(n40554), .B(n40555), .Z(n40552) );
  IV U40424 ( .A(n40550), .Z(n40554) );
  XNOR U40425 ( .A(n40556), .B(n40557), .Z(n40549) );
  NOR U40426 ( .A(n40558), .B(n40559), .Z(n40557) );
  XNOR U40427 ( .A(n40556), .B(n40560), .Z(n40558) );
  XOR U40428 ( .A(n40480), .B(n40479), .Z(n40470) );
  XNOR U40429 ( .A(n40561), .B(n40476), .Z(n40479) );
  XOR U40430 ( .A(n40562), .B(n40563), .Z(n40476) );
  AND U40431 ( .A(n40564), .B(n40565), .Z(n40563) );
  XNOR U40432 ( .A(n40566), .B(n40567), .Z(n40564) );
  IV U40433 ( .A(n40562), .Z(n40566) );
  XNOR U40434 ( .A(n40568), .B(n40569), .Z(n40561) );
  NOR U40435 ( .A(n40570), .B(n40571), .Z(n40569) );
  XNOR U40436 ( .A(n40568), .B(n40572), .Z(n40570) );
  XOR U40437 ( .A(n40573), .B(n40574), .Z(n40480) );
  NOR U40438 ( .A(n40575), .B(n40576), .Z(n40574) );
  XNOR U40439 ( .A(n40573), .B(n40577), .Z(n40575) );
  XNOR U40440 ( .A(n40372), .B(n40486), .Z(n40488) );
  XNOR U40441 ( .A(n40578), .B(n40579), .Z(n40372) );
  AND U40442 ( .A(n781), .B(n40580), .Z(n40579) );
  XNOR U40443 ( .A(n40581), .B(n40582), .Z(n40580) );
  AND U40444 ( .A(n40378), .B(n40381), .Z(n40486) );
  XOR U40445 ( .A(n40583), .B(n40537), .Z(n40381) );
  XNOR U40446 ( .A(p_input[1088]), .B(p_input[2048]), .Z(n40537) );
  XNOR U40447 ( .A(n40513), .B(n40512), .Z(n40583) );
  XNOR U40448 ( .A(n40584), .B(n40524), .Z(n40512) );
  XOR U40449 ( .A(n40498), .B(n40496), .Z(n40524) );
  XNOR U40450 ( .A(n40585), .B(n40503), .Z(n40496) );
  XOR U40451 ( .A(p_input[1112]), .B(p_input[2072]), .Z(n40503) );
  XOR U40452 ( .A(n40493), .B(n40502), .Z(n40585) );
  XOR U40453 ( .A(n40586), .B(n40499), .Z(n40502) );
  XOR U40454 ( .A(p_input[1110]), .B(p_input[2070]), .Z(n40499) );
  XOR U40455 ( .A(p_input[1111]), .B(n29410), .Z(n40586) );
  XOR U40456 ( .A(p_input[1106]), .B(p_input[2066]), .Z(n40493) );
  XNOR U40457 ( .A(n40508), .B(n40507), .Z(n40498) );
  XOR U40458 ( .A(n40587), .B(n40504), .Z(n40507) );
  XOR U40459 ( .A(p_input[1107]), .B(p_input[2067]), .Z(n40504) );
  XOR U40460 ( .A(p_input[1108]), .B(n29412), .Z(n40587) );
  XOR U40461 ( .A(p_input[1109]), .B(p_input[2069]), .Z(n40508) );
  XOR U40462 ( .A(n40523), .B(n40588), .Z(n40584) );
  IV U40463 ( .A(n40509), .Z(n40588) );
  XOR U40464 ( .A(p_input[1089]), .B(p_input[2049]), .Z(n40509) );
  XNOR U40465 ( .A(n40589), .B(n40531), .Z(n40523) );
  XNOR U40466 ( .A(n40519), .B(n40518), .Z(n40531) );
  XNOR U40467 ( .A(n40590), .B(n40515), .Z(n40518) );
  XNOR U40468 ( .A(p_input[1114]), .B(p_input[2074]), .Z(n40515) );
  XOR U40469 ( .A(p_input[1115]), .B(n29415), .Z(n40590) );
  XOR U40470 ( .A(p_input[1116]), .B(p_input[2076]), .Z(n40519) );
  XOR U40471 ( .A(n40529), .B(n40591), .Z(n40589) );
  IV U40472 ( .A(n40520), .Z(n40591) );
  XOR U40473 ( .A(p_input[1105]), .B(p_input[2065]), .Z(n40520) );
  XNOR U40474 ( .A(n40592), .B(n40536), .Z(n40529) );
  XNOR U40475 ( .A(p_input[1119]), .B(n29418), .Z(n40536) );
  XOR U40476 ( .A(n40526), .B(n40535), .Z(n40592) );
  XOR U40477 ( .A(n40593), .B(n40532), .Z(n40535) );
  XOR U40478 ( .A(p_input[1117]), .B(p_input[2077]), .Z(n40532) );
  XOR U40479 ( .A(p_input[1118]), .B(n29420), .Z(n40593) );
  XOR U40480 ( .A(p_input[1113]), .B(p_input[2073]), .Z(n40526) );
  XOR U40481 ( .A(n40548), .B(n40547), .Z(n40513) );
  XNOR U40482 ( .A(n40594), .B(n40555), .Z(n40547) );
  XNOR U40483 ( .A(n40543), .B(n40542), .Z(n40555) );
  XNOR U40484 ( .A(n40595), .B(n40539), .Z(n40542) );
  XNOR U40485 ( .A(p_input[1099]), .B(p_input[2059]), .Z(n40539) );
  XOR U40486 ( .A(p_input[1100]), .B(n28329), .Z(n40595) );
  XOR U40487 ( .A(p_input[1101]), .B(p_input[2061]), .Z(n40543) );
  XOR U40488 ( .A(n40553), .B(n40596), .Z(n40594) );
  IV U40489 ( .A(n40544), .Z(n40596) );
  XOR U40490 ( .A(p_input[1090]), .B(p_input[2050]), .Z(n40544) );
  XNOR U40491 ( .A(n40597), .B(n40560), .Z(n40553) );
  XNOR U40492 ( .A(p_input[1104]), .B(n28332), .Z(n40560) );
  XOR U40493 ( .A(n40550), .B(n40559), .Z(n40597) );
  XOR U40494 ( .A(n40598), .B(n40556), .Z(n40559) );
  XOR U40495 ( .A(p_input[1102]), .B(p_input[2062]), .Z(n40556) );
  XOR U40496 ( .A(p_input[1103]), .B(n28334), .Z(n40598) );
  XOR U40497 ( .A(p_input[1098]), .B(p_input[2058]), .Z(n40550) );
  XOR U40498 ( .A(n40567), .B(n40565), .Z(n40548) );
  XNOR U40499 ( .A(n40599), .B(n40572), .Z(n40565) );
  XOR U40500 ( .A(p_input[1097]), .B(p_input[2057]), .Z(n40572) );
  XOR U40501 ( .A(n40562), .B(n40571), .Z(n40599) );
  XOR U40502 ( .A(n40600), .B(n40568), .Z(n40571) );
  XOR U40503 ( .A(p_input[1095]), .B(p_input[2055]), .Z(n40568) );
  XOR U40504 ( .A(p_input[1096]), .B(n29427), .Z(n40600) );
  XOR U40505 ( .A(p_input[1091]), .B(p_input[2051]), .Z(n40562) );
  XNOR U40506 ( .A(n40577), .B(n40576), .Z(n40567) );
  XOR U40507 ( .A(n40601), .B(n40573), .Z(n40576) );
  XOR U40508 ( .A(p_input[1092]), .B(p_input[2052]), .Z(n40573) );
  XOR U40509 ( .A(p_input[1093]), .B(n29429), .Z(n40601) );
  XOR U40510 ( .A(p_input[1094]), .B(p_input[2054]), .Z(n40577) );
  XNOR U40511 ( .A(n40602), .B(n40603), .Z(n40378) );
  AND U40512 ( .A(n781), .B(n40604), .Z(n40603) );
  XNOR U40513 ( .A(n40605), .B(n40606), .Z(n781) );
  AND U40514 ( .A(n40607), .B(n40608), .Z(n40606) );
  XOR U40515 ( .A(n40392), .B(n40605), .Z(n40608) );
  XNOR U40516 ( .A(n40609), .B(n40605), .Z(n40607) );
  XOR U40517 ( .A(n40610), .B(n40611), .Z(n40605) );
  AND U40518 ( .A(n40612), .B(n40613), .Z(n40611) );
  XOR U40519 ( .A(n40407), .B(n40610), .Z(n40613) );
  XOR U40520 ( .A(n40610), .B(n40408), .Z(n40612) );
  XOR U40521 ( .A(n40614), .B(n40615), .Z(n40610) );
  AND U40522 ( .A(n40616), .B(n40617), .Z(n40615) );
  XOR U40523 ( .A(n40435), .B(n40614), .Z(n40617) );
  XOR U40524 ( .A(n40614), .B(n40436), .Z(n40616) );
  XOR U40525 ( .A(n40618), .B(n40619), .Z(n40614) );
  AND U40526 ( .A(n40620), .B(n40621), .Z(n40619) );
  XOR U40527 ( .A(n40484), .B(n40618), .Z(n40621) );
  XOR U40528 ( .A(n40618), .B(n40485), .Z(n40620) );
  XOR U40529 ( .A(n40622), .B(n40623), .Z(n40618) );
  AND U40530 ( .A(n40624), .B(n40625), .Z(n40623) );
  XOR U40531 ( .A(n40622), .B(n40581), .Z(n40625) );
  XNOR U40532 ( .A(n40626), .B(n40627), .Z(n40328) );
  AND U40533 ( .A(n785), .B(n40628), .Z(n40627) );
  XNOR U40534 ( .A(n40629), .B(n40630), .Z(n785) );
  AND U40535 ( .A(n40631), .B(n40632), .Z(n40630) );
  XOR U40536 ( .A(n40629), .B(n40338), .Z(n40632) );
  XNOR U40537 ( .A(n40629), .B(n40288), .Z(n40631) );
  XOR U40538 ( .A(n40633), .B(n40634), .Z(n40629) );
  AND U40539 ( .A(n40635), .B(n40636), .Z(n40634) );
  XNOR U40540 ( .A(n40348), .B(n40633), .Z(n40636) );
  XOR U40541 ( .A(n40633), .B(n40298), .Z(n40635) );
  XOR U40542 ( .A(n40637), .B(n40638), .Z(n40633) );
  AND U40543 ( .A(n40639), .B(n40640), .Z(n40638) );
  XNOR U40544 ( .A(n40358), .B(n40637), .Z(n40640) );
  XOR U40545 ( .A(n40637), .B(n40307), .Z(n40639) );
  XOR U40546 ( .A(n40641), .B(n40642), .Z(n40637) );
  AND U40547 ( .A(n40643), .B(n40644), .Z(n40642) );
  XOR U40548 ( .A(n40641), .B(n40315), .Z(n40643) );
  XOR U40549 ( .A(n40645), .B(n40646), .Z(n40279) );
  AND U40550 ( .A(n789), .B(n40628), .Z(n40646) );
  XNOR U40551 ( .A(n40626), .B(n40645), .Z(n40628) );
  XNOR U40552 ( .A(n40647), .B(n40648), .Z(n789) );
  AND U40553 ( .A(n40649), .B(n40650), .Z(n40648) );
  XNOR U40554 ( .A(n40651), .B(n40647), .Z(n40650) );
  IV U40555 ( .A(n40338), .Z(n40651) );
  XOR U40556 ( .A(n40609), .B(n40652), .Z(n40338) );
  AND U40557 ( .A(n792), .B(n40653), .Z(n40652) );
  XOR U40558 ( .A(n40391), .B(n40388), .Z(n40653) );
  IV U40559 ( .A(n40609), .Z(n40391) );
  XNOR U40560 ( .A(n40288), .B(n40647), .Z(n40649) );
  XOR U40561 ( .A(n40654), .B(n40655), .Z(n40288) );
  AND U40562 ( .A(n808), .B(n40656), .Z(n40655) );
  XOR U40563 ( .A(n40657), .B(n40658), .Z(n40647) );
  AND U40564 ( .A(n40659), .B(n40660), .Z(n40658) );
  XNOR U40565 ( .A(n40657), .B(n40348), .Z(n40660) );
  XOR U40566 ( .A(n40408), .B(n40661), .Z(n40348) );
  AND U40567 ( .A(n792), .B(n40662), .Z(n40661) );
  XOR U40568 ( .A(n40404), .B(n40408), .Z(n40662) );
  XNOR U40569 ( .A(n40663), .B(n40657), .Z(n40659) );
  IV U40570 ( .A(n40298), .Z(n40663) );
  XOR U40571 ( .A(n40664), .B(n40665), .Z(n40298) );
  AND U40572 ( .A(n808), .B(n40666), .Z(n40665) );
  XOR U40573 ( .A(n40667), .B(n40668), .Z(n40657) );
  AND U40574 ( .A(n40669), .B(n40670), .Z(n40668) );
  XNOR U40575 ( .A(n40667), .B(n40358), .Z(n40670) );
  XOR U40576 ( .A(n40436), .B(n40671), .Z(n40358) );
  AND U40577 ( .A(n792), .B(n40672), .Z(n40671) );
  XOR U40578 ( .A(n40432), .B(n40436), .Z(n40672) );
  XOR U40579 ( .A(n40307), .B(n40667), .Z(n40669) );
  XOR U40580 ( .A(n40673), .B(n40674), .Z(n40307) );
  AND U40581 ( .A(n808), .B(n40675), .Z(n40674) );
  XOR U40582 ( .A(n40641), .B(n40676), .Z(n40667) );
  AND U40583 ( .A(n40677), .B(n40644), .Z(n40676) );
  XNOR U40584 ( .A(n40368), .B(n40641), .Z(n40644) );
  XOR U40585 ( .A(n40485), .B(n40678), .Z(n40368) );
  AND U40586 ( .A(n792), .B(n40679), .Z(n40678) );
  XOR U40587 ( .A(n40481), .B(n40485), .Z(n40679) );
  XNOR U40588 ( .A(n40680), .B(n40641), .Z(n40677) );
  IV U40589 ( .A(n40315), .Z(n40680) );
  XOR U40590 ( .A(n40681), .B(n40682), .Z(n40315) );
  AND U40591 ( .A(n808), .B(n40683), .Z(n40682) );
  XOR U40592 ( .A(n40684), .B(n40685), .Z(n40641) );
  AND U40593 ( .A(n40686), .B(n40687), .Z(n40685) );
  XNOR U40594 ( .A(n40684), .B(n40376), .Z(n40687) );
  XOR U40595 ( .A(n40582), .B(n40688), .Z(n40376) );
  AND U40596 ( .A(n792), .B(n40689), .Z(n40688) );
  XOR U40597 ( .A(n40578), .B(n40582), .Z(n40689) );
  XNOR U40598 ( .A(n40690), .B(n40684), .Z(n40686) );
  IV U40599 ( .A(n40325), .Z(n40690) );
  XOR U40600 ( .A(n40691), .B(n40692), .Z(n40325) );
  AND U40601 ( .A(n808), .B(n40693), .Z(n40692) );
  AND U40602 ( .A(n40645), .B(n40626), .Z(n40684) );
  XNOR U40603 ( .A(n40694), .B(n40695), .Z(n40626) );
  AND U40604 ( .A(n792), .B(n40604), .Z(n40695) );
  XNOR U40605 ( .A(n40602), .B(n40694), .Z(n40604) );
  XNOR U40606 ( .A(n40696), .B(n40697), .Z(n792) );
  AND U40607 ( .A(n40698), .B(n40699), .Z(n40697) );
  XNOR U40608 ( .A(n40696), .B(n40388), .Z(n40699) );
  IV U40609 ( .A(n40392), .Z(n40388) );
  XOR U40610 ( .A(n40700), .B(n40701), .Z(n40392) );
  AND U40611 ( .A(n796), .B(n40702), .Z(n40701) );
  XOR U40612 ( .A(n40703), .B(n40700), .Z(n40702) );
  XNOR U40613 ( .A(n40696), .B(n40609), .Z(n40698) );
  XOR U40614 ( .A(n40704), .B(n40705), .Z(n40609) );
  AND U40615 ( .A(n804), .B(n40656), .Z(n40705) );
  XOR U40616 ( .A(n40654), .B(n40704), .Z(n40656) );
  XOR U40617 ( .A(n40706), .B(n40707), .Z(n40696) );
  AND U40618 ( .A(n40708), .B(n40709), .Z(n40707) );
  XNOR U40619 ( .A(n40706), .B(n40404), .Z(n40709) );
  IV U40620 ( .A(n40407), .Z(n40404) );
  XOR U40621 ( .A(n40710), .B(n40711), .Z(n40407) );
  AND U40622 ( .A(n796), .B(n40712), .Z(n40711) );
  XOR U40623 ( .A(n40713), .B(n40710), .Z(n40712) );
  XOR U40624 ( .A(n40408), .B(n40706), .Z(n40708) );
  XOR U40625 ( .A(n40714), .B(n40715), .Z(n40408) );
  AND U40626 ( .A(n804), .B(n40666), .Z(n40715) );
  XOR U40627 ( .A(n40714), .B(n40664), .Z(n40666) );
  XOR U40628 ( .A(n40716), .B(n40717), .Z(n40706) );
  AND U40629 ( .A(n40718), .B(n40719), .Z(n40717) );
  XNOR U40630 ( .A(n40716), .B(n40432), .Z(n40719) );
  IV U40631 ( .A(n40435), .Z(n40432) );
  XOR U40632 ( .A(n40720), .B(n40721), .Z(n40435) );
  AND U40633 ( .A(n796), .B(n40722), .Z(n40721) );
  XNOR U40634 ( .A(n40723), .B(n40720), .Z(n40722) );
  XOR U40635 ( .A(n40436), .B(n40716), .Z(n40718) );
  XOR U40636 ( .A(n40724), .B(n40725), .Z(n40436) );
  AND U40637 ( .A(n804), .B(n40675), .Z(n40725) );
  XOR U40638 ( .A(n40724), .B(n40673), .Z(n40675) );
  XOR U40639 ( .A(n40726), .B(n40727), .Z(n40716) );
  AND U40640 ( .A(n40728), .B(n40729), .Z(n40727) );
  XNOR U40641 ( .A(n40726), .B(n40481), .Z(n40729) );
  IV U40642 ( .A(n40484), .Z(n40481) );
  XOR U40643 ( .A(n40730), .B(n40731), .Z(n40484) );
  AND U40644 ( .A(n796), .B(n40732), .Z(n40731) );
  XOR U40645 ( .A(n40733), .B(n40730), .Z(n40732) );
  XOR U40646 ( .A(n40485), .B(n40726), .Z(n40728) );
  XOR U40647 ( .A(n40734), .B(n40735), .Z(n40485) );
  AND U40648 ( .A(n804), .B(n40683), .Z(n40735) );
  XOR U40649 ( .A(n40734), .B(n40681), .Z(n40683) );
  XOR U40650 ( .A(n40622), .B(n40736), .Z(n40726) );
  AND U40651 ( .A(n40624), .B(n40737), .Z(n40736) );
  XNOR U40652 ( .A(n40622), .B(n40578), .Z(n40737) );
  IV U40653 ( .A(n40581), .Z(n40578) );
  XOR U40654 ( .A(n40738), .B(n40739), .Z(n40581) );
  AND U40655 ( .A(n796), .B(n40740), .Z(n40739) );
  XNOR U40656 ( .A(n40741), .B(n40738), .Z(n40740) );
  XOR U40657 ( .A(n40582), .B(n40622), .Z(n40624) );
  XOR U40658 ( .A(n40742), .B(n40743), .Z(n40582) );
  AND U40659 ( .A(n804), .B(n40693), .Z(n40743) );
  XOR U40660 ( .A(n40742), .B(n40691), .Z(n40693) );
  AND U40661 ( .A(n40694), .B(n40602), .Z(n40622) );
  XNOR U40662 ( .A(n40744), .B(n40745), .Z(n40602) );
  AND U40663 ( .A(n796), .B(n40746), .Z(n40745) );
  XNOR U40664 ( .A(n40747), .B(n40744), .Z(n40746) );
  XNOR U40665 ( .A(n40748), .B(n40749), .Z(n796) );
  AND U40666 ( .A(n40750), .B(n40751), .Z(n40749) );
  XOR U40667 ( .A(n40703), .B(n40748), .Z(n40751) );
  AND U40668 ( .A(n40752), .B(n40753), .Z(n40703) );
  XNOR U40669 ( .A(n40700), .B(n40748), .Z(n40750) );
  XNOR U40670 ( .A(n40754), .B(n40755), .Z(n40700) );
  AND U40671 ( .A(n800), .B(n40756), .Z(n40755) );
  XNOR U40672 ( .A(n40757), .B(n40758), .Z(n40756) );
  XOR U40673 ( .A(n40759), .B(n40760), .Z(n40748) );
  AND U40674 ( .A(n40761), .B(n40762), .Z(n40760) );
  XNOR U40675 ( .A(n40759), .B(n40752), .Z(n40762) );
  IV U40676 ( .A(n40713), .Z(n40752) );
  XOR U40677 ( .A(n40763), .B(n40764), .Z(n40713) );
  XOR U40678 ( .A(n40765), .B(n40753), .Z(n40764) );
  AND U40679 ( .A(n40723), .B(n40766), .Z(n40753) );
  AND U40680 ( .A(n40767), .B(n40768), .Z(n40765) );
  XOR U40681 ( .A(n40769), .B(n40763), .Z(n40767) );
  XNOR U40682 ( .A(n40710), .B(n40759), .Z(n40761) );
  XNOR U40683 ( .A(n40770), .B(n40771), .Z(n40710) );
  AND U40684 ( .A(n800), .B(n40772), .Z(n40771) );
  XNOR U40685 ( .A(n40773), .B(n40774), .Z(n40772) );
  XOR U40686 ( .A(n40775), .B(n40776), .Z(n40759) );
  AND U40687 ( .A(n40777), .B(n40778), .Z(n40776) );
  XNOR U40688 ( .A(n40775), .B(n40723), .Z(n40778) );
  XOR U40689 ( .A(n40779), .B(n40768), .Z(n40723) );
  XNOR U40690 ( .A(n40780), .B(n40763), .Z(n40768) );
  XOR U40691 ( .A(n40781), .B(n40782), .Z(n40763) );
  AND U40692 ( .A(n40783), .B(n40784), .Z(n40782) );
  XOR U40693 ( .A(n40785), .B(n40781), .Z(n40783) );
  XNOR U40694 ( .A(n40786), .B(n40787), .Z(n40780) );
  AND U40695 ( .A(n40788), .B(n40789), .Z(n40787) );
  XOR U40696 ( .A(n40786), .B(n40790), .Z(n40788) );
  XNOR U40697 ( .A(n40769), .B(n40766), .Z(n40779) );
  AND U40698 ( .A(n40791), .B(n40792), .Z(n40766) );
  XOR U40699 ( .A(n40793), .B(n40794), .Z(n40769) );
  AND U40700 ( .A(n40795), .B(n40796), .Z(n40794) );
  XOR U40701 ( .A(n40793), .B(n40797), .Z(n40795) );
  XNOR U40702 ( .A(n40720), .B(n40775), .Z(n40777) );
  XNOR U40703 ( .A(n40798), .B(n40799), .Z(n40720) );
  AND U40704 ( .A(n800), .B(n40800), .Z(n40799) );
  XNOR U40705 ( .A(n40801), .B(n40802), .Z(n40800) );
  XOR U40706 ( .A(n40803), .B(n40804), .Z(n40775) );
  AND U40707 ( .A(n40805), .B(n40806), .Z(n40804) );
  XNOR U40708 ( .A(n40803), .B(n40791), .Z(n40806) );
  IV U40709 ( .A(n40733), .Z(n40791) );
  XNOR U40710 ( .A(n40807), .B(n40784), .Z(n40733) );
  XNOR U40711 ( .A(n40808), .B(n40790), .Z(n40784) );
  XOR U40712 ( .A(n40809), .B(n40810), .Z(n40790) );
  AND U40713 ( .A(n40811), .B(n40812), .Z(n40810) );
  XOR U40714 ( .A(n40809), .B(n40813), .Z(n40811) );
  XNOR U40715 ( .A(n40789), .B(n40781), .Z(n40808) );
  XOR U40716 ( .A(n40814), .B(n40815), .Z(n40781) );
  AND U40717 ( .A(n40816), .B(n40817), .Z(n40815) );
  XNOR U40718 ( .A(n40818), .B(n40814), .Z(n40816) );
  XNOR U40719 ( .A(n40819), .B(n40786), .Z(n40789) );
  XOR U40720 ( .A(n40820), .B(n40821), .Z(n40786) );
  AND U40721 ( .A(n40822), .B(n40823), .Z(n40821) );
  XOR U40722 ( .A(n40820), .B(n40824), .Z(n40822) );
  XNOR U40723 ( .A(n40825), .B(n40826), .Z(n40819) );
  AND U40724 ( .A(n40827), .B(n40828), .Z(n40826) );
  XNOR U40725 ( .A(n40825), .B(n40829), .Z(n40827) );
  XNOR U40726 ( .A(n40785), .B(n40792), .Z(n40807) );
  AND U40727 ( .A(n40741), .B(n40830), .Z(n40792) );
  XOR U40728 ( .A(n40797), .B(n40796), .Z(n40785) );
  XNOR U40729 ( .A(n40831), .B(n40793), .Z(n40796) );
  XOR U40730 ( .A(n40832), .B(n40833), .Z(n40793) );
  AND U40731 ( .A(n40834), .B(n40835), .Z(n40833) );
  XOR U40732 ( .A(n40832), .B(n40836), .Z(n40834) );
  XNOR U40733 ( .A(n40837), .B(n40838), .Z(n40831) );
  AND U40734 ( .A(n40839), .B(n40840), .Z(n40838) );
  XOR U40735 ( .A(n40837), .B(n40841), .Z(n40839) );
  XOR U40736 ( .A(n40842), .B(n40843), .Z(n40797) );
  AND U40737 ( .A(n40844), .B(n40845), .Z(n40843) );
  XOR U40738 ( .A(n40842), .B(n40846), .Z(n40844) );
  XNOR U40739 ( .A(n40730), .B(n40803), .Z(n40805) );
  XNOR U40740 ( .A(n40847), .B(n40848), .Z(n40730) );
  AND U40741 ( .A(n800), .B(n40849), .Z(n40848) );
  XNOR U40742 ( .A(n40850), .B(n40851), .Z(n40849) );
  XOR U40743 ( .A(n40852), .B(n40853), .Z(n40803) );
  AND U40744 ( .A(n40854), .B(n40855), .Z(n40853) );
  XNOR U40745 ( .A(n40852), .B(n40741), .Z(n40855) );
  XOR U40746 ( .A(n40856), .B(n40817), .Z(n40741) );
  XNOR U40747 ( .A(n40857), .B(n40824), .Z(n40817) );
  XOR U40748 ( .A(n40813), .B(n40812), .Z(n40824) );
  XNOR U40749 ( .A(n40858), .B(n40809), .Z(n40812) );
  XOR U40750 ( .A(n40859), .B(n40860), .Z(n40809) );
  AND U40751 ( .A(n40861), .B(n40862), .Z(n40860) );
  XNOR U40752 ( .A(n40863), .B(n40864), .Z(n40861) );
  IV U40753 ( .A(n40859), .Z(n40863) );
  XNOR U40754 ( .A(n40865), .B(n40866), .Z(n40858) );
  NOR U40755 ( .A(n40867), .B(n40868), .Z(n40866) );
  XNOR U40756 ( .A(n40865), .B(n40869), .Z(n40867) );
  XOR U40757 ( .A(n40870), .B(n40871), .Z(n40813) );
  NOR U40758 ( .A(n40872), .B(n40873), .Z(n40871) );
  XNOR U40759 ( .A(n40870), .B(n40874), .Z(n40872) );
  XNOR U40760 ( .A(n40823), .B(n40814), .Z(n40857) );
  XOR U40761 ( .A(n40875), .B(n40876), .Z(n40814) );
  AND U40762 ( .A(n40877), .B(n40878), .Z(n40876) );
  XOR U40763 ( .A(n40875), .B(n40879), .Z(n40877) );
  XOR U40764 ( .A(n40880), .B(n40829), .Z(n40823) );
  XOR U40765 ( .A(n40881), .B(n40882), .Z(n40829) );
  NOR U40766 ( .A(n40883), .B(n40884), .Z(n40882) );
  XOR U40767 ( .A(n40881), .B(n40885), .Z(n40883) );
  XNOR U40768 ( .A(n40828), .B(n40820), .Z(n40880) );
  XOR U40769 ( .A(n40886), .B(n40887), .Z(n40820) );
  AND U40770 ( .A(n40888), .B(n40889), .Z(n40887) );
  XOR U40771 ( .A(n40886), .B(n40890), .Z(n40888) );
  XNOR U40772 ( .A(n40891), .B(n40825), .Z(n40828) );
  XOR U40773 ( .A(n40892), .B(n40893), .Z(n40825) );
  AND U40774 ( .A(n40894), .B(n40895), .Z(n40893) );
  XNOR U40775 ( .A(n40896), .B(n40897), .Z(n40894) );
  IV U40776 ( .A(n40892), .Z(n40896) );
  XNOR U40777 ( .A(n40898), .B(n40899), .Z(n40891) );
  NOR U40778 ( .A(n40900), .B(n40901), .Z(n40899) );
  XNOR U40779 ( .A(n40898), .B(n40902), .Z(n40900) );
  XOR U40780 ( .A(n40818), .B(n40830), .Z(n40856) );
  NOR U40781 ( .A(n40747), .B(n40903), .Z(n40830) );
  XNOR U40782 ( .A(n40836), .B(n40835), .Z(n40818) );
  XNOR U40783 ( .A(n40904), .B(n40841), .Z(n40835) );
  XNOR U40784 ( .A(n40905), .B(n40906), .Z(n40841) );
  NOR U40785 ( .A(n40907), .B(n40908), .Z(n40906) );
  XOR U40786 ( .A(n40905), .B(n40909), .Z(n40907) );
  XNOR U40787 ( .A(n40840), .B(n40832), .Z(n40904) );
  XOR U40788 ( .A(n40910), .B(n40911), .Z(n40832) );
  AND U40789 ( .A(n40912), .B(n40913), .Z(n40911) );
  XOR U40790 ( .A(n40910), .B(n40914), .Z(n40912) );
  XNOR U40791 ( .A(n40915), .B(n40837), .Z(n40840) );
  XOR U40792 ( .A(n40916), .B(n40917), .Z(n40837) );
  AND U40793 ( .A(n40918), .B(n40919), .Z(n40917) );
  XNOR U40794 ( .A(n40920), .B(n40921), .Z(n40918) );
  IV U40795 ( .A(n40916), .Z(n40920) );
  XNOR U40796 ( .A(n40922), .B(n40923), .Z(n40915) );
  NOR U40797 ( .A(n40924), .B(n40925), .Z(n40923) );
  XNOR U40798 ( .A(n40922), .B(n40926), .Z(n40924) );
  XOR U40799 ( .A(n40846), .B(n40845), .Z(n40836) );
  XNOR U40800 ( .A(n40927), .B(n40842), .Z(n40845) );
  XOR U40801 ( .A(n40928), .B(n40929), .Z(n40842) );
  AND U40802 ( .A(n40930), .B(n40931), .Z(n40929) );
  XNOR U40803 ( .A(n40932), .B(n40933), .Z(n40930) );
  IV U40804 ( .A(n40928), .Z(n40932) );
  XNOR U40805 ( .A(n40934), .B(n40935), .Z(n40927) );
  NOR U40806 ( .A(n40936), .B(n40937), .Z(n40935) );
  XNOR U40807 ( .A(n40934), .B(n40938), .Z(n40936) );
  XOR U40808 ( .A(n40939), .B(n40940), .Z(n40846) );
  NOR U40809 ( .A(n40941), .B(n40942), .Z(n40940) );
  XNOR U40810 ( .A(n40939), .B(n40943), .Z(n40941) );
  XNOR U40811 ( .A(n40738), .B(n40852), .Z(n40854) );
  XNOR U40812 ( .A(n40944), .B(n40945), .Z(n40738) );
  AND U40813 ( .A(n800), .B(n40946), .Z(n40945) );
  XNOR U40814 ( .A(n40947), .B(n40948), .Z(n40946) );
  AND U40815 ( .A(n40744), .B(n40747), .Z(n40852) );
  XOR U40816 ( .A(n40949), .B(n40903), .Z(n40747) );
  XNOR U40817 ( .A(p_input[1120]), .B(p_input[2048]), .Z(n40903) );
  XNOR U40818 ( .A(n40879), .B(n40878), .Z(n40949) );
  XNOR U40819 ( .A(n40950), .B(n40890), .Z(n40878) );
  XOR U40820 ( .A(n40864), .B(n40862), .Z(n40890) );
  XNOR U40821 ( .A(n40951), .B(n40869), .Z(n40862) );
  XOR U40822 ( .A(p_input[1144]), .B(p_input[2072]), .Z(n40869) );
  XOR U40823 ( .A(n40859), .B(n40868), .Z(n40951) );
  XOR U40824 ( .A(n40952), .B(n40865), .Z(n40868) );
  XOR U40825 ( .A(p_input[1142]), .B(p_input[2070]), .Z(n40865) );
  XOR U40826 ( .A(p_input[1143]), .B(n29410), .Z(n40952) );
  XOR U40827 ( .A(p_input[1138]), .B(p_input[2066]), .Z(n40859) );
  XNOR U40828 ( .A(n40874), .B(n40873), .Z(n40864) );
  XOR U40829 ( .A(n40953), .B(n40870), .Z(n40873) );
  XOR U40830 ( .A(p_input[1139]), .B(p_input[2067]), .Z(n40870) );
  XOR U40831 ( .A(p_input[1140]), .B(n29412), .Z(n40953) );
  XOR U40832 ( .A(p_input[1141]), .B(p_input[2069]), .Z(n40874) );
  XOR U40833 ( .A(n40889), .B(n40954), .Z(n40950) );
  IV U40834 ( .A(n40875), .Z(n40954) );
  XOR U40835 ( .A(p_input[1121]), .B(p_input[2049]), .Z(n40875) );
  XNOR U40836 ( .A(n40955), .B(n40897), .Z(n40889) );
  XNOR U40837 ( .A(n40885), .B(n40884), .Z(n40897) );
  XNOR U40838 ( .A(n40956), .B(n40881), .Z(n40884) );
  XNOR U40839 ( .A(p_input[1146]), .B(p_input[2074]), .Z(n40881) );
  XOR U40840 ( .A(p_input[1147]), .B(n29415), .Z(n40956) );
  XOR U40841 ( .A(p_input[1148]), .B(p_input[2076]), .Z(n40885) );
  XOR U40842 ( .A(n40895), .B(n40957), .Z(n40955) );
  IV U40843 ( .A(n40886), .Z(n40957) );
  XOR U40844 ( .A(p_input[1137]), .B(p_input[2065]), .Z(n40886) );
  XNOR U40845 ( .A(n40958), .B(n40902), .Z(n40895) );
  XNOR U40846 ( .A(p_input[1151]), .B(n29418), .Z(n40902) );
  XOR U40847 ( .A(n40892), .B(n40901), .Z(n40958) );
  XOR U40848 ( .A(n40959), .B(n40898), .Z(n40901) );
  XOR U40849 ( .A(p_input[1149]), .B(p_input[2077]), .Z(n40898) );
  XOR U40850 ( .A(p_input[1150]), .B(n29420), .Z(n40959) );
  XOR U40851 ( .A(p_input[1145]), .B(p_input[2073]), .Z(n40892) );
  XOR U40852 ( .A(n40914), .B(n40913), .Z(n40879) );
  XNOR U40853 ( .A(n40960), .B(n40921), .Z(n40913) );
  XNOR U40854 ( .A(n40909), .B(n40908), .Z(n40921) );
  XNOR U40855 ( .A(n40961), .B(n40905), .Z(n40908) );
  XNOR U40856 ( .A(p_input[1131]), .B(p_input[2059]), .Z(n40905) );
  XOR U40857 ( .A(p_input[1132]), .B(n28329), .Z(n40961) );
  XOR U40858 ( .A(p_input[1133]), .B(p_input[2061]), .Z(n40909) );
  XOR U40859 ( .A(n40919), .B(n40962), .Z(n40960) );
  IV U40860 ( .A(n40910), .Z(n40962) );
  XOR U40861 ( .A(p_input[1122]), .B(p_input[2050]), .Z(n40910) );
  XNOR U40862 ( .A(n40963), .B(n40926), .Z(n40919) );
  XNOR U40863 ( .A(p_input[1136]), .B(n28332), .Z(n40926) );
  XOR U40864 ( .A(n40916), .B(n40925), .Z(n40963) );
  XOR U40865 ( .A(n40964), .B(n40922), .Z(n40925) );
  XOR U40866 ( .A(p_input[1134]), .B(p_input[2062]), .Z(n40922) );
  XOR U40867 ( .A(p_input[1135]), .B(n28334), .Z(n40964) );
  XOR U40868 ( .A(p_input[1130]), .B(p_input[2058]), .Z(n40916) );
  XOR U40869 ( .A(n40933), .B(n40931), .Z(n40914) );
  XNOR U40870 ( .A(n40965), .B(n40938), .Z(n40931) );
  XOR U40871 ( .A(p_input[1129]), .B(p_input[2057]), .Z(n40938) );
  XOR U40872 ( .A(n40928), .B(n40937), .Z(n40965) );
  XOR U40873 ( .A(n40966), .B(n40934), .Z(n40937) );
  XOR U40874 ( .A(p_input[1127]), .B(p_input[2055]), .Z(n40934) );
  XOR U40875 ( .A(p_input[1128]), .B(n29427), .Z(n40966) );
  XOR U40876 ( .A(p_input[1123]), .B(p_input[2051]), .Z(n40928) );
  XNOR U40877 ( .A(n40943), .B(n40942), .Z(n40933) );
  XOR U40878 ( .A(n40967), .B(n40939), .Z(n40942) );
  XOR U40879 ( .A(p_input[1124]), .B(p_input[2052]), .Z(n40939) );
  XOR U40880 ( .A(p_input[1125]), .B(n29429), .Z(n40967) );
  XOR U40881 ( .A(p_input[1126]), .B(p_input[2054]), .Z(n40943) );
  XNOR U40882 ( .A(n40968), .B(n40969), .Z(n40744) );
  AND U40883 ( .A(n800), .B(n40970), .Z(n40969) );
  XNOR U40884 ( .A(n40971), .B(n40972), .Z(n800) );
  AND U40885 ( .A(n40973), .B(n40974), .Z(n40972) );
  XOR U40886 ( .A(n40758), .B(n40971), .Z(n40974) );
  XNOR U40887 ( .A(n40975), .B(n40971), .Z(n40973) );
  XOR U40888 ( .A(n40976), .B(n40977), .Z(n40971) );
  AND U40889 ( .A(n40978), .B(n40979), .Z(n40977) );
  XOR U40890 ( .A(n40773), .B(n40976), .Z(n40979) );
  XOR U40891 ( .A(n40976), .B(n40774), .Z(n40978) );
  XOR U40892 ( .A(n40980), .B(n40981), .Z(n40976) );
  AND U40893 ( .A(n40982), .B(n40983), .Z(n40981) );
  XOR U40894 ( .A(n40801), .B(n40980), .Z(n40983) );
  XOR U40895 ( .A(n40980), .B(n40802), .Z(n40982) );
  XOR U40896 ( .A(n40984), .B(n40985), .Z(n40980) );
  AND U40897 ( .A(n40986), .B(n40987), .Z(n40985) );
  XOR U40898 ( .A(n40850), .B(n40984), .Z(n40987) );
  XOR U40899 ( .A(n40984), .B(n40851), .Z(n40986) );
  XOR U40900 ( .A(n40988), .B(n40989), .Z(n40984) );
  AND U40901 ( .A(n40990), .B(n40991), .Z(n40989) );
  XOR U40902 ( .A(n40988), .B(n40947), .Z(n40991) );
  XNOR U40903 ( .A(n40992), .B(n40993), .Z(n40694) );
  AND U40904 ( .A(n804), .B(n40994), .Z(n40993) );
  XNOR U40905 ( .A(n40995), .B(n40996), .Z(n804) );
  AND U40906 ( .A(n40997), .B(n40998), .Z(n40996) );
  XOR U40907 ( .A(n40995), .B(n40704), .Z(n40998) );
  XNOR U40908 ( .A(n40995), .B(n40654), .Z(n40997) );
  XOR U40909 ( .A(n40999), .B(n41000), .Z(n40995) );
  AND U40910 ( .A(n41001), .B(n41002), .Z(n41000) );
  XNOR U40911 ( .A(n40714), .B(n40999), .Z(n41002) );
  XOR U40912 ( .A(n40999), .B(n40664), .Z(n41001) );
  XOR U40913 ( .A(n41003), .B(n41004), .Z(n40999) );
  AND U40914 ( .A(n41005), .B(n41006), .Z(n41004) );
  XNOR U40915 ( .A(n40724), .B(n41003), .Z(n41006) );
  XOR U40916 ( .A(n41003), .B(n40673), .Z(n41005) );
  XOR U40917 ( .A(n41007), .B(n41008), .Z(n41003) );
  AND U40918 ( .A(n41009), .B(n41010), .Z(n41008) );
  XOR U40919 ( .A(n41007), .B(n40681), .Z(n41009) );
  XOR U40920 ( .A(n41011), .B(n41012), .Z(n40645) );
  AND U40921 ( .A(n808), .B(n40994), .Z(n41012) );
  XNOR U40922 ( .A(n40992), .B(n41011), .Z(n40994) );
  XNOR U40923 ( .A(n41013), .B(n41014), .Z(n808) );
  AND U40924 ( .A(n41015), .B(n41016), .Z(n41014) );
  XNOR U40925 ( .A(n41017), .B(n41013), .Z(n41016) );
  IV U40926 ( .A(n40704), .Z(n41017) );
  XOR U40927 ( .A(n40975), .B(n41018), .Z(n40704) );
  AND U40928 ( .A(n811), .B(n41019), .Z(n41018) );
  XOR U40929 ( .A(n40757), .B(n40754), .Z(n41019) );
  IV U40930 ( .A(n40975), .Z(n40757) );
  XNOR U40931 ( .A(n40654), .B(n41013), .Z(n41015) );
  XOR U40932 ( .A(n41020), .B(n41021), .Z(n40654) );
  AND U40933 ( .A(n827), .B(n41022), .Z(n41021) );
  XOR U40934 ( .A(n41023), .B(n41024), .Z(n41013) );
  AND U40935 ( .A(n41025), .B(n41026), .Z(n41024) );
  XNOR U40936 ( .A(n41023), .B(n40714), .Z(n41026) );
  XOR U40937 ( .A(n40774), .B(n41027), .Z(n40714) );
  AND U40938 ( .A(n811), .B(n41028), .Z(n41027) );
  XOR U40939 ( .A(n40770), .B(n40774), .Z(n41028) );
  XNOR U40940 ( .A(n41029), .B(n41023), .Z(n41025) );
  IV U40941 ( .A(n40664), .Z(n41029) );
  XOR U40942 ( .A(n41030), .B(n41031), .Z(n40664) );
  AND U40943 ( .A(n827), .B(n41032), .Z(n41031) );
  XOR U40944 ( .A(n41033), .B(n41034), .Z(n41023) );
  AND U40945 ( .A(n41035), .B(n41036), .Z(n41034) );
  XNOR U40946 ( .A(n41033), .B(n40724), .Z(n41036) );
  XOR U40947 ( .A(n40802), .B(n41037), .Z(n40724) );
  AND U40948 ( .A(n811), .B(n41038), .Z(n41037) );
  XOR U40949 ( .A(n40798), .B(n40802), .Z(n41038) );
  XOR U40950 ( .A(n40673), .B(n41033), .Z(n41035) );
  XOR U40951 ( .A(n41039), .B(n41040), .Z(n40673) );
  AND U40952 ( .A(n827), .B(n41041), .Z(n41040) );
  XOR U40953 ( .A(n41007), .B(n41042), .Z(n41033) );
  AND U40954 ( .A(n41043), .B(n41010), .Z(n41042) );
  XNOR U40955 ( .A(n40734), .B(n41007), .Z(n41010) );
  XOR U40956 ( .A(n40851), .B(n41044), .Z(n40734) );
  AND U40957 ( .A(n811), .B(n41045), .Z(n41044) );
  XOR U40958 ( .A(n40847), .B(n40851), .Z(n41045) );
  XNOR U40959 ( .A(n41046), .B(n41007), .Z(n41043) );
  IV U40960 ( .A(n40681), .Z(n41046) );
  XOR U40961 ( .A(n41047), .B(n41048), .Z(n40681) );
  AND U40962 ( .A(n827), .B(n41049), .Z(n41048) );
  XOR U40963 ( .A(n41050), .B(n41051), .Z(n41007) );
  AND U40964 ( .A(n41052), .B(n41053), .Z(n41051) );
  XNOR U40965 ( .A(n41050), .B(n40742), .Z(n41053) );
  XOR U40966 ( .A(n40948), .B(n41054), .Z(n40742) );
  AND U40967 ( .A(n811), .B(n41055), .Z(n41054) );
  XOR U40968 ( .A(n40944), .B(n40948), .Z(n41055) );
  XNOR U40969 ( .A(n41056), .B(n41050), .Z(n41052) );
  IV U40970 ( .A(n40691), .Z(n41056) );
  XOR U40971 ( .A(n41057), .B(n41058), .Z(n40691) );
  AND U40972 ( .A(n827), .B(n41059), .Z(n41058) );
  AND U40973 ( .A(n41011), .B(n40992), .Z(n41050) );
  XNOR U40974 ( .A(n41060), .B(n41061), .Z(n40992) );
  AND U40975 ( .A(n811), .B(n40970), .Z(n41061) );
  XNOR U40976 ( .A(n40968), .B(n41060), .Z(n40970) );
  XNOR U40977 ( .A(n41062), .B(n41063), .Z(n811) );
  AND U40978 ( .A(n41064), .B(n41065), .Z(n41063) );
  XNOR U40979 ( .A(n41062), .B(n40754), .Z(n41065) );
  IV U40980 ( .A(n40758), .Z(n40754) );
  XOR U40981 ( .A(n41066), .B(n41067), .Z(n40758) );
  AND U40982 ( .A(n815), .B(n41068), .Z(n41067) );
  XOR U40983 ( .A(n41069), .B(n41066), .Z(n41068) );
  XNOR U40984 ( .A(n41062), .B(n40975), .Z(n41064) );
  XOR U40985 ( .A(n41070), .B(n41071), .Z(n40975) );
  AND U40986 ( .A(n823), .B(n41022), .Z(n41071) );
  XOR U40987 ( .A(n41020), .B(n41070), .Z(n41022) );
  XOR U40988 ( .A(n41072), .B(n41073), .Z(n41062) );
  AND U40989 ( .A(n41074), .B(n41075), .Z(n41073) );
  XNOR U40990 ( .A(n41072), .B(n40770), .Z(n41075) );
  IV U40991 ( .A(n40773), .Z(n40770) );
  XOR U40992 ( .A(n41076), .B(n41077), .Z(n40773) );
  AND U40993 ( .A(n815), .B(n41078), .Z(n41077) );
  XOR U40994 ( .A(n41079), .B(n41076), .Z(n41078) );
  XOR U40995 ( .A(n40774), .B(n41072), .Z(n41074) );
  XOR U40996 ( .A(n41080), .B(n41081), .Z(n40774) );
  AND U40997 ( .A(n823), .B(n41032), .Z(n41081) );
  XOR U40998 ( .A(n41080), .B(n41030), .Z(n41032) );
  XOR U40999 ( .A(n41082), .B(n41083), .Z(n41072) );
  AND U41000 ( .A(n41084), .B(n41085), .Z(n41083) );
  XNOR U41001 ( .A(n41082), .B(n40798), .Z(n41085) );
  IV U41002 ( .A(n40801), .Z(n40798) );
  XOR U41003 ( .A(n41086), .B(n41087), .Z(n40801) );
  AND U41004 ( .A(n815), .B(n41088), .Z(n41087) );
  XNOR U41005 ( .A(n41089), .B(n41086), .Z(n41088) );
  XOR U41006 ( .A(n40802), .B(n41082), .Z(n41084) );
  XOR U41007 ( .A(n41090), .B(n41091), .Z(n40802) );
  AND U41008 ( .A(n823), .B(n41041), .Z(n41091) );
  XOR U41009 ( .A(n41090), .B(n41039), .Z(n41041) );
  XOR U41010 ( .A(n41092), .B(n41093), .Z(n41082) );
  AND U41011 ( .A(n41094), .B(n41095), .Z(n41093) );
  XNOR U41012 ( .A(n41092), .B(n40847), .Z(n41095) );
  IV U41013 ( .A(n40850), .Z(n40847) );
  XOR U41014 ( .A(n41096), .B(n41097), .Z(n40850) );
  AND U41015 ( .A(n815), .B(n41098), .Z(n41097) );
  XOR U41016 ( .A(n41099), .B(n41096), .Z(n41098) );
  XOR U41017 ( .A(n40851), .B(n41092), .Z(n41094) );
  XOR U41018 ( .A(n41100), .B(n41101), .Z(n40851) );
  AND U41019 ( .A(n823), .B(n41049), .Z(n41101) );
  XOR U41020 ( .A(n41100), .B(n41047), .Z(n41049) );
  XOR U41021 ( .A(n40988), .B(n41102), .Z(n41092) );
  AND U41022 ( .A(n40990), .B(n41103), .Z(n41102) );
  XNOR U41023 ( .A(n40988), .B(n40944), .Z(n41103) );
  IV U41024 ( .A(n40947), .Z(n40944) );
  XOR U41025 ( .A(n41104), .B(n41105), .Z(n40947) );
  AND U41026 ( .A(n815), .B(n41106), .Z(n41105) );
  XNOR U41027 ( .A(n41107), .B(n41104), .Z(n41106) );
  XOR U41028 ( .A(n40948), .B(n40988), .Z(n40990) );
  XOR U41029 ( .A(n41108), .B(n41109), .Z(n40948) );
  AND U41030 ( .A(n823), .B(n41059), .Z(n41109) );
  XOR U41031 ( .A(n41108), .B(n41057), .Z(n41059) );
  AND U41032 ( .A(n41060), .B(n40968), .Z(n40988) );
  XNOR U41033 ( .A(n41110), .B(n41111), .Z(n40968) );
  AND U41034 ( .A(n815), .B(n41112), .Z(n41111) );
  XNOR U41035 ( .A(n41113), .B(n41110), .Z(n41112) );
  XNOR U41036 ( .A(n41114), .B(n41115), .Z(n815) );
  AND U41037 ( .A(n41116), .B(n41117), .Z(n41115) );
  XOR U41038 ( .A(n41069), .B(n41114), .Z(n41117) );
  AND U41039 ( .A(n41118), .B(n41119), .Z(n41069) );
  XNOR U41040 ( .A(n41066), .B(n41114), .Z(n41116) );
  XNOR U41041 ( .A(n41120), .B(n41121), .Z(n41066) );
  AND U41042 ( .A(n819), .B(n41122), .Z(n41121) );
  XNOR U41043 ( .A(n41123), .B(n41124), .Z(n41122) );
  XOR U41044 ( .A(n41125), .B(n41126), .Z(n41114) );
  AND U41045 ( .A(n41127), .B(n41128), .Z(n41126) );
  XNOR U41046 ( .A(n41125), .B(n41118), .Z(n41128) );
  IV U41047 ( .A(n41079), .Z(n41118) );
  XOR U41048 ( .A(n41129), .B(n41130), .Z(n41079) );
  XOR U41049 ( .A(n41131), .B(n41119), .Z(n41130) );
  AND U41050 ( .A(n41089), .B(n41132), .Z(n41119) );
  AND U41051 ( .A(n41133), .B(n41134), .Z(n41131) );
  XOR U41052 ( .A(n41135), .B(n41129), .Z(n41133) );
  XNOR U41053 ( .A(n41076), .B(n41125), .Z(n41127) );
  XNOR U41054 ( .A(n41136), .B(n41137), .Z(n41076) );
  AND U41055 ( .A(n819), .B(n41138), .Z(n41137) );
  XNOR U41056 ( .A(n41139), .B(n41140), .Z(n41138) );
  XOR U41057 ( .A(n41141), .B(n41142), .Z(n41125) );
  AND U41058 ( .A(n41143), .B(n41144), .Z(n41142) );
  XNOR U41059 ( .A(n41141), .B(n41089), .Z(n41144) );
  XOR U41060 ( .A(n41145), .B(n41134), .Z(n41089) );
  XNOR U41061 ( .A(n41146), .B(n41129), .Z(n41134) );
  XOR U41062 ( .A(n41147), .B(n41148), .Z(n41129) );
  AND U41063 ( .A(n41149), .B(n41150), .Z(n41148) );
  XOR U41064 ( .A(n41151), .B(n41147), .Z(n41149) );
  XNOR U41065 ( .A(n41152), .B(n41153), .Z(n41146) );
  AND U41066 ( .A(n41154), .B(n41155), .Z(n41153) );
  XOR U41067 ( .A(n41152), .B(n41156), .Z(n41154) );
  XNOR U41068 ( .A(n41135), .B(n41132), .Z(n41145) );
  AND U41069 ( .A(n41157), .B(n41158), .Z(n41132) );
  XOR U41070 ( .A(n41159), .B(n41160), .Z(n41135) );
  AND U41071 ( .A(n41161), .B(n41162), .Z(n41160) );
  XOR U41072 ( .A(n41159), .B(n41163), .Z(n41161) );
  XNOR U41073 ( .A(n41086), .B(n41141), .Z(n41143) );
  XNOR U41074 ( .A(n41164), .B(n41165), .Z(n41086) );
  AND U41075 ( .A(n819), .B(n41166), .Z(n41165) );
  XNOR U41076 ( .A(n41167), .B(n41168), .Z(n41166) );
  XOR U41077 ( .A(n41169), .B(n41170), .Z(n41141) );
  AND U41078 ( .A(n41171), .B(n41172), .Z(n41170) );
  XNOR U41079 ( .A(n41169), .B(n41157), .Z(n41172) );
  IV U41080 ( .A(n41099), .Z(n41157) );
  XNOR U41081 ( .A(n41173), .B(n41150), .Z(n41099) );
  XNOR U41082 ( .A(n41174), .B(n41156), .Z(n41150) );
  XOR U41083 ( .A(n41175), .B(n41176), .Z(n41156) );
  AND U41084 ( .A(n41177), .B(n41178), .Z(n41176) );
  XOR U41085 ( .A(n41175), .B(n41179), .Z(n41177) );
  XNOR U41086 ( .A(n41155), .B(n41147), .Z(n41174) );
  XOR U41087 ( .A(n41180), .B(n41181), .Z(n41147) );
  AND U41088 ( .A(n41182), .B(n41183), .Z(n41181) );
  XNOR U41089 ( .A(n41184), .B(n41180), .Z(n41182) );
  XNOR U41090 ( .A(n41185), .B(n41152), .Z(n41155) );
  XOR U41091 ( .A(n41186), .B(n41187), .Z(n41152) );
  AND U41092 ( .A(n41188), .B(n41189), .Z(n41187) );
  XOR U41093 ( .A(n41186), .B(n41190), .Z(n41188) );
  XNOR U41094 ( .A(n41191), .B(n41192), .Z(n41185) );
  AND U41095 ( .A(n41193), .B(n41194), .Z(n41192) );
  XNOR U41096 ( .A(n41191), .B(n41195), .Z(n41193) );
  XNOR U41097 ( .A(n41151), .B(n41158), .Z(n41173) );
  AND U41098 ( .A(n41107), .B(n41196), .Z(n41158) );
  XOR U41099 ( .A(n41163), .B(n41162), .Z(n41151) );
  XNOR U41100 ( .A(n41197), .B(n41159), .Z(n41162) );
  XOR U41101 ( .A(n41198), .B(n41199), .Z(n41159) );
  AND U41102 ( .A(n41200), .B(n41201), .Z(n41199) );
  XOR U41103 ( .A(n41198), .B(n41202), .Z(n41200) );
  XNOR U41104 ( .A(n41203), .B(n41204), .Z(n41197) );
  AND U41105 ( .A(n41205), .B(n41206), .Z(n41204) );
  XOR U41106 ( .A(n41203), .B(n41207), .Z(n41205) );
  XOR U41107 ( .A(n41208), .B(n41209), .Z(n41163) );
  AND U41108 ( .A(n41210), .B(n41211), .Z(n41209) );
  XOR U41109 ( .A(n41208), .B(n41212), .Z(n41210) );
  XNOR U41110 ( .A(n41096), .B(n41169), .Z(n41171) );
  XNOR U41111 ( .A(n41213), .B(n41214), .Z(n41096) );
  AND U41112 ( .A(n819), .B(n41215), .Z(n41214) );
  XNOR U41113 ( .A(n41216), .B(n41217), .Z(n41215) );
  XOR U41114 ( .A(n41218), .B(n41219), .Z(n41169) );
  AND U41115 ( .A(n41220), .B(n41221), .Z(n41219) );
  XNOR U41116 ( .A(n41218), .B(n41107), .Z(n41221) );
  XOR U41117 ( .A(n41222), .B(n41183), .Z(n41107) );
  XNOR U41118 ( .A(n41223), .B(n41190), .Z(n41183) );
  XOR U41119 ( .A(n41179), .B(n41178), .Z(n41190) );
  XNOR U41120 ( .A(n41224), .B(n41175), .Z(n41178) );
  XOR U41121 ( .A(n41225), .B(n41226), .Z(n41175) );
  AND U41122 ( .A(n41227), .B(n41228), .Z(n41226) );
  XNOR U41123 ( .A(n41229), .B(n41230), .Z(n41227) );
  IV U41124 ( .A(n41225), .Z(n41229) );
  XNOR U41125 ( .A(n41231), .B(n41232), .Z(n41224) );
  NOR U41126 ( .A(n41233), .B(n41234), .Z(n41232) );
  XNOR U41127 ( .A(n41231), .B(n41235), .Z(n41233) );
  XOR U41128 ( .A(n41236), .B(n41237), .Z(n41179) );
  NOR U41129 ( .A(n41238), .B(n41239), .Z(n41237) );
  XNOR U41130 ( .A(n41236), .B(n41240), .Z(n41238) );
  XNOR U41131 ( .A(n41189), .B(n41180), .Z(n41223) );
  XOR U41132 ( .A(n41241), .B(n41242), .Z(n41180) );
  AND U41133 ( .A(n41243), .B(n41244), .Z(n41242) );
  XOR U41134 ( .A(n41241), .B(n41245), .Z(n41243) );
  XOR U41135 ( .A(n41246), .B(n41195), .Z(n41189) );
  XOR U41136 ( .A(n41247), .B(n41248), .Z(n41195) );
  NOR U41137 ( .A(n41249), .B(n41250), .Z(n41248) );
  XOR U41138 ( .A(n41247), .B(n41251), .Z(n41249) );
  XNOR U41139 ( .A(n41194), .B(n41186), .Z(n41246) );
  XOR U41140 ( .A(n41252), .B(n41253), .Z(n41186) );
  AND U41141 ( .A(n41254), .B(n41255), .Z(n41253) );
  XOR U41142 ( .A(n41252), .B(n41256), .Z(n41254) );
  XNOR U41143 ( .A(n41257), .B(n41191), .Z(n41194) );
  XOR U41144 ( .A(n41258), .B(n41259), .Z(n41191) );
  AND U41145 ( .A(n41260), .B(n41261), .Z(n41259) );
  XNOR U41146 ( .A(n41262), .B(n41263), .Z(n41260) );
  IV U41147 ( .A(n41258), .Z(n41262) );
  XNOR U41148 ( .A(n41264), .B(n41265), .Z(n41257) );
  NOR U41149 ( .A(n41266), .B(n41267), .Z(n41265) );
  XNOR U41150 ( .A(n41264), .B(n41268), .Z(n41266) );
  XOR U41151 ( .A(n41184), .B(n41196), .Z(n41222) );
  NOR U41152 ( .A(n41113), .B(n41269), .Z(n41196) );
  XNOR U41153 ( .A(n41202), .B(n41201), .Z(n41184) );
  XNOR U41154 ( .A(n41270), .B(n41207), .Z(n41201) );
  XNOR U41155 ( .A(n41271), .B(n41272), .Z(n41207) );
  NOR U41156 ( .A(n41273), .B(n41274), .Z(n41272) );
  XOR U41157 ( .A(n41271), .B(n41275), .Z(n41273) );
  XNOR U41158 ( .A(n41206), .B(n41198), .Z(n41270) );
  XOR U41159 ( .A(n41276), .B(n41277), .Z(n41198) );
  AND U41160 ( .A(n41278), .B(n41279), .Z(n41277) );
  XOR U41161 ( .A(n41276), .B(n41280), .Z(n41278) );
  XNOR U41162 ( .A(n41281), .B(n41203), .Z(n41206) );
  XOR U41163 ( .A(n41282), .B(n41283), .Z(n41203) );
  AND U41164 ( .A(n41284), .B(n41285), .Z(n41283) );
  XNOR U41165 ( .A(n41286), .B(n41287), .Z(n41284) );
  IV U41166 ( .A(n41282), .Z(n41286) );
  XNOR U41167 ( .A(n41288), .B(n41289), .Z(n41281) );
  NOR U41168 ( .A(n41290), .B(n41291), .Z(n41289) );
  XNOR U41169 ( .A(n41288), .B(n41292), .Z(n41290) );
  XOR U41170 ( .A(n41212), .B(n41211), .Z(n41202) );
  XNOR U41171 ( .A(n41293), .B(n41208), .Z(n41211) );
  XOR U41172 ( .A(n41294), .B(n41295), .Z(n41208) );
  AND U41173 ( .A(n41296), .B(n41297), .Z(n41295) );
  XNOR U41174 ( .A(n41298), .B(n41299), .Z(n41296) );
  IV U41175 ( .A(n41294), .Z(n41298) );
  XNOR U41176 ( .A(n41300), .B(n41301), .Z(n41293) );
  NOR U41177 ( .A(n41302), .B(n41303), .Z(n41301) );
  XNOR U41178 ( .A(n41300), .B(n41304), .Z(n41302) );
  XOR U41179 ( .A(n41305), .B(n41306), .Z(n41212) );
  NOR U41180 ( .A(n41307), .B(n41308), .Z(n41306) );
  XNOR U41181 ( .A(n41305), .B(n41309), .Z(n41307) );
  XNOR U41182 ( .A(n41104), .B(n41218), .Z(n41220) );
  XNOR U41183 ( .A(n41310), .B(n41311), .Z(n41104) );
  AND U41184 ( .A(n819), .B(n41312), .Z(n41311) );
  XNOR U41185 ( .A(n41313), .B(n41314), .Z(n41312) );
  AND U41186 ( .A(n41110), .B(n41113), .Z(n41218) );
  XOR U41187 ( .A(n41315), .B(n41269), .Z(n41113) );
  XNOR U41188 ( .A(p_input[1152]), .B(p_input[2048]), .Z(n41269) );
  XNOR U41189 ( .A(n41245), .B(n41244), .Z(n41315) );
  XNOR U41190 ( .A(n41316), .B(n41256), .Z(n41244) );
  XOR U41191 ( .A(n41230), .B(n41228), .Z(n41256) );
  XNOR U41192 ( .A(n41317), .B(n41235), .Z(n41228) );
  XOR U41193 ( .A(p_input[1176]), .B(p_input[2072]), .Z(n41235) );
  XOR U41194 ( .A(n41225), .B(n41234), .Z(n41317) );
  XOR U41195 ( .A(n41318), .B(n41231), .Z(n41234) );
  XOR U41196 ( .A(p_input[1174]), .B(p_input[2070]), .Z(n41231) );
  XOR U41197 ( .A(p_input[1175]), .B(n29410), .Z(n41318) );
  XOR U41198 ( .A(p_input[1170]), .B(p_input[2066]), .Z(n41225) );
  XNOR U41199 ( .A(n41240), .B(n41239), .Z(n41230) );
  XOR U41200 ( .A(n41319), .B(n41236), .Z(n41239) );
  XOR U41201 ( .A(p_input[1171]), .B(p_input[2067]), .Z(n41236) );
  XOR U41202 ( .A(p_input[1172]), .B(n29412), .Z(n41319) );
  XOR U41203 ( .A(p_input[1173]), .B(p_input[2069]), .Z(n41240) );
  XOR U41204 ( .A(n41255), .B(n41320), .Z(n41316) );
  IV U41205 ( .A(n41241), .Z(n41320) );
  XOR U41206 ( .A(p_input[1153]), .B(p_input[2049]), .Z(n41241) );
  XNOR U41207 ( .A(n41321), .B(n41263), .Z(n41255) );
  XNOR U41208 ( .A(n41251), .B(n41250), .Z(n41263) );
  XNOR U41209 ( .A(n41322), .B(n41247), .Z(n41250) );
  XNOR U41210 ( .A(p_input[1178]), .B(p_input[2074]), .Z(n41247) );
  XOR U41211 ( .A(p_input[1179]), .B(n29415), .Z(n41322) );
  XOR U41212 ( .A(p_input[1180]), .B(p_input[2076]), .Z(n41251) );
  XOR U41213 ( .A(n41261), .B(n41323), .Z(n41321) );
  IV U41214 ( .A(n41252), .Z(n41323) );
  XOR U41215 ( .A(p_input[1169]), .B(p_input[2065]), .Z(n41252) );
  XNOR U41216 ( .A(n41324), .B(n41268), .Z(n41261) );
  XNOR U41217 ( .A(p_input[1183]), .B(n29418), .Z(n41268) );
  XOR U41218 ( .A(n41258), .B(n41267), .Z(n41324) );
  XOR U41219 ( .A(n41325), .B(n41264), .Z(n41267) );
  XOR U41220 ( .A(p_input[1181]), .B(p_input[2077]), .Z(n41264) );
  XOR U41221 ( .A(p_input[1182]), .B(n29420), .Z(n41325) );
  XOR U41222 ( .A(p_input[1177]), .B(p_input[2073]), .Z(n41258) );
  XOR U41223 ( .A(n41280), .B(n41279), .Z(n41245) );
  XNOR U41224 ( .A(n41326), .B(n41287), .Z(n41279) );
  XNOR U41225 ( .A(n41275), .B(n41274), .Z(n41287) );
  XNOR U41226 ( .A(n41327), .B(n41271), .Z(n41274) );
  XNOR U41227 ( .A(p_input[1163]), .B(p_input[2059]), .Z(n41271) );
  XOR U41228 ( .A(p_input[1164]), .B(n28329), .Z(n41327) );
  XOR U41229 ( .A(p_input[1165]), .B(p_input[2061]), .Z(n41275) );
  XOR U41230 ( .A(n41285), .B(n41328), .Z(n41326) );
  IV U41231 ( .A(n41276), .Z(n41328) );
  XOR U41232 ( .A(p_input[1154]), .B(p_input[2050]), .Z(n41276) );
  XNOR U41233 ( .A(n41329), .B(n41292), .Z(n41285) );
  XNOR U41234 ( .A(p_input[1168]), .B(n28332), .Z(n41292) );
  XOR U41235 ( .A(n41282), .B(n41291), .Z(n41329) );
  XOR U41236 ( .A(n41330), .B(n41288), .Z(n41291) );
  XOR U41237 ( .A(p_input[1166]), .B(p_input[2062]), .Z(n41288) );
  XOR U41238 ( .A(p_input[1167]), .B(n28334), .Z(n41330) );
  XOR U41239 ( .A(p_input[1162]), .B(p_input[2058]), .Z(n41282) );
  XOR U41240 ( .A(n41299), .B(n41297), .Z(n41280) );
  XNOR U41241 ( .A(n41331), .B(n41304), .Z(n41297) );
  XOR U41242 ( .A(p_input[1161]), .B(p_input[2057]), .Z(n41304) );
  XOR U41243 ( .A(n41294), .B(n41303), .Z(n41331) );
  XOR U41244 ( .A(n41332), .B(n41300), .Z(n41303) );
  XOR U41245 ( .A(p_input[1159]), .B(p_input[2055]), .Z(n41300) );
  XOR U41246 ( .A(p_input[1160]), .B(n29427), .Z(n41332) );
  XOR U41247 ( .A(p_input[1155]), .B(p_input[2051]), .Z(n41294) );
  XNOR U41248 ( .A(n41309), .B(n41308), .Z(n41299) );
  XOR U41249 ( .A(n41333), .B(n41305), .Z(n41308) );
  XOR U41250 ( .A(p_input[1156]), .B(p_input[2052]), .Z(n41305) );
  XOR U41251 ( .A(p_input[1157]), .B(n29429), .Z(n41333) );
  XOR U41252 ( .A(p_input[1158]), .B(p_input[2054]), .Z(n41309) );
  XNOR U41253 ( .A(n41334), .B(n41335), .Z(n41110) );
  AND U41254 ( .A(n819), .B(n41336), .Z(n41335) );
  XNOR U41255 ( .A(n41337), .B(n41338), .Z(n819) );
  AND U41256 ( .A(n41339), .B(n41340), .Z(n41338) );
  XOR U41257 ( .A(n41124), .B(n41337), .Z(n41340) );
  XNOR U41258 ( .A(n41341), .B(n41337), .Z(n41339) );
  XOR U41259 ( .A(n41342), .B(n41343), .Z(n41337) );
  AND U41260 ( .A(n41344), .B(n41345), .Z(n41343) );
  XOR U41261 ( .A(n41139), .B(n41342), .Z(n41345) );
  XOR U41262 ( .A(n41342), .B(n41140), .Z(n41344) );
  XOR U41263 ( .A(n41346), .B(n41347), .Z(n41342) );
  AND U41264 ( .A(n41348), .B(n41349), .Z(n41347) );
  XOR U41265 ( .A(n41167), .B(n41346), .Z(n41349) );
  XOR U41266 ( .A(n41346), .B(n41168), .Z(n41348) );
  XOR U41267 ( .A(n41350), .B(n41351), .Z(n41346) );
  AND U41268 ( .A(n41352), .B(n41353), .Z(n41351) );
  XOR U41269 ( .A(n41216), .B(n41350), .Z(n41353) );
  XOR U41270 ( .A(n41350), .B(n41217), .Z(n41352) );
  XOR U41271 ( .A(n41354), .B(n41355), .Z(n41350) );
  AND U41272 ( .A(n41356), .B(n41357), .Z(n41355) );
  XOR U41273 ( .A(n41354), .B(n41313), .Z(n41357) );
  XNOR U41274 ( .A(n41358), .B(n41359), .Z(n41060) );
  AND U41275 ( .A(n823), .B(n41360), .Z(n41359) );
  XNOR U41276 ( .A(n41361), .B(n41362), .Z(n823) );
  AND U41277 ( .A(n41363), .B(n41364), .Z(n41362) );
  XOR U41278 ( .A(n41361), .B(n41070), .Z(n41364) );
  XNOR U41279 ( .A(n41361), .B(n41020), .Z(n41363) );
  XOR U41280 ( .A(n41365), .B(n41366), .Z(n41361) );
  AND U41281 ( .A(n41367), .B(n41368), .Z(n41366) );
  XNOR U41282 ( .A(n41080), .B(n41365), .Z(n41368) );
  XOR U41283 ( .A(n41365), .B(n41030), .Z(n41367) );
  XOR U41284 ( .A(n41369), .B(n41370), .Z(n41365) );
  AND U41285 ( .A(n41371), .B(n41372), .Z(n41370) );
  XNOR U41286 ( .A(n41090), .B(n41369), .Z(n41372) );
  XOR U41287 ( .A(n41369), .B(n41039), .Z(n41371) );
  XOR U41288 ( .A(n41373), .B(n41374), .Z(n41369) );
  AND U41289 ( .A(n41375), .B(n41376), .Z(n41374) );
  XOR U41290 ( .A(n41373), .B(n41047), .Z(n41375) );
  XOR U41291 ( .A(n41377), .B(n41378), .Z(n41011) );
  AND U41292 ( .A(n827), .B(n41360), .Z(n41378) );
  XNOR U41293 ( .A(n41358), .B(n41377), .Z(n41360) );
  XNOR U41294 ( .A(n41379), .B(n41380), .Z(n827) );
  AND U41295 ( .A(n41381), .B(n41382), .Z(n41380) );
  XNOR U41296 ( .A(n41383), .B(n41379), .Z(n41382) );
  IV U41297 ( .A(n41070), .Z(n41383) );
  XOR U41298 ( .A(n41341), .B(n41384), .Z(n41070) );
  AND U41299 ( .A(n830), .B(n41385), .Z(n41384) );
  XOR U41300 ( .A(n41123), .B(n41120), .Z(n41385) );
  IV U41301 ( .A(n41341), .Z(n41123) );
  XNOR U41302 ( .A(n41020), .B(n41379), .Z(n41381) );
  XOR U41303 ( .A(n41386), .B(n41387), .Z(n41020) );
  AND U41304 ( .A(n846), .B(n41388), .Z(n41387) );
  XOR U41305 ( .A(n41389), .B(n41390), .Z(n41379) );
  AND U41306 ( .A(n41391), .B(n41392), .Z(n41390) );
  XNOR U41307 ( .A(n41389), .B(n41080), .Z(n41392) );
  XOR U41308 ( .A(n41140), .B(n41393), .Z(n41080) );
  AND U41309 ( .A(n830), .B(n41394), .Z(n41393) );
  XOR U41310 ( .A(n41136), .B(n41140), .Z(n41394) );
  XNOR U41311 ( .A(n41395), .B(n41389), .Z(n41391) );
  IV U41312 ( .A(n41030), .Z(n41395) );
  XOR U41313 ( .A(n41396), .B(n41397), .Z(n41030) );
  AND U41314 ( .A(n846), .B(n41398), .Z(n41397) );
  XOR U41315 ( .A(n41399), .B(n41400), .Z(n41389) );
  AND U41316 ( .A(n41401), .B(n41402), .Z(n41400) );
  XNOR U41317 ( .A(n41399), .B(n41090), .Z(n41402) );
  XOR U41318 ( .A(n41168), .B(n41403), .Z(n41090) );
  AND U41319 ( .A(n830), .B(n41404), .Z(n41403) );
  XOR U41320 ( .A(n41164), .B(n41168), .Z(n41404) );
  XOR U41321 ( .A(n41039), .B(n41399), .Z(n41401) );
  XOR U41322 ( .A(n41405), .B(n41406), .Z(n41039) );
  AND U41323 ( .A(n846), .B(n41407), .Z(n41406) );
  XOR U41324 ( .A(n41373), .B(n41408), .Z(n41399) );
  AND U41325 ( .A(n41409), .B(n41376), .Z(n41408) );
  XNOR U41326 ( .A(n41100), .B(n41373), .Z(n41376) );
  XOR U41327 ( .A(n41217), .B(n41410), .Z(n41100) );
  AND U41328 ( .A(n830), .B(n41411), .Z(n41410) );
  XOR U41329 ( .A(n41213), .B(n41217), .Z(n41411) );
  XNOR U41330 ( .A(n41412), .B(n41373), .Z(n41409) );
  IV U41331 ( .A(n41047), .Z(n41412) );
  XOR U41332 ( .A(n41413), .B(n41414), .Z(n41047) );
  AND U41333 ( .A(n846), .B(n41415), .Z(n41414) );
  XOR U41334 ( .A(n41416), .B(n41417), .Z(n41373) );
  AND U41335 ( .A(n41418), .B(n41419), .Z(n41417) );
  XNOR U41336 ( .A(n41416), .B(n41108), .Z(n41419) );
  XOR U41337 ( .A(n41314), .B(n41420), .Z(n41108) );
  AND U41338 ( .A(n830), .B(n41421), .Z(n41420) );
  XOR U41339 ( .A(n41310), .B(n41314), .Z(n41421) );
  XNOR U41340 ( .A(n41422), .B(n41416), .Z(n41418) );
  IV U41341 ( .A(n41057), .Z(n41422) );
  XOR U41342 ( .A(n41423), .B(n41424), .Z(n41057) );
  AND U41343 ( .A(n846), .B(n41425), .Z(n41424) );
  AND U41344 ( .A(n41377), .B(n41358), .Z(n41416) );
  XNOR U41345 ( .A(n41426), .B(n41427), .Z(n41358) );
  AND U41346 ( .A(n830), .B(n41336), .Z(n41427) );
  XNOR U41347 ( .A(n41334), .B(n41426), .Z(n41336) );
  XNOR U41348 ( .A(n41428), .B(n41429), .Z(n830) );
  AND U41349 ( .A(n41430), .B(n41431), .Z(n41429) );
  XNOR U41350 ( .A(n41428), .B(n41120), .Z(n41431) );
  IV U41351 ( .A(n41124), .Z(n41120) );
  XOR U41352 ( .A(n41432), .B(n41433), .Z(n41124) );
  AND U41353 ( .A(n834), .B(n41434), .Z(n41433) );
  XOR U41354 ( .A(n41435), .B(n41432), .Z(n41434) );
  XNOR U41355 ( .A(n41428), .B(n41341), .Z(n41430) );
  XOR U41356 ( .A(n41436), .B(n41437), .Z(n41341) );
  AND U41357 ( .A(n842), .B(n41388), .Z(n41437) );
  XOR U41358 ( .A(n41386), .B(n41436), .Z(n41388) );
  XOR U41359 ( .A(n41438), .B(n41439), .Z(n41428) );
  AND U41360 ( .A(n41440), .B(n41441), .Z(n41439) );
  XNOR U41361 ( .A(n41438), .B(n41136), .Z(n41441) );
  IV U41362 ( .A(n41139), .Z(n41136) );
  XOR U41363 ( .A(n41442), .B(n41443), .Z(n41139) );
  AND U41364 ( .A(n834), .B(n41444), .Z(n41443) );
  XOR U41365 ( .A(n41445), .B(n41442), .Z(n41444) );
  XOR U41366 ( .A(n41140), .B(n41438), .Z(n41440) );
  XOR U41367 ( .A(n41446), .B(n41447), .Z(n41140) );
  AND U41368 ( .A(n842), .B(n41398), .Z(n41447) );
  XOR U41369 ( .A(n41446), .B(n41396), .Z(n41398) );
  XOR U41370 ( .A(n41448), .B(n41449), .Z(n41438) );
  AND U41371 ( .A(n41450), .B(n41451), .Z(n41449) );
  XNOR U41372 ( .A(n41448), .B(n41164), .Z(n41451) );
  IV U41373 ( .A(n41167), .Z(n41164) );
  XOR U41374 ( .A(n41452), .B(n41453), .Z(n41167) );
  AND U41375 ( .A(n834), .B(n41454), .Z(n41453) );
  XNOR U41376 ( .A(n41455), .B(n41452), .Z(n41454) );
  XOR U41377 ( .A(n41168), .B(n41448), .Z(n41450) );
  XOR U41378 ( .A(n41456), .B(n41457), .Z(n41168) );
  AND U41379 ( .A(n842), .B(n41407), .Z(n41457) );
  XOR U41380 ( .A(n41456), .B(n41405), .Z(n41407) );
  XOR U41381 ( .A(n41458), .B(n41459), .Z(n41448) );
  AND U41382 ( .A(n41460), .B(n41461), .Z(n41459) );
  XNOR U41383 ( .A(n41458), .B(n41213), .Z(n41461) );
  IV U41384 ( .A(n41216), .Z(n41213) );
  XOR U41385 ( .A(n41462), .B(n41463), .Z(n41216) );
  AND U41386 ( .A(n834), .B(n41464), .Z(n41463) );
  XOR U41387 ( .A(n41465), .B(n41462), .Z(n41464) );
  XOR U41388 ( .A(n41217), .B(n41458), .Z(n41460) );
  XOR U41389 ( .A(n41466), .B(n41467), .Z(n41217) );
  AND U41390 ( .A(n842), .B(n41415), .Z(n41467) );
  XOR U41391 ( .A(n41466), .B(n41413), .Z(n41415) );
  XOR U41392 ( .A(n41354), .B(n41468), .Z(n41458) );
  AND U41393 ( .A(n41356), .B(n41469), .Z(n41468) );
  XNOR U41394 ( .A(n41354), .B(n41310), .Z(n41469) );
  IV U41395 ( .A(n41313), .Z(n41310) );
  XOR U41396 ( .A(n41470), .B(n41471), .Z(n41313) );
  AND U41397 ( .A(n834), .B(n41472), .Z(n41471) );
  XNOR U41398 ( .A(n41473), .B(n41470), .Z(n41472) );
  XOR U41399 ( .A(n41314), .B(n41354), .Z(n41356) );
  XOR U41400 ( .A(n41474), .B(n41475), .Z(n41314) );
  AND U41401 ( .A(n842), .B(n41425), .Z(n41475) );
  XOR U41402 ( .A(n41474), .B(n41423), .Z(n41425) );
  AND U41403 ( .A(n41426), .B(n41334), .Z(n41354) );
  XNOR U41404 ( .A(n41476), .B(n41477), .Z(n41334) );
  AND U41405 ( .A(n834), .B(n41478), .Z(n41477) );
  XNOR U41406 ( .A(n41479), .B(n41476), .Z(n41478) );
  XNOR U41407 ( .A(n41480), .B(n41481), .Z(n834) );
  AND U41408 ( .A(n41482), .B(n41483), .Z(n41481) );
  XOR U41409 ( .A(n41435), .B(n41480), .Z(n41483) );
  AND U41410 ( .A(n41484), .B(n41485), .Z(n41435) );
  XNOR U41411 ( .A(n41432), .B(n41480), .Z(n41482) );
  XNOR U41412 ( .A(n41486), .B(n41487), .Z(n41432) );
  AND U41413 ( .A(n838), .B(n41488), .Z(n41487) );
  XNOR U41414 ( .A(n41489), .B(n41490), .Z(n41488) );
  XOR U41415 ( .A(n41491), .B(n41492), .Z(n41480) );
  AND U41416 ( .A(n41493), .B(n41494), .Z(n41492) );
  XNOR U41417 ( .A(n41491), .B(n41484), .Z(n41494) );
  IV U41418 ( .A(n41445), .Z(n41484) );
  XOR U41419 ( .A(n41495), .B(n41496), .Z(n41445) );
  XOR U41420 ( .A(n41497), .B(n41485), .Z(n41496) );
  AND U41421 ( .A(n41455), .B(n41498), .Z(n41485) );
  AND U41422 ( .A(n41499), .B(n41500), .Z(n41497) );
  XOR U41423 ( .A(n41501), .B(n41495), .Z(n41499) );
  XNOR U41424 ( .A(n41442), .B(n41491), .Z(n41493) );
  XNOR U41425 ( .A(n41502), .B(n41503), .Z(n41442) );
  AND U41426 ( .A(n838), .B(n41504), .Z(n41503) );
  XNOR U41427 ( .A(n41505), .B(n41506), .Z(n41504) );
  XOR U41428 ( .A(n41507), .B(n41508), .Z(n41491) );
  AND U41429 ( .A(n41509), .B(n41510), .Z(n41508) );
  XNOR U41430 ( .A(n41507), .B(n41455), .Z(n41510) );
  XOR U41431 ( .A(n41511), .B(n41500), .Z(n41455) );
  XNOR U41432 ( .A(n41512), .B(n41495), .Z(n41500) );
  XOR U41433 ( .A(n41513), .B(n41514), .Z(n41495) );
  AND U41434 ( .A(n41515), .B(n41516), .Z(n41514) );
  XOR U41435 ( .A(n41517), .B(n41513), .Z(n41515) );
  XNOR U41436 ( .A(n41518), .B(n41519), .Z(n41512) );
  AND U41437 ( .A(n41520), .B(n41521), .Z(n41519) );
  XOR U41438 ( .A(n41518), .B(n41522), .Z(n41520) );
  XNOR U41439 ( .A(n41501), .B(n41498), .Z(n41511) );
  AND U41440 ( .A(n41523), .B(n41524), .Z(n41498) );
  XOR U41441 ( .A(n41525), .B(n41526), .Z(n41501) );
  AND U41442 ( .A(n41527), .B(n41528), .Z(n41526) );
  XOR U41443 ( .A(n41525), .B(n41529), .Z(n41527) );
  XNOR U41444 ( .A(n41452), .B(n41507), .Z(n41509) );
  XNOR U41445 ( .A(n41530), .B(n41531), .Z(n41452) );
  AND U41446 ( .A(n838), .B(n41532), .Z(n41531) );
  XNOR U41447 ( .A(n41533), .B(n41534), .Z(n41532) );
  XOR U41448 ( .A(n41535), .B(n41536), .Z(n41507) );
  AND U41449 ( .A(n41537), .B(n41538), .Z(n41536) );
  XNOR U41450 ( .A(n41535), .B(n41523), .Z(n41538) );
  IV U41451 ( .A(n41465), .Z(n41523) );
  XNOR U41452 ( .A(n41539), .B(n41516), .Z(n41465) );
  XNOR U41453 ( .A(n41540), .B(n41522), .Z(n41516) );
  XOR U41454 ( .A(n41541), .B(n41542), .Z(n41522) );
  AND U41455 ( .A(n41543), .B(n41544), .Z(n41542) );
  XOR U41456 ( .A(n41541), .B(n41545), .Z(n41543) );
  XNOR U41457 ( .A(n41521), .B(n41513), .Z(n41540) );
  XOR U41458 ( .A(n41546), .B(n41547), .Z(n41513) );
  AND U41459 ( .A(n41548), .B(n41549), .Z(n41547) );
  XNOR U41460 ( .A(n41550), .B(n41546), .Z(n41548) );
  XNOR U41461 ( .A(n41551), .B(n41518), .Z(n41521) );
  XOR U41462 ( .A(n41552), .B(n41553), .Z(n41518) );
  AND U41463 ( .A(n41554), .B(n41555), .Z(n41553) );
  XOR U41464 ( .A(n41552), .B(n41556), .Z(n41554) );
  XNOR U41465 ( .A(n41557), .B(n41558), .Z(n41551) );
  AND U41466 ( .A(n41559), .B(n41560), .Z(n41558) );
  XNOR U41467 ( .A(n41557), .B(n41561), .Z(n41559) );
  XNOR U41468 ( .A(n41517), .B(n41524), .Z(n41539) );
  AND U41469 ( .A(n41473), .B(n41562), .Z(n41524) );
  XOR U41470 ( .A(n41529), .B(n41528), .Z(n41517) );
  XNOR U41471 ( .A(n41563), .B(n41525), .Z(n41528) );
  XOR U41472 ( .A(n41564), .B(n41565), .Z(n41525) );
  AND U41473 ( .A(n41566), .B(n41567), .Z(n41565) );
  XOR U41474 ( .A(n41564), .B(n41568), .Z(n41566) );
  XNOR U41475 ( .A(n41569), .B(n41570), .Z(n41563) );
  AND U41476 ( .A(n41571), .B(n41572), .Z(n41570) );
  XOR U41477 ( .A(n41569), .B(n41573), .Z(n41571) );
  XOR U41478 ( .A(n41574), .B(n41575), .Z(n41529) );
  AND U41479 ( .A(n41576), .B(n41577), .Z(n41575) );
  XOR U41480 ( .A(n41574), .B(n41578), .Z(n41576) );
  XNOR U41481 ( .A(n41462), .B(n41535), .Z(n41537) );
  XNOR U41482 ( .A(n41579), .B(n41580), .Z(n41462) );
  AND U41483 ( .A(n838), .B(n41581), .Z(n41580) );
  XNOR U41484 ( .A(n41582), .B(n41583), .Z(n41581) );
  XOR U41485 ( .A(n41584), .B(n41585), .Z(n41535) );
  AND U41486 ( .A(n41586), .B(n41587), .Z(n41585) );
  XNOR U41487 ( .A(n41584), .B(n41473), .Z(n41587) );
  XOR U41488 ( .A(n41588), .B(n41549), .Z(n41473) );
  XNOR U41489 ( .A(n41589), .B(n41556), .Z(n41549) );
  XOR U41490 ( .A(n41545), .B(n41544), .Z(n41556) );
  XNOR U41491 ( .A(n41590), .B(n41541), .Z(n41544) );
  XOR U41492 ( .A(n41591), .B(n41592), .Z(n41541) );
  AND U41493 ( .A(n41593), .B(n41594), .Z(n41592) );
  XNOR U41494 ( .A(n41595), .B(n41596), .Z(n41593) );
  IV U41495 ( .A(n41591), .Z(n41595) );
  XNOR U41496 ( .A(n41597), .B(n41598), .Z(n41590) );
  NOR U41497 ( .A(n41599), .B(n41600), .Z(n41598) );
  XNOR U41498 ( .A(n41597), .B(n41601), .Z(n41599) );
  XOR U41499 ( .A(n41602), .B(n41603), .Z(n41545) );
  NOR U41500 ( .A(n41604), .B(n41605), .Z(n41603) );
  XNOR U41501 ( .A(n41602), .B(n41606), .Z(n41604) );
  XNOR U41502 ( .A(n41555), .B(n41546), .Z(n41589) );
  XOR U41503 ( .A(n41607), .B(n41608), .Z(n41546) );
  AND U41504 ( .A(n41609), .B(n41610), .Z(n41608) );
  XOR U41505 ( .A(n41607), .B(n41611), .Z(n41609) );
  XOR U41506 ( .A(n41612), .B(n41561), .Z(n41555) );
  XOR U41507 ( .A(n41613), .B(n41614), .Z(n41561) );
  NOR U41508 ( .A(n41615), .B(n41616), .Z(n41614) );
  XOR U41509 ( .A(n41613), .B(n41617), .Z(n41615) );
  XNOR U41510 ( .A(n41560), .B(n41552), .Z(n41612) );
  XOR U41511 ( .A(n41618), .B(n41619), .Z(n41552) );
  AND U41512 ( .A(n41620), .B(n41621), .Z(n41619) );
  XOR U41513 ( .A(n41618), .B(n41622), .Z(n41620) );
  XNOR U41514 ( .A(n41623), .B(n41557), .Z(n41560) );
  XOR U41515 ( .A(n41624), .B(n41625), .Z(n41557) );
  AND U41516 ( .A(n41626), .B(n41627), .Z(n41625) );
  XNOR U41517 ( .A(n41628), .B(n41629), .Z(n41626) );
  IV U41518 ( .A(n41624), .Z(n41628) );
  XNOR U41519 ( .A(n41630), .B(n41631), .Z(n41623) );
  NOR U41520 ( .A(n41632), .B(n41633), .Z(n41631) );
  XNOR U41521 ( .A(n41630), .B(n41634), .Z(n41632) );
  XOR U41522 ( .A(n41550), .B(n41562), .Z(n41588) );
  NOR U41523 ( .A(n41479), .B(n41635), .Z(n41562) );
  XNOR U41524 ( .A(n41568), .B(n41567), .Z(n41550) );
  XNOR U41525 ( .A(n41636), .B(n41573), .Z(n41567) );
  XNOR U41526 ( .A(n41637), .B(n41638), .Z(n41573) );
  NOR U41527 ( .A(n41639), .B(n41640), .Z(n41638) );
  XOR U41528 ( .A(n41637), .B(n41641), .Z(n41639) );
  XNOR U41529 ( .A(n41572), .B(n41564), .Z(n41636) );
  XOR U41530 ( .A(n41642), .B(n41643), .Z(n41564) );
  AND U41531 ( .A(n41644), .B(n41645), .Z(n41643) );
  XOR U41532 ( .A(n41642), .B(n41646), .Z(n41644) );
  XNOR U41533 ( .A(n41647), .B(n41569), .Z(n41572) );
  XOR U41534 ( .A(n41648), .B(n41649), .Z(n41569) );
  AND U41535 ( .A(n41650), .B(n41651), .Z(n41649) );
  XNOR U41536 ( .A(n41652), .B(n41653), .Z(n41650) );
  IV U41537 ( .A(n41648), .Z(n41652) );
  XNOR U41538 ( .A(n41654), .B(n41655), .Z(n41647) );
  NOR U41539 ( .A(n41656), .B(n41657), .Z(n41655) );
  XNOR U41540 ( .A(n41654), .B(n41658), .Z(n41656) );
  XOR U41541 ( .A(n41578), .B(n41577), .Z(n41568) );
  XNOR U41542 ( .A(n41659), .B(n41574), .Z(n41577) );
  XOR U41543 ( .A(n41660), .B(n41661), .Z(n41574) );
  AND U41544 ( .A(n41662), .B(n41663), .Z(n41661) );
  XNOR U41545 ( .A(n41664), .B(n41665), .Z(n41662) );
  IV U41546 ( .A(n41660), .Z(n41664) );
  XNOR U41547 ( .A(n41666), .B(n41667), .Z(n41659) );
  NOR U41548 ( .A(n41668), .B(n41669), .Z(n41667) );
  XNOR U41549 ( .A(n41666), .B(n41670), .Z(n41668) );
  XOR U41550 ( .A(n41671), .B(n41672), .Z(n41578) );
  NOR U41551 ( .A(n41673), .B(n41674), .Z(n41672) );
  XNOR U41552 ( .A(n41671), .B(n41675), .Z(n41673) );
  XNOR U41553 ( .A(n41470), .B(n41584), .Z(n41586) );
  XNOR U41554 ( .A(n41676), .B(n41677), .Z(n41470) );
  AND U41555 ( .A(n838), .B(n41678), .Z(n41677) );
  XNOR U41556 ( .A(n41679), .B(n41680), .Z(n41678) );
  AND U41557 ( .A(n41476), .B(n41479), .Z(n41584) );
  XOR U41558 ( .A(n41681), .B(n41635), .Z(n41479) );
  XNOR U41559 ( .A(p_input[1184]), .B(p_input[2048]), .Z(n41635) );
  XNOR U41560 ( .A(n41611), .B(n41610), .Z(n41681) );
  XNOR U41561 ( .A(n41682), .B(n41622), .Z(n41610) );
  XOR U41562 ( .A(n41596), .B(n41594), .Z(n41622) );
  XNOR U41563 ( .A(n41683), .B(n41601), .Z(n41594) );
  XOR U41564 ( .A(p_input[1208]), .B(p_input[2072]), .Z(n41601) );
  XOR U41565 ( .A(n41591), .B(n41600), .Z(n41683) );
  XOR U41566 ( .A(n41684), .B(n41597), .Z(n41600) );
  XOR U41567 ( .A(p_input[1206]), .B(p_input[2070]), .Z(n41597) );
  XOR U41568 ( .A(p_input[1207]), .B(n29410), .Z(n41684) );
  XOR U41569 ( .A(p_input[1202]), .B(p_input[2066]), .Z(n41591) );
  XNOR U41570 ( .A(n41606), .B(n41605), .Z(n41596) );
  XOR U41571 ( .A(n41685), .B(n41602), .Z(n41605) );
  XOR U41572 ( .A(p_input[1203]), .B(p_input[2067]), .Z(n41602) );
  XOR U41573 ( .A(p_input[1204]), .B(n29412), .Z(n41685) );
  XOR U41574 ( .A(p_input[1205]), .B(p_input[2069]), .Z(n41606) );
  XOR U41575 ( .A(n41621), .B(n41686), .Z(n41682) );
  IV U41576 ( .A(n41607), .Z(n41686) );
  XOR U41577 ( .A(p_input[1185]), .B(p_input[2049]), .Z(n41607) );
  XNOR U41578 ( .A(n41687), .B(n41629), .Z(n41621) );
  XNOR U41579 ( .A(n41617), .B(n41616), .Z(n41629) );
  XNOR U41580 ( .A(n41688), .B(n41613), .Z(n41616) );
  XNOR U41581 ( .A(p_input[1210]), .B(p_input[2074]), .Z(n41613) );
  XOR U41582 ( .A(p_input[1211]), .B(n29415), .Z(n41688) );
  XOR U41583 ( .A(p_input[1212]), .B(p_input[2076]), .Z(n41617) );
  XOR U41584 ( .A(n41627), .B(n41689), .Z(n41687) );
  IV U41585 ( .A(n41618), .Z(n41689) );
  XOR U41586 ( .A(p_input[1201]), .B(p_input[2065]), .Z(n41618) );
  XNOR U41587 ( .A(n41690), .B(n41634), .Z(n41627) );
  XNOR U41588 ( .A(p_input[1215]), .B(n29418), .Z(n41634) );
  XOR U41589 ( .A(n41624), .B(n41633), .Z(n41690) );
  XOR U41590 ( .A(n41691), .B(n41630), .Z(n41633) );
  XOR U41591 ( .A(p_input[1213]), .B(p_input[2077]), .Z(n41630) );
  XOR U41592 ( .A(p_input[1214]), .B(n29420), .Z(n41691) );
  XOR U41593 ( .A(p_input[1209]), .B(p_input[2073]), .Z(n41624) );
  XOR U41594 ( .A(n41646), .B(n41645), .Z(n41611) );
  XNOR U41595 ( .A(n41692), .B(n41653), .Z(n41645) );
  XNOR U41596 ( .A(n41641), .B(n41640), .Z(n41653) );
  XNOR U41597 ( .A(n41693), .B(n41637), .Z(n41640) );
  XNOR U41598 ( .A(p_input[1195]), .B(p_input[2059]), .Z(n41637) );
  XOR U41599 ( .A(p_input[1196]), .B(n28329), .Z(n41693) );
  XOR U41600 ( .A(p_input[1197]), .B(p_input[2061]), .Z(n41641) );
  XOR U41601 ( .A(n41651), .B(n41694), .Z(n41692) );
  IV U41602 ( .A(n41642), .Z(n41694) );
  XOR U41603 ( .A(p_input[1186]), .B(p_input[2050]), .Z(n41642) );
  XNOR U41604 ( .A(n41695), .B(n41658), .Z(n41651) );
  XNOR U41605 ( .A(p_input[1200]), .B(n28332), .Z(n41658) );
  XOR U41606 ( .A(n41648), .B(n41657), .Z(n41695) );
  XOR U41607 ( .A(n41696), .B(n41654), .Z(n41657) );
  XOR U41608 ( .A(p_input[1198]), .B(p_input[2062]), .Z(n41654) );
  XOR U41609 ( .A(p_input[1199]), .B(n28334), .Z(n41696) );
  XOR U41610 ( .A(p_input[1194]), .B(p_input[2058]), .Z(n41648) );
  XOR U41611 ( .A(n41665), .B(n41663), .Z(n41646) );
  XNOR U41612 ( .A(n41697), .B(n41670), .Z(n41663) );
  XOR U41613 ( .A(p_input[1193]), .B(p_input[2057]), .Z(n41670) );
  XOR U41614 ( .A(n41660), .B(n41669), .Z(n41697) );
  XOR U41615 ( .A(n41698), .B(n41666), .Z(n41669) );
  XOR U41616 ( .A(p_input[1191]), .B(p_input[2055]), .Z(n41666) );
  XOR U41617 ( .A(p_input[1192]), .B(n29427), .Z(n41698) );
  XOR U41618 ( .A(p_input[1187]), .B(p_input[2051]), .Z(n41660) );
  XNOR U41619 ( .A(n41675), .B(n41674), .Z(n41665) );
  XOR U41620 ( .A(n41699), .B(n41671), .Z(n41674) );
  XOR U41621 ( .A(p_input[1188]), .B(p_input[2052]), .Z(n41671) );
  XOR U41622 ( .A(p_input[1189]), .B(n29429), .Z(n41699) );
  XOR U41623 ( .A(p_input[1190]), .B(p_input[2054]), .Z(n41675) );
  XNOR U41624 ( .A(n41700), .B(n41701), .Z(n41476) );
  AND U41625 ( .A(n838), .B(n41702), .Z(n41701) );
  XNOR U41626 ( .A(n41703), .B(n41704), .Z(n838) );
  AND U41627 ( .A(n41705), .B(n41706), .Z(n41704) );
  XOR U41628 ( .A(n41490), .B(n41703), .Z(n41706) );
  XNOR U41629 ( .A(n41707), .B(n41703), .Z(n41705) );
  XOR U41630 ( .A(n41708), .B(n41709), .Z(n41703) );
  AND U41631 ( .A(n41710), .B(n41711), .Z(n41709) );
  XOR U41632 ( .A(n41505), .B(n41708), .Z(n41711) );
  XOR U41633 ( .A(n41708), .B(n41506), .Z(n41710) );
  XOR U41634 ( .A(n41712), .B(n41713), .Z(n41708) );
  AND U41635 ( .A(n41714), .B(n41715), .Z(n41713) );
  XOR U41636 ( .A(n41533), .B(n41712), .Z(n41715) );
  XOR U41637 ( .A(n41712), .B(n41534), .Z(n41714) );
  XOR U41638 ( .A(n41716), .B(n41717), .Z(n41712) );
  AND U41639 ( .A(n41718), .B(n41719), .Z(n41717) );
  XOR U41640 ( .A(n41582), .B(n41716), .Z(n41719) );
  XOR U41641 ( .A(n41716), .B(n41583), .Z(n41718) );
  XOR U41642 ( .A(n41720), .B(n41721), .Z(n41716) );
  AND U41643 ( .A(n41722), .B(n41723), .Z(n41721) );
  XOR U41644 ( .A(n41720), .B(n41679), .Z(n41723) );
  XNOR U41645 ( .A(n41724), .B(n41725), .Z(n41426) );
  AND U41646 ( .A(n842), .B(n41726), .Z(n41725) );
  XNOR U41647 ( .A(n41727), .B(n41728), .Z(n842) );
  AND U41648 ( .A(n41729), .B(n41730), .Z(n41728) );
  XOR U41649 ( .A(n41727), .B(n41436), .Z(n41730) );
  XNOR U41650 ( .A(n41727), .B(n41386), .Z(n41729) );
  XOR U41651 ( .A(n41731), .B(n41732), .Z(n41727) );
  AND U41652 ( .A(n41733), .B(n41734), .Z(n41732) );
  XNOR U41653 ( .A(n41446), .B(n41731), .Z(n41734) );
  XOR U41654 ( .A(n41731), .B(n41396), .Z(n41733) );
  XOR U41655 ( .A(n41735), .B(n41736), .Z(n41731) );
  AND U41656 ( .A(n41737), .B(n41738), .Z(n41736) );
  XNOR U41657 ( .A(n41456), .B(n41735), .Z(n41738) );
  XOR U41658 ( .A(n41735), .B(n41405), .Z(n41737) );
  XOR U41659 ( .A(n41739), .B(n41740), .Z(n41735) );
  AND U41660 ( .A(n41741), .B(n41742), .Z(n41740) );
  XOR U41661 ( .A(n41739), .B(n41413), .Z(n41741) );
  XOR U41662 ( .A(n41743), .B(n41744), .Z(n41377) );
  AND U41663 ( .A(n846), .B(n41726), .Z(n41744) );
  XNOR U41664 ( .A(n41724), .B(n41743), .Z(n41726) );
  XNOR U41665 ( .A(n41745), .B(n41746), .Z(n846) );
  AND U41666 ( .A(n41747), .B(n41748), .Z(n41746) );
  XNOR U41667 ( .A(n41749), .B(n41745), .Z(n41748) );
  IV U41668 ( .A(n41436), .Z(n41749) );
  XOR U41669 ( .A(n41707), .B(n41750), .Z(n41436) );
  AND U41670 ( .A(n849), .B(n41751), .Z(n41750) );
  XOR U41671 ( .A(n41489), .B(n41486), .Z(n41751) );
  IV U41672 ( .A(n41707), .Z(n41489) );
  XNOR U41673 ( .A(n41386), .B(n41745), .Z(n41747) );
  XOR U41674 ( .A(n41752), .B(n41753), .Z(n41386) );
  AND U41675 ( .A(n865), .B(n41754), .Z(n41753) );
  XOR U41676 ( .A(n41755), .B(n41756), .Z(n41745) );
  AND U41677 ( .A(n41757), .B(n41758), .Z(n41756) );
  XNOR U41678 ( .A(n41755), .B(n41446), .Z(n41758) );
  XOR U41679 ( .A(n41506), .B(n41759), .Z(n41446) );
  AND U41680 ( .A(n849), .B(n41760), .Z(n41759) );
  XOR U41681 ( .A(n41502), .B(n41506), .Z(n41760) );
  XNOR U41682 ( .A(n41761), .B(n41755), .Z(n41757) );
  IV U41683 ( .A(n41396), .Z(n41761) );
  XOR U41684 ( .A(n41762), .B(n41763), .Z(n41396) );
  AND U41685 ( .A(n865), .B(n41764), .Z(n41763) );
  XOR U41686 ( .A(n41765), .B(n41766), .Z(n41755) );
  AND U41687 ( .A(n41767), .B(n41768), .Z(n41766) );
  XNOR U41688 ( .A(n41765), .B(n41456), .Z(n41768) );
  XOR U41689 ( .A(n41534), .B(n41769), .Z(n41456) );
  AND U41690 ( .A(n849), .B(n41770), .Z(n41769) );
  XOR U41691 ( .A(n41530), .B(n41534), .Z(n41770) );
  XOR U41692 ( .A(n41405), .B(n41765), .Z(n41767) );
  XOR U41693 ( .A(n41771), .B(n41772), .Z(n41405) );
  AND U41694 ( .A(n865), .B(n41773), .Z(n41772) );
  XOR U41695 ( .A(n41739), .B(n41774), .Z(n41765) );
  AND U41696 ( .A(n41775), .B(n41742), .Z(n41774) );
  XNOR U41697 ( .A(n41466), .B(n41739), .Z(n41742) );
  XOR U41698 ( .A(n41583), .B(n41776), .Z(n41466) );
  AND U41699 ( .A(n849), .B(n41777), .Z(n41776) );
  XOR U41700 ( .A(n41579), .B(n41583), .Z(n41777) );
  XNOR U41701 ( .A(n41778), .B(n41739), .Z(n41775) );
  IV U41702 ( .A(n41413), .Z(n41778) );
  XOR U41703 ( .A(n41779), .B(n41780), .Z(n41413) );
  AND U41704 ( .A(n865), .B(n41781), .Z(n41780) );
  XOR U41705 ( .A(n41782), .B(n41783), .Z(n41739) );
  AND U41706 ( .A(n41784), .B(n41785), .Z(n41783) );
  XNOR U41707 ( .A(n41782), .B(n41474), .Z(n41785) );
  XOR U41708 ( .A(n41680), .B(n41786), .Z(n41474) );
  AND U41709 ( .A(n849), .B(n41787), .Z(n41786) );
  XOR U41710 ( .A(n41676), .B(n41680), .Z(n41787) );
  XNOR U41711 ( .A(n41788), .B(n41782), .Z(n41784) );
  IV U41712 ( .A(n41423), .Z(n41788) );
  XOR U41713 ( .A(n41789), .B(n41790), .Z(n41423) );
  AND U41714 ( .A(n865), .B(n41791), .Z(n41790) );
  AND U41715 ( .A(n41743), .B(n41724), .Z(n41782) );
  XNOR U41716 ( .A(n41792), .B(n41793), .Z(n41724) );
  AND U41717 ( .A(n849), .B(n41702), .Z(n41793) );
  XNOR U41718 ( .A(n41700), .B(n41792), .Z(n41702) );
  XNOR U41719 ( .A(n41794), .B(n41795), .Z(n849) );
  AND U41720 ( .A(n41796), .B(n41797), .Z(n41795) );
  XNOR U41721 ( .A(n41794), .B(n41486), .Z(n41797) );
  IV U41722 ( .A(n41490), .Z(n41486) );
  XOR U41723 ( .A(n41798), .B(n41799), .Z(n41490) );
  AND U41724 ( .A(n853), .B(n41800), .Z(n41799) );
  XOR U41725 ( .A(n41801), .B(n41798), .Z(n41800) );
  XNOR U41726 ( .A(n41794), .B(n41707), .Z(n41796) );
  XOR U41727 ( .A(n41802), .B(n41803), .Z(n41707) );
  AND U41728 ( .A(n861), .B(n41754), .Z(n41803) );
  XOR U41729 ( .A(n41752), .B(n41802), .Z(n41754) );
  XOR U41730 ( .A(n41804), .B(n41805), .Z(n41794) );
  AND U41731 ( .A(n41806), .B(n41807), .Z(n41805) );
  XNOR U41732 ( .A(n41804), .B(n41502), .Z(n41807) );
  IV U41733 ( .A(n41505), .Z(n41502) );
  XOR U41734 ( .A(n41808), .B(n41809), .Z(n41505) );
  AND U41735 ( .A(n853), .B(n41810), .Z(n41809) );
  XOR U41736 ( .A(n41811), .B(n41808), .Z(n41810) );
  XOR U41737 ( .A(n41506), .B(n41804), .Z(n41806) );
  XOR U41738 ( .A(n41812), .B(n41813), .Z(n41506) );
  AND U41739 ( .A(n861), .B(n41764), .Z(n41813) );
  XOR U41740 ( .A(n41812), .B(n41762), .Z(n41764) );
  XOR U41741 ( .A(n41814), .B(n41815), .Z(n41804) );
  AND U41742 ( .A(n41816), .B(n41817), .Z(n41815) );
  XNOR U41743 ( .A(n41814), .B(n41530), .Z(n41817) );
  IV U41744 ( .A(n41533), .Z(n41530) );
  XOR U41745 ( .A(n41818), .B(n41819), .Z(n41533) );
  AND U41746 ( .A(n853), .B(n41820), .Z(n41819) );
  XNOR U41747 ( .A(n41821), .B(n41818), .Z(n41820) );
  XOR U41748 ( .A(n41534), .B(n41814), .Z(n41816) );
  XOR U41749 ( .A(n41822), .B(n41823), .Z(n41534) );
  AND U41750 ( .A(n861), .B(n41773), .Z(n41823) );
  XOR U41751 ( .A(n41822), .B(n41771), .Z(n41773) );
  XOR U41752 ( .A(n41824), .B(n41825), .Z(n41814) );
  AND U41753 ( .A(n41826), .B(n41827), .Z(n41825) );
  XNOR U41754 ( .A(n41824), .B(n41579), .Z(n41827) );
  IV U41755 ( .A(n41582), .Z(n41579) );
  XOR U41756 ( .A(n41828), .B(n41829), .Z(n41582) );
  AND U41757 ( .A(n853), .B(n41830), .Z(n41829) );
  XOR U41758 ( .A(n41831), .B(n41828), .Z(n41830) );
  XOR U41759 ( .A(n41583), .B(n41824), .Z(n41826) );
  XOR U41760 ( .A(n41832), .B(n41833), .Z(n41583) );
  AND U41761 ( .A(n861), .B(n41781), .Z(n41833) );
  XOR U41762 ( .A(n41832), .B(n41779), .Z(n41781) );
  XOR U41763 ( .A(n41720), .B(n41834), .Z(n41824) );
  AND U41764 ( .A(n41722), .B(n41835), .Z(n41834) );
  XNOR U41765 ( .A(n41720), .B(n41676), .Z(n41835) );
  IV U41766 ( .A(n41679), .Z(n41676) );
  XOR U41767 ( .A(n41836), .B(n41837), .Z(n41679) );
  AND U41768 ( .A(n853), .B(n41838), .Z(n41837) );
  XNOR U41769 ( .A(n41839), .B(n41836), .Z(n41838) );
  XOR U41770 ( .A(n41680), .B(n41720), .Z(n41722) );
  XOR U41771 ( .A(n41840), .B(n41841), .Z(n41680) );
  AND U41772 ( .A(n861), .B(n41791), .Z(n41841) );
  XOR U41773 ( .A(n41840), .B(n41789), .Z(n41791) );
  AND U41774 ( .A(n41792), .B(n41700), .Z(n41720) );
  XNOR U41775 ( .A(n41842), .B(n41843), .Z(n41700) );
  AND U41776 ( .A(n853), .B(n41844), .Z(n41843) );
  XNOR U41777 ( .A(n41845), .B(n41842), .Z(n41844) );
  XNOR U41778 ( .A(n41846), .B(n41847), .Z(n853) );
  AND U41779 ( .A(n41848), .B(n41849), .Z(n41847) );
  XOR U41780 ( .A(n41801), .B(n41846), .Z(n41849) );
  AND U41781 ( .A(n41850), .B(n41851), .Z(n41801) );
  XNOR U41782 ( .A(n41798), .B(n41846), .Z(n41848) );
  XNOR U41783 ( .A(n41852), .B(n41853), .Z(n41798) );
  AND U41784 ( .A(n857), .B(n41854), .Z(n41853) );
  XNOR U41785 ( .A(n41855), .B(n41856), .Z(n41854) );
  XOR U41786 ( .A(n41857), .B(n41858), .Z(n41846) );
  AND U41787 ( .A(n41859), .B(n41860), .Z(n41858) );
  XNOR U41788 ( .A(n41857), .B(n41850), .Z(n41860) );
  IV U41789 ( .A(n41811), .Z(n41850) );
  XOR U41790 ( .A(n41861), .B(n41862), .Z(n41811) );
  XOR U41791 ( .A(n41863), .B(n41851), .Z(n41862) );
  AND U41792 ( .A(n41821), .B(n41864), .Z(n41851) );
  AND U41793 ( .A(n41865), .B(n41866), .Z(n41863) );
  XOR U41794 ( .A(n41867), .B(n41861), .Z(n41865) );
  XNOR U41795 ( .A(n41808), .B(n41857), .Z(n41859) );
  XNOR U41796 ( .A(n41868), .B(n41869), .Z(n41808) );
  AND U41797 ( .A(n857), .B(n41870), .Z(n41869) );
  XNOR U41798 ( .A(n41871), .B(n41872), .Z(n41870) );
  XOR U41799 ( .A(n41873), .B(n41874), .Z(n41857) );
  AND U41800 ( .A(n41875), .B(n41876), .Z(n41874) );
  XNOR U41801 ( .A(n41873), .B(n41821), .Z(n41876) );
  XOR U41802 ( .A(n41877), .B(n41866), .Z(n41821) );
  XNOR U41803 ( .A(n41878), .B(n41861), .Z(n41866) );
  XOR U41804 ( .A(n41879), .B(n41880), .Z(n41861) );
  AND U41805 ( .A(n41881), .B(n41882), .Z(n41880) );
  XOR U41806 ( .A(n41883), .B(n41879), .Z(n41881) );
  XNOR U41807 ( .A(n41884), .B(n41885), .Z(n41878) );
  AND U41808 ( .A(n41886), .B(n41887), .Z(n41885) );
  XOR U41809 ( .A(n41884), .B(n41888), .Z(n41886) );
  XNOR U41810 ( .A(n41867), .B(n41864), .Z(n41877) );
  AND U41811 ( .A(n41889), .B(n41890), .Z(n41864) );
  XOR U41812 ( .A(n41891), .B(n41892), .Z(n41867) );
  AND U41813 ( .A(n41893), .B(n41894), .Z(n41892) );
  XOR U41814 ( .A(n41891), .B(n41895), .Z(n41893) );
  XNOR U41815 ( .A(n41818), .B(n41873), .Z(n41875) );
  XNOR U41816 ( .A(n41896), .B(n41897), .Z(n41818) );
  AND U41817 ( .A(n857), .B(n41898), .Z(n41897) );
  XNOR U41818 ( .A(n41899), .B(n41900), .Z(n41898) );
  XOR U41819 ( .A(n41901), .B(n41902), .Z(n41873) );
  AND U41820 ( .A(n41903), .B(n41904), .Z(n41902) );
  XNOR U41821 ( .A(n41901), .B(n41889), .Z(n41904) );
  IV U41822 ( .A(n41831), .Z(n41889) );
  XNOR U41823 ( .A(n41905), .B(n41882), .Z(n41831) );
  XNOR U41824 ( .A(n41906), .B(n41888), .Z(n41882) );
  XOR U41825 ( .A(n41907), .B(n41908), .Z(n41888) );
  AND U41826 ( .A(n41909), .B(n41910), .Z(n41908) );
  XOR U41827 ( .A(n41907), .B(n41911), .Z(n41909) );
  XNOR U41828 ( .A(n41887), .B(n41879), .Z(n41906) );
  XOR U41829 ( .A(n41912), .B(n41913), .Z(n41879) );
  AND U41830 ( .A(n41914), .B(n41915), .Z(n41913) );
  XNOR U41831 ( .A(n41916), .B(n41912), .Z(n41914) );
  XNOR U41832 ( .A(n41917), .B(n41884), .Z(n41887) );
  XOR U41833 ( .A(n41918), .B(n41919), .Z(n41884) );
  AND U41834 ( .A(n41920), .B(n41921), .Z(n41919) );
  XOR U41835 ( .A(n41918), .B(n41922), .Z(n41920) );
  XNOR U41836 ( .A(n41923), .B(n41924), .Z(n41917) );
  AND U41837 ( .A(n41925), .B(n41926), .Z(n41924) );
  XNOR U41838 ( .A(n41923), .B(n41927), .Z(n41925) );
  XNOR U41839 ( .A(n41883), .B(n41890), .Z(n41905) );
  AND U41840 ( .A(n41839), .B(n41928), .Z(n41890) );
  XOR U41841 ( .A(n41895), .B(n41894), .Z(n41883) );
  XNOR U41842 ( .A(n41929), .B(n41891), .Z(n41894) );
  XOR U41843 ( .A(n41930), .B(n41931), .Z(n41891) );
  AND U41844 ( .A(n41932), .B(n41933), .Z(n41931) );
  XOR U41845 ( .A(n41930), .B(n41934), .Z(n41932) );
  XNOR U41846 ( .A(n41935), .B(n41936), .Z(n41929) );
  AND U41847 ( .A(n41937), .B(n41938), .Z(n41936) );
  XOR U41848 ( .A(n41935), .B(n41939), .Z(n41937) );
  XOR U41849 ( .A(n41940), .B(n41941), .Z(n41895) );
  AND U41850 ( .A(n41942), .B(n41943), .Z(n41941) );
  XOR U41851 ( .A(n41940), .B(n41944), .Z(n41942) );
  XNOR U41852 ( .A(n41828), .B(n41901), .Z(n41903) );
  XNOR U41853 ( .A(n41945), .B(n41946), .Z(n41828) );
  AND U41854 ( .A(n857), .B(n41947), .Z(n41946) );
  XNOR U41855 ( .A(n41948), .B(n41949), .Z(n41947) );
  XOR U41856 ( .A(n41950), .B(n41951), .Z(n41901) );
  AND U41857 ( .A(n41952), .B(n41953), .Z(n41951) );
  XNOR U41858 ( .A(n41950), .B(n41839), .Z(n41953) );
  XOR U41859 ( .A(n41954), .B(n41915), .Z(n41839) );
  XNOR U41860 ( .A(n41955), .B(n41922), .Z(n41915) );
  XOR U41861 ( .A(n41911), .B(n41910), .Z(n41922) );
  XNOR U41862 ( .A(n41956), .B(n41907), .Z(n41910) );
  XOR U41863 ( .A(n41957), .B(n41958), .Z(n41907) );
  AND U41864 ( .A(n41959), .B(n41960), .Z(n41958) );
  XNOR U41865 ( .A(n41961), .B(n41962), .Z(n41959) );
  IV U41866 ( .A(n41957), .Z(n41961) );
  XNOR U41867 ( .A(n41963), .B(n41964), .Z(n41956) );
  NOR U41868 ( .A(n41965), .B(n41966), .Z(n41964) );
  XNOR U41869 ( .A(n41963), .B(n41967), .Z(n41965) );
  XOR U41870 ( .A(n41968), .B(n41969), .Z(n41911) );
  NOR U41871 ( .A(n41970), .B(n41971), .Z(n41969) );
  XNOR U41872 ( .A(n41968), .B(n41972), .Z(n41970) );
  XNOR U41873 ( .A(n41921), .B(n41912), .Z(n41955) );
  XOR U41874 ( .A(n41973), .B(n41974), .Z(n41912) );
  AND U41875 ( .A(n41975), .B(n41976), .Z(n41974) );
  XOR U41876 ( .A(n41973), .B(n41977), .Z(n41975) );
  XOR U41877 ( .A(n41978), .B(n41927), .Z(n41921) );
  XOR U41878 ( .A(n41979), .B(n41980), .Z(n41927) );
  NOR U41879 ( .A(n41981), .B(n41982), .Z(n41980) );
  XOR U41880 ( .A(n41979), .B(n41983), .Z(n41981) );
  XNOR U41881 ( .A(n41926), .B(n41918), .Z(n41978) );
  XOR U41882 ( .A(n41984), .B(n41985), .Z(n41918) );
  AND U41883 ( .A(n41986), .B(n41987), .Z(n41985) );
  XOR U41884 ( .A(n41984), .B(n41988), .Z(n41986) );
  XNOR U41885 ( .A(n41989), .B(n41923), .Z(n41926) );
  XOR U41886 ( .A(n41990), .B(n41991), .Z(n41923) );
  AND U41887 ( .A(n41992), .B(n41993), .Z(n41991) );
  XNOR U41888 ( .A(n41994), .B(n41995), .Z(n41992) );
  IV U41889 ( .A(n41990), .Z(n41994) );
  XNOR U41890 ( .A(n41996), .B(n41997), .Z(n41989) );
  NOR U41891 ( .A(n41998), .B(n41999), .Z(n41997) );
  XNOR U41892 ( .A(n41996), .B(n42000), .Z(n41998) );
  XOR U41893 ( .A(n41916), .B(n41928), .Z(n41954) );
  NOR U41894 ( .A(n41845), .B(n42001), .Z(n41928) );
  XNOR U41895 ( .A(n41934), .B(n41933), .Z(n41916) );
  XNOR U41896 ( .A(n42002), .B(n41939), .Z(n41933) );
  XNOR U41897 ( .A(n42003), .B(n42004), .Z(n41939) );
  NOR U41898 ( .A(n42005), .B(n42006), .Z(n42004) );
  XOR U41899 ( .A(n42003), .B(n42007), .Z(n42005) );
  XNOR U41900 ( .A(n41938), .B(n41930), .Z(n42002) );
  XOR U41901 ( .A(n42008), .B(n42009), .Z(n41930) );
  AND U41902 ( .A(n42010), .B(n42011), .Z(n42009) );
  XOR U41903 ( .A(n42008), .B(n42012), .Z(n42010) );
  XNOR U41904 ( .A(n42013), .B(n41935), .Z(n41938) );
  XOR U41905 ( .A(n42014), .B(n42015), .Z(n41935) );
  AND U41906 ( .A(n42016), .B(n42017), .Z(n42015) );
  XNOR U41907 ( .A(n42018), .B(n42019), .Z(n42016) );
  IV U41908 ( .A(n42014), .Z(n42018) );
  XNOR U41909 ( .A(n42020), .B(n42021), .Z(n42013) );
  NOR U41910 ( .A(n42022), .B(n42023), .Z(n42021) );
  XNOR U41911 ( .A(n42020), .B(n42024), .Z(n42022) );
  XOR U41912 ( .A(n41944), .B(n41943), .Z(n41934) );
  XNOR U41913 ( .A(n42025), .B(n41940), .Z(n41943) );
  XOR U41914 ( .A(n42026), .B(n42027), .Z(n41940) );
  AND U41915 ( .A(n42028), .B(n42029), .Z(n42027) );
  XNOR U41916 ( .A(n42030), .B(n42031), .Z(n42028) );
  IV U41917 ( .A(n42026), .Z(n42030) );
  XNOR U41918 ( .A(n42032), .B(n42033), .Z(n42025) );
  NOR U41919 ( .A(n42034), .B(n42035), .Z(n42033) );
  XNOR U41920 ( .A(n42032), .B(n42036), .Z(n42034) );
  XOR U41921 ( .A(n42037), .B(n42038), .Z(n41944) );
  NOR U41922 ( .A(n42039), .B(n42040), .Z(n42038) );
  XNOR U41923 ( .A(n42037), .B(n42041), .Z(n42039) );
  XNOR U41924 ( .A(n41836), .B(n41950), .Z(n41952) );
  XNOR U41925 ( .A(n42042), .B(n42043), .Z(n41836) );
  AND U41926 ( .A(n857), .B(n42044), .Z(n42043) );
  XNOR U41927 ( .A(n42045), .B(n42046), .Z(n42044) );
  AND U41928 ( .A(n41842), .B(n41845), .Z(n41950) );
  XOR U41929 ( .A(n42047), .B(n42001), .Z(n41845) );
  XNOR U41930 ( .A(p_input[1216]), .B(p_input[2048]), .Z(n42001) );
  XNOR U41931 ( .A(n41977), .B(n41976), .Z(n42047) );
  XNOR U41932 ( .A(n42048), .B(n41988), .Z(n41976) );
  XOR U41933 ( .A(n41962), .B(n41960), .Z(n41988) );
  XNOR U41934 ( .A(n42049), .B(n41967), .Z(n41960) );
  XOR U41935 ( .A(p_input[1240]), .B(p_input[2072]), .Z(n41967) );
  XOR U41936 ( .A(n41957), .B(n41966), .Z(n42049) );
  XOR U41937 ( .A(n42050), .B(n41963), .Z(n41966) );
  XOR U41938 ( .A(p_input[1238]), .B(p_input[2070]), .Z(n41963) );
  XOR U41939 ( .A(p_input[1239]), .B(n29410), .Z(n42050) );
  XOR U41940 ( .A(p_input[1234]), .B(p_input[2066]), .Z(n41957) );
  XNOR U41941 ( .A(n41972), .B(n41971), .Z(n41962) );
  XOR U41942 ( .A(n42051), .B(n41968), .Z(n41971) );
  XOR U41943 ( .A(p_input[1235]), .B(p_input[2067]), .Z(n41968) );
  XOR U41944 ( .A(p_input[1236]), .B(n29412), .Z(n42051) );
  XOR U41945 ( .A(p_input[1237]), .B(p_input[2069]), .Z(n41972) );
  XOR U41946 ( .A(n41987), .B(n42052), .Z(n42048) );
  IV U41947 ( .A(n41973), .Z(n42052) );
  XOR U41948 ( .A(p_input[1217]), .B(p_input[2049]), .Z(n41973) );
  XNOR U41949 ( .A(n42053), .B(n41995), .Z(n41987) );
  XNOR U41950 ( .A(n41983), .B(n41982), .Z(n41995) );
  XNOR U41951 ( .A(n42054), .B(n41979), .Z(n41982) );
  XNOR U41952 ( .A(p_input[1242]), .B(p_input[2074]), .Z(n41979) );
  XOR U41953 ( .A(p_input[1243]), .B(n29415), .Z(n42054) );
  XOR U41954 ( .A(p_input[1244]), .B(p_input[2076]), .Z(n41983) );
  XOR U41955 ( .A(n41993), .B(n42055), .Z(n42053) );
  IV U41956 ( .A(n41984), .Z(n42055) );
  XOR U41957 ( .A(p_input[1233]), .B(p_input[2065]), .Z(n41984) );
  XNOR U41958 ( .A(n42056), .B(n42000), .Z(n41993) );
  XNOR U41959 ( .A(p_input[1247]), .B(n29418), .Z(n42000) );
  XOR U41960 ( .A(n41990), .B(n41999), .Z(n42056) );
  XOR U41961 ( .A(n42057), .B(n41996), .Z(n41999) );
  XOR U41962 ( .A(p_input[1245]), .B(p_input[2077]), .Z(n41996) );
  XOR U41963 ( .A(p_input[1246]), .B(n29420), .Z(n42057) );
  XOR U41964 ( .A(p_input[1241]), .B(p_input[2073]), .Z(n41990) );
  XOR U41965 ( .A(n42012), .B(n42011), .Z(n41977) );
  XNOR U41966 ( .A(n42058), .B(n42019), .Z(n42011) );
  XNOR U41967 ( .A(n42007), .B(n42006), .Z(n42019) );
  XNOR U41968 ( .A(n42059), .B(n42003), .Z(n42006) );
  XNOR U41969 ( .A(p_input[1227]), .B(p_input[2059]), .Z(n42003) );
  XOR U41970 ( .A(p_input[1228]), .B(n28329), .Z(n42059) );
  XOR U41971 ( .A(p_input[1229]), .B(p_input[2061]), .Z(n42007) );
  XOR U41972 ( .A(n42017), .B(n42060), .Z(n42058) );
  IV U41973 ( .A(n42008), .Z(n42060) );
  XOR U41974 ( .A(p_input[1218]), .B(p_input[2050]), .Z(n42008) );
  XNOR U41975 ( .A(n42061), .B(n42024), .Z(n42017) );
  XNOR U41976 ( .A(p_input[1232]), .B(n28332), .Z(n42024) );
  XOR U41977 ( .A(n42014), .B(n42023), .Z(n42061) );
  XOR U41978 ( .A(n42062), .B(n42020), .Z(n42023) );
  XOR U41979 ( .A(p_input[1230]), .B(p_input[2062]), .Z(n42020) );
  XOR U41980 ( .A(p_input[1231]), .B(n28334), .Z(n42062) );
  XOR U41981 ( .A(p_input[1226]), .B(p_input[2058]), .Z(n42014) );
  XOR U41982 ( .A(n42031), .B(n42029), .Z(n42012) );
  XNOR U41983 ( .A(n42063), .B(n42036), .Z(n42029) );
  XOR U41984 ( .A(p_input[1225]), .B(p_input[2057]), .Z(n42036) );
  XOR U41985 ( .A(n42026), .B(n42035), .Z(n42063) );
  XOR U41986 ( .A(n42064), .B(n42032), .Z(n42035) );
  XOR U41987 ( .A(p_input[1223]), .B(p_input[2055]), .Z(n42032) );
  XOR U41988 ( .A(p_input[1224]), .B(n29427), .Z(n42064) );
  XOR U41989 ( .A(p_input[1219]), .B(p_input[2051]), .Z(n42026) );
  XNOR U41990 ( .A(n42041), .B(n42040), .Z(n42031) );
  XOR U41991 ( .A(n42065), .B(n42037), .Z(n42040) );
  XOR U41992 ( .A(p_input[1220]), .B(p_input[2052]), .Z(n42037) );
  XOR U41993 ( .A(p_input[1221]), .B(n29429), .Z(n42065) );
  XOR U41994 ( .A(p_input[1222]), .B(p_input[2054]), .Z(n42041) );
  XNOR U41995 ( .A(n42066), .B(n42067), .Z(n41842) );
  AND U41996 ( .A(n857), .B(n42068), .Z(n42067) );
  XNOR U41997 ( .A(n42069), .B(n42070), .Z(n857) );
  AND U41998 ( .A(n42071), .B(n42072), .Z(n42070) );
  XOR U41999 ( .A(n41856), .B(n42069), .Z(n42072) );
  XNOR U42000 ( .A(n42073), .B(n42069), .Z(n42071) );
  XOR U42001 ( .A(n42074), .B(n42075), .Z(n42069) );
  AND U42002 ( .A(n42076), .B(n42077), .Z(n42075) );
  XOR U42003 ( .A(n41871), .B(n42074), .Z(n42077) );
  XOR U42004 ( .A(n42074), .B(n41872), .Z(n42076) );
  XOR U42005 ( .A(n42078), .B(n42079), .Z(n42074) );
  AND U42006 ( .A(n42080), .B(n42081), .Z(n42079) );
  XOR U42007 ( .A(n41899), .B(n42078), .Z(n42081) );
  XOR U42008 ( .A(n42078), .B(n41900), .Z(n42080) );
  XOR U42009 ( .A(n42082), .B(n42083), .Z(n42078) );
  AND U42010 ( .A(n42084), .B(n42085), .Z(n42083) );
  XOR U42011 ( .A(n41948), .B(n42082), .Z(n42085) );
  XOR U42012 ( .A(n42082), .B(n41949), .Z(n42084) );
  XOR U42013 ( .A(n42086), .B(n42087), .Z(n42082) );
  AND U42014 ( .A(n42088), .B(n42089), .Z(n42087) );
  XOR U42015 ( .A(n42086), .B(n42045), .Z(n42089) );
  XNOR U42016 ( .A(n42090), .B(n42091), .Z(n41792) );
  AND U42017 ( .A(n861), .B(n42092), .Z(n42091) );
  XNOR U42018 ( .A(n42093), .B(n42094), .Z(n861) );
  AND U42019 ( .A(n42095), .B(n42096), .Z(n42094) );
  XOR U42020 ( .A(n42093), .B(n41802), .Z(n42096) );
  XNOR U42021 ( .A(n42093), .B(n41752), .Z(n42095) );
  XOR U42022 ( .A(n42097), .B(n42098), .Z(n42093) );
  AND U42023 ( .A(n42099), .B(n42100), .Z(n42098) );
  XNOR U42024 ( .A(n41812), .B(n42097), .Z(n42100) );
  XOR U42025 ( .A(n42097), .B(n41762), .Z(n42099) );
  XOR U42026 ( .A(n42101), .B(n42102), .Z(n42097) );
  AND U42027 ( .A(n42103), .B(n42104), .Z(n42102) );
  XNOR U42028 ( .A(n41822), .B(n42101), .Z(n42104) );
  XOR U42029 ( .A(n42101), .B(n41771), .Z(n42103) );
  XOR U42030 ( .A(n42105), .B(n42106), .Z(n42101) );
  AND U42031 ( .A(n42107), .B(n42108), .Z(n42106) );
  XOR U42032 ( .A(n42105), .B(n41779), .Z(n42107) );
  XOR U42033 ( .A(n42109), .B(n42110), .Z(n41743) );
  AND U42034 ( .A(n865), .B(n42092), .Z(n42110) );
  XNOR U42035 ( .A(n42090), .B(n42109), .Z(n42092) );
  XNOR U42036 ( .A(n42111), .B(n42112), .Z(n865) );
  AND U42037 ( .A(n42113), .B(n42114), .Z(n42112) );
  XNOR U42038 ( .A(n42115), .B(n42111), .Z(n42114) );
  IV U42039 ( .A(n41802), .Z(n42115) );
  XOR U42040 ( .A(n42073), .B(n42116), .Z(n41802) );
  AND U42041 ( .A(n868), .B(n42117), .Z(n42116) );
  XOR U42042 ( .A(n41855), .B(n41852), .Z(n42117) );
  IV U42043 ( .A(n42073), .Z(n41855) );
  XNOR U42044 ( .A(n41752), .B(n42111), .Z(n42113) );
  XOR U42045 ( .A(n42118), .B(n42119), .Z(n41752) );
  AND U42046 ( .A(n884), .B(n42120), .Z(n42119) );
  XOR U42047 ( .A(n42121), .B(n42122), .Z(n42111) );
  AND U42048 ( .A(n42123), .B(n42124), .Z(n42122) );
  XNOR U42049 ( .A(n42121), .B(n41812), .Z(n42124) );
  XOR U42050 ( .A(n41872), .B(n42125), .Z(n41812) );
  AND U42051 ( .A(n868), .B(n42126), .Z(n42125) );
  XOR U42052 ( .A(n41868), .B(n41872), .Z(n42126) );
  XNOR U42053 ( .A(n42127), .B(n42121), .Z(n42123) );
  IV U42054 ( .A(n41762), .Z(n42127) );
  XOR U42055 ( .A(n42128), .B(n42129), .Z(n41762) );
  AND U42056 ( .A(n884), .B(n42130), .Z(n42129) );
  XOR U42057 ( .A(n42131), .B(n42132), .Z(n42121) );
  AND U42058 ( .A(n42133), .B(n42134), .Z(n42132) );
  XNOR U42059 ( .A(n42131), .B(n41822), .Z(n42134) );
  XOR U42060 ( .A(n41900), .B(n42135), .Z(n41822) );
  AND U42061 ( .A(n868), .B(n42136), .Z(n42135) );
  XOR U42062 ( .A(n41896), .B(n41900), .Z(n42136) );
  XOR U42063 ( .A(n41771), .B(n42131), .Z(n42133) );
  XOR U42064 ( .A(n42137), .B(n42138), .Z(n41771) );
  AND U42065 ( .A(n884), .B(n42139), .Z(n42138) );
  XOR U42066 ( .A(n42105), .B(n42140), .Z(n42131) );
  AND U42067 ( .A(n42141), .B(n42108), .Z(n42140) );
  XNOR U42068 ( .A(n41832), .B(n42105), .Z(n42108) );
  XOR U42069 ( .A(n41949), .B(n42142), .Z(n41832) );
  AND U42070 ( .A(n868), .B(n42143), .Z(n42142) );
  XOR U42071 ( .A(n41945), .B(n41949), .Z(n42143) );
  XNOR U42072 ( .A(n42144), .B(n42105), .Z(n42141) );
  IV U42073 ( .A(n41779), .Z(n42144) );
  XOR U42074 ( .A(n42145), .B(n42146), .Z(n41779) );
  AND U42075 ( .A(n884), .B(n42147), .Z(n42146) );
  XOR U42076 ( .A(n42148), .B(n42149), .Z(n42105) );
  AND U42077 ( .A(n42150), .B(n42151), .Z(n42149) );
  XNOR U42078 ( .A(n42148), .B(n41840), .Z(n42151) );
  XOR U42079 ( .A(n42046), .B(n42152), .Z(n41840) );
  AND U42080 ( .A(n868), .B(n42153), .Z(n42152) );
  XOR U42081 ( .A(n42042), .B(n42046), .Z(n42153) );
  XNOR U42082 ( .A(n42154), .B(n42148), .Z(n42150) );
  IV U42083 ( .A(n41789), .Z(n42154) );
  XOR U42084 ( .A(n42155), .B(n42156), .Z(n41789) );
  AND U42085 ( .A(n884), .B(n42157), .Z(n42156) );
  AND U42086 ( .A(n42109), .B(n42090), .Z(n42148) );
  XNOR U42087 ( .A(n42158), .B(n42159), .Z(n42090) );
  AND U42088 ( .A(n868), .B(n42068), .Z(n42159) );
  XNOR U42089 ( .A(n42066), .B(n42158), .Z(n42068) );
  XNOR U42090 ( .A(n42160), .B(n42161), .Z(n868) );
  AND U42091 ( .A(n42162), .B(n42163), .Z(n42161) );
  XNOR U42092 ( .A(n42160), .B(n41852), .Z(n42163) );
  IV U42093 ( .A(n41856), .Z(n41852) );
  XOR U42094 ( .A(n42164), .B(n42165), .Z(n41856) );
  AND U42095 ( .A(n872), .B(n42166), .Z(n42165) );
  XOR U42096 ( .A(n42167), .B(n42164), .Z(n42166) );
  XNOR U42097 ( .A(n42160), .B(n42073), .Z(n42162) );
  XOR U42098 ( .A(n42168), .B(n42169), .Z(n42073) );
  AND U42099 ( .A(n880), .B(n42120), .Z(n42169) );
  XOR U42100 ( .A(n42118), .B(n42168), .Z(n42120) );
  XOR U42101 ( .A(n42170), .B(n42171), .Z(n42160) );
  AND U42102 ( .A(n42172), .B(n42173), .Z(n42171) );
  XNOR U42103 ( .A(n42170), .B(n41868), .Z(n42173) );
  IV U42104 ( .A(n41871), .Z(n41868) );
  XOR U42105 ( .A(n42174), .B(n42175), .Z(n41871) );
  AND U42106 ( .A(n872), .B(n42176), .Z(n42175) );
  XOR U42107 ( .A(n42177), .B(n42174), .Z(n42176) );
  XOR U42108 ( .A(n41872), .B(n42170), .Z(n42172) );
  XOR U42109 ( .A(n42178), .B(n42179), .Z(n41872) );
  AND U42110 ( .A(n880), .B(n42130), .Z(n42179) );
  XOR U42111 ( .A(n42178), .B(n42128), .Z(n42130) );
  XOR U42112 ( .A(n42180), .B(n42181), .Z(n42170) );
  AND U42113 ( .A(n42182), .B(n42183), .Z(n42181) );
  XNOR U42114 ( .A(n42180), .B(n41896), .Z(n42183) );
  IV U42115 ( .A(n41899), .Z(n41896) );
  XOR U42116 ( .A(n42184), .B(n42185), .Z(n41899) );
  AND U42117 ( .A(n872), .B(n42186), .Z(n42185) );
  XNOR U42118 ( .A(n42187), .B(n42184), .Z(n42186) );
  XOR U42119 ( .A(n41900), .B(n42180), .Z(n42182) );
  XOR U42120 ( .A(n42188), .B(n42189), .Z(n41900) );
  AND U42121 ( .A(n880), .B(n42139), .Z(n42189) );
  XOR U42122 ( .A(n42188), .B(n42137), .Z(n42139) );
  XOR U42123 ( .A(n42190), .B(n42191), .Z(n42180) );
  AND U42124 ( .A(n42192), .B(n42193), .Z(n42191) );
  XNOR U42125 ( .A(n42190), .B(n41945), .Z(n42193) );
  IV U42126 ( .A(n41948), .Z(n41945) );
  XOR U42127 ( .A(n42194), .B(n42195), .Z(n41948) );
  AND U42128 ( .A(n872), .B(n42196), .Z(n42195) );
  XOR U42129 ( .A(n42197), .B(n42194), .Z(n42196) );
  XOR U42130 ( .A(n41949), .B(n42190), .Z(n42192) );
  XOR U42131 ( .A(n42198), .B(n42199), .Z(n41949) );
  AND U42132 ( .A(n880), .B(n42147), .Z(n42199) );
  XOR U42133 ( .A(n42198), .B(n42145), .Z(n42147) );
  XOR U42134 ( .A(n42086), .B(n42200), .Z(n42190) );
  AND U42135 ( .A(n42088), .B(n42201), .Z(n42200) );
  XNOR U42136 ( .A(n42086), .B(n42042), .Z(n42201) );
  IV U42137 ( .A(n42045), .Z(n42042) );
  XOR U42138 ( .A(n42202), .B(n42203), .Z(n42045) );
  AND U42139 ( .A(n872), .B(n42204), .Z(n42203) );
  XNOR U42140 ( .A(n42205), .B(n42202), .Z(n42204) );
  XOR U42141 ( .A(n42046), .B(n42086), .Z(n42088) );
  XOR U42142 ( .A(n42206), .B(n42207), .Z(n42046) );
  AND U42143 ( .A(n880), .B(n42157), .Z(n42207) );
  XOR U42144 ( .A(n42206), .B(n42155), .Z(n42157) );
  AND U42145 ( .A(n42158), .B(n42066), .Z(n42086) );
  XNOR U42146 ( .A(n42208), .B(n42209), .Z(n42066) );
  AND U42147 ( .A(n872), .B(n42210), .Z(n42209) );
  XNOR U42148 ( .A(n42211), .B(n42208), .Z(n42210) );
  XNOR U42149 ( .A(n42212), .B(n42213), .Z(n872) );
  AND U42150 ( .A(n42214), .B(n42215), .Z(n42213) );
  XOR U42151 ( .A(n42167), .B(n42212), .Z(n42215) );
  AND U42152 ( .A(n42216), .B(n42217), .Z(n42167) );
  XNOR U42153 ( .A(n42164), .B(n42212), .Z(n42214) );
  XNOR U42154 ( .A(n42218), .B(n42219), .Z(n42164) );
  AND U42155 ( .A(n876), .B(n42220), .Z(n42219) );
  XNOR U42156 ( .A(n42221), .B(n42222), .Z(n42220) );
  XOR U42157 ( .A(n42223), .B(n42224), .Z(n42212) );
  AND U42158 ( .A(n42225), .B(n42226), .Z(n42224) );
  XNOR U42159 ( .A(n42223), .B(n42216), .Z(n42226) );
  IV U42160 ( .A(n42177), .Z(n42216) );
  XOR U42161 ( .A(n42227), .B(n42228), .Z(n42177) );
  XOR U42162 ( .A(n42229), .B(n42217), .Z(n42228) );
  AND U42163 ( .A(n42187), .B(n42230), .Z(n42217) );
  AND U42164 ( .A(n42231), .B(n42232), .Z(n42229) );
  XOR U42165 ( .A(n42233), .B(n42227), .Z(n42231) );
  XNOR U42166 ( .A(n42174), .B(n42223), .Z(n42225) );
  XNOR U42167 ( .A(n42234), .B(n42235), .Z(n42174) );
  AND U42168 ( .A(n876), .B(n42236), .Z(n42235) );
  XNOR U42169 ( .A(n42237), .B(n42238), .Z(n42236) );
  XOR U42170 ( .A(n42239), .B(n42240), .Z(n42223) );
  AND U42171 ( .A(n42241), .B(n42242), .Z(n42240) );
  XNOR U42172 ( .A(n42239), .B(n42187), .Z(n42242) );
  XOR U42173 ( .A(n42243), .B(n42232), .Z(n42187) );
  XNOR U42174 ( .A(n42244), .B(n42227), .Z(n42232) );
  XOR U42175 ( .A(n42245), .B(n42246), .Z(n42227) );
  AND U42176 ( .A(n42247), .B(n42248), .Z(n42246) );
  XOR U42177 ( .A(n42249), .B(n42245), .Z(n42247) );
  XNOR U42178 ( .A(n42250), .B(n42251), .Z(n42244) );
  AND U42179 ( .A(n42252), .B(n42253), .Z(n42251) );
  XOR U42180 ( .A(n42250), .B(n42254), .Z(n42252) );
  XNOR U42181 ( .A(n42233), .B(n42230), .Z(n42243) );
  AND U42182 ( .A(n42255), .B(n42256), .Z(n42230) );
  XOR U42183 ( .A(n42257), .B(n42258), .Z(n42233) );
  AND U42184 ( .A(n42259), .B(n42260), .Z(n42258) );
  XOR U42185 ( .A(n42257), .B(n42261), .Z(n42259) );
  XNOR U42186 ( .A(n42184), .B(n42239), .Z(n42241) );
  XNOR U42187 ( .A(n42262), .B(n42263), .Z(n42184) );
  AND U42188 ( .A(n876), .B(n42264), .Z(n42263) );
  XNOR U42189 ( .A(n42265), .B(n42266), .Z(n42264) );
  XOR U42190 ( .A(n42267), .B(n42268), .Z(n42239) );
  AND U42191 ( .A(n42269), .B(n42270), .Z(n42268) );
  XNOR U42192 ( .A(n42267), .B(n42255), .Z(n42270) );
  IV U42193 ( .A(n42197), .Z(n42255) );
  XNOR U42194 ( .A(n42271), .B(n42248), .Z(n42197) );
  XNOR U42195 ( .A(n42272), .B(n42254), .Z(n42248) );
  XOR U42196 ( .A(n42273), .B(n42274), .Z(n42254) );
  AND U42197 ( .A(n42275), .B(n42276), .Z(n42274) );
  XOR U42198 ( .A(n42273), .B(n42277), .Z(n42275) );
  XNOR U42199 ( .A(n42253), .B(n42245), .Z(n42272) );
  XOR U42200 ( .A(n42278), .B(n42279), .Z(n42245) );
  AND U42201 ( .A(n42280), .B(n42281), .Z(n42279) );
  XNOR U42202 ( .A(n42282), .B(n42278), .Z(n42280) );
  XNOR U42203 ( .A(n42283), .B(n42250), .Z(n42253) );
  XOR U42204 ( .A(n42284), .B(n42285), .Z(n42250) );
  AND U42205 ( .A(n42286), .B(n42287), .Z(n42285) );
  XOR U42206 ( .A(n42284), .B(n42288), .Z(n42286) );
  XNOR U42207 ( .A(n42289), .B(n42290), .Z(n42283) );
  AND U42208 ( .A(n42291), .B(n42292), .Z(n42290) );
  XNOR U42209 ( .A(n42289), .B(n42293), .Z(n42291) );
  XNOR U42210 ( .A(n42249), .B(n42256), .Z(n42271) );
  AND U42211 ( .A(n42205), .B(n42294), .Z(n42256) );
  XOR U42212 ( .A(n42261), .B(n42260), .Z(n42249) );
  XNOR U42213 ( .A(n42295), .B(n42257), .Z(n42260) );
  XOR U42214 ( .A(n42296), .B(n42297), .Z(n42257) );
  AND U42215 ( .A(n42298), .B(n42299), .Z(n42297) );
  XOR U42216 ( .A(n42296), .B(n42300), .Z(n42298) );
  XNOR U42217 ( .A(n42301), .B(n42302), .Z(n42295) );
  AND U42218 ( .A(n42303), .B(n42304), .Z(n42302) );
  XOR U42219 ( .A(n42301), .B(n42305), .Z(n42303) );
  XOR U42220 ( .A(n42306), .B(n42307), .Z(n42261) );
  AND U42221 ( .A(n42308), .B(n42309), .Z(n42307) );
  XOR U42222 ( .A(n42306), .B(n42310), .Z(n42308) );
  XNOR U42223 ( .A(n42194), .B(n42267), .Z(n42269) );
  XNOR U42224 ( .A(n42311), .B(n42312), .Z(n42194) );
  AND U42225 ( .A(n876), .B(n42313), .Z(n42312) );
  XNOR U42226 ( .A(n42314), .B(n42315), .Z(n42313) );
  XOR U42227 ( .A(n42316), .B(n42317), .Z(n42267) );
  AND U42228 ( .A(n42318), .B(n42319), .Z(n42317) );
  XNOR U42229 ( .A(n42316), .B(n42205), .Z(n42319) );
  XOR U42230 ( .A(n42320), .B(n42281), .Z(n42205) );
  XNOR U42231 ( .A(n42321), .B(n42288), .Z(n42281) );
  XOR U42232 ( .A(n42277), .B(n42276), .Z(n42288) );
  XNOR U42233 ( .A(n42322), .B(n42273), .Z(n42276) );
  XOR U42234 ( .A(n42323), .B(n42324), .Z(n42273) );
  AND U42235 ( .A(n42325), .B(n42326), .Z(n42324) );
  XNOR U42236 ( .A(n42327), .B(n42328), .Z(n42325) );
  IV U42237 ( .A(n42323), .Z(n42327) );
  XNOR U42238 ( .A(n42329), .B(n42330), .Z(n42322) );
  NOR U42239 ( .A(n42331), .B(n42332), .Z(n42330) );
  XNOR U42240 ( .A(n42329), .B(n42333), .Z(n42331) );
  XOR U42241 ( .A(n42334), .B(n42335), .Z(n42277) );
  NOR U42242 ( .A(n42336), .B(n42337), .Z(n42335) );
  XNOR U42243 ( .A(n42334), .B(n42338), .Z(n42336) );
  XNOR U42244 ( .A(n42287), .B(n42278), .Z(n42321) );
  XOR U42245 ( .A(n42339), .B(n42340), .Z(n42278) );
  AND U42246 ( .A(n42341), .B(n42342), .Z(n42340) );
  XOR U42247 ( .A(n42339), .B(n42343), .Z(n42341) );
  XOR U42248 ( .A(n42344), .B(n42293), .Z(n42287) );
  XOR U42249 ( .A(n42345), .B(n42346), .Z(n42293) );
  NOR U42250 ( .A(n42347), .B(n42348), .Z(n42346) );
  XOR U42251 ( .A(n42345), .B(n42349), .Z(n42347) );
  XNOR U42252 ( .A(n42292), .B(n42284), .Z(n42344) );
  XOR U42253 ( .A(n42350), .B(n42351), .Z(n42284) );
  AND U42254 ( .A(n42352), .B(n42353), .Z(n42351) );
  XOR U42255 ( .A(n42350), .B(n42354), .Z(n42352) );
  XNOR U42256 ( .A(n42355), .B(n42289), .Z(n42292) );
  XOR U42257 ( .A(n42356), .B(n42357), .Z(n42289) );
  AND U42258 ( .A(n42358), .B(n42359), .Z(n42357) );
  XNOR U42259 ( .A(n42360), .B(n42361), .Z(n42358) );
  IV U42260 ( .A(n42356), .Z(n42360) );
  XNOR U42261 ( .A(n42362), .B(n42363), .Z(n42355) );
  NOR U42262 ( .A(n42364), .B(n42365), .Z(n42363) );
  XNOR U42263 ( .A(n42362), .B(n42366), .Z(n42364) );
  XOR U42264 ( .A(n42282), .B(n42294), .Z(n42320) );
  NOR U42265 ( .A(n42211), .B(n42367), .Z(n42294) );
  XNOR U42266 ( .A(n42300), .B(n42299), .Z(n42282) );
  XNOR U42267 ( .A(n42368), .B(n42305), .Z(n42299) );
  XNOR U42268 ( .A(n42369), .B(n42370), .Z(n42305) );
  NOR U42269 ( .A(n42371), .B(n42372), .Z(n42370) );
  XOR U42270 ( .A(n42369), .B(n42373), .Z(n42371) );
  XNOR U42271 ( .A(n42304), .B(n42296), .Z(n42368) );
  XOR U42272 ( .A(n42374), .B(n42375), .Z(n42296) );
  AND U42273 ( .A(n42376), .B(n42377), .Z(n42375) );
  XOR U42274 ( .A(n42374), .B(n42378), .Z(n42376) );
  XNOR U42275 ( .A(n42379), .B(n42301), .Z(n42304) );
  XOR U42276 ( .A(n42380), .B(n42381), .Z(n42301) );
  AND U42277 ( .A(n42382), .B(n42383), .Z(n42381) );
  XNOR U42278 ( .A(n42384), .B(n42385), .Z(n42382) );
  IV U42279 ( .A(n42380), .Z(n42384) );
  XNOR U42280 ( .A(n42386), .B(n42387), .Z(n42379) );
  NOR U42281 ( .A(n42388), .B(n42389), .Z(n42387) );
  XNOR U42282 ( .A(n42386), .B(n42390), .Z(n42388) );
  XOR U42283 ( .A(n42310), .B(n42309), .Z(n42300) );
  XNOR U42284 ( .A(n42391), .B(n42306), .Z(n42309) );
  XOR U42285 ( .A(n42392), .B(n42393), .Z(n42306) );
  AND U42286 ( .A(n42394), .B(n42395), .Z(n42393) );
  XNOR U42287 ( .A(n42396), .B(n42397), .Z(n42394) );
  IV U42288 ( .A(n42392), .Z(n42396) );
  XNOR U42289 ( .A(n42398), .B(n42399), .Z(n42391) );
  NOR U42290 ( .A(n42400), .B(n42401), .Z(n42399) );
  XNOR U42291 ( .A(n42398), .B(n42402), .Z(n42400) );
  XOR U42292 ( .A(n42403), .B(n42404), .Z(n42310) );
  NOR U42293 ( .A(n42405), .B(n42406), .Z(n42404) );
  XNOR U42294 ( .A(n42403), .B(n42407), .Z(n42405) );
  XNOR U42295 ( .A(n42202), .B(n42316), .Z(n42318) );
  XNOR U42296 ( .A(n42408), .B(n42409), .Z(n42202) );
  AND U42297 ( .A(n876), .B(n42410), .Z(n42409) );
  XNOR U42298 ( .A(n42411), .B(n42412), .Z(n42410) );
  AND U42299 ( .A(n42208), .B(n42211), .Z(n42316) );
  XOR U42300 ( .A(n42413), .B(n42367), .Z(n42211) );
  XNOR U42301 ( .A(p_input[1248]), .B(p_input[2048]), .Z(n42367) );
  XNOR U42302 ( .A(n42343), .B(n42342), .Z(n42413) );
  XNOR U42303 ( .A(n42414), .B(n42354), .Z(n42342) );
  XOR U42304 ( .A(n42328), .B(n42326), .Z(n42354) );
  XNOR U42305 ( .A(n42415), .B(n42333), .Z(n42326) );
  XOR U42306 ( .A(p_input[1272]), .B(p_input[2072]), .Z(n42333) );
  XOR U42307 ( .A(n42323), .B(n42332), .Z(n42415) );
  XOR U42308 ( .A(n42416), .B(n42329), .Z(n42332) );
  XOR U42309 ( .A(p_input[1270]), .B(p_input[2070]), .Z(n42329) );
  XOR U42310 ( .A(p_input[1271]), .B(n29410), .Z(n42416) );
  XOR U42311 ( .A(p_input[1266]), .B(p_input[2066]), .Z(n42323) );
  XNOR U42312 ( .A(n42338), .B(n42337), .Z(n42328) );
  XOR U42313 ( .A(n42417), .B(n42334), .Z(n42337) );
  XOR U42314 ( .A(p_input[1267]), .B(p_input[2067]), .Z(n42334) );
  XOR U42315 ( .A(p_input[1268]), .B(n29412), .Z(n42417) );
  XOR U42316 ( .A(p_input[1269]), .B(p_input[2069]), .Z(n42338) );
  XOR U42317 ( .A(n42353), .B(n42418), .Z(n42414) );
  IV U42318 ( .A(n42339), .Z(n42418) );
  XOR U42319 ( .A(p_input[1249]), .B(p_input[2049]), .Z(n42339) );
  XNOR U42320 ( .A(n42419), .B(n42361), .Z(n42353) );
  XNOR U42321 ( .A(n42349), .B(n42348), .Z(n42361) );
  XNOR U42322 ( .A(n42420), .B(n42345), .Z(n42348) );
  XNOR U42323 ( .A(p_input[1274]), .B(p_input[2074]), .Z(n42345) );
  XOR U42324 ( .A(p_input[1275]), .B(n29415), .Z(n42420) );
  XOR U42325 ( .A(p_input[1276]), .B(p_input[2076]), .Z(n42349) );
  XOR U42326 ( .A(n42359), .B(n42421), .Z(n42419) );
  IV U42327 ( .A(n42350), .Z(n42421) );
  XOR U42328 ( .A(p_input[1265]), .B(p_input[2065]), .Z(n42350) );
  XNOR U42329 ( .A(n42422), .B(n42366), .Z(n42359) );
  XNOR U42330 ( .A(p_input[1279]), .B(n29418), .Z(n42366) );
  XOR U42331 ( .A(n42356), .B(n42365), .Z(n42422) );
  XOR U42332 ( .A(n42423), .B(n42362), .Z(n42365) );
  XOR U42333 ( .A(p_input[1277]), .B(p_input[2077]), .Z(n42362) );
  XOR U42334 ( .A(p_input[1278]), .B(n29420), .Z(n42423) );
  XOR U42335 ( .A(p_input[1273]), .B(p_input[2073]), .Z(n42356) );
  XOR U42336 ( .A(n42378), .B(n42377), .Z(n42343) );
  XNOR U42337 ( .A(n42424), .B(n42385), .Z(n42377) );
  XNOR U42338 ( .A(n42373), .B(n42372), .Z(n42385) );
  XNOR U42339 ( .A(n42425), .B(n42369), .Z(n42372) );
  XNOR U42340 ( .A(p_input[1259]), .B(p_input[2059]), .Z(n42369) );
  XOR U42341 ( .A(p_input[1260]), .B(n28329), .Z(n42425) );
  XOR U42342 ( .A(p_input[1261]), .B(p_input[2061]), .Z(n42373) );
  XOR U42343 ( .A(n42383), .B(n42426), .Z(n42424) );
  IV U42344 ( .A(n42374), .Z(n42426) );
  XOR U42345 ( .A(p_input[1250]), .B(p_input[2050]), .Z(n42374) );
  XNOR U42346 ( .A(n42427), .B(n42390), .Z(n42383) );
  XNOR U42347 ( .A(p_input[1264]), .B(n28332), .Z(n42390) );
  XOR U42348 ( .A(n42380), .B(n42389), .Z(n42427) );
  XOR U42349 ( .A(n42428), .B(n42386), .Z(n42389) );
  XOR U42350 ( .A(p_input[1262]), .B(p_input[2062]), .Z(n42386) );
  XOR U42351 ( .A(p_input[1263]), .B(n28334), .Z(n42428) );
  XOR U42352 ( .A(p_input[1258]), .B(p_input[2058]), .Z(n42380) );
  XOR U42353 ( .A(n42397), .B(n42395), .Z(n42378) );
  XNOR U42354 ( .A(n42429), .B(n42402), .Z(n42395) );
  XOR U42355 ( .A(p_input[1257]), .B(p_input[2057]), .Z(n42402) );
  XOR U42356 ( .A(n42392), .B(n42401), .Z(n42429) );
  XOR U42357 ( .A(n42430), .B(n42398), .Z(n42401) );
  XOR U42358 ( .A(p_input[1255]), .B(p_input[2055]), .Z(n42398) );
  XOR U42359 ( .A(p_input[1256]), .B(n29427), .Z(n42430) );
  XOR U42360 ( .A(p_input[1251]), .B(p_input[2051]), .Z(n42392) );
  XNOR U42361 ( .A(n42407), .B(n42406), .Z(n42397) );
  XOR U42362 ( .A(n42431), .B(n42403), .Z(n42406) );
  XOR U42363 ( .A(p_input[1252]), .B(p_input[2052]), .Z(n42403) );
  XOR U42364 ( .A(p_input[1253]), .B(n29429), .Z(n42431) );
  XOR U42365 ( .A(p_input[1254]), .B(p_input[2054]), .Z(n42407) );
  XNOR U42366 ( .A(n42432), .B(n42433), .Z(n42208) );
  AND U42367 ( .A(n876), .B(n42434), .Z(n42433) );
  XNOR U42368 ( .A(n42435), .B(n42436), .Z(n876) );
  AND U42369 ( .A(n42437), .B(n42438), .Z(n42436) );
  XOR U42370 ( .A(n42222), .B(n42435), .Z(n42438) );
  XNOR U42371 ( .A(n42439), .B(n42435), .Z(n42437) );
  XOR U42372 ( .A(n42440), .B(n42441), .Z(n42435) );
  AND U42373 ( .A(n42442), .B(n42443), .Z(n42441) );
  XOR U42374 ( .A(n42237), .B(n42440), .Z(n42443) );
  XOR U42375 ( .A(n42440), .B(n42238), .Z(n42442) );
  XOR U42376 ( .A(n42444), .B(n42445), .Z(n42440) );
  AND U42377 ( .A(n42446), .B(n42447), .Z(n42445) );
  XOR U42378 ( .A(n42265), .B(n42444), .Z(n42447) );
  XOR U42379 ( .A(n42444), .B(n42266), .Z(n42446) );
  XOR U42380 ( .A(n42448), .B(n42449), .Z(n42444) );
  AND U42381 ( .A(n42450), .B(n42451), .Z(n42449) );
  XOR U42382 ( .A(n42314), .B(n42448), .Z(n42451) );
  XOR U42383 ( .A(n42448), .B(n42315), .Z(n42450) );
  XOR U42384 ( .A(n42452), .B(n42453), .Z(n42448) );
  AND U42385 ( .A(n42454), .B(n42455), .Z(n42453) );
  XOR U42386 ( .A(n42452), .B(n42411), .Z(n42455) );
  XNOR U42387 ( .A(n42456), .B(n42457), .Z(n42158) );
  AND U42388 ( .A(n880), .B(n42458), .Z(n42457) );
  XNOR U42389 ( .A(n42459), .B(n42460), .Z(n880) );
  AND U42390 ( .A(n42461), .B(n42462), .Z(n42460) );
  XOR U42391 ( .A(n42459), .B(n42168), .Z(n42462) );
  XNOR U42392 ( .A(n42459), .B(n42118), .Z(n42461) );
  XOR U42393 ( .A(n42463), .B(n42464), .Z(n42459) );
  AND U42394 ( .A(n42465), .B(n42466), .Z(n42464) );
  XNOR U42395 ( .A(n42178), .B(n42463), .Z(n42466) );
  XOR U42396 ( .A(n42463), .B(n42128), .Z(n42465) );
  XOR U42397 ( .A(n42467), .B(n42468), .Z(n42463) );
  AND U42398 ( .A(n42469), .B(n42470), .Z(n42468) );
  XNOR U42399 ( .A(n42188), .B(n42467), .Z(n42470) );
  XOR U42400 ( .A(n42467), .B(n42137), .Z(n42469) );
  XOR U42401 ( .A(n42471), .B(n42472), .Z(n42467) );
  AND U42402 ( .A(n42473), .B(n42474), .Z(n42472) );
  XOR U42403 ( .A(n42471), .B(n42145), .Z(n42473) );
  XOR U42404 ( .A(n42475), .B(n42476), .Z(n42109) );
  AND U42405 ( .A(n884), .B(n42458), .Z(n42476) );
  XNOR U42406 ( .A(n42456), .B(n42475), .Z(n42458) );
  XNOR U42407 ( .A(n42477), .B(n42478), .Z(n884) );
  AND U42408 ( .A(n42479), .B(n42480), .Z(n42478) );
  XNOR U42409 ( .A(n42481), .B(n42477), .Z(n42480) );
  IV U42410 ( .A(n42168), .Z(n42481) );
  XOR U42411 ( .A(n42439), .B(n42482), .Z(n42168) );
  AND U42412 ( .A(n887), .B(n42483), .Z(n42482) );
  XOR U42413 ( .A(n42221), .B(n42218), .Z(n42483) );
  IV U42414 ( .A(n42439), .Z(n42221) );
  XNOR U42415 ( .A(n42118), .B(n42477), .Z(n42479) );
  XOR U42416 ( .A(n42484), .B(n42485), .Z(n42118) );
  AND U42417 ( .A(n903), .B(n42486), .Z(n42485) );
  XOR U42418 ( .A(n42487), .B(n42488), .Z(n42477) );
  AND U42419 ( .A(n42489), .B(n42490), .Z(n42488) );
  XNOR U42420 ( .A(n42487), .B(n42178), .Z(n42490) );
  XOR U42421 ( .A(n42238), .B(n42491), .Z(n42178) );
  AND U42422 ( .A(n887), .B(n42492), .Z(n42491) );
  XOR U42423 ( .A(n42234), .B(n42238), .Z(n42492) );
  XNOR U42424 ( .A(n42493), .B(n42487), .Z(n42489) );
  IV U42425 ( .A(n42128), .Z(n42493) );
  XOR U42426 ( .A(n42494), .B(n42495), .Z(n42128) );
  AND U42427 ( .A(n903), .B(n42496), .Z(n42495) );
  XOR U42428 ( .A(n42497), .B(n42498), .Z(n42487) );
  AND U42429 ( .A(n42499), .B(n42500), .Z(n42498) );
  XNOR U42430 ( .A(n42497), .B(n42188), .Z(n42500) );
  XOR U42431 ( .A(n42266), .B(n42501), .Z(n42188) );
  AND U42432 ( .A(n887), .B(n42502), .Z(n42501) );
  XOR U42433 ( .A(n42262), .B(n42266), .Z(n42502) );
  XOR U42434 ( .A(n42137), .B(n42497), .Z(n42499) );
  XOR U42435 ( .A(n42503), .B(n42504), .Z(n42137) );
  AND U42436 ( .A(n903), .B(n42505), .Z(n42504) );
  XOR U42437 ( .A(n42471), .B(n42506), .Z(n42497) );
  AND U42438 ( .A(n42507), .B(n42474), .Z(n42506) );
  XNOR U42439 ( .A(n42198), .B(n42471), .Z(n42474) );
  XOR U42440 ( .A(n42315), .B(n42508), .Z(n42198) );
  AND U42441 ( .A(n887), .B(n42509), .Z(n42508) );
  XOR U42442 ( .A(n42311), .B(n42315), .Z(n42509) );
  XNOR U42443 ( .A(n42510), .B(n42471), .Z(n42507) );
  IV U42444 ( .A(n42145), .Z(n42510) );
  XOR U42445 ( .A(n42511), .B(n42512), .Z(n42145) );
  AND U42446 ( .A(n903), .B(n42513), .Z(n42512) );
  XOR U42447 ( .A(n42514), .B(n42515), .Z(n42471) );
  AND U42448 ( .A(n42516), .B(n42517), .Z(n42515) );
  XNOR U42449 ( .A(n42514), .B(n42206), .Z(n42517) );
  XOR U42450 ( .A(n42412), .B(n42518), .Z(n42206) );
  AND U42451 ( .A(n887), .B(n42519), .Z(n42518) );
  XOR U42452 ( .A(n42408), .B(n42412), .Z(n42519) );
  XNOR U42453 ( .A(n42520), .B(n42514), .Z(n42516) );
  IV U42454 ( .A(n42155), .Z(n42520) );
  XOR U42455 ( .A(n42521), .B(n42522), .Z(n42155) );
  AND U42456 ( .A(n903), .B(n42523), .Z(n42522) );
  AND U42457 ( .A(n42475), .B(n42456), .Z(n42514) );
  XNOR U42458 ( .A(n42524), .B(n42525), .Z(n42456) );
  AND U42459 ( .A(n887), .B(n42434), .Z(n42525) );
  XNOR U42460 ( .A(n42432), .B(n42524), .Z(n42434) );
  XNOR U42461 ( .A(n42526), .B(n42527), .Z(n887) );
  AND U42462 ( .A(n42528), .B(n42529), .Z(n42527) );
  XNOR U42463 ( .A(n42526), .B(n42218), .Z(n42529) );
  IV U42464 ( .A(n42222), .Z(n42218) );
  XOR U42465 ( .A(n42530), .B(n42531), .Z(n42222) );
  AND U42466 ( .A(n891), .B(n42532), .Z(n42531) );
  XOR U42467 ( .A(n42533), .B(n42530), .Z(n42532) );
  XNOR U42468 ( .A(n42526), .B(n42439), .Z(n42528) );
  XOR U42469 ( .A(n42534), .B(n42535), .Z(n42439) );
  AND U42470 ( .A(n899), .B(n42486), .Z(n42535) );
  XOR U42471 ( .A(n42484), .B(n42534), .Z(n42486) );
  XOR U42472 ( .A(n42536), .B(n42537), .Z(n42526) );
  AND U42473 ( .A(n42538), .B(n42539), .Z(n42537) );
  XNOR U42474 ( .A(n42536), .B(n42234), .Z(n42539) );
  IV U42475 ( .A(n42237), .Z(n42234) );
  XOR U42476 ( .A(n42540), .B(n42541), .Z(n42237) );
  AND U42477 ( .A(n891), .B(n42542), .Z(n42541) );
  XOR U42478 ( .A(n42543), .B(n42540), .Z(n42542) );
  XOR U42479 ( .A(n42238), .B(n42536), .Z(n42538) );
  XOR U42480 ( .A(n42544), .B(n42545), .Z(n42238) );
  AND U42481 ( .A(n899), .B(n42496), .Z(n42545) );
  XOR U42482 ( .A(n42544), .B(n42494), .Z(n42496) );
  XOR U42483 ( .A(n42546), .B(n42547), .Z(n42536) );
  AND U42484 ( .A(n42548), .B(n42549), .Z(n42547) );
  XNOR U42485 ( .A(n42546), .B(n42262), .Z(n42549) );
  IV U42486 ( .A(n42265), .Z(n42262) );
  XOR U42487 ( .A(n42550), .B(n42551), .Z(n42265) );
  AND U42488 ( .A(n891), .B(n42552), .Z(n42551) );
  XNOR U42489 ( .A(n42553), .B(n42550), .Z(n42552) );
  XOR U42490 ( .A(n42266), .B(n42546), .Z(n42548) );
  XOR U42491 ( .A(n42554), .B(n42555), .Z(n42266) );
  AND U42492 ( .A(n899), .B(n42505), .Z(n42555) );
  XOR U42493 ( .A(n42554), .B(n42503), .Z(n42505) );
  XOR U42494 ( .A(n42556), .B(n42557), .Z(n42546) );
  AND U42495 ( .A(n42558), .B(n42559), .Z(n42557) );
  XNOR U42496 ( .A(n42556), .B(n42311), .Z(n42559) );
  IV U42497 ( .A(n42314), .Z(n42311) );
  XOR U42498 ( .A(n42560), .B(n42561), .Z(n42314) );
  AND U42499 ( .A(n891), .B(n42562), .Z(n42561) );
  XOR U42500 ( .A(n42563), .B(n42560), .Z(n42562) );
  XOR U42501 ( .A(n42315), .B(n42556), .Z(n42558) );
  XOR U42502 ( .A(n42564), .B(n42565), .Z(n42315) );
  AND U42503 ( .A(n899), .B(n42513), .Z(n42565) );
  XOR U42504 ( .A(n42564), .B(n42511), .Z(n42513) );
  XOR U42505 ( .A(n42452), .B(n42566), .Z(n42556) );
  AND U42506 ( .A(n42454), .B(n42567), .Z(n42566) );
  XNOR U42507 ( .A(n42452), .B(n42408), .Z(n42567) );
  IV U42508 ( .A(n42411), .Z(n42408) );
  XOR U42509 ( .A(n42568), .B(n42569), .Z(n42411) );
  AND U42510 ( .A(n891), .B(n42570), .Z(n42569) );
  XNOR U42511 ( .A(n42571), .B(n42568), .Z(n42570) );
  XOR U42512 ( .A(n42412), .B(n42452), .Z(n42454) );
  XOR U42513 ( .A(n42572), .B(n42573), .Z(n42412) );
  AND U42514 ( .A(n899), .B(n42523), .Z(n42573) );
  XOR U42515 ( .A(n42572), .B(n42521), .Z(n42523) );
  AND U42516 ( .A(n42524), .B(n42432), .Z(n42452) );
  XNOR U42517 ( .A(n42574), .B(n42575), .Z(n42432) );
  AND U42518 ( .A(n891), .B(n42576), .Z(n42575) );
  XNOR U42519 ( .A(n42577), .B(n42574), .Z(n42576) );
  XNOR U42520 ( .A(n42578), .B(n42579), .Z(n891) );
  AND U42521 ( .A(n42580), .B(n42581), .Z(n42579) );
  XOR U42522 ( .A(n42533), .B(n42578), .Z(n42581) );
  AND U42523 ( .A(n42582), .B(n42583), .Z(n42533) );
  XNOR U42524 ( .A(n42530), .B(n42578), .Z(n42580) );
  XNOR U42525 ( .A(n42584), .B(n42585), .Z(n42530) );
  AND U42526 ( .A(n895), .B(n42586), .Z(n42585) );
  XNOR U42527 ( .A(n42587), .B(n42588), .Z(n42586) );
  XOR U42528 ( .A(n42589), .B(n42590), .Z(n42578) );
  AND U42529 ( .A(n42591), .B(n42592), .Z(n42590) );
  XNOR U42530 ( .A(n42589), .B(n42582), .Z(n42592) );
  IV U42531 ( .A(n42543), .Z(n42582) );
  XOR U42532 ( .A(n42593), .B(n42594), .Z(n42543) );
  XOR U42533 ( .A(n42595), .B(n42583), .Z(n42594) );
  AND U42534 ( .A(n42553), .B(n42596), .Z(n42583) );
  AND U42535 ( .A(n42597), .B(n42598), .Z(n42595) );
  XOR U42536 ( .A(n42599), .B(n42593), .Z(n42597) );
  XNOR U42537 ( .A(n42540), .B(n42589), .Z(n42591) );
  XNOR U42538 ( .A(n42600), .B(n42601), .Z(n42540) );
  AND U42539 ( .A(n895), .B(n42602), .Z(n42601) );
  XNOR U42540 ( .A(n42603), .B(n42604), .Z(n42602) );
  XOR U42541 ( .A(n42605), .B(n42606), .Z(n42589) );
  AND U42542 ( .A(n42607), .B(n42608), .Z(n42606) );
  XNOR U42543 ( .A(n42605), .B(n42553), .Z(n42608) );
  XOR U42544 ( .A(n42609), .B(n42598), .Z(n42553) );
  XNOR U42545 ( .A(n42610), .B(n42593), .Z(n42598) );
  XOR U42546 ( .A(n42611), .B(n42612), .Z(n42593) );
  AND U42547 ( .A(n42613), .B(n42614), .Z(n42612) );
  XOR U42548 ( .A(n42615), .B(n42611), .Z(n42613) );
  XNOR U42549 ( .A(n42616), .B(n42617), .Z(n42610) );
  AND U42550 ( .A(n42618), .B(n42619), .Z(n42617) );
  XOR U42551 ( .A(n42616), .B(n42620), .Z(n42618) );
  XNOR U42552 ( .A(n42599), .B(n42596), .Z(n42609) );
  AND U42553 ( .A(n42621), .B(n42622), .Z(n42596) );
  XOR U42554 ( .A(n42623), .B(n42624), .Z(n42599) );
  AND U42555 ( .A(n42625), .B(n42626), .Z(n42624) );
  XOR U42556 ( .A(n42623), .B(n42627), .Z(n42625) );
  XNOR U42557 ( .A(n42550), .B(n42605), .Z(n42607) );
  XNOR U42558 ( .A(n42628), .B(n42629), .Z(n42550) );
  AND U42559 ( .A(n895), .B(n42630), .Z(n42629) );
  XNOR U42560 ( .A(n42631), .B(n42632), .Z(n42630) );
  XOR U42561 ( .A(n42633), .B(n42634), .Z(n42605) );
  AND U42562 ( .A(n42635), .B(n42636), .Z(n42634) );
  XNOR U42563 ( .A(n42633), .B(n42621), .Z(n42636) );
  IV U42564 ( .A(n42563), .Z(n42621) );
  XNOR U42565 ( .A(n42637), .B(n42614), .Z(n42563) );
  XNOR U42566 ( .A(n42638), .B(n42620), .Z(n42614) );
  XOR U42567 ( .A(n42639), .B(n42640), .Z(n42620) );
  AND U42568 ( .A(n42641), .B(n42642), .Z(n42640) );
  XOR U42569 ( .A(n42639), .B(n42643), .Z(n42641) );
  XNOR U42570 ( .A(n42619), .B(n42611), .Z(n42638) );
  XOR U42571 ( .A(n42644), .B(n42645), .Z(n42611) );
  AND U42572 ( .A(n42646), .B(n42647), .Z(n42645) );
  XNOR U42573 ( .A(n42648), .B(n42644), .Z(n42646) );
  XNOR U42574 ( .A(n42649), .B(n42616), .Z(n42619) );
  XOR U42575 ( .A(n42650), .B(n42651), .Z(n42616) );
  AND U42576 ( .A(n42652), .B(n42653), .Z(n42651) );
  XOR U42577 ( .A(n42650), .B(n42654), .Z(n42652) );
  XNOR U42578 ( .A(n42655), .B(n42656), .Z(n42649) );
  AND U42579 ( .A(n42657), .B(n42658), .Z(n42656) );
  XNOR U42580 ( .A(n42655), .B(n42659), .Z(n42657) );
  XNOR U42581 ( .A(n42615), .B(n42622), .Z(n42637) );
  AND U42582 ( .A(n42571), .B(n42660), .Z(n42622) );
  XOR U42583 ( .A(n42627), .B(n42626), .Z(n42615) );
  XNOR U42584 ( .A(n42661), .B(n42623), .Z(n42626) );
  XOR U42585 ( .A(n42662), .B(n42663), .Z(n42623) );
  AND U42586 ( .A(n42664), .B(n42665), .Z(n42663) );
  XOR U42587 ( .A(n42662), .B(n42666), .Z(n42664) );
  XNOR U42588 ( .A(n42667), .B(n42668), .Z(n42661) );
  AND U42589 ( .A(n42669), .B(n42670), .Z(n42668) );
  XOR U42590 ( .A(n42667), .B(n42671), .Z(n42669) );
  XOR U42591 ( .A(n42672), .B(n42673), .Z(n42627) );
  AND U42592 ( .A(n42674), .B(n42675), .Z(n42673) );
  XOR U42593 ( .A(n42672), .B(n42676), .Z(n42674) );
  XNOR U42594 ( .A(n42560), .B(n42633), .Z(n42635) );
  XNOR U42595 ( .A(n42677), .B(n42678), .Z(n42560) );
  AND U42596 ( .A(n895), .B(n42679), .Z(n42678) );
  XNOR U42597 ( .A(n42680), .B(n42681), .Z(n42679) );
  XOR U42598 ( .A(n42682), .B(n42683), .Z(n42633) );
  AND U42599 ( .A(n42684), .B(n42685), .Z(n42683) );
  XNOR U42600 ( .A(n42682), .B(n42571), .Z(n42685) );
  XOR U42601 ( .A(n42686), .B(n42647), .Z(n42571) );
  XNOR U42602 ( .A(n42687), .B(n42654), .Z(n42647) );
  XOR U42603 ( .A(n42643), .B(n42642), .Z(n42654) );
  XNOR U42604 ( .A(n42688), .B(n42639), .Z(n42642) );
  XOR U42605 ( .A(n42689), .B(n42690), .Z(n42639) );
  AND U42606 ( .A(n42691), .B(n42692), .Z(n42690) );
  XNOR U42607 ( .A(n42693), .B(n42694), .Z(n42691) );
  IV U42608 ( .A(n42689), .Z(n42693) );
  XNOR U42609 ( .A(n42695), .B(n42696), .Z(n42688) );
  NOR U42610 ( .A(n42697), .B(n42698), .Z(n42696) );
  XNOR U42611 ( .A(n42695), .B(n42699), .Z(n42697) );
  XOR U42612 ( .A(n42700), .B(n42701), .Z(n42643) );
  NOR U42613 ( .A(n42702), .B(n42703), .Z(n42701) );
  XNOR U42614 ( .A(n42700), .B(n42704), .Z(n42702) );
  XNOR U42615 ( .A(n42653), .B(n42644), .Z(n42687) );
  XOR U42616 ( .A(n42705), .B(n42706), .Z(n42644) );
  AND U42617 ( .A(n42707), .B(n42708), .Z(n42706) );
  XOR U42618 ( .A(n42705), .B(n42709), .Z(n42707) );
  XOR U42619 ( .A(n42710), .B(n42659), .Z(n42653) );
  XOR U42620 ( .A(n42711), .B(n42712), .Z(n42659) );
  NOR U42621 ( .A(n42713), .B(n42714), .Z(n42712) );
  XOR U42622 ( .A(n42711), .B(n42715), .Z(n42713) );
  XNOR U42623 ( .A(n42658), .B(n42650), .Z(n42710) );
  XOR U42624 ( .A(n42716), .B(n42717), .Z(n42650) );
  AND U42625 ( .A(n42718), .B(n42719), .Z(n42717) );
  XOR U42626 ( .A(n42716), .B(n42720), .Z(n42718) );
  XNOR U42627 ( .A(n42721), .B(n42655), .Z(n42658) );
  XOR U42628 ( .A(n42722), .B(n42723), .Z(n42655) );
  AND U42629 ( .A(n42724), .B(n42725), .Z(n42723) );
  XNOR U42630 ( .A(n42726), .B(n42727), .Z(n42724) );
  IV U42631 ( .A(n42722), .Z(n42726) );
  XNOR U42632 ( .A(n42728), .B(n42729), .Z(n42721) );
  NOR U42633 ( .A(n42730), .B(n42731), .Z(n42729) );
  XNOR U42634 ( .A(n42728), .B(n42732), .Z(n42730) );
  XOR U42635 ( .A(n42648), .B(n42660), .Z(n42686) );
  NOR U42636 ( .A(n42577), .B(n42733), .Z(n42660) );
  XNOR U42637 ( .A(n42666), .B(n42665), .Z(n42648) );
  XNOR U42638 ( .A(n42734), .B(n42671), .Z(n42665) );
  XNOR U42639 ( .A(n42735), .B(n42736), .Z(n42671) );
  NOR U42640 ( .A(n42737), .B(n42738), .Z(n42736) );
  XOR U42641 ( .A(n42735), .B(n42739), .Z(n42737) );
  XNOR U42642 ( .A(n42670), .B(n42662), .Z(n42734) );
  XOR U42643 ( .A(n42740), .B(n42741), .Z(n42662) );
  AND U42644 ( .A(n42742), .B(n42743), .Z(n42741) );
  XOR U42645 ( .A(n42740), .B(n42744), .Z(n42742) );
  XNOR U42646 ( .A(n42745), .B(n42667), .Z(n42670) );
  XOR U42647 ( .A(n42746), .B(n42747), .Z(n42667) );
  AND U42648 ( .A(n42748), .B(n42749), .Z(n42747) );
  XNOR U42649 ( .A(n42750), .B(n42751), .Z(n42748) );
  IV U42650 ( .A(n42746), .Z(n42750) );
  XNOR U42651 ( .A(n42752), .B(n42753), .Z(n42745) );
  NOR U42652 ( .A(n42754), .B(n42755), .Z(n42753) );
  XNOR U42653 ( .A(n42752), .B(n42756), .Z(n42754) );
  XOR U42654 ( .A(n42676), .B(n42675), .Z(n42666) );
  XNOR U42655 ( .A(n42757), .B(n42672), .Z(n42675) );
  XOR U42656 ( .A(n42758), .B(n42759), .Z(n42672) );
  AND U42657 ( .A(n42760), .B(n42761), .Z(n42759) );
  XNOR U42658 ( .A(n42762), .B(n42763), .Z(n42760) );
  IV U42659 ( .A(n42758), .Z(n42762) );
  XNOR U42660 ( .A(n42764), .B(n42765), .Z(n42757) );
  NOR U42661 ( .A(n42766), .B(n42767), .Z(n42765) );
  XNOR U42662 ( .A(n42764), .B(n42768), .Z(n42766) );
  XOR U42663 ( .A(n42769), .B(n42770), .Z(n42676) );
  NOR U42664 ( .A(n42771), .B(n42772), .Z(n42770) );
  XNOR U42665 ( .A(n42769), .B(n42773), .Z(n42771) );
  XNOR U42666 ( .A(n42568), .B(n42682), .Z(n42684) );
  XNOR U42667 ( .A(n42774), .B(n42775), .Z(n42568) );
  AND U42668 ( .A(n895), .B(n42776), .Z(n42775) );
  XNOR U42669 ( .A(n42777), .B(n42778), .Z(n42776) );
  AND U42670 ( .A(n42574), .B(n42577), .Z(n42682) );
  XOR U42671 ( .A(n42779), .B(n42733), .Z(n42577) );
  XNOR U42672 ( .A(p_input[1280]), .B(p_input[2048]), .Z(n42733) );
  XNOR U42673 ( .A(n42709), .B(n42708), .Z(n42779) );
  XNOR U42674 ( .A(n42780), .B(n42720), .Z(n42708) );
  XOR U42675 ( .A(n42694), .B(n42692), .Z(n42720) );
  XNOR U42676 ( .A(n42781), .B(n42699), .Z(n42692) );
  XOR U42677 ( .A(p_input[1304]), .B(p_input[2072]), .Z(n42699) );
  XOR U42678 ( .A(n42689), .B(n42698), .Z(n42781) );
  XOR U42679 ( .A(n42782), .B(n42695), .Z(n42698) );
  XOR U42680 ( .A(p_input[1302]), .B(p_input[2070]), .Z(n42695) );
  XOR U42681 ( .A(p_input[1303]), .B(n29410), .Z(n42782) );
  XOR U42682 ( .A(p_input[1298]), .B(p_input[2066]), .Z(n42689) );
  XNOR U42683 ( .A(n42704), .B(n42703), .Z(n42694) );
  XOR U42684 ( .A(n42783), .B(n42700), .Z(n42703) );
  XOR U42685 ( .A(p_input[1299]), .B(p_input[2067]), .Z(n42700) );
  XOR U42686 ( .A(p_input[1300]), .B(n29412), .Z(n42783) );
  XOR U42687 ( .A(p_input[1301]), .B(p_input[2069]), .Z(n42704) );
  XOR U42688 ( .A(n42719), .B(n42784), .Z(n42780) );
  IV U42689 ( .A(n42705), .Z(n42784) );
  XOR U42690 ( .A(p_input[1281]), .B(p_input[2049]), .Z(n42705) );
  XNOR U42691 ( .A(n42785), .B(n42727), .Z(n42719) );
  XNOR U42692 ( .A(n42715), .B(n42714), .Z(n42727) );
  XNOR U42693 ( .A(n42786), .B(n42711), .Z(n42714) );
  XNOR U42694 ( .A(p_input[1306]), .B(p_input[2074]), .Z(n42711) );
  XOR U42695 ( .A(p_input[1307]), .B(n29415), .Z(n42786) );
  XOR U42696 ( .A(p_input[1308]), .B(p_input[2076]), .Z(n42715) );
  XOR U42697 ( .A(n42725), .B(n42787), .Z(n42785) );
  IV U42698 ( .A(n42716), .Z(n42787) );
  XOR U42699 ( .A(p_input[1297]), .B(p_input[2065]), .Z(n42716) );
  XNOR U42700 ( .A(n42788), .B(n42732), .Z(n42725) );
  XNOR U42701 ( .A(p_input[1311]), .B(n29418), .Z(n42732) );
  XOR U42702 ( .A(n42722), .B(n42731), .Z(n42788) );
  XOR U42703 ( .A(n42789), .B(n42728), .Z(n42731) );
  XOR U42704 ( .A(p_input[1309]), .B(p_input[2077]), .Z(n42728) );
  XOR U42705 ( .A(p_input[1310]), .B(n29420), .Z(n42789) );
  XOR U42706 ( .A(p_input[1305]), .B(p_input[2073]), .Z(n42722) );
  XOR U42707 ( .A(n42744), .B(n42743), .Z(n42709) );
  XNOR U42708 ( .A(n42790), .B(n42751), .Z(n42743) );
  XNOR U42709 ( .A(n42739), .B(n42738), .Z(n42751) );
  XNOR U42710 ( .A(n42791), .B(n42735), .Z(n42738) );
  XNOR U42711 ( .A(p_input[1291]), .B(p_input[2059]), .Z(n42735) );
  XOR U42712 ( .A(p_input[1292]), .B(n28329), .Z(n42791) );
  XOR U42713 ( .A(p_input[1293]), .B(p_input[2061]), .Z(n42739) );
  XOR U42714 ( .A(n42749), .B(n42792), .Z(n42790) );
  IV U42715 ( .A(n42740), .Z(n42792) );
  XOR U42716 ( .A(p_input[1282]), .B(p_input[2050]), .Z(n42740) );
  XNOR U42717 ( .A(n42793), .B(n42756), .Z(n42749) );
  XNOR U42718 ( .A(p_input[1296]), .B(n28332), .Z(n42756) );
  XOR U42719 ( .A(n42746), .B(n42755), .Z(n42793) );
  XOR U42720 ( .A(n42794), .B(n42752), .Z(n42755) );
  XOR U42721 ( .A(p_input[1294]), .B(p_input[2062]), .Z(n42752) );
  XOR U42722 ( .A(p_input[1295]), .B(n28334), .Z(n42794) );
  XOR U42723 ( .A(p_input[1290]), .B(p_input[2058]), .Z(n42746) );
  XOR U42724 ( .A(n42763), .B(n42761), .Z(n42744) );
  XNOR U42725 ( .A(n42795), .B(n42768), .Z(n42761) );
  XOR U42726 ( .A(p_input[1289]), .B(p_input[2057]), .Z(n42768) );
  XOR U42727 ( .A(n42758), .B(n42767), .Z(n42795) );
  XOR U42728 ( .A(n42796), .B(n42764), .Z(n42767) );
  XOR U42729 ( .A(p_input[1287]), .B(p_input[2055]), .Z(n42764) );
  XOR U42730 ( .A(p_input[1288]), .B(n29427), .Z(n42796) );
  XOR U42731 ( .A(p_input[1283]), .B(p_input[2051]), .Z(n42758) );
  XNOR U42732 ( .A(n42773), .B(n42772), .Z(n42763) );
  XOR U42733 ( .A(n42797), .B(n42769), .Z(n42772) );
  XOR U42734 ( .A(p_input[1284]), .B(p_input[2052]), .Z(n42769) );
  XOR U42735 ( .A(p_input[1285]), .B(n29429), .Z(n42797) );
  XOR U42736 ( .A(p_input[1286]), .B(p_input[2054]), .Z(n42773) );
  XNOR U42737 ( .A(n42798), .B(n42799), .Z(n42574) );
  AND U42738 ( .A(n895), .B(n42800), .Z(n42799) );
  XNOR U42739 ( .A(n42801), .B(n42802), .Z(n895) );
  AND U42740 ( .A(n42803), .B(n42804), .Z(n42802) );
  XOR U42741 ( .A(n42588), .B(n42801), .Z(n42804) );
  XNOR U42742 ( .A(n42805), .B(n42801), .Z(n42803) );
  XOR U42743 ( .A(n42806), .B(n42807), .Z(n42801) );
  AND U42744 ( .A(n42808), .B(n42809), .Z(n42807) );
  XOR U42745 ( .A(n42603), .B(n42806), .Z(n42809) );
  XOR U42746 ( .A(n42806), .B(n42604), .Z(n42808) );
  XOR U42747 ( .A(n42810), .B(n42811), .Z(n42806) );
  AND U42748 ( .A(n42812), .B(n42813), .Z(n42811) );
  XOR U42749 ( .A(n42631), .B(n42810), .Z(n42813) );
  XOR U42750 ( .A(n42810), .B(n42632), .Z(n42812) );
  XOR U42751 ( .A(n42814), .B(n42815), .Z(n42810) );
  AND U42752 ( .A(n42816), .B(n42817), .Z(n42815) );
  XOR U42753 ( .A(n42680), .B(n42814), .Z(n42817) );
  XOR U42754 ( .A(n42814), .B(n42681), .Z(n42816) );
  XOR U42755 ( .A(n42818), .B(n42819), .Z(n42814) );
  AND U42756 ( .A(n42820), .B(n42821), .Z(n42819) );
  XOR U42757 ( .A(n42818), .B(n42777), .Z(n42821) );
  XNOR U42758 ( .A(n42822), .B(n42823), .Z(n42524) );
  AND U42759 ( .A(n899), .B(n42824), .Z(n42823) );
  XNOR U42760 ( .A(n42825), .B(n42826), .Z(n899) );
  AND U42761 ( .A(n42827), .B(n42828), .Z(n42826) );
  XOR U42762 ( .A(n42825), .B(n42534), .Z(n42828) );
  XNOR U42763 ( .A(n42825), .B(n42484), .Z(n42827) );
  XOR U42764 ( .A(n42829), .B(n42830), .Z(n42825) );
  AND U42765 ( .A(n42831), .B(n42832), .Z(n42830) );
  XNOR U42766 ( .A(n42544), .B(n42829), .Z(n42832) );
  XOR U42767 ( .A(n42829), .B(n42494), .Z(n42831) );
  XOR U42768 ( .A(n42833), .B(n42834), .Z(n42829) );
  AND U42769 ( .A(n42835), .B(n42836), .Z(n42834) );
  XNOR U42770 ( .A(n42554), .B(n42833), .Z(n42836) );
  XOR U42771 ( .A(n42833), .B(n42503), .Z(n42835) );
  XOR U42772 ( .A(n42837), .B(n42838), .Z(n42833) );
  AND U42773 ( .A(n42839), .B(n42840), .Z(n42838) );
  XOR U42774 ( .A(n42837), .B(n42511), .Z(n42839) );
  XOR U42775 ( .A(n42841), .B(n42842), .Z(n42475) );
  AND U42776 ( .A(n903), .B(n42824), .Z(n42842) );
  XNOR U42777 ( .A(n42822), .B(n42841), .Z(n42824) );
  XNOR U42778 ( .A(n42843), .B(n42844), .Z(n903) );
  AND U42779 ( .A(n42845), .B(n42846), .Z(n42844) );
  XNOR U42780 ( .A(n42847), .B(n42843), .Z(n42846) );
  IV U42781 ( .A(n42534), .Z(n42847) );
  XOR U42782 ( .A(n42805), .B(n42848), .Z(n42534) );
  AND U42783 ( .A(n906), .B(n42849), .Z(n42848) );
  XOR U42784 ( .A(n42587), .B(n42584), .Z(n42849) );
  IV U42785 ( .A(n42805), .Z(n42587) );
  XNOR U42786 ( .A(n42484), .B(n42843), .Z(n42845) );
  XOR U42787 ( .A(n42850), .B(n42851), .Z(n42484) );
  AND U42788 ( .A(n922), .B(n42852), .Z(n42851) );
  XOR U42789 ( .A(n42853), .B(n42854), .Z(n42843) );
  AND U42790 ( .A(n42855), .B(n42856), .Z(n42854) );
  XNOR U42791 ( .A(n42853), .B(n42544), .Z(n42856) );
  XOR U42792 ( .A(n42604), .B(n42857), .Z(n42544) );
  AND U42793 ( .A(n906), .B(n42858), .Z(n42857) );
  XOR U42794 ( .A(n42600), .B(n42604), .Z(n42858) );
  XNOR U42795 ( .A(n42859), .B(n42853), .Z(n42855) );
  IV U42796 ( .A(n42494), .Z(n42859) );
  XOR U42797 ( .A(n42860), .B(n42861), .Z(n42494) );
  AND U42798 ( .A(n922), .B(n42862), .Z(n42861) );
  XOR U42799 ( .A(n42863), .B(n42864), .Z(n42853) );
  AND U42800 ( .A(n42865), .B(n42866), .Z(n42864) );
  XNOR U42801 ( .A(n42863), .B(n42554), .Z(n42866) );
  XOR U42802 ( .A(n42632), .B(n42867), .Z(n42554) );
  AND U42803 ( .A(n906), .B(n42868), .Z(n42867) );
  XOR U42804 ( .A(n42628), .B(n42632), .Z(n42868) );
  XOR U42805 ( .A(n42503), .B(n42863), .Z(n42865) );
  XOR U42806 ( .A(n42869), .B(n42870), .Z(n42503) );
  AND U42807 ( .A(n922), .B(n42871), .Z(n42870) );
  XOR U42808 ( .A(n42837), .B(n42872), .Z(n42863) );
  AND U42809 ( .A(n42873), .B(n42840), .Z(n42872) );
  XNOR U42810 ( .A(n42564), .B(n42837), .Z(n42840) );
  XOR U42811 ( .A(n42681), .B(n42874), .Z(n42564) );
  AND U42812 ( .A(n906), .B(n42875), .Z(n42874) );
  XOR U42813 ( .A(n42677), .B(n42681), .Z(n42875) );
  XNOR U42814 ( .A(n42876), .B(n42837), .Z(n42873) );
  IV U42815 ( .A(n42511), .Z(n42876) );
  XOR U42816 ( .A(n42877), .B(n42878), .Z(n42511) );
  AND U42817 ( .A(n922), .B(n42879), .Z(n42878) );
  XOR U42818 ( .A(n42880), .B(n42881), .Z(n42837) );
  AND U42819 ( .A(n42882), .B(n42883), .Z(n42881) );
  XNOR U42820 ( .A(n42880), .B(n42572), .Z(n42883) );
  XOR U42821 ( .A(n42778), .B(n42884), .Z(n42572) );
  AND U42822 ( .A(n906), .B(n42885), .Z(n42884) );
  XOR U42823 ( .A(n42774), .B(n42778), .Z(n42885) );
  XNOR U42824 ( .A(n42886), .B(n42880), .Z(n42882) );
  IV U42825 ( .A(n42521), .Z(n42886) );
  XOR U42826 ( .A(n42887), .B(n42888), .Z(n42521) );
  AND U42827 ( .A(n922), .B(n42889), .Z(n42888) );
  AND U42828 ( .A(n42841), .B(n42822), .Z(n42880) );
  XNOR U42829 ( .A(n42890), .B(n42891), .Z(n42822) );
  AND U42830 ( .A(n906), .B(n42800), .Z(n42891) );
  XNOR U42831 ( .A(n42798), .B(n42890), .Z(n42800) );
  XNOR U42832 ( .A(n42892), .B(n42893), .Z(n906) );
  AND U42833 ( .A(n42894), .B(n42895), .Z(n42893) );
  XNOR U42834 ( .A(n42892), .B(n42584), .Z(n42895) );
  IV U42835 ( .A(n42588), .Z(n42584) );
  XOR U42836 ( .A(n42896), .B(n42897), .Z(n42588) );
  AND U42837 ( .A(n910), .B(n42898), .Z(n42897) );
  XOR U42838 ( .A(n42899), .B(n42896), .Z(n42898) );
  XNOR U42839 ( .A(n42892), .B(n42805), .Z(n42894) );
  XOR U42840 ( .A(n42900), .B(n42901), .Z(n42805) );
  AND U42841 ( .A(n918), .B(n42852), .Z(n42901) );
  XOR U42842 ( .A(n42850), .B(n42900), .Z(n42852) );
  XOR U42843 ( .A(n42902), .B(n42903), .Z(n42892) );
  AND U42844 ( .A(n42904), .B(n42905), .Z(n42903) );
  XNOR U42845 ( .A(n42902), .B(n42600), .Z(n42905) );
  IV U42846 ( .A(n42603), .Z(n42600) );
  XOR U42847 ( .A(n42906), .B(n42907), .Z(n42603) );
  AND U42848 ( .A(n910), .B(n42908), .Z(n42907) );
  XOR U42849 ( .A(n42909), .B(n42906), .Z(n42908) );
  XOR U42850 ( .A(n42604), .B(n42902), .Z(n42904) );
  XOR U42851 ( .A(n42910), .B(n42911), .Z(n42604) );
  AND U42852 ( .A(n918), .B(n42862), .Z(n42911) );
  XOR U42853 ( .A(n42910), .B(n42860), .Z(n42862) );
  XOR U42854 ( .A(n42912), .B(n42913), .Z(n42902) );
  AND U42855 ( .A(n42914), .B(n42915), .Z(n42913) );
  XNOR U42856 ( .A(n42912), .B(n42628), .Z(n42915) );
  IV U42857 ( .A(n42631), .Z(n42628) );
  XOR U42858 ( .A(n42916), .B(n42917), .Z(n42631) );
  AND U42859 ( .A(n910), .B(n42918), .Z(n42917) );
  XNOR U42860 ( .A(n42919), .B(n42916), .Z(n42918) );
  XOR U42861 ( .A(n42632), .B(n42912), .Z(n42914) );
  XOR U42862 ( .A(n42920), .B(n42921), .Z(n42632) );
  AND U42863 ( .A(n918), .B(n42871), .Z(n42921) );
  XOR U42864 ( .A(n42920), .B(n42869), .Z(n42871) );
  XOR U42865 ( .A(n42922), .B(n42923), .Z(n42912) );
  AND U42866 ( .A(n42924), .B(n42925), .Z(n42923) );
  XNOR U42867 ( .A(n42922), .B(n42677), .Z(n42925) );
  IV U42868 ( .A(n42680), .Z(n42677) );
  XOR U42869 ( .A(n42926), .B(n42927), .Z(n42680) );
  AND U42870 ( .A(n910), .B(n42928), .Z(n42927) );
  XOR U42871 ( .A(n42929), .B(n42926), .Z(n42928) );
  XOR U42872 ( .A(n42681), .B(n42922), .Z(n42924) );
  XOR U42873 ( .A(n42930), .B(n42931), .Z(n42681) );
  AND U42874 ( .A(n918), .B(n42879), .Z(n42931) );
  XOR U42875 ( .A(n42930), .B(n42877), .Z(n42879) );
  XOR U42876 ( .A(n42818), .B(n42932), .Z(n42922) );
  AND U42877 ( .A(n42820), .B(n42933), .Z(n42932) );
  XNOR U42878 ( .A(n42818), .B(n42774), .Z(n42933) );
  IV U42879 ( .A(n42777), .Z(n42774) );
  XOR U42880 ( .A(n42934), .B(n42935), .Z(n42777) );
  AND U42881 ( .A(n910), .B(n42936), .Z(n42935) );
  XNOR U42882 ( .A(n42937), .B(n42934), .Z(n42936) );
  XOR U42883 ( .A(n42778), .B(n42818), .Z(n42820) );
  XOR U42884 ( .A(n42938), .B(n42939), .Z(n42778) );
  AND U42885 ( .A(n918), .B(n42889), .Z(n42939) );
  XOR U42886 ( .A(n42938), .B(n42887), .Z(n42889) );
  AND U42887 ( .A(n42890), .B(n42798), .Z(n42818) );
  XNOR U42888 ( .A(n42940), .B(n42941), .Z(n42798) );
  AND U42889 ( .A(n910), .B(n42942), .Z(n42941) );
  XNOR U42890 ( .A(n42943), .B(n42940), .Z(n42942) );
  XNOR U42891 ( .A(n42944), .B(n42945), .Z(n910) );
  AND U42892 ( .A(n42946), .B(n42947), .Z(n42945) );
  XOR U42893 ( .A(n42899), .B(n42944), .Z(n42947) );
  AND U42894 ( .A(n42948), .B(n42949), .Z(n42899) );
  XNOR U42895 ( .A(n42896), .B(n42944), .Z(n42946) );
  XNOR U42896 ( .A(n42950), .B(n42951), .Z(n42896) );
  AND U42897 ( .A(n914), .B(n42952), .Z(n42951) );
  XNOR U42898 ( .A(n42953), .B(n42954), .Z(n42952) );
  XOR U42899 ( .A(n42955), .B(n42956), .Z(n42944) );
  AND U42900 ( .A(n42957), .B(n42958), .Z(n42956) );
  XNOR U42901 ( .A(n42955), .B(n42948), .Z(n42958) );
  IV U42902 ( .A(n42909), .Z(n42948) );
  XOR U42903 ( .A(n42959), .B(n42960), .Z(n42909) );
  XOR U42904 ( .A(n42961), .B(n42949), .Z(n42960) );
  AND U42905 ( .A(n42919), .B(n42962), .Z(n42949) );
  AND U42906 ( .A(n42963), .B(n42964), .Z(n42961) );
  XOR U42907 ( .A(n42965), .B(n42959), .Z(n42963) );
  XNOR U42908 ( .A(n42906), .B(n42955), .Z(n42957) );
  XNOR U42909 ( .A(n42966), .B(n42967), .Z(n42906) );
  AND U42910 ( .A(n914), .B(n42968), .Z(n42967) );
  XNOR U42911 ( .A(n42969), .B(n42970), .Z(n42968) );
  XOR U42912 ( .A(n42971), .B(n42972), .Z(n42955) );
  AND U42913 ( .A(n42973), .B(n42974), .Z(n42972) );
  XNOR U42914 ( .A(n42971), .B(n42919), .Z(n42974) );
  XOR U42915 ( .A(n42975), .B(n42964), .Z(n42919) );
  XNOR U42916 ( .A(n42976), .B(n42959), .Z(n42964) );
  XOR U42917 ( .A(n42977), .B(n42978), .Z(n42959) );
  AND U42918 ( .A(n42979), .B(n42980), .Z(n42978) );
  XOR U42919 ( .A(n42981), .B(n42977), .Z(n42979) );
  XNOR U42920 ( .A(n42982), .B(n42983), .Z(n42976) );
  AND U42921 ( .A(n42984), .B(n42985), .Z(n42983) );
  XOR U42922 ( .A(n42982), .B(n42986), .Z(n42984) );
  XNOR U42923 ( .A(n42965), .B(n42962), .Z(n42975) );
  AND U42924 ( .A(n42987), .B(n42988), .Z(n42962) );
  XOR U42925 ( .A(n42989), .B(n42990), .Z(n42965) );
  AND U42926 ( .A(n42991), .B(n42992), .Z(n42990) );
  XOR U42927 ( .A(n42989), .B(n42993), .Z(n42991) );
  XNOR U42928 ( .A(n42916), .B(n42971), .Z(n42973) );
  XNOR U42929 ( .A(n42994), .B(n42995), .Z(n42916) );
  AND U42930 ( .A(n914), .B(n42996), .Z(n42995) );
  XNOR U42931 ( .A(n42997), .B(n42998), .Z(n42996) );
  XOR U42932 ( .A(n42999), .B(n43000), .Z(n42971) );
  AND U42933 ( .A(n43001), .B(n43002), .Z(n43000) );
  XNOR U42934 ( .A(n42999), .B(n42987), .Z(n43002) );
  IV U42935 ( .A(n42929), .Z(n42987) );
  XNOR U42936 ( .A(n43003), .B(n42980), .Z(n42929) );
  XNOR U42937 ( .A(n43004), .B(n42986), .Z(n42980) );
  XOR U42938 ( .A(n43005), .B(n43006), .Z(n42986) );
  AND U42939 ( .A(n43007), .B(n43008), .Z(n43006) );
  XOR U42940 ( .A(n43005), .B(n43009), .Z(n43007) );
  XNOR U42941 ( .A(n42985), .B(n42977), .Z(n43004) );
  XOR U42942 ( .A(n43010), .B(n43011), .Z(n42977) );
  AND U42943 ( .A(n43012), .B(n43013), .Z(n43011) );
  XNOR U42944 ( .A(n43014), .B(n43010), .Z(n43012) );
  XNOR U42945 ( .A(n43015), .B(n42982), .Z(n42985) );
  XOR U42946 ( .A(n43016), .B(n43017), .Z(n42982) );
  AND U42947 ( .A(n43018), .B(n43019), .Z(n43017) );
  XOR U42948 ( .A(n43016), .B(n43020), .Z(n43018) );
  XNOR U42949 ( .A(n43021), .B(n43022), .Z(n43015) );
  AND U42950 ( .A(n43023), .B(n43024), .Z(n43022) );
  XNOR U42951 ( .A(n43021), .B(n43025), .Z(n43023) );
  XNOR U42952 ( .A(n42981), .B(n42988), .Z(n43003) );
  AND U42953 ( .A(n42937), .B(n43026), .Z(n42988) );
  XOR U42954 ( .A(n42993), .B(n42992), .Z(n42981) );
  XNOR U42955 ( .A(n43027), .B(n42989), .Z(n42992) );
  XOR U42956 ( .A(n43028), .B(n43029), .Z(n42989) );
  AND U42957 ( .A(n43030), .B(n43031), .Z(n43029) );
  XOR U42958 ( .A(n43028), .B(n43032), .Z(n43030) );
  XNOR U42959 ( .A(n43033), .B(n43034), .Z(n43027) );
  AND U42960 ( .A(n43035), .B(n43036), .Z(n43034) );
  XOR U42961 ( .A(n43033), .B(n43037), .Z(n43035) );
  XOR U42962 ( .A(n43038), .B(n43039), .Z(n42993) );
  AND U42963 ( .A(n43040), .B(n43041), .Z(n43039) );
  XOR U42964 ( .A(n43038), .B(n43042), .Z(n43040) );
  XNOR U42965 ( .A(n42926), .B(n42999), .Z(n43001) );
  XNOR U42966 ( .A(n43043), .B(n43044), .Z(n42926) );
  AND U42967 ( .A(n914), .B(n43045), .Z(n43044) );
  XNOR U42968 ( .A(n43046), .B(n43047), .Z(n43045) );
  XOR U42969 ( .A(n43048), .B(n43049), .Z(n42999) );
  AND U42970 ( .A(n43050), .B(n43051), .Z(n43049) );
  XNOR U42971 ( .A(n43048), .B(n42937), .Z(n43051) );
  XOR U42972 ( .A(n43052), .B(n43013), .Z(n42937) );
  XNOR U42973 ( .A(n43053), .B(n43020), .Z(n43013) );
  XOR U42974 ( .A(n43009), .B(n43008), .Z(n43020) );
  XNOR U42975 ( .A(n43054), .B(n43005), .Z(n43008) );
  XOR U42976 ( .A(n43055), .B(n43056), .Z(n43005) );
  AND U42977 ( .A(n43057), .B(n43058), .Z(n43056) );
  XNOR U42978 ( .A(n43059), .B(n43060), .Z(n43057) );
  IV U42979 ( .A(n43055), .Z(n43059) );
  XNOR U42980 ( .A(n43061), .B(n43062), .Z(n43054) );
  NOR U42981 ( .A(n43063), .B(n43064), .Z(n43062) );
  XNOR U42982 ( .A(n43061), .B(n43065), .Z(n43063) );
  XOR U42983 ( .A(n43066), .B(n43067), .Z(n43009) );
  NOR U42984 ( .A(n43068), .B(n43069), .Z(n43067) );
  XNOR U42985 ( .A(n43066), .B(n43070), .Z(n43068) );
  XNOR U42986 ( .A(n43019), .B(n43010), .Z(n43053) );
  XOR U42987 ( .A(n43071), .B(n43072), .Z(n43010) );
  AND U42988 ( .A(n43073), .B(n43074), .Z(n43072) );
  XOR U42989 ( .A(n43071), .B(n43075), .Z(n43073) );
  XOR U42990 ( .A(n43076), .B(n43025), .Z(n43019) );
  XOR U42991 ( .A(n43077), .B(n43078), .Z(n43025) );
  NOR U42992 ( .A(n43079), .B(n43080), .Z(n43078) );
  XOR U42993 ( .A(n43077), .B(n43081), .Z(n43079) );
  XNOR U42994 ( .A(n43024), .B(n43016), .Z(n43076) );
  XOR U42995 ( .A(n43082), .B(n43083), .Z(n43016) );
  AND U42996 ( .A(n43084), .B(n43085), .Z(n43083) );
  XOR U42997 ( .A(n43082), .B(n43086), .Z(n43084) );
  XNOR U42998 ( .A(n43087), .B(n43021), .Z(n43024) );
  XOR U42999 ( .A(n43088), .B(n43089), .Z(n43021) );
  AND U43000 ( .A(n43090), .B(n43091), .Z(n43089) );
  XNOR U43001 ( .A(n43092), .B(n43093), .Z(n43090) );
  IV U43002 ( .A(n43088), .Z(n43092) );
  XNOR U43003 ( .A(n43094), .B(n43095), .Z(n43087) );
  NOR U43004 ( .A(n43096), .B(n43097), .Z(n43095) );
  XNOR U43005 ( .A(n43094), .B(n43098), .Z(n43096) );
  XOR U43006 ( .A(n43014), .B(n43026), .Z(n43052) );
  NOR U43007 ( .A(n42943), .B(n43099), .Z(n43026) );
  XNOR U43008 ( .A(n43032), .B(n43031), .Z(n43014) );
  XNOR U43009 ( .A(n43100), .B(n43037), .Z(n43031) );
  XNOR U43010 ( .A(n43101), .B(n43102), .Z(n43037) );
  NOR U43011 ( .A(n43103), .B(n43104), .Z(n43102) );
  XOR U43012 ( .A(n43101), .B(n43105), .Z(n43103) );
  XNOR U43013 ( .A(n43036), .B(n43028), .Z(n43100) );
  XOR U43014 ( .A(n43106), .B(n43107), .Z(n43028) );
  AND U43015 ( .A(n43108), .B(n43109), .Z(n43107) );
  XOR U43016 ( .A(n43106), .B(n43110), .Z(n43108) );
  XNOR U43017 ( .A(n43111), .B(n43033), .Z(n43036) );
  XOR U43018 ( .A(n43112), .B(n43113), .Z(n43033) );
  AND U43019 ( .A(n43114), .B(n43115), .Z(n43113) );
  XNOR U43020 ( .A(n43116), .B(n43117), .Z(n43114) );
  IV U43021 ( .A(n43112), .Z(n43116) );
  XNOR U43022 ( .A(n43118), .B(n43119), .Z(n43111) );
  NOR U43023 ( .A(n43120), .B(n43121), .Z(n43119) );
  XNOR U43024 ( .A(n43118), .B(n43122), .Z(n43120) );
  XOR U43025 ( .A(n43042), .B(n43041), .Z(n43032) );
  XNOR U43026 ( .A(n43123), .B(n43038), .Z(n43041) );
  XOR U43027 ( .A(n43124), .B(n43125), .Z(n43038) );
  AND U43028 ( .A(n43126), .B(n43127), .Z(n43125) );
  XNOR U43029 ( .A(n43128), .B(n43129), .Z(n43126) );
  IV U43030 ( .A(n43124), .Z(n43128) );
  XNOR U43031 ( .A(n43130), .B(n43131), .Z(n43123) );
  NOR U43032 ( .A(n43132), .B(n43133), .Z(n43131) );
  XNOR U43033 ( .A(n43130), .B(n43134), .Z(n43132) );
  XOR U43034 ( .A(n43135), .B(n43136), .Z(n43042) );
  NOR U43035 ( .A(n43137), .B(n43138), .Z(n43136) );
  XNOR U43036 ( .A(n43135), .B(n43139), .Z(n43137) );
  XNOR U43037 ( .A(n42934), .B(n43048), .Z(n43050) );
  XNOR U43038 ( .A(n43140), .B(n43141), .Z(n42934) );
  AND U43039 ( .A(n914), .B(n43142), .Z(n43141) );
  XNOR U43040 ( .A(n43143), .B(n43144), .Z(n43142) );
  AND U43041 ( .A(n42940), .B(n42943), .Z(n43048) );
  XOR U43042 ( .A(n43145), .B(n43099), .Z(n42943) );
  XNOR U43043 ( .A(p_input[1312]), .B(p_input[2048]), .Z(n43099) );
  XNOR U43044 ( .A(n43075), .B(n43074), .Z(n43145) );
  XNOR U43045 ( .A(n43146), .B(n43086), .Z(n43074) );
  XOR U43046 ( .A(n43060), .B(n43058), .Z(n43086) );
  XNOR U43047 ( .A(n43147), .B(n43065), .Z(n43058) );
  XOR U43048 ( .A(p_input[1336]), .B(p_input[2072]), .Z(n43065) );
  XOR U43049 ( .A(n43055), .B(n43064), .Z(n43147) );
  XOR U43050 ( .A(n43148), .B(n43061), .Z(n43064) );
  XOR U43051 ( .A(p_input[1334]), .B(p_input[2070]), .Z(n43061) );
  XOR U43052 ( .A(p_input[1335]), .B(n29410), .Z(n43148) );
  XOR U43053 ( .A(p_input[1330]), .B(p_input[2066]), .Z(n43055) );
  XNOR U43054 ( .A(n43070), .B(n43069), .Z(n43060) );
  XOR U43055 ( .A(n43149), .B(n43066), .Z(n43069) );
  XOR U43056 ( .A(p_input[1331]), .B(p_input[2067]), .Z(n43066) );
  XOR U43057 ( .A(p_input[1332]), .B(n29412), .Z(n43149) );
  XOR U43058 ( .A(p_input[1333]), .B(p_input[2069]), .Z(n43070) );
  XOR U43059 ( .A(n43085), .B(n43150), .Z(n43146) );
  IV U43060 ( .A(n43071), .Z(n43150) );
  XOR U43061 ( .A(p_input[1313]), .B(p_input[2049]), .Z(n43071) );
  XNOR U43062 ( .A(n43151), .B(n43093), .Z(n43085) );
  XNOR U43063 ( .A(n43081), .B(n43080), .Z(n43093) );
  XNOR U43064 ( .A(n43152), .B(n43077), .Z(n43080) );
  XNOR U43065 ( .A(p_input[1338]), .B(p_input[2074]), .Z(n43077) );
  XOR U43066 ( .A(p_input[1339]), .B(n29415), .Z(n43152) );
  XOR U43067 ( .A(p_input[1340]), .B(p_input[2076]), .Z(n43081) );
  XOR U43068 ( .A(n43091), .B(n43153), .Z(n43151) );
  IV U43069 ( .A(n43082), .Z(n43153) );
  XOR U43070 ( .A(p_input[1329]), .B(p_input[2065]), .Z(n43082) );
  XNOR U43071 ( .A(n43154), .B(n43098), .Z(n43091) );
  XNOR U43072 ( .A(p_input[1343]), .B(n29418), .Z(n43098) );
  XOR U43073 ( .A(n43088), .B(n43097), .Z(n43154) );
  XOR U43074 ( .A(n43155), .B(n43094), .Z(n43097) );
  XOR U43075 ( .A(p_input[1341]), .B(p_input[2077]), .Z(n43094) );
  XOR U43076 ( .A(p_input[1342]), .B(n29420), .Z(n43155) );
  XOR U43077 ( .A(p_input[1337]), .B(p_input[2073]), .Z(n43088) );
  XOR U43078 ( .A(n43110), .B(n43109), .Z(n43075) );
  XNOR U43079 ( .A(n43156), .B(n43117), .Z(n43109) );
  XNOR U43080 ( .A(n43105), .B(n43104), .Z(n43117) );
  XNOR U43081 ( .A(n43157), .B(n43101), .Z(n43104) );
  XNOR U43082 ( .A(p_input[1323]), .B(p_input[2059]), .Z(n43101) );
  XOR U43083 ( .A(p_input[1324]), .B(n28329), .Z(n43157) );
  XOR U43084 ( .A(p_input[1325]), .B(p_input[2061]), .Z(n43105) );
  XOR U43085 ( .A(n43115), .B(n43158), .Z(n43156) );
  IV U43086 ( .A(n43106), .Z(n43158) );
  XOR U43087 ( .A(p_input[1314]), .B(p_input[2050]), .Z(n43106) );
  XNOR U43088 ( .A(n43159), .B(n43122), .Z(n43115) );
  XNOR U43089 ( .A(p_input[1328]), .B(n28332), .Z(n43122) );
  XOR U43090 ( .A(n43112), .B(n43121), .Z(n43159) );
  XOR U43091 ( .A(n43160), .B(n43118), .Z(n43121) );
  XOR U43092 ( .A(p_input[1326]), .B(p_input[2062]), .Z(n43118) );
  XOR U43093 ( .A(p_input[1327]), .B(n28334), .Z(n43160) );
  XOR U43094 ( .A(p_input[1322]), .B(p_input[2058]), .Z(n43112) );
  XOR U43095 ( .A(n43129), .B(n43127), .Z(n43110) );
  XNOR U43096 ( .A(n43161), .B(n43134), .Z(n43127) );
  XOR U43097 ( .A(p_input[1321]), .B(p_input[2057]), .Z(n43134) );
  XOR U43098 ( .A(n43124), .B(n43133), .Z(n43161) );
  XOR U43099 ( .A(n43162), .B(n43130), .Z(n43133) );
  XOR U43100 ( .A(p_input[1319]), .B(p_input[2055]), .Z(n43130) );
  XOR U43101 ( .A(p_input[1320]), .B(n29427), .Z(n43162) );
  XOR U43102 ( .A(p_input[1315]), .B(p_input[2051]), .Z(n43124) );
  XNOR U43103 ( .A(n43139), .B(n43138), .Z(n43129) );
  XOR U43104 ( .A(n43163), .B(n43135), .Z(n43138) );
  XOR U43105 ( .A(p_input[1316]), .B(p_input[2052]), .Z(n43135) );
  XOR U43106 ( .A(p_input[1317]), .B(n29429), .Z(n43163) );
  XOR U43107 ( .A(p_input[1318]), .B(p_input[2054]), .Z(n43139) );
  XNOR U43108 ( .A(n43164), .B(n43165), .Z(n42940) );
  AND U43109 ( .A(n914), .B(n43166), .Z(n43165) );
  XNOR U43110 ( .A(n43167), .B(n43168), .Z(n914) );
  AND U43111 ( .A(n43169), .B(n43170), .Z(n43168) );
  XOR U43112 ( .A(n42954), .B(n43167), .Z(n43170) );
  XNOR U43113 ( .A(n43171), .B(n43167), .Z(n43169) );
  XOR U43114 ( .A(n43172), .B(n43173), .Z(n43167) );
  AND U43115 ( .A(n43174), .B(n43175), .Z(n43173) );
  XOR U43116 ( .A(n42969), .B(n43172), .Z(n43175) );
  XOR U43117 ( .A(n43172), .B(n42970), .Z(n43174) );
  XOR U43118 ( .A(n43176), .B(n43177), .Z(n43172) );
  AND U43119 ( .A(n43178), .B(n43179), .Z(n43177) );
  XOR U43120 ( .A(n42997), .B(n43176), .Z(n43179) );
  XOR U43121 ( .A(n43176), .B(n42998), .Z(n43178) );
  XOR U43122 ( .A(n43180), .B(n43181), .Z(n43176) );
  AND U43123 ( .A(n43182), .B(n43183), .Z(n43181) );
  XOR U43124 ( .A(n43046), .B(n43180), .Z(n43183) );
  XOR U43125 ( .A(n43180), .B(n43047), .Z(n43182) );
  XOR U43126 ( .A(n43184), .B(n43185), .Z(n43180) );
  AND U43127 ( .A(n43186), .B(n43187), .Z(n43185) );
  XOR U43128 ( .A(n43184), .B(n43143), .Z(n43187) );
  XNOR U43129 ( .A(n43188), .B(n43189), .Z(n42890) );
  AND U43130 ( .A(n918), .B(n43190), .Z(n43189) );
  XNOR U43131 ( .A(n43191), .B(n43192), .Z(n918) );
  AND U43132 ( .A(n43193), .B(n43194), .Z(n43192) );
  XOR U43133 ( .A(n43191), .B(n42900), .Z(n43194) );
  XNOR U43134 ( .A(n43191), .B(n42850), .Z(n43193) );
  XOR U43135 ( .A(n43195), .B(n43196), .Z(n43191) );
  AND U43136 ( .A(n43197), .B(n43198), .Z(n43196) );
  XNOR U43137 ( .A(n42910), .B(n43195), .Z(n43198) );
  XOR U43138 ( .A(n43195), .B(n42860), .Z(n43197) );
  XOR U43139 ( .A(n43199), .B(n43200), .Z(n43195) );
  AND U43140 ( .A(n43201), .B(n43202), .Z(n43200) );
  XNOR U43141 ( .A(n42920), .B(n43199), .Z(n43202) );
  XOR U43142 ( .A(n43199), .B(n42869), .Z(n43201) );
  XOR U43143 ( .A(n43203), .B(n43204), .Z(n43199) );
  AND U43144 ( .A(n43205), .B(n43206), .Z(n43204) );
  XOR U43145 ( .A(n43203), .B(n42877), .Z(n43205) );
  XOR U43146 ( .A(n43207), .B(n43208), .Z(n42841) );
  AND U43147 ( .A(n922), .B(n43190), .Z(n43208) );
  XNOR U43148 ( .A(n43188), .B(n43207), .Z(n43190) );
  XNOR U43149 ( .A(n43209), .B(n43210), .Z(n922) );
  AND U43150 ( .A(n43211), .B(n43212), .Z(n43210) );
  XNOR U43151 ( .A(n43213), .B(n43209), .Z(n43212) );
  IV U43152 ( .A(n42900), .Z(n43213) );
  XOR U43153 ( .A(n43171), .B(n43214), .Z(n42900) );
  AND U43154 ( .A(n925), .B(n43215), .Z(n43214) );
  XOR U43155 ( .A(n42953), .B(n42950), .Z(n43215) );
  IV U43156 ( .A(n43171), .Z(n42953) );
  XNOR U43157 ( .A(n42850), .B(n43209), .Z(n43211) );
  XOR U43158 ( .A(n43216), .B(n43217), .Z(n42850) );
  AND U43159 ( .A(n941), .B(n43218), .Z(n43217) );
  XOR U43160 ( .A(n43219), .B(n43220), .Z(n43209) );
  AND U43161 ( .A(n43221), .B(n43222), .Z(n43220) );
  XNOR U43162 ( .A(n43219), .B(n42910), .Z(n43222) );
  XOR U43163 ( .A(n42970), .B(n43223), .Z(n42910) );
  AND U43164 ( .A(n925), .B(n43224), .Z(n43223) );
  XOR U43165 ( .A(n42966), .B(n42970), .Z(n43224) );
  XNOR U43166 ( .A(n43225), .B(n43219), .Z(n43221) );
  IV U43167 ( .A(n42860), .Z(n43225) );
  XOR U43168 ( .A(n43226), .B(n43227), .Z(n42860) );
  AND U43169 ( .A(n941), .B(n43228), .Z(n43227) );
  XOR U43170 ( .A(n43229), .B(n43230), .Z(n43219) );
  AND U43171 ( .A(n43231), .B(n43232), .Z(n43230) );
  XNOR U43172 ( .A(n43229), .B(n42920), .Z(n43232) );
  XOR U43173 ( .A(n42998), .B(n43233), .Z(n42920) );
  AND U43174 ( .A(n925), .B(n43234), .Z(n43233) );
  XOR U43175 ( .A(n42994), .B(n42998), .Z(n43234) );
  XOR U43176 ( .A(n42869), .B(n43229), .Z(n43231) );
  XOR U43177 ( .A(n43235), .B(n43236), .Z(n42869) );
  AND U43178 ( .A(n941), .B(n43237), .Z(n43236) );
  XOR U43179 ( .A(n43203), .B(n43238), .Z(n43229) );
  AND U43180 ( .A(n43239), .B(n43206), .Z(n43238) );
  XNOR U43181 ( .A(n42930), .B(n43203), .Z(n43206) );
  XOR U43182 ( .A(n43047), .B(n43240), .Z(n42930) );
  AND U43183 ( .A(n925), .B(n43241), .Z(n43240) );
  XOR U43184 ( .A(n43043), .B(n43047), .Z(n43241) );
  XNOR U43185 ( .A(n43242), .B(n43203), .Z(n43239) );
  IV U43186 ( .A(n42877), .Z(n43242) );
  XOR U43187 ( .A(n43243), .B(n43244), .Z(n42877) );
  AND U43188 ( .A(n941), .B(n43245), .Z(n43244) );
  XOR U43189 ( .A(n43246), .B(n43247), .Z(n43203) );
  AND U43190 ( .A(n43248), .B(n43249), .Z(n43247) );
  XNOR U43191 ( .A(n43246), .B(n42938), .Z(n43249) );
  XOR U43192 ( .A(n43144), .B(n43250), .Z(n42938) );
  AND U43193 ( .A(n925), .B(n43251), .Z(n43250) );
  XOR U43194 ( .A(n43140), .B(n43144), .Z(n43251) );
  XNOR U43195 ( .A(n43252), .B(n43246), .Z(n43248) );
  IV U43196 ( .A(n42887), .Z(n43252) );
  XOR U43197 ( .A(n43253), .B(n43254), .Z(n42887) );
  AND U43198 ( .A(n941), .B(n43255), .Z(n43254) );
  AND U43199 ( .A(n43207), .B(n43188), .Z(n43246) );
  XNOR U43200 ( .A(n43256), .B(n43257), .Z(n43188) );
  AND U43201 ( .A(n925), .B(n43166), .Z(n43257) );
  XNOR U43202 ( .A(n43164), .B(n43256), .Z(n43166) );
  XNOR U43203 ( .A(n43258), .B(n43259), .Z(n925) );
  AND U43204 ( .A(n43260), .B(n43261), .Z(n43259) );
  XNOR U43205 ( .A(n43258), .B(n42950), .Z(n43261) );
  IV U43206 ( .A(n42954), .Z(n42950) );
  XOR U43207 ( .A(n43262), .B(n43263), .Z(n42954) );
  AND U43208 ( .A(n929), .B(n43264), .Z(n43263) );
  XOR U43209 ( .A(n43265), .B(n43262), .Z(n43264) );
  XNOR U43210 ( .A(n43258), .B(n43171), .Z(n43260) );
  XOR U43211 ( .A(n43266), .B(n43267), .Z(n43171) );
  AND U43212 ( .A(n937), .B(n43218), .Z(n43267) );
  XOR U43213 ( .A(n43216), .B(n43266), .Z(n43218) );
  XOR U43214 ( .A(n43268), .B(n43269), .Z(n43258) );
  AND U43215 ( .A(n43270), .B(n43271), .Z(n43269) );
  XNOR U43216 ( .A(n43268), .B(n42966), .Z(n43271) );
  IV U43217 ( .A(n42969), .Z(n42966) );
  XOR U43218 ( .A(n43272), .B(n43273), .Z(n42969) );
  AND U43219 ( .A(n929), .B(n43274), .Z(n43273) );
  XOR U43220 ( .A(n43275), .B(n43272), .Z(n43274) );
  XOR U43221 ( .A(n42970), .B(n43268), .Z(n43270) );
  XOR U43222 ( .A(n43276), .B(n43277), .Z(n42970) );
  AND U43223 ( .A(n937), .B(n43228), .Z(n43277) );
  XOR U43224 ( .A(n43276), .B(n43226), .Z(n43228) );
  XOR U43225 ( .A(n43278), .B(n43279), .Z(n43268) );
  AND U43226 ( .A(n43280), .B(n43281), .Z(n43279) );
  XNOR U43227 ( .A(n43278), .B(n42994), .Z(n43281) );
  IV U43228 ( .A(n42997), .Z(n42994) );
  XOR U43229 ( .A(n43282), .B(n43283), .Z(n42997) );
  AND U43230 ( .A(n929), .B(n43284), .Z(n43283) );
  XNOR U43231 ( .A(n43285), .B(n43282), .Z(n43284) );
  XOR U43232 ( .A(n42998), .B(n43278), .Z(n43280) );
  XOR U43233 ( .A(n43286), .B(n43287), .Z(n42998) );
  AND U43234 ( .A(n937), .B(n43237), .Z(n43287) );
  XOR U43235 ( .A(n43286), .B(n43235), .Z(n43237) );
  XOR U43236 ( .A(n43288), .B(n43289), .Z(n43278) );
  AND U43237 ( .A(n43290), .B(n43291), .Z(n43289) );
  XNOR U43238 ( .A(n43288), .B(n43043), .Z(n43291) );
  IV U43239 ( .A(n43046), .Z(n43043) );
  XOR U43240 ( .A(n43292), .B(n43293), .Z(n43046) );
  AND U43241 ( .A(n929), .B(n43294), .Z(n43293) );
  XOR U43242 ( .A(n43295), .B(n43292), .Z(n43294) );
  XOR U43243 ( .A(n43047), .B(n43288), .Z(n43290) );
  XOR U43244 ( .A(n43296), .B(n43297), .Z(n43047) );
  AND U43245 ( .A(n937), .B(n43245), .Z(n43297) );
  XOR U43246 ( .A(n43296), .B(n43243), .Z(n43245) );
  XOR U43247 ( .A(n43184), .B(n43298), .Z(n43288) );
  AND U43248 ( .A(n43186), .B(n43299), .Z(n43298) );
  XNOR U43249 ( .A(n43184), .B(n43140), .Z(n43299) );
  IV U43250 ( .A(n43143), .Z(n43140) );
  XOR U43251 ( .A(n43300), .B(n43301), .Z(n43143) );
  AND U43252 ( .A(n929), .B(n43302), .Z(n43301) );
  XNOR U43253 ( .A(n43303), .B(n43300), .Z(n43302) );
  XOR U43254 ( .A(n43144), .B(n43184), .Z(n43186) );
  XOR U43255 ( .A(n43304), .B(n43305), .Z(n43144) );
  AND U43256 ( .A(n937), .B(n43255), .Z(n43305) );
  XOR U43257 ( .A(n43304), .B(n43253), .Z(n43255) );
  AND U43258 ( .A(n43256), .B(n43164), .Z(n43184) );
  XNOR U43259 ( .A(n43306), .B(n43307), .Z(n43164) );
  AND U43260 ( .A(n929), .B(n43308), .Z(n43307) );
  XNOR U43261 ( .A(n43309), .B(n43306), .Z(n43308) );
  XNOR U43262 ( .A(n43310), .B(n43311), .Z(n929) );
  AND U43263 ( .A(n43312), .B(n43313), .Z(n43311) );
  XOR U43264 ( .A(n43265), .B(n43310), .Z(n43313) );
  AND U43265 ( .A(n43314), .B(n43315), .Z(n43265) );
  XNOR U43266 ( .A(n43262), .B(n43310), .Z(n43312) );
  XNOR U43267 ( .A(n43316), .B(n43317), .Z(n43262) );
  AND U43268 ( .A(n933), .B(n43318), .Z(n43317) );
  XNOR U43269 ( .A(n43319), .B(n43320), .Z(n43318) );
  XOR U43270 ( .A(n43321), .B(n43322), .Z(n43310) );
  AND U43271 ( .A(n43323), .B(n43324), .Z(n43322) );
  XNOR U43272 ( .A(n43321), .B(n43314), .Z(n43324) );
  IV U43273 ( .A(n43275), .Z(n43314) );
  XOR U43274 ( .A(n43325), .B(n43326), .Z(n43275) );
  XOR U43275 ( .A(n43327), .B(n43315), .Z(n43326) );
  AND U43276 ( .A(n43285), .B(n43328), .Z(n43315) );
  AND U43277 ( .A(n43329), .B(n43330), .Z(n43327) );
  XOR U43278 ( .A(n43331), .B(n43325), .Z(n43329) );
  XNOR U43279 ( .A(n43272), .B(n43321), .Z(n43323) );
  XNOR U43280 ( .A(n43332), .B(n43333), .Z(n43272) );
  AND U43281 ( .A(n933), .B(n43334), .Z(n43333) );
  XNOR U43282 ( .A(n43335), .B(n43336), .Z(n43334) );
  XOR U43283 ( .A(n43337), .B(n43338), .Z(n43321) );
  AND U43284 ( .A(n43339), .B(n43340), .Z(n43338) );
  XNOR U43285 ( .A(n43337), .B(n43285), .Z(n43340) );
  XOR U43286 ( .A(n43341), .B(n43330), .Z(n43285) );
  XNOR U43287 ( .A(n43342), .B(n43325), .Z(n43330) );
  XOR U43288 ( .A(n43343), .B(n43344), .Z(n43325) );
  AND U43289 ( .A(n43345), .B(n43346), .Z(n43344) );
  XOR U43290 ( .A(n43347), .B(n43343), .Z(n43345) );
  XNOR U43291 ( .A(n43348), .B(n43349), .Z(n43342) );
  AND U43292 ( .A(n43350), .B(n43351), .Z(n43349) );
  XOR U43293 ( .A(n43348), .B(n43352), .Z(n43350) );
  XNOR U43294 ( .A(n43331), .B(n43328), .Z(n43341) );
  AND U43295 ( .A(n43353), .B(n43354), .Z(n43328) );
  XOR U43296 ( .A(n43355), .B(n43356), .Z(n43331) );
  AND U43297 ( .A(n43357), .B(n43358), .Z(n43356) );
  XOR U43298 ( .A(n43355), .B(n43359), .Z(n43357) );
  XNOR U43299 ( .A(n43282), .B(n43337), .Z(n43339) );
  XNOR U43300 ( .A(n43360), .B(n43361), .Z(n43282) );
  AND U43301 ( .A(n933), .B(n43362), .Z(n43361) );
  XNOR U43302 ( .A(n43363), .B(n43364), .Z(n43362) );
  XOR U43303 ( .A(n43365), .B(n43366), .Z(n43337) );
  AND U43304 ( .A(n43367), .B(n43368), .Z(n43366) );
  XNOR U43305 ( .A(n43365), .B(n43353), .Z(n43368) );
  IV U43306 ( .A(n43295), .Z(n43353) );
  XNOR U43307 ( .A(n43369), .B(n43346), .Z(n43295) );
  XNOR U43308 ( .A(n43370), .B(n43352), .Z(n43346) );
  XOR U43309 ( .A(n43371), .B(n43372), .Z(n43352) );
  AND U43310 ( .A(n43373), .B(n43374), .Z(n43372) );
  XOR U43311 ( .A(n43371), .B(n43375), .Z(n43373) );
  XNOR U43312 ( .A(n43351), .B(n43343), .Z(n43370) );
  XOR U43313 ( .A(n43376), .B(n43377), .Z(n43343) );
  AND U43314 ( .A(n43378), .B(n43379), .Z(n43377) );
  XNOR U43315 ( .A(n43380), .B(n43376), .Z(n43378) );
  XNOR U43316 ( .A(n43381), .B(n43348), .Z(n43351) );
  XOR U43317 ( .A(n43382), .B(n43383), .Z(n43348) );
  AND U43318 ( .A(n43384), .B(n43385), .Z(n43383) );
  XOR U43319 ( .A(n43382), .B(n43386), .Z(n43384) );
  XNOR U43320 ( .A(n43387), .B(n43388), .Z(n43381) );
  AND U43321 ( .A(n43389), .B(n43390), .Z(n43388) );
  XNOR U43322 ( .A(n43387), .B(n43391), .Z(n43389) );
  XNOR U43323 ( .A(n43347), .B(n43354), .Z(n43369) );
  AND U43324 ( .A(n43303), .B(n43392), .Z(n43354) );
  XOR U43325 ( .A(n43359), .B(n43358), .Z(n43347) );
  XNOR U43326 ( .A(n43393), .B(n43355), .Z(n43358) );
  XOR U43327 ( .A(n43394), .B(n43395), .Z(n43355) );
  AND U43328 ( .A(n43396), .B(n43397), .Z(n43395) );
  XOR U43329 ( .A(n43394), .B(n43398), .Z(n43396) );
  XNOR U43330 ( .A(n43399), .B(n43400), .Z(n43393) );
  AND U43331 ( .A(n43401), .B(n43402), .Z(n43400) );
  XOR U43332 ( .A(n43399), .B(n43403), .Z(n43401) );
  XOR U43333 ( .A(n43404), .B(n43405), .Z(n43359) );
  AND U43334 ( .A(n43406), .B(n43407), .Z(n43405) );
  XOR U43335 ( .A(n43404), .B(n43408), .Z(n43406) );
  XNOR U43336 ( .A(n43292), .B(n43365), .Z(n43367) );
  XNOR U43337 ( .A(n43409), .B(n43410), .Z(n43292) );
  AND U43338 ( .A(n933), .B(n43411), .Z(n43410) );
  XNOR U43339 ( .A(n43412), .B(n43413), .Z(n43411) );
  XOR U43340 ( .A(n43414), .B(n43415), .Z(n43365) );
  AND U43341 ( .A(n43416), .B(n43417), .Z(n43415) );
  XNOR U43342 ( .A(n43414), .B(n43303), .Z(n43417) );
  XOR U43343 ( .A(n43418), .B(n43379), .Z(n43303) );
  XNOR U43344 ( .A(n43419), .B(n43386), .Z(n43379) );
  XOR U43345 ( .A(n43375), .B(n43374), .Z(n43386) );
  XNOR U43346 ( .A(n43420), .B(n43371), .Z(n43374) );
  XOR U43347 ( .A(n43421), .B(n43422), .Z(n43371) );
  AND U43348 ( .A(n43423), .B(n43424), .Z(n43422) );
  XNOR U43349 ( .A(n43425), .B(n43426), .Z(n43423) );
  IV U43350 ( .A(n43421), .Z(n43425) );
  XNOR U43351 ( .A(n43427), .B(n43428), .Z(n43420) );
  NOR U43352 ( .A(n43429), .B(n43430), .Z(n43428) );
  XNOR U43353 ( .A(n43427), .B(n43431), .Z(n43429) );
  XOR U43354 ( .A(n43432), .B(n43433), .Z(n43375) );
  NOR U43355 ( .A(n43434), .B(n43435), .Z(n43433) );
  XNOR U43356 ( .A(n43432), .B(n43436), .Z(n43434) );
  XNOR U43357 ( .A(n43385), .B(n43376), .Z(n43419) );
  XOR U43358 ( .A(n43437), .B(n43438), .Z(n43376) );
  AND U43359 ( .A(n43439), .B(n43440), .Z(n43438) );
  XOR U43360 ( .A(n43437), .B(n43441), .Z(n43439) );
  XOR U43361 ( .A(n43442), .B(n43391), .Z(n43385) );
  XOR U43362 ( .A(n43443), .B(n43444), .Z(n43391) );
  NOR U43363 ( .A(n43445), .B(n43446), .Z(n43444) );
  XOR U43364 ( .A(n43443), .B(n43447), .Z(n43445) );
  XNOR U43365 ( .A(n43390), .B(n43382), .Z(n43442) );
  XOR U43366 ( .A(n43448), .B(n43449), .Z(n43382) );
  AND U43367 ( .A(n43450), .B(n43451), .Z(n43449) );
  XOR U43368 ( .A(n43448), .B(n43452), .Z(n43450) );
  XNOR U43369 ( .A(n43453), .B(n43387), .Z(n43390) );
  XOR U43370 ( .A(n43454), .B(n43455), .Z(n43387) );
  AND U43371 ( .A(n43456), .B(n43457), .Z(n43455) );
  XNOR U43372 ( .A(n43458), .B(n43459), .Z(n43456) );
  IV U43373 ( .A(n43454), .Z(n43458) );
  XNOR U43374 ( .A(n43460), .B(n43461), .Z(n43453) );
  NOR U43375 ( .A(n43462), .B(n43463), .Z(n43461) );
  XNOR U43376 ( .A(n43460), .B(n43464), .Z(n43462) );
  XOR U43377 ( .A(n43380), .B(n43392), .Z(n43418) );
  NOR U43378 ( .A(n43309), .B(n43465), .Z(n43392) );
  XNOR U43379 ( .A(n43398), .B(n43397), .Z(n43380) );
  XNOR U43380 ( .A(n43466), .B(n43403), .Z(n43397) );
  XNOR U43381 ( .A(n43467), .B(n43468), .Z(n43403) );
  NOR U43382 ( .A(n43469), .B(n43470), .Z(n43468) );
  XOR U43383 ( .A(n43467), .B(n43471), .Z(n43469) );
  XNOR U43384 ( .A(n43402), .B(n43394), .Z(n43466) );
  XOR U43385 ( .A(n43472), .B(n43473), .Z(n43394) );
  AND U43386 ( .A(n43474), .B(n43475), .Z(n43473) );
  XOR U43387 ( .A(n43472), .B(n43476), .Z(n43474) );
  XNOR U43388 ( .A(n43477), .B(n43399), .Z(n43402) );
  XOR U43389 ( .A(n43478), .B(n43479), .Z(n43399) );
  AND U43390 ( .A(n43480), .B(n43481), .Z(n43479) );
  XNOR U43391 ( .A(n43482), .B(n43483), .Z(n43480) );
  IV U43392 ( .A(n43478), .Z(n43482) );
  XNOR U43393 ( .A(n43484), .B(n43485), .Z(n43477) );
  NOR U43394 ( .A(n43486), .B(n43487), .Z(n43485) );
  XNOR U43395 ( .A(n43484), .B(n43488), .Z(n43486) );
  XOR U43396 ( .A(n43408), .B(n43407), .Z(n43398) );
  XNOR U43397 ( .A(n43489), .B(n43404), .Z(n43407) );
  XOR U43398 ( .A(n43490), .B(n43491), .Z(n43404) );
  AND U43399 ( .A(n43492), .B(n43493), .Z(n43491) );
  XNOR U43400 ( .A(n43494), .B(n43495), .Z(n43492) );
  IV U43401 ( .A(n43490), .Z(n43494) );
  XNOR U43402 ( .A(n43496), .B(n43497), .Z(n43489) );
  NOR U43403 ( .A(n43498), .B(n43499), .Z(n43497) );
  XNOR U43404 ( .A(n43496), .B(n43500), .Z(n43498) );
  XOR U43405 ( .A(n43501), .B(n43502), .Z(n43408) );
  NOR U43406 ( .A(n43503), .B(n43504), .Z(n43502) );
  XNOR U43407 ( .A(n43501), .B(n43505), .Z(n43503) );
  XNOR U43408 ( .A(n43300), .B(n43414), .Z(n43416) );
  XNOR U43409 ( .A(n43506), .B(n43507), .Z(n43300) );
  AND U43410 ( .A(n933), .B(n43508), .Z(n43507) );
  XNOR U43411 ( .A(n43509), .B(n43510), .Z(n43508) );
  AND U43412 ( .A(n43306), .B(n43309), .Z(n43414) );
  XOR U43413 ( .A(n43511), .B(n43465), .Z(n43309) );
  XNOR U43414 ( .A(p_input[1344]), .B(p_input[2048]), .Z(n43465) );
  XNOR U43415 ( .A(n43441), .B(n43440), .Z(n43511) );
  XNOR U43416 ( .A(n43512), .B(n43452), .Z(n43440) );
  XOR U43417 ( .A(n43426), .B(n43424), .Z(n43452) );
  XNOR U43418 ( .A(n43513), .B(n43431), .Z(n43424) );
  XOR U43419 ( .A(p_input[1368]), .B(p_input[2072]), .Z(n43431) );
  XOR U43420 ( .A(n43421), .B(n43430), .Z(n43513) );
  XOR U43421 ( .A(n43514), .B(n43427), .Z(n43430) );
  XOR U43422 ( .A(p_input[1366]), .B(p_input[2070]), .Z(n43427) );
  XOR U43423 ( .A(p_input[1367]), .B(n29410), .Z(n43514) );
  XOR U43424 ( .A(p_input[1362]), .B(p_input[2066]), .Z(n43421) );
  XNOR U43425 ( .A(n43436), .B(n43435), .Z(n43426) );
  XOR U43426 ( .A(n43515), .B(n43432), .Z(n43435) );
  XOR U43427 ( .A(p_input[1363]), .B(p_input[2067]), .Z(n43432) );
  XOR U43428 ( .A(p_input[1364]), .B(n29412), .Z(n43515) );
  XOR U43429 ( .A(p_input[1365]), .B(p_input[2069]), .Z(n43436) );
  XOR U43430 ( .A(n43451), .B(n43516), .Z(n43512) );
  IV U43431 ( .A(n43437), .Z(n43516) );
  XOR U43432 ( .A(p_input[1345]), .B(p_input[2049]), .Z(n43437) );
  XNOR U43433 ( .A(n43517), .B(n43459), .Z(n43451) );
  XNOR U43434 ( .A(n43447), .B(n43446), .Z(n43459) );
  XNOR U43435 ( .A(n43518), .B(n43443), .Z(n43446) );
  XNOR U43436 ( .A(p_input[1370]), .B(p_input[2074]), .Z(n43443) );
  XOR U43437 ( .A(p_input[1371]), .B(n29415), .Z(n43518) );
  XOR U43438 ( .A(p_input[1372]), .B(p_input[2076]), .Z(n43447) );
  XOR U43439 ( .A(n43457), .B(n43519), .Z(n43517) );
  IV U43440 ( .A(n43448), .Z(n43519) );
  XOR U43441 ( .A(p_input[1361]), .B(p_input[2065]), .Z(n43448) );
  XNOR U43442 ( .A(n43520), .B(n43464), .Z(n43457) );
  XNOR U43443 ( .A(p_input[1375]), .B(n29418), .Z(n43464) );
  XOR U43444 ( .A(n43454), .B(n43463), .Z(n43520) );
  XOR U43445 ( .A(n43521), .B(n43460), .Z(n43463) );
  XOR U43446 ( .A(p_input[1373]), .B(p_input[2077]), .Z(n43460) );
  XOR U43447 ( .A(p_input[1374]), .B(n29420), .Z(n43521) );
  XOR U43448 ( .A(p_input[1369]), .B(p_input[2073]), .Z(n43454) );
  XOR U43449 ( .A(n43476), .B(n43475), .Z(n43441) );
  XNOR U43450 ( .A(n43522), .B(n43483), .Z(n43475) );
  XNOR U43451 ( .A(n43471), .B(n43470), .Z(n43483) );
  XNOR U43452 ( .A(n43523), .B(n43467), .Z(n43470) );
  XNOR U43453 ( .A(p_input[1355]), .B(p_input[2059]), .Z(n43467) );
  XOR U43454 ( .A(p_input[1356]), .B(n28329), .Z(n43523) );
  XOR U43455 ( .A(p_input[1357]), .B(p_input[2061]), .Z(n43471) );
  XOR U43456 ( .A(n43481), .B(n43524), .Z(n43522) );
  IV U43457 ( .A(n43472), .Z(n43524) );
  XOR U43458 ( .A(p_input[1346]), .B(p_input[2050]), .Z(n43472) );
  XNOR U43459 ( .A(n43525), .B(n43488), .Z(n43481) );
  XNOR U43460 ( .A(p_input[1360]), .B(n28332), .Z(n43488) );
  XOR U43461 ( .A(n43478), .B(n43487), .Z(n43525) );
  XOR U43462 ( .A(n43526), .B(n43484), .Z(n43487) );
  XOR U43463 ( .A(p_input[1358]), .B(p_input[2062]), .Z(n43484) );
  XOR U43464 ( .A(p_input[1359]), .B(n28334), .Z(n43526) );
  XOR U43465 ( .A(p_input[1354]), .B(p_input[2058]), .Z(n43478) );
  XOR U43466 ( .A(n43495), .B(n43493), .Z(n43476) );
  XNOR U43467 ( .A(n43527), .B(n43500), .Z(n43493) );
  XOR U43468 ( .A(p_input[1353]), .B(p_input[2057]), .Z(n43500) );
  XOR U43469 ( .A(n43490), .B(n43499), .Z(n43527) );
  XOR U43470 ( .A(n43528), .B(n43496), .Z(n43499) );
  XOR U43471 ( .A(p_input[1351]), .B(p_input[2055]), .Z(n43496) );
  XOR U43472 ( .A(p_input[1352]), .B(n29427), .Z(n43528) );
  XOR U43473 ( .A(p_input[1347]), .B(p_input[2051]), .Z(n43490) );
  XNOR U43474 ( .A(n43505), .B(n43504), .Z(n43495) );
  XOR U43475 ( .A(n43529), .B(n43501), .Z(n43504) );
  XOR U43476 ( .A(p_input[1348]), .B(p_input[2052]), .Z(n43501) );
  XOR U43477 ( .A(p_input[1349]), .B(n29429), .Z(n43529) );
  XOR U43478 ( .A(p_input[1350]), .B(p_input[2054]), .Z(n43505) );
  XNOR U43479 ( .A(n43530), .B(n43531), .Z(n43306) );
  AND U43480 ( .A(n933), .B(n43532), .Z(n43531) );
  XNOR U43481 ( .A(n43533), .B(n43534), .Z(n933) );
  AND U43482 ( .A(n43535), .B(n43536), .Z(n43534) );
  XOR U43483 ( .A(n43320), .B(n43533), .Z(n43536) );
  XNOR U43484 ( .A(n43537), .B(n43533), .Z(n43535) );
  XOR U43485 ( .A(n43538), .B(n43539), .Z(n43533) );
  AND U43486 ( .A(n43540), .B(n43541), .Z(n43539) );
  XOR U43487 ( .A(n43335), .B(n43538), .Z(n43541) );
  XOR U43488 ( .A(n43538), .B(n43336), .Z(n43540) );
  XOR U43489 ( .A(n43542), .B(n43543), .Z(n43538) );
  AND U43490 ( .A(n43544), .B(n43545), .Z(n43543) );
  XOR U43491 ( .A(n43363), .B(n43542), .Z(n43545) );
  XOR U43492 ( .A(n43542), .B(n43364), .Z(n43544) );
  XOR U43493 ( .A(n43546), .B(n43547), .Z(n43542) );
  AND U43494 ( .A(n43548), .B(n43549), .Z(n43547) );
  XOR U43495 ( .A(n43412), .B(n43546), .Z(n43549) );
  XOR U43496 ( .A(n43546), .B(n43413), .Z(n43548) );
  XOR U43497 ( .A(n43550), .B(n43551), .Z(n43546) );
  AND U43498 ( .A(n43552), .B(n43553), .Z(n43551) );
  XOR U43499 ( .A(n43550), .B(n43509), .Z(n43553) );
  XNOR U43500 ( .A(n43554), .B(n43555), .Z(n43256) );
  AND U43501 ( .A(n937), .B(n43556), .Z(n43555) );
  XNOR U43502 ( .A(n43557), .B(n43558), .Z(n937) );
  AND U43503 ( .A(n43559), .B(n43560), .Z(n43558) );
  XOR U43504 ( .A(n43557), .B(n43266), .Z(n43560) );
  XNOR U43505 ( .A(n43557), .B(n43216), .Z(n43559) );
  XOR U43506 ( .A(n43561), .B(n43562), .Z(n43557) );
  AND U43507 ( .A(n43563), .B(n43564), .Z(n43562) );
  XNOR U43508 ( .A(n43276), .B(n43561), .Z(n43564) );
  XOR U43509 ( .A(n43561), .B(n43226), .Z(n43563) );
  XOR U43510 ( .A(n43565), .B(n43566), .Z(n43561) );
  AND U43511 ( .A(n43567), .B(n43568), .Z(n43566) );
  XNOR U43512 ( .A(n43286), .B(n43565), .Z(n43568) );
  XOR U43513 ( .A(n43565), .B(n43235), .Z(n43567) );
  XOR U43514 ( .A(n43569), .B(n43570), .Z(n43565) );
  AND U43515 ( .A(n43571), .B(n43572), .Z(n43570) );
  XOR U43516 ( .A(n43569), .B(n43243), .Z(n43571) );
  XOR U43517 ( .A(n43573), .B(n43574), .Z(n43207) );
  AND U43518 ( .A(n941), .B(n43556), .Z(n43574) );
  XNOR U43519 ( .A(n43554), .B(n43573), .Z(n43556) );
  XNOR U43520 ( .A(n43575), .B(n43576), .Z(n941) );
  AND U43521 ( .A(n43577), .B(n43578), .Z(n43576) );
  XNOR U43522 ( .A(n43579), .B(n43575), .Z(n43578) );
  IV U43523 ( .A(n43266), .Z(n43579) );
  XOR U43524 ( .A(n43537), .B(n43580), .Z(n43266) );
  AND U43525 ( .A(n944), .B(n43581), .Z(n43580) );
  XOR U43526 ( .A(n43319), .B(n43316), .Z(n43581) );
  IV U43527 ( .A(n43537), .Z(n43319) );
  XNOR U43528 ( .A(n43216), .B(n43575), .Z(n43577) );
  XOR U43529 ( .A(n43582), .B(n43583), .Z(n43216) );
  AND U43530 ( .A(n960), .B(n43584), .Z(n43583) );
  XOR U43531 ( .A(n43585), .B(n43586), .Z(n43575) );
  AND U43532 ( .A(n43587), .B(n43588), .Z(n43586) );
  XNOR U43533 ( .A(n43585), .B(n43276), .Z(n43588) );
  XOR U43534 ( .A(n43336), .B(n43589), .Z(n43276) );
  AND U43535 ( .A(n944), .B(n43590), .Z(n43589) );
  XOR U43536 ( .A(n43332), .B(n43336), .Z(n43590) );
  XNOR U43537 ( .A(n43591), .B(n43585), .Z(n43587) );
  IV U43538 ( .A(n43226), .Z(n43591) );
  XOR U43539 ( .A(n43592), .B(n43593), .Z(n43226) );
  AND U43540 ( .A(n960), .B(n43594), .Z(n43593) );
  XOR U43541 ( .A(n43595), .B(n43596), .Z(n43585) );
  AND U43542 ( .A(n43597), .B(n43598), .Z(n43596) );
  XNOR U43543 ( .A(n43595), .B(n43286), .Z(n43598) );
  XOR U43544 ( .A(n43364), .B(n43599), .Z(n43286) );
  AND U43545 ( .A(n944), .B(n43600), .Z(n43599) );
  XOR U43546 ( .A(n43360), .B(n43364), .Z(n43600) );
  XOR U43547 ( .A(n43235), .B(n43595), .Z(n43597) );
  XOR U43548 ( .A(n43601), .B(n43602), .Z(n43235) );
  AND U43549 ( .A(n960), .B(n43603), .Z(n43602) );
  XOR U43550 ( .A(n43569), .B(n43604), .Z(n43595) );
  AND U43551 ( .A(n43605), .B(n43572), .Z(n43604) );
  XNOR U43552 ( .A(n43296), .B(n43569), .Z(n43572) );
  XOR U43553 ( .A(n43413), .B(n43606), .Z(n43296) );
  AND U43554 ( .A(n944), .B(n43607), .Z(n43606) );
  XOR U43555 ( .A(n43409), .B(n43413), .Z(n43607) );
  XNOR U43556 ( .A(n43608), .B(n43569), .Z(n43605) );
  IV U43557 ( .A(n43243), .Z(n43608) );
  XOR U43558 ( .A(n43609), .B(n43610), .Z(n43243) );
  AND U43559 ( .A(n960), .B(n43611), .Z(n43610) );
  XOR U43560 ( .A(n43612), .B(n43613), .Z(n43569) );
  AND U43561 ( .A(n43614), .B(n43615), .Z(n43613) );
  XNOR U43562 ( .A(n43612), .B(n43304), .Z(n43615) );
  XOR U43563 ( .A(n43510), .B(n43616), .Z(n43304) );
  AND U43564 ( .A(n944), .B(n43617), .Z(n43616) );
  XOR U43565 ( .A(n43506), .B(n43510), .Z(n43617) );
  XNOR U43566 ( .A(n43618), .B(n43612), .Z(n43614) );
  IV U43567 ( .A(n43253), .Z(n43618) );
  XOR U43568 ( .A(n43619), .B(n43620), .Z(n43253) );
  AND U43569 ( .A(n960), .B(n43621), .Z(n43620) );
  AND U43570 ( .A(n43573), .B(n43554), .Z(n43612) );
  XNOR U43571 ( .A(n43622), .B(n43623), .Z(n43554) );
  AND U43572 ( .A(n944), .B(n43532), .Z(n43623) );
  XNOR U43573 ( .A(n43530), .B(n43622), .Z(n43532) );
  XNOR U43574 ( .A(n43624), .B(n43625), .Z(n944) );
  AND U43575 ( .A(n43626), .B(n43627), .Z(n43625) );
  XNOR U43576 ( .A(n43624), .B(n43316), .Z(n43627) );
  IV U43577 ( .A(n43320), .Z(n43316) );
  XOR U43578 ( .A(n43628), .B(n43629), .Z(n43320) );
  AND U43579 ( .A(n948), .B(n43630), .Z(n43629) );
  XOR U43580 ( .A(n43631), .B(n43628), .Z(n43630) );
  XNOR U43581 ( .A(n43624), .B(n43537), .Z(n43626) );
  XOR U43582 ( .A(n43632), .B(n43633), .Z(n43537) );
  AND U43583 ( .A(n956), .B(n43584), .Z(n43633) );
  XOR U43584 ( .A(n43582), .B(n43632), .Z(n43584) );
  XOR U43585 ( .A(n43634), .B(n43635), .Z(n43624) );
  AND U43586 ( .A(n43636), .B(n43637), .Z(n43635) );
  XNOR U43587 ( .A(n43634), .B(n43332), .Z(n43637) );
  IV U43588 ( .A(n43335), .Z(n43332) );
  XOR U43589 ( .A(n43638), .B(n43639), .Z(n43335) );
  AND U43590 ( .A(n948), .B(n43640), .Z(n43639) );
  XOR U43591 ( .A(n43641), .B(n43638), .Z(n43640) );
  XOR U43592 ( .A(n43336), .B(n43634), .Z(n43636) );
  XOR U43593 ( .A(n43642), .B(n43643), .Z(n43336) );
  AND U43594 ( .A(n956), .B(n43594), .Z(n43643) );
  XOR U43595 ( .A(n43642), .B(n43592), .Z(n43594) );
  XOR U43596 ( .A(n43644), .B(n43645), .Z(n43634) );
  AND U43597 ( .A(n43646), .B(n43647), .Z(n43645) );
  XNOR U43598 ( .A(n43644), .B(n43360), .Z(n43647) );
  IV U43599 ( .A(n43363), .Z(n43360) );
  XOR U43600 ( .A(n43648), .B(n43649), .Z(n43363) );
  AND U43601 ( .A(n948), .B(n43650), .Z(n43649) );
  XNOR U43602 ( .A(n43651), .B(n43648), .Z(n43650) );
  XOR U43603 ( .A(n43364), .B(n43644), .Z(n43646) );
  XOR U43604 ( .A(n43652), .B(n43653), .Z(n43364) );
  AND U43605 ( .A(n956), .B(n43603), .Z(n43653) );
  XOR U43606 ( .A(n43652), .B(n43601), .Z(n43603) );
  XOR U43607 ( .A(n43654), .B(n43655), .Z(n43644) );
  AND U43608 ( .A(n43656), .B(n43657), .Z(n43655) );
  XNOR U43609 ( .A(n43654), .B(n43409), .Z(n43657) );
  IV U43610 ( .A(n43412), .Z(n43409) );
  XOR U43611 ( .A(n43658), .B(n43659), .Z(n43412) );
  AND U43612 ( .A(n948), .B(n43660), .Z(n43659) );
  XOR U43613 ( .A(n43661), .B(n43658), .Z(n43660) );
  XOR U43614 ( .A(n43413), .B(n43654), .Z(n43656) );
  XOR U43615 ( .A(n43662), .B(n43663), .Z(n43413) );
  AND U43616 ( .A(n956), .B(n43611), .Z(n43663) );
  XOR U43617 ( .A(n43662), .B(n43609), .Z(n43611) );
  XOR U43618 ( .A(n43550), .B(n43664), .Z(n43654) );
  AND U43619 ( .A(n43552), .B(n43665), .Z(n43664) );
  XNOR U43620 ( .A(n43550), .B(n43506), .Z(n43665) );
  IV U43621 ( .A(n43509), .Z(n43506) );
  XOR U43622 ( .A(n43666), .B(n43667), .Z(n43509) );
  AND U43623 ( .A(n948), .B(n43668), .Z(n43667) );
  XNOR U43624 ( .A(n43669), .B(n43666), .Z(n43668) );
  XOR U43625 ( .A(n43510), .B(n43550), .Z(n43552) );
  XOR U43626 ( .A(n43670), .B(n43671), .Z(n43510) );
  AND U43627 ( .A(n956), .B(n43621), .Z(n43671) );
  XOR U43628 ( .A(n43670), .B(n43619), .Z(n43621) );
  AND U43629 ( .A(n43622), .B(n43530), .Z(n43550) );
  XNOR U43630 ( .A(n43672), .B(n43673), .Z(n43530) );
  AND U43631 ( .A(n948), .B(n43674), .Z(n43673) );
  XNOR U43632 ( .A(n43675), .B(n43672), .Z(n43674) );
  XNOR U43633 ( .A(n43676), .B(n43677), .Z(n948) );
  AND U43634 ( .A(n43678), .B(n43679), .Z(n43677) );
  XOR U43635 ( .A(n43631), .B(n43676), .Z(n43679) );
  AND U43636 ( .A(n43680), .B(n43681), .Z(n43631) );
  XNOR U43637 ( .A(n43628), .B(n43676), .Z(n43678) );
  XNOR U43638 ( .A(n43682), .B(n43683), .Z(n43628) );
  AND U43639 ( .A(n952), .B(n43684), .Z(n43683) );
  XNOR U43640 ( .A(n43685), .B(n43686), .Z(n43684) );
  XOR U43641 ( .A(n43687), .B(n43688), .Z(n43676) );
  AND U43642 ( .A(n43689), .B(n43690), .Z(n43688) );
  XNOR U43643 ( .A(n43687), .B(n43680), .Z(n43690) );
  IV U43644 ( .A(n43641), .Z(n43680) );
  XOR U43645 ( .A(n43691), .B(n43692), .Z(n43641) );
  XOR U43646 ( .A(n43693), .B(n43681), .Z(n43692) );
  AND U43647 ( .A(n43651), .B(n43694), .Z(n43681) );
  AND U43648 ( .A(n43695), .B(n43696), .Z(n43693) );
  XOR U43649 ( .A(n43697), .B(n43691), .Z(n43695) );
  XNOR U43650 ( .A(n43638), .B(n43687), .Z(n43689) );
  XNOR U43651 ( .A(n43698), .B(n43699), .Z(n43638) );
  AND U43652 ( .A(n952), .B(n43700), .Z(n43699) );
  XNOR U43653 ( .A(n43701), .B(n43702), .Z(n43700) );
  XOR U43654 ( .A(n43703), .B(n43704), .Z(n43687) );
  AND U43655 ( .A(n43705), .B(n43706), .Z(n43704) );
  XNOR U43656 ( .A(n43703), .B(n43651), .Z(n43706) );
  XOR U43657 ( .A(n43707), .B(n43696), .Z(n43651) );
  XNOR U43658 ( .A(n43708), .B(n43691), .Z(n43696) );
  XOR U43659 ( .A(n43709), .B(n43710), .Z(n43691) );
  AND U43660 ( .A(n43711), .B(n43712), .Z(n43710) );
  XOR U43661 ( .A(n43713), .B(n43709), .Z(n43711) );
  XNOR U43662 ( .A(n43714), .B(n43715), .Z(n43708) );
  AND U43663 ( .A(n43716), .B(n43717), .Z(n43715) );
  XOR U43664 ( .A(n43714), .B(n43718), .Z(n43716) );
  XNOR U43665 ( .A(n43697), .B(n43694), .Z(n43707) );
  AND U43666 ( .A(n43719), .B(n43720), .Z(n43694) );
  XOR U43667 ( .A(n43721), .B(n43722), .Z(n43697) );
  AND U43668 ( .A(n43723), .B(n43724), .Z(n43722) );
  XOR U43669 ( .A(n43721), .B(n43725), .Z(n43723) );
  XNOR U43670 ( .A(n43648), .B(n43703), .Z(n43705) );
  XNOR U43671 ( .A(n43726), .B(n43727), .Z(n43648) );
  AND U43672 ( .A(n952), .B(n43728), .Z(n43727) );
  XNOR U43673 ( .A(n43729), .B(n43730), .Z(n43728) );
  XOR U43674 ( .A(n43731), .B(n43732), .Z(n43703) );
  AND U43675 ( .A(n43733), .B(n43734), .Z(n43732) );
  XNOR U43676 ( .A(n43731), .B(n43719), .Z(n43734) );
  IV U43677 ( .A(n43661), .Z(n43719) );
  XNOR U43678 ( .A(n43735), .B(n43712), .Z(n43661) );
  XNOR U43679 ( .A(n43736), .B(n43718), .Z(n43712) );
  XOR U43680 ( .A(n43737), .B(n43738), .Z(n43718) );
  AND U43681 ( .A(n43739), .B(n43740), .Z(n43738) );
  XOR U43682 ( .A(n43737), .B(n43741), .Z(n43739) );
  XNOR U43683 ( .A(n43717), .B(n43709), .Z(n43736) );
  XOR U43684 ( .A(n43742), .B(n43743), .Z(n43709) );
  AND U43685 ( .A(n43744), .B(n43745), .Z(n43743) );
  XNOR U43686 ( .A(n43746), .B(n43742), .Z(n43744) );
  XNOR U43687 ( .A(n43747), .B(n43714), .Z(n43717) );
  XOR U43688 ( .A(n43748), .B(n43749), .Z(n43714) );
  AND U43689 ( .A(n43750), .B(n43751), .Z(n43749) );
  XOR U43690 ( .A(n43748), .B(n43752), .Z(n43750) );
  XNOR U43691 ( .A(n43753), .B(n43754), .Z(n43747) );
  AND U43692 ( .A(n43755), .B(n43756), .Z(n43754) );
  XNOR U43693 ( .A(n43753), .B(n43757), .Z(n43755) );
  XNOR U43694 ( .A(n43713), .B(n43720), .Z(n43735) );
  AND U43695 ( .A(n43669), .B(n43758), .Z(n43720) );
  XOR U43696 ( .A(n43725), .B(n43724), .Z(n43713) );
  XNOR U43697 ( .A(n43759), .B(n43721), .Z(n43724) );
  XOR U43698 ( .A(n43760), .B(n43761), .Z(n43721) );
  AND U43699 ( .A(n43762), .B(n43763), .Z(n43761) );
  XOR U43700 ( .A(n43760), .B(n43764), .Z(n43762) );
  XNOR U43701 ( .A(n43765), .B(n43766), .Z(n43759) );
  AND U43702 ( .A(n43767), .B(n43768), .Z(n43766) );
  XOR U43703 ( .A(n43765), .B(n43769), .Z(n43767) );
  XOR U43704 ( .A(n43770), .B(n43771), .Z(n43725) );
  AND U43705 ( .A(n43772), .B(n43773), .Z(n43771) );
  XOR U43706 ( .A(n43770), .B(n43774), .Z(n43772) );
  XNOR U43707 ( .A(n43658), .B(n43731), .Z(n43733) );
  XNOR U43708 ( .A(n43775), .B(n43776), .Z(n43658) );
  AND U43709 ( .A(n952), .B(n43777), .Z(n43776) );
  XNOR U43710 ( .A(n43778), .B(n43779), .Z(n43777) );
  XOR U43711 ( .A(n43780), .B(n43781), .Z(n43731) );
  AND U43712 ( .A(n43782), .B(n43783), .Z(n43781) );
  XNOR U43713 ( .A(n43780), .B(n43669), .Z(n43783) );
  XOR U43714 ( .A(n43784), .B(n43745), .Z(n43669) );
  XNOR U43715 ( .A(n43785), .B(n43752), .Z(n43745) );
  XOR U43716 ( .A(n43741), .B(n43740), .Z(n43752) );
  XNOR U43717 ( .A(n43786), .B(n43737), .Z(n43740) );
  XOR U43718 ( .A(n43787), .B(n43788), .Z(n43737) );
  AND U43719 ( .A(n43789), .B(n43790), .Z(n43788) );
  XNOR U43720 ( .A(n43791), .B(n43792), .Z(n43789) );
  IV U43721 ( .A(n43787), .Z(n43791) );
  XNOR U43722 ( .A(n43793), .B(n43794), .Z(n43786) );
  NOR U43723 ( .A(n43795), .B(n43796), .Z(n43794) );
  XNOR U43724 ( .A(n43793), .B(n43797), .Z(n43795) );
  XOR U43725 ( .A(n43798), .B(n43799), .Z(n43741) );
  NOR U43726 ( .A(n43800), .B(n43801), .Z(n43799) );
  XNOR U43727 ( .A(n43798), .B(n43802), .Z(n43800) );
  XNOR U43728 ( .A(n43751), .B(n43742), .Z(n43785) );
  XOR U43729 ( .A(n43803), .B(n43804), .Z(n43742) );
  AND U43730 ( .A(n43805), .B(n43806), .Z(n43804) );
  XOR U43731 ( .A(n43803), .B(n43807), .Z(n43805) );
  XOR U43732 ( .A(n43808), .B(n43757), .Z(n43751) );
  XOR U43733 ( .A(n43809), .B(n43810), .Z(n43757) );
  NOR U43734 ( .A(n43811), .B(n43812), .Z(n43810) );
  XOR U43735 ( .A(n43809), .B(n43813), .Z(n43811) );
  XNOR U43736 ( .A(n43756), .B(n43748), .Z(n43808) );
  XOR U43737 ( .A(n43814), .B(n43815), .Z(n43748) );
  AND U43738 ( .A(n43816), .B(n43817), .Z(n43815) );
  XOR U43739 ( .A(n43814), .B(n43818), .Z(n43816) );
  XNOR U43740 ( .A(n43819), .B(n43753), .Z(n43756) );
  XOR U43741 ( .A(n43820), .B(n43821), .Z(n43753) );
  AND U43742 ( .A(n43822), .B(n43823), .Z(n43821) );
  XNOR U43743 ( .A(n43824), .B(n43825), .Z(n43822) );
  IV U43744 ( .A(n43820), .Z(n43824) );
  XNOR U43745 ( .A(n43826), .B(n43827), .Z(n43819) );
  NOR U43746 ( .A(n43828), .B(n43829), .Z(n43827) );
  XNOR U43747 ( .A(n43826), .B(n43830), .Z(n43828) );
  XOR U43748 ( .A(n43746), .B(n43758), .Z(n43784) );
  NOR U43749 ( .A(n43675), .B(n43831), .Z(n43758) );
  XNOR U43750 ( .A(n43764), .B(n43763), .Z(n43746) );
  XNOR U43751 ( .A(n43832), .B(n43769), .Z(n43763) );
  XNOR U43752 ( .A(n43833), .B(n43834), .Z(n43769) );
  NOR U43753 ( .A(n43835), .B(n43836), .Z(n43834) );
  XOR U43754 ( .A(n43833), .B(n43837), .Z(n43835) );
  XNOR U43755 ( .A(n43768), .B(n43760), .Z(n43832) );
  XOR U43756 ( .A(n43838), .B(n43839), .Z(n43760) );
  AND U43757 ( .A(n43840), .B(n43841), .Z(n43839) );
  XOR U43758 ( .A(n43838), .B(n43842), .Z(n43840) );
  XNOR U43759 ( .A(n43843), .B(n43765), .Z(n43768) );
  XOR U43760 ( .A(n43844), .B(n43845), .Z(n43765) );
  AND U43761 ( .A(n43846), .B(n43847), .Z(n43845) );
  XNOR U43762 ( .A(n43848), .B(n43849), .Z(n43846) );
  IV U43763 ( .A(n43844), .Z(n43848) );
  XNOR U43764 ( .A(n43850), .B(n43851), .Z(n43843) );
  NOR U43765 ( .A(n43852), .B(n43853), .Z(n43851) );
  XNOR U43766 ( .A(n43850), .B(n43854), .Z(n43852) );
  XOR U43767 ( .A(n43774), .B(n43773), .Z(n43764) );
  XNOR U43768 ( .A(n43855), .B(n43770), .Z(n43773) );
  XOR U43769 ( .A(n43856), .B(n43857), .Z(n43770) );
  AND U43770 ( .A(n43858), .B(n43859), .Z(n43857) );
  XNOR U43771 ( .A(n43860), .B(n43861), .Z(n43858) );
  IV U43772 ( .A(n43856), .Z(n43860) );
  XNOR U43773 ( .A(n43862), .B(n43863), .Z(n43855) );
  NOR U43774 ( .A(n43864), .B(n43865), .Z(n43863) );
  XNOR U43775 ( .A(n43862), .B(n43866), .Z(n43864) );
  XOR U43776 ( .A(n43867), .B(n43868), .Z(n43774) );
  NOR U43777 ( .A(n43869), .B(n43870), .Z(n43868) );
  XNOR U43778 ( .A(n43867), .B(n43871), .Z(n43869) );
  XNOR U43779 ( .A(n43666), .B(n43780), .Z(n43782) );
  XNOR U43780 ( .A(n43872), .B(n43873), .Z(n43666) );
  AND U43781 ( .A(n952), .B(n43874), .Z(n43873) );
  XNOR U43782 ( .A(n43875), .B(n43876), .Z(n43874) );
  AND U43783 ( .A(n43672), .B(n43675), .Z(n43780) );
  XOR U43784 ( .A(n43877), .B(n43831), .Z(n43675) );
  XNOR U43785 ( .A(p_input[1376]), .B(p_input[2048]), .Z(n43831) );
  XNOR U43786 ( .A(n43807), .B(n43806), .Z(n43877) );
  XNOR U43787 ( .A(n43878), .B(n43818), .Z(n43806) );
  XOR U43788 ( .A(n43792), .B(n43790), .Z(n43818) );
  XNOR U43789 ( .A(n43879), .B(n43797), .Z(n43790) );
  XOR U43790 ( .A(p_input[1400]), .B(p_input[2072]), .Z(n43797) );
  XOR U43791 ( .A(n43787), .B(n43796), .Z(n43879) );
  XOR U43792 ( .A(n43880), .B(n43793), .Z(n43796) );
  XOR U43793 ( .A(p_input[1398]), .B(p_input[2070]), .Z(n43793) );
  XOR U43794 ( .A(p_input[1399]), .B(n29410), .Z(n43880) );
  XOR U43795 ( .A(p_input[1394]), .B(p_input[2066]), .Z(n43787) );
  XNOR U43796 ( .A(n43802), .B(n43801), .Z(n43792) );
  XOR U43797 ( .A(n43881), .B(n43798), .Z(n43801) );
  XOR U43798 ( .A(p_input[1395]), .B(p_input[2067]), .Z(n43798) );
  XOR U43799 ( .A(p_input[1396]), .B(n29412), .Z(n43881) );
  XOR U43800 ( .A(p_input[1397]), .B(p_input[2069]), .Z(n43802) );
  XOR U43801 ( .A(n43817), .B(n43882), .Z(n43878) );
  IV U43802 ( .A(n43803), .Z(n43882) );
  XOR U43803 ( .A(p_input[1377]), .B(p_input[2049]), .Z(n43803) );
  XNOR U43804 ( .A(n43883), .B(n43825), .Z(n43817) );
  XNOR U43805 ( .A(n43813), .B(n43812), .Z(n43825) );
  XNOR U43806 ( .A(n43884), .B(n43809), .Z(n43812) );
  XNOR U43807 ( .A(p_input[1402]), .B(p_input[2074]), .Z(n43809) );
  XOR U43808 ( .A(p_input[1403]), .B(n29415), .Z(n43884) );
  XOR U43809 ( .A(p_input[1404]), .B(p_input[2076]), .Z(n43813) );
  XOR U43810 ( .A(n43823), .B(n43885), .Z(n43883) );
  IV U43811 ( .A(n43814), .Z(n43885) );
  XOR U43812 ( .A(p_input[1393]), .B(p_input[2065]), .Z(n43814) );
  XNOR U43813 ( .A(n43886), .B(n43830), .Z(n43823) );
  XNOR U43814 ( .A(p_input[1407]), .B(n29418), .Z(n43830) );
  XOR U43815 ( .A(n43820), .B(n43829), .Z(n43886) );
  XOR U43816 ( .A(n43887), .B(n43826), .Z(n43829) );
  XOR U43817 ( .A(p_input[1405]), .B(p_input[2077]), .Z(n43826) );
  XOR U43818 ( .A(p_input[1406]), .B(n29420), .Z(n43887) );
  XOR U43819 ( .A(p_input[1401]), .B(p_input[2073]), .Z(n43820) );
  XOR U43820 ( .A(n43842), .B(n43841), .Z(n43807) );
  XNOR U43821 ( .A(n43888), .B(n43849), .Z(n43841) );
  XNOR U43822 ( .A(n43837), .B(n43836), .Z(n43849) );
  XNOR U43823 ( .A(n43889), .B(n43833), .Z(n43836) );
  XNOR U43824 ( .A(p_input[1387]), .B(p_input[2059]), .Z(n43833) );
  XOR U43825 ( .A(p_input[1388]), .B(n28329), .Z(n43889) );
  XOR U43826 ( .A(p_input[1389]), .B(p_input[2061]), .Z(n43837) );
  XOR U43827 ( .A(n43847), .B(n43890), .Z(n43888) );
  IV U43828 ( .A(n43838), .Z(n43890) );
  XOR U43829 ( .A(p_input[1378]), .B(p_input[2050]), .Z(n43838) );
  XNOR U43830 ( .A(n43891), .B(n43854), .Z(n43847) );
  XNOR U43831 ( .A(p_input[1392]), .B(n28332), .Z(n43854) );
  XOR U43832 ( .A(n43844), .B(n43853), .Z(n43891) );
  XOR U43833 ( .A(n43892), .B(n43850), .Z(n43853) );
  XOR U43834 ( .A(p_input[1390]), .B(p_input[2062]), .Z(n43850) );
  XOR U43835 ( .A(p_input[1391]), .B(n28334), .Z(n43892) );
  XOR U43836 ( .A(p_input[1386]), .B(p_input[2058]), .Z(n43844) );
  XOR U43837 ( .A(n43861), .B(n43859), .Z(n43842) );
  XNOR U43838 ( .A(n43893), .B(n43866), .Z(n43859) );
  XOR U43839 ( .A(p_input[1385]), .B(p_input[2057]), .Z(n43866) );
  XOR U43840 ( .A(n43856), .B(n43865), .Z(n43893) );
  XOR U43841 ( .A(n43894), .B(n43862), .Z(n43865) );
  XOR U43842 ( .A(p_input[1383]), .B(p_input[2055]), .Z(n43862) );
  XOR U43843 ( .A(p_input[1384]), .B(n29427), .Z(n43894) );
  XOR U43844 ( .A(p_input[1379]), .B(p_input[2051]), .Z(n43856) );
  XNOR U43845 ( .A(n43871), .B(n43870), .Z(n43861) );
  XOR U43846 ( .A(n43895), .B(n43867), .Z(n43870) );
  XOR U43847 ( .A(p_input[1380]), .B(p_input[2052]), .Z(n43867) );
  XOR U43848 ( .A(p_input[1381]), .B(n29429), .Z(n43895) );
  XOR U43849 ( .A(p_input[1382]), .B(p_input[2054]), .Z(n43871) );
  XNOR U43850 ( .A(n43896), .B(n43897), .Z(n43672) );
  AND U43851 ( .A(n952), .B(n43898), .Z(n43897) );
  XNOR U43852 ( .A(n43899), .B(n43900), .Z(n952) );
  AND U43853 ( .A(n43901), .B(n43902), .Z(n43900) );
  XOR U43854 ( .A(n43686), .B(n43899), .Z(n43902) );
  XNOR U43855 ( .A(n43903), .B(n43899), .Z(n43901) );
  XOR U43856 ( .A(n43904), .B(n43905), .Z(n43899) );
  AND U43857 ( .A(n43906), .B(n43907), .Z(n43905) );
  XOR U43858 ( .A(n43701), .B(n43904), .Z(n43907) );
  XOR U43859 ( .A(n43904), .B(n43702), .Z(n43906) );
  XOR U43860 ( .A(n43908), .B(n43909), .Z(n43904) );
  AND U43861 ( .A(n43910), .B(n43911), .Z(n43909) );
  XOR U43862 ( .A(n43729), .B(n43908), .Z(n43911) );
  XOR U43863 ( .A(n43908), .B(n43730), .Z(n43910) );
  XOR U43864 ( .A(n43912), .B(n43913), .Z(n43908) );
  AND U43865 ( .A(n43914), .B(n43915), .Z(n43913) );
  XOR U43866 ( .A(n43778), .B(n43912), .Z(n43915) );
  XOR U43867 ( .A(n43912), .B(n43779), .Z(n43914) );
  XOR U43868 ( .A(n43916), .B(n43917), .Z(n43912) );
  AND U43869 ( .A(n43918), .B(n43919), .Z(n43917) );
  XOR U43870 ( .A(n43916), .B(n43875), .Z(n43919) );
  XNOR U43871 ( .A(n43920), .B(n43921), .Z(n43622) );
  AND U43872 ( .A(n956), .B(n43922), .Z(n43921) );
  XNOR U43873 ( .A(n43923), .B(n43924), .Z(n956) );
  AND U43874 ( .A(n43925), .B(n43926), .Z(n43924) );
  XOR U43875 ( .A(n43923), .B(n43632), .Z(n43926) );
  XNOR U43876 ( .A(n43923), .B(n43582), .Z(n43925) );
  XOR U43877 ( .A(n43927), .B(n43928), .Z(n43923) );
  AND U43878 ( .A(n43929), .B(n43930), .Z(n43928) );
  XNOR U43879 ( .A(n43642), .B(n43927), .Z(n43930) );
  XOR U43880 ( .A(n43927), .B(n43592), .Z(n43929) );
  XOR U43881 ( .A(n43931), .B(n43932), .Z(n43927) );
  AND U43882 ( .A(n43933), .B(n43934), .Z(n43932) );
  XNOR U43883 ( .A(n43652), .B(n43931), .Z(n43934) );
  XOR U43884 ( .A(n43931), .B(n43601), .Z(n43933) );
  XOR U43885 ( .A(n43935), .B(n43936), .Z(n43931) );
  AND U43886 ( .A(n43937), .B(n43938), .Z(n43936) );
  XOR U43887 ( .A(n43935), .B(n43609), .Z(n43937) );
  XOR U43888 ( .A(n43939), .B(n43940), .Z(n43573) );
  AND U43889 ( .A(n960), .B(n43922), .Z(n43940) );
  XNOR U43890 ( .A(n43920), .B(n43939), .Z(n43922) );
  XNOR U43891 ( .A(n43941), .B(n43942), .Z(n960) );
  AND U43892 ( .A(n43943), .B(n43944), .Z(n43942) );
  XNOR U43893 ( .A(n43945), .B(n43941), .Z(n43944) );
  IV U43894 ( .A(n43632), .Z(n43945) );
  XOR U43895 ( .A(n43903), .B(n43946), .Z(n43632) );
  AND U43896 ( .A(n963), .B(n43947), .Z(n43946) );
  XOR U43897 ( .A(n43685), .B(n43682), .Z(n43947) );
  IV U43898 ( .A(n43903), .Z(n43685) );
  XNOR U43899 ( .A(n43582), .B(n43941), .Z(n43943) );
  XOR U43900 ( .A(n43948), .B(n43949), .Z(n43582) );
  AND U43901 ( .A(n979), .B(n43950), .Z(n43949) );
  XOR U43902 ( .A(n43951), .B(n43952), .Z(n43941) );
  AND U43903 ( .A(n43953), .B(n43954), .Z(n43952) );
  XNOR U43904 ( .A(n43951), .B(n43642), .Z(n43954) );
  XOR U43905 ( .A(n43702), .B(n43955), .Z(n43642) );
  AND U43906 ( .A(n963), .B(n43956), .Z(n43955) );
  XOR U43907 ( .A(n43698), .B(n43702), .Z(n43956) );
  XNOR U43908 ( .A(n43957), .B(n43951), .Z(n43953) );
  IV U43909 ( .A(n43592), .Z(n43957) );
  XOR U43910 ( .A(n43958), .B(n43959), .Z(n43592) );
  AND U43911 ( .A(n979), .B(n43960), .Z(n43959) );
  XOR U43912 ( .A(n43961), .B(n43962), .Z(n43951) );
  AND U43913 ( .A(n43963), .B(n43964), .Z(n43962) );
  XNOR U43914 ( .A(n43961), .B(n43652), .Z(n43964) );
  XOR U43915 ( .A(n43730), .B(n43965), .Z(n43652) );
  AND U43916 ( .A(n963), .B(n43966), .Z(n43965) );
  XOR U43917 ( .A(n43726), .B(n43730), .Z(n43966) );
  XOR U43918 ( .A(n43601), .B(n43961), .Z(n43963) );
  XOR U43919 ( .A(n43967), .B(n43968), .Z(n43601) );
  AND U43920 ( .A(n979), .B(n43969), .Z(n43968) );
  XOR U43921 ( .A(n43935), .B(n43970), .Z(n43961) );
  AND U43922 ( .A(n43971), .B(n43938), .Z(n43970) );
  XNOR U43923 ( .A(n43662), .B(n43935), .Z(n43938) );
  XOR U43924 ( .A(n43779), .B(n43972), .Z(n43662) );
  AND U43925 ( .A(n963), .B(n43973), .Z(n43972) );
  XOR U43926 ( .A(n43775), .B(n43779), .Z(n43973) );
  XNOR U43927 ( .A(n43974), .B(n43935), .Z(n43971) );
  IV U43928 ( .A(n43609), .Z(n43974) );
  XOR U43929 ( .A(n43975), .B(n43976), .Z(n43609) );
  AND U43930 ( .A(n979), .B(n43977), .Z(n43976) );
  XOR U43931 ( .A(n43978), .B(n43979), .Z(n43935) );
  AND U43932 ( .A(n43980), .B(n43981), .Z(n43979) );
  XNOR U43933 ( .A(n43978), .B(n43670), .Z(n43981) );
  XOR U43934 ( .A(n43876), .B(n43982), .Z(n43670) );
  AND U43935 ( .A(n963), .B(n43983), .Z(n43982) );
  XOR U43936 ( .A(n43872), .B(n43876), .Z(n43983) );
  XNOR U43937 ( .A(n43984), .B(n43978), .Z(n43980) );
  IV U43938 ( .A(n43619), .Z(n43984) );
  XOR U43939 ( .A(n43985), .B(n43986), .Z(n43619) );
  AND U43940 ( .A(n979), .B(n43987), .Z(n43986) );
  AND U43941 ( .A(n43939), .B(n43920), .Z(n43978) );
  XNOR U43942 ( .A(n43988), .B(n43989), .Z(n43920) );
  AND U43943 ( .A(n963), .B(n43898), .Z(n43989) );
  XNOR U43944 ( .A(n43896), .B(n43988), .Z(n43898) );
  XNOR U43945 ( .A(n43990), .B(n43991), .Z(n963) );
  AND U43946 ( .A(n43992), .B(n43993), .Z(n43991) );
  XNOR U43947 ( .A(n43990), .B(n43682), .Z(n43993) );
  IV U43948 ( .A(n43686), .Z(n43682) );
  XOR U43949 ( .A(n43994), .B(n43995), .Z(n43686) );
  AND U43950 ( .A(n967), .B(n43996), .Z(n43995) );
  XOR U43951 ( .A(n43997), .B(n43994), .Z(n43996) );
  XNOR U43952 ( .A(n43990), .B(n43903), .Z(n43992) );
  XOR U43953 ( .A(n43998), .B(n43999), .Z(n43903) );
  AND U43954 ( .A(n975), .B(n43950), .Z(n43999) );
  XOR U43955 ( .A(n43948), .B(n43998), .Z(n43950) );
  XOR U43956 ( .A(n44000), .B(n44001), .Z(n43990) );
  AND U43957 ( .A(n44002), .B(n44003), .Z(n44001) );
  XNOR U43958 ( .A(n44000), .B(n43698), .Z(n44003) );
  IV U43959 ( .A(n43701), .Z(n43698) );
  XOR U43960 ( .A(n44004), .B(n44005), .Z(n43701) );
  AND U43961 ( .A(n967), .B(n44006), .Z(n44005) );
  XOR U43962 ( .A(n44007), .B(n44004), .Z(n44006) );
  XOR U43963 ( .A(n43702), .B(n44000), .Z(n44002) );
  XOR U43964 ( .A(n44008), .B(n44009), .Z(n43702) );
  AND U43965 ( .A(n975), .B(n43960), .Z(n44009) );
  XOR U43966 ( .A(n44008), .B(n43958), .Z(n43960) );
  XOR U43967 ( .A(n44010), .B(n44011), .Z(n44000) );
  AND U43968 ( .A(n44012), .B(n44013), .Z(n44011) );
  XNOR U43969 ( .A(n44010), .B(n43726), .Z(n44013) );
  IV U43970 ( .A(n43729), .Z(n43726) );
  XOR U43971 ( .A(n44014), .B(n44015), .Z(n43729) );
  AND U43972 ( .A(n967), .B(n44016), .Z(n44015) );
  XNOR U43973 ( .A(n44017), .B(n44014), .Z(n44016) );
  XOR U43974 ( .A(n43730), .B(n44010), .Z(n44012) );
  XOR U43975 ( .A(n44018), .B(n44019), .Z(n43730) );
  AND U43976 ( .A(n975), .B(n43969), .Z(n44019) );
  XOR U43977 ( .A(n44018), .B(n43967), .Z(n43969) );
  XOR U43978 ( .A(n44020), .B(n44021), .Z(n44010) );
  AND U43979 ( .A(n44022), .B(n44023), .Z(n44021) );
  XNOR U43980 ( .A(n44020), .B(n43775), .Z(n44023) );
  IV U43981 ( .A(n43778), .Z(n43775) );
  XOR U43982 ( .A(n44024), .B(n44025), .Z(n43778) );
  AND U43983 ( .A(n967), .B(n44026), .Z(n44025) );
  XOR U43984 ( .A(n44027), .B(n44024), .Z(n44026) );
  XOR U43985 ( .A(n43779), .B(n44020), .Z(n44022) );
  XOR U43986 ( .A(n44028), .B(n44029), .Z(n43779) );
  AND U43987 ( .A(n975), .B(n43977), .Z(n44029) );
  XOR U43988 ( .A(n44028), .B(n43975), .Z(n43977) );
  XOR U43989 ( .A(n43916), .B(n44030), .Z(n44020) );
  AND U43990 ( .A(n43918), .B(n44031), .Z(n44030) );
  XNOR U43991 ( .A(n43916), .B(n43872), .Z(n44031) );
  IV U43992 ( .A(n43875), .Z(n43872) );
  XOR U43993 ( .A(n44032), .B(n44033), .Z(n43875) );
  AND U43994 ( .A(n967), .B(n44034), .Z(n44033) );
  XNOR U43995 ( .A(n44035), .B(n44032), .Z(n44034) );
  XOR U43996 ( .A(n43876), .B(n43916), .Z(n43918) );
  XOR U43997 ( .A(n44036), .B(n44037), .Z(n43876) );
  AND U43998 ( .A(n975), .B(n43987), .Z(n44037) );
  XOR U43999 ( .A(n44036), .B(n43985), .Z(n43987) );
  AND U44000 ( .A(n43988), .B(n43896), .Z(n43916) );
  XNOR U44001 ( .A(n44038), .B(n44039), .Z(n43896) );
  AND U44002 ( .A(n967), .B(n44040), .Z(n44039) );
  XNOR U44003 ( .A(n44041), .B(n44038), .Z(n44040) );
  XNOR U44004 ( .A(n44042), .B(n44043), .Z(n967) );
  AND U44005 ( .A(n44044), .B(n44045), .Z(n44043) );
  XOR U44006 ( .A(n43997), .B(n44042), .Z(n44045) );
  AND U44007 ( .A(n44046), .B(n44047), .Z(n43997) );
  XNOR U44008 ( .A(n43994), .B(n44042), .Z(n44044) );
  XNOR U44009 ( .A(n44048), .B(n44049), .Z(n43994) );
  AND U44010 ( .A(n971), .B(n44050), .Z(n44049) );
  XNOR U44011 ( .A(n44051), .B(n44052), .Z(n44050) );
  XOR U44012 ( .A(n44053), .B(n44054), .Z(n44042) );
  AND U44013 ( .A(n44055), .B(n44056), .Z(n44054) );
  XNOR U44014 ( .A(n44053), .B(n44046), .Z(n44056) );
  IV U44015 ( .A(n44007), .Z(n44046) );
  XOR U44016 ( .A(n44057), .B(n44058), .Z(n44007) );
  XOR U44017 ( .A(n44059), .B(n44047), .Z(n44058) );
  AND U44018 ( .A(n44017), .B(n44060), .Z(n44047) );
  AND U44019 ( .A(n44061), .B(n44062), .Z(n44059) );
  XOR U44020 ( .A(n44063), .B(n44057), .Z(n44061) );
  XNOR U44021 ( .A(n44004), .B(n44053), .Z(n44055) );
  XNOR U44022 ( .A(n44064), .B(n44065), .Z(n44004) );
  AND U44023 ( .A(n971), .B(n44066), .Z(n44065) );
  XNOR U44024 ( .A(n44067), .B(n44068), .Z(n44066) );
  XOR U44025 ( .A(n44069), .B(n44070), .Z(n44053) );
  AND U44026 ( .A(n44071), .B(n44072), .Z(n44070) );
  XNOR U44027 ( .A(n44069), .B(n44017), .Z(n44072) );
  XOR U44028 ( .A(n44073), .B(n44062), .Z(n44017) );
  XNOR U44029 ( .A(n44074), .B(n44057), .Z(n44062) );
  XOR U44030 ( .A(n44075), .B(n44076), .Z(n44057) );
  AND U44031 ( .A(n44077), .B(n44078), .Z(n44076) );
  XOR U44032 ( .A(n44079), .B(n44075), .Z(n44077) );
  XNOR U44033 ( .A(n44080), .B(n44081), .Z(n44074) );
  AND U44034 ( .A(n44082), .B(n44083), .Z(n44081) );
  XOR U44035 ( .A(n44080), .B(n44084), .Z(n44082) );
  XNOR U44036 ( .A(n44063), .B(n44060), .Z(n44073) );
  AND U44037 ( .A(n44085), .B(n44086), .Z(n44060) );
  XOR U44038 ( .A(n44087), .B(n44088), .Z(n44063) );
  AND U44039 ( .A(n44089), .B(n44090), .Z(n44088) );
  XOR U44040 ( .A(n44087), .B(n44091), .Z(n44089) );
  XNOR U44041 ( .A(n44014), .B(n44069), .Z(n44071) );
  XNOR U44042 ( .A(n44092), .B(n44093), .Z(n44014) );
  AND U44043 ( .A(n971), .B(n44094), .Z(n44093) );
  XNOR U44044 ( .A(n44095), .B(n44096), .Z(n44094) );
  XOR U44045 ( .A(n44097), .B(n44098), .Z(n44069) );
  AND U44046 ( .A(n44099), .B(n44100), .Z(n44098) );
  XNOR U44047 ( .A(n44097), .B(n44085), .Z(n44100) );
  IV U44048 ( .A(n44027), .Z(n44085) );
  XNOR U44049 ( .A(n44101), .B(n44078), .Z(n44027) );
  XNOR U44050 ( .A(n44102), .B(n44084), .Z(n44078) );
  XOR U44051 ( .A(n44103), .B(n44104), .Z(n44084) );
  AND U44052 ( .A(n44105), .B(n44106), .Z(n44104) );
  XOR U44053 ( .A(n44103), .B(n44107), .Z(n44105) );
  XNOR U44054 ( .A(n44083), .B(n44075), .Z(n44102) );
  XOR U44055 ( .A(n44108), .B(n44109), .Z(n44075) );
  AND U44056 ( .A(n44110), .B(n44111), .Z(n44109) );
  XNOR U44057 ( .A(n44112), .B(n44108), .Z(n44110) );
  XNOR U44058 ( .A(n44113), .B(n44080), .Z(n44083) );
  XOR U44059 ( .A(n44114), .B(n44115), .Z(n44080) );
  AND U44060 ( .A(n44116), .B(n44117), .Z(n44115) );
  XOR U44061 ( .A(n44114), .B(n44118), .Z(n44116) );
  XNOR U44062 ( .A(n44119), .B(n44120), .Z(n44113) );
  AND U44063 ( .A(n44121), .B(n44122), .Z(n44120) );
  XNOR U44064 ( .A(n44119), .B(n44123), .Z(n44121) );
  XNOR U44065 ( .A(n44079), .B(n44086), .Z(n44101) );
  AND U44066 ( .A(n44035), .B(n44124), .Z(n44086) );
  XOR U44067 ( .A(n44091), .B(n44090), .Z(n44079) );
  XNOR U44068 ( .A(n44125), .B(n44087), .Z(n44090) );
  XOR U44069 ( .A(n44126), .B(n44127), .Z(n44087) );
  AND U44070 ( .A(n44128), .B(n44129), .Z(n44127) );
  XOR U44071 ( .A(n44126), .B(n44130), .Z(n44128) );
  XNOR U44072 ( .A(n44131), .B(n44132), .Z(n44125) );
  AND U44073 ( .A(n44133), .B(n44134), .Z(n44132) );
  XOR U44074 ( .A(n44131), .B(n44135), .Z(n44133) );
  XOR U44075 ( .A(n44136), .B(n44137), .Z(n44091) );
  AND U44076 ( .A(n44138), .B(n44139), .Z(n44137) );
  XOR U44077 ( .A(n44136), .B(n44140), .Z(n44138) );
  XNOR U44078 ( .A(n44024), .B(n44097), .Z(n44099) );
  XNOR U44079 ( .A(n44141), .B(n44142), .Z(n44024) );
  AND U44080 ( .A(n971), .B(n44143), .Z(n44142) );
  XNOR U44081 ( .A(n44144), .B(n44145), .Z(n44143) );
  XOR U44082 ( .A(n44146), .B(n44147), .Z(n44097) );
  AND U44083 ( .A(n44148), .B(n44149), .Z(n44147) );
  XNOR U44084 ( .A(n44146), .B(n44035), .Z(n44149) );
  XOR U44085 ( .A(n44150), .B(n44111), .Z(n44035) );
  XNOR U44086 ( .A(n44151), .B(n44118), .Z(n44111) );
  XOR U44087 ( .A(n44107), .B(n44106), .Z(n44118) );
  XNOR U44088 ( .A(n44152), .B(n44103), .Z(n44106) );
  XOR U44089 ( .A(n44153), .B(n44154), .Z(n44103) );
  AND U44090 ( .A(n44155), .B(n44156), .Z(n44154) );
  XNOR U44091 ( .A(n44157), .B(n44158), .Z(n44155) );
  IV U44092 ( .A(n44153), .Z(n44157) );
  XNOR U44093 ( .A(n44159), .B(n44160), .Z(n44152) );
  NOR U44094 ( .A(n44161), .B(n44162), .Z(n44160) );
  XNOR U44095 ( .A(n44159), .B(n44163), .Z(n44161) );
  XOR U44096 ( .A(n44164), .B(n44165), .Z(n44107) );
  NOR U44097 ( .A(n44166), .B(n44167), .Z(n44165) );
  XNOR U44098 ( .A(n44164), .B(n44168), .Z(n44166) );
  XNOR U44099 ( .A(n44117), .B(n44108), .Z(n44151) );
  XOR U44100 ( .A(n44169), .B(n44170), .Z(n44108) );
  AND U44101 ( .A(n44171), .B(n44172), .Z(n44170) );
  XOR U44102 ( .A(n44169), .B(n44173), .Z(n44171) );
  XOR U44103 ( .A(n44174), .B(n44123), .Z(n44117) );
  XOR U44104 ( .A(n44175), .B(n44176), .Z(n44123) );
  NOR U44105 ( .A(n44177), .B(n44178), .Z(n44176) );
  XOR U44106 ( .A(n44175), .B(n44179), .Z(n44177) );
  XNOR U44107 ( .A(n44122), .B(n44114), .Z(n44174) );
  XOR U44108 ( .A(n44180), .B(n44181), .Z(n44114) );
  AND U44109 ( .A(n44182), .B(n44183), .Z(n44181) );
  XOR U44110 ( .A(n44180), .B(n44184), .Z(n44182) );
  XNOR U44111 ( .A(n44185), .B(n44119), .Z(n44122) );
  XOR U44112 ( .A(n44186), .B(n44187), .Z(n44119) );
  AND U44113 ( .A(n44188), .B(n44189), .Z(n44187) );
  XNOR U44114 ( .A(n44190), .B(n44191), .Z(n44188) );
  IV U44115 ( .A(n44186), .Z(n44190) );
  XNOR U44116 ( .A(n44192), .B(n44193), .Z(n44185) );
  NOR U44117 ( .A(n44194), .B(n44195), .Z(n44193) );
  XNOR U44118 ( .A(n44192), .B(n44196), .Z(n44194) );
  XOR U44119 ( .A(n44112), .B(n44124), .Z(n44150) );
  NOR U44120 ( .A(n44041), .B(n44197), .Z(n44124) );
  XNOR U44121 ( .A(n44130), .B(n44129), .Z(n44112) );
  XNOR U44122 ( .A(n44198), .B(n44135), .Z(n44129) );
  XNOR U44123 ( .A(n44199), .B(n44200), .Z(n44135) );
  NOR U44124 ( .A(n44201), .B(n44202), .Z(n44200) );
  XOR U44125 ( .A(n44199), .B(n44203), .Z(n44201) );
  XNOR U44126 ( .A(n44134), .B(n44126), .Z(n44198) );
  XOR U44127 ( .A(n44204), .B(n44205), .Z(n44126) );
  AND U44128 ( .A(n44206), .B(n44207), .Z(n44205) );
  XOR U44129 ( .A(n44204), .B(n44208), .Z(n44206) );
  XNOR U44130 ( .A(n44209), .B(n44131), .Z(n44134) );
  XOR U44131 ( .A(n44210), .B(n44211), .Z(n44131) );
  AND U44132 ( .A(n44212), .B(n44213), .Z(n44211) );
  XNOR U44133 ( .A(n44214), .B(n44215), .Z(n44212) );
  IV U44134 ( .A(n44210), .Z(n44214) );
  XNOR U44135 ( .A(n44216), .B(n44217), .Z(n44209) );
  NOR U44136 ( .A(n44218), .B(n44219), .Z(n44217) );
  XNOR U44137 ( .A(n44216), .B(n44220), .Z(n44218) );
  XOR U44138 ( .A(n44140), .B(n44139), .Z(n44130) );
  XNOR U44139 ( .A(n44221), .B(n44136), .Z(n44139) );
  XOR U44140 ( .A(n44222), .B(n44223), .Z(n44136) );
  AND U44141 ( .A(n44224), .B(n44225), .Z(n44223) );
  XNOR U44142 ( .A(n44226), .B(n44227), .Z(n44224) );
  IV U44143 ( .A(n44222), .Z(n44226) );
  XNOR U44144 ( .A(n44228), .B(n44229), .Z(n44221) );
  NOR U44145 ( .A(n44230), .B(n44231), .Z(n44229) );
  XNOR U44146 ( .A(n44228), .B(n44232), .Z(n44230) );
  XOR U44147 ( .A(n44233), .B(n44234), .Z(n44140) );
  NOR U44148 ( .A(n44235), .B(n44236), .Z(n44234) );
  XNOR U44149 ( .A(n44233), .B(n44237), .Z(n44235) );
  XNOR U44150 ( .A(n44032), .B(n44146), .Z(n44148) );
  XNOR U44151 ( .A(n44238), .B(n44239), .Z(n44032) );
  AND U44152 ( .A(n971), .B(n44240), .Z(n44239) );
  XNOR U44153 ( .A(n44241), .B(n44242), .Z(n44240) );
  AND U44154 ( .A(n44038), .B(n44041), .Z(n44146) );
  XOR U44155 ( .A(n44243), .B(n44197), .Z(n44041) );
  XNOR U44156 ( .A(p_input[1408]), .B(p_input[2048]), .Z(n44197) );
  XNOR U44157 ( .A(n44173), .B(n44172), .Z(n44243) );
  XNOR U44158 ( .A(n44244), .B(n44184), .Z(n44172) );
  XOR U44159 ( .A(n44158), .B(n44156), .Z(n44184) );
  XNOR U44160 ( .A(n44245), .B(n44163), .Z(n44156) );
  XOR U44161 ( .A(p_input[1432]), .B(p_input[2072]), .Z(n44163) );
  XOR U44162 ( .A(n44153), .B(n44162), .Z(n44245) );
  XOR U44163 ( .A(n44246), .B(n44159), .Z(n44162) );
  XOR U44164 ( .A(p_input[1430]), .B(p_input[2070]), .Z(n44159) );
  XOR U44165 ( .A(p_input[1431]), .B(n29410), .Z(n44246) );
  XOR U44166 ( .A(p_input[1426]), .B(p_input[2066]), .Z(n44153) );
  XNOR U44167 ( .A(n44168), .B(n44167), .Z(n44158) );
  XOR U44168 ( .A(n44247), .B(n44164), .Z(n44167) );
  XOR U44169 ( .A(p_input[1427]), .B(p_input[2067]), .Z(n44164) );
  XOR U44170 ( .A(p_input[1428]), .B(n29412), .Z(n44247) );
  XOR U44171 ( .A(p_input[1429]), .B(p_input[2069]), .Z(n44168) );
  XOR U44172 ( .A(n44183), .B(n44248), .Z(n44244) );
  IV U44173 ( .A(n44169), .Z(n44248) );
  XOR U44174 ( .A(p_input[1409]), .B(p_input[2049]), .Z(n44169) );
  XNOR U44175 ( .A(n44249), .B(n44191), .Z(n44183) );
  XNOR U44176 ( .A(n44179), .B(n44178), .Z(n44191) );
  XNOR U44177 ( .A(n44250), .B(n44175), .Z(n44178) );
  XNOR U44178 ( .A(p_input[1434]), .B(p_input[2074]), .Z(n44175) );
  XOR U44179 ( .A(p_input[1435]), .B(n29415), .Z(n44250) );
  XOR U44180 ( .A(p_input[1436]), .B(p_input[2076]), .Z(n44179) );
  XOR U44181 ( .A(n44189), .B(n44251), .Z(n44249) );
  IV U44182 ( .A(n44180), .Z(n44251) );
  XOR U44183 ( .A(p_input[1425]), .B(p_input[2065]), .Z(n44180) );
  XNOR U44184 ( .A(n44252), .B(n44196), .Z(n44189) );
  XNOR U44185 ( .A(p_input[1439]), .B(n29418), .Z(n44196) );
  XOR U44186 ( .A(n44186), .B(n44195), .Z(n44252) );
  XOR U44187 ( .A(n44253), .B(n44192), .Z(n44195) );
  XOR U44188 ( .A(p_input[1437]), .B(p_input[2077]), .Z(n44192) );
  XOR U44189 ( .A(p_input[1438]), .B(n29420), .Z(n44253) );
  XOR U44190 ( .A(p_input[1433]), .B(p_input[2073]), .Z(n44186) );
  XOR U44191 ( .A(n44208), .B(n44207), .Z(n44173) );
  XNOR U44192 ( .A(n44254), .B(n44215), .Z(n44207) );
  XNOR U44193 ( .A(n44203), .B(n44202), .Z(n44215) );
  XNOR U44194 ( .A(n44255), .B(n44199), .Z(n44202) );
  XNOR U44195 ( .A(p_input[1419]), .B(p_input[2059]), .Z(n44199) );
  XOR U44196 ( .A(p_input[1420]), .B(n28329), .Z(n44255) );
  XOR U44197 ( .A(p_input[1421]), .B(p_input[2061]), .Z(n44203) );
  XOR U44198 ( .A(n44213), .B(n44256), .Z(n44254) );
  IV U44199 ( .A(n44204), .Z(n44256) );
  XOR U44200 ( .A(p_input[1410]), .B(p_input[2050]), .Z(n44204) );
  XNOR U44201 ( .A(n44257), .B(n44220), .Z(n44213) );
  XNOR U44202 ( .A(p_input[1424]), .B(n28332), .Z(n44220) );
  XOR U44203 ( .A(n44210), .B(n44219), .Z(n44257) );
  XOR U44204 ( .A(n44258), .B(n44216), .Z(n44219) );
  XOR U44205 ( .A(p_input[1422]), .B(p_input[2062]), .Z(n44216) );
  XOR U44206 ( .A(p_input[1423]), .B(n28334), .Z(n44258) );
  XOR U44207 ( .A(p_input[1418]), .B(p_input[2058]), .Z(n44210) );
  XOR U44208 ( .A(n44227), .B(n44225), .Z(n44208) );
  XNOR U44209 ( .A(n44259), .B(n44232), .Z(n44225) );
  XOR U44210 ( .A(p_input[1417]), .B(p_input[2057]), .Z(n44232) );
  XOR U44211 ( .A(n44222), .B(n44231), .Z(n44259) );
  XOR U44212 ( .A(n44260), .B(n44228), .Z(n44231) );
  XOR U44213 ( .A(p_input[1415]), .B(p_input[2055]), .Z(n44228) );
  XOR U44214 ( .A(p_input[1416]), .B(n29427), .Z(n44260) );
  XOR U44215 ( .A(p_input[1411]), .B(p_input[2051]), .Z(n44222) );
  XNOR U44216 ( .A(n44237), .B(n44236), .Z(n44227) );
  XOR U44217 ( .A(n44261), .B(n44233), .Z(n44236) );
  XOR U44218 ( .A(p_input[1412]), .B(p_input[2052]), .Z(n44233) );
  XOR U44219 ( .A(p_input[1413]), .B(n29429), .Z(n44261) );
  XOR U44220 ( .A(p_input[1414]), .B(p_input[2054]), .Z(n44237) );
  XNOR U44221 ( .A(n44262), .B(n44263), .Z(n44038) );
  AND U44222 ( .A(n971), .B(n44264), .Z(n44263) );
  XNOR U44223 ( .A(n44265), .B(n44266), .Z(n971) );
  AND U44224 ( .A(n44267), .B(n44268), .Z(n44266) );
  XOR U44225 ( .A(n44052), .B(n44265), .Z(n44268) );
  XNOR U44226 ( .A(n44269), .B(n44265), .Z(n44267) );
  XOR U44227 ( .A(n44270), .B(n44271), .Z(n44265) );
  AND U44228 ( .A(n44272), .B(n44273), .Z(n44271) );
  XOR U44229 ( .A(n44067), .B(n44270), .Z(n44273) );
  XOR U44230 ( .A(n44270), .B(n44068), .Z(n44272) );
  XOR U44231 ( .A(n44274), .B(n44275), .Z(n44270) );
  AND U44232 ( .A(n44276), .B(n44277), .Z(n44275) );
  XOR U44233 ( .A(n44095), .B(n44274), .Z(n44277) );
  XOR U44234 ( .A(n44274), .B(n44096), .Z(n44276) );
  XOR U44235 ( .A(n44278), .B(n44279), .Z(n44274) );
  AND U44236 ( .A(n44280), .B(n44281), .Z(n44279) );
  XOR U44237 ( .A(n44144), .B(n44278), .Z(n44281) );
  XOR U44238 ( .A(n44278), .B(n44145), .Z(n44280) );
  XOR U44239 ( .A(n44282), .B(n44283), .Z(n44278) );
  AND U44240 ( .A(n44284), .B(n44285), .Z(n44283) );
  XOR U44241 ( .A(n44282), .B(n44241), .Z(n44285) );
  XNOR U44242 ( .A(n44286), .B(n44287), .Z(n43988) );
  AND U44243 ( .A(n975), .B(n44288), .Z(n44287) );
  XNOR U44244 ( .A(n44289), .B(n44290), .Z(n975) );
  AND U44245 ( .A(n44291), .B(n44292), .Z(n44290) );
  XOR U44246 ( .A(n44289), .B(n43998), .Z(n44292) );
  XNOR U44247 ( .A(n44289), .B(n43948), .Z(n44291) );
  XOR U44248 ( .A(n44293), .B(n44294), .Z(n44289) );
  AND U44249 ( .A(n44295), .B(n44296), .Z(n44294) );
  XNOR U44250 ( .A(n44008), .B(n44293), .Z(n44296) );
  XOR U44251 ( .A(n44293), .B(n43958), .Z(n44295) );
  XOR U44252 ( .A(n44297), .B(n44298), .Z(n44293) );
  AND U44253 ( .A(n44299), .B(n44300), .Z(n44298) );
  XNOR U44254 ( .A(n44018), .B(n44297), .Z(n44300) );
  XOR U44255 ( .A(n44297), .B(n43967), .Z(n44299) );
  XOR U44256 ( .A(n44301), .B(n44302), .Z(n44297) );
  AND U44257 ( .A(n44303), .B(n44304), .Z(n44302) );
  XOR U44258 ( .A(n44301), .B(n43975), .Z(n44303) );
  XOR U44259 ( .A(n44305), .B(n44306), .Z(n43939) );
  AND U44260 ( .A(n979), .B(n44288), .Z(n44306) );
  XNOR U44261 ( .A(n44286), .B(n44305), .Z(n44288) );
  XNOR U44262 ( .A(n44307), .B(n44308), .Z(n979) );
  AND U44263 ( .A(n44309), .B(n44310), .Z(n44308) );
  XNOR U44264 ( .A(n44311), .B(n44307), .Z(n44310) );
  IV U44265 ( .A(n43998), .Z(n44311) );
  XOR U44266 ( .A(n44269), .B(n44312), .Z(n43998) );
  AND U44267 ( .A(n982), .B(n44313), .Z(n44312) );
  XOR U44268 ( .A(n44051), .B(n44048), .Z(n44313) );
  IV U44269 ( .A(n44269), .Z(n44051) );
  XNOR U44270 ( .A(n43948), .B(n44307), .Z(n44309) );
  XOR U44271 ( .A(n44314), .B(n44315), .Z(n43948) );
  AND U44272 ( .A(n998), .B(n44316), .Z(n44315) );
  XOR U44273 ( .A(n44317), .B(n44318), .Z(n44307) );
  AND U44274 ( .A(n44319), .B(n44320), .Z(n44318) );
  XNOR U44275 ( .A(n44317), .B(n44008), .Z(n44320) );
  XOR U44276 ( .A(n44068), .B(n44321), .Z(n44008) );
  AND U44277 ( .A(n982), .B(n44322), .Z(n44321) );
  XOR U44278 ( .A(n44064), .B(n44068), .Z(n44322) );
  XNOR U44279 ( .A(n44323), .B(n44317), .Z(n44319) );
  IV U44280 ( .A(n43958), .Z(n44323) );
  XOR U44281 ( .A(n44324), .B(n44325), .Z(n43958) );
  AND U44282 ( .A(n998), .B(n44326), .Z(n44325) );
  XOR U44283 ( .A(n44327), .B(n44328), .Z(n44317) );
  AND U44284 ( .A(n44329), .B(n44330), .Z(n44328) );
  XNOR U44285 ( .A(n44327), .B(n44018), .Z(n44330) );
  XOR U44286 ( .A(n44096), .B(n44331), .Z(n44018) );
  AND U44287 ( .A(n982), .B(n44332), .Z(n44331) );
  XOR U44288 ( .A(n44092), .B(n44096), .Z(n44332) );
  XOR U44289 ( .A(n43967), .B(n44327), .Z(n44329) );
  XOR U44290 ( .A(n44333), .B(n44334), .Z(n43967) );
  AND U44291 ( .A(n998), .B(n44335), .Z(n44334) );
  XOR U44292 ( .A(n44301), .B(n44336), .Z(n44327) );
  AND U44293 ( .A(n44337), .B(n44304), .Z(n44336) );
  XNOR U44294 ( .A(n44028), .B(n44301), .Z(n44304) );
  XOR U44295 ( .A(n44145), .B(n44338), .Z(n44028) );
  AND U44296 ( .A(n982), .B(n44339), .Z(n44338) );
  XOR U44297 ( .A(n44141), .B(n44145), .Z(n44339) );
  XNOR U44298 ( .A(n44340), .B(n44301), .Z(n44337) );
  IV U44299 ( .A(n43975), .Z(n44340) );
  XOR U44300 ( .A(n44341), .B(n44342), .Z(n43975) );
  AND U44301 ( .A(n998), .B(n44343), .Z(n44342) );
  XOR U44302 ( .A(n44344), .B(n44345), .Z(n44301) );
  AND U44303 ( .A(n44346), .B(n44347), .Z(n44345) );
  XNOR U44304 ( .A(n44344), .B(n44036), .Z(n44347) );
  XOR U44305 ( .A(n44242), .B(n44348), .Z(n44036) );
  AND U44306 ( .A(n982), .B(n44349), .Z(n44348) );
  XOR U44307 ( .A(n44238), .B(n44242), .Z(n44349) );
  XNOR U44308 ( .A(n44350), .B(n44344), .Z(n44346) );
  IV U44309 ( .A(n43985), .Z(n44350) );
  XOR U44310 ( .A(n44351), .B(n44352), .Z(n43985) );
  AND U44311 ( .A(n998), .B(n44353), .Z(n44352) );
  AND U44312 ( .A(n44305), .B(n44286), .Z(n44344) );
  XNOR U44313 ( .A(n44354), .B(n44355), .Z(n44286) );
  AND U44314 ( .A(n982), .B(n44264), .Z(n44355) );
  XNOR U44315 ( .A(n44262), .B(n44354), .Z(n44264) );
  XNOR U44316 ( .A(n44356), .B(n44357), .Z(n982) );
  AND U44317 ( .A(n44358), .B(n44359), .Z(n44357) );
  XNOR U44318 ( .A(n44356), .B(n44048), .Z(n44359) );
  IV U44319 ( .A(n44052), .Z(n44048) );
  XOR U44320 ( .A(n44360), .B(n44361), .Z(n44052) );
  AND U44321 ( .A(n986), .B(n44362), .Z(n44361) );
  XOR U44322 ( .A(n44363), .B(n44360), .Z(n44362) );
  XNOR U44323 ( .A(n44356), .B(n44269), .Z(n44358) );
  XOR U44324 ( .A(n44364), .B(n44365), .Z(n44269) );
  AND U44325 ( .A(n994), .B(n44316), .Z(n44365) );
  XOR U44326 ( .A(n44314), .B(n44364), .Z(n44316) );
  XOR U44327 ( .A(n44366), .B(n44367), .Z(n44356) );
  AND U44328 ( .A(n44368), .B(n44369), .Z(n44367) );
  XNOR U44329 ( .A(n44366), .B(n44064), .Z(n44369) );
  IV U44330 ( .A(n44067), .Z(n44064) );
  XOR U44331 ( .A(n44370), .B(n44371), .Z(n44067) );
  AND U44332 ( .A(n986), .B(n44372), .Z(n44371) );
  XOR U44333 ( .A(n44373), .B(n44370), .Z(n44372) );
  XOR U44334 ( .A(n44068), .B(n44366), .Z(n44368) );
  XOR U44335 ( .A(n44374), .B(n44375), .Z(n44068) );
  AND U44336 ( .A(n994), .B(n44326), .Z(n44375) );
  XOR U44337 ( .A(n44374), .B(n44324), .Z(n44326) );
  XOR U44338 ( .A(n44376), .B(n44377), .Z(n44366) );
  AND U44339 ( .A(n44378), .B(n44379), .Z(n44377) );
  XNOR U44340 ( .A(n44376), .B(n44092), .Z(n44379) );
  IV U44341 ( .A(n44095), .Z(n44092) );
  XOR U44342 ( .A(n44380), .B(n44381), .Z(n44095) );
  AND U44343 ( .A(n986), .B(n44382), .Z(n44381) );
  XNOR U44344 ( .A(n44383), .B(n44380), .Z(n44382) );
  XOR U44345 ( .A(n44096), .B(n44376), .Z(n44378) );
  XOR U44346 ( .A(n44384), .B(n44385), .Z(n44096) );
  AND U44347 ( .A(n994), .B(n44335), .Z(n44385) );
  XOR U44348 ( .A(n44384), .B(n44333), .Z(n44335) );
  XOR U44349 ( .A(n44386), .B(n44387), .Z(n44376) );
  AND U44350 ( .A(n44388), .B(n44389), .Z(n44387) );
  XNOR U44351 ( .A(n44386), .B(n44141), .Z(n44389) );
  IV U44352 ( .A(n44144), .Z(n44141) );
  XOR U44353 ( .A(n44390), .B(n44391), .Z(n44144) );
  AND U44354 ( .A(n986), .B(n44392), .Z(n44391) );
  XOR U44355 ( .A(n44393), .B(n44390), .Z(n44392) );
  XOR U44356 ( .A(n44145), .B(n44386), .Z(n44388) );
  XOR U44357 ( .A(n44394), .B(n44395), .Z(n44145) );
  AND U44358 ( .A(n994), .B(n44343), .Z(n44395) );
  XOR U44359 ( .A(n44394), .B(n44341), .Z(n44343) );
  XOR U44360 ( .A(n44282), .B(n44396), .Z(n44386) );
  AND U44361 ( .A(n44284), .B(n44397), .Z(n44396) );
  XNOR U44362 ( .A(n44282), .B(n44238), .Z(n44397) );
  IV U44363 ( .A(n44241), .Z(n44238) );
  XOR U44364 ( .A(n44398), .B(n44399), .Z(n44241) );
  AND U44365 ( .A(n986), .B(n44400), .Z(n44399) );
  XNOR U44366 ( .A(n44401), .B(n44398), .Z(n44400) );
  XOR U44367 ( .A(n44242), .B(n44282), .Z(n44284) );
  XOR U44368 ( .A(n44402), .B(n44403), .Z(n44242) );
  AND U44369 ( .A(n994), .B(n44353), .Z(n44403) );
  XOR U44370 ( .A(n44402), .B(n44351), .Z(n44353) );
  AND U44371 ( .A(n44354), .B(n44262), .Z(n44282) );
  XNOR U44372 ( .A(n44404), .B(n44405), .Z(n44262) );
  AND U44373 ( .A(n986), .B(n44406), .Z(n44405) );
  XNOR U44374 ( .A(n44407), .B(n44404), .Z(n44406) );
  XNOR U44375 ( .A(n44408), .B(n44409), .Z(n986) );
  AND U44376 ( .A(n44410), .B(n44411), .Z(n44409) );
  XOR U44377 ( .A(n44363), .B(n44408), .Z(n44411) );
  AND U44378 ( .A(n44412), .B(n44413), .Z(n44363) );
  XNOR U44379 ( .A(n44360), .B(n44408), .Z(n44410) );
  XNOR U44380 ( .A(n44414), .B(n44415), .Z(n44360) );
  AND U44381 ( .A(n990), .B(n44416), .Z(n44415) );
  XNOR U44382 ( .A(n44417), .B(n44418), .Z(n44416) );
  XOR U44383 ( .A(n44419), .B(n44420), .Z(n44408) );
  AND U44384 ( .A(n44421), .B(n44422), .Z(n44420) );
  XNOR U44385 ( .A(n44419), .B(n44412), .Z(n44422) );
  IV U44386 ( .A(n44373), .Z(n44412) );
  XOR U44387 ( .A(n44423), .B(n44424), .Z(n44373) );
  XOR U44388 ( .A(n44425), .B(n44413), .Z(n44424) );
  AND U44389 ( .A(n44383), .B(n44426), .Z(n44413) );
  AND U44390 ( .A(n44427), .B(n44428), .Z(n44425) );
  XOR U44391 ( .A(n44429), .B(n44423), .Z(n44427) );
  XNOR U44392 ( .A(n44370), .B(n44419), .Z(n44421) );
  XNOR U44393 ( .A(n44430), .B(n44431), .Z(n44370) );
  AND U44394 ( .A(n990), .B(n44432), .Z(n44431) );
  XNOR U44395 ( .A(n44433), .B(n44434), .Z(n44432) );
  XOR U44396 ( .A(n44435), .B(n44436), .Z(n44419) );
  AND U44397 ( .A(n44437), .B(n44438), .Z(n44436) );
  XNOR U44398 ( .A(n44435), .B(n44383), .Z(n44438) );
  XOR U44399 ( .A(n44439), .B(n44428), .Z(n44383) );
  XNOR U44400 ( .A(n44440), .B(n44423), .Z(n44428) );
  XOR U44401 ( .A(n44441), .B(n44442), .Z(n44423) );
  AND U44402 ( .A(n44443), .B(n44444), .Z(n44442) );
  XOR U44403 ( .A(n44445), .B(n44441), .Z(n44443) );
  XNOR U44404 ( .A(n44446), .B(n44447), .Z(n44440) );
  AND U44405 ( .A(n44448), .B(n44449), .Z(n44447) );
  XOR U44406 ( .A(n44446), .B(n44450), .Z(n44448) );
  XNOR U44407 ( .A(n44429), .B(n44426), .Z(n44439) );
  AND U44408 ( .A(n44451), .B(n44452), .Z(n44426) );
  XOR U44409 ( .A(n44453), .B(n44454), .Z(n44429) );
  AND U44410 ( .A(n44455), .B(n44456), .Z(n44454) );
  XOR U44411 ( .A(n44453), .B(n44457), .Z(n44455) );
  XNOR U44412 ( .A(n44380), .B(n44435), .Z(n44437) );
  XNOR U44413 ( .A(n44458), .B(n44459), .Z(n44380) );
  AND U44414 ( .A(n990), .B(n44460), .Z(n44459) );
  XNOR U44415 ( .A(n44461), .B(n44462), .Z(n44460) );
  XOR U44416 ( .A(n44463), .B(n44464), .Z(n44435) );
  AND U44417 ( .A(n44465), .B(n44466), .Z(n44464) );
  XNOR U44418 ( .A(n44463), .B(n44451), .Z(n44466) );
  IV U44419 ( .A(n44393), .Z(n44451) );
  XNOR U44420 ( .A(n44467), .B(n44444), .Z(n44393) );
  XNOR U44421 ( .A(n44468), .B(n44450), .Z(n44444) );
  XOR U44422 ( .A(n44469), .B(n44470), .Z(n44450) );
  AND U44423 ( .A(n44471), .B(n44472), .Z(n44470) );
  XOR U44424 ( .A(n44469), .B(n44473), .Z(n44471) );
  XNOR U44425 ( .A(n44449), .B(n44441), .Z(n44468) );
  XOR U44426 ( .A(n44474), .B(n44475), .Z(n44441) );
  AND U44427 ( .A(n44476), .B(n44477), .Z(n44475) );
  XNOR U44428 ( .A(n44478), .B(n44474), .Z(n44476) );
  XNOR U44429 ( .A(n44479), .B(n44446), .Z(n44449) );
  XOR U44430 ( .A(n44480), .B(n44481), .Z(n44446) );
  AND U44431 ( .A(n44482), .B(n44483), .Z(n44481) );
  XOR U44432 ( .A(n44480), .B(n44484), .Z(n44482) );
  XNOR U44433 ( .A(n44485), .B(n44486), .Z(n44479) );
  AND U44434 ( .A(n44487), .B(n44488), .Z(n44486) );
  XNOR U44435 ( .A(n44485), .B(n44489), .Z(n44487) );
  XNOR U44436 ( .A(n44445), .B(n44452), .Z(n44467) );
  AND U44437 ( .A(n44401), .B(n44490), .Z(n44452) );
  XOR U44438 ( .A(n44457), .B(n44456), .Z(n44445) );
  XNOR U44439 ( .A(n44491), .B(n44453), .Z(n44456) );
  XOR U44440 ( .A(n44492), .B(n44493), .Z(n44453) );
  AND U44441 ( .A(n44494), .B(n44495), .Z(n44493) );
  XOR U44442 ( .A(n44492), .B(n44496), .Z(n44494) );
  XNOR U44443 ( .A(n44497), .B(n44498), .Z(n44491) );
  AND U44444 ( .A(n44499), .B(n44500), .Z(n44498) );
  XOR U44445 ( .A(n44497), .B(n44501), .Z(n44499) );
  XOR U44446 ( .A(n44502), .B(n44503), .Z(n44457) );
  AND U44447 ( .A(n44504), .B(n44505), .Z(n44503) );
  XOR U44448 ( .A(n44502), .B(n44506), .Z(n44504) );
  XNOR U44449 ( .A(n44390), .B(n44463), .Z(n44465) );
  XNOR U44450 ( .A(n44507), .B(n44508), .Z(n44390) );
  AND U44451 ( .A(n990), .B(n44509), .Z(n44508) );
  XNOR U44452 ( .A(n44510), .B(n44511), .Z(n44509) );
  XOR U44453 ( .A(n44512), .B(n44513), .Z(n44463) );
  AND U44454 ( .A(n44514), .B(n44515), .Z(n44513) );
  XNOR U44455 ( .A(n44512), .B(n44401), .Z(n44515) );
  XOR U44456 ( .A(n44516), .B(n44477), .Z(n44401) );
  XNOR U44457 ( .A(n44517), .B(n44484), .Z(n44477) );
  XOR U44458 ( .A(n44473), .B(n44472), .Z(n44484) );
  XNOR U44459 ( .A(n44518), .B(n44469), .Z(n44472) );
  XOR U44460 ( .A(n44519), .B(n44520), .Z(n44469) );
  AND U44461 ( .A(n44521), .B(n44522), .Z(n44520) );
  XNOR U44462 ( .A(n44523), .B(n44524), .Z(n44521) );
  IV U44463 ( .A(n44519), .Z(n44523) );
  XNOR U44464 ( .A(n44525), .B(n44526), .Z(n44518) );
  NOR U44465 ( .A(n44527), .B(n44528), .Z(n44526) );
  XNOR U44466 ( .A(n44525), .B(n44529), .Z(n44527) );
  XOR U44467 ( .A(n44530), .B(n44531), .Z(n44473) );
  NOR U44468 ( .A(n44532), .B(n44533), .Z(n44531) );
  XNOR U44469 ( .A(n44530), .B(n44534), .Z(n44532) );
  XNOR U44470 ( .A(n44483), .B(n44474), .Z(n44517) );
  XOR U44471 ( .A(n44535), .B(n44536), .Z(n44474) );
  AND U44472 ( .A(n44537), .B(n44538), .Z(n44536) );
  XOR U44473 ( .A(n44535), .B(n44539), .Z(n44537) );
  XOR U44474 ( .A(n44540), .B(n44489), .Z(n44483) );
  XOR U44475 ( .A(n44541), .B(n44542), .Z(n44489) );
  NOR U44476 ( .A(n44543), .B(n44544), .Z(n44542) );
  XOR U44477 ( .A(n44541), .B(n44545), .Z(n44543) );
  XNOR U44478 ( .A(n44488), .B(n44480), .Z(n44540) );
  XOR U44479 ( .A(n44546), .B(n44547), .Z(n44480) );
  AND U44480 ( .A(n44548), .B(n44549), .Z(n44547) );
  XOR U44481 ( .A(n44546), .B(n44550), .Z(n44548) );
  XNOR U44482 ( .A(n44551), .B(n44485), .Z(n44488) );
  XOR U44483 ( .A(n44552), .B(n44553), .Z(n44485) );
  AND U44484 ( .A(n44554), .B(n44555), .Z(n44553) );
  XNOR U44485 ( .A(n44556), .B(n44557), .Z(n44554) );
  IV U44486 ( .A(n44552), .Z(n44556) );
  XNOR U44487 ( .A(n44558), .B(n44559), .Z(n44551) );
  NOR U44488 ( .A(n44560), .B(n44561), .Z(n44559) );
  XNOR U44489 ( .A(n44558), .B(n44562), .Z(n44560) );
  XOR U44490 ( .A(n44478), .B(n44490), .Z(n44516) );
  NOR U44491 ( .A(n44407), .B(n44563), .Z(n44490) );
  XNOR U44492 ( .A(n44496), .B(n44495), .Z(n44478) );
  XNOR U44493 ( .A(n44564), .B(n44501), .Z(n44495) );
  XNOR U44494 ( .A(n44565), .B(n44566), .Z(n44501) );
  NOR U44495 ( .A(n44567), .B(n44568), .Z(n44566) );
  XOR U44496 ( .A(n44565), .B(n44569), .Z(n44567) );
  XNOR U44497 ( .A(n44500), .B(n44492), .Z(n44564) );
  XOR U44498 ( .A(n44570), .B(n44571), .Z(n44492) );
  AND U44499 ( .A(n44572), .B(n44573), .Z(n44571) );
  XOR U44500 ( .A(n44570), .B(n44574), .Z(n44572) );
  XNOR U44501 ( .A(n44575), .B(n44497), .Z(n44500) );
  XOR U44502 ( .A(n44576), .B(n44577), .Z(n44497) );
  AND U44503 ( .A(n44578), .B(n44579), .Z(n44577) );
  XNOR U44504 ( .A(n44580), .B(n44581), .Z(n44578) );
  IV U44505 ( .A(n44576), .Z(n44580) );
  XNOR U44506 ( .A(n44582), .B(n44583), .Z(n44575) );
  NOR U44507 ( .A(n44584), .B(n44585), .Z(n44583) );
  XNOR U44508 ( .A(n44582), .B(n44586), .Z(n44584) );
  XOR U44509 ( .A(n44506), .B(n44505), .Z(n44496) );
  XNOR U44510 ( .A(n44587), .B(n44502), .Z(n44505) );
  XOR U44511 ( .A(n44588), .B(n44589), .Z(n44502) );
  AND U44512 ( .A(n44590), .B(n44591), .Z(n44589) );
  XNOR U44513 ( .A(n44592), .B(n44593), .Z(n44590) );
  IV U44514 ( .A(n44588), .Z(n44592) );
  XNOR U44515 ( .A(n44594), .B(n44595), .Z(n44587) );
  NOR U44516 ( .A(n44596), .B(n44597), .Z(n44595) );
  XNOR U44517 ( .A(n44594), .B(n44598), .Z(n44596) );
  XOR U44518 ( .A(n44599), .B(n44600), .Z(n44506) );
  NOR U44519 ( .A(n44601), .B(n44602), .Z(n44600) );
  XNOR U44520 ( .A(n44599), .B(n44603), .Z(n44601) );
  XNOR U44521 ( .A(n44398), .B(n44512), .Z(n44514) );
  XNOR U44522 ( .A(n44604), .B(n44605), .Z(n44398) );
  AND U44523 ( .A(n990), .B(n44606), .Z(n44605) );
  XNOR U44524 ( .A(n44607), .B(n44608), .Z(n44606) );
  AND U44525 ( .A(n44404), .B(n44407), .Z(n44512) );
  XOR U44526 ( .A(n44609), .B(n44563), .Z(n44407) );
  XNOR U44527 ( .A(p_input[1440]), .B(p_input[2048]), .Z(n44563) );
  XNOR U44528 ( .A(n44539), .B(n44538), .Z(n44609) );
  XNOR U44529 ( .A(n44610), .B(n44550), .Z(n44538) );
  XOR U44530 ( .A(n44524), .B(n44522), .Z(n44550) );
  XNOR U44531 ( .A(n44611), .B(n44529), .Z(n44522) );
  XOR U44532 ( .A(p_input[1464]), .B(p_input[2072]), .Z(n44529) );
  XOR U44533 ( .A(n44519), .B(n44528), .Z(n44611) );
  XOR U44534 ( .A(n44612), .B(n44525), .Z(n44528) );
  XOR U44535 ( .A(p_input[1462]), .B(p_input[2070]), .Z(n44525) );
  XOR U44536 ( .A(p_input[1463]), .B(n29410), .Z(n44612) );
  XOR U44537 ( .A(p_input[1458]), .B(p_input[2066]), .Z(n44519) );
  XNOR U44538 ( .A(n44534), .B(n44533), .Z(n44524) );
  XOR U44539 ( .A(n44613), .B(n44530), .Z(n44533) );
  XOR U44540 ( .A(p_input[1459]), .B(p_input[2067]), .Z(n44530) );
  XOR U44541 ( .A(p_input[1460]), .B(n29412), .Z(n44613) );
  XOR U44542 ( .A(p_input[1461]), .B(p_input[2069]), .Z(n44534) );
  XOR U44543 ( .A(n44549), .B(n44614), .Z(n44610) );
  IV U44544 ( .A(n44535), .Z(n44614) );
  XOR U44545 ( .A(p_input[1441]), .B(p_input[2049]), .Z(n44535) );
  XNOR U44546 ( .A(n44615), .B(n44557), .Z(n44549) );
  XNOR U44547 ( .A(n44545), .B(n44544), .Z(n44557) );
  XNOR U44548 ( .A(n44616), .B(n44541), .Z(n44544) );
  XNOR U44549 ( .A(p_input[1466]), .B(p_input[2074]), .Z(n44541) );
  XOR U44550 ( .A(p_input[1467]), .B(n29415), .Z(n44616) );
  XOR U44551 ( .A(p_input[1468]), .B(p_input[2076]), .Z(n44545) );
  XOR U44552 ( .A(n44555), .B(n44617), .Z(n44615) );
  IV U44553 ( .A(n44546), .Z(n44617) );
  XOR U44554 ( .A(p_input[1457]), .B(p_input[2065]), .Z(n44546) );
  XNOR U44555 ( .A(n44618), .B(n44562), .Z(n44555) );
  XNOR U44556 ( .A(p_input[1471]), .B(n29418), .Z(n44562) );
  XOR U44557 ( .A(n44552), .B(n44561), .Z(n44618) );
  XOR U44558 ( .A(n44619), .B(n44558), .Z(n44561) );
  XOR U44559 ( .A(p_input[1469]), .B(p_input[2077]), .Z(n44558) );
  XOR U44560 ( .A(p_input[1470]), .B(n29420), .Z(n44619) );
  XOR U44561 ( .A(p_input[1465]), .B(p_input[2073]), .Z(n44552) );
  XOR U44562 ( .A(n44574), .B(n44573), .Z(n44539) );
  XNOR U44563 ( .A(n44620), .B(n44581), .Z(n44573) );
  XNOR U44564 ( .A(n44569), .B(n44568), .Z(n44581) );
  XNOR U44565 ( .A(n44621), .B(n44565), .Z(n44568) );
  XNOR U44566 ( .A(p_input[1451]), .B(p_input[2059]), .Z(n44565) );
  XOR U44567 ( .A(p_input[1452]), .B(n28329), .Z(n44621) );
  XOR U44568 ( .A(p_input[1453]), .B(p_input[2061]), .Z(n44569) );
  XOR U44569 ( .A(n44579), .B(n44622), .Z(n44620) );
  IV U44570 ( .A(n44570), .Z(n44622) );
  XOR U44571 ( .A(p_input[1442]), .B(p_input[2050]), .Z(n44570) );
  XNOR U44572 ( .A(n44623), .B(n44586), .Z(n44579) );
  XNOR U44573 ( .A(p_input[1456]), .B(n28332), .Z(n44586) );
  XOR U44574 ( .A(n44576), .B(n44585), .Z(n44623) );
  XOR U44575 ( .A(n44624), .B(n44582), .Z(n44585) );
  XOR U44576 ( .A(p_input[1454]), .B(p_input[2062]), .Z(n44582) );
  XOR U44577 ( .A(p_input[1455]), .B(n28334), .Z(n44624) );
  XOR U44578 ( .A(p_input[1450]), .B(p_input[2058]), .Z(n44576) );
  XOR U44579 ( .A(n44593), .B(n44591), .Z(n44574) );
  XNOR U44580 ( .A(n44625), .B(n44598), .Z(n44591) );
  XOR U44581 ( .A(p_input[1449]), .B(p_input[2057]), .Z(n44598) );
  XOR U44582 ( .A(n44588), .B(n44597), .Z(n44625) );
  XOR U44583 ( .A(n44626), .B(n44594), .Z(n44597) );
  XOR U44584 ( .A(p_input[1447]), .B(p_input[2055]), .Z(n44594) );
  XOR U44585 ( .A(p_input[1448]), .B(n29427), .Z(n44626) );
  XOR U44586 ( .A(p_input[1443]), .B(p_input[2051]), .Z(n44588) );
  XNOR U44587 ( .A(n44603), .B(n44602), .Z(n44593) );
  XOR U44588 ( .A(n44627), .B(n44599), .Z(n44602) );
  XOR U44589 ( .A(p_input[1444]), .B(p_input[2052]), .Z(n44599) );
  XOR U44590 ( .A(p_input[1445]), .B(n29429), .Z(n44627) );
  XOR U44591 ( .A(p_input[1446]), .B(p_input[2054]), .Z(n44603) );
  XNOR U44592 ( .A(n44628), .B(n44629), .Z(n44404) );
  AND U44593 ( .A(n990), .B(n44630), .Z(n44629) );
  XNOR U44594 ( .A(n44631), .B(n44632), .Z(n990) );
  AND U44595 ( .A(n44633), .B(n44634), .Z(n44632) );
  XOR U44596 ( .A(n44418), .B(n44631), .Z(n44634) );
  XNOR U44597 ( .A(n44635), .B(n44631), .Z(n44633) );
  XOR U44598 ( .A(n44636), .B(n44637), .Z(n44631) );
  AND U44599 ( .A(n44638), .B(n44639), .Z(n44637) );
  XOR U44600 ( .A(n44433), .B(n44636), .Z(n44639) );
  XOR U44601 ( .A(n44636), .B(n44434), .Z(n44638) );
  XOR U44602 ( .A(n44640), .B(n44641), .Z(n44636) );
  AND U44603 ( .A(n44642), .B(n44643), .Z(n44641) );
  XOR U44604 ( .A(n44461), .B(n44640), .Z(n44643) );
  XOR U44605 ( .A(n44640), .B(n44462), .Z(n44642) );
  XOR U44606 ( .A(n44644), .B(n44645), .Z(n44640) );
  AND U44607 ( .A(n44646), .B(n44647), .Z(n44645) );
  XOR U44608 ( .A(n44510), .B(n44644), .Z(n44647) );
  XOR U44609 ( .A(n44644), .B(n44511), .Z(n44646) );
  XOR U44610 ( .A(n44648), .B(n44649), .Z(n44644) );
  AND U44611 ( .A(n44650), .B(n44651), .Z(n44649) );
  XOR U44612 ( .A(n44648), .B(n44607), .Z(n44651) );
  XNOR U44613 ( .A(n44652), .B(n44653), .Z(n44354) );
  AND U44614 ( .A(n994), .B(n44654), .Z(n44653) );
  XNOR U44615 ( .A(n44655), .B(n44656), .Z(n994) );
  AND U44616 ( .A(n44657), .B(n44658), .Z(n44656) );
  XOR U44617 ( .A(n44655), .B(n44364), .Z(n44658) );
  XNOR U44618 ( .A(n44655), .B(n44314), .Z(n44657) );
  XOR U44619 ( .A(n44659), .B(n44660), .Z(n44655) );
  AND U44620 ( .A(n44661), .B(n44662), .Z(n44660) );
  XNOR U44621 ( .A(n44374), .B(n44659), .Z(n44662) );
  XOR U44622 ( .A(n44659), .B(n44324), .Z(n44661) );
  XOR U44623 ( .A(n44663), .B(n44664), .Z(n44659) );
  AND U44624 ( .A(n44665), .B(n44666), .Z(n44664) );
  XNOR U44625 ( .A(n44384), .B(n44663), .Z(n44666) );
  XOR U44626 ( .A(n44663), .B(n44333), .Z(n44665) );
  XOR U44627 ( .A(n44667), .B(n44668), .Z(n44663) );
  AND U44628 ( .A(n44669), .B(n44670), .Z(n44668) );
  XOR U44629 ( .A(n44667), .B(n44341), .Z(n44669) );
  XOR U44630 ( .A(n44671), .B(n44672), .Z(n44305) );
  AND U44631 ( .A(n998), .B(n44654), .Z(n44672) );
  XNOR U44632 ( .A(n44652), .B(n44671), .Z(n44654) );
  XNOR U44633 ( .A(n44673), .B(n44674), .Z(n998) );
  AND U44634 ( .A(n44675), .B(n44676), .Z(n44674) );
  XNOR U44635 ( .A(n44677), .B(n44673), .Z(n44676) );
  IV U44636 ( .A(n44364), .Z(n44677) );
  XOR U44637 ( .A(n44635), .B(n44678), .Z(n44364) );
  AND U44638 ( .A(n1001), .B(n44679), .Z(n44678) );
  XOR U44639 ( .A(n44417), .B(n44414), .Z(n44679) );
  IV U44640 ( .A(n44635), .Z(n44417) );
  XNOR U44641 ( .A(n44314), .B(n44673), .Z(n44675) );
  XOR U44642 ( .A(n44680), .B(n44681), .Z(n44314) );
  AND U44643 ( .A(n1017), .B(n44682), .Z(n44681) );
  XOR U44644 ( .A(n44683), .B(n44684), .Z(n44673) );
  AND U44645 ( .A(n44685), .B(n44686), .Z(n44684) );
  XNOR U44646 ( .A(n44683), .B(n44374), .Z(n44686) );
  XOR U44647 ( .A(n44434), .B(n44687), .Z(n44374) );
  AND U44648 ( .A(n1001), .B(n44688), .Z(n44687) );
  XOR U44649 ( .A(n44430), .B(n44434), .Z(n44688) );
  XNOR U44650 ( .A(n44689), .B(n44683), .Z(n44685) );
  IV U44651 ( .A(n44324), .Z(n44689) );
  XOR U44652 ( .A(n44690), .B(n44691), .Z(n44324) );
  AND U44653 ( .A(n1017), .B(n44692), .Z(n44691) );
  XOR U44654 ( .A(n44693), .B(n44694), .Z(n44683) );
  AND U44655 ( .A(n44695), .B(n44696), .Z(n44694) );
  XNOR U44656 ( .A(n44693), .B(n44384), .Z(n44696) );
  XOR U44657 ( .A(n44462), .B(n44697), .Z(n44384) );
  AND U44658 ( .A(n1001), .B(n44698), .Z(n44697) );
  XOR U44659 ( .A(n44458), .B(n44462), .Z(n44698) );
  XOR U44660 ( .A(n44333), .B(n44693), .Z(n44695) );
  XOR U44661 ( .A(n44699), .B(n44700), .Z(n44333) );
  AND U44662 ( .A(n1017), .B(n44701), .Z(n44700) );
  XOR U44663 ( .A(n44667), .B(n44702), .Z(n44693) );
  AND U44664 ( .A(n44703), .B(n44670), .Z(n44702) );
  XNOR U44665 ( .A(n44394), .B(n44667), .Z(n44670) );
  XOR U44666 ( .A(n44511), .B(n44704), .Z(n44394) );
  AND U44667 ( .A(n1001), .B(n44705), .Z(n44704) );
  XOR U44668 ( .A(n44507), .B(n44511), .Z(n44705) );
  XNOR U44669 ( .A(n44706), .B(n44667), .Z(n44703) );
  IV U44670 ( .A(n44341), .Z(n44706) );
  XOR U44671 ( .A(n44707), .B(n44708), .Z(n44341) );
  AND U44672 ( .A(n1017), .B(n44709), .Z(n44708) );
  XOR U44673 ( .A(n44710), .B(n44711), .Z(n44667) );
  AND U44674 ( .A(n44712), .B(n44713), .Z(n44711) );
  XNOR U44675 ( .A(n44710), .B(n44402), .Z(n44713) );
  XOR U44676 ( .A(n44608), .B(n44714), .Z(n44402) );
  AND U44677 ( .A(n1001), .B(n44715), .Z(n44714) );
  XOR U44678 ( .A(n44604), .B(n44608), .Z(n44715) );
  XNOR U44679 ( .A(n44716), .B(n44710), .Z(n44712) );
  IV U44680 ( .A(n44351), .Z(n44716) );
  XOR U44681 ( .A(n44717), .B(n44718), .Z(n44351) );
  AND U44682 ( .A(n1017), .B(n44719), .Z(n44718) );
  AND U44683 ( .A(n44671), .B(n44652), .Z(n44710) );
  XNOR U44684 ( .A(n44720), .B(n44721), .Z(n44652) );
  AND U44685 ( .A(n1001), .B(n44630), .Z(n44721) );
  XNOR U44686 ( .A(n44628), .B(n44720), .Z(n44630) );
  XNOR U44687 ( .A(n44722), .B(n44723), .Z(n1001) );
  AND U44688 ( .A(n44724), .B(n44725), .Z(n44723) );
  XNOR U44689 ( .A(n44722), .B(n44414), .Z(n44725) );
  IV U44690 ( .A(n44418), .Z(n44414) );
  XOR U44691 ( .A(n44726), .B(n44727), .Z(n44418) );
  AND U44692 ( .A(n1005), .B(n44728), .Z(n44727) );
  XOR U44693 ( .A(n44729), .B(n44726), .Z(n44728) );
  XNOR U44694 ( .A(n44722), .B(n44635), .Z(n44724) );
  XOR U44695 ( .A(n44730), .B(n44731), .Z(n44635) );
  AND U44696 ( .A(n1013), .B(n44682), .Z(n44731) );
  XOR U44697 ( .A(n44680), .B(n44730), .Z(n44682) );
  XOR U44698 ( .A(n44732), .B(n44733), .Z(n44722) );
  AND U44699 ( .A(n44734), .B(n44735), .Z(n44733) );
  XNOR U44700 ( .A(n44732), .B(n44430), .Z(n44735) );
  IV U44701 ( .A(n44433), .Z(n44430) );
  XOR U44702 ( .A(n44736), .B(n44737), .Z(n44433) );
  AND U44703 ( .A(n1005), .B(n44738), .Z(n44737) );
  XOR U44704 ( .A(n44739), .B(n44736), .Z(n44738) );
  XOR U44705 ( .A(n44434), .B(n44732), .Z(n44734) );
  XOR U44706 ( .A(n44740), .B(n44741), .Z(n44434) );
  AND U44707 ( .A(n1013), .B(n44692), .Z(n44741) );
  XOR U44708 ( .A(n44740), .B(n44690), .Z(n44692) );
  XOR U44709 ( .A(n44742), .B(n44743), .Z(n44732) );
  AND U44710 ( .A(n44744), .B(n44745), .Z(n44743) );
  XNOR U44711 ( .A(n44742), .B(n44458), .Z(n44745) );
  IV U44712 ( .A(n44461), .Z(n44458) );
  XOR U44713 ( .A(n44746), .B(n44747), .Z(n44461) );
  AND U44714 ( .A(n1005), .B(n44748), .Z(n44747) );
  XNOR U44715 ( .A(n44749), .B(n44746), .Z(n44748) );
  XOR U44716 ( .A(n44462), .B(n44742), .Z(n44744) );
  XOR U44717 ( .A(n44750), .B(n44751), .Z(n44462) );
  AND U44718 ( .A(n1013), .B(n44701), .Z(n44751) );
  XOR U44719 ( .A(n44750), .B(n44699), .Z(n44701) );
  XOR U44720 ( .A(n44752), .B(n44753), .Z(n44742) );
  AND U44721 ( .A(n44754), .B(n44755), .Z(n44753) );
  XNOR U44722 ( .A(n44752), .B(n44507), .Z(n44755) );
  IV U44723 ( .A(n44510), .Z(n44507) );
  XOR U44724 ( .A(n44756), .B(n44757), .Z(n44510) );
  AND U44725 ( .A(n1005), .B(n44758), .Z(n44757) );
  XOR U44726 ( .A(n44759), .B(n44756), .Z(n44758) );
  XOR U44727 ( .A(n44511), .B(n44752), .Z(n44754) );
  XOR U44728 ( .A(n44760), .B(n44761), .Z(n44511) );
  AND U44729 ( .A(n1013), .B(n44709), .Z(n44761) );
  XOR U44730 ( .A(n44760), .B(n44707), .Z(n44709) );
  XOR U44731 ( .A(n44648), .B(n44762), .Z(n44752) );
  AND U44732 ( .A(n44650), .B(n44763), .Z(n44762) );
  XNOR U44733 ( .A(n44648), .B(n44604), .Z(n44763) );
  IV U44734 ( .A(n44607), .Z(n44604) );
  XOR U44735 ( .A(n44764), .B(n44765), .Z(n44607) );
  AND U44736 ( .A(n1005), .B(n44766), .Z(n44765) );
  XNOR U44737 ( .A(n44767), .B(n44764), .Z(n44766) );
  XOR U44738 ( .A(n44608), .B(n44648), .Z(n44650) );
  XOR U44739 ( .A(n44768), .B(n44769), .Z(n44608) );
  AND U44740 ( .A(n1013), .B(n44719), .Z(n44769) );
  XOR U44741 ( .A(n44768), .B(n44717), .Z(n44719) );
  AND U44742 ( .A(n44720), .B(n44628), .Z(n44648) );
  XNOR U44743 ( .A(n44770), .B(n44771), .Z(n44628) );
  AND U44744 ( .A(n1005), .B(n44772), .Z(n44771) );
  XNOR U44745 ( .A(n44773), .B(n44770), .Z(n44772) );
  XNOR U44746 ( .A(n44774), .B(n44775), .Z(n1005) );
  AND U44747 ( .A(n44776), .B(n44777), .Z(n44775) );
  XOR U44748 ( .A(n44729), .B(n44774), .Z(n44777) );
  AND U44749 ( .A(n44778), .B(n44779), .Z(n44729) );
  XNOR U44750 ( .A(n44726), .B(n44774), .Z(n44776) );
  XNOR U44751 ( .A(n44780), .B(n44781), .Z(n44726) );
  AND U44752 ( .A(n1009), .B(n44782), .Z(n44781) );
  XNOR U44753 ( .A(n44783), .B(n44784), .Z(n44782) );
  XOR U44754 ( .A(n44785), .B(n44786), .Z(n44774) );
  AND U44755 ( .A(n44787), .B(n44788), .Z(n44786) );
  XNOR U44756 ( .A(n44785), .B(n44778), .Z(n44788) );
  IV U44757 ( .A(n44739), .Z(n44778) );
  XOR U44758 ( .A(n44789), .B(n44790), .Z(n44739) );
  XOR U44759 ( .A(n44791), .B(n44779), .Z(n44790) );
  AND U44760 ( .A(n44749), .B(n44792), .Z(n44779) );
  AND U44761 ( .A(n44793), .B(n44794), .Z(n44791) );
  XOR U44762 ( .A(n44795), .B(n44789), .Z(n44793) );
  XNOR U44763 ( .A(n44736), .B(n44785), .Z(n44787) );
  XNOR U44764 ( .A(n44796), .B(n44797), .Z(n44736) );
  AND U44765 ( .A(n1009), .B(n44798), .Z(n44797) );
  XNOR U44766 ( .A(n44799), .B(n44800), .Z(n44798) );
  XOR U44767 ( .A(n44801), .B(n44802), .Z(n44785) );
  AND U44768 ( .A(n44803), .B(n44804), .Z(n44802) );
  XNOR U44769 ( .A(n44801), .B(n44749), .Z(n44804) );
  XOR U44770 ( .A(n44805), .B(n44794), .Z(n44749) );
  XNOR U44771 ( .A(n44806), .B(n44789), .Z(n44794) );
  XOR U44772 ( .A(n44807), .B(n44808), .Z(n44789) );
  AND U44773 ( .A(n44809), .B(n44810), .Z(n44808) );
  XOR U44774 ( .A(n44811), .B(n44807), .Z(n44809) );
  XNOR U44775 ( .A(n44812), .B(n44813), .Z(n44806) );
  AND U44776 ( .A(n44814), .B(n44815), .Z(n44813) );
  XOR U44777 ( .A(n44812), .B(n44816), .Z(n44814) );
  XNOR U44778 ( .A(n44795), .B(n44792), .Z(n44805) );
  AND U44779 ( .A(n44817), .B(n44818), .Z(n44792) );
  XOR U44780 ( .A(n44819), .B(n44820), .Z(n44795) );
  AND U44781 ( .A(n44821), .B(n44822), .Z(n44820) );
  XOR U44782 ( .A(n44819), .B(n44823), .Z(n44821) );
  XNOR U44783 ( .A(n44746), .B(n44801), .Z(n44803) );
  XNOR U44784 ( .A(n44824), .B(n44825), .Z(n44746) );
  AND U44785 ( .A(n1009), .B(n44826), .Z(n44825) );
  XNOR U44786 ( .A(n44827), .B(n44828), .Z(n44826) );
  XOR U44787 ( .A(n44829), .B(n44830), .Z(n44801) );
  AND U44788 ( .A(n44831), .B(n44832), .Z(n44830) );
  XNOR U44789 ( .A(n44829), .B(n44817), .Z(n44832) );
  IV U44790 ( .A(n44759), .Z(n44817) );
  XNOR U44791 ( .A(n44833), .B(n44810), .Z(n44759) );
  XNOR U44792 ( .A(n44834), .B(n44816), .Z(n44810) );
  XOR U44793 ( .A(n44835), .B(n44836), .Z(n44816) );
  AND U44794 ( .A(n44837), .B(n44838), .Z(n44836) );
  XOR U44795 ( .A(n44835), .B(n44839), .Z(n44837) );
  XNOR U44796 ( .A(n44815), .B(n44807), .Z(n44834) );
  XOR U44797 ( .A(n44840), .B(n44841), .Z(n44807) );
  AND U44798 ( .A(n44842), .B(n44843), .Z(n44841) );
  XNOR U44799 ( .A(n44844), .B(n44840), .Z(n44842) );
  XNOR U44800 ( .A(n44845), .B(n44812), .Z(n44815) );
  XOR U44801 ( .A(n44846), .B(n44847), .Z(n44812) );
  AND U44802 ( .A(n44848), .B(n44849), .Z(n44847) );
  XOR U44803 ( .A(n44846), .B(n44850), .Z(n44848) );
  XNOR U44804 ( .A(n44851), .B(n44852), .Z(n44845) );
  AND U44805 ( .A(n44853), .B(n44854), .Z(n44852) );
  XNOR U44806 ( .A(n44851), .B(n44855), .Z(n44853) );
  XNOR U44807 ( .A(n44811), .B(n44818), .Z(n44833) );
  AND U44808 ( .A(n44767), .B(n44856), .Z(n44818) );
  XOR U44809 ( .A(n44823), .B(n44822), .Z(n44811) );
  XNOR U44810 ( .A(n44857), .B(n44819), .Z(n44822) );
  XOR U44811 ( .A(n44858), .B(n44859), .Z(n44819) );
  AND U44812 ( .A(n44860), .B(n44861), .Z(n44859) );
  XOR U44813 ( .A(n44858), .B(n44862), .Z(n44860) );
  XNOR U44814 ( .A(n44863), .B(n44864), .Z(n44857) );
  AND U44815 ( .A(n44865), .B(n44866), .Z(n44864) );
  XOR U44816 ( .A(n44863), .B(n44867), .Z(n44865) );
  XOR U44817 ( .A(n44868), .B(n44869), .Z(n44823) );
  AND U44818 ( .A(n44870), .B(n44871), .Z(n44869) );
  XOR U44819 ( .A(n44868), .B(n44872), .Z(n44870) );
  XNOR U44820 ( .A(n44756), .B(n44829), .Z(n44831) );
  XNOR U44821 ( .A(n44873), .B(n44874), .Z(n44756) );
  AND U44822 ( .A(n1009), .B(n44875), .Z(n44874) );
  XNOR U44823 ( .A(n44876), .B(n44877), .Z(n44875) );
  XOR U44824 ( .A(n44878), .B(n44879), .Z(n44829) );
  AND U44825 ( .A(n44880), .B(n44881), .Z(n44879) );
  XNOR U44826 ( .A(n44878), .B(n44767), .Z(n44881) );
  XOR U44827 ( .A(n44882), .B(n44843), .Z(n44767) );
  XNOR U44828 ( .A(n44883), .B(n44850), .Z(n44843) );
  XOR U44829 ( .A(n44839), .B(n44838), .Z(n44850) );
  XNOR U44830 ( .A(n44884), .B(n44835), .Z(n44838) );
  XOR U44831 ( .A(n44885), .B(n44886), .Z(n44835) );
  AND U44832 ( .A(n44887), .B(n44888), .Z(n44886) );
  XNOR U44833 ( .A(n44889), .B(n44890), .Z(n44887) );
  IV U44834 ( .A(n44885), .Z(n44889) );
  XNOR U44835 ( .A(n44891), .B(n44892), .Z(n44884) );
  NOR U44836 ( .A(n44893), .B(n44894), .Z(n44892) );
  XNOR U44837 ( .A(n44891), .B(n44895), .Z(n44893) );
  XOR U44838 ( .A(n44896), .B(n44897), .Z(n44839) );
  NOR U44839 ( .A(n44898), .B(n44899), .Z(n44897) );
  XNOR U44840 ( .A(n44896), .B(n44900), .Z(n44898) );
  XNOR U44841 ( .A(n44849), .B(n44840), .Z(n44883) );
  XOR U44842 ( .A(n44901), .B(n44902), .Z(n44840) );
  AND U44843 ( .A(n44903), .B(n44904), .Z(n44902) );
  XOR U44844 ( .A(n44901), .B(n44905), .Z(n44903) );
  XOR U44845 ( .A(n44906), .B(n44855), .Z(n44849) );
  XOR U44846 ( .A(n44907), .B(n44908), .Z(n44855) );
  NOR U44847 ( .A(n44909), .B(n44910), .Z(n44908) );
  XOR U44848 ( .A(n44907), .B(n44911), .Z(n44909) );
  XNOR U44849 ( .A(n44854), .B(n44846), .Z(n44906) );
  XOR U44850 ( .A(n44912), .B(n44913), .Z(n44846) );
  AND U44851 ( .A(n44914), .B(n44915), .Z(n44913) );
  XOR U44852 ( .A(n44912), .B(n44916), .Z(n44914) );
  XNOR U44853 ( .A(n44917), .B(n44851), .Z(n44854) );
  XOR U44854 ( .A(n44918), .B(n44919), .Z(n44851) );
  AND U44855 ( .A(n44920), .B(n44921), .Z(n44919) );
  XNOR U44856 ( .A(n44922), .B(n44923), .Z(n44920) );
  IV U44857 ( .A(n44918), .Z(n44922) );
  XNOR U44858 ( .A(n44924), .B(n44925), .Z(n44917) );
  NOR U44859 ( .A(n44926), .B(n44927), .Z(n44925) );
  XNOR U44860 ( .A(n44924), .B(n44928), .Z(n44926) );
  XOR U44861 ( .A(n44844), .B(n44856), .Z(n44882) );
  NOR U44862 ( .A(n44773), .B(n44929), .Z(n44856) );
  XNOR U44863 ( .A(n44862), .B(n44861), .Z(n44844) );
  XNOR U44864 ( .A(n44930), .B(n44867), .Z(n44861) );
  XNOR U44865 ( .A(n44931), .B(n44932), .Z(n44867) );
  NOR U44866 ( .A(n44933), .B(n44934), .Z(n44932) );
  XOR U44867 ( .A(n44931), .B(n44935), .Z(n44933) );
  XNOR U44868 ( .A(n44866), .B(n44858), .Z(n44930) );
  XOR U44869 ( .A(n44936), .B(n44937), .Z(n44858) );
  AND U44870 ( .A(n44938), .B(n44939), .Z(n44937) );
  XOR U44871 ( .A(n44936), .B(n44940), .Z(n44938) );
  XNOR U44872 ( .A(n44941), .B(n44863), .Z(n44866) );
  XOR U44873 ( .A(n44942), .B(n44943), .Z(n44863) );
  AND U44874 ( .A(n44944), .B(n44945), .Z(n44943) );
  XNOR U44875 ( .A(n44946), .B(n44947), .Z(n44944) );
  IV U44876 ( .A(n44942), .Z(n44946) );
  XNOR U44877 ( .A(n44948), .B(n44949), .Z(n44941) );
  NOR U44878 ( .A(n44950), .B(n44951), .Z(n44949) );
  XNOR U44879 ( .A(n44948), .B(n44952), .Z(n44950) );
  XOR U44880 ( .A(n44872), .B(n44871), .Z(n44862) );
  XNOR U44881 ( .A(n44953), .B(n44868), .Z(n44871) );
  XOR U44882 ( .A(n44954), .B(n44955), .Z(n44868) );
  AND U44883 ( .A(n44956), .B(n44957), .Z(n44955) );
  XNOR U44884 ( .A(n44958), .B(n44959), .Z(n44956) );
  IV U44885 ( .A(n44954), .Z(n44958) );
  XNOR U44886 ( .A(n44960), .B(n44961), .Z(n44953) );
  NOR U44887 ( .A(n44962), .B(n44963), .Z(n44961) );
  XNOR U44888 ( .A(n44960), .B(n44964), .Z(n44962) );
  XOR U44889 ( .A(n44965), .B(n44966), .Z(n44872) );
  NOR U44890 ( .A(n44967), .B(n44968), .Z(n44966) );
  XNOR U44891 ( .A(n44965), .B(n44969), .Z(n44967) );
  XNOR U44892 ( .A(n44764), .B(n44878), .Z(n44880) );
  XNOR U44893 ( .A(n44970), .B(n44971), .Z(n44764) );
  AND U44894 ( .A(n1009), .B(n44972), .Z(n44971) );
  XNOR U44895 ( .A(n44973), .B(n44974), .Z(n44972) );
  AND U44896 ( .A(n44770), .B(n44773), .Z(n44878) );
  XOR U44897 ( .A(n44975), .B(n44929), .Z(n44773) );
  XNOR U44898 ( .A(p_input[1472]), .B(p_input[2048]), .Z(n44929) );
  XNOR U44899 ( .A(n44905), .B(n44904), .Z(n44975) );
  XNOR U44900 ( .A(n44976), .B(n44916), .Z(n44904) );
  XOR U44901 ( .A(n44890), .B(n44888), .Z(n44916) );
  XNOR U44902 ( .A(n44977), .B(n44895), .Z(n44888) );
  XOR U44903 ( .A(p_input[1496]), .B(p_input[2072]), .Z(n44895) );
  XOR U44904 ( .A(n44885), .B(n44894), .Z(n44977) );
  XOR U44905 ( .A(n44978), .B(n44891), .Z(n44894) );
  XOR U44906 ( .A(p_input[1494]), .B(p_input[2070]), .Z(n44891) );
  XOR U44907 ( .A(p_input[1495]), .B(n29410), .Z(n44978) );
  XOR U44908 ( .A(p_input[1490]), .B(p_input[2066]), .Z(n44885) );
  XNOR U44909 ( .A(n44900), .B(n44899), .Z(n44890) );
  XOR U44910 ( .A(n44979), .B(n44896), .Z(n44899) );
  XOR U44911 ( .A(p_input[1491]), .B(p_input[2067]), .Z(n44896) );
  XOR U44912 ( .A(p_input[1492]), .B(n29412), .Z(n44979) );
  XOR U44913 ( .A(p_input[1493]), .B(p_input[2069]), .Z(n44900) );
  XOR U44914 ( .A(n44915), .B(n44980), .Z(n44976) );
  IV U44915 ( .A(n44901), .Z(n44980) );
  XOR U44916 ( .A(p_input[1473]), .B(p_input[2049]), .Z(n44901) );
  XNOR U44917 ( .A(n44981), .B(n44923), .Z(n44915) );
  XNOR U44918 ( .A(n44911), .B(n44910), .Z(n44923) );
  XNOR U44919 ( .A(n44982), .B(n44907), .Z(n44910) );
  XNOR U44920 ( .A(p_input[1498]), .B(p_input[2074]), .Z(n44907) );
  XOR U44921 ( .A(p_input[1499]), .B(n29415), .Z(n44982) );
  XOR U44922 ( .A(p_input[1500]), .B(p_input[2076]), .Z(n44911) );
  XOR U44923 ( .A(n44921), .B(n44983), .Z(n44981) );
  IV U44924 ( .A(n44912), .Z(n44983) );
  XOR U44925 ( .A(p_input[1489]), .B(p_input[2065]), .Z(n44912) );
  XNOR U44926 ( .A(n44984), .B(n44928), .Z(n44921) );
  XNOR U44927 ( .A(p_input[1503]), .B(n29418), .Z(n44928) );
  XOR U44928 ( .A(n44918), .B(n44927), .Z(n44984) );
  XOR U44929 ( .A(n44985), .B(n44924), .Z(n44927) );
  XOR U44930 ( .A(p_input[1501]), .B(p_input[2077]), .Z(n44924) );
  XOR U44931 ( .A(p_input[1502]), .B(n29420), .Z(n44985) );
  XOR U44932 ( .A(p_input[1497]), .B(p_input[2073]), .Z(n44918) );
  XOR U44933 ( .A(n44940), .B(n44939), .Z(n44905) );
  XNOR U44934 ( .A(n44986), .B(n44947), .Z(n44939) );
  XNOR U44935 ( .A(n44935), .B(n44934), .Z(n44947) );
  XNOR U44936 ( .A(n44987), .B(n44931), .Z(n44934) );
  XNOR U44937 ( .A(p_input[1483]), .B(p_input[2059]), .Z(n44931) );
  XOR U44938 ( .A(p_input[1484]), .B(n28329), .Z(n44987) );
  XOR U44939 ( .A(p_input[1485]), .B(p_input[2061]), .Z(n44935) );
  XOR U44940 ( .A(n44945), .B(n44988), .Z(n44986) );
  IV U44941 ( .A(n44936), .Z(n44988) );
  XOR U44942 ( .A(p_input[1474]), .B(p_input[2050]), .Z(n44936) );
  XNOR U44943 ( .A(n44989), .B(n44952), .Z(n44945) );
  XNOR U44944 ( .A(p_input[1488]), .B(n28332), .Z(n44952) );
  XOR U44945 ( .A(n44942), .B(n44951), .Z(n44989) );
  XOR U44946 ( .A(n44990), .B(n44948), .Z(n44951) );
  XOR U44947 ( .A(p_input[1486]), .B(p_input[2062]), .Z(n44948) );
  XOR U44948 ( .A(p_input[1487]), .B(n28334), .Z(n44990) );
  XOR U44949 ( .A(p_input[1482]), .B(p_input[2058]), .Z(n44942) );
  XOR U44950 ( .A(n44959), .B(n44957), .Z(n44940) );
  XNOR U44951 ( .A(n44991), .B(n44964), .Z(n44957) );
  XOR U44952 ( .A(p_input[1481]), .B(p_input[2057]), .Z(n44964) );
  XOR U44953 ( .A(n44954), .B(n44963), .Z(n44991) );
  XOR U44954 ( .A(n44992), .B(n44960), .Z(n44963) );
  XOR U44955 ( .A(p_input[1479]), .B(p_input[2055]), .Z(n44960) );
  XOR U44956 ( .A(p_input[1480]), .B(n29427), .Z(n44992) );
  XOR U44957 ( .A(p_input[1475]), .B(p_input[2051]), .Z(n44954) );
  XNOR U44958 ( .A(n44969), .B(n44968), .Z(n44959) );
  XOR U44959 ( .A(n44993), .B(n44965), .Z(n44968) );
  XOR U44960 ( .A(p_input[1476]), .B(p_input[2052]), .Z(n44965) );
  XOR U44961 ( .A(p_input[1477]), .B(n29429), .Z(n44993) );
  XOR U44962 ( .A(p_input[1478]), .B(p_input[2054]), .Z(n44969) );
  XNOR U44963 ( .A(n44994), .B(n44995), .Z(n44770) );
  AND U44964 ( .A(n1009), .B(n44996), .Z(n44995) );
  XNOR U44965 ( .A(n44997), .B(n44998), .Z(n1009) );
  AND U44966 ( .A(n44999), .B(n45000), .Z(n44998) );
  XOR U44967 ( .A(n44784), .B(n44997), .Z(n45000) );
  XNOR U44968 ( .A(n45001), .B(n44997), .Z(n44999) );
  XOR U44969 ( .A(n45002), .B(n45003), .Z(n44997) );
  AND U44970 ( .A(n45004), .B(n45005), .Z(n45003) );
  XOR U44971 ( .A(n44799), .B(n45002), .Z(n45005) );
  XOR U44972 ( .A(n45002), .B(n44800), .Z(n45004) );
  XOR U44973 ( .A(n45006), .B(n45007), .Z(n45002) );
  AND U44974 ( .A(n45008), .B(n45009), .Z(n45007) );
  XOR U44975 ( .A(n44827), .B(n45006), .Z(n45009) );
  XOR U44976 ( .A(n45006), .B(n44828), .Z(n45008) );
  XOR U44977 ( .A(n45010), .B(n45011), .Z(n45006) );
  AND U44978 ( .A(n45012), .B(n45013), .Z(n45011) );
  XOR U44979 ( .A(n44876), .B(n45010), .Z(n45013) );
  XOR U44980 ( .A(n45010), .B(n44877), .Z(n45012) );
  XOR U44981 ( .A(n45014), .B(n45015), .Z(n45010) );
  AND U44982 ( .A(n45016), .B(n45017), .Z(n45015) );
  XOR U44983 ( .A(n45014), .B(n44973), .Z(n45017) );
  XNOR U44984 ( .A(n45018), .B(n45019), .Z(n44720) );
  AND U44985 ( .A(n1013), .B(n45020), .Z(n45019) );
  XNOR U44986 ( .A(n45021), .B(n45022), .Z(n1013) );
  AND U44987 ( .A(n45023), .B(n45024), .Z(n45022) );
  XOR U44988 ( .A(n45021), .B(n44730), .Z(n45024) );
  XNOR U44989 ( .A(n45021), .B(n44680), .Z(n45023) );
  XOR U44990 ( .A(n45025), .B(n45026), .Z(n45021) );
  AND U44991 ( .A(n45027), .B(n45028), .Z(n45026) );
  XNOR U44992 ( .A(n44740), .B(n45025), .Z(n45028) );
  XOR U44993 ( .A(n45025), .B(n44690), .Z(n45027) );
  XOR U44994 ( .A(n45029), .B(n45030), .Z(n45025) );
  AND U44995 ( .A(n45031), .B(n45032), .Z(n45030) );
  XNOR U44996 ( .A(n44750), .B(n45029), .Z(n45032) );
  XOR U44997 ( .A(n45029), .B(n44699), .Z(n45031) );
  XOR U44998 ( .A(n45033), .B(n45034), .Z(n45029) );
  AND U44999 ( .A(n45035), .B(n45036), .Z(n45034) );
  XOR U45000 ( .A(n45033), .B(n44707), .Z(n45035) );
  XOR U45001 ( .A(n45037), .B(n45038), .Z(n44671) );
  AND U45002 ( .A(n1017), .B(n45020), .Z(n45038) );
  XNOR U45003 ( .A(n45018), .B(n45037), .Z(n45020) );
  XNOR U45004 ( .A(n45039), .B(n45040), .Z(n1017) );
  AND U45005 ( .A(n45041), .B(n45042), .Z(n45040) );
  XNOR U45006 ( .A(n45043), .B(n45039), .Z(n45042) );
  IV U45007 ( .A(n44730), .Z(n45043) );
  XOR U45008 ( .A(n45001), .B(n45044), .Z(n44730) );
  AND U45009 ( .A(n1020), .B(n45045), .Z(n45044) );
  XOR U45010 ( .A(n44783), .B(n44780), .Z(n45045) );
  IV U45011 ( .A(n45001), .Z(n44783) );
  XNOR U45012 ( .A(n44680), .B(n45039), .Z(n45041) );
  XOR U45013 ( .A(n45046), .B(n45047), .Z(n44680) );
  AND U45014 ( .A(n1036), .B(n45048), .Z(n45047) );
  XOR U45015 ( .A(n45049), .B(n45050), .Z(n45039) );
  AND U45016 ( .A(n45051), .B(n45052), .Z(n45050) );
  XNOR U45017 ( .A(n45049), .B(n44740), .Z(n45052) );
  XOR U45018 ( .A(n44800), .B(n45053), .Z(n44740) );
  AND U45019 ( .A(n1020), .B(n45054), .Z(n45053) );
  XOR U45020 ( .A(n44796), .B(n44800), .Z(n45054) );
  XNOR U45021 ( .A(n45055), .B(n45049), .Z(n45051) );
  IV U45022 ( .A(n44690), .Z(n45055) );
  XOR U45023 ( .A(n45056), .B(n45057), .Z(n44690) );
  AND U45024 ( .A(n1036), .B(n45058), .Z(n45057) );
  XOR U45025 ( .A(n45059), .B(n45060), .Z(n45049) );
  AND U45026 ( .A(n45061), .B(n45062), .Z(n45060) );
  XNOR U45027 ( .A(n45059), .B(n44750), .Z(n45062) );
  XOR U45028 ( .A(n44828), .B(n45063), .Z(n44750) );
  AND U45029 ( .A(n1020), .B(n45064), .Z(n45063) );
  XOR U45030 ( .A(n44824), .B(n44828), .Z(n45064) );
  XOR U45031 ( .A(n44699), .B(n45059), .Z(n45061) );
  XOR U45032 ( .A(n45065), .B(n45066), .Z(n44699) );
  AND U45033 ( .A(n1036), .B(n45067), .Z(n45066) );
  XOR U45034 ( .A(n45033), .B(n45068), .Z(n45059) );
  AND U45035 ( .A(n45069), .B(n45036), .Z(n45068) );
  XNOR U45036 ( .A(n44760), .B(n45033), .Z(n45036) );
  XOR U45037 ( .A(n44877), .B(n45070), .Z(n44760) );
  AND U45038 ( .A(n1020), .B(n45071), .Z(n45070) );
  XOR U45039 ( .A(n44873), .B(n44877), .Z(n45071) );
  XNOR U45040 ( .A(n45072), .B(n45033), .Z(n45069) );
  IV U45041 ( .A(n44707), .Z(n45072) );
  XOR U45042 ( .A(n45073), .B(n45074), .Z(n44707) );
  AND U45043 ( .A(n1036), .B(n45075), .Z(n45074) );
  XOR U45044 ( .A(n45076), .B(n45077), .Z(n45033) );
  AND U45045 ( .A(n45078), .B(n45079), .Z(n45077) );
  XNOR U45046 ( .A(n45076), .B(n44768), .Z(n45079) );
  XOR U45047 ( .A(n44974), .B(n45080), .Z(n44768) );
  AND U45048 ( .A(n1020), .B(n45081), .Z(n45080) );
  XOR U45049 ( .A(n44970), .B(n44974), .Z(n45081) );
  XNOR U45050 ( .A(n45082), .B(n45076), .Z(n45078) );
  IV U45051 ( .A(n44717), .Z(n45082) );
  XOR U45052 ( .A(n45083), .B(n45084), .Z(n44717) );
  AND U45053 ( .A(n1036), .B(n45085), .Z(n45084) );
  AND U45054 ( .A(n45037), .B(n45018), .Z(n45076) );
  XNOR U45055 ( .A(n45086), .B(n45087), .Z(n45018) );
  AND U45056 ( .A(n1020), .B(n44996), .Z(n45087) );
  XNOR U45057 ( .A(n44994), .B(n45086), .Z(n44996) );
  XNOR U45058 ( .A(n45088), .B(n45089), .Z(n1020) );
  AND U45059 ( .A(n45090), .B(n45091), .Z(n45089) );
  XNOR U45060 ( .A(n45088), .B(n44780), .Z(n45091) );
  IV U45061 ( .A(n44784), .Z(n44780) );
  XOR U45062 ( .A(n45092), .B(n45093), .Z(n44784) );
  AND U45063 ( .A(n1024), .B(n45094), .Z(n45093) );
  XOR U45064 ( .A(n45095), .B(n45092), .Z(n45094) );
  XNOR U45065 ( .A(n45088), .B(n45001), .Z(n45090) );
  XOR U45066 ( .A(n45096), .B(n45097), .Z(n45001) );
  AND U45067 ( .A(n1032), .B(n45048), .Z(n45097) );
  XOR U45068 ( .A(n45046), .B(n45096), .Z(n45048) );
  XOR U45069 ( .A(n45098), .B(n45099), .Z(n45088) );
  AND U45070 ( .A(n45100), .B(n45101), .Z(n45099) );
  XNOR U45071 ( .A(n45098), .B(n44796), .Z(n45101) );
  IV U45072 ( .A(n44799), .Z(n44796) );
  XOR U45073 ( .A(n45102), .B(n45103), .Z(n44799) );
  AND U45074 ( .A(n1024), .B(n45104), .Z(n45103) );
  XOR U45075 ( .A(n45105), .B(n45102), .Z(n45104) );
  XOR U45076 ( .A(n44800), .B(n45098), .Z(n45100) );
  XOR U45077 ( .A(n45106), .B(n45107), .Z(n44800) );
  AND U45078 ( .A(n1032), .B(n45058), .Z(n45107) );
  XOR U45079 ( .A(n45106), .B(n45056), .Z(n45058) );
  XOR U45080 ( .A(n45108), .B(n45109), .Z(n45098) );
  AND U45081 ( .A(n45110), .B(n45111), .Z(n45109) );
  XNOR U45082 ( .A(n45108), .B(n44824), .Z(n45111) );
  IV U45083 ( .A(n44827), .Z(n44824) );
  XOR U45084 ( .A(n45112), .B(n45113), .Z(n44827) );
  AND U45085 ( .A(n1024), .B(n45114), .Z(n45113) );
  XNOR U45086 ( .A(n45115), .B(n45112), .Z(n45114) );
  XOR U45087 ( .A(n44828), .B(n45108), .Z(n45110) );
  XOR U45088 ( .A(n45116), .B(n45117), .Z(n44828) );
  AND U45089 ( .A(n1032), .B(n45067), .Z(n45117) );
  XOR U45090 ( .A(n45116), .B(n45065), .Z(n45067) );
  XOR U45091 ( .A(n45118), .B(n45119), .Z(n45108) );
  AND U45092 ( .A(n45120), .B(n45121), .Z(n45119) );
  XNOR U45093 ( .A(n45118), .B(n44873), .Z(n45121) );
  IV U45094 ( .A(n44876), .Z(n44873) );
  XOR U45095 ( .A(n45122), .B(n45123), .Z(n44876) );
  AND U45096 ( .A(n1024), .B(n45124), .Z(n45123) );
  XOR U45097 ( .A(n45125), .B(n45122), .Z(n45124) );
  XOR U45098 ( .A(n44877), .B(n45118), .Z(n45120) );
  XOR U45099 ( .A(n45126), .B(n45127), .Z(n44877) );
  AND U45100 ( .A(n1032), .B(n45075), .Z(n45127) );
  XOR U45101 ( .A(n45126), .B(n45073), .Z(n45075) );
  XOR U45102 ( .A(n45014), .B(n45128), .Z(n45118) );
  AND U45103 ( .A(n45016), .B(n45129), .Z(n45128) );
  XNOR U45104 ( .A(n45014), .B(n44970), .Z(n45129) );
  IV U45105 ( .A(n44973), .Z(n44970) );
  XOR U45106 ( .A(n45130), .B(n45131), .Z(n44973) );
  AND U45107 ( .A(n1024), .B(n45132), .Z(n45131) );
  XNOR U45108 ( .A(n45133), .B(n45130), .Z(n45132) );
  XOR U45109 ( .A(n44974), .B(n45014), .Z(n45016) );
  XOR U45110 ( .A(n45134), .B(n45135), .Z(n44974) );
  AND U45111 ( .A(n1032), .B(n45085), .Z(n45135) );
  XOR U45112 ( .A(n45134), .B(n45083), .Z(n45085) );
  AND U45113 ( .A(n45086), .B(n44994), .Z(n45014) );
  XNOR U45114 ( .A(n45136), .B(n45137), .Z(n44994) );
  AND U45115 ( .A(n1024), .B(n45138), .Z(n45137) );
  XNOR U45116 ( .A(n45139), .B(n45136), .Z(n45138) );
  XNOR U45117 ( .A(n45140), .B(n45141), .Z(n1024) );
  AND U45118 ( .A(n45142), .B(n45143), .Z(n45141) );
  XOR U45119 ( .A(n45095), .B(n45140), .Z(n45143) );
  AND U45120 ( .A(n45144), .B(n45145), .Z(n45095) );
  XNOR U45121 ( .A(n45092), .B(n45140), .Z(n45142) );
  XNOR U45122 ( .A(n45146), .B(n45147), .Z(n45092) );
  AND U45123 ( .A(n1028), .B(n45148), .Z(n45147) );
  XNOR U45124 ( .A(n45149), .B(n45150), .Z(n45148) );
  XOR U45125 ( .A(n45151), .B(n45152), .Z(n45140) );
  AND U45126 ( .A(n45153), .B(n45154), .Z(n45152) );
  XNOR U45127 ( .A(n45151), .B(n45144), .Z(n45154) );
  IV U45128 ( .A(n45105), .Z(n45144) );
  XOR U45129 ( .A(n45155), .B(n45156), .Z(n45105) );
  XOR U45130 ( .A(n45157), .B(n45145), .Z(n45156) );
  AND U45131 ( .A(n45115), .B(n45158), .Z(n45145) );
  AND U45132 ( .A(n45159), .B(n45160), .Z(n45157) );
  XOR U45133 ( .A(n45161), .B(n45155), .Z(n45159) );
  XNOR U45134 ( .A(n45102), .B(n45151), .Z(n45153) );
  XNOR U45135 ( .A(n45162), .B(n45163), .Z(n45102) );
  AND U45136 ( .A(n1028), .B(n45164), .Z(n45163) );
  XNOR U45137 ( .A(n45165), .B(n45166), .Z(n45164) );
  XOR U45138 ( .A(n45167), .B(n45168), .Z(n45151) );
  AND U45139 ( .A(n45169), .B(n45170), .Z(n45168) );
  XNOR U45140 ( .A(n45167), .B(n45115), .Z(n45170) );
  XOR U45141 ( .A(n45171), .B(n45160), .Z(n45115) );
  XNOR U45142 ( .A(n45172), .B(n45155), .Z(n45160) );
  XOR U45143 ( .A(n45173), .B(n45174), .Z(n45155) );
  AND U45144 ( .A(n45175), .B(n45176), .Z(n45174) );
  XOR U45145 ( .A(n45177), .B(n45173), .Z(n45175) );
  XNOR U45146 ( .A(n45178), .B(n45179), .Z(n45172) );
  AND U45147 ( .A(n45180), .B(n45181), .Z(n45179) );
  XOR U45148 ( .A(n45178), .B(n45182), .Z(n45180) );
  XNOR U45149 ( .A(n45161), .B(n45158), .Z(n45171) );
  AND U45150 ( .A(n45183), .B(n45184), .Z(n45158) );
  XOR U45151 ( .A(n45185), .B(n45186), .Z(n45161) );
  AND U45152 ( .A(n45187), .B(n45188), .Z(n45186) );
  XOR U45153 ( .A(n45185), .B(n45189), .Z(n45187) );
  XNOR U45154 ( .A(n45112), .B(n45167), .Z(n45169) );
  XNOR U45155 ( .A(n45190), .B(n45191), .Z(n45112) );
  AND U45156 ( .A(n1028), .B(n45192), .Z(n45191) );
  XNOR U45157 ( .A(n45193), .B(n45194), .Z(n45192) );
  XOR U45158 ( .A(n45195), .B(n45196), .Z(n45167) );
  AND U45159 ( .A(n45197), .B(n45198), .Z(n45196) );
  XNOR U45160 ( .A(n45195), .B(n45183), .Z(n45198) );
  IV U45161 ( .A(n45125), .Z(n45183) );
  XNOR U45162 ( .A(n45199), .B(n45176), .Z(n45125) );
  XNOR U45163 ( .A(n45200), .B(n45182), .Z(n45176) );
  XOR U45164 ( .A(n45201), .B(n45202), .Z(n45182) );
  AND U45165 ( .A(n45203), .B(n45204), .Z(n45202) );
  XOR U45166 ( .A(n45201), .B(n45205), .Z(n45203) );
  XNOR U45167 ( .A(n45181), .B(n45173), .Z(n45200) );
  XOR U45168 ( .A(n45206), .B(n45207), .Z(n45173) );
  AND U45169 ( .A(n45208), .B(n45209), .Z(n45207) );
  XNOR U45170 ( .A(n45210), .B(n45206), .Z(n45208) );
  XNOR U45171 ( .A(n45211), .B(n45178), .Z(n45181) );
  XOR U45172 ( .A(n45212), .B(n45213), .Z(n45178) );
  AND U45173 ( .A(n45214), .B(n45215), .Z(n45213) );
  XOR U45174 ( .A(n45212), .B(n45216), .Z(n45214) );
  XNOR U45175 ( .A(n45217), .B(n45218), .Z(n45211) );
  AND U45176 ( .A(n45219), .B(n45220), .Z(n45218) );
  XNOR U45177 ( .A(n45217), .B(n45221), .Z(n45219) );
  XNOR U45178 ( .A(n45177), .B(n45184), .Z(n45199) );
  AND U45179 ( .A(n45133), .B(n45222), .Z(n45184) );
  XOR U45180 ( .A(n45189), .B(n45188), .Z(n45177) );
  XNOR U45181 ( .A(n45223), .B(n45185), .Z(n45188) );
  XOR U45182 ( .A(n45224), .B(n45225), .Z(n45185) );
  AND U45183 ( .A(n45226), .B(n45227), .Z(n45225) );
  XOR U45184 ( .A(n45224), .B(n45228), .Z(n45226) );
  XNOR U45185 ( .A(n45229), .B(n45230), .Z(n45223) );
  AND U45186 ( .A(n45231), .B(n45232), .Z(n45230) );
  XOR U45187 ( .A(n45229), .B(n45233), .Z(n45231) );
  XOR U45188 ( .A(n45234), .B(n45235), .Z(n45189) );
  AND U45189 ( .A(n45236), .B(n45237), .Z(n45235) );
  XOR U45190 ( .A(n45234), .B(n45238), .Z(n45236) );
  XNOR U45191 ( .A(n45122), .B(n45195), .Z(n45197) );
  XNOR U45192 ( .A(n45239), .B(n45240), .Z(n45122) );
  AND U45193 ( .A(n1028), .B(n45241), .Z(n45240) );
  XNOR U45194 ( .A(n45242), .B(n45243), .Z(n45241) );
  XOR U45195 ( .A(n45244), .B(n45245), .Z(n45195) );
  AND U45196 ( .A(n45246), .B(n45247), .Z(n45245) );
  XNOR U45197 ( .A(n45244), .B(n45133), .Z(n45247) );
  XOR U45198 ( .A(n45248), .B(n45209), .Z(n45133) );
  XNOR U45199 ( .A(n45249), .B(n45216), .Z(n45209) );
  XOR U45200 ( .A(n45205), .B(n45204), .Z(n45216) );
  XNOR U45201 ( .A(n45250), .B(n45201), .Z(n45204) );
  XOR U45202 ( .A(n45251), .B(n45252), .Z(n45201) );
  AND U45203 ( .A(n45253), .B(n45254), .Z(n45252) );
  XNOR U45204 ( .A(n45255), .B(n45256), .Z(n45253) );
  IV U45205 ( .A(n45251), .Z(n45255) );
  XNOR U45206 ( .A(n45257), .B(n45258), .Z(n45250) );
  NOR U45207 ( .A(n45259), .B(n45260), .Z(n45258) );
  XNOR U45208 ( .A(n45257), .B(n45261), .Z(n45259) );
  XOR U45209 ( .A(n45262), .B(n45263), .Z(n45205) );
  NOR U45210 ( .A(n45264), .B(n45265), .Z(n45263) );
  XNOR U45211 ( .A(n45262), .B(n45266), .Z(n45264) );
  XNOR U45212 ( .A(n45215), .B(n45206), .Z(n45249) );
  XOR U45213 ( .A(n45267), .B(n45268), .Z(n45206) );
  AND U45214 ( .A(n45269), .B(n45270), .Z(n45268) );
  XOR U45215 ( .A(n45267), .B(n45271), .Z(n45269) );
  XOR U45216 ( .A(n45272), .B(n45221), .Z(n45215) );
  XOR U45217 ( .A(n45273), .B(n45274), .Z(n45221) );
  NOR U45218 ( .A(n45275), .B(n45276), .Z(n45274) );
  XOR U45219 ( .A(n45273), .B(n45277), .Z(n45275) );
  XNOR U45220 ( .A(n45220), .B(n45212), .Z(n45272) );
  XOR U45221 ( .A(n45278), .B(n45279), .Z(n45212) );
  AND U45222 ( .A(n45280), .B(n45281), .Z(n45279) );
  XOR U45223 ( .A(n45278), .B(n45282), .Z(n45280) );
  XNOR U45224 ( .A(n45283), .B(n45217), .Z(n45220) );
  XOR U45225 ( .A(n45284), .B(n45285), .Z(n45217) );
  AND U45226 ( .A(n45286), .B(n45287), .Z(n45285) );
  XNOR U45227 ( .A(n45288), .B(n45289), .Z(n45286) );
  IV U45228 ( .A(n45284), .Z(n45288) );
  XNOR U45229 ( .A(n45290), .B(n45291), .Z(n45283) );
  NOR U45230 ( .A(n45292), .B(n45293), .Z(n45291) );
  XNOR U45231 ( .A(n45290), .B(n45294), .Z(n45292) );
  XOR U45232 ( .A(n45210), .B(n45222), .Z(n45248) );
  NOR U45233 ( .A(n45139), .B(n45295), .Z(n45222) );
  XNOR U45234 ( .A(n45228), .B(n45227), .Z(n45210) );
  XNOR U45235 ( .A(n45296), .B(n45233), .Z(n45227) );
  XNOR U45236 ( .A(n45297), .B(n45298), .Z(n45233) );
  NOR U45237 ( .A(n45299), .B(n45300), .Z(n45298) );
  XOR U45238 ( .A(n45297), .B(n45301), .Z(n45299) );
  XNOR U45239 ( .A(n45232), .B(n45224), .Z(n45296) );
  XOR U45240 ( .A(n45302), .B(n45303), .Z(n45224) );
  AND U45241 ( .A(n45304), .B(n45305), .Z(n45303) );
  XOR U45242 ( .A(n45302), .B(n45306), .Z(n45304) );
  XNOR U45243 ( .A(n45307), .B(n45229), .Z(n45232) );
  XOR U45244 ( .A(n45308), .B(n45309), .Z(n45229) );
  AND U45245 ( .A(n45310), .B(n45311), .Z(n45309) );
  XNOR U45246 ( .A(n45312), .B(n45313), .Z(n45310) );
  IV U45247 ( .A(n45308), .Z(n45312) );
  XNOR U45248 ( .A(n45314), .B(n45315), .Z(n45307) );
  NOR U45249 ( .A(n45316), .B(n45317), .Z(n45315) );
  XNOR U45250 ( .A(n45314), .B(n45318), .Z(n45316) );
  XOR U45251 ( .A(n45238), .B(n45237), .Z(n45228) );
  XNOR U45252 ( .A(n45319), .B(n45234), .Z(n45237) );
  XOR U45253 ( .A(n45320), .B(n45321), .Z(n45234) );
  AND U45254 ( .A(n45322), .B(n45323), .Z(n45321) );
  XNOR U45255 ( .A(n45324), .B(n45325), .Z(n45322) );
  IV U45256 ( .A(n45320), .Z(n45324) );
  XNOR U45257 ( .A(n45326), .B(n45327), .Z(n45319) );
  NOR U45258 ( .A(n45328), .B(n45329), .Z(n45327) );
  XNOR U45259 ( .A(n45326), .B(n45330), .Z(n45328) );
  XOR U45260 ( .A(n45331), .B(n45332), .Z(n45238) );
  NOR U45261 ( .A(n45333), .B(n45334), .Z(n45332) );
  XNOR U45262 ( .A(n45331), .B(n45335), .Z(n45333) );
  XNOR U45263 ( .A(n45130), .B(n45244), .Z(n45246) );
  XNOR U45264 ( .A(n45336), .B(n45337), .Z(n45130) );
  AND U45265 ( .A(n1028), .B(n45338), .Z(n45337) );
  XNOR U45266 ( .A(n45339), .B(n45340), .Z(n45338) );
  AND U45267 ( .A(n45136), .B(n45139), .Z(n45244) );
  XOR U45268 ( .A(n45341), .B(n45295), .Z(n45139) );
  XNOR U45269 ( .A(p_input[1504]), .B(p_input[2048]), .Z(n45295) );
  XNOR U45270 ( .A(n45271), .B(n45270), .Z(n45341) );
  XNOR U45271 ( .A(n45342), .B(n45282), .Z(n45270) );
  XOR U45272 ( .A(n45256), .B(n45254), .Z(n45282) );
  XNOR U45273 ( .A(n45343), .B(n45261), .Z(n45254) );
  XOR U45274 ( .A(p_input[1528]), .B(p_input[2072]), .Z(n45261) );
  XOR U45275 ( .A(n45251), .B(n45260), .Z(n45343) );
  XOR U45276 ( .A(n45344), .B(n45257), .Z(n45260) );
  XOR U45277 ( .A(p_input[1526]), .B(p_input[2070]), .Z(n45257) );
  XOR U45278 ( .A(p_input[1527]), .B(n29410), .Z(n45344) );
  XOR U45279 ( .A(p_input[1522]), .B(p_input[2066]), .Z(n45251) );
  XNOR U45280 ( .A(n45266), .B(n45265), .Z(n45256) );
  XOR U45281 ( .A(n45345), .B(n45262), .Z(n45265) );
  XOR U45282 ( .A(p_input[1523]), .B(p_input[2067]), .Z(n45262) );
  XOR U45283 ( .A(p_input[1524]), .B(n29412), .Z(n45345) );
  XOR U45284 ( .A(p_input[1525]), .B(p_input[2069]), .Z(n45266) );
  XOR U45285 ( .A(n45281), .B(n45346), .Z(n45342) );
  IV U45286 ( .A(n45267), .Z(n45346) );
  XOR U45287 ( .A(p_input[1505]), .B(p_input[2049]), .Z(n45267) );
  XNOR U45288 ( .A(n45347), .B(n45289), .Z(n45281) );
  XNOR U45289 ( .A(n45277), .B(n45276), .Z(n45289) );
  XNOR U45290 ( .A(n45348), .B(n45273), .Z(n45276) );
  XNOR U45291 ( .A(p_input[1530]), .B(p_input[2074]), .Z(n45273) );
  XOR U45292 ( .A(p_input[1531]), .B(n29415), .Z(n45348) );
  XOR U45293 ( .A(p_input[1532]), .B(p_input[2076]), .Z(n45277) );
  XOR U45294 ( .A(n45287), .B(n45349), .Z(n45347) );
  IV U45295 ( .A(n45278), .Z(n45349) );
  XOR U45296 ( .A(p_input[1521]), .B(p_input[2065]), .Z(n45278) );
  XNOR U45297 ( .A(n45350), .B(n45294), .Z(n45287) );
  XNOR U45298 ( .A(p_input[1535]), .B(n29418), .Z(n45294) );
  XOR U45299 ( .A(n45284), .B(n45293), .Z(n45350) );
  XOR U45300 ( .A(n45351), .B(n45290), .Z(n45293) );
  XOR U45301 ( .A(p_input[1533]), .B(p_input[2077]), .Z(n45290) );
  XOR U45302 ( .A(p_input[1534]), .B(n29420), .Z(n45351) );
  XOR U45303 ( .A(p_input[1529]), .B(p_input[2073]), .Z(n45284) );
  XOR U45304 ( .A(n45306), .B(n45305), .Z(n45271) );
  XNOR U45305 ( .A(n45352), .B(n45313), .Z(n45305) );
  XNOR U45306 ( .A(n45301), .B(n45300), .Z(n45313) );
  XNOR U45307 ( .A(n45353), .B(n45297), .Z(n45300) );
  XNOR U45308 ( .A(p_input[1515]), .B(p_input[2059]), .Z(n45297) );
  XOR U45309 ( .A(p_input[1516]), .B(n28329), .Z(n45353) );
  XOR U45310 ( .A(p_input[1517]), .B(p_input[2061]), .Z(n45301) );
  XOR U45311 ( .A(n45311), .B(n45354), .Z(n45352) );
  IV U45312 ( .A(n45302), .Z(n45354) );
  XOR U45313 ( .A(p_input[1506]), .B(p_input[2050]), .Z(n45302) );
  XNOR U45314 ( .A(n45355), .B(n45318), .Z(n45311) );
  XNOR U45315 ( .A(p_input[1520]), .B(n28332), .Z(n45318) );
  XOR U45316 ( .A(n45308), .B(n45317), .Z(n45355) );
  XOR U45317 ( .A(n45356), .B(n45314), .Z(n45317) );
  XOR U45318 ( .A(p_input[1518]), .B(p_input[2062]), .Z(n45314) );
  XOR U45319 ( .A(p_input[1519]), .B(n28334), .Z(n45356) );
  XOR U45320 ( .A(p_input[1514]), .B(p_input[2058]), .Z(n45308) );
  XOR U45321 ( .A(n45325), .B(n45323), .Z(n45306) );
  XNOR U45322 ( .A(n45357), .B(n45330), .Z(n45323) );
  XOR U45323 ( .A(p_input[1513]), .B(p_input[2057]), .Z(n45330) );
  XOR U45324 ( .A(n45320), .B(n45329), .Z(n45357) );
  XOR U45325 ( .A(n45358), .B(n45326), .Z(n45329) );
  XOR U45326 ( .A(p_input[1511]), .B(p_input[2055]), .Z(n45326) );
  XOR U45327 ( .A(p_input[1512]), .B(n29427), .Z(n45358) );
  XOR U45328 ( .A(p_input[1507]), .B(p_input[2051]), .Z(n45320) );
  XNOR U45329 ( .A(n45335), .B(n45334), .Z(n45325) );
  XOR U45330 ( .A(n45359), .B(n45331), .Z(n45334) );
  XOR U45331 ( .A(p_input[1508]), .B(p_input[2052]), .Z(n45331) );
  XOR U45332 ( .A(p_input[1509]), .B(n29429), .Z(n45359) );
  XOR U45333 ( .A(p_input[1510]), .B(p_input[2054]), .Z(n45335) );
  XNOR U45334 ( .A(n45360), .B(n45361), .Z(n45136) );
  AND U45335 ( .A(n1028), .B(n45362), .Z(n45361) );
  XNOR U45336 ( .A(n45363), .B(n45364), .Z(n1028) );
  AND U45337 ( .A(n45365), .B(n45366), .Z(n45364) );
  XOR U45338 ( .A(n45150), .B(n45363), .Z(n45366) );
  XNOR U45339 ( .A(n45367), .B(n45363), .Z(n45365) );
  XOR U45340 ( .A(n45368), .B(n45369), .Z(n45363) );
  AND U45341 ( .A(n45370), .B(n45371), .Z(n45369) );
  XOR U45342 ( .A(n45165), .B(n45368), .Z(n45371) );
  XOR U45343 ( .A(n45368), .B(n45166), .Z(n45370) );
  XOR U45344 ( .A(n45372), .B(n45373), .Z(n45368) );
  AND U45345 ( .A(n45374), .B(n45375), .Z(n45373) );
  XOR U45346 ( .A(n45193), .B(n45372), .Z(n45375) );
  XOR U45347 ( .A(n45372), .B(n45194), .Z(n45374) );
  XOR U45348 ( .A(n45376), .B(n45377), .Z(n45372) );
  AND U45349 ( .A(n45378), .B(n45379), .Z(n45377) );
  XOR U45350 ( .A(n45242), .B(n45376), .Z(n45379) );
  XOR U45351 ( .A(n45376), .B(n45243), .Z(n45378) );
  XOR U45352 ( .A(n45380), .B(n45381), .Z(n45376) );
  AND U45353 ( .A(n45382), .B(n45383), .Z(n45381) );
  XOR U45354 ( .A(n45380), .B(n45339), .Z(n45383) );
  XNOR U45355 ( .A(n45384), .B(n45385), .Z(n45086) );
  AND U45356 ( .A(n1032), .B(n45386), .Z(n45385) );
  XNOR U45357 ( .A(n45387), .B(n45388), .Z(n1032) );
  AND U45358 ( .A(n45389), .B(n45390), .Z(n45388) );
  XOR U45359 ( .A(n45387), .B(n45096), .Z(n45390) );
  XNOR U45360 ( .A(n45387), .B(n45046), .Z(n45389) );
  XOR U45361 ( .A(n45391), .B(n45392), .Z(n45387) );
  AND U45362 ( .A(n45393), .B(n45394), .Z(n45392) );
  XNOR U45363 ( .A(n45106), .B(n45391), .Z(n45394) );
  XOR U45364 ( .A(n45391), .B(n45056), .Z(n45393) );
  XOR U45365 ( .A(n45395), .B(n45396), .Z(n45391) );
  AND U45366 ( .A(n45397), .B(n45398), .Z(n45396) );
  XNOR U45367 ( .A(n45116), .B(n45395), .Z(n45398) );
  XOR U45368 ( .A(n45395), .B(n45065), .Z(n45397) );
  XOR U45369 ( .A(n45399), .B(n45400), .Z(n45395) );
  AND U45370 ( .A(n45401), .B(n45402), .Z(n45400) );
  XOR U45371 ( .A(n45399), .B(n45073), .Z(n45401) );
  XOR U45372 ( .A(n45403), .B(n45404), .Z(n45037) );
  AND U45373 ( .A(n1036), .B(n45386), .Z(n45404) );
  XNOR U45374 ( .A(n45384), .B(n45403), .Z(n45386) );
  XNOR U45375 ( .A(n45405), .B(n45406), .Z(n1036) );
  AND U45376 ( .A(n45407), .B(n45408), .Z(n45406) );
  XNOR U45377 ( .A(n45409), .B(n45405), .Z(n45408) );
  IV U45378 ( .A(n45096), .Z(n45409) );
  XOR U45379 ( .A(n45367), .B(n45410), .Z(n45096) );
  AND U45380 ( .A(n1039), .B(n45411), .Z(n45410) );
  XOR U45381 ( .A(n45149), .B(n45146), .Z(n45411) );
  IV U45382 ( .A(n45367), .Z(n45149) );
  XNOR U45383 ( .A(n45046), .B(n45405), .Z(n45407) );
  XOR U45384 ( .A(n45412), .B(n45413), .Z(n45046) );
  AND U45385 ( .A(n1055), .B(n45414), .Z(n45413) );
  XOR U45386 ( .A(n45415), .B(n45416), .Z(n45405) );
  AND U45387 ( .A(n45417), .B(n45418), .Z(n45416) );
  XNOR U45388 ( .A(n45415), .B(n45106), .Z(n45418) );
  XOR U45389 ( .A(n45166), .B(n45419), .Z(n45106) );
  AND U45390 ( .A(n1039), .B(n45420), .Z(n45419) );
  XOR U45391 ( .A(n45162), .B(n45166), .Z(n45420) );
  XNOR U45392 ( .A(n45421), .B(n45415), .Z(n45417) );
  IV U45393 ( .A(n45056), .Z(n45421) );
  XOR U45394 ( .A(n45422), .B(n45423), .Z(n45056) );
  AND U45395 ( .A(n1055), .B(n45424), .Z(n45423) );
  XOR U45396 ( .A(n45425), .B(n45426), .Z(n45415) );
  AND U45397 ( .A(n45427), .B(n45428), .Z(n45426) );
  XNOR U45398 ( .A(n45425), .B(n45116), .Z(n45428) );
  XOR U45399 ( .A(n45194), .B(n45429), .Z(n45116) );
  AND U45400 ( .A(n1039), .B(n45430), .Z(n45429) );
  XOR U45401 ( .A(n45190), .B(n45194), .Z(n45430) );
  XOR U45402 ( .A(n45065), .B(n45425), .Z(n45427) );
  XOR U45403 ( .A(n45431), .B(n45432), .Z(n45065) );
  AND U45404 ( .A(n1055), .B(n45433), .Z(n45432) );
  XOR U45405 ( .A(n45399), .B(n45434), .Z(n45425) );
  AND U45406 ( .A(n45435), .B(n45402), .Z(n45434) );
  XNOR U45407 ( .A(n45126), .B(n45399), .Z(n45402) );
  XOR U45408 ( .A(n45243), .B(n45436), .Z(n45126) );
  AND U45409 ( .A(n1039), .B(n45437), .Z(n45436) );
  XOR U45410 ( .A(n45239), .B(n45243), .Z(n45437) );
  XNOR U45411 ( .A(n45438), .B(n45399), .Z(n45435) );
  IV U45412 ( .A(n45073), .Z(n45438) );
  XOR U45413 ( .A(n45439), .B(n45440), .Z(n45073) );
  AND U45414 ( .A(n1055), .B(n45441), .Z(n45440) );
  XOR U45415 ( .A(n45442), .B(n45443), .Z(n45399) );
  AND U45416 ( .A(n45444), .B(n45445), .Z(n45443) );
  XNOR U45417 ( .A(n45442), .B(n45134), .Z(n45445) );
  XOR U45418 ( .A(n45340), .B(n45446), .Z(n45134) );
  AND U45419 ( .A(n1039), .B(n45447), .Z(n45446) );
  XOR U45420 ( .A(n45336), .B(n45340), .Z(n45447) );
  XNOR U45421 ( .A(n45448), .B(n45442), .Z(n45444) );
  IV U45422 ( .A(n45083), .Z(n45448) );
  XOR U45423 ( .A(n45449), .B(n45450), .Z(n45083) );
  AND U45424 ( .A(n1055), .B(n45451), .Z(n45450) );
  AND U45425 ( .A(n45403), .B(n45384), .Z(n45442) );
  XNOR U45426 ( .A(n45452), .B(n45453), .Z(n45384) );
  AND U45427 ( .A(n1039), .B(n45362), .Z(n45453) );
  XNOR U45428 ( .A(n45360), .B(n45452), .Z(n45362) );
  XNOR U45429 ( .A(n45454), .B(n45455), .Z(n1039) );
  AND U45430 ( .A(n45456), .B(n45457), .Z(n45455) );
  XNOR U45431 ( .A(n45454), .B(n45146), .Z(n45457) );
  IV U45432 ( .A(n45150), .Z(n45146) );
  XOR U45433 ( .A(n45458), .B(n45459), .Z(n45150) );
  AND U45434 ( .A(n1043), .B(n45460), .Z(n45459) );
  XOR U45435 ( .A(n45461), .B(n45458), .Z(n45460) );
  XNOR U45436 ( .A(n45454), .B(n45367), .Z(n45456) );
  XOR U45437 ( .A(n45462), .B(n45463), .Z(n45367) );
  AND U45438 ( .A(n1051), .B(n45414), .Z(n45463) );
  XOR U45439 ( .A(n45412), .B(n45462), .Z(n45414) );
  XOR U45440 ( .A(n45464), .B(n45465), .Z(n45454) );
  AND U45441 ( .A(n45466), .B(n45467), .Z(n45465) );
  XNOR U45442 ( .A(n45464), .B(n45162), .Z(n45467) );
  IV U45443 ( .A(n45165), .Z(n45162) );
  XOR U45444 ( .A(n45468), .B(n45469), .Z(n45165) );
  AND U45445 ( .A(n1043), .B(n45470), .Z(n45469) );
  XOR U45446 ( .A(n45471), .B(n45468), .Z(n45470) );
  XOR U45447 ( .A(n45166), .B(n45464), .Z(n45466) );
  XOR U45448 ( .A(n45472), .B(n45473), .Z(n45166) );
  AND U45449 ( .A(n1051), .B(n45424), .Z(n45473) );
  XOR U45450 ( .A(n45472), .B(n45422), .Z(n45424) );
  XOR U45451 ( .A(n45474), .B(n45475), .Z(n45464) );
  AND U45452 ( .A(n45476), .B(n45477), .Z(n45475) );
  XNOR U45453 ( .A(n45474), .B(n45190), .Z(n45477) );
  IV U45454 ( .A(n45193), .Z(n45190) );
  XOR U45455 ( .A(n45478), .B(n45479), .Z(n45193) );
  AND U45456 ( .A(n1043), .B(n45480), .Z(n45479) );
  XNOR U45457 ( .A(n45481), .B(n45478), .Z(n45480) );
  XOR U45458 ( .A(n45194), .B(n45474), .Z(n45476) );
  XOR U45459 ( .A(n45482), .B(n45483), .Z(n45194) );
  AND U45460 ( .A(n1051), .B(n45433), .Z(n45483) );
  XOR U45461 ( .A(n45482), .B(n45431), .Z(n45433) );
  XOR U45462 ( .A(n45484), .B(n45485), .Z(n45474) );
  AND U45463 ( .A(n45486), .B(n45487), .Z(n45485) );
  XNOR U45464 ( .A(n45484), .B(n45239), .Z(n45487) );
  IV U45465 ( .A(n45242), .Z(n45239) );
  XOR U45466 ( .A(n45488), .B(n45489), .Z(n45242) );
  AND U45467 ( .A(n1043), .B(n45490), .Z(n45489) );
  XOR U45468 ( .A(n45491), .B(n45488), .Z(n45490) );
  XOR U45469 ( .A(n45243), .B(n45484), .Z(n45486) );
  XOR U45470 ( .A(n45492), .B(n45493), .Z(n45243) );
  AND U45471 ( .A(n1051), .B(n45441), .Z(n45493) );
  XOR U45472 ( .A(n45492), .B(n45439), .Z(n45441) );
  XOR U45473 ( .A(n45380), .B(n45494), .Z(n45484) );
  AND U45474 ( .A(n45382), .B(n45495), .Z(n45494) );
  XNOR U45475 ( .A(n45380), .B(n45336), .Z(n45495) );
  IV U45476 ( .A(n45339), .Z(n45336) );
  XOR U45477 ( .A(n45496), .B(n45497), .Z(n45339) );
  AND U45478 ( .A(n1043), .B(n45498), .Z(n45497) );
  XNOR U45479 ( .A(n45499), .B(n45496), .Z(n45498) );
  XOR U45480 ( .A(n45340), .B(n45380), .Z(n45382) );
  XOR U45481 ( .A(n45500), .B(n45501), .Z(n45340) );
  AND U45482 ( .A(n1051), .B(n45451), .Z(n45501) );
  XOR U45483 ( .A(n45500), .B(n45449), .Z(n45451) );
  AND U45484 ( .A(n45452), .B(n45360), .Z(n45380) );
  XNOR U45485 ( .A(n45502), .B(n45503), .Z(n45360) );
  AND U45486 ( .A(n1043), .B(n45504), .Z(n45503) );
  XNOR U45487 ( .A(n45505), .B(n45502), .Z(n45504) );
  XNOR U45488 ( .A(n45506), .B(n45507), .Z(n1043) );
  AND U45489 ( .A(n45508), .B(n45509), .Z(n45507) );
  XOR U45490 ( .A(n45461), .B(n45506), .Z(n45509) );
  AND U45491 ( .A(n45510), .B(n45511), .Z(n45461) );
  XNOR U45492 ( .A(n45458), .B(n45506), .Z(n45508) );
  XNOR U45493 ( .A(n45512), .B(n45513), .Z(n45458) );
  AND U45494 ( .A(n1047), .B(n45514), .Z(n45513) );
  XNOR U45495 ( .A(n45515), .B(n45516), .Z(n45514) );
  XOR U45496 ( .A(n45517), .B(n45518), .Z(n45506) );
  AND U45497 ( .A(n45519), .B(n45520), .Z(n45518) );
  XNOR U45498 ( .A(n45517), .B(n45510), .Z(n45520) );
  IV U45499 ( .A(n45471), .Z(n45510) );
  XOR U45500 ( .A(n45521), .B(n45522), .Z(n45471) );
  XOR U45501 ( .A(n45523), .B(n45511), .Z(n45522) );
  AND U45502 ( .A(n45481), .B(n45524), .Z(n45511) );
  AND U45503 ( .A(n45525), .B(n45526), .Z(n45523) );
  XOR U45504 ( .A(n45527), .B(n45521), .Z(n45525) );
  XNOR U45505 ( .A(n45468), .B(n45517), .Z(n45519) );
  XNOR U45506 ( .A(n45528), .B(n45529), .Z(n45468) );
  AND U45507 ( .A(n1047), .B(n45530), .Z(n45529) );
  XNOR U45508 ( .A(n45531), .B(n45532), .Z(n45530) );
  XOR U45509 ( .A(n45533), .B(n45534), .Z(n45517) );
  AND U45510 ( .A(n45535), .B(n45536), .Z(n45534) );
  XNOR U45511 ( .A(n45533), .B(n45481), .Z(n45536) );
  XOR U45512 ( .A(n45537), .B(n45526), .Z(n45481) );
  XNOR U45513 ( .A(n45538), .B(n45521), .Z(n45526) );
  XOR U45514 ( .A(n45539), .B(n45540), .Z(n45521) );
  AND U45515 ( .A(n45541), .B(n45542), .Z(n45540) );
  XOR U45516 ( .A(n45543), .B(n45539), .Z(n45541) );
  XNOR U45517 ( .A(n45544), .B(n45545), .Z(n45538) );
  AND U45518 ( .A(n45546), .B(n45547), .Z(n45545) );
  XOR U45519 ( .A(n45544), .B(n45548), .Z(n45546) );
  XNOR U45520 ( .A(n45527), .B(n45524), .Z(n45537) );
  AND U45521 ( .A(n45549), .B(n45550), .Z(n45524) );
  XOR U45522 ( .A(n45551), .B(n45552), .Z(n45527) );
  AND U45523 ( .A(n45553), .B(n45554), .Z(n45552) );
  XOR U45524 ( .A(n45551), .B(n45555), .Z(n45553) );
  XNOR U45525 ( .A(n45478), .B(n45533), .Z(n45535) );
  XNOR U45526 ( .A(n45556), .B(n45557), .Z(n45478) );
  AND U45527 ( .A(n1047), .B(n45558), .Z(n45557) );
  XNOR U45528 ( .A(n45559), .B(n45560), .Z(n45558) );
  XOR U45529 ( .A(n45561), .B(n45562), .Z(n45533) );
  AND U45530 ( .A(n45563), .B(n45564), .Z(n45562) );
  XNOR U45531 ( .A(n45561), .B(n45549), .Z(n45564) );
  IV U45532 ( .A(n45491), .Z(n45549) );
  XNOR U45533 ( .A(n45565), .B(n45542), .Z(n45491) );
  XNOR U45534 ( .A(n45566), .B(n45548), .Z(n45542) );
  XOR U45535 ( .A(n45567), .B(n45568), .Z(n45548) );
  AND U45536 ( .A(n45569), .B(n45570), .Z(n45568) );
  XOR U45537 ( .A(n45567), .B(n45571), .Z(n45569) );
  XNOR U45538 ( .A(n45547), .B(n45539), .Z(n45566) );
  XOR U45539 ( .A(n45572), .B(n45573), .Z(n45539) );
  AND U45540 ( .A(n45574), .B(n45575), .Z(n45573) );
  XNOR U45541 ( .A(n45576), .B(n45572), .Z(n45574) );
  XNOR U45542 ( .A(n45577), .B(n45544), .Z(n45547) );
  XOR U45543 ( .A(n45578), .B(n45579), .Z(n45544) );
  AND U45544 ( .A(n45580), .B(n45581), .Z(n45579) );
  XOR U45545 ( .A(n45578), .B(n45582), .Z(n45580) );
  XNOR U45546 ( .A(n45583), .B(n45584), .Z(n45577) );
  AND U45547 ( .A(n45585), .B(n45586), .Z(n45584) );
  XNOR U45548 ( .A(n45583), .B(n45587), .Z(n45585) );
  XNOR U45549 ( .A(n45543), .B(n45550), .Z(n45565) );
  AND U45550 ( .A(n45499), .B(n45588), .Z(n45550) );
  XOR U45551 ( .A(n45555), .B(n45554), .Z(n45543) );
  XNOR U45552 ( .A(n45589), .B(n45551), .Z(n45554) );
  XOR U45553 ( .A(n45590), .B(n45591), .Z(n45551) );
  AND U45554 ( .A(n45592), .B(n45593), .Z(n45591) );
  XOR U45555 ( .A(n45590), .B(n45594), .Z(n45592) );
  XNOR U45556 ( .A(n45595), .B(n45596), .Z(n45589) );
  AND U45557 ( .A(n45597), .B(n45598), .Z(n45596) );
  XOR U45558 ( .A(n45595), .B(n45599), .Z(n45597) );
  XOR U45559 ( .A(n45600), .B(n45601), .Z(n45555) );
  AND U45560 ( .A(n45602), .B(n45603), .Z(n45601) );
  XOR U45561 ( .A(n45600), .B(n45604), .Z(n45602) );
  XNOR U45562 ( .A(n45488), .B(n45561), .Z(n45563) );
  XNOR U45563 ( .A(n45605), .B(n45606), .Z(n45488) );
  AND U45564 ( .A(n1047), .B(n45607), .Z(n45606) );
  XNOR U45565 ( .A(n45608), .B(n45609), .Z(n45607) );
  XOR U45566 ( .A(n45610), .B(n45611), .Z(n45561) );
  AND U45567 ( .A(n45612), .B(n45613), .Z(n45611) );
  XNOR U45568 ( .A(n45610), .B(n45499), .Z(n45613) );
  XOR U45569 ( .A(n45614), .B(n45575), .Z(n45499) );
  XNOR U45570 ( .A(n45615), .B(n45582), .Z(n45575) );
  XOR U45571 ( .A(n45571), .B(n45570), .Z(n45582) );
  XNOR U45572 ( .A(n45616), .B(n45567), .Z(n45570) );
  XOR U45573 ( .A(n45617), .B(n45618), .Z(n45567) );
  AND U45574 ( .A(n45619), .B(n45620), .Z(n45618) );
  XNOR U45575 ( .A(n45621), .B(n45622), .Z(n45619) );
  IV U45576 ( .A(n45617), .Z(n45621) );
  XNOR U45577 ( .A(n45623), .B(n45624), .Z(n45616) );
  NOR U45578 ( .A(n45625), .B(n45626), .Z(n45624) );
  XNOR U45579 ( .A(n45623), .B(n45627), .Z(n45625) );
  XOR U45580 ( .A(n45628), .B(n45629), .Z(n45571) );
  NOR U45581 ( .A(n45630), .B(n45631), .Z(n45629) );
  XNOR U45582 ( .A(n45628), .B(n45632), .Z(n45630) );
  XNOR U45583 ( .A(n45581), .B(n45572), .Z(n45615) );
  XOR U45584 ( .A(n45633), .B(n45634), .Z(n45572) );
  AND U45585 ( .A(n45635), .B(n45636), .Z(n45634) );
  XOR U45586 ( .A(n45633), .B(n45637), .Z(n45635) );
  XOR U45587 ( .A(n45638), .B(n45587), .Z(n45581) );
  XOR U45588 ( .A(n45639), .B(n45640), .Z(n45587) );
  NOR U45589 ( .A(n45641), .B(n45642), .Z(n45640) );
  XOR U45590 ( .A(n45639), .B(n45643), .Z(n45641) );
  XNOR U45591 ( .A(n45586), .B(n45578), .Z(n45638) );
  XOR U45592 ( .A(n45644), .B(n45645), .Z(n45578) );
  AND U45593 ( .A(n45646), .B(n45647), .Z(n45645) );
  XOR U45594 ( .A(n45644), .B(n45648), .Z(n45646) );
  XNOR U45595 ( .A(n45649), .B(n45583), .Z(n45586) );
  XOR U45596 ( .A(n45650), .B(n45651), .Z(n45583) );
  AND U45597 ( .A(n45652), .B(n45653), .Z(n45651) );
  XNOR U45598 ( .A(n45654), .B(n45655), .Z(n45652) );
  IV U45599 ( .A(n45650), .Z(n45654) );
  XNOR U45600 ( .A(n45656), .B(n45657), .Z(n45649) );
  NOR U45601 ( .A(n45658), .B(n45659), .Z(n45657) );
  XNOR U45602 ( .A(n45656), .B(n45660), .Z(n45658) );
  XOR U45603 ( .A(n45576), .B(n45588), .Z(n45614) );
  NOR U45604 ( .A(n45505), .B(n45661), .Z(n45588) );
  XNOR U45605 ( .A(n45594), .B(n45593), .Z(n45576) );
  XNOR U45606 ( .A(n45662), .B(n45599), .Z(n45593) );
  XNOR U45607 ( .A(n45663), .B(n45664), .Z(n45599) );
  NOR U45608 ( .A(n45665), .B(n45666), .Z(n45664) );
  XOR U45609 ( .A(n45663), .B(n45667), .Z(n45665) );
  XNOR U45610 ( .A(n45598), .B(n45590), .Z(n45662) );
  XOR U45611 ( .A(n45668), .B(n45669), .Z(n45590) );
  AND U45612 ( .A(n45670), .B(n45671), .Z(n45669) );
  XOR U45613 ( .A(n45668), .B(n45672), .Z(n45670) );
  XNOR U45614 ( .A(n45673), .B(n45595), .Z(n45598) );
  XOR U45615 ( .A(n45674), .B(n45675), .Z(n45595) );
  AND U45616 ( .A(n45676), .B(n45677), .Z(n45675) );
  XNOR U45617 ( .A(n45678), .B(n45679), .Z(n45676) );
  IV U45618 ( .A(n45674), .Z(n45678) );
  XNOR U45619 ( .A(n45680), .B(n45681), .Z(n45673) );
  NOR U45620 ( .A(n45682), .B(n45683), .Z(n45681) );
  XNOR U45621 ( .A(n45680), .B(n45684), .Z(n45682) );
  XOR U45622 ( .A(n45604), .B(n45603), .Z(n45594) );
  XNOR U45623 ( .A(n45685), .B(n45600), .Z(n45603) );
  XOR U45624 ( .A(n45686), .B(n45687), .Z(n45600) );
  AND U45625 ( .A(n45688), .B(n45689), .Z(n45687) );
  XNOR U45626 ( .A(n45690), .B(n45691), .Z(n45688) );
  IV U45627 ( .A(n45686), .Z(n45690) );
  XNOR U45628 ( .A(n45692), .B(n45693), .Z(n45685) );
  NOR U45629 ( .A(n45694), .B(n45695), .Z(n45693) );
  XNOR U45630 ( .A(n45692), .B(n45696), .Z(n45694) );
  XOR U45631 ( .A(n45697), .B(n45698), .Z(n45604) );
  NOR U45632 ( .A(n45699), .B(n45700), .Z(n45698) );
  XNOR U45633 ( .A(n45697), .B(n45701), .Z(n45699) );
  XNOR U45634 ( .A(n45496), .B(n45610), .Z(n45612) );
  XNOR U45635 ( .A(n45702), .B(n45703), .Z(n45496) );
  AND U45636 ( .A(n1047), .B(n45704), .Z(n45703) );
  XNOR U45637 ( .A(n45705), .B(n45706), .Z(n45704) );
  AND U45638 ( .A(n45502), .B(n45505), .Z(n45610) );
  XOR U45639 ( .A(n45707), .B(n45661), .Z(n45505) );
  XNOR U45640 ( .A(p_input[1536]), .B(p_input[2048]), .Z(n45661) );
  XNOR U45641 ( .A(n45637), .B(n45636), .Z(n45707) );
  XNOR U45642 ( .A(n45708), .B(n45648), .Z(n45636) );
  XOR U45643 ( .A(n45622), .B(n45620), .Z(n45648) );
  XNOR U45644 ( .A(n45709), .B(n45627), .Z(n45620) );
  XOR U45645 ( .A(p_input[1560]), .B(p_input[2072]), .Z(n45627) );
  XOR U45646 ( .A(n45617), .B(n45626), .Z(n45709) );
  XOR U45647 ( .A(n45710), .B(n45623), .Z(n45626) );
  XOR U45648 ( .A(p_input[1558]), .B(p_input[2070]), .Z(n45623) );
  XOR U45649 ( .A(p_input[1559]), .B(n29410), .Z(n45710) );
  XOR U45650 ( .A(p_input[1554]), .B(p_input[2066]), .Z(n45617) );
  XNOR U45651 ( .A(n45632), .B(n45631), .Z(n45622) );
  XOR U45652 ( .A(n45711), .B(n45628), .Z(n45631) );
  XOR U45653 ( .A(p_input[1555]), .B(p_input[2067]), .Z(n45628) );
  XOR U45654 ( .A(p_input[1556]), .B(n29412), .Z(n45711) );
  XOR U45655 ( .A(p_input[1557]), .B(p_input[2069]), .Z(n45632) );
  XOR U45656 ( .A(n45647), .B(n45712), .Z(n45708) );
  IV U45657 ( .A(n45633), .Z(n45712) );
  XOR U45658 ( .A(p_input[1537]), .B(p_input[2049]), .Z(n45633) );
  XNOR U45659 ( .A(n45713), .B(n45655), .Z(n45647) );
  XNOR U45660 ( .A(n45643), .B(n45642), .Z(n45655) );
  XNOR U45661 ( .A(n45714), .B(n45639), .Z(n45642) );
  XNOR U45662 ( .A(p_input[1562]), .B(p_input[2074]), .Z(n45639) );
  XOR U45663 ( .A(p_input[1563]), .B(n29415), .Z(n45714) );
  XOR U45664 ( .A(p_input[1564]), .B(p_input[2076]), .Z(n45643) );
  XOR U45665 ( .A(n45653), .B(n45715), .Z(n45713) );
  IV U45666 ( .A(n45644), .Z(n45715) );
  XOR U45667 ( .A(p_input[1553]), .B(p_input[2065]), .Z(n45644) );
  XNOR U45668 ( .A(n45716), .B(n45660), .Z(n45653) );
  XNOR U45669 ( .A(p_input[1567]), .B(n29418), .Z(n45660) );
  XOR U45670 ( .A(n45650), .B(n45659), .Z(n45716) );
  XOR U45671 ( .A(n45717), .B(n45656), .Z(n45659) );
  XOR U45672 ( .A(p_input[1565]), .B(p_input[2077]), .Z(n45656) );
  XOR U45673 ( .A(p_input[1566]), .B(n29420), .Z(n45717) );
  XOR U45674 ( .A(p_input[1561]), .B(p_input[2073]), .Z(n45650) );
  XOR U45675 ( .A(n45672), .B(n45671), .Z(n45637) );
  XNOR U45676 ( .A(n45718), .B(n45679), .Z(n45671) );
  XNOR U45677 ( .A(n45667), .B(n45666), .Z(n45679) );
  XNOR U45678 ( .A(n45719), .B(n45663), .Z(n45666) );
  XNOR U45679 ( .A(p_input[1547]), .B(p_input[2059]), .Z(n45663) );
  XOR U45680 ( .A(p_input[1548]), .B(n28329), .Z(n45719) );
  XOR U45681 ( .A(p_input[1549]), .B(p_input[2061]), .Z(n45667) );
  XOR U45682 ( .A(n45677), .B(n45720), .Z(n45718) );
  IV U45683 ( .A(n45668), .Z(n45720) );
  XOR U45684 ( .A(p_input[1538]), .B(p_input[2050]), .Z(n45668) );
  XNOR U45685 ( .A(n45721), .B(n45684), .Z(n45677) );
  XNOR U45686 ( .A(p_input[1552]), .B(n28332), .Z(n45684) );
  XOR U45687 ( .A(n45674), .B(n45683), .Z(n45721) );
  XOR U45688 ( .A(n45722), .B(n45680), .Z(n45683) );
  XOR U45689 ( .A(p_input[1550]), .B(p_input[2062]), .Z(n45680) );
  XOR U45690 ( .A(p_input[1551]), .B(n28334), .Z(n45722) );
  XOR U45691 ( .A(p_input[1546]), .B(p_input[2058]), .Z(n45674) );
  XOR U45692 ( .A(n45691), .B(n45689), .Z(n45672) );
  XNOR U45693 ( .A(n45723), .B(n45696), .Z(n45689) );
  XOR U45694 ( .A(p_input[1545]), .B(p_input[2057]), .Z(n45696) );
  XOR U45695 ( .A(n45686), .B(n45695), .Z(n45723) );
  XOR U45696 ( .A(n45724), .B(n45692), .Z(n45695) );
  XOR U45697 ( .A(p_input[1543]), .B(p_input[2055]), .Z(n45692) );
  XOR U45698 ( .A(p_input[1544]), .B(n29427), .Z(n45724) );
  XOR U45699 ( .A(p_input[1539]), .B(p_input[2051]), .Z(n45686) );
  XNOR U45700 ( .A(n45701), .B(n45700), .Z(n45691) );
  XOR U45701 ( .A(n45725), .B(n45697), .Z(n45700) );
  XOR U45702 ( .A(p_input[1540]), .B(p_input[2052]), .Z(n45697) );
  XOR U45703 ( .A(p_input[1541]), .B(n29429), .Z(n45725) );
  XOR U45704 ( .A(p_input[1542]), .B(p_input[2054]), .Z(n45701) );
  XNOR U45705 ( .A(n45726), .B(n45727), .Z(n45502) );
  AND U45706 ( .A(n1047), .B(n45728), .Z(n45727) );
  XNOR U45707 ( .A(n45729), .B(n45730), .Z(n1047) );
  AND U45708 ( .A(n45731), .B(n45732), .Z(n45730) );
  XOR U45709 ( .A(n45516), .B(n45729), .Z(n45732) );
  XNOR U45710 ( .A(n45733), .B(n45729), .Z(n45731) );
  XOR U45711 ( .A(n45734), .B(n45735), .Z(n45729) );
  AND U45712 ( .A(n45736), .B(n45737), .Z(n45735) );
  XOR U45713 ( .A(n45531), .B(n45734), .Z(n45737) );
  XOR U45714 ( .A(n45734), .B(n45532), .Z(n45736) );
  XOR U45715 ( .A(n45738), .B(n45739), .Z(n45734) );
  AND U45716 ( .A(n45740), .B(n45741), .Z(n45739) );
  XOR U45717 ( .A(n45559), .B(n45738), .Z(n45741) );
  XOR U45718 ( .A(n45738), .B(n45560), .Z(n45740) );
  XOR U45719 ( .A(n45742), .B(n45743), .Z(n45738) );
  AND U45720 ( .A(n45744), .B(n45745), .Z(n45743) );
  XOR U45721 ( .A(n45608), .B(n45742), .Z(n45745) );
  XOR U45722 ( .A(n45742), .B(n45609), .Z(n45744) );
  XOR U45723 ( .A(n45746), .B(n45747), .Z(n45742) );
  AND U45724 ( .A(n45748), .B(n45749), .Z(n45747) );
  XOR U45725 ( .A(n45746), .B(n45705), .Z(n45749) );
  XNOR U45726 ( .A(n45750), .B(n45751), .Z(n45452) );
  AND U45727 ( .A(n1051), .B(n45752), .Z(n45751) );
  XNOR U45728 ( .A(n45753), .B(n45754), .Z(n1051) );
  AND U45729 ( .A(n45755), .B(n45756), .Z(n45754) );
  XOR U45730 ( .A(n45753), .B(n45462), .Z(n45756) );
  XNOR U45731 ( .A(n45753), .B(n45412), .Z(n45755) );
  XOR U45732 ( .A(n45757), .B(n45758), .Z(n45753) );
  AND U45733 ( .A(n45759), .B(n45760), .Z(n45758) );
  XNOR U45734 ( .A(n45472), .B(n45757), .Z(n45760) );
  XOR U45735 ( .A(n45757), .B(n45422), .Z(n45759) );
  XOR U45736 ( .A(n45761), .B(n45762), .Z(n45757) );
  AND U45737 ( .A(n45763), .B(n45764), .Z(n45762) );
  XNOR U45738 ( .A(n45482), .B(n45761), .Z(n45764) );
  XOR U45739 ( .A(n45761), .B(n45431), .Z(n45763) );
  XOR U45740 ( .A(n45765), .B(n45766), .Z(n45761) );
  AND U45741 ( .A(n45767), .B(n45768), .Z(n45766) );
  XOR U45742 ( .A(n45765), .B(n45439), .Z(n45767) );
  XOR U45743 ( .A(n45769), .B(n45770), .Z(n45403) );
  AND U45744 ( .A(n1055), .B(n45752), .Z(n45770) );
  XNOR U45745 ( .A(n45750), .B(n45769), .Z(n45752) );
  XNOR U45746 ( .A(n45771), .B(n45772), .Z(n1055) );
  AND U45747 ( .A(n45773), .B(n45774), .Z(n45772) );
  XNOR U45748 ( .A(n45775), .B(n45771), .Z(n45774) );
  IV U45749 ( .A(n45462), .Z(n45775) );
  XOR U45750 ( .A(n45733), .B(n45776), .Z(n45462) );
  AND U45751 ( .A(n1058), .B(n45777), .Z(n45776) );
  XOR U45752 ( .A(n45515), .B(n45512), .Z(n45777) );
  IV U45753 ( .A(n45733), .Z(n45515) );
  XNOR U45754 ( .A(n45412), .B(n45771), .Z(n45773) );
  XOR U45755 ( .A(n45778), .B(n45779), .Z(n45412) );
  AND U45756 ( .A(n1074), .B(n45780), .Z(n45779) );
  XOR U45757 ( .A(n45781), .B(n45782), .Z(n45771) );
  AND U45758 ( .A(n45783), .B(n45784), .Z(n45782) );
  XNOR U45759 ( .A(n45781), .B(n45472), .Z(n45784) );
  XOR U45760 ( .A(n45532), .B(n45785), .Z(n45472) );
  AND U45761 ( .A(n1058), .B(n45786), .Z(n45785) );
  XOR U45762 ( .A(n45528), .B(n45532), .Z(n45786) );
  XNOR U45763 ( .A(n45787), .B(n45781), .Z(n45783) );
  IV U45764 ( .A(n45422), .Z(n45787) );
  XOR U45765 ( .A(n45788), .B(n45789), .Z(n45422) );
  AND U45766 ( .A(n1074), .B(n45790), .Z(n45789) );
  XOR U45767 ( .A(n45791), .B(n45792), .Z(n45781) );
  AND U45768 ( .A(n45793), .B(n45794), .Z(n45792) );
  XNOR U45769 ( .A(n45791), .B(n45482), .Z(n45794) );
  XOR U45770 ( .A(n45560), .B(n45795), .Z(n45482) );
  AND U45771 ( .A(n1058), .B(n45796), .Z(n45795) );
  XOR U45772 ( .A(n45556), .B(n45560), .Z(n45796) );
  XOR U45773 ( .A(n45431), .B(n45791), .Z(n45793) );
  XOR U45774 ( .A(n45797), .B(n45798), .Z(n45431) );
  AND U45775 ( .A(n1074), .B(n45799), .Z(n45798) );
  XOR U45776 ( .A(n45765), .B(n45800), .Z(n45791) );
  AND U45777 ( .A(n45801), .B(n45768), .Z(n45800) );
  XNOR U45778 ( .A(n45492), .B(n45765), .Z(n45768) );
  XOR U45779 ( .A(n45609), .B(n45802), .Z(n45492) );
  AND U45780 ( .A(n1058), .B(n45803), .Z(n45802) );
  XOR U45781 ( .A(n45605), .B(n45609), .Z(n45803) );
  XNOR U45782 ( .A(n45804), .B(n45765), .Z(n45801) );
  IV U45783 ( .A(n45439), .Z(n45804) );
  XOR U45784 ( .A(n45805), .B(n45806), .Z(n45439) );
  AND U45785 ( .A(n1074), .B(n45807), .Z(n45806) );
  XOR U45786 ( .A(n45808), .B(n45809), .Z(n45765) );
  AND U45787 ( .A(n45810), .B(n45811), .Z(n45809) );
  XNOR U45788 ( .A(n45808), .B(n45500), .Z(n45811) );
  XOR U45789 ( .A(n45706), .B(n45812), .Z(n45500) );
  AND U45790 ( .A(n1058), .B(n45813), .Z(n45812) );
  XOR U45791 ( .A(n45702), .B(n45706), .Z(n45813) );
  XNOR U45792 ( .A(n45814), .B(n45808), .Z(n45810) );
  IV U45793 ( .A(n45449), .Z(n45814) );
  XOR U45794 ( .A(n45815), .B(n45816), .Z(n45449) );
  AND U45795 ( .A(n1074), .B(n45817), .Z(n45816) );
  AND U45796 ( .A(n45769), .B(n45750), .Z(n45808) );
  XNOR U45797 ( .A(n45818), .B(n45819), .Z(n45750) );
  AND U45798 ( .A(n1058), .B(n45728), .Z(n45819) );
  XNOR U45799 ( .A(n45726), .B(n45818), .Z(n45728) );
  XNOR U45800 ( .A(n45820), .B(n45821), .Z(n1058) );
  AND U45801 ( .A(n45822), .B(n45823), .Z(n45821) );
  XNOR U45802 ( .A(n45820), .B(n45512), .Z(n45823) );
  IV U45803 ( .A(n45516), .Z(n45512) );
  XOR U45804 ( .A(n45824), .B(n45825), .Z(n45516) );
  AND U45805 ( .A(n1062), .B(n45826), .Z(n45825) );
  XOR U45806 ( .A(n45827), .B(n45824), .Z(n45826) );
  XNOR U45807 ( .A(n45820), .B(n45733), .Z(n45822) );
  XOR U45808 ( .A(n45828), .B(n45829), .Z(n45733) );
  AND U45809 ( .A(n1070), .B(n45780), .Z(n45829) );
  XOR U45810 ( .A(n45778), .B(n45828), .Z(n45780) );
  XOR U45811 ( .A(n45830), .B(n45831), .Z(n45820) );
  AND U45812 ( .A(n45832), .B(n45833), .Z(n45831) );
  XNOR U45813 ( .A(n45830), .B(n45528), .Z(n45833) );
  IV U45814 ( .A(n45531), .Z(n45528) );
  XOR U45815 ( .A(n45834), .B(n45835), .Z(n45531) );
  AND U45816 ( .A(n1062), .B(n45836), .Z(n45835) );
  XOR U45817 ( .A(n45837), .B(n45834), .Z(n45836) );
  XOR U45818 ( .A(n45532), .B(n45830), .Z(n45832) );
  XOR U45819 ( .A(n45838), .B(n45839), .Z(n45532) );
  AND U45820 ( .A(n1070), .B(n45790), .Z(n45839) );
  XOR U45821 ( .A(n45838), .B(n45788), .Z(n45790) );
  XOR U45822 ( .A(n45840), .B(n45841), .Z(n45830) );
  AND U45823 ( .A(n45842), .B(n45843), .Z(n45841) );
  XNOR U45824 ( .A(n45840), .B(n45556), .Z(n45843) );
  IV U45825 ( .A(n45559), .Z(n45556) );
  XOR U45826 ( .A(n45844), .B(n45845), .Z(n45559) );
  AND U45827 ( .A(n1062), .B(n45846), .Z(n45845) );
  XNOR U45828 ( .A(n45847), .B(n45844), .Z(n45846) );
  XOR U45829 ( .A(n45560), .B(n45840), .Z(n45842) );
  XOR U45830 ( .A(n45848), .B(n45849), .Z(n45560) );
  AND U45831 ( .A(n1070), .B(n45799), .Z(n45849) );
  XOR U45832 ( .A(n45848), .B(n45797), .Z(n45799) );
  XOR U45833 ( .A(n45850), .B(n45851), .Z(n45840) );
  AND U45834 ( .A(n45852), .B(n45853), .Z(n45851) );
  XNOR U45835 ( .A(n45850), .B(n45605), .Z(n45853) );
  IV U45836 ( .A(n45608), .Z(n45605) );
  XOR U45837 ( .A(n45854), .B(n45855), .Z(n45608) );
  AND U45838 ( .A(n1062), .B(n45856), .Z(n45855) );
  XOR U45839 ( .A(n45857), .B(n45854), .Z(n45856) );
  XOR U45840 ( .A(n45609), .B(n45850), .Z(n45852) );
  XOR U45841 ( .A(n45858), .B(n45859), .Z(n45609) );
  AND U45842 ( .A(n1070), .B(n45807), .Z(n45859) );
  XOR U45843 ( .A(n45858), .B(n45805), .Z(n45807) );
  XOR U45844 ( .A(n45746), .B(n45860), .Z(n45850) );
  AND U45845 ( .A(n45748), .B(n45861), .Z(n45860) );
  XNOR U45846 ( .A(n45746), .B(n45702), .Z(n45861) );
  IV U45847 ( .A(n45705), .Z(n45702) );
  XOR U45848 ( .A(n45862), .B(n45863), .Z(n45705) );
  AND U45849 ( .A(n1062), .B(n45864), .Z(n45863) );
  XNOR U45850 ( .A(n45865), .B(n45862), .Z(n45864) );
  XOR U45851 ( .A(n45706), .B(n45746), .Z(n45748) );
  XOR U45852 ( .A(n45866), .B(n45867), .Z(n45706) );
  AND U45853 ( .A(n1070), .B(n45817), .Z(n45867) );
  XOR U45854 ( .A(n45866), .B(n45815), .Z(n45817) );
  AND U45855 ( .A(n45818), .B(n45726), .Z(n45746) );
  XNOR U45856 ( .A(n45868), .B(n45869), .Z(n45726) );
  AND U45857 ( .A(n1062), .B(n45870), .Z(n45869) );
  XNOR U45858 ( .A(n45871), .B(n45868), .Z(n45870) );
  XNOR U45859 ( .A(n45872), .B(n45873), .Z(n1062) );
  AND U45860 ( .A(n45874), .B(n45875), .Z(n45873) );
  XOR U45861 ( .A(n45827), .B(n45872), .Z(n45875) );
  AND U45862 ( .A(n45876), .B(n45877), .Z(n45827) );
  XNOR U45863 ( .A(n45824), .B(n45872), .Z(n45874) );
  XNOR U45864 ( .A(n45878), .B(n45879), .Z(n45824) );
  AND U45865 ( .A(n1066), .B(n45880), .Z(n45879) );
  XNOR U45866 ( .A(n45881), .B(n45882), .Z(n45880) );
  XOR U45867 ( .A(n45883), .B(n45884), .Z(n45872) );
  AND U45868 ( .A(n45885), .B(n45886), .Z(n45884) );
  XNOR U45869 ( .A(n45883), .B(n45876), .Z(n45886) );
  IV U45870 ( .A(n45837), .Z(n45876) );
  XOR U45871 ( .A(n45887), .B(n45888), .Z(n45837) );
  XOR U45872 ( .A(n45889), .B(n45877), .Z(n45888) );
  AND U45873 ( .A(n45847), .B(n45890), .Z(n45877) );
  AND U45874 ( .A(n45891), .B(n45892), .Z(n45889) );
  XOR U45875 ( .A(n45893), .B(n45887), .Z(n45891) );
  XNOR U45876 ( .A(n45834), .B(n45883), .Z(n45885) );
  XNOR U45877 ( .A(n45894), .B(n45895), .Z(n45834) );
  AND U45878 ( .A(n1066), .B(n45896), .Z(n45895) );
  XNOR U45879 ( .A(n45897), .B(n45898), .Z(n45896) );
  XOR U45880 ( .A(n45899), .B(n45900), .Z(n45883) );
  AND U45881 ( .A(n45901), .B(n45902), .Z(n45900) );
  XNOR U45882 ( .A(n45899), .B(n45847), .Z(n45902) );
  XOR U45883 ( .A(n45903), .B(n45892), .Z(n45847) );
  XNOR U45884 ( .A(n45904), .B(n45887), .Z(n45892) );
  XOR U45885 ( .A(n45905), .B(n45906), .Z(n45887) );
  AND U45886 ( .A(n45907), .B(n45908), .Z(n45906) );
  XOR U45887 ( .A(n45909), .B(n45905), .Z(n45907) );
  XNOR U45888 ( .A(n45910), .B(n45911), .Z(n45904) );
  AND U45889 ( .A(n45912), .B(n45913), .Z(n45911) );
  XOR U45890 ( .A(n45910), .B(n45914), .Z(n45912) );
  XNOR U45891 ( .A(n45893), .B(n45890), .Z(n45903) );
  AND U45892 ( .A(n45915), .B(n45916), .Z(n45890) );
  XOR U45893 ( .A(n45917), .B(n45918), .Z(n45893) );
  AND U45894 ( .A(n45919), .B(n45920), .Z(n45918) );
  XOR U45895 ( .A(n45917), .B(n45921), .Z(n45919) );
  XNOR U45896 ( .A(n45844), .B(n45899), .Z(n45901) );
  XNOR U45897 ( .A(n45922), .B(n45923), .Z(n45844) );
  AND U45898 ( .A(n1066), .B(n45924), .Z(n45923) );
  XNOR U45899 ( .A(n45925), .B(n45926), .Z(n45924) );
  XOR U45900 ( .A(n45927), .B(n45928), .Z(n45899) );
  AND U45901 ( .A(n45929), .B(n45930), .Z(n45928) );
  XNOR U45902 ( .A(n45927), .B(n45915), .Z(n45930) );
  IV U45903 ( .A(n45857), .Z(n45915) );
  XNOR U45904 ( .A(n45931), .B(n45908), .Z(n45857) );
  XNOR U45905 ( .A(n45932), .B(n45914), .Z(n45908) );
  XOR U45906 ( .A(n45933), .B(n45934), .Z(n45914) );
  AND U45907 ( .A(n45935), .B(n45936), .Z(n45934) );
  XOR U45908 ( .A(n45933), .B(n45937), .Z(n45935) );
  XNOR U45909 ( .A(n45913), .B(n45905), .Z(n45932) );
  XOR U45910 ( .A(n45938), .B(n45939), .Z(n45905) );
  AND U45911 ( .A(n45940), .B(n45941), .Z(n45939) );
  XNOR U45912 ( .A(n45942), .B(n45938), .Z(n45940) );
  XNOR U45913 ( .A(n45943), .B(n45910), .Z(n45913) );
  XOR U45914 ( .A(n45944), .B(n45945), .Z(n45910) );
  AND U45915 ( .A(n45946), .B(n45947), .Z(n45945) );
  XOR U45916 ( .A(n45944), .B(n45948), .Z(n45946) );
  XNOR U45917 ( .A(n45949), .B(n45950), .Z(n45943) );
  AND U45918 ( .A(n45951), .B(n45952), .Z(n45950) );
  XNOR U45919 ( .A(n45949), .B(n45953), .Z(n45951) );
  XNOR U45920 ( .A(n45909), .B(n45916), .Z(n45931) );
  AND U45921 ( .A(n45865), .B(n45954), .Z(n45916) );
  XOR U45922 ( .A(n45921), .B(n45920), .Z(n45909) );
  XNOR U45923 ( .A(n45955), .B(n45917), .Z(n45920) );
  XOR U45924 ( .A(n45956), .B(n45957), .Z(n45917) );
  AND U45925 ( .A(n45958), .B(n45959), .Z(n45957) );
  XOR U45926 ( .A(n45956), .B(n45960), .Z(n45958) );
  XNOR U45927 ( .A(n45961), .B(n45962), .Z(n45955) );
  AND U45928 ( .A(n45963), .B(n45964), .Z(n45962) );
  XOR U45929 ( .A(n45961), .B(n45965), .Z(n45963) );
  XOR U45930 ( .A(n45966), .B(n45967), .Z(n45921) );
  AND U45931 ( .A(n45968), .B(n45969), .Z(n45967) );
  XOR U45932 ( .A(n45966), .B(n45970), .Z(n45968) );
  XNOR U45933 ( .A(n45854), .B(n45927), .Z(n45929) );
  XNOR U45934 ( .A(n45971), .B(n45972), .Z(n45854) );
  AND U45935 ( .A(n1066), .B(n45973), .Z(n45972) );
  XNOR U45936 ( .A(n45974), .B(n45975), .Z(n45973) );
  XOR U45937 ( .A(n45976), .B(n45977), .Z(n45927) );
  AND U45938 ( .A(n45978), .B(n45979), .Z(n45977) );
  XNOR U45939 ( .A(n45976), .B(n45865), .Z(n45979) );
  XOR U45940 ( .A(n45980), .B(n45941), .Z(n45865) );
  XNOR U45941 ( .A(n45981), .B(n45948), .Z(n45941) );
  XOR U45942 ( .A(n45937), .B(n45936), .Z(n45948) );
  XNOR U45943 ( .A(n45982), .B(n45933), .Z(n45936) );
  XOR U45944 ( .A(n45983), .B(n45984), .Z(n45933) );
  AND U45945 ( .A(n45985), .B(n45986), .Z(n45984) );
  XNOR U45946 ( .A(n45987), .B(n45988), .Z(n45985) );
  IV U45947 ( .A(n45983), .Z(n45987) );
  XNOR U45948 ( .A(n45989), .B(n45990), .Z(n45982) );
  NOR U45949 ( .A(n45991), .B(n45992), .Z(n45990) );
  XNOR U45950 ( .A(n45989), .B(n45993), .Z(n45991) );
  XOR U45951 ( .A(n45994), .B(n45995), .Z(n45937) );
  NOR U45952 ( .A(n45996), .B(n45997), .Z(n45995) );
  XNOR U45953 ( .A(n45994), .B(n45998), .Z(n45996) );
  XNOR U45954 ( .A(n45947), .B(n45938), .Z(n45981) );
  XOR U45955 ( .A(n45999), .B(n46000), .Z(n45938) );
  AND U45956 ( .A(n46001), .B(n46002), .Z(n46000) );
  XOR U45957 ( .A(n45999), .B(n46003), .Z(n46001) );
  XOR U45958 ( .A(n46004), .B(n45953), .Z(n45947) );
  XOR U45959 ( .A(n46005), .B(n46006), .Z(n45953) );
  NOR U45960 ( .A(n46007), .B(n46008), .Z(n46006) );
  XOR U45961 ( .A(n46005), .B(n46009), .Z(n46007) );
  XNOR U45962 ( .A(n45952), .B(n45944), .Z(n46004) );
  XOR U45963 ( .A(n46010), .B(n46011), .Z(n45944) );
  AND U45964 ( .A(n46012), .B(n46013), .Z(n46011) );
  XOR U45965 ( .A(n46010), .B(n46014), .Z(n46012) );
  XNOR U45966 ( .A(n46015), .B(n45949), .Z(n45952) );
  XOR U45967 ( .A(n46016), .B(n46017), .Z(n45949) );
  AND U45968 ( .A(n46018), .B(n46019), .Z(n46017) );
  XNOR U45969 ( .A(n46020), .B(n46021), .Z(n46018) );
  IV U45970 ( .A(n46016), .Z(n46020) );
  XNOR U45971 ( .A(n46022), .B(n46023), .Z(n46015) );
  NOR U45972 ( .A(n46024), .B(n46025), .Z(n46023) );
  XNOR U45973 ( .A(n46022), .B(n46026), .Z(n46024) );
  XOR U45974 ( .A(n45942), .B(n45954), .Z(n45980) );
  NOR U45975 ( .A(n45871), .B(n46027), .Z(n45954) );
  XNOR U45976 ( .A(n45960), .B(n45959), .Z(n45942) );
  XNOR U45977 ( .A(n46028), .B(n45965), .Z(n45959) );
  XNOR U45978 ( .A(n46029), .B(n46030), .Z(n45965) );
  NOR U45979 ( .A(n46031), .B(n46032), .Z(n46030) );
  XOR U45980 ( .A(n46029), .B(n46033), .Z(n46031) );
  XNOR U45981 ( .A(n45964), .B(n45956), .Z(n46028) );
  XOR U45982 ( .A(n46034), .B(n46035), .Z(n45956) );
  AND U45983 ( .A(n46036), .B(n46037), .Z(n46035) );
  XOR U45984 ( .A(n46034), .B(n46038), .Z(n46036) );
  XNOR U45985 ( .A(n46039), .B(n45961), .Z(n45964) );
  XOR U45986 ( .A(n46040), .B(n46041), .Z(n45961) );
  AND U45987 ( .A(n46042), .B(n46043), .Z(n46041) );
  XNOR U45988 ( .A(n46044), .B(n46045), .Z(n46042) );
  IV U45989 ( .A(n46040), .Z(n46044) );
  XNOR U45990 ( .A(n46046), .B(n46047), .Z(n46039) );
  NOR U45991 ( .A(n46048), .B(n46049), .Z(n46047) );
  XNOR U45992 ( .A(n46046), .B(n46050), .Z(n46048) );
  XOR U45993 ( .A(n45970), .B(n45969), .Z(n45960) );
  XNOR U45994 ( .A(n46051), .B(n45966), .Z(n45969) );
  XOR U45995 ( .A(n46052), .B(n46053), .Z(n45966) );
  AND U45996 ( .A(n46054), .B(n46055), .Z(n46053) );
  XNOR U45997 ( .A(n46056), .B(n46057), .Z(n46054) );
  IV U45998 ( .A(n46052), .Z(n46056) );
  XNOR U45999 ( .A(n46058), .B(n46059), .Z(n46051) );
  NOR U46000 ( .A(n46060), .B(n46061), .Z(n46059) );
  XNOR U46001 ( .A(n46058), .B(n46062), .Z(n46060) );
  XOR U46002 ( .A(n46063), .B(n46064), .Z(n45970) );
  NOR U46003 ( .A(n46065), .B(n46066), .Z(n46064) );
  XNOR U46004 ( .A(n46063), .B(n46067), .Z(n46065) );
  XNOR U46005 ( .A(n45862), .B(n45976), .Z(n45978) );
  XNOR U46006 ( .A(n46068), .B(n46069), .Z(n45862) );
  AND U46007 ( .A(n1066), .B(n46070), .Z(n46069) );
  XNOR U46008 ( .A(n46071), .B(n46072), .Z(n46070) );
  AND U46009 ( .A(n45868), .B(n45871), .Z(n45976) );
  XOR U46010 ( .A(n46073), .B(n46027), .Z(n45871) );
  XNOR U46011 ( .A(p_input[1568]), .B(p_input[2048]), .Z(n46027) );
  XNOR U46012 ( .A(n46003), .B(n46002), .Z(n46073) );
  XNOR U46013 ( .A(n46074), .B(n46014), .Z(n46002) );
  XOR U46014 ( .A(n45988), .B(n45986), .Z(n46014) );
  XNOR U46015 ( .A(n46075), .B(n45993), .Z(n45986) );
  XOR U46016 ( .A(p_input[1592]), .B(p_input[2072]), .Z(n45993) );
  XOR U46017 ( .A(n45983), .B(n45992), .Z(n46075) );
  XOR U46018 ( .A(n46076), .B(n45989), .Z(n45992) );
  XOR U46019 ( .A(p_input[1590]), .B(p_input[2070]), .Z(n45989) );
  XOR U46020 ( .A(p_input[1591]), .B(n29410), .Z(n46076) );
  XOR U46021 ( .A(p_input[1586]), .B(p_input[2066]), .Z(n45983) );
  XNOR U46022 ( .A(n45998), .B(n45997), .Z(n45988) );
  XOR U46023 ( .A(n46077), .B(n45994), .Z(n45997) );
  XOR U46024 ( .A(p_input[1587]), .B(p_input[2067]), .Z(n45994) );
  XOR U46025 ( .A(p_input[1588]), .B(n29412), .Z(n46077) );
  XOR U46026 ( .A(p_input[1589]), .B(p_input[2069]), .Z(n45998) );
  XOR U46027 ( .A(n46013), .B(n46078), .Z(n46074) );
  IV U46028 ( .A(n45999), .Z(n46078) );
  XOR U46029 ( .A(p_input[1569]), .B(p_input[2049]), .Z(n45999) );
  XNOR U46030 ( .A(n46079), .B(n46021), .Z(n46013) );
  XNOR U46031 ( .A(n46009), .B(n46008), .Z(n46021) );
  XNOR U46032 ( .A(n46080), .B(n46005), .Z(n46008) );
  XNOR U46033 ( .A(p_input[1594]), .B(p_input[2074]), .Z(n46005) );
  XOR U46034 ( .A(p_input[1595]), .B(n29415), .Z(n46080) );
  XOR U46035 ( .A(p_input[1596]), .B(p_input[2076]), .Z(n46009) );
  XOR U46036 ( .A(n46019), .B(n46081), .Z(n46079) );
  IV U46037 ( .A(n46010), .Z(n46081) );
  XOR U46038 ( .A(p_input[1585]), .B(p_input[2065]), .Z(n46010) );
  XNOR U46039 ( .A(n46082), .B(n46026), .Z(n46019) );
  XNOR U46040 ( .A(p_input[1599]), .B(n29418), .Z(n46026) );
  XOR U46041 ( .A(n46016), .B(n46025), .Z(n46082) );
  XOR U46042 ( .A(n46083), .B(n46022), .Z(n46025) );
  XOR U46043 ( .A(p_input[1597]), .B(p_input[2077]), .Z(n46022) );
  XOR U46044 ( .A(p_input[1598]), .B(n29420), .Z(n46083) );
  XOR U46045 ( .A(p_input[1593]), .B(p_input[2073]), .Z(n46016) );
  XOR U46046 ( .A(n46038), .B(n46037), .Z(n46003) );
  XNOR U46047 ( .A(n46084), .B(n46045), .Z(n46037) );
  XNOR U46048 ( .A(n46033), .B(n46032), .Z(n46045) );
  XNOR U46049 ( .A(n46085), .B(n46029), .Z(n46032) );
  XNOR U46050 ( .A(p_input[1579]), .B(p_input[2059]), .Z(n46029) );
  XOR U46051 ( .A(p_input[1580]), .B(n28329), .Z(n46085) );
  XOR U46052 ( .A(p_input[1581]), .B(p_input[2061]), .Z(n46033) );
  XOR U46053 ( .A(n46043), .B(n46086), .Z(n46084) );
  IV U46054 ( .A(n46034), .Z(n46086) );
  XOR U46055 ( .A(p_input[1570]), .B(p_input[2050]), .Z(n46034) );
  XNOR U46056 ( .A(n46087), .B(n46050), .Z(n46043) );
  XNOR U46057 ( .A(p_input[1584]), .B(n28332), .Z(n46050) );
  XOR U46058 ( .A(n46040), .B(n46049), .Z(n46087) );
  XOR U46059 ( .A(n46088), .B(n46046), .Z(n46049) );
  XOR U46060 ( .A(p_input[1582]), .B(p_input[2062]), .Z(n46046) );
  XOR U46061 ( .A(p_input[1583]), .B(n28334), .Z(n46088) );
  XOR U46062 ( .A(p_input[1578]), .B(p_input[2058]), .Z(n46040) );
  XOR U46063 ( .A(n46057), .B(n46055), .Z(n46038) );
  XNOR U46064 ( .A(n46089), .B(n46062), .Z(n46055) );
  XOR U46065 ( .A(p_input[1577]), .B(p_input[2057]), .Z(n46062) );
  XOR U46066 ( .A(n46052), .B(n46061), .Z(n46089) );
  XOR U46067 ( .A(n46090), .B(n46058), .Z(n46061) );
  XOR U46068 ( .A(p_input[1575]), .B(p_input[2055]), .Z(n46058) );
  XOR U46069 ( .A(p_input[1576]), .B(n29427), .Z(n46090) );
  XOR U46070 ( .A(p_input[1571]), .B(p_input[2051]), .Z(n46052) );
  XNOR U46071 ( .A(n46067), .B(n46066), .Z(n46057) );
  XOR U46072 ( .A(n46091), .B(n46063), .Z(n46066) );
  XOR U46073 ( .A(p_input[1572]), .B(p_input[2052]), .Z(n46063) );
  XOR U46074 ( .A(p_input[1573]), .B(n29429), .Z(n46091) );
  XOR U46075 ( .A(p_input[1574]), .B(p_input[2054]), .Z(n46067) );
  XNOR U46076 ( .A(n46092), .B(n46093), .Z(n45868) );
  AND U46077 ( .A(n1066), .B(n46094), .Z(n46093) );
  XNOR U46078 ( .A(n46095), .B(n46096), .Z(n1066) );
  AND U46079 ( .A(n46097), .B(n46098), .Z(n46096) );
  XOR U46080 ( .A(n45882), .B(n46095), .Z(n46098) );
  XNOR U46081 ( .A(n46099), .B(n46095), .Z(n46097) );
  XOR U46082 ( .A(n46100), .B(n46101), .Z(n46095) );
  AND U46083 ( .A(n46102), .B(n46103), .Z(n46101) );
  XOR U46084 ( .A(n45897), .B(n46100), .Z(n46103) );
  XOR U46085 ( .A(n46100), .B(n45898), .Z(n46102) );
  XOR U46086 ( .A(n46104), .B(n46105), .Z(n46100) );
  AND U46087 ( .A(n46106), .B(n46107), .Z(n46105) );
  XOR U46088 ( .A(n45925), .B(n46104), .Z(n46107) );
  XOR U46089 ( .A(n46104), .B(n45926), .Z(n46106) );
  XOR U46090 ( .A(n46108), .B(n46109), .Z(n46104) );
  AND U46091 ( .A(n46110), .B(n46111), .Z(n46109) );
  XOR U46092 ( .A(n45974), .B(n46108), .Z(n46111) );
  XOR U46093 ( .A(n46108), .B(n45975), .Z(n46110) );
  XOR U46094 ( .A(n46112), .B(n46113), .Z(n46108) );
  AND U46095 ( .A(n46114), .B(n46115), .Z(n46113) );
  XOR U46096 ( .A(n46112), .B(n46071), .Z(n46115) );
  XNOR U46097 ( .A(n46116), .B(n46117), .Z(n45818) );
  AND U46098 ( .A(n1070), .B(n46118), .Z(n46117) );
  XNOR U46099 ( .A(n46119), .B(n46120), .Z(n1070) );
  AND U46100 ( .A(n46121), .B(n46122), .Z(n46120) );
  XOR U46101 ( .A(n46119), .B(n45828), .Z(n46122) );
  XNOR U46102 ( .A(n46119), .B(n45778), .Z(n46121) );
  XOR U46103 ( .A(n46123), .B(n46124), .Z(n46119) );
  AND U46104 ( .A(n46125), .B(n46126), .Z(n46124) );
  XNOR U46105 ( .A(n45838), .B(n46123), .Z(n46126) );
  XOR U46106 ( .A(n46123), .B(n45788), .Z(n46125) );
  XOR U46107 ( .A(n46127), .B(n46128), .Z(n46123) );
  AND U46108 ( .A(n46129), .B(n46130), .Z(n46128) );
  XNOR U46109 ( .A(n45848), .B(n46127), .Z(n46130) );
  XOR U46110 ( .A(n46127), .B(n45797), .Z(n46129) );
  XOR U46111 ( .A(n46131), .B(n46132), .Z(n46127) );
  AND U46112 ( .A(n46133), .B(n46134), .Z(n46132) );
  XOR U46113 ( .A(n46131), .B(n45805), .Z(n46133) );
  XOR U46114 ( .A(n46135), .B(n46136), .Z(n45769) );
  AND U46115 ( .A(n1074), .B(n46118), .Z(n46136) );
  XNOR U46116 ( .A(n46116), .B(n46135), .Z(n46118) );
  XNOR U46117 ( .A(n46137), .B(n46138), .Z(n1074) );
  AND U46118 ( .A(n46139), .B(n46140), .Z(n46138) );
  XNOR U46119 ( .A(n46141), .B(n46137), .Z(n46140) );
  IV U46120 ( .A(n45828), .Z(n46141) );
  XOR U46121 ( .A(n46099), .B(n46142), .Z(n45828) );
  AND U46122 ( .A(n1077), .B(n46143), .Z(n46142) );
  XOR U46123 ( .A(n45881), .B(n45878), .Z(n46143) );
  IV U46124 ( .A(n46099), .Z(n45881) );
  XNOR U46125 ( .A(n45778), .B(n46137), .Z(n46139) );
  XOR U46126 ( .A(n46144), .B(n46145), .Z(n45778) );
  AND U46127 ( .A(n1093), .B(n46146), .Z(n46145) );
  XOR U46128 ( .A(n46147), .B(n46148), .Z(n46137) );
  AND U46129 ( .A(n46149), .B(n46150), .Z(n46148) );
  XNOR U46130 ( .A(n46147), .B(n45838), .Z(n46150) );
  XOR U46131 ( .A(n45898), .B(n46151), .Z(n45838) );
  AND U46132 ( .A(n1077), .B(n46152), .Z(n46151) );
  XOR U46133 ( .A(n45894), .B(n45898), .Z(n46152) );
  XNOR U46134 ( .A(n46153), .B(n46147), .Z(n46149) );
  IV U46135 ( .A(n45788), .Z(n46153) );
  XOR U46136 ( .A(n46154), .B(n46155), .Z(n45788) );
  AND U46137 ( .A(n1093), .B(n46156), .Z(n46155) );
  XOR U46138 ( .A(n46157), .B(n46158), .Z(n46147) );
  AND U46139 ( .A(n46159), .B(n46160), .Z(n46158) );
  XNOR U46140 ( .A(n46157), .B(n45848), .Z(n46160) );
  XOR U46141 ( .A(n45926), .B(n46161), .Z(n45848) );
  AND U46142 ( .A(n1077), .B(n46162), .Z(n46161) );
  XOR U46143 ( .A(n45922), .B(n45926), .Z(n46162) );
  XOR U46144 ( .A(n45797), .B(n46157), .Z(n46159) );
  XOR U46145 ( .A(n46163), .B(n46164), .Z(n45797) );
  AND U46146 ( .A(n1093), .B(n46165), .Z(n46164) );
  XOR U46147 ( .A(n46131), .B(n46166), .Z(n46157) );
  AND U46148 ( .A(n46167), .B(n46134), .Z(n46166) );
  XNOR U46149 ( .A(n45858), .B(n46131), .Z(n46134) );
  XOR U46150 ( .A(n45975), .B(n46168), .Z(n45858) );
  AND U46151 ( .A(n1077), .B(n46169), .Z(n46168) );
  XOR U46152 ( .A(n45971), .B(n45975), .Z(n46169) );
  XNOR U46153 ( .A(n46170), .B(n46131), .Z(n46167) );
  IV U46154 ( .A(n45805), .Z(n46170) );
  XOR U46155 ( .A(n46171), .B(n46172), .Z(n45805) );
  AND U46156 ( .A(n1093), .B(n46173), .Z(n46172) );
  XOR U46157 ( .A(n46174), .B(n46175), .Z(n46131) );
  AND U46158 ( .A(n46176), .B(n46177), .Z(n46175) );
  XNOR U46159 ( .A(n46174), .B(n45866), .Z(n46177) );
  XOR U46160 ( .A(n46072), .B(n46178), .Z(n45866) );
  AND U46161 ( .A(n1077), .B(n46179), .Z(n46178) );
  XOR U46162 ( .A(n46068), .B(n46072), .Z(n46179) );
  XNOR U46163 ( .A(n46180), .B(n46174), .Z(n46176) );
  IV U46164 ( .A(n45815), .Z(n46180) );
  XOR U46165 ( .A(n46181), .B(n46182), .Z(n45815) );
  AND U46166 ( .A(n1093), .B(n46183), .Z(n46182) );
  AND U46167 ( .A(n46135), .B(n46116), .Z(n46174) );
  XNOR U46168 ( .A(n46184), .B(n46185), .Z(n46116) );
  AND U46169 ( .A(n1077), .B(n46094), .Z(n46185) );
  XNOR U46170 ( .A(n46092), .B(n46184), .Z(n46094) );
  XNOR U46171 ( .A(n46186), .B(n46187), .Z(n1077) );
  AND U46172 ( .A(n46188), .B(n46189), .Z(n46187) );
  XNOR U46173 ( .A(n46186), .B(n45878), .Z(n46189) );
  IV U46174 ( .A(n45882), .Z(n45878) );
  XOR U46175 ( .A(n46190), .B(n46191), .Z(n45882) );
  AND U46176 ( .A(n1081), .B(n46192), .Z(n46191) );
  XOR U46177 ( .A(n46193), .B(n46190), .Z(n46192) );
  XNOR U46178 ( .A(n46186), .B(n46099), .Z(n46188) );
  XOR U46179 ( .A(n46194), .B(n46195), .Z(n46099) );
  AND U46180 ( .A(n1089), .B(n46146), .Z(n46195) );
  XOR U46181 ( .A(n46144), .B(n46194), .Z(n46146) );
  XOR U46182 ( .A(n46196), .B(n46197), .Z(n46186) );
  AND U46183 ( .A(n46198), .B(n46199), .Z(n46197) );
  XNOR U46184 ( .A(n46196), .B(n45894), .Z(n46199) );
  IV U46185 ( .A(n45897), .Z(n45894) );
  XOR U46186 ( .A(n46200), .B(n46201), .Z(n45897) );
  AND U46187 ( .A(n1081), .B(n46202), .Z(n46201) );
  XOR U46188 ( .A(n46203), .B(n46200), .Z(n46202) );
  XOR U46189 ( .A(n45898), .B(n46196), .Z(n46198) );
  XOR U46190 ( .A(n46204), .B(n46205), .Z(n45898) );
  AND U46191 ( .A(n1089), .B(n46156), .Z(n46205) );
  XOR U46192 ( .A(n46204), .B(n46154), .Z(n46156) );
  XOR U46193 ( .A(n46206), .B(n46207), .Z(n46196) );
  AND U46194 ( .A(n46208), .B(n46209), .Z(n46207) );
  XNOR U46195 ( .A(n46206), .B(n45922), .Z(n46209) );
  IV U46196 ( .A(n45925), .Z(n45922) );
  XOR U46197 ( .A(n46210), .B(n46211), .Z(n45925) );
  AND U46198 ( .A(n1081), .B(n46212), .Z(n46211) );
  XNOR U46199 ( .A(n46213), .B(n46210), .Z(n46212) );
  XOR U46200 ( .A(n45926), .B(n46206), .Z(n46208) );
  XOR U46201 ( .A(n46214), .B(n46215), .Z(n45926) );
  AND U46202 ( .A(n1089), .B(n46165), .Z(n46215) );
  XOR U46203 ( .A(n46214), .B(n46163), .Z(n46165) );
  XOR U46204 ( .A(n46216), .B(n46217), .Z(n46206) );
  AND U46205 ( .A(n46218), .B(n46219), .Z(n46217) );
  XNOR U46206 ( .A(n46216), .B(n45971), .Z(n46219) );
  IV U46207 ( .A(n45974), .Z(n45971) );
  XOR U46208 ( .A(n46220), .B(n46221), .Z(n45974) );
  AND U46209 ( .A(n1081), .B(n46222), .Z(n46221) );
  XOR U46210 ( .A(n46223), .B(n46220), .Z(n46222) );
  XOR U46211 ( .A(n45975), .B(n46216), .Z(n46218) );
  XOR U46212 ( .A(n46224), .B(n46225), .Z(n45975) );
  AND U46213 ( .A(n1089), .B(n46173), .Z(n46225) );
  XOR U46214 ( .A(n46224), .B(n46171), .Z(n46173) );
  XOR U46215 ( .A(n46112), .B(n46226), .Z(n46216) );
  AND U46216 ( .A(n46114), .B(n46227), .Z(n46226) );
  XNOR U46217 ( .A(n46112), .B(n46068), .Z(n46227) );
  IV U46218 ( .A(n46071), .Z(n46068) );
  XOR U46219 ( .A(n46228), .B(n46229), .Z(n46071) );
  AND U46220 ( .A(n1081), .B(n46230), .Z(n46229) );
  XNOR U46221 ( .A(n46231), .B(n46228), .Z(n46230) );
  XOR U46222 ( .A(n46072), .B(n46112), .Z(n46114) );
  XOR U46223 ( .A(n46232), .B(n46233), .Z(n46072) );
  AND U46224 ( .A(n1089), .B(n46183), .Z(n46233) );
  XOR U46225 ( .A(n46232), .B(n46181), .Z(n46183) );
  AND U46226 ( .A(n46184), .B(n46092), .Z(n46112) );
  XNOR U46227 ( .A(n46234), .B(n46235), .Z(n46092) );
  AND U46228 ( .A(n1081), .B(n46236), .Z(n46235) );
  XNOR U46229 ( .A(n46237), .B(n46234), .Z(n46236) );
  XNOR U46230 ( .A(n46238), .B(n46239), .Z(n1081) );
  AND U46231 ( .A(n46240), .B(n46241), .Z(n46239) );
  XOR U46232 ( .A(n46193), .B(n46238), .Z(n46241) );
  AND U46233 ( .A(n46242), .B(n46243), .Z(n46193) );
  XNOR U46234 ( .A(n46190), .B(n46238), .Z(n46240) );
  XNOR U46235 ( .A(n46244), .B(n46245), .Z(n46190) );
  AND U46236 ( .A(n1085), .B(n46246), .Z(n46245) );
  XNOR U46237 ( .A(n46247), .B(n46248), .Z(n46246) );
  XOR U46238 ( .A(n46249), .B(n46250), .Z(n46238) );
  AND U46239 ( .A(n46251), .B(n46252), .Z(n46250) );
  XNOR U46240 ( .A(n46249), .B(n46242), .Z(n46252) );
  IV U46241 ( .A(n46203), .Z(n46242) );
  XOR U46242 ( .A(n46253), .B(n46254), .Z(n46203) );
  XOR U46243 ( .A(n46255), .B(n46243), .Z(n46254) );
  AND U46244 ( .A(n46213), .B(n46256), .Z(n46243) );
  AND U46245 ( .A(n46257), .B(n46258), .Z(n46255) );
  XOR U46246 ( .A(n46259), .B(n46253), .Z(n46257) );
  XNOR U46247 ( .A(n46200), .B(n46249), .Z(n46251) );
  XNOR U46248 ( .A(n46260), .B(n46261), .Z(n46200) );
  AND U46249 ( .A(n1085), .B(n46262), .Z(n46261) );
  XNOR U46250 ( .A(n46263), .B(n46264), .Z(n46262) );
  XOR U46251 ( .A(n46265), .B(n46266), .Z(n46249) );
  AND U46252 ( .A(n46267), .B(n46268), .Z(n46266) );
  XNOR U46253 ( .A(n46265), .B(n46213), .Z(n46268) );
  XOR U46254 ( .A(n46269), .B(n46258), .Z(n46213) );
  XNOR U46255 ( .A(n46270), .B(n46253), .Z(n46258) );
  XOR U46256 ( .A(n46271), .B(n46272), .Z(n46253) );
  AND U46257 ( .A(n46273), .B(n46274), .Z(n46272) );
  XOR U46258 ( .A(n46275), .B(n46271), .Z(n46273) );
  XNOR U46259 ( .A(n46276), .B(n46277), .Z(n46270) );
  AND U46260 ( .A(n46278), .B(n46279), .Z(n46277) );
  XOR U46261 ( .A(n46276), .B(n46280), .Z(n46278) );
  XNOR U46262 ( .A(n46259), .B(n46256), .Z(n46269) );
  AND U46263 ( .A(n46281), .B(n46282), .Z(n46256) );
  XOR U46264 ( .A(n46283), .B(n46284), .Z(n46259) );
  AND U46265 ( .A(n46285), .B(n46286), .Z(n46284) );
  XOR U46266 ( .A(n46283), .B(n46287), .Z(n46285) );
  XNOR U46267 ( .A(n46210), .B(n46265), .Z(n46267) );
  XNOR U46268 ( .A(n46288), .B(n46289), .Z(n46210) );
  AND U46269 ( .A(n1085), .B(n46290), .Z(n46289) );
  XNOR U46270 ( .A(n46291), .B(n46292), .Z(n46290) );
  XOR U46271 ( .A(n46293), .B(n46294), .Z(n46265) );
  AND U46272 ( .A(n46295), .B(n46296), .Z(n46294) );
  XNOR U46273 ( .A(n46293), .B(n46281), .Z(n46296) );
  IV U46274 ( .A(n46223), .Z(n46281) );
  XNOR U46275 ( .A(n46297), .B(n46274), .Z(n46223) );
  XNOR U46276 ( .A(n46298), .B(n46280), .Z(n46274) );
  XOR U46277 ( .A(n46299), .B(n46300), .Z(n46280) );
  AND U46278 ( .A(n46301), .B(n46302), .Z(n46300) );
  XOR U46279 ( .A(n46299), .B(n46303), .Z(n46301) );
  XNOR U46280 ( .A(n46279), .B(n46271), .Z(n46298) );
  XOR U46281 ( .A(n46304), .B(n46305), .Z(n46271) );
  AND U46282 ( .A(n46306), .B(n46307), .Z(n46305) );
  XNOR U46283 ( .A(n46308), .B(n46304), .Z(n46306) );
  XNOR U46284 ( .A(n46309), .B(n46276), .Z(n46279) );
  XOR U46285 ( .A(n46310), .B(n46311), .Z(n46276) );
  AND U46286 ( .A(n46312), .B(n46313), .Z(n46311) );
  XOR U46287 ( .A(n46310), .B(n46314), .Z(n46312) );
  XNOR U46288 ( .A(n46315), .B(n46316), .Z(n46309) );
  AND U46289 ( .A(n46317), .B(n46318), .Z(n46316) );
  XNOR U46290 ( .A(n46315), .B(n46319), .Z(n46317) );
  XNOR U46291 ( .A(n46275), .B(n46282), .Z(n46297) );
  AND U46292 ( .A(n46231), .B(n46320), .Z(n46282) );
  XOR U46293 ( .A(n46287), .B(n46286), .Z(n46275) );
  XNOR U46294 ( .A(n46321), .B(n46283), .Z(n46286) );
  XOR U46295 ( .A(n46322), .B(n46323), .Z(n46283) );
  AND U46296 ( .A(n46324), .B(n46325), .Z(n46323) );
  XOR U46297 ( .A(n46322), .B(n46326), .Z(n46324) );
  XNOR U46298 ( .A(n46327), .B(n46328), .Z(n46321) );
  AND U46299 ( .A(n46329), .B(n46330), .Z(n46328) );
  XOR U46300 ( .A(n46327), .B(n46331), .Z(n46329) );
  XOR U46301 ( .A(n46332), .B(n46333), .Z(n46287) );
  AND U46302 ( .A(n46334), .B(n46335), .Z(n46333) );
  XOR U46303 ( .A(n46332), .B(n46336), .Z(n46334) );
  XNOR U46304 ( .A(n46220), .B(n46293), .Z(n46295) );
  XNOR U46305 ( .A(n46337), .B(n46338), .Z(n46220) );
  AND U46306 ( .A(n1085), .B(n46339), .Z(n46338) );
  XNOR U46307 ( .A(n46340), .B(n46341), .Z(n46339) );
  XOR U46308 ( .A(n46342), .B(n46343), .Z(n46293) );
  AND U46309 ( .A(n46344), .B(n46345), .Z(n46343) );
  XNOR U46310 ( .A(n46342), .B(n46231), .Z(n46345) );
  XOR U46311 ( .A(n46346), .B(n46307), .Z(n46231) );
  XNOR U46312 ( .A(n46347), .B(n46314), .Z(n46307) );
  XOR U46313 ( .A(n46303), .B(n46302), .Z(n46314) );
  XNOR U46314 ( .A(n46348), .B(n46299), .Z(n46302) );
  XOR U46315 ( .A(n46349), .B(n46350), .Z(n46299) );
  AND U46316 ( .A(n46351), .B(n46352), .Z(n46350) );
  XNOR U46317 ( .A(n46353), .B(n46354), .Z(n46351) );
  IV U46318 ( .A(n46349), .Z(n46353) );
  XNOR U46319 ( .A(n46355), .B(n46356), .Z(n46348) );
  NOR U46320 ( .A(n46357), .B(n46358), .Z(n46356) );
  XNOR U46321 ( .A(n46355), .B(n46359), .Z(n46357) );
  XOR U46322 ( .A(n46360), .B(n46361), .Z(n46303) );
  NOR U46323 ( .A(n46362), .B(n46363), .Z(n46361) );
  XNOR U46324 ( .A(n46360), .B(n46364), .Z(n46362) );
  XNOR U46325 ( .A(n46313), .B(n46304), .Z(n46347) );
  XOR U46326 ( .A(n46365), .B(n46366), .Z(n46304) );
  AND U46327 ( .A(n46367), .B(n46368), .Z(n46366) );
  XOR U46328 ( .A(n46365), .B(n46369), .Z(n46367) );
  XOR U46329 ( .A(n46370), .B(n46319), .Z(n46313) );
  XOR U46330 ( .A(n46371), .B(n46372), .Z(n46319) );
  NOR U46331 ( .A(n46373), .B(n46374), .Z(n46372) );
  XOR U46332 ( .A(n46371), .B(n46375), .Z(n46373) );
  XNOR U46333 ( .A(n46318), .B(n46310), .Z(n46370) );
  XOR U46334 ( .A(n46376), .B(n46377), .Z(n46310) );
  AND U46335 ( .A(n46378), .B(n46379), .Z(n46377) );
  XOR U46336 ( .A(n46376), .B(n46380), .Z(n46378) );
  XNOR U46337 ( .A(n46381), .B(n46315), .Z(n46318) );
  XOR U46338 ( .A(n46382), .B(n46383), .Z(n46315) );
  AND U46339 ( .A(n46384), .B(n46385), .Z(n46383) );
  XNOR U46340 ( .A(n46386), .B(n46387), .Z(n46384) );
  IV U46341 ( .A(n46382), .Z(n46386) );
  XNOR U46342 ( .A(n46388), .B(n46389), .Z(n46381) );
  NOR U46343 ( .A(n46390), .B(n46391), .Z(n46389) );
  XNOR U46344 ( .A(n46388), .B(n46392), .Z(n46390) );
  XOR U46345 ( .A(n46308), .B(n46320), .Z(n46346) );
  NOR U46346 ( .A(n46237), .B(n46393), .Z(n46320) );
  XNOR U46347 ( .A(n46326), .B(n46325), .Z(n46308) );
  XNOR U46348 ( .A(n46394), .B(n46331), .Z(n46325) );
  XNOR U46349 ( .A(n46395), .B(n46396), .Z(n46331) );
  NOR U46350 ( .A(n46397), .B(n46398), .Z(n46396) );
  XOR U46351 ( .A(n46395), .B(n46399), .Z(n46397) );
  XNOR U46352 ( .A(n46330), .B(n46322), .Z(n46394) );
  XOR U46353 ( .A(n46400), .B(n46401), .Z(n46322) );
  AND U46354 ( .A(n46402), .B(n46403), .Z(n46401) );
  XOR U46355 ( .A(n46400), .B(n46404), .Z(n46402) );
  XNOR U46356 ( .A(n46405), .B(n46327), .Z(n46330) );
  XOR U46357 ( .A(n46406), .B(n46407), .Z(n46327) );
  AND U46358 ( .A(n46408), .B(n46409), .Z(n46407) );
  XNOR U46359 ( .A(n46410), .B(n46411), .Z(n46408) );
  IV U46360 ( .A(n46406), .Z(n46410) );
  XNOR U46361 ( .A(n46412), .B(n46413), .Z(n46405) );
  NOR U46362 ( .A(n46414), .B(n46415), .Z(n46413) );
  XNOR U46363 ( .A(n46412), .B(n46416), .Z(n46414) );
  XOR U46364 ( .A(n46336), .B(n46335), .Z(n46326) );
  XNOR U46365 ( .A(n46417), .B(n46332), .Z(n46335) );
  XOR U46366 ( .A(n46418), .B(n46419), .Z(n46332) );
  AND U46367 ( .A(n46420), .B(n46421), .Z(n46419) );
  XNOR U46368 ( .A(n46422), .B(n46423), .Z(n46420) );
  IV U46369 ( .A(n46418), .Z(n46422) );
  XNOR U46370 ( .A(n46424), .B(n46425), .Z(n46417) );
  NOR U46371 ( .A(n46426), .B(n46427), .Z(n46425) );
  XNOR U46372 ( .A(n46424), .B(n46428), .Z(n46426) );
  XOR U46373 ( .A(n46429), .B(n46430), .Z(n46336) );
  NOR U46374 ( .A(n46431), .B(n46432), .Z(n46430) );
  XNOR U46375 ( .A(n46429), .B(n46433), .Z(n46431) );
  XNOR U46376 ( .A(n46228), .B(n46342), .Z(n46344) );
  XNOR U46377 ( .A(n46434), .B(n46435), .Z(n46228) );
  AND U46378 ( .A(n1085), .B(n46436), .Z(n46435) );
  XNOR U46379 ( .A(n46437), .B(n46438), .Z(n46436) );
  AND U46380 ( .A(n46234), .B(n46237), .Z(n46342) );
  XOR U46381 ( .A(n46439), .B(n46393), .Z(n46237) );
  XNOR U46382 ( .A(p_input[1600]), .B(p_input[2048]), .Z(n46393) );
  XNOR U46383 ( .A(n46369), .B(n46368), .Z(n46439) );
  XNOR U46384 ( .A(n46440), .B(n46380), .Z(n46368) );
  XOR U46385 ( .A(n46354), .B(n46352), .Z(n46380) );
  XNOR U46386 ( .A(n46441), .B(n46359), .Z(n46352) );
  XOR U46387 ( .A(p_input[1624]), .B(p_input[2072]), .Z(n46359) );
  XOR U46388 ( .A(n46349), .B(n46358), .Z(n46441) );
  XOR U46389 ( .A(n46442), .B(n46355), .Z(n46358) );
  XOR U46390 ( .A(p_input[1622]), .B(p_input[2070]), .Z(n46355) );
  XOR U46391 ( .A(p_input[1623]), .B(n29410), .Z(n46442) );
  XOR U46392 ( .A(p_input[1618]), .B(p_input[2066]), .Z(n46349) );
  XNOR U46393 ( .A(n46364), .B(n46363), .Z(n46354) );
  XOR U46394 ( .A(n46443), .B(n46360), .Z(n46363) );
  XOR U46395 ( .A(p_input[1619]), .B(p_input[2067]), .Z(n46360) );
  XOR U46396 ( .A(p_input[1620]), .B(n29412), .Z(n46443) );
  XOR U46397 ( .A(p_input[1621]), .B(p_input[2069]), .Z(n46364) );
  XOR U46398 ( .A(n46379), .B(n46444), .Z(n46440) );
  IV U46399 ( .A(n46365), .Z(n46444) );
  XOR U46400 ( .A(p_input[1601]), .B(p_input[2049]), .Z(n46365) );
  XNOR U46401 ( .A(n46445), .B(n46387), .Z(n46379) );
  XNOR U46402 ( .A(n46375), .B(n46374), .Z(n46387) );
  XNOR U46403 ( .A(n46446), .B(n46371), .Z(n46374) );
  XNOR U46404 ( .A(p_input[1626]), .B(p_input[2074]), .Z(n46371) );
  XOR U46405 ( .A(p_input[1627]), .B(n29415), .Z(n46446) );
  XOR U46406 ( .A(p_input[1628]), .B(p_input[2076]), .Z(n46375) );
  XOR U46407 ( .A(n46385), .B(n46447), .Z(n46445) );
  IV U46408 ( .A(n46376), .Z(n46447) );
  XOR U46409 ( .A(p_input[1617]), .B(p_input[2065]), .Z(n46376) );
  XNOR U46410 ( .A(n46448), .B(n46392), .Z(n46385) );
  XNOR U46411 ( .A(p_input[1631]), .B(n29418), .Z(n46392) );
  XOR U46412 ( .A(n46382), .B(n46391), .Z(n46448) );
  XOR U46413 ( .A(n46449), .B(n46388), .Z(n46391) );
  XOR U46414 ( .A(p_input[1629]), .B(p_input[2077]), .Z(n46388) );
  XOR U46415 ( .A(p_input[1630]), .B(n29420), .Z(n46449) );
  XOR U46416 ( .A(p_input[1625]), .B(p_input[2073]), .Z(n46382) );
  XOR U46417 ( .A(n46404), .B(n46403), .Z(n46369) );
  XNOR U46418 ( .A(n46450), .B(n46411), .Z(n46403) );
  XNOR U46419 ( .A(n46399), .B(n46398), .Z(n46411) );
  XNOR U46420 ( .A(n46451), .B(n46395), .Z(n46398) );
  XNOR U46421 ( .A(p_input[1611]), .B(p_input[2059]), .Z(n46395) );
  XOR U46422 ( .A(p_input[1612]), .B(n28329), .Z(n46451) );
  XOR U46423 ( .A(p_input[1613]), .B(p_input[2061]), .Z(n46399) );
  XOR U46424 ( .A(n46409), .B(n46452), .Z(n46450) );
  IV U46425 ( .A(n46400), .Z(n46452) );
  XOR U46426 ( .A(p_input[1602]), .B(p_input[2050]), .Z(n46400) );
  XNOR U46427 ( .A(n46453), .B(n46416), .Z(n46409) );
  XNOR U46428 ( .A(p_input[1616]), .B(n28332), .Z(n46416) );
  XOR U46429 ( .A(n46406), .B(n46415), .Z(n46453) );
  XOR U46430 ( .A(n46454), .B(n46412), .Z(n46415) );
  XOR U46431 ( .A(p_input[1614]), .B(p_input[2062]), .Z(n46412) );
  XOR U46432 ( .A(p_input[1615]), .B(n28334), .Z(n46454) );
  XOR U46433 ( .A(p_input[1610]), .B(p_input[2058]), .Z(n46406) );
  XOR U46434 ( .A(n46423), .B(n46421), .Z(n46404) );
  XNOR U46435 ( .A(n46455), .B(n46428), .Z(n46421) );
  XOR U46436 ( .A(p_input[1609]), .B(p_input[2057]), .Z(n46428) );
  XOR U46437 ( .A(n46418), .B(n46427), .Z(n46455) );
  XOR U46438 ( .A(n46456), .B(n46424), .Z(n46427) );
  XOR U46439 ( .A(p_input[1607]), .B(p_input[2055]), .Z(n46424) );
  XOR U46440 ( .A(p_input[1608]), .B(n29427), .Z(n46456) );
  XOR U46441 ( .A(p_input[1603]), .B(p_input[2051]), .Z(n46418) );
  XNOR U46442 ( .A(n46433), .B(n46432), .Z(n46423) );
  XOR U46443 ( .A(n46457), .B(n46429), .Z(n46432) );
  XOR U46444 ( .A(p_input[1604]), .B(p_input[2052]), .Z(n46429) );
  XOR U46445 ( .A(p_input[1605]), .B(n29429), .Z(n46457) );
  XOR U46446 ( .A(p_input[1606]), .B(p_input[2054]), .Z(n46433) );
  XNOR U46447 ( .A(n46458), .B(n46459), .Z(n46234) );
  AND U46448 ( .A(n1085), .B(n46460), .Z(n46459) );
  XNOR U46449 ( .A(n46461), .B(n46462), .Z(n1085) );
  AND U46450 ( .A(n46463), .B(n46464), .Z(n46462) );
  XOR U46451 ( .A(n46248), .B(n46461), .Z(n46464) );
  XNOR U46452 ( .A(n46465), .B(n46461), .Z(n46463) );
  XOR U46453 ( .A(n46466), .B(n46467), .Z(n46461) );
  AND U46454 ( .A(n46468), .B(n46469), .Z(n46467) );
  XOR U46455 ( .A(n46263), .B(n46466), .Z(n46469) );
  XOR U46456 ( .A(n46466), .B(n46264), .Z(n46468) );
  XOR U46457 ( .A(n46470), .B(n46471), .Z(n46466) );
  AND U46458 ( .A(n46472), .B(n46473), .Z(n46471) );
  XOR U46459 ( .A(n46291), .B(n46470), .Z(n46473) );
  XOR U46460 ( .A(n46470), .B(n46292), .Z(n46472) );
  XOR U46461 ( .A(n46474), .B(n46475), .Z(n46470) );
  AND U46462 ( .A(n46476), .B(n46477), .Z(n46475) );
  XOR U46463 ( .A(n46340), .B(n46474), .Z(n46477) );
  XOR U46464 ( .A(n46474), .B(n46341), .Z(n46476) );
  XOR U46465 ( .A(n46478), .B(n46479), .Z(n46474) );
  AND U46466 ( .A(n46480), .B(n46481), .Z(n46479) );
  XOR U46467 ( .A(n46478), .B(n46437), .Z(n46481) );
  XNOR U46468 ( .A(n46482), .B(n46483), .Z(n46184) );
  AND U46469 ( .A(n1089), .B(n46484), .Z(n46483) );
  XNOR U46470 ( .A(n46485), .B(n46486), .Z(n1089) );
  AND U46471 ( .A(n46487), .B(n46488), .Z(n46486) );
  XOR U46472 ( .A(n46485), .B(n46194), .Z(n46488) );
  XNOR U46473 ( .A(n46485), .B(n46144), .Z(n46487) );
  XOR U46474 ( .A(n46489), .B(n46490), .Z(n46485) );
  AND U46475 ( .A(n46491), .B(n46492), .Z(n46490) );
  XNOR U46476 ( .A(n46204), .B(n46489), .Z(n46492) );
  XOR U46477 ( .A(n46489), .B(n46154), .Z(n46491) );
  XOR U46478 ( .A(n46493), .B(n46494), .Z(n46489) );
  AND U46479 ( .A(n46495), .B(n46496), .Z(n46494) );
  XNOR U46480 ( .A(n46214), .B(n46493), .Z(n46496) );
  XOR U46481 ( .A(n46493), .B(n46163), .Z(n46495) );
  XOR U46482 ( .A(n46497), .B(n46498), .Z(n46493) );
  AND U46483 ( .A(n46499), .B(n46500), .Z(n46498) );
  XOR U46484 ( .A(n46497), .B(n46171), .Z(n46499) );
  XOR U46485 ( .A(n46501), .B(n46502), .Z(n46135) );
  AND U46486 ( .A(n1093), .B(n46484), .Z(n46502) );
  XNOR U46487 ( .A(n46482), .B(n46501), .Z(n46484) );
  XNOR U46488 ( .A(n46503), .B(n46504), .Z(n1093) );
  AND U46489 ( .A(n46505), .B(n46506), .Z(n46504) );
  XNOR U46490 ( .A(n46507), .B(n46503), .Z(n46506) );
  IV U46491 ( .A(n46194), .Z(n46507) );
  XOR U46492 ( .A(n46465), .B(n46508), .Z(n46194) );
  AND U46493 ( .A(n1096), .B(n46509), .Z(n46508) );
  XOR U46494 ( .A(n46247), .B(n46244), .Z(n46509) );
  IV U46495 ( .A(n46465), .Z(n46247) );
  XNOR U46496 ( .A(n46144), .B(n46503), .Z(n46505) );
  XOR U46497 ( .A(n46510), .B(n46511), .Z(n46144) );
  AND U46498 ( .A(n1112), .B(n46512), .Z(n46511) );
  XOR U46499 ( .A(n46513), .B(n46514), .Z(n46503) );
  AND U46500 ( .A(n46515), .B(n46516), .Z(n46514) );
  XNOR U46501 ( .A(n46513), .B(n46204), .Z(n46516) );
  XOR U46502 ( .A(n46264), .B(n46517), .Z(n46204) );
  AND U46503 ( .A(n1096), .B(n46518), .Z(n46517) );
  XOR U46504 ( .A(n46260), .B(n46264), .Z(n46518) );
  XNOR U46505 ( .A(n46519), .B(n46513), .Z(n46515) );
  IV U46506 ( .A(n46154), .Z(n46519) );
  XOR U46507 ( .A(n46520), .B(n46521), .Z(n46154) );
  AND U46508 ( .A(n1112), .B(n46522), .Z(n46521) );
  XOR U46509 ( .A(n46523), .B(n46524), .Z(n46513) );
  AND U46510 ( .A(n46525), .B(n46526), .Z(n46524) );
  XNOR U46511 ( .A(n46523), .B(n46214), .Z(n46526) );
  XOR U46512 ( .A(n46292), .B(n46527), .Z(n46214) );
  AND U46513 ( .A(n1096), .B(n46528), .Z(n46527) );
  XOR U46514 ( .A(n46288), .B(n46292), .Z(n46528) );
  XOR U46515 ( .A(n46163), .B(n46523), .Z(n46525) );
  XOR U46516 ( .A(n46529), .B(n46530), .Z(n46163) );
  AND U46517 ( .A(n1112), .B(n46531), .Z(n46530) );
  XOR U46518 ( .A(n46497), .B(n46532), .Z(n46523) );
  AND U46519 ( .A(n46533), .B(n46500), .Z(n46532) );
  XNOR U46520 ( .A(n46224), .B(n46497), .Z(n46500) );
  XOR U46521 ( .A(n46341), .B(n46534), .Z(n46224) );
  AND U46522 ( .A(n1096), .B(n46535), .Z(n46534) );
  XOR U46523 ( .A(n46337), .B(n46341), .Z(n46535) );
  XNOR U46524 ( .A(n46536), .B(n46497), .Z(n46533) );
  IV U46525 ( .A(n46171), .Z(n46536) );
  XOR U46526 ( .A(n46537), .B(n46538), .Z(n46171) );
  AND U46527 ( .A(n1112), .B(n46539), .Z(n46538) );
  XOR U46528 ( .A(n46540), .B(n46541), .Z(n46497) );
  AND U46529 ( .A(n46542), .B(n46543), .Z(n46541) );
  XNOR U46530 ( .A(n46540), .B(n46232), .Z(n46543) );
  XOR U46531 ( .A(n46438), .B(n46544), .Z(n46232) );
  AND U46532 ( .A(n1096), .B(n46545), .Z(n46544) );
  XOR U46533 ( .A(n46434), .B(n46438), .Z(n46545) );
  XNOR U46534 ( .A(n46546), .B(n46540), .Z(n46542) );
  IV U46535 ( .A(n46181), .Z(n46546) );
  XOR U46536 ( .A(n46547), .B(n46548), .Z(n46181) );
  AND U46537 ( .A(n1112), .B(n46549), .Z(n46548) );
  AND U46538 ( .A(n46501), .B(n46482), .Z(n46540) );
  XNOR U46539 ( .A(n46550), .B(n46551), .Z(n46482) );
  AND U46540 ( .A(n1096), .B(n46460), .Z(n46551) );
  XNOR U46541 ( .A(n46458), .B(n46550), .Z(n46460) );
  XNOR U46542 ( .A(n46552), .B(n46553), .Z(n1096) );
  AND U46543 ( .A(n46554), .B(n46555), .Z(n46553) );
  XNOR U46544 ( .A(n46552), .B(n46244), .Z(n46555) );
  IV U46545 ( .A(n46248), .Z(n46244) );
  XOR U46546 ( .A(n46556), .B(n46557), .Z(n46248) );
  AND U46547 ( .A(n1100), .B(n46558), .Z(n46557) );
  XOR U46548 ( .A(n46559), .B(n46556), .Z(n46558) );
  XNOR U46549 ( .A(n46552), .B(n46465), .Z(n46554) );
  XOR U46550 ( .A(n46560), .B(n46561), .Z(n46465) );
  AND U46551 ( .A(n1108), .B(n46512), .Z(n46561) );
  XOR U46552 ( .A(n46510), .B(n46560), .Z(n46512) );
  XOR U46553 ( .A(n46562), .B(n46563), .Z(n46552) );
  AND U46554 ( .A(n46564), .B(n46565), .Z(n46563) );
  XNOR U46555 ( .A(n46562), .B(n46260), .Z(n46565) );
  IV U46556 ( .A(n46263), .Z(n46260) );
  XOR U46557 ( .A(n46566), .B(n46567), .Z(n46263) );
  AND U46558 ( .A(n1100), .B(n46568), .Z(n46567) );
  XOR U46559 ( .A(n46569), .B(n46566), .Z(n46568) );
  XOR U46560 ( .A(n46264), .B(n46562), .Z(n46564) );
  XOR U46561 ( .A(n46570), .B(n46571), .Z(n46264) );
  AND U46562 ( .A(n1108), .B(n46522), .Z(n46571) );
  XOR U46563 ( .A(n46570), .B(n46520), .Z(n46522) );
  XOR U46564 ( .A(n46572), .B(n46573), .Z(n46562) );
  AND U46565 ( .A(n46574), .B(n46575), .Z(n46573) );
  XNOR U46566 ( .A(n46572), .B(n46288), .Z(n46575) );
  IV U46567 ( .A(n46291), .Z(n46288) );
  XOR U46568 ( .A(n46576), .B(n46577), .Z(n46291) );
  AND U46569 ( .A(n1100), .B(n46578), .Z(n46577) );
  XNOR U46570 ( .A(n46579), .B(n46576), .Z(n46578) );
  XOR U46571 ( .A(n46292), .B(n46572), .Z(n46574) );
  XOR U46572 ( .A(n46580), .B(n46581), .Z(n46292) );
  AND U46573 ( .A(n1108), .B(n46531), .Z(n46581) );
  XOR U46574 ( .A(n46580), .B(n46529), .Z(n46531) );
  XOR U46575 ( .A(n46582), .B(n46583), .Z(n46572) );
  AND U46576 ( .A(n46584), .B(n46585), .Z(n46583) );
  XNOR U46577 ( .A(n46582), .B(n46337), .Z(n46585) );
  IV U46578 ( .A(n46340), .Z(n46337) );
  XOR U46579 ( .A(n46586), .B(n46587), .Z(n46340) );
  AND U46580 ( .A(n1100), .B(n46588), .Z(n46587) );
  XOR U46581 ( .A(n46589), .B(n46586), .Z(n46588) );
  XOR U46582 ( .A(n46341), .B(n46582), .Z(n46584) );
  XOR U46583 ( .A(n46590), .B(n46591), .Z(n46341) );
  AND U46584 ( .A(n1108), .B(n46539), .Z(n46591) );
  XOR U46585 ( .A(n46590), .B(n46537), .Z(n46539) );
  XOR U46586 ( .A(n46478), .B(n46592), .Z(n46582) );
  AND U46587 ( .A(n46480), .B(n46593), .Z(n46592) );
  XNOR U46588 ( .A(n46478), .B(n46434), .Z(n46593) );
  IV U46589 ( .A(n46437), .Z(n46434) );
  XOR U46590 ( .A(n46594), .B(n46595), .Z(n46437) );
  AND U46591 ( .A(n1100), .B(n46596), .Z(n46595) );
  XNOR U46592 ( .A(n46597), .B(n46594), .Z(n46596) );
  XOR U46593 ( .A(n46438), .B(n46478), .Z(n46480) );
  XOR U46594 ( .A(n46598), .B(n46599), .Z(n46438) );
  AND U46595 ( .A(n1108), .B(n46549), .Z(n46599) );
  XOR U46596 ( .A(n46598), .B(n46547), .Z(n46549) );
  AND U46597 ( .A(n46550), .B(n46458), .Z(n46478) );
  XNOR U46598 ( .A(n46600), .B(n46601), .Z(n46458) );
  AND U46599 ( .A(n1100), .B(n46602), .Z(n46601) );
  XNOR U46600 ( .A(n46603), .B(n46600), .Z(n46602) );
  XNOR U46601 ( .A(n46604), .B(n46605), .Z(n1100) );
  AND U46602 ( .A(n46606), .B(n46607), .Z(n46605) );
  XOR U46603 ( .A(n46559), .B(n46604), .Z(n46607) );
  AND U46604 ( .A(n46608), .B(n46609), .Z(n46559) );
  XNOR U46605 ( .A(n46556), .B(n46604), .Z(n46606) );
  XNOR U46606 ( .A(n46610), .B(n46611), .Z(n46556) );
  AND U46607 ( .A(n1104), .B(n46612), .Z(n46611) );
  XNOR U46608 ( .A(n46613), .B(n46614), .Z(n46612) );
  XOR U46609 ( .A(n46615), .B(n46616), .Z(n46604) );
  AND U46610 ( .A(n46617), .B(n46618), .Z(n46616) );
  XNOR U46611 ( .A(n46615), .B(n46608), .Z(n46618) );
  IV U46612 ( .A(n46569), .Z(n46608) );
  XOR U46613 ( .A(n46619), .B(n46620), .Z(n46569) );
  XOR U46614 ( .A(n46621), .B(n46609), .Z(n46620) );
  AND U46615 ( .A(n46579), .B(n46622), .Z(n46609) );
  AND U46616 ( .A(n46623), .B(n46624), .Z(n46621) );
  XOR U46617 ( .A(n46625), .B(n46619), .Z(n46623) );
  XNOR U46618 ( .A(n46566), .B(n46615), .Z(n46617) );
  XNOR U46619 ( .A(n46626), .B(n46627), .Z(n46566) );
  AND U46620 ( .A(n1104), .B(n46628), .Z(n46627) );
  XNOR U46621 ( .A(n46629), .B(n46630), .Z(n46628) );
  XOR U46622 ( .A(n46631), .B(n46632), .Z(n46615) );
  AND U46623 ( .A(n46633), .B(n46634), .Z(n46632) );
  XNOR U46624 ( .A(n46631), .B(n46579), .Z(n46634) );
  XOR U46625 ( .A(n46635), .B(n46624), .Z(n46579) );
  XNOR U46626 ( .A(n46636), .B(n46619), .Z(n46624) );
  XOR U46627 ( .A(n46637), .B(n46638), .Z(n46619) );
  AND U46628 ( .A(n46639), .B(n46640), .Z(n46638) );
  XOR U46629 ( .A(n46641), .B(n46637), .Z(n46639) );
  XNOR U46630 ( .A(n46642), .B(n46643), .Z(n46636) );
  AND U46631 ( .A(n46644), .B(n46645), .Z(n46643) );
  XOR U46632 ( .A(n46642), .B(n46646), .Z(n46644) );
  XNOR U46633 ( .A(n46625), .B(n46622), .Z(n46635) );
  AND U46634 ( .A(n46647), .B(n46648), .Z(n46622) );
  XOR U46635 ( .A(n46649), .B(n46650), .Z(n46625) );
  AND U46636 ( .A(n46651), .B(n46652), .Z(n46650) );
  XOR U46637 ( .A(n46649), .B(n46653), .Z(n46651) );
  XNOR U46638 ( .A(n46576), .B(n46631), .Z(n46633) );
  XNOR U46639 ( .A(n46654), .B(n46655), .Z(n46576) );
  AND U46640 ( .A(n1104), .B(n46656), .Z(n46655) );
  XNOR U46641 ( .A(n46657), .B(n46658), .Z(n46656) );
  XOR U46642 ( .A(n46659), .B(n46660), .Z(n46631) );
  AND U46643 ( .A(n46661), .B(n46662), .Z(n46660) );
  XNOR U46644 ( .A(n46659), .B(n46647), .Z(n46662) );
  IV U46645 ( .A(n46589), .Z(n46647) );
  XNOR U46646 ( .A(n46663), .B(n46640), .Z(n46589) );
  XNOR U46647 ( .A(n46664), .B(n46646), .Z(n46640) );
  XOR U46648 ( .A(n46665), .B(n46666), .Z(n46646) );
  AND U46649 ( .A(n46667), .B(n46668), .Z(n46666) );
  XOR U46650 ( .A(n46665), .B(n46669), .Z(n46667) );
  XNOR U46651 ( .A(n46645), .B(n46637), .Z(n46664) );
  XOR U46652 ( .A(n46670), .B(n46671), .Z(n46637) );
  AND U46653 ( .A(n46672), .B(n46673), .Z(n46671) );
  XNOR U46654 ( .A(n46674), .B(n46670), .Z(n46672) );
  XNOR U46655 ( .A(n46675), .B(n46642), .Z(n46645) );
  XOR U46656 ( .A(n46676), .B(n46677), .Z(n46642) );
  AND U46657 ( .A(n46678), .B(n46679), .Z(n46677) );
  XOR U46658 ( .A(n46676), .B(n46680), .Z(n46678) );
  XNOR U46659 ( .A(n46681), .B(n46682), .Z(n46675) );
  AND U46660 ( .A(n46683), .B(n46684), .Z(n46682) );
  XNOR U46661 ( .A(n46681), .B(n46685), .Z(n46683) );
  XNOR U46662 ( .A(n46641), .B(n46648), .Z(n46663) );
  AND U46663 ( .A(n46597), .B(n46686), .Z(n46648) );
  XOR U46664 ( .A(n46653), .B(n46652), .Z(n46641) );
  XNOR U46665 ( .A(n46687), .B(n46649), .Z(n46652) );
  XOR U46666 ( .A(n46688), .B(n46689), .Z(n46649) );
  AND U46667 ( .A(n46690), .B(n46691), .Z(n46689) );
  XOR U46668 ( .A(n46688), .B(n46692), .Z(n46690) );
  XNOR U46669 ( .A(n46693), .B(n46694), .Z(n46687) );
  AND U46670 ( .A(n46695), .B(n46696), .Z(n46694) );
  XOR U46671 ( .A(n46693), .B(n46697), .Z(n46695) );
  XOR U46672 ( .A(n46698), .B(n46699), .Z(n46653) );
  AND U46673 ( .A(n46700), .B(n46701), .Z(n46699) );
  XOR U46674 ( .A(n46698), .B(n46702), .Z(n46700) );
  XNOR U46675 ( .A(n46586), .B(n46659), .Z(n46661) );
  XNOR U46676 ( .A(n46703), .B(n46704), .Z(n46586) );
  AND U46677 ( .A(n1104), .B(n46705), .Z(n46704) );
  XNOR U46678 ( .A(n46706), .B(n46707), .Z(n46705) );
  XOR U46679 ( .A(n46708), .B(n46709), .Z(n46659) );
  AND U46680 ( .A(n46710), .B(n46711), .Z(n46709) );
  XNOR U46681 ( .A(n46708), .B(n46597), .Z(n46711) );
  XOR U46682 ( .A(n46712), .B(n46673), .Z(n46597) );
  XNOR U46683 ( .A(n46713), .B(n46680), .Z(n46673) );
  XOR U46684 ( .A(n46669), .B(n46668), .Z(n46680) );
  XNOR U46685 ( .A(n46714), .B(n46665), .Z(n46668) );
  XOR U46686 ( .A(n46715), .B(n46716), .Z(n46665) );
  AND U46687 ( .A(n46717), .B(n46718), .Z(n46716) );
  XNOR U46688 ( .A(n46719), .B(n46720), .Z(n46717) );
  IV U46689 ( .A(n46715), .Z(n46719) );
  XNOR U46690 ( .A(n46721), .B(n46722), .Z(n46714) );
  NOR U46691 ( .A(n46723), .B(n46724), .Z(n46722) );
  XNOR U46692 ( .A(n46721), .B(n46725), .Z(n46723) );
  XOR U46693 ( .A(n46726), .B(n46727), .Z(n46669) );
  NOR U46694 ( .A(n46728), .B(n46729), .Z(n46727) );
  XNOR U46695 ( .A(n46726), .B(n46730), .Z(n46728) );
  XNOR U46696 ( .A(n46679), .B(n46670), .Z(n46713) );
  XOR U46697 ( .A(n46731), .B(n46732), .Z(n46670) );
  AND U46698 ( .A(n46733), .B(n46734), .Z(n46732) );
  XOR U46699 ( .A(n46731), .B(n46735), .Z(n46733) );
  XOR U46700 ( .A(n46736), .B(n46685), .Z(n46679) );
  XOR U46701 ( .A(n46737), .B(n46738), .Z(n46685) );
  NOR U46702 ( .A(n46739), .B(n46740), .Z(n46738) );
  XOR U46703 ( .A(n46737), .B(n46741), .Z(n46739) );
  XNOR U46704 ( .A(n46684), .B(n46676), .Z(n46736) );
  XOR U46705 ( .A(n46742), .B(n46743), .Z(n46676) );
  AND U46706 ( .A(n46744), .B(n46745), .Z(n46743) );
  XOR U46707 ( .A(n46742), .B(n46746), .Z(n46744) );
  XNOR U46708 ( .A(n46747), .B(n46681), .Z(n46684) );
  XOR U46709 ( .A(n46748), .B(n46749), .Z(n46681) );
  AND U46710 ( .A(n46750), .B(n46751), .Z(n46749) );
  XNOR U46711 ( .A(n46752), .B(n46753), .Z(n46750) );
  IV U46712 ( .A(n46748), .Z(n46752) );
  XNOR U46713 ( .A(n46754), .B(n46755), .Z(n46747) );
  NOR U46714 ( .A(n46756), .B(n46757), .Z(n46755) );
  XNOR U46715 ( .A(n46754), .B(n46758), .Z(n46756) );
  XOR U46716 ( .A(n46674), .B(n46686), .Z(n46712) );
  NOR U46717 ( .A(n46603), .B(n46759), .Z(n46686) );
  XNOR U46718 ( .A(n46692), .B(n46691), .Z(n46674) );
  XNOR U46719 ( .A(n46760), .B(n46697), .Z(n46691) );
  XNOR U46720 ( .A(n46761), .B(n46762), .Z(n46697) );
  NOR U46721 ( .A(n46763), .B(n46764), .Z(n46762) );
  XOR U46722 ( .A(n46761), .B(n46765), .Z(n46763) );
  XNOR U46723 ( .A(n46696), .B(n46688), .Z(n46760) );
  XOR U46724 ( .A(n46766), .B(n46767), .Z(n46688) );
  AND U46725 ( .A(n46768), .B(n46769), .Z(n46767) );
  XOR U46726 ( .A(n46766), .B(n46770), .Z(n46768) );
  XNOR U46727 ( .A(n46771), .B(n46693), .Z(n46696) );
  XOR U46728 ( .A(n46772), .B(n46773), .Z(n46693) );
  AND U46729 ( .A(n46774), .B(n46775), .Z(n46773) );
  XNOR U46730 ( .A(n46776), .B(n46777), .Z(n46774) );
  IV U46731 ( .A(n46772), .Z(n46776) );
  XNOR U46732 ( .A(n46778), .B(n46779), .Z(n46771) );
  NOR U46733 ( .A(n46780), .B(n46781), .Z(n46779) );
  XNOR U46734 ( .A(n46778), .B(n46782), .Z(n46780) );
  XOR U46735 ( .A(n46702), .B(n46701), .Z(n46692) );
  XNOR U46736 ( .A(n46783), .B(n46698), .Z(n46701) );
  XOR U46737 ( .A(n46784), .B(n46785), .Z(n46698) );
  AND U46738 ( .A(n46786), .B(n46787), .Z(n46785) );
  XNOR U46739 ( .A(n46788), .B(n46789), .Z(n46786) );
  IV U46740 ( .A(n46784), .Z(n46788) );
  XNOR U46741 ( .A(n46790), .B(n46791), .Z(n46783) );
  NOR U46742 ( .A(n46792), .B(n46793), .Z(n46791) );
  XNOR U46743 ( .A(n46790), .B(n46794), .Z(n46792) );
  XOR U46744 ( .A(n46795), .B(n46796), .Z(n46702) );
  NOR U46745 ( .A(n46797), .B(n46798), .Z(n46796) );
  XNOR U46746 ( .A(n46795), .B(n46799), .Z(n46797) );
  XNOR U46747 ( .A(n46594), .B(n46708), .Z(n46710) );
  XNOR U46748 ( .A(n46800), .B(n46801), .Z(n46594) );
  AND U46749 ( .A(n1104), .B(n46802), .Z(n46801) );
  XNOR U46750 ( .A(n46803), .B(n46804), .Z(n46802) );
  AND U46751 ( .A(n46600), .B(n46603), .Z(n46708) );
  XOR U46752 ( .A(n46805), .B(n46759), .Z(n46603) );
  XNOR U46753 ( .A(p_input[1632]), .B(p_input[2048]), .Z(n46759) );
  XNOR U46754 ( .A(n46735), .B(n46734), .Z(n46805) );
  XNOR U46755 ( .A(n46806), .B(n46746), .Z(n46734) );
  XOR U46756 ( .A(n46720), .B(n46718), .Z(n46746) );
  XNOR U46757 ( .A(n46807), .B(n46725), .Z(n46718) );
  XOR U46758 ( .A(p_input[1656]), .B(p_input[2072]), .Z(n46725) );
  XOR U46759 ( .A(n46715), .B(n46724), .Z(n46807) );
  XOR U46760 ( .A(n46808), .B(n46721), .Z(n46724) );
  XOR U46761 ( .A(p_input[1654]), .B(p_input[2070]), .Z(n46721) );
  XOR U46762 ( .A(p_input[1655]), .B(n29410), .Z(n46808) );
  XOR U46763 ( .A(p_input[1650]), .B(p_input[2066]), .Z(n46715) );
  XNOR U46764 ( .A(n46730), .B(n46729), .Z(n46720) );
  XOR U46765 ( .A(n46809), .B(n46726), .Z(n46729) );
  XOR U46766 ( .A(p_input[1651]), .B(p_input[2067]), .Z(n46726) );
  XOR U46767 ( .A(p_input[1652]), .B(n29412), .Z(n46809) );
  XOR U46768 ( .A(p_input[1653]), .B(p_input[2069]), .Z(n46730) );
  XOR U46769 ( .A(n46745), .B(n46810), .Z(n46806) );
  IV U46770 ( .A(n46731), .Z(n46810) );
  XOR U46771 ( .A(p_input[1633]), .B(p_input[2049]), .Z(n46731) );
  XNOR U46772 ( .A(n46811), .B(n46753), .Z(n46745) );
  XNOR U46773 ( .A(n46741), .B(n46740), .Z(n46753) );
  XNOR U46774 ( .A(n46812), .B(n46737), .Z(n46740) );
  XNOR U46775 ( .A(p_input[1658]), .B(p_input[2074]), .Z(n46737) );
  XOR U46776 ( .A(p_input[1659]), .B(n29415), .Z(n46812) );
  XOR U46777 ( .A(p_input[1660]), .B(p_input[2076]), .Z(n46741) );
  XOR U46778 ( .A(n46751), .B(n46813), .Z(n46811) );
  IV U46779 ( .A(n46742), .Z(n46813) );
  XOR U46780 ( .A(p_input[1649]), .B(p_input[2065]), .Z(n46742) );
  XNOR U46781 ( .A(n46814), .B(n46758), .Z(n46751) );
  XNOR U46782 ( .A(p_input[1663]), .B(n29418), .Z(n46758) );
  XOR U46783 ( .A(n46748), .B(n46757), .Z(n46814) );
  XOR U46784 ( .A(n46815), .B(n46754), .Z(n46757) );
  XOR U46785 ( .A(p_input[1661]), .B(p_input[2077]), .Z(n46754) );
  XOR U46786 ( .A(p_input[1662]), .B(n29420), .Z(n46815) );
  XOR U46787 ( .A(p_input[1657]), .B(p_input[2073]), .Z(n46748) );
  XOR U46788 ( .A(n46770), .B(n46769), .Z(n46735) );
  XNOR U46789 ( .A(n46816), .B(n46777), .Z(n46769) );
  XNOR U46790 ( .A(n46765), .B(n46764), .Z(n46777) );
  XNOR U46791 ( .A(n46817), .B(n46761), .Z(n46764) );
  XNOR U46792 ( .A(p_input[1643]), .B(p_input[2059]), .Z(n46761) );
  XOR U46793 ( .A(p_input[1644]), .B(n28329), .Z(n46817) );
  XOR U46794 ( .A(p_input[1645]), .B(p_input[2061]), .Z(n46765) );
  XOR U46795 ( .A(n46775), .B(n46818), .Z(n46816) );
  IV U46796 ( .A(n46766), .Z(n46818) );
  XOR U46797 ( .A(p_input[1634]), .B(p_input[2050]), .Z(n46766) );
  XNOR U46798 ( .A(n46819), .B(n46782), .Z(n46775) );
  XNOR U46799 ( .A(p_input[1648]), .B(n28332), .Z(n46782) );
  XOR U46800 ( .A(n46772), .B(n46781), .Z(n46819) );
  XOR U46801 ( .A(n46820), .B(n46778), .Z(n46781) );
  XOR U46802 ( .A(p_input[1646]), .B(p_input[2062]), .Z(n46778) );
  XOR U46803 ( .A(p_input[1647]), .B(n28334), .Z(n46820) );
  XOR U46804 ( .A(p_input[1642]), .B(p_input[2058]), .Z(n46772) );
  XOR U46805 ( .A(n46789), .B(n46787), .Z(n46770) );
  XNOR U46806 ( .A(n46821), .B(n46794), .Z(n46787) );
  XOR U46807 ( .A(p_input[1641]), .B(p_input[2057]), .Z(n46794) );
  XOR U46808 ( .A(n46784), .B(n46793), .Z(n46821) );
  XOR U46809 ( .A(n46822), .B(n46790), .Z(n46793) );
  XOR U46810 ( .A(p_input[1639]), .B(p_input[2055]), .Z(n46790) );
  XOR U46811 ( .A(p_input[1640]), .B(n29427), .Z(n46822) );
  XOR U46812 ( .A(p_input[1635]), .B(p_input[2051]), .Z(n46784) );
  XNOR U46813 ( .A(n46799), .B(n46798), .Z(n46789) );
  XOR U46814 ( .A(n46823), .B(n46795), .Z(n46798) );
  XOR U46815 ( .A(p_input[1636]), .B(p_input[2052]), .Z(n46795) );
  XOR U46816 ( .A(p_input[1637]), .B(n29429), .Z(n46823) );
  XOR U46817 ( .A(p_input[1638]), .B(p_input[2054]), .Z(n46799) );
  XNOR U46818 ( .A(n46824), .B(n46825), .Z(n46600) );
  AND U46819 ( .A(n1104), .B(n46826), .Z(n46825) );
  XNOR U46820 ( .A(n46827), .B(n46828), .Z(n1104) );
  AND U46821 ( .A(n46829), .B(n46830), .Z(n46828) );
  XOR U46822 ( .A(n46614), .B(n46827), .Z(n46830) );
  XNOR U46823 ( .A(n46831), .B(n46827), .Z(n46829) );
  XOR U46824 ( .A(n46832), .B(n46833), .Z(n46827) );
  AND U46825 ( .A(n46834), .B(n46835), .Z(n46833) );
  XOR U46826 ( .A(n46629), .B(n46832), .Z(n46835) );
  XOR U46827 ( .A(n46832), .B(n46630), .Z(n46834) );
  XOR U46828 ( .A(n46836), .B(n46837), .Z(n46832) );
  AND U46829 ( .A(n46838), .B(n46839), .Z(n46837) );
  XOR U46830 ( .A(n46657), .B(n46836), .Z(n46839) );
  XOR U46831 ( .A(n46836), .B(n46658), .Z(n46838) );
  XOR U46832 ( .A(n46840), .B(n46841), .Z(n46836) );
  AND U46833 ( .A(n46842), .B(n46843), .Z(n46841) );
  XOR U46834 ( .A(n46706), .B(n46840), .Z(n46843) );
  XOR U46835 ( .A(n46840), .B(n46707), .Z(n46842) );
  XOR U46836 ( .A(n46844), .B(n46845), .Z(n46840) );
  AND U46837 ( .A(n46846), .B(n46847), .Z(n46845) );
  XOR U46838 ( .A(n46844), .B(n46803), .Z(n46847) );
  XNOR U46839 ( .A(n46848), .B(n46849), .Z(n46550) );
  AND U46840 ( .A(n1108), .B(n46850), .Z(n46849) );
  XNOR U46841 ( .A(n46851), .B(n46852), .Z(n1108) );
  AND U46842 ( .A(n46853), .B(n46854), .Z(n46852) );
  XOR U46843 ( .A(n46851), .B(n46560), .Z(n46854) );
  XNOR U46844 ( .A(n46851), .B(n46510), .Z(n46853) );
  XOR U46845 ( .A(n46855), .B(n46856), .Z(n46851) );
  AND U46846 ( .A(n46857), .B(n46858), .Z(n46856) );
  XNOR U46847 ( .A(n46570), .B(n46855), .Z(n46858) );
  XOR U46848 ( .A(n46855), .B(n46520), .Z(n46857) );
  XOR U46849 ( .A(n46859), .B(n46860), .Z(n46855) );
  AND U46850 ( .A(n46861), .B(n46862), .Z(n46860) );
  XNOR U46851 ( .A(n46580), .B(n46859), .Z(n46862) );
  XOR U46852 ( .A(n46859), .B(n46529), .Z(n46861) );
  XOR U46853 ( .A(n46863), .B(n46864), .Z(n46859) );
  AND U46854 ( .A(n46865), .B(n46866), .Z(n46864) );
  XOR U46855 ( .A(n46863), .B(n46537), .Z(n46865) );
  XOR U46856 ( .A(n46867), .B(n46868), .Z(n46501) );
  AND U46857 ( .A(n1112), .B(n46850), .Z(n46868) );
  XNOR U46858 ( .A(n46848), .B(n46867), .Z(n46850) );
  XNOR U46859 ( .A(n46869), .B(n46870), .Z(n1112) );
  AND U46860 ( .A(n46871), .B(n46872), .Z(n46870) );
  XNOR U46861 ( .A(n46873), .B(n46869), .Z(n46872) );
  IV U46862 ( .A(n46560), .Z(n46873) );
  XOR U46863 ( .A(n46831), .B(n46874), .Z(n46560) );
  AND U46864 ( .A(n1115), .B(n46875), .Z(n46874) );
  XOR U46865 ( .A(n46613), .B(n46610), .Z(n46875) );
  IV U46866 ( .A(n46831), .Z(n46613) );
  XNOR U46867 ( .A(n46510), .B(n46869), .Z(n46871) );
  XOR U46868 ( .A(n46876), .B(n46877), .Z(n46510) );
  AND U46869 ( .A(n1131), .B(n46878), .Z(n46877) );
  XOR U46870 ( .A(n46879), .B(n46880), .Z(n46869) );
  AND U46871 ( .A(n46881), .B(n46882), .Z(n46880) );
  XNOR U46872 ( .A(n46879), .B(n46570), .Z(n46882) );
  XOR U46873 ( .A(n46630), .B(n46883), .Z(n46570) );
  AND U46874 ( .A(n1115), .B(n46884), .Z(n46883) );
  XOR U46875 ( .A(n46626), .B(n46630), .Z(n46884) );
  XNOR U46876 ( .A(n46885), .B(n46879), .Z(n46881) );
  IV U46877 ( .A(n46520), .Z(n46885) );
  XOR U46878 ( .A(n46886), .B(n46887), .Z(n46520) );
  AND U46879 ( .A(n1131), .B(n46888), .Z(n46887) );
  XOR U46880 ( .A(n46889), .B(n46890), .Z(n46879) );
  AND U46881 ( .A(n46891), .B(n46892), .Z(n46890) );
  XNOR U46882 ( .A(n46889), .B(n46580), .Z(n46892) );
  XOR U46883 ( .A(n46658), .B(n46893), .Z(n46580) );
  AND U46884 ( .A(n1115), .B(n46894), .Z(n46893) );
  XOR U46885 ( .A(n46654), .B(n46658), .Z(n46894) );
  XOR U46886 ( .A(n46529), .B(n46889), .Z(n46891) );
  XOR U46887 ( .A(n46895), .B(n46896), .Z(n46529) );
  AND U46888 ( .A(n1131), .B(n46897), .Z(n46896) );
  XOR U46889 ( .A(n46863), .B(n46898), .Z(n46889) );
  AND U46890 ( .A(n46899), .B(n46866), .Z(n46898) );
  XNOR U46891 ( .A(n46590), .B(n46863), .Z(n46866) );
  XOR U46892 ( .A(n46707), .B(n46900), .Z(n46590) );
  AND U46893 ( .A(n1115), .B(n46901), .Z(n46900) );
  XOR U46894 ( .A(n46703), .B(n46707), .Z(n46901) );
  XNOR U46895 ( .A(n46902), .B(n46863), .Z(n46899) );
  IV U46896 ( .A(n46537), .Z(n46902) );
  XOR U46897 ( .A(n46903), .B(n46904), .Z(n46537) );
  AND U46898 ( .A(n1131), .B(n46905), .Z(n46904) );
  XOR U46899 ( .A(n46906), .B(n46907), .Z(n46863) );
  AND U46900 ( .A(n46908), .B(n46909), .Z(n46907) );
  XNOR U46901 ( .A(n46906), .B(n46598), .Z(n46909) );
  XOR U46902 ( .A(n46804), .B(n46910), .Z(n46598) );
  AND U46903 ( .A(n1115), .B(n46911), .Z(n46910) );
  XOR U46904 ( .A(n46800), .B(n46804), .Z(n46911) );
  XNOR U46905 ( .A(n46912), .B(n46906), .Z(n46908) );
  IV U46906 ( .A(n46547), .Z(n46912) );
  XOR U46907 ( .A(n46913), .B(n46914), .Z(n46547) );
  AND U46908 ( .A(n1131), .B(n46915), .Z(n46914) );
  AND U46909 ( .A(n46867), .B(n46848), .Z(n46906) );
  XNOR U46910 ( .A(n46916), .B(n46917), .Z(n46848) );
  AND U46911 ( .A(n1115), .B(n46826), .Z(n46917) );
  XNOR U46912 ( .A(n46824), .B(n46916), .Z(n46826) );
  XNOR U46913 ( .A(n46918), .B(n46919), .Z(n1115) );
  AND U46914 ( .A(n46920), .B(n46921), .Z(n46919) );
  XNOR U46915 ( .A(n46918), .B(n46610), .Z(n46921) );
  IV U46916 ( .A(n46614), .Z(n46610) );
  XOR U46917 ( .A(n46922), .B(n46923), .Z(n46614) );
  AND U46918 ( .A(n1119), .B(n46924), .Z(n46923) );
  XOR U46919 ( .A(n46925), .B(n46922), .Z(n46924) );
  XNOR U46920 ( .A(n46918), .B(n46831), .Z(n46920) );
  XOR U46921 ( .A(n46926), .B(n46927), .Z(n46831) );
  AND U46922 ( .A(n1127), .B(n46878), .Z(n46927) );
  XOR U46923 ( .A(n46876), .B(n46926), .Z(n46878) );
  XOR U46924 ( .A(n46928), .B(n46929), .Z(n46918) );
  AND U46925 ( .A(n46930), .B(n46931), .Z(n46929) );
  XNOR U46926 ( .A(n46928), .B(n46626), .Z(n46931) );
  IV U46927 ( .A(n46629), .Z(n46626) );
  XOR U46928 ( .A(n46932), .B(n46933), .Z(n46629) );
  AND U46929 ( .A(n1119), .B(n46934), .Z(n46933) );
  XOR U46930 ( .A(n46935), .B(n46932), .Z(n46934) );
  XOR U46931 ( .A(n46630), .B(n46928), .Z(n46930) );
  XOR U46932 ( .A(n46936), .B(n46937), .Z(n46630) );
  AND U46933 ( .A(n1127), .B(n46888), .Z(n46937) );
  XOR U46934 ( .A(n46936), .B(n46886), .Z(n46888) );
  XOR U46935 ( .A(n46938), .B(n46939), .Z(n46928) );
  AND U46936 ( .A(n46940), .B(n46941), .Z(n46939) );
  XNOR U46937 ( .A(n46938), .B(n46654), .Z(n46941) );
  IV U46938 ( .A(n46657), .Z(n46654) );
  XOR U46939 ( .A(n46942), .B(n46943), .Z(n46657) );
  AND U46940 ( .A(n1119), .B(n46944), .Z(n46943) );
  XNOR U46941 ( .A(n46945), .B(n46942), .Z(n46944) );
  XOR U46942 ( .A(n46658), .B(n46938), .Z(n46940) );
  XOR U46943 ( .A(n46946), .B(n46947), .Z(n46658) );
  AND U46944 ( .A(n1127), .B(n46897), .Z(n46947) );
  XOR U46945 ( .A(n46946), .B(n46895), .Z(n46897) );
  XOR U46946 ( .A(n46948), .B(n46949), .Z(n46938) );
  AND U46947 ( .A(n46950), .B(n46951), .Z(n46949) );
  XNOR U46948 ( .A(n46948), .B(n46703), .Z(n46951) );
  IV U46949 ( .A(n46706), .Z(n46703) );
  XOR U46950 ( .A(n46952), .B(n46953), .Z(n46706) );
  AND U46951 ( .A(n1119), .B(n46954), .Z(n46953) );
  XOR U46952 ( .A(n46955), .B(n46952), .Z(n46954) );
  XOR U46953 ( .A(n46707), .B(n46948), .Z(n46950) );
  XOR U46954 ( .A(n46956), .B(n46957), .Z(n46707) );
  AND U46955 ( .A(n1127), .B(n46905), .Z(n46957) );
  XOR U46956 ( .A(n46956), .B(n46903), .Z(n46905) );
  XOR U46957 ( .A(n46844), .B(n46958), .Z(n46948) );
  AND U46958 ( .A(n46846), .B(n46959), .Z(n46958) );
  XNOR U46959 ( .A(n46844), .B(n46800), .Z(n46959) );
  IV U46960 ( .A(n46803), .Z(n46800) );
  XOR U46961 ( .A(n46960), .B(n46961), .Z(n46803) );
  AND U46962 ( .A(n1119), .B(n46962), .Z(n46961) );
  XNOR U46963 ( .A(n46963), .B(n46960), .Z(n46962) );
  XOR U46964 ( .A(n46804), .B(n46844), .Z(n46846) );
  XOR U46965 ( .A(n46964), .B(n46965), .Z(n46804) );
  AND U46966 ( .A(n1127), .B(n46915), .Z(n46965) );
  XOR U46967 ( .A(n46964), .B(n46913), .Z(n46915) );
  AND U46968 ( .A(n46916), .B(n46824), .Z(n46844) );
  XNOR U46969 ( .A(n46966), .B(n46967), .Z(n46824) );
  AND U46970 ( .A(n1119), .B(n46968), .Z(n46967) );
  XNOR U46971 ( .A(n46969), .B(n46966), .Z(n46968) );
  XNOR U46972 ( .A(n46970), .B(n46971), .Z(n1119) );
  AND U46973 ( .A(n46972), .B(n46973), .Z(n46971) );
  XOR U46974 ( .A(n46925), .B(n46970), .Z(n46973) );
  AND U46975 ( .A(n46974), .B(n46975), .Z(n46925) );
  XNOR U46976 ( .A(n46922), .B(n46970), .Z(n46972) );
  XNOR U46977 ( .A(n46976), .B(n46977), .Z(n46922) );
  AND U46978 ( .A(n1123), .B(n46978), .Z(n46977) );
  XNOR U46979 ( .A(n46979), .B(n46980), .Z(n46978) );
  XOR U46980 ( .A(n46981), .B(n46982), .Z(n46970) );
  AND U46981 ( .A(n46983), .B(n46984), .Z(n46982) );
  XNOR U46982 ( .A(n46981), .B(n46974), .Z(n46984) );
  IV U46983 ( .A(n46935), .Z(n46974) );
  XOR U46984 ( .A(n46985), .B(n46986), .Z(n46935) );
  XOR U46985 ( .A(n46987), .B(n46975), .Z(n46986) );
  AND U46986 ( .A(n46945), .B(n46988), .Z(n46975) );
  AND U46987 ( .A(n46989), .B(n46990), .Z(n46987) );
  XOR U46988 ( .A(n46991), .B(n46985), .Z(n46989) );
  XNOR U46989 ( .A(n46932), .B(n46981), .Z(n46983) );
  XNOR U46990 ( .A(n46992), .B(n46993), .Z(n46932) );
  AND U46991 ( .A(n1123), .B(n46994), .Z(n46993) );
  XNOR U46992 ( .A(n46995), .B(n46996), .Z(n46994) );
  XOR U46993 ( .A(n46997), .B(n46998), .Z(n46981) );
  AND U46994 ( .A(n46999), .B(n47000), .Z(n46998) );
  XNOR U46995 ( .A(n46997), .B(n46945), .Z(n47000) );
  XOR U46996 ( .A(n47001), .B(n46990), .Z(n46945) );
  XNOR U46997 ( .A(n47002), .B(n46985), .Z(n46990) );
  XOR U46998 ( .A(n47003), .B(n47004), .Z(n46985) );
  AND U46999 ( .A(n47005), .B(n47006), .Z(n47004) );
  XOR U47000 ( .A(n47007), .B(n47003), .Z(n47005) );
  XNOR U47001 ( .A(n47008), .B(n47009), .Z(n47002) );
  AND U47002 ( .A(n47010), .B(n47011), .Z(n47009) );
  XOR U47003 ( .A(n47008), .B(n47012), .Z(n47010) );
  XNOR U47004 ( .A(n46991), .B(n46988), .Z(n47001) );
  AND U47005 ( .A(n47013), .B(n47014), .Z(n46988) );
  XOR U47006 ( .A(n47015), .B(n47016), .Z(n46991) );
  AND U47007 ( .A(n47017), .B(n47018), .Z(n47016) );
  XOR U47008 ( .A(n47015), .B(n47019), .Z(n47017) );
  XNOR U47009 ( .A(n46942), .B(n46997), .Z(n46999) );
  XNOR U47010 ( .A(n47020), .B(n47021), .Z(n46942) );
  AND U47011 ( .A(n1123), .B(n47022), .Z(n47021) );
  XNOR U47012 ( .A(n47023), .B(n47024), .Z(n47022) );
  XOR U47013 ( .A(n47025), .B(n47026), .Z(n46997) );
  AND U47014 ( .A(n47027), .B(n47028), .Z(n47026) );
  XNOR U47015 ( .A(n47025), .B(n47013), .Z(n47028) );
  IV U47016 ( .A(n46955), .Z(n47013) );
  XNOR U47017 ( .A(n47029), .B(n47006), .Z(n46955) );
  XNOR U47018 ( .A(n47030), .B(n47012), .Z(n47006) );
  XOR U47019 ( .A(n47031), .B(n47032), .Z(n47012) );
  AND U47020 ( .A(n47033), .B(n47034), .Z(n47032) );
  XOR U47021 ( .A(n47031), .B(n47035), .Z(n47033) );
  XNOR U47022 ( .A(n47011), .B(n47003), .Z(n47030) );
  XOR U47023 ( .A(n47036), .B(n47037), .Z(n47003) );
  AND U47024 ( .A(n47038), .B(n47039), .Z(n47037) );
  XNOR U47025 ( .A(n47040), .B(n47036), .Z(n47038) );
  XNOR U47026 ( .A(n47041), .B(n47008), .Z(n47011) );
  XOR U47027 ( .A(n47042), .B(n47043), .Z(n47008) );
  AND U47028 ( .A(n47044), .B(n47045), .Z(n47043) );
  XOR U47029 ( .A(n47042), .B(n47046), .Z(n47044) );
  XNOR U47030 ( .A(n47047), .B(n47048), .Z(n47041) );
  AND U47031 ( .A(n47049), .B(n47050), .Z(n47048) );
  XNOR U47032 ( .A(n47047), .B(n47051), .Z(n47049) );
  XNOR U47033 ( .A(n47007), .B(n47014), .Z(n47029) );
  AND U47034 ( .A(n46963), .B(n47052), .Z(n47014) );
  XOR U47035 ( .A(n47019), .B(n47018), .Z(n47007) );
  XNOR U47036 ( .A(n47053), .B(n47015), .Z(n47018) );
  XOR U47037 ( .A(n47054), .B(n47055), .Z(n47015) );
  AND U47038 ( .A(n47056), .B(n47057), .Z(n47055) );
  XOR U47039 ( .A(n47054), .B(n47058), .Z(n47056) );
  XNOR U47040 ( .A(n47059), .B(n47060), .Z(n47053) );
  AND U47041 ( .A(n47061), .B(n47062), .Z(n47060) );
  XOR U47042 ( .A(n47059), .B(n47063), .Z(n47061) );
  XOR U47043 ( .A(n47064), .B(n47065), .Z(n47019) );
  AND U47044 ( .A(n47066), .B(n47067), .Z(n47065) );
  XOR U47045 ( .A(n47064), .B(n47068), .Z(n47066) );
  XNOR U47046 ( .A(n46952), .B(n47025), .Z(n47027) );
  XNOR U47047 ( .A(n47069), .B(n47070), .Z(n46952) );
  AND U47048 ( .A(n1123), .B(n47071), .Z(n47070) );
  XNOR U47049 ( .A(n47072), .B(n47073), .Z(n47071) );
  XOR U47050 ( .A(n47074), .B(n47075), .Z(n47025) );
  AND U47051 ( .A(n47076), .B(n47077), .Z(n47075) );
  XNOR U47052 ( .A(n47074), .B(n46963), .Z(n47077) );
  XOR U47053 ( .A(n47078), .B(n47039), .Z(n46963) );
  XNOR U47054 ( .A(n47079), .B(n47046), .Z(n47039) );
  XOR U47055 ( .A(n47035), .B(n47034), .Z(n47046) );
  XNOR U47056 ( .A(n47080), .B(n47031), .Z(n47034) );
  XOR U47057 ( .A(n47081), .B(n47082), .Z(n47031) );
  AND U47058 ( .A(n47083), .B(n47084), .Z(n47082) );
  XNOR U47059 ( .A(n47085), .B(n47086), .Z(n47083) );
  IV U47060 ( .A(n47081), .Z(n47085) );
  XNOR U47061 ( .A(n47087), .B(n47088), .Z(n47080) );
  NOR U47062 ( .A(n47089), .B(n47090), .Z(n47088) );
  XNOR U47063 ( .A(n47087), .B(n47091), .Z(n47089) );
  XOR U47064 ( .A(n47092), .B(n47093), .Z(n47035) );
  NOR U47065 ( .A(n47094), .B(n47095), .Z(n47093) );
  XNOR U47066 ( .A(n47092), .B(n47096), .Z(n47094) );
  XNOR U47067 ( .A(n47045), .B(n47036), .Z(n47079) );
  XOR U47068 ( .A(n47097), .B(n47098), .Z(n47036) );
  AND U47069 ( .A(n47099), .B(n47100), .Z(n47098) );
  XOR U47070 ( .A(n47097), .B(n47101), .Z(n47099) );
  XOR U47071 ( .A(n47102), .B(n47051), .Z(n47045) );
  XOR U47072 ( .A(n47103), .B(n47104), .Z(n47051) );
  NOR U47073 ( .A(n47105), .B(n47106), .Z(n47104) );
  XOR U47074 ( .A(n47103), .B(n47107), .Z(n47105) );
  XNOR U47075 ( .A(n47050), .B(n47042), .Z(n47102) );
  XOR U47076 ( .A(n47108), .B(n47109), .Z(n47042) );
  AND U47077 ( .A(n47110), .B(n47111), .Z(n47109) );
  XOR U47078 ( .A(n47108), .B(n47112), .Z(n47110) );
  XNOR U47079 ( .A(n47113), .B(n47047), .Z(n47050) );
  XOR U47080 ( .A(n47114), .B(n47115), .Z(n47047) );
  AND U47081 ( .A(n47116), .B(n47117), .Z(n47115) );
  XNOR U47082 ( .A(n47118), .B(n47119), .Z(n47116) );
  IV U47083 ( .A(n47114), .Z(n47118) );
  XNOR U47084 ( .A(n47120), .B(n47121), .Z(n47113) );
  NOR U47085 ( .A(n47122), .B(n47123), .Z(n47121) );
  XNOR U47086 ( .A(n47120), .B(n47124), .Z(n47122) );
  XOR U47087 ( .A(n47040), .B(n47052), .Z(n47078) );
  NOR U47088 ( .A(n46969), .B(n47125), .Z(n47052) );
  XNOR U47089 ( .A(n47058), .B(n47057), .Z(n47040) );
  XNOR U47090 ( .A(n47126), .B(n47063), .Z(n47057) );
  XNOR U47091 ( .A(n47127), .B(n47128), .Z(n47063) );
  NOR U47092 ( .A(n47129), .B(n47130), .Z(n47128) );
  XOR U47093 ( .A(n47127), .B(n47131), .Z(n47129) );
  XNOR U47094 ( .A(n47062), .B(n47054), .Z(n47126) );
  XOR U47095 ( .A(n47132), .B(n47133), .Z(n47054) );
  AND U47096 ( .A(n47134), .B(n47135), .Z(n47133) );
  XOR U47097 ( .A(n47132), .B(n47136), .Z(n47134) );
  XNOR U47098 ( .A(n47137), .B(n47059), .Z(n47062) );
  XOR U47099 ( .A(n47138), .B(n47139), .Z(n47059) );
  AND U47100 ( .A(n47140), .B(n47141), .Z(n47139) );
  XNOR U47101 ( .A(n47142), .B(n47143), .Z(n47140) );
  IV U47102 ( .A(n47138), .Z(n47142) );
  XNOR U47103 ( .A(n47144), .B(n47145), .Z(n47137) );
  NOR U47104 ( .A(n47146), .B(n47147), .Z(n47145) );
  XNOR U47105 ( .A(n47144), .B(n47148), .Z(n47146) );
  XOR U47106 ( .A(n47068), .B(n47067), .Z(n47058) );
  XNOR U47107 ( .A(n47149), .B(n47064), .Z(n47067) );
  XOR U47108 ( .A(n47150), .B(n47151), .Z(n47064) );
  AND U47109 ( .A(n47152), .B(n47153), .Z(n47151) );
  XNOR U47110 ( .A(n47154), .B(n47155), .Z(n47152) );
  IV U47111 ( .A(n47150), .Z(n47154) );
  XNOR U47112 ( .A(n47156), .B(n47157), .Z(n47149) );
  NOR U47113 ( .A(n47158), .B(n47159), .Z(n47157) );
  XNOR U47114 ( .A(n47156), .B(n47160), .Z(n47158) );
  XOR U47115 ( .A(n47161), .B(n47162), .Z(n47068) );
  NOR U47116 ( .A(n47163), .B(n47164), .Z(n47162) );
  XNOR U47117 ( .A(n47161), .B(n47165), .Z(n47163) );
  XNOR U47118 ( .A(n46960), .B(n47074), .Z(n47076) );
  XNOR U47119 ( .A(n47166), .B(n47167), .Z(n46960) );
  AND U47120 ( .A(n1123), .B(n47168), .Z(n47167) );
  XNOR U47121 ( .A(n47169), .B(n47170), .Z(n47168) );
  AND U47122 ( .A(n46966), .B(n46969), .Z(n47074) );
  XOR U47123 ( .A(n47171), .B(n47125), .Z(n46969) );
  XNOR U47124 ( .A(p_input[1664]), .B(p_input[2048]), .Z(n47125) );
  XNOR U47125 ( .A(n47101), .B(n47100), .Z(n47171) );
  XNOR U47126 ( .A(n47172), .B(n47112), .Z(n47100) );
  XOR U47127 ( .A(n47086), .B(n47084), .Z(n47112) );
  XNOR U47128 ( .A(n47173), .B(n47091), .Z(n47084) );
  XOR U47129 ( .A(p_input[1688]), .B(p_input[2072]), .Z(n47091) );
  XOR U47130 ( .A(n47081), .B(n47090), .Z(n47173) );
  XOR U47131 ( .A(n47174), .B(n47087), .Z(n47090) );
  XOR U47132 ( .A(p_input[1686]), .B(p_input[2070]), .Z(n47087) );
  XOR U47133 ( .A(p_input[1687]), .B(n29410), .Z(n47174) );
  XOR U47134 ( .A(p_input[1682]), .B(p_input[2066]), .Z(n47081) );
  XNOR U47135 ( .A(n47096), .B(n47095), .Z(n47086) );
  XOR U47136 ( .A(n47175), .B(n47092), .Z(n47095) );
  XOR U47137 ( .A(p_input[1683]), .B(p_input[2067]), .Z(n47092) );
  XOR U47138 ( .A(p_input[1684]), .B(n29412), .Z(n47175) );
  XOR U47139 ( .A(p_input[1685]), .B(p_input[2069]), .Z(n47096) );
  XOR U47140 ( .A(n47111), .B(n47176), .Z(n47172) );
  IV U47141 ( .A(n47097), .Z(n47176) );
  XOR U47142 ( .A(p_input[1665]), .B(p_input[2049]), .Z(n47097) );
  XNOR U47143 ( .A(n47177), .B(n47119), .Z(n47111) );
  XNOR U47144 ( .A(n47107), .B(n47106), .Z(n47119) );
  XNOR U47145 ( .A(n47178), .B(n47103), .Z(n47106) );
  XNOR U47146 ( .A(p_input[1690]), .B(p_input[2074]), .Z(n47103) );
  XOR U47147 ( .A(p_input[1691]), .B(n29415), .Z(n47178) );
  XOR U47148 ( .A(p_input[1692]), .B(p_input[2076]), .Z(n47107) );
  XOR U47149 ( .A(n47117), .B(n47179), .Z(n47177) );
  IV U47150 ( .A(n47108), .Z(n47179) );
  XOR U47151 ( .A(p_input[1681]), .B(p_input[2065]), .Z(n47108) );
  XNOR U47152 ( .A(n47180), .B(n47124), .Z(n47117) );
  XNOR U47153 ( .A(p_input[1695]), .B(n29418), .Z(n47124) );
  XOR U47154 ( .A(n47114), .B(n47123), .Z(n47180) );
  XOR U47155 ( .A(n47181), .B(n47120), .Z(n47123) );
  XOR U47156 ( .A(p_input[1693]), .B(p_input[2077]), .Z(n47120) );
  XOR U47157 ( .A(p_input[1694]), .B(n29420), .Z(n47181) );
  XOR U47158 ( .A(p_input[1689]), .B(p_input[2073]), .Z(n47114) );
  XOR U47159 ( .A(n47136), .B(n47135), .Z(n47101) );
  XNOR U47160 ( .A(n47182), .B(n47143), .Z(n47135) );
  XNOR U47161 ( .A(n47131), .B(n47130), .Z(n47143) );
  XNOR U47162 ( .A(n47183), .B(n47127), .Z(n47130) );
  XNOR U47163 ( .A(p_input[1675]), .B(p_input[2059]), .Z(n47127) );
  XOR U47164 ( .A(p_input[1676]), .B(n28329), .Z(n47183) );
  XOR U47165 ( .A(p_input[1677]), .B(p_input[2061]), .Z(n47131) );
  XOR U47166 ( .A(n47141), .B(n47184), .Z(n47182) );
  IV U47167 ( .A(n47132), .Z(n47184) );
  XOR U47168 ( .A(p_input[1666]), .B(p_input[2050]), .Z(n47132) );
  XNOR U47169 ( .A(n47185), .B(n47148), .Z(n47141) );
  XNOR U47170 ( .A(p_input[1680]), .B(n28332), .Z(n47148) );
  XOR U47171 ( .A(n47138), .B(n47147), .Z(n47185) );
  XOR U47172 ( .A(n47186), .B(n47144), .Z(n47147) );
  XOR U47173 ( .A(p_input[1678]), .B(p_input[2062]), .Z(n47144) );
  XOR U47174 ( .A(p_input[1679]), .B(n28334), .Z(n47186) );
  XOR U47175 ( .A(p_input[1674]), .B(p_input[2058]), .Z(n47138) );
  XOR U47176 ( .A(n47155), .B(n47153), .Z(n47136) );
  XNOR U47177 ( .A(n47187), .B(n47160), .Z(n47153) );
  XOR U47178 ( .A(p_input[1673]), .B(p_input[2057]), .Z(n47160) );
  XOR U47179 ( .A(n47150), .B(n47159), .Z(n47187) );
  XOR U47180 ( .A(n47188), .B(n47156), .Z(n47159) );
  XOR U47181 ( .A(p_input[1671]), .B(p_input[2055]), .Z(n47156) );
  XOR U47182 ( .A(p_input[1672]), .B(n29427), .Z(n47188) );
  XOR U47183 ( .A(p_input[1667]), .B(p_input[2051]), .Z(n47150) );
  XNOR U47184 ( .A(n47165), .B(n47164), .Z(n47155) );
  XOR U47185 ( .A(n47189), .B(n47161), .Z(n47164) );
  XOR U47186 ( .A(p_input[1668]), .B(p_input[2052]), .Z(n47161) );
  XOR U47187 ( .A(p_input[1669]), .B(n29429), .Z(n47189) );
  XOR U47188 ( .A(p_input[1670]), .B(p_input[2054]), .Z(n47165) );
  XNOR U47189 ( .A(n47190), .B(n47191), .Z(n46966) );
  AND U47190 ( .A(n1123), .B(n47192), .Z(n47191) );
  XNOR U47191 ( .A(n47193), .B(n47194), .Z(n1123) );
  AND U47192 ( .A(n47195), .B(n47196), .Z(n47194) );
  XOR U47193 ( .A(n46980), .B(n47193), .Z(n47196) );
  XNOR U47194 ( .A(n47197), .B(n47193), .Z(n47195) );
  XOR U47195 ( .A(n47198), .B(n47199), .Z(n47193) );
  AND U47196 ( .A(n47200), .B(n47201), .Z(n47199) );
  XOR U47197 ( .A(n46995), .B(n47198), .Z(n47201) );
  XOR U47198 ( .A(n47198), .B(n46996), .Z(n47200) );
  XOR U47199 ( .A(n47202), .B(n47203), .Z(n47198) );
  AND U47200 ( .A(n47204), .B(n47205), .Z(n47203) );
  XOR U47201 ( .A(n47023), .B(n47202), .Z(n47205) );
  XOR U47202 ( .A(n47202), .B(n47024), .Z(n47204) );
  XOR U47203 ( .A(n47206), .B(n47207), .Z(n47202) );
  AND U47204 ( .A(n47208), .B(n47209), .Z(n47207) );
  XOR U47205 ( .A(n47072), .B(n47206), .Z(n47209) );
  XOR U47206 ( .A(n47206), .B(n47073), .Z(n47208) );
  XOR U47207 ( .A(n47210), .B(n47211), .Z(n47206) );
  AND U47208 ( .A(n47212), .B(n47213), .Z(n47211) );
  XOR U47209 ( .A(n47210), .B(n47169), .Z(n47213) );
  XNOR U47210 ( .A(n47214), .B(n47215), .Z(n46916) );
  AND U47211 ( .A(n1127), .B(n47216), .Z(n47215) );
  XNOR U47212 ( .A(n47217), .B(n47218), .Z(n1127) );
  AND U47213 ( .A(n47219), .B(n47220), .Z(n47218) );
  XOR U47214 ( .A(n47217), .B(n46926), .Z(n47220) );
  XNOR U47215 ( .A(n47217), .B(n46876), .Z(n47219) );
  XOR U47216 ( .A(n47221), .B(n47222), .Z(n47217) );
  AND U47217 ( .A(n47223), .B(n47224), .Z(n47222) );
  XNOR U47218 ( .A(n46936), .B(n47221), .Z(n47224) );
  XOR U47219 ( .A(n47221), .B(n46886), .Z(n47223) );
  XOR U47220 ( .A(n47225), .B(n47226), .Z(n47221) );
  AND U47221 ( .A(n47227), .B(n47228), .Z(n47226) );
  XNOR U47222 ( .A(n46946), .B(n47225), .Z(n47228) );
  XOR U47223 ( .A(n47225), .B(n46895), .Z(n47227) );
  XOR U47224 ( .A(n47229), .B(n47230), .Z(n47225) );
  AND U47225 ( .A(n47231), .B(n47232), .Z(n47230) );
  XOR U47226 ( .A(n47229), .B(n46903), .Z(n47231) );
  XOR U47227 ( .A(n47233), .B(n47234), .Z(n46867) );
  AND U47228 ( .A(n1131), .B(n47216), .Z(n47234) );
  XNOR U47229 ( .A(n47214), .B(n47233), .Z(n47216) );
  XNOR U47230 ( .A(n47235), .B(n47236), .Z(n1131) );
  AND U47231 ( .A(n47237), .B(n47238), .Z(n47236) );
  XNOR U47232 ( .A(n47239), .B(n47235), .Z(n47238) );
  IV U47233 ( .A(n46926), .Z(n47239) );
  XOR U47234 ( .A(n47197), .B(n47240), .Z(n46926) );
  AND U47235 ( .A(n1134), .B(n47241), .Z(n47240) );
  XOR U47236 ( .A(n46979), .B(n46976), .Z(n47241) );
  IV U47237 ( .A(n47197), .Z(n46979) );
  XNOR U47238 ( .A(n46876), .B(n47235), .Z(n47237) );
  XOR U47239 ( .A(n47242), .B(n47243), .Z(n46876) );
  AND U47240 ( .A(n1150), .B(n47244), .Z(n47243) );
  XOR U47241 ( .A(n47245), .B(n47246), .Z(n47235) );
  AND U47242 ( .A(n47247), .B(n47248), .Z(n47246) );
  XNOR U47243 ( .A(n47245), .B(n46936), .Z(n47248) );
  XOR U47244 ( .A(n46996), .B(n47249), .Z(n46936) );
  AND U47245 ( .A(n1134), .B(n47250), .Z(n47249) );
  XOR U47246 ( .A(n46992), .B(n46996), .Z(n47250) );
  XNOR U47247 ( .A(n47251), .B(n47245), .Z(n47247) );
  IV U47248 ( .A(n46886), .Z(n47251) );
  XOR U47249 ( .A(n47252), .B(n47253), .Z(n46886) );
  AND U47250 ( .A(n1150), .B(n47254), .Z(n47253) );
  XOR U47251 ( .A(n47255), .B(n47256), .Z(n47245) );
  AND U47252 ( .A(n47257), .B(n47258), .Z(n47256) );
  XNOR U47253 ( .A(n47255), .B(n46946), .Z(n47258) );
  XOR U47254 ( .A(n47024), .B(n47259), .Z(n46946) );
  AND U47255 ( .A(n1134), .B(n47260), .Z(n47259) );
  XOR U47256 ( .A(n47020), .B(n47024), .Z(n47260) );
  XOR U47257 ( .A(n46895), .B(n47255), .Z(n47257) );
  XOR U47258 ( .A(n47261), .B(n47262), .Z(n46895) );
  AND U47259 ( .A(n1150), .B(n47263), .Z(n47262) );
  XOR U47260 ( .A(n47229), .B(n47264), .Z(n47255) );
  AND U47261 ( .A(n47265), .B(n47232), .Z(n47264) );
  XNOR U47262 ( .A(n46956), .B(n47229), .Z(n47232) );
  XOR U47263 ( .A(n47073), .B(n47266), .Z(n46956) );
  AND U47264 ( .A(n1134), .B(n47267), .Z(n47266) );
  XOR U47265 ( .A(n47069), .B(n47073), .Z(n47267) );
  XNOR U47266 ( .A(n47268), .B(n47229), .Z(n47265) );
  IV U47267 ( .A(n46903), .Z(n47268) );
  XOR U47268 ( .A(n47269), .B(n47270), .Z(n46903) );
  AND U47269 ( .A(n1150), .B(n47271), .Z(n47270) );
  XOR U47270 ( .A(n47272), .B(n47273), .Z(n47229) );
  AND U47271 ( .A(n47274), .B(n47275), .Z(n47273) );
  XNOR U47272 ( .A(n47272), .B(n46964), .Z(n47275) );
  XOR U47273 ( .A(n47170), .B(n47276), .Z(n46964) );
  AND U47274 ( .A(n1134), .B(n47277), .Z(n47276) );
  XOR U47275 ( .A(n47166), .B(n47170), .Z(n47277) );
  XNOR U47276 ( .A(n47278), .B(n47272), .Z(n47274) );
  IV U47277 ( .A(n46913), .Z(n47278) );
  XOR U47278 ( .A(n47279), .B(n47280), .Z(n46913) );
  AND U47279 ( .A(n1150), .B(n47281), .Z(n47280) );
  AND U47280 ( .A(n47233), .B(n47214), .Z(n47272) );
  XNOR U47281 ( .A(n47282), .B(n47283), .Z(n47214) );
  AND U47282 ( .A(n1134), .B(n47192), .Z(n47283) );
  XNOR U47283 ( .A(n47190), .B(n47282), .Z(n47192) );
  XNOR U47284 ( .A(n47284), .B(n47285), .Z(n1134) );
  AND U47285 ( .A(n47286), .B(n47287), .Z(n47285) );
  XNOR U47286 ( .A(n47284), .B(n46976), .Z(n47287) );
  IV U47287 ( .A(n46980), .Z(n46976) );
  XOR U47288 ( .A(n47288), .B(n47289), .Z(n46980) );
  AND U47289 ( .A(n1138), .B(n47290), .Z(n47289) );
  XOR U47290 ( .A(n47291), .B(n47288), .Z(n47290) );
  XNOR U47291 ( .A(n47284), .B(n47197), .Z(n47286) );
  XOR U47292 ( .A(n47292), .B(n47293), .Z(n47197) );
  AND U47293 ( .A(n1146), .B(n47244), .Z(n47293) );
  XOR U47294 ( .A(n47242), .B(n47292), .Z(n47244) );
  XOR U47295 ( .A(n47294), .B(n47295), .Z(n47284) );
  AND U47296 ( .A(n47296), .B(n47297), .Z(n47295) );
  XNOR U47297 ( .A(n47294), .B(n46992), .Z(n47297) );
  IV U47298 ( .A(n46995), .Z(n46992) );
  XOR U47299 ( .A(n47298), .B(n47299), .Z(n46995) );
  AND U47300 ( .A(n1138), .B(n47300), .Z(n47299) );
  XOR U47301 ( .A(n47301), .B(n47298), .Z(n47300) );
  XOR U47302 ( .A(n46996), .B(n47294), .Z(n47296) );
  XOR U47303 ( .A(n47302), .B(n47303), .Z(n46996) );
  AND U47304 ( .A(n1146), .B(n47254), .Z(n47303) );
  XOR U47305 ( .A(n47302), .B(n47252), .Z(n47254) );
  XOR U47306 ( .A(n47304), .B(n47305), .Z(n47294) );
  AND U47307 ( .A(n47306), .B(n47307), .Z(n47305) );
  XNOR U47308 ( .A(n47304), .B(n47020), .Z(n47307) );
  IV U47309 ( .A(n47023), .Z(n47020) );
  XOR U47310 ( .A(n47308), .B(n47309), .Z(n47023) );
  AND U47311 ( .A(n1138), .B(n47310), .Z(n47309) );
  XNOR U47312 ( .A(n47311), .B(n47308), .Z(n47310) );
  XOR U47313 ( .A(n47024), .B(n47304), .Z(n47306) );
  XOR U47314 ( .A(n47312), .B(n47313), .Z(n47024) );
  AND U47315 ( .A(n1146), .B(n47263), .Z(n47313) );
  XOR U47316 ( .A(n47312), .B(n47261), .Z(n47263) );
  XOR U47317 ( .A(n47314), .B(n47315), .Z(n47304) );
  AND U47318 ( .A(n47316), .B(n47317), .Z(n47315) );
  XNOR U47319 ( .A(n47314), .B(n47069), .Z(n47317) );
  IV U47320 ( .A(n47072), .Z(n47069) );
  XOR U47321 ( .A(n47318), .B(n47319), .Z(n47072) );
  AND U47322 ( .A(n1138), .B(n47320), .Z(n47319) );
  XOR U47323 ( .A(n47321), .B(n47318), .Z(n47320) );
  XOR U47324 ( .A(n47073), .B(n47314), .Z(n47316) );
  XOR U47325 ( .A(n47322), .B(n47323), .Z(n47073) );
  AND U47326 ( .A(n1146), .B(n47271), .Z(n47323) );
  XOR U47327 ( .A(n47322), .B(n47269), .Z(n47271) );
  XOR U47328 ( .A(n47210), .B(n47324), .Z(n47314) );
  AND U47329 ( .A(n47212), .B(n47325), .Z(n47324) );
  XNOR U47330 ( .A(n47210), .B(n47166), .Z(n47325) );
  IV U47331 ( .A(n47169), .Z(n47166) );
  XOR U47332 ( .A(n47326), .B(n47327), .Z(n47169) );
  AND U47333 ( .A(n1138), .B(n47328), .Z(n47327) );
  XNOR U47334 ( .A(n47329), .B(n47326), .Z(n47328) );
  XOR U47335 ( .A(n47170), .B(n47210), .Z(n47212) );
  XOR U47336 ( .A(n47330), .B(n47331), .Z(n47170) );
  AND U47337 ( .A(n1146), .B(n47281), .Z(n47331) );
  XOR U47338 ( .A(n47330), .B(n47279), .Z(n47281) );
  AND U47339 ( .A(n47282), .B(n47190), .Z(n47210) );
  XNOR U47340 ( .A(n47332), .B(n47333), .Z(n47190) );
  AND U47341 ( .A(n1138), .B(n47334), .Z(n47333) );
  XNOR U47342 ( .A(n47335), .B(n47332), .Z(n47334) );
  XNOR U47343 ( .A(n47336), .B(n47337), .Z(n1138) );
  AND U47344 ( .A(n47338), .B(n47339), .Z(n47337) );
  XOR U47345 ( .A(n47291), .B(n47336), .Z(n47339) );
  AND U47346 ( .A(n47340), .B(n47341), .Z(n47291) );
  XNOR U47347 ( .A(n47288), .B(n47336), .Z(n47338) );
  XNOR U47348 ( .A(n47342), .B(n47343), .Z(n47288) );
  AND U47349 ( .A(n1142), .B(n47344), .Z(n47343) );
  XNOR U47350 ( .A(n47345), .B(n47346), .Z(n47344) );
  XOR U47351 ( .A(n47347), .B(n47348), .Z(n47336) );
  AND U47352 ( .A(n47349), .B(n47350), .Z(n47348) );
  XNOR U47353 ( .A(n47347), .B(n47340), .Z(n47350) );
  IV U47354 ( .A(n47301), .Z(n47340) );
  XOR U47355 ( .A(n47351), .B(n47352), .Z(n47301) );
  XOR U47356 ( .A(n47353), .B(n47341), .Z(n47352) );
  AND U47357 ( .A(n47311), .B(n47354), .Z(n47341) );
  AND U47358 ( .A(n47355), .B(n47356), .Z(n47353) );
  XOR U47359 ( .A(n47357), .B(n47351), .Z(n47355) );
  XNOR U47360 ( .A(n47298), .B(n47347), .Z(n47349) );
  XNOR U47361 ( .A(n47358), .B(n47359), .Z(n47298) );
  AND U47362 ( .A(n1142), .B(n47360), .Z(n47359) );
  XNOR U47363 ( .A(n47361), .B(n47362), .Z(n47360) );
  XOR U47364 ( .A(n47363), .B(n47364), .Z(n47347) );
  AND U47365 ( .A(n47365), .B(n47366), .Z(n47364) );
  XNOR U47366 ( .A(n47363), .B(n47311), .Z(n47366) );
  XOR U47367 ( .A(n47367), .B(n47356), .Z(n47311) );
  XNOR U47368 ( .A(n47368), .B(n47351), .Z(n47356) );
  XOR U47369 ( .A(n47369), .B(n47370), .Z(n47351) );
  AND U47370 ( .A(n47371), .B(n47372), .Z(n47370) );
  XOR U47371 ( .A(n47373), .B(n47369), .Z(n47371) );
  XNOR U47372 ( .A(n47374), .B(n47375), .Z(n47368) );
  AND U47373 ( .A(n47376), .B(n47377), .Z(n47375) );
  XOR U47374 ( .A(n47374), .B(n47378), .Z(n47376) );
  XNOR U47375 ( .A(n47357), .B(n47354), .Z(n47367) );
  AND U47376 ( .A(n47379), .B(n47380), .Z(n47354) );
  XOR U47377 ( .A(n47381), .B(n47382), .Z(n47357) );
  AND U47378 ( .A(n47383), .B(n47384), .Z(n47382) );
  XOR U47379 ( .A(n47381), .B(n47385), .Z(n47383) );
  XNOR U47380 ( .A(n47308), .B(n47363), .Z(n47365) );
  XNOR U47381 ( .A(n47386), .B(n47387), .Z(n47308) );
  AND U47382 ( .A(n1142), .B(n47388), .Z(n47387) );
  XNOR U47383 ( .A(n47389), .B(n47390), .Z(n47388) );
  XOR U47384 ( .A(n47391), .B(n47392), .Z(n47363) );
  AND U47385 ( .A(n47393), .B(n47394), .Z(n47392) );
  XNOR U47386 ( .A(n47391), .B(n47379), .Z(n47394) );
  IV U47387 ( .A(n47321), .Z(n47379) );
  XNOR U47388 ( .A(n47395), .B(n47372), .Z(n47321) );
  XNOR U47389 ( .A(n47396), .B(n47378), .Z(n47372) );
  XOR U47390 ( .A(n47397), .B(n47398), .Z(n47378) );
  AND U47391 ( .A(n47399), .B(n47400), .Z(n47398) );
  XOR U47392 ( .A(n47397), .B(n47401), .Z(n47399) );
  XNOR U47393 ( .A(n47377), .B(n47369), .Z(n47396) );
  XOR U47394 ( .A(n47402), .B(n47403), .Z(n47369) );
  AND U47395 ( .A(n47404), .B(n47405), .Z(n47403) );
  XNOR U47396 ( .A(n47406), .B(n47402), .Z(n47404) );
  XNOR U47397 ( .A(n47407), .B(n47374), .Z(n47377) );
  XOR U47398 ( .A(n47408), .B(n47409), .Z(n47374) );
  AND U47399 ( .A(n47410), .B(n47411), .Z(n47409) );
  XOR U47400 ( .A(n47408), .B(n47412), .Z(n47410) );
  XNOR U47401 ( .A(n47413), .B(n47414), .Z(n47407) );
  AND U47402 ( .A(n47415), .B(n47416), .Z(n47414) );
  XNOR U47403 ( .A(n47413), .B(n47417), .Z(n47415) );
  XNOR U47404 ( .A(n47373), .B(n47380), .Z(n47395) );
  AND U47405 ( .A(n47329), .B(n47418), .Z(n47380) );
  XOR U47406 ( .A(n47385), .B(n47384), .Z(n47373) );
  XNOR U47407 ( .A(n47419), .B(n47381), .Z(n47384) );
  XOR U47408 ( .A(n47420), .B(n47421), .Z(n47381) );
  AND U47409 ( .A(n47422), .B(n47423), .Z(n47421) );
  XOR U47410 ( .A(n47420), .B(n47424), .Z(n47422) );
  XNOR U47411 ( .A(n47425), .B(n47426), .Z(n47419) );
  AND U47412 ( .A(n47427), .B(n47428), .Z(n47426) );
  XOR U47413 ( .A(n47425), .B(n47429), .Z(n47427) );
  XOR U47414 ( .A(n47430), .B(n47431), .Z(n47385) );
  AND U47415 ( .A(n47432), .B(n47433), .Z(n47431) );
  XOR U47416 ( .A(n47430), .B(n47434), .Z(n47432) );
  XNOR U47417 ( .A(n47318), .B(n47391), .Z(n47393) );
  XNOR U47418 ( .A(n47435), .B(n47436), .Z(n47318) );
  AND U47419 ( .A(n1142), .B(n47437), .Z(n47436) );
  XNOR U47420 ( .A(n47438), .B(n47439), .Z(n47437) );
  XOR U47421 ( .A(n47440), .B(n47441), .Z(n47391) );
  AND U47422 ( .A(n47442), .B(n47443), .Z(n47441) );
  XNOR U47423 ( .A(n47440), .B(n47329), .Z(n47443) );
  XOR U47424 ( .A(n47444), .B(n47405), .Z(n47329) );
  XNOR U47425 ( .A(n47445), .B(n47412), .Z(n47405) );
  XOR U47426 ( .A(n47401), .B(n47400), .Z(n47412) );
  XNOR U47427 ( .A(n47446), .B(n47397), .Z(n47400) );
  XOR U47428 ( .A(n47447), .B(n47448), .Z(n47397) );
  AND U47429 ( .A(n47449), .B(n47450), .Z(n47448) );
  XNOR U47430 ( .A(n47451), .B(n47452), .Z(n47449) );
  IV U47431 ( .A(n47447), .Z(n47451) );
  XNOR U47432 ( .A(n47453), .B(n47454), .Z(n47446) );
  NOR U47433 ( .A(n47455), .B(n47456), .Z(n47454) );
  XNOR U47434 ( .A(n47453), .B(n47457), .Z(n47455) );
  XOR U47435 ( .A(n47458), .B(n47459), .Z(n47401) );
  NOR U47436 ( .A(n47460), .B(n47461), .Z(n47459) );
  XNOR U47437 ( .A(n47458), .B(n47462), .Z(n47460) );
  XNOR U47438 ( .A(n47411), .B(n47402), .Z(n47445) );
  XOR U47439 ( .A(n47463), .B(n47464), .Z(n47402) );
  AND U47440 ( .A(n47465), .B(n47466), .Z(n47464) );
  XOR U47441 ( .A(n47463), .B(n47467), .Z(n47465) );
  XOR U47442 ( .A(n47468), .B(n47417), .Z(n47411) );
  XOR U47443 ( .A(n47469), .B(n47470), .Z(n47417) );
  NOR U47444 ( .A(n47471), .B(n47472), .Z(n47470) );
  XOR U47445 ( .A(n47469), .B(n47473), .Z(n47471) );
  XNOR U47446 ( .A(n47416), .B(n47408), .Z(n47468) );
  XOR U47447 ( .A(n47474), .B(n47475), .Z(n47408) );
  AND U47448 ( .A(n47476), .B(n47477), .Z(n47475) );
  XOR U47449 ( .A(n47474), .B(n47478), .Z(n47476) );
  XNOR U47450 ( .A(n47479), .B(n47413), .Z(n47416) );
  XOR U47451 ( .A(n47480), .B(n47481), .Z(n47413) );
  AND U47452 ( .A(n47482), .B(n47483), .Z(n47481) );
  XNOR U47453 ( .A(n47484), .B(n47485), .Z(n47482) );
  IV U47454 ( .A(n47480), .Z(n47484) );
  XNOR U47455 ( .A(n47486), .B(n47487), .Z(n47479) );
  NOR U47456 ( .A(n47488), .B(n47489), .Z(n47487) );
  XNOR U47457 ( .A(n47486), .B(n47490), .Z(n47488) );
  XOR U47458 ( .A(n47406), .B(n47418), .Z(n47444) );
  NOR U47459 ( .A(n47335), .B(n47491), .Z(n47418) );
  XNOR U47460 ( .A(n47424), .B(n47423), .Z(n47406) );
  XNOR U47461 ( .A(n47492), .B(n47429), .Z(n47423) );
  XNOR U47462 ( .A(n47493), .B(n47494), .Z(n47429) );
  NOR U47463 ( .A(n47495), .B(n47496), .Z(n47494) );
  XOR U47464 ( .A(n47493), .B(n47497), .Z(n47495) );
  XNOR U47465 ( .A(n47428), .B(n47420), .Z(n47492) );
  XOR U47466 ( .A(n47498), .B(n47499), .Z(n47420) );
  AND U47467 ( .A(n47500), .B(n47501), .Z(n47499) );
  XOR U47468 ( .A(n47498), .B(n47502), .Z(n47500) );
  XNOR U47469 ( .A(n47503), .B(n47425), .Z(n47428) );
  XOR U47470 ( .A(n47504), .B(n47505), .Z(n47425) );
  AND U47471 ( .A(n47506), .B(n47507), .Z(n47505) );
  XNOR U47472 ( .A(n47508), .B(n47509), .Z(n47506) );
  IV U47473 ( .A(n47504), .Z(n47508) );
  XNOR U47474 ( .A(n47510), .B(n47511), .Z(n47503) );
  NOR U47475 ( .A(n47512), .B(n47513), .Z(n47511) );
  XNOR U47476 ( .A(n47510), .B(n47514), .Z(n47512) );
  XOR U47477 ( .A(n47434), .B(n47433), .Z(n47424) );
  XNOR U47478 ( .A(n47515), .B(n47430), .Z(n47433) );
  XOR U47479 ( .A(n47516), .B(n47517), .Z(n47430) );
  AND U47480 ( .A(n47518), .B(n47519), .Z(n47517) );
  XNOR U47481 ( .A(n47520), .B(n47521), .Z(n47518) );
  IV U47482 ( .A(n47516), .Z(n47520) );
  XNOR U47483 ( .A(n47522), .B(n47523), .Z(n47515) );
  NOR U47484 ( .A(n47524), .B(n47525), .Z(n47523) );
  XNOR U47485 ( .A(n47522), .B(n47526), .Z(n47524) );
  XOR U47486 ( .A(n47527), .B(n47528), .Z(n47434) );
  NOR U47487 ( .A(n47529), .B(n47530), .Z(n47528) );
  XNOR U47488 ( .A(n47527), .B(n47531), .Z(n47529) );
  XNOR U47489 ( .A(n47326), .B(n47440), .Z(n47442) );
  XNOR U47490 ( .A(n47532), .B(n47533), .Z(n47326) );
  AND U47491 ( .A(n1142), .B(n47534), .Z(n47533) );
  XNOR U47492 ( .A(n47535), .B(n47536), .Z(n47534) );
  AND U47493 ( .A(n47332), .B(n47335), .Z(n47440) );
  XOR U47494 ( .A(n47537), .B(n47491), .Z(n47335) );
  XNOR U47495 ( .A(p_input[1696]), .B(p_input[2048]), .Z(n47491) );
  XNOR U47496 ( .A(n47467), .B(n47466), .Z(n47537) );
  XNOR U47497 ( .A(n47538), .B(n47478), .Z(n47466) );
  XOR U47498 ( .A(n47452), .B(n47450), .Z(n47478) );
  XNOR U47499 ( .A(n47539), .B(n47457), .Z(n47450) );
  XOR U47500 ( .A(p_input[1720]), .B(p_input[2072]), .Z(n47457) );
  XOR U47501 ( .A(n47447), .B(n47456), .Z(n47539) );
  XOR U47502 ( .A(n47540), .B(n47453), .Z(n47456) );
  XOR U47503 ( .A(p_input[1718]), .B(p_input[2070]), .Z(n47453) );
  XOR U47504 ( .A(p_input[1719]), .B(n29410), .Z(n47540) );
  XOR U47505 ( .A(p_input[1714]), .B(p_input[2066]), .Z(n47447) );
  XNOR U47506 ( .A(n47462), .B(n47461), .Z(n47452) );
  XOR U47507 ( .A(n47541), .B(n47458), .Z(n47461) );
  XOR U47508 ( .A(p_input[1715]), .B(p_input[2067]), .Z(n47458) );
  XOR U47509 ( .A(p_input[1716]), .B(n29412), .Z(n47541) );
  XOR U47510 ( .A(p_input[1717]), .B(p_input[2069]), .Z(n47462) );
  XOR U47511 ( .A(n47477), .B(n47542), .Z(n47538) );
  IV U47512 ( .A(n47463), .Z(n47542) );
  XOR U47513 ( .A(p_input[1697]), .B(p_input[2049]), .Z(n47463) );
  XNOR U47514 ( .A(n47543), .B(n47485), .Z(n47477) );
  XNOR U47515 ( .A(n47473), .B(n47472), .Z(n47485) );
  XNOR U47516 ( .A(n47544), .B(n47469), .Z(n47472) );
  XNOR U47517 ( .A(p_input[1722]), .B(p_input[2074]), .Z(n47469) );
  XOR U47518 ( .A(p_input[1723]), .B(n29415), .Z(n47544) );
  XOR U47519 ( .A(p_input[1724]), .B(p_input[2076]), .Z(n47473) );
  XOR U47520 ( .A(n47483), .B(n47545), .Z(n47543) );
  IV U47521 ( .A(n47474), .Z(n47545) );
  XOR U47522 ( .A(p_input[1713]), .B(p_input[2065]), .Z(n47474) );
  XNOR U47523 ( .A(n47546), .B(n47490), .Z(n47483) );
  XNOR U47524 ( .A(p_input[1727]), .B(n29418), .Z(n47490) );
  XOR U47525 ( .A(n47480), .B(n47489), .Z(n47546) );
  XOR U47526 ( .A(n47547), .B(n47486), .Z(n47489) );
  XOR U47527 ( .A(p_input[1725]), .B(p_input[2077]), .Z(n47486) );
  XOR U47528 ( .A(p_input[1726]), .B(n29420), .Z(n47547) );
  XOR U47529 ( .A(p_input[1721]), .B(p_input[2073]), .Z(n47480) );
  XOR U47530 ( .A(n47502), .B(n47501), .Z(n47467) );
  XNOR U47531 ( .A(n47548), .B(n47509), .Z(n47501) );
  XNOR U47532 ( .A(n47497), .B(n47496), .Z(n47509) );
  XNOR U47533 ( .A(n47549), .B(n47493), .Z(n47496) );
  XNOR U47534 ( .A(p_input[1707]), .B(p_input[2059]), .Z(n47493) );
  XOR U47535 ( .A(p_input[1708]), .B(n28329), .Z(n47549) );
  XOR U47536 ( .A(p_input[1709]), .B(p_input[2061]), .Z(n47497) );
  XOR U47537 ( .A(n47507), .B(n47550), .Z(n47548) );
  IV U47538 ( .A(n47498), .Z(n47550) );
  XOR U47539 ( .A(p_input[1698]), .B(p_input[2050]), .Z(n47498) );
  XNOR U47540 ( .A(n47551), .B(n47514), .Z(n47507) );
  XNOR U47541 ( .A(p_input[1712]), .B(n28332), .Z(n47514) );
  XOR U47542 ( .A(n47504), .B(n47513), .Z(n47551) );
  XOR U47543 ( .A(n47552), .B(n47510), .Z(n47513) );
  XOR U47544 ( .A(p_input[1710]), .B(p_input[2062]), .Z(n47510) );
  XOR U47545 ( .A(p_input[1711]), .B(n28334), .Z(n47552) );
  XOR U47546 ( .A(p_input[1706]), .B(p_input[2058]), .Z(n47504) );
  XOR U47547 ( .A(n47521), .B(n47519), .Z(n47502) );
  XNOR U47548 ( .A(n47553), .B(n47526), .Z(n47519) );
  XOR U47549 ( .A(p_input[1705]), .B(p_input[2057]), .Z(n47526) );
  XOR U47550 ( .A(n47516), .B(n47525), .Z(n47553) );
  XOR U47551 ( .A(n47554), .B(n47522), .Z(n47525) );
  XOR U47552 ( .A(p_input[1703]), .B(p_input[2055]), .Z(n47522) );
  XOR U47553 ( .A(p_input[1704]), .B(n29427), .Z(n47554) );
  XOR U47554 ( .A(p_input[1699]), .B(p_input[2051]), .Z(n47516) );
  XNOR U47555 ( .A(n47531), .B(n47530), .Z(n47521) );
  XOR U47556 ( .A(n47555), .B(n47527), .Z(n47530) );
  XOR U47557 ( .A(p_input[1700]), .B(p_input[2052]), .Z(n47527) );
  XOR U47558 ( .A(p_input[1701]), .B(n29429), .Z(n47555) );
  XOR U47559 ( .A(p_input[1702]), .B(p_input[2054]), .Z(n47531) );
  XNOR U47560 ( .A(n47556), .B(n47557), .Z(n47332) );
  AND U47561 ( .A(n1142), .B(n47558), .Z(n47557) );
  XNOR U47562 ( .A(n47559), .B(n47560), .Z(n1142) );
  AND U47563 ( .A(n47561), .B(n47562), .Z(n47560) );
  XOR U47564 ( .A(n47346), .B(n47559), .Z(n47562) );
  XNOR U47565 ( .A(n47563), .B(n47559), .Z(n47561) );
  XOR U47566 ( .A(n47564), .B(n47565), .Z(n47559) );
  AND U47567 ( .A(n47566), .B(n47567), .Z(n47565) );
  XOR U47568 ( .A(n47361), .B(n47564), .Z(n47567) );
  XOR U47569 ( .A(n47564), .B(n47362), .Z(n47566) );
  XOR U47570 ( .A(n47568), .B(n47569), .Z(n47564) );
  AND U47571 ( .A(n47570), .B(n47571), .Z(n47569) );
  XOR U47572 ( .A(n47389), .B(n47568), .Z(n47571) );
  XOR U47573 ( .A(n47568), .B(n47390), .Z(n47570) );
  XOR U47574 ( .A(n47572), .B(n47573), .Z(n47568) );
  AND U47575 ( .A(n47574), .B(n47575), .Z(n47573) );
  XOR U47576 ( .A(n47438), .B(n47572), .Z(n47575) );
  XOR U47577 ( .A(n47572), .B(n47439), .Z(n47574) );
  XOR U47578 ( .A(n47576), .B(n47577), .Z(n47572) );
  AND U47579 ( .A(n47578), .B(n47579), .Z(n47577) );
  XOR U47580 ( .A(n47576), .B(n47535), .Z(n47579) );
  XNOR U47581 ( .A(n47580), .B(n47581), .Z(n47282) );
  AND U47582 ( .A(n1146), .B(n47582), .Z(n47581) );
  XNOR U47583 ( .A(n47583), .B(n47584), .Z(n1146) );
  AND U47584 ( .A(n47585), .B(n47586), .Z(n47584) );
  XOR U47585 ( .A(n47583), .B(n47292), .Z(n47586) );
  XNOR U47586 ( .A(n47583), .B(n47242), .Z(n47585) );
  XOR U47587 ( .A(n47587), .B(n47588), .Z(n47583) );
  AND U47588 ( .A(n47589), .B(n47590), .Z(n47588) );
  XNOR U47589 ( .A(n47302), .B(n47587), .Z(n47590) );
  XOR U47590 ( .A(n47587), .B(n47252), .Z(n47589) );
  XOR U47591 ( .A(n47591), .B(n47592), .Z(n47587) );
  AND U47592 ( .A(n47593), .B(n47594), .Z(n47592) );
  XNOR U47593 ( .A(n47312), .B(n47591), .Z(n47594) );
  XOR U47594 ( .A(n47591), .B(n47261), .Z(n47593) );
  XOR U47595 ( .A(n47595), .B(n47596), .Z(n47591) );
  AND U47596 ( .A(n47597), .B(n47598), .Z(n47596) );
  XOR U47597 ( .A(n47595), .B(n47269), .Z(n47597) );
  XOR U47598 ( .A(n47599), .B(n47600), .Z(n47233) );
  AND U47599 ( .A(n1150), .B(n47582), .Z(n47600) );
  XNOR U47600 ( .A(n47580), .B(n47599), .Z(n47582) );
  XNOR U47601 ( .A(n47601), .B(n47602), .Z(n1150) );
  AND U47602 ( .A(n47603), .B(n47604), .Z(n47602) );
  XNOR U47603 ( .A(n47605), .B(n47601), .Z(n47604) );
  IV U47604 ( .A(n47292), .Z(n47605) );
  XOR U47605 ( .A(n47563), .B(n47606), .Z(n47292) );
  AND U47606 ( .A(n1153), .B(n47607), .Z(n47606) );
  XOR U47607 ( .A(n47345), .B(n47342), .Z(n47607) );
  IV U47608 ( .A(n47563), .Z(n47345) );
  XNOR U47609 ( .A(n47242), .B(n47601), .Z(n47603) );
  XOR U47610 ( .A(n47608), .B(n47609), .Z(n47242) );
  AND U47611 ( .A(n1169), .B(n47610), .Z(n47609) );
  XOR U47612 ( .A(n47611), .B(n47612), .Z(n47601) );
  AND U47613 ( .A(n47613), .B(n47614), .Z(n47612) );
  XNOR U47614 ( .A(n47611), .B(n47302), .Z(n47614) );
  XOR U47615 ( .A(n47362), .B(n47615), .Z(n47302) );
  AND U47616 ( .A(n1153), .B(n47616), .Z(n47615) );
  XOR U47617 ( .A(n47358), .B(n47362), .Z(n47616) );
  XNOR U47618 ( .A(n47617), .B(n47611), .Z(n47613) );
  IV U47619 ( .A(n47252), .Z(n47617) );
  XOR U47620 ( .A(n47618), .B(n47619), .Z(n47252) );
  AND U47621 ( .A(n1169), .B(n47620), .Z(n47619) );
  XOR U47622 ( .A(n47621), .B(n47622), .Z(n47611) );
  AND U47623 ( .A(n47623), .B(n47624), .Z(n47622) );
  XNOR U47624 ( .A(n47621), .B(n47312), .Z(n47624) );
  XOR U47625 ( .A(n47390), .B(n47625), .Z(n47312) );
  AND U47626 ( .A(n1153), .B(n47626), .Z(n47625) );
  XOR U47627 ( .A(n47386), .B(n47390), .Z(n47626) );
  XOR U47628 ( .A(n47261), .B(n47621), .Z(n47623) );
  XOR U47629 ( .A(n47627), .B(n47628), .Z(n47261) );
  AND U47630 ( .A(n1169), .B(n47629), .Z(n47628) );
  XOR U47631 ( .A(n47595), .B(n47630), .Z(n47621) );
  AND U47632 ( .A(n47631), .B(n47598), .Z(n47630) );
  XNOR U47633 ( .A(n47322), .B(n47595), .Z(n47598) );
  XOR U47634 ( .A(n47439), .B(n47632), .Z(n47322) );
  AND U47635 ( .A(n1153), .B(n47633), .Z(n47632) );
  XOR U47636 ( .A(n47435), .B(n47439), .Z(n47633) );
  XNOR U47637 ( .A(n47634), .B(n47595), .Z(n47631) );
  IV U47638 ( .A(n47269), .Z(n47634) );
  XOR U47639 ( .A(n47635), .B(n47636), .Z(n47269) );
  AND U47640 ( .A(n1169), .B(n47637), .Z(n47636) );
  XOR U47641 ( .A(n47638), .B(n47639), .Z(n47595) );
  AND U47642 ( .A(n47640), .B(n47641), .Z(n47639) );
  XNOR U47643 ( .A(n47638), .B(n47330), .Z(n47641) );
  XOR U47644 ( .A(n47536), .B(n47642), .Z(n47330) );
  AND U47645 ( .A(n1153), .B(n47643), .Z(n47642) );
  XOR U47646 ( .A(n47532), .B(n47536), .Z(n47643) );
  XNOR U47647 ( .A(n47644), .B(n47638), .Z(n47640) );
  IV U47648 ( .A(n47279), .Z(n47644) );
  XOR U47649 ( .A(n47645), .B(n47646), .Z(n47279) );
  AND U47650 ( .A(n1169), .B(n47647), .Z(n47646) );
  AND U47651 ( .A(n47599), .B(n47580), .Z(n47638) );
  XNOR U47652 ( .A(n47648), .B(n47649), .Z(n47580) );
  AND U47653 ( .A(n1153), .B(n47558), .Z(n47649) );
  XNOR U47654 ( .A(n47556), .B(n47648), .Z(n47558) );
  XNOR U47655 ( .A(n47650), .B(n47651), .Z(n1153) );
  AND U47656 ( .A(n47652), .B(n47653), .Z(n47651) );
  XNOR U47657 ( .A(n47650), .B(n47342), .Z(n47653) );
  IV U47658 ( .A(n47346), .Z(n47342) );
  XOR U47659 ( .A(n47654), .B(n47655), .Z(n47346) );
  AND U47660 ( .A(n1157), .B(n47656), .Z(n47655) );
  XOR U47661 ( .A(n47657), .B(n47654), .Z(n47656) );
  XNOR U47662 ( .A(n47650), .B(n47563), .Z(n47652) );
  XOR U47663 ( .A(n47658), .B(n47659), .Z(n47563) );
  AND U47664 ( .A(n1165), .B(n47610), .Z(n47659) );
  XOR U47665 ( .A(n47608), .B(n47658), .Z(n47610) );
  XOR U47666 ( .A(n47660), .B(n47661), .Z(n47650) );
  AND U47667 ( .A(n47662), .B(n47663), .Z(n47661) );
  XNOR U47668 ( .A(n47660), .B(n47358), .Z(n47663) );
  IV U47669 ( .A(n47361), .Z(n47358) );
  XOR U47670 ( .A(n47664), .B(n47665), .Z(n47361) );
  AND U47671 ( .A(n1157), .B(n47666), .Z(n47665) );
  XOR U47672 ( .A(n47667), .B(n47664), .Z(n47666) );
  XOR U47673 ( .A(n47362), .B(n47660), .Z(n47662) );
  XOR U47674 ( .A(n47668), .B(n47669), .Z(n47362) );
  AND U47675 ( .A(n1165), .B(n47620), .Z(n47669) );
  XOR U47676 ( .A(n47668), .B(n47618), .Z(n47620) );
  XOR U47677 ( .A(n47670), .B(n47671), .Z(n47660) );
  AND U47678 ( .A(n47672), .B(n47673), .Z(n47671) );
  XNOR U47679 ( .A(n47670), .B(n47386), .Z(n47673) );
  IV U47680 ( .A(n47389), .Z(n47386) );
  XOR U47681 ( .A(n47674), .B(n47675), .Z(n47389) );
  AND U47682 ( .A(n1157), .B(n47676), .Z(n47675) );
  XNOR U47683 ( .A(n47677), .B(n47674), .Z(n47676) );
  XOR U47684 ( .A(n47390), .B(n47670), .Z(n47672) );
  XOR U47685 ( .A(n47678), .B(n47679), .Z(n47390) );
  AND U47686 ( .A(n1165), .B(n47629), .Z(n47679) );
  XOR U47687 ( .A(n47678), .B(n47627), .Z(n47629) );
  XOR U47688 ( .A(n47680), .B(n47681), .Z(n47670) );
  AND U47689 ( .A(n47682), .B(n47683), .Z(n47681) );
  XNOR U47690 ( .A(n47680), .B(n47435), .Z(n47683) );
  IV U47691 ( .A(n47438), .Z(n47435) );
  XOR U47692 ( .A(n47684), .B(n47685), .Z(n47438) );
  AND U47693 ( .A(n1157), .B(n47686), .Z(n47685) );
  XOR U47694 ( .A(n47687), .B(n47684), .Z(n47686) );
  XOR U47695 ( .A(n47439), .B(n47680), .Z(n47682) );
  XOR U47696 ( .A(n47688), .B(n47689), .Z(n47439) );
  AND U47697 ( .A(n1165), .B(n47637), .Z(n47689) );
  XOR U47698 ( .A(n47688), .B(n47635), .Z(n47637) );
  XOR U47699 ( .A(n47576), .B(n47690), .Z(n47680) );
  AND U47700 ( .A(n47578), .B(n47691), .Z(n47690) );
  XNOR U47701 ( .A(n47576), .B(n47532), .Z(n47691) );
  IV U47702 ( .A(n47535), .Z(n47532) );
  XOR U47703 ( .A(n47692), .B(n47693), .Z(n47535) );
  AND U47704 ( .A(n1157), .B(n47694), .Z(n47693) );
  XNOR U47705 ( .A(n47695), .B(n47692), .Z(n47694) );
  XOR U47706 ( .A(n47536), .B(n47576), .Z(n47578) );
  XOR U47707 ( .A(n47696), .B(n47697), .Z(n47536) );
  AND U47708 ( .A(n1165), .B(n47647), .Z(n47697) );
  XOR U47709 ( .A(n47696), .B(n47645), .Z(n47647) );
  AND U47710 ( .A(n47648), .B(n47556), .Z(n47576) );
  XNOR U47711 ( .A(n47698), .B(n47699), .Z(n47556) );
  AND U47712 ( .A(n1157), .B(n47700), .Z(n47699) );
  XNOR U47713 ( .A(n47701), .B(n47698), .Z(n47700) );
  XNOR U47714 ( .A(n47702), .B(n47703), .Z(n1157) );
  AND U47715 ( .A(n47704), .B(n47705), .Z(n47703) );
  XOR U47716 ( .A(n47657), .B(n47702), .Z(n47705) );
  AND U47717 ( .A(n47706), .B(n47707), .Z(n47657) );
  XNOR U47718 ( .A(n47654), .B(n47702), .Z(n47704) );
  XNOR U47719 ( .A(n47708), .B(n47709), .Z(n47654) );
  AND U47720 ( .A(n1161), .B(n47710), .Z(n47709) );
  XNOR U47721 ( .A(n47711), .B(n47712), .Z(n47710) );
  XOR U47722 ( .A(n47713), .B(n47714), .Z(n47702) );
  AND U47723 ( .A(n47715), .B(n47716), .Z(n47714) );
  XNOR U47724 ( .A(n47713), .B(n47706), .Z(n47716) );
  IV U47725 ( .A(n47667), .Z(n47706) );
  XOR U47726 ( .A(n47717), .B(n47718), .Z(n47667) );
  XOR U47727 ( .A(n47719), .B(n47707), .Z(n47718) );
  AND U47728 ( .A(n47677), .B(n47720), .Z(n47707) );
  AND U47729 ( .A(n47721), .B(n47722), .Z(n47719) );
  XOR U47730 ( .A(n47723), .B(n47717), .Z(n47721) );
  XNOR U47731 ( .A(n47664), .B(n47713), .Z(n47715) );
  XNOR U47732 ( .A(n47724), .B(n47725), .Z(n47664) );
  AND U47733 ( .A(n1161), .B(n47726), .Z(n47725) );
  XNOR U47734 ( .A(n47727), .B(n47728), .Z(n47726) );
  XOR U47735 ( .A(n47729), .B(n47730), .Z(n47713) );
  AND U47736 ( .A(n47731), .B(n47732), .Z(n47730) );
  XNOR U47737 ( .A(n47729), .B(n47677), .Z(n47732) );
  XOR U47738 ( .A(n47733), .B(n47722), .Z(n47677) );
  XNOR U47739 ( .A(n47734), .B(n47717), .Z(n47722) );
  XOR U47740 ( .A(n47735), .B(n47736), .Z(n47717) );
  AND U47741 ( .A(n47737), .B(n47738), .Z(n47736) );
  XOR U47742 ( .A(n47739), .B(n47735), .Z(n47737) );
  XNOR U47743 ( .A(n47740), .B(n47741), .Z(n47734) );
  AND U47744 ( .A(n47742), .B(n47743), .Z(n47741) );
  XOR U47745 ( .A(n47740), .B(n47744), .Z(n47742) );
  XNOR U47746 ( .A(n47723), .B(n47720), .Z(n47733) );
  AND U47747 ( .A(n47745), .B(n47746), .Z(n47720) );
  XOR U47748 ( .A(n47747), .B(n47748), .Z(n47723) );
  AND U47749 ( .A(n47749), .B(n47750), .Z(n47748) );
  XOR U47750 ( .A(n47747), .B(n47751), .Z(n47749) );
  XNOR U47751 ( .A(n47674), .B(n47729), .Z(n47731) );
  XNOR U47752 ( .A(n47752), .B(n47753), .Z(n47674) );
  AND U47753 ( .A(n1161), .B(n47754), .Z(n47753) );
  XNOR U47754 ( .A(n47755), .B(n47756), .Z(n47754) );
  XOR U47755 ( .A(n47757), .B(n47758), .Z(n47729) );
  AND U47756 ( .A(n47759), .B(n47760), .Z(n47758) );
  XNOR U47757 ( .A(n47757), .B(n47745), .Z(n47760) );
  IV U47758 ( .A(n47687), .Z(n47745) );
  XNOR U47759 ( .A(n47761), .B(n47738), .Z(n47687) );
  XNOR U47760 ( .A(n47762), .B(n47744), .Z(n47738) );
  XOR U47761 ( .A(n47763), .B(n47764), .Z(n47744) );
  AND U47762 ( .A(n47765), .B(n47766), .Z(n47764) );
  XOR U47763 ( .A(n47763), .B(n47767), .Z(n47765) );
  XNOR U47764 ( .A(n47743), .B(n47735), .Z(n47762) );
  XOR U47765 ( .A(n47768), .B(n47769), .Z(n47735) );
  AND U47766 ( .A(n47770), .B(n47771), .Z(n47769) );
  XNOR U47767 ( .A(n47772), .B(n47768), .Z(n47770) );
  XNOR U47768 ( .A(n47773), .B(n47740), .Z(n47743) );
  XOR U47769 ( .A(n47774), .B(n47775), .Z(n47740) );
  AND U47770 ( .A(n47776), .B(n47777), .Z(n47775) );
  XOR U47771 ( .A(n47774), .B(n47778), .Z(n47776) );
  XNOR U47772 ( .A(n47779), .B(n47780), .Z(n47773) );
  AND U47773 ( .A(n47781), .B(n47782), .Z(n47780) );
  XNOR U47774 ( .A(n47779), .B(n47783), .Z(n47781) );
  XNOR U47775 ( .A(n47739), .B(n47746), .Z(n47761) );
  AND U47776 ( .A(n47695), .B(n47784), .Z(n47746) );
  XOR U47777 ( .A(n47751), .B(n47750), .Z(n47739) );
  XNOR U47778 ( .A(n47785), .B(n47747), .Z(n47750) );
  XOR U47779 ( .A(n47786), .B(n47787), .Z(n47747) );
  AND U47780 ( .A(n47788), .B(n47789), .Z(n47787) );
  XOR U47781 ( .A(n47786), .B(n47790), .Z(n47788) );
  XNOR U47782 ( .A(n47791), .B(n47792), .Z(n47785) );
  AND U47783 ( .A(n47793), .B(n47794), .Z(n47792) );
  XOR U47784 ( .A(n47791), .B(n47795), .Z(n47793) );
  XOR U47785 ( .A(n47796), .B(n47797), .Z(n47751) );
  AND U47786 ( .A(n47798), .B(n47799), .Z(n47797) );
  XOR U47787 ( .A(n47796), .B(n47800), .Z(n47798) );
  XNOR U47788 ( .A(n47684), .B(n47757), .Z(n47759) );
  XNOR U47789 ( .A(n47801), .B(n47802), .Z(n47684) );
  AND U47790 ( .A(n1161), .B(n47803), .Z(n47802) );
  XNOR U47791 ( .A(n47804), .B(n47805), .Z(n47803) );
  XOR U47792 ( .A(n47806), .B(n47807), .Z(n47757) );
  AND U47793 ( .A(n47808), .B(n47809), .Z(n47807) );
  XNOR U47794 ( .A(n47806), .B(n47695), .Z(n47809) );
  XOR U47795 ( .A(n47810), .B(n47771), .Z(n47695) );
  XNOR U47796 ( .A(n47811), .B(n47778), .Z(n47771) );
  XOR U47797 ( .A(n47767), .B(n47766), .Z(n47778) );
  XNOR U47798 ( .A(n47812), .B(n47763), .Z(n47766) );
  XOR U47799 ( .A(n47813), .B(n47814), .Z(n47763) );
  AND U47800 ( .A(n47815), .B(n47816), .Z(n47814) );
  XNOR U47801 ( .A(n47817), .B(n47818), .Z(n47815) );
  IV U47802 ( .A(n47813), .Z(n47817) );
  XNOR U47803 ( .A(n47819), .B(n47820), .Z(n47812) );
  NOR U47804 ( .A(n47821), .B(n47822), .Z(n47820) );
  XNOR U47805 ( .A(n47819), .B(n47823), .Z(n47821) );
  XOR U47806 ( .A(n47824), .B(n47825), .Z(n47767) );
  NOR U47807 ( .A(n47826), .B(n47827), .Z(n47825) );
  XNOR U47808 ( .A(n47824), .B(n47828), .Z(n47826) );
  XNOR U47809 ( .A(n47777), .B(n47768), .Z(n47811) );
  XOR U47810 ( .A(n47829), .B(n47830), .Z(n47768) );
  AND U47811 ( .A(n47831), .B(n47832), .Z(n47830) );
  XOR U47812 ( .A(n47829), .B(n47833), .Z(n47831) );
  XOR U47813 ( .A(n47834), .B(n47783), .Z(n47777) );
  XOR U47814 ( .A(n47835), .B(n47836), .Z(n47783) );
  NOR U47815 ( .A(n47837), .B(n47838), .Z(n47836) );
  XOR U47816 ( .A(n47835), .B(n47839), .Z(n47837) );
  XNOR U47817 ( .A(n47782), .B(n47774), .Z(n47834) );
  XOR U47818 ( .A(n47840), .B(n47841), .Z(n47774) );
  AND U47819 ( .A(n47842), .B(n47843), .Z(n47841) );
  XOR U47820 ( .A(n47840), .B(n47844), .Z(n47842) );
  XNOR U47821 ( .A(n47845), .B(n47779), .Z(n47782) );
  XOR U47822 ( .A(n47846), .B(n47847), .Z(n47779) );
  AND U47823 ( .A(n47848), .B(n47849), .Z(n47847) );
  XNOR U47824 ( .A(n47850), .B(n47851), .Z(n47848) );
  IV U47825 ( .A(n47846), .Z(n47850) );
  XNOR U47826 ( .A(n47852), .B(n47853), .Z(n47845) );
  NOR U47827 ( .A(n47854), .B(n47855), .Z(n47853) );
  XNOR U47828 ( .A(n47852), .B(n47856), .Z(n47854) );
  XOR U47829 ( .A(n47772), .B(n47784), .Z(n47810) );
  NOR U47830 ( .A(n47701), .B(n47857), .Z(n47784) );
  XNOR U47831 ( .A(n47790), .B(n47789), .Z(n47772) );
  XNOR U47832 ( .A(n47858), .B(n47795), .Z(n47789) );
  XNOR U47833 ( .A(n47859), .B(n47860), .Z(n47795) );
  NOR U47834 ( .A(n47861), .B(n47862), .Z(n47860) );
  XOR U47835 ( .A(n47859), .B(n47863), .Z(n47861) );
  XNOR U47836 ( .A(n47794), .B(n47786), .Z(n47858) );
  XOR U47837 ( .A(n47864), .B(n47865), .Z(n47786) );
  AND U47838 ( .A(n47866), .B(n47867), .Z(n47865) );
  XOR U47839 ( .A(n47864), .B(n47868), .Z(n47866) );
  XNOR U47840 ( .A(n47869), .B(n47791), .Z(n47794) );
  XOR U47841 ( .A(n47870), .B(n47871), .Z(n47791) );
  AND U47842 ( .A(n47872), .B(n47873), .Z(n47871) );
  XNOR U47843 ( .A(n47874), .B(n47875), .Z(n47872) );
  IV U47844 ( .A(n47870), .Z(n47874) );
  XNOR U47845 ( .A(n47876), .B(n47877), .Z(n47869) );
  NOR U47846 ( .A(n47878), .B(n47879), .Z(n47877) );
  XNOR U47847 ( .A(n47876), .B(n47880), .Z(n47878) );
  XOR U47848 ( .A(n47800), .B(n47799), .Z(n47790) );
  XNOR U47849 ( .A(n47881), .B(n47796), .Z(n47799) );
  XOR U47850 ( .A(n47882), .B(n47883), .Z(n47796) );
  AND U47851 ( .A(n47884), .B(n47885), .Z(n47883) );
  XNOR U47852 ( .A(n47886), .B(n47887), .Z(n47884) );
  IV U47853 ( .A(n47882), .Z(n47886) );
  XNOR U47854 ( .A(n47888), .B(n47889), .Z(n47881) );
  NOR U47855 ( .A(n47890), .B(n47891), .Z(n47889) );
  XNOR U47856 ( .A(n47888), .B(n47892), .Z(n47890) );
  XOR U47857 ( .A(n47893), .B(n47894), .Z(n47800) );
  NOR U47858 ( .A(n47895), .B(n47896), .Z(n47894) );
  XNOR U47859 ( .A(n47893), .B(n47897), .Z(n47895) );
  XNOR U47860 ( .A(n47692), .B(n47806), .Z(n47808) );
  XNOR U47861 ( .A(n47898), .B(n47899), .Z(n47692) );
  AND U47862 ( .A(n1161), .B(n47900), .Z(n47899) );
  XNOR U47863 ( .A(n47901), .B(n47902), .Z(n47900) );
  AND U47864 ( .A(n47698), .B(n47701), .Z(n47806) );
  XOR U47865 ( .A(n47903), .B(n47857), .Z(n47701) );
  XNOR U47866 ( .A(p_input[1728]), .B(p_input[2048]), .Z(n47857) );
  XNOR U47867 ( .A(n47833), .B(n47832), .Z(n47903) );
  XNOR U47868 ( .A(n47904), .B(n47844), .Z(n47832) );
  XOR U47869 ( .A(n47818), .B(n47816), .Z(n47844) );
  XNOR U47870 ( .A(n47905), .B(n47823), .Z(n47816) );
  XOR U47871 ( .A(p_input[1752]), .B(p_input[2072]), .Z(n47823) );
  XOR U47872 ( .A(n47813), .B(n47822), .Z(n47905) );
  XOR U47873 ( .A(n47906), .B(n47819), .Z(n47822) );
  XOR U47874 ( .A(p_input[1750]), .B(p_input[2070]), .Z(n47819) );
  XOR U47875 ( .A(p_input[1751]), .B(n29410), .Z(n47906) );
  XOR U47876 ( .A(p_input[1746]), .B(p_input[2066]), .Z(n47813) );
  XNOR U47877 ( .A(n47828), .B(n47827), .Z(n47818) );
  XOR U47878 ( .A(n47907), .B(n47824), .Z(n47827) );
  XOR U47879 ( .A(p_input[1747]), .B(p_input[2067]), .Z(n47824) );
  XOR U47880 ( .A(p_input[1748]), .B(n29412), .Z(n47907) );
  XOR U47881 ( .A(p_input[1749]), .B(p_input[2069]), .Z(n47828) );
  XOR U47882 ( .A(n47843), .B(n47908), .Z(n47904) );
  IV U47883 ( .A(n47829), .Z(n47908) );
  XOR U47884 ( .A(p_input[1729]), .B(p_input[2049]), .Z(n47829) );
  XNOR U47885 ( .A(n47909), .B(n47851), .Z(n47843) );
  XNOR U47886 ( .A(n47839), .B(n47838), .Z(n47851) );
  XNOR U47887 ( .A(n47910), .B(n47835), .Z(n47838) );
  XNOR U47888 ( .A(p_input[1754]), .B(p_input[2074]), .Z(n47835) );
  XOR U47889 ( .A(p_input[1755]), .B(n29415), .Z(n47910) );
  XOR U47890 ( .A(p_input[1756]), .B(p_input[2076]), .Z(n47839) );
  XOR U47891 ( .A(n47849), .B(n47911), .Z(n47909) );
  IV U47892 ( .A(n47840), .Z(n47911) );
  XOR U47893 ( .A(p_input[1745]), .B(p_input[2065]), .Z(n47840) );
  XNOR U47894 ( .A(n47912), .B(n47856), .Z(n47849) );
  XNOR U47895 ( .A(p_input[1759]), .B(n29418), .Z(n47856) );
  XOR U47896 ( .A(n47846), .B(n47855), .Z(n47912) );
  XOR U47897 ( .A(n47913), .B(n47852), .Z(n47855) );
  XOR U47898 ( .A(p_input[1757]), .B(p_input[2077]), .Z(n47852) );
  XOR U47899 ( .A(p_input[1758]), .B(n29420), .Z(n47913) );
  XOR U47900 ( .A(p_input[1753]), .B(p_input[2073]), .Z(n47846) );
  XOR U47901 ( .A(n47868), .B(n47867), .Z(n47833) );
  XNOR U47902 ( .A(n47914), .B(n47875), .Z(n47867) );
  XNOR U47903 ( .A(n47863), .B(n47862), .Z(n47875) );
  XNOR U47904 ( .A(n47915), .B(n47859), .Z(n47862) );
  XNOR U47905 ( .A(p_input[1739]), .B(p_input[2059]), .Z(n47859) );
  XOR U47906 ( .A(p_input[1740]), .B(n28329), .Z(n47915) );
  XOR U47907 ( .A(p_input[1741]), .B(p_input[2061]), .Z(n47863) );
  XOR U47908 ( .A(n47873), .B(n47916), .Z(n47914) );
  IV U47909 ( .A(n47864), .Z(n47916) );
  XOR U47910 ( .A(p_input[1730]), .B(p_input[2050]), .Z(n47864) );
  XNOR U47911 ( .A(n47917), .B(n47880), .Z(n47873) );
  XNOR U47912 ( .A(p_input[1744]), .B(n28332), .Z(n47880) );
  XOR U47913 ( .A(n47870), .B(n47879), .Z(n47917) );
  XOR U47914 ( .A(n47918), .B(n47876), .Z(n47879) );
  XOR U47915 ( .A(p_input[1742]), .B(p_input[2062]), .Z(n47876) );
  XOR U47916 ( .A(p_input[1743]), .B(n28334), .Z(n47918) );
  XOR U47917 ( .A(p_input[1738]), .B(p_input[2058]), .Z(n47870) );
  XOR U47918 ( .A(n47887), .B(n47885), .Z(n47868) );
  XNOR U47919 ( .A(n47919), .B(n47892), .Z(n47885) );
  XOR U47920 ( .A(p_input[1737]), .B(p_input[2057]), .Z(n47892) );
  XOR U47921 ( .A(n47882), .B(n47891), .Z(n47919) );
  XOR U47922 ( .A(n47920), .B(n47888), .Z(n47891) );
  XOR U47923 ( .A(p_input[1735]), .B(p_input[2055]), .Z(n47888) );
  XOR U47924 ( .A(p_input[1736]), .B(n29427), .Z(n47920) );
  XOR U47925 ( .A(p_input[1731]), .B(p_input[2051]), .Z(n47882) );
  XNOR U47926 ( .A(n47897), .B(n47896), .Z(n47887) );
  XOR U47927 ( .A(n47921), .B(n47893), .Z(n47896) );
  XOR U47928 ( .A(p_input[1732]), .B(p_input[2052]), .Z(n47893) );
  XOR U47929 ( .A(p_input[1733]), .B(n29429), .Z(n47921) );
  XOR U47930 ( .A(p_input[1734]), .B(p_input[2054]), .Z(n47897) );
  XNOR U47931 ( .A(n47922), .B(n47923), .Z(n47698) );
  AND U47932 ( .A(n1161), .B(n47924), .Z(n47923) );
  XNOR U47933 ( .A(n47925), .B(n47926), .Z(n1161) );
  AND U47934 ( .A(n47927), .B(n47928), .Z(n47926) );
  XOR U47935 ( .A(n47712), .B(n47925), .Z(n47928) );
  XNOR U47936 ( .A(n47929), .B(n47925), .Z(n47927) );
  XOR U47937 ( .A(n47930), .B(n47931), .Z(n47925) );
  AND U47938 ( .A(n47932), .B(n47933), .Z(n47931) );
  XOR U47939 ( .A(n47727), .B(n47930), .Z(n47933) );
  XOR U47940 ( .A(n47930), .B(n47728), .Z(n47932) );
  XOR U47941 ( .A(n47934), .B(n47935), .Z(n47930) );
  AND U47942 ( .A(n47936), .B(n47937), .Z(n47935) );
  XOR U47943 ( .A(n47755), .B(n47934), .Z(n47937) );
  XOR U47944 ( .A(n47934), .B(n47756), .Z(n47936) );
  XOR U47945 ( .A(n47938), .B(n47939), .Z(n47934) );
  AND U47946 ( .A(n47940), .B(n47941), .Z(n47939) );
  XOR U47947 ( .A(n47804), .B(n47938), .Z(n47941) );
  XOR U47948 ( .A(n47938), .B(n47805), .Z(n47940) );
  XOR U47949 ( .A(n47942), .B(n47943), .Z(n47938) );
  AND U47950 ( .A(n47944), .B(n47945), .Z(n47943) );
  XOR U47951 ( .A(n47942), .B(n47901), .Z(n47945) );
  XNOR U47952 ( .A(n47946), .B(n47947), .Z(n47648) );
  AND U47953 ( .A(n1165), .B(n47948), .Z(n47947) );
  XNOR U47954 ( .A(n47949), .B(n47950), .Z(n1165) );
  AND U47955 ( .A(n47951), .B(n47952), .Z(n47950) );
  XOR U47956 ( .A(n47949), .B(n47658), .Z(n47952) );
  XNOR U47957 ( .A(n47949), .B(n47608), .Z(n47951) );
  XOR U47958 ( .A(n47953), .B(n47954), .Z(n47949) );
  AND U47959 ( .A(n47955), .B(n47956), .Z(n47954) );
  XNOR U47960 ( .A(n47668), .B(n47953), .Z(n47956) );
  XOR U47961 ( .A(n47953), .B(n47618), .Z(n47955) );
  XOR U47962 ( .A(n47957), .B(n47958), .Z(n47953) );
  AND U47963 ( .A(n47959), .B(n47960), .Z(n47958) );
  XNOR U47964 ( .A(n47678), .B(n47957), .Z(n47960) );
  XOR U47965 ( .A(n47957), .B(n47627), .Z(n47959) );
  XOR U47966 ( .A(n47961), .B(n47962), .Z(n47957) );
  AND U47967 ( .A(n47963), .B(n47964), .Z(n47962) );
  XOR U47968 ( .A(n47961), .B(n47635), .Z(n47963) );
  XOR U47969 ( .A(n47965), .B(n47966), .Z(n47599) );
  AND U47970 ( .A(n1169), .B(n47948), .Z(n47966) );
  XNOR U47971 ( .A(n47946), .B(n47965), .Z(n47948) );
  XNOR U47972 ( .A(n47967), .B(n47968), .Z(n1169) );
  AND U47973 ( .A(n47969), .B(n47970), .Z(n47968) );
  XNOR U47974 ( .A(n47971), .B(n47967), .Z(n47970) );
  IV U47975 ( .A(n47658), .Z(n47971) );
  XOR U47976 ( .A(n47929), .B(n47972), .Z(n47658) );
  AND U47977 ( .A(n1172), .B(n47973), .Z(n47972) );
  XOR U47978 ( .A(n47711), .B(n47708), .Z(n47973) );
  IV U47979 ( .A(n47929), .Z(n47711) );
  XNOR U47980 ( .A(n47608), .B(n47967), .Z(n47969) );
  XOR U47981 ( .A(n47974), .B(n47975), .Z(n47608) );
  AND U47982 ( .A(n1188), .B(n47976), .Z(n47975) );
  XOR U47983 ( .A(n47977), .B(n47978), .Z(n47967) );
  AND U47984 ( .A(n47979), .B(n47980), .Z(n47978) );
  XNOR U47985 ( .A(n47977), .B(n47668), .Z(n47980) );
  XOR U47986 ( .A(n47728), .B(n47981), .Z(n47668) );
  AND U47987 ( .A(n1172), .B(n47982), .Z(n47981) );
  XOR U47988 ( .A(n47724), .B(n47728), .Z(n47982) );
  XNOR U47989 ( .A(n47983), .B(n47977), .Z(n47979) );
  IV U47990 ( .A(n47618), .Z(n47983) );
  XOR U47991 ( .A(n47984), .B(n47985), .Z(n47618) );
  AND U47992 ( .A(n1188), .B(n47986), .Z(n47985) );
  XOR U47993 ( .A(n47987), .B(n47988), .Z(n47977) );
  AND U47994 ( .A(n47989), .B(n47990), .Z(n47988) );
  XNOR U47995 ( .A(n47987), .B(n47678), .Z(n47990) );
  XOR U47996 ( .A(n47756), .B(n47991), .Z(n47678) );
  AND U47997 ( .A(n1172), .B(n47992), .Z(n47991) );
  XOR U47998 ( .A(n47752), .B(n47756), .Z(n47992) );
  XOR U47999 ( .A(n47627), .B(n47987), .Z(n47989) );
  XOR U48000 ( .A(n47993), .B(n47994), .Z(n47627) );
  AND U48001 ( .A(n1188), .B(n47995), .Z(n47994) );
  XOR U48002 ( .A(n47961), .B(n47996), .Z(n47987) );
  AND U48003 ( .A(n47997), .B(n47964), .Z(n47996) );
  XNOR U48004 ( .A(n47688), .B(n47961), .Z(n47964) );
  XOR U48005 ( .A(n47805), .B(n47998), .Z(n47688) );
  AND U48006 ( .A(n1172), .B(n47999), .Z(n47998) );
  XOR U48007 ( .A(n47801), .B(n47805), .Z(n47999) );
  XNOR U48008 ( .A(n48000), .B(n47961), .Z(n47997) );
  IV U48009 ( .A(n47635), .Z(n48000) );
  XOR U48010 ( .A(n48001), .B(n48002), .Z(n47635) );
  AND U48011 ( .A(n1188), .B(n48003), .Z(n48002) );
  XOR U48012 ( .A(n48004), .B(n48005), .Z(n47961) );
  AND U48013 ( .A(n48006), .B(n48007), .Z(n48005) );
  XNOR U48014 ( .A(n48004), .B(n47696), .Z(n48007) );
  XOR U48015 ( .A(n47902), .B(n48008), .Z(n47696) );
  AND U48016 ( .A(n1172), .B(n48009), .Z(n48008) );
  XOR U48017 ( .A(n47898), .B(n47902), .Z(n48009) );
  XNOR U48018 ( .A(n48010), .B(n48004), .Z(n48006) );
  IV U48019 ( .A(n47645), .Z(n48010) );
  XOR U48020 ( .A(n48011), .B(n48012), .Z(n47645) );
  AND U48021 ( .A(n1188), .B(n48013), .Z(n48012) );
  AND U48022 ( .A(n47965), .B(n47946), .Z(n48004) );
  XNOR U48023 ( .A(n48014), .B(n48015), .Z(n47946) );
  AND U48024 ( .A(n1172), .B(n47924), .Z(n48015) );
  XNOR U48025 ( .A(n47922), .B(n48014), .Z(n47924) );
  XNOR U48026 ( .A(n48016), .B(n48017), .Z(n1172) );
  AND U48027 ( .A(n48018), .B(n48019), .Z(n48017) );
  XNOR U48028 ( .A(n48016), .B(n47708), .Z(n48019) );
  IV U48029 ( .A(n47712), .Z(n47708) );
  XOR U48030 ( .A(n48020), .B(n48021), .Z(n47712) );
  AND U48031 ( .A(n1176), .B(n48022), .Z(n48021) );
  XOR U48032 ( .A(n48023), .B(n48020), .Z(n48022) );
  XNOR U48033 ( .A(n48016), .B(n47929), .Z(n48018) );
  XOR U48034 ( .A(n48024), .B(n48025), .Z(n47929) );
  AND U48035 ( .A(n1184), .B(n47976), .Z(n48025) );
  XOR U48036 ( .A(n47974), .B(n48024), .Z(n47976) );
  XOR U48037 ( .A(n48026), .B(n48027), .Z(n48016) );
  AND U48038 ( .A(n48028), .B(n48029), .Z(n48027) );
  XNOR U48039 ( .A(n48026), .B(n47724), .Z(n48029) );
  IV U48040 ( .A(n47727), .Z(n47724) );
  XOR U48041 ( .A(n48030), .B(n48031), .Z(n47727) );
  AND U48042 ( .A(n1176), .B(n48032), .Z(n48031) );
  XOR U48043 ( .A(n48033), .B(n48030), .Z(n48032) );
  XOR U48044 ( .A(n47728), .B(n48026), .Z(n48028) );
  XOR U48045 ( .A(n48034), .B(n48035), .Z(n47728) );
  AND U48046 ( .A(n1184), .B(n47986), .Z(n48035) );
  XOR U48047 ( .A(n48034), .B(n47984), .Z(n47986) );
  XOR U48048 ( .A(n48036), .B(n48037), .Z(n48026) );
  AND U48049 ( .A(n48038), .B(n48039), .Z(n48037) );
  XNOR U48050 ( .A(n48036), .B(n47752), .Z(n48039) );
  IV U48051 ( .A(n47755), .Z(n47752) );
  XOR U48052 ( .A(n48040), .B(n48041), .Z(n47755) );
  AND U48053 ( .A(n1176), .B(n48042), .Z(n48041) );
  XNOR U48054 ( .A(n48043), .B(n48040), .Z(n48042) );
  XOR U48055 ( .A(n47756), .B(n48036), .Z(n48038) );
  XOR U48056 ( .A(n48044), .B(n48045), .Z(n47756) );
  AND U48057 ( .A(n1184), .B(n47995), .Z(n48045) );
  XOR U48058 ( .A(n48044), .B(n47993), .Z(n47995) );
  XOR U48059 ( .A(n48046), .B(n48047), .Z(n48036) );
  AND U48060 ( .A(n48048), .B(n48049), .Z(n48047) );
  XNOR U48061 ( .A(n48046), .B(n47801), .Z(n48049) );
  IV U48062 ( .A(n47804), .Z(n47801) );
  XOR U48063 ( .A(n48050), .B(n48051), .Z(n47804) );
  AND U48064 ( .A(n1176), .B(n48052), .Z(n48051) );
  XOR U48065 ( .A(n48053), .B(n48050), .Z(n48052) );
  XOR U48066 ( .A(n47805), .B(n48046), .Z(n48048) );
  XOR U48067 ( .A(n48054), .B(n48055), .Z(n47805) );
  AND U48068 ( .A(n1184), .B(n48003), .Z(n48055) );
  XOR U48069 ( .A(n48054), .B(n48001), .Z(n48003) );
  XOR U48070 ( .A(n47942), .B(n48056), .Z(n48046) );
  AND U48071 ( .A(n47944), .B(n48057), .Z(n48056) );
  XNOR U48072 ( .A(n47942), .B(n47898), .Z(n48057) );
  IV U48073 ( .A(n47901), .Z(n47898) );
  XOR U48074 ( .A(n48058), .B(n48059), .Z(n47901) );
  AND U48075 ( .A(n1176), .B(n48060), .Z(n48059) );
  XNOR U48076 ( .A(n48061), .B(n48058), .Z(n48060) );
  XOR U48077 ( .A(n47902), .B(n47942), .Z(n47944) );
  XOR U48078 ( .A(n48062), .B(n48063), .Z(n47902) );
  AND U48079 ( .A(n1184), .B(n48013), .Z(n48063) );
  XOR U48080 ( .A(n48062), .B(n48011), .Z(n48013) );
  AND U48081 ( .A(n48014), .B(n47922), .Z(n47942) );
  XNOR U48082 ( .A(n48064), .B(n48065), .Z(n47922) );
  AND U48083 ( .A(n1176), .B(n48066), .Z(n48065) );
  XNOR U48084 ( .A(n48067), .B(n48064), .Z(n48066) );
  XNOR U48085 ( .A(n48068), .B(n48069), .Z(n1176) );
  AND U48086 ( .A(n48070), .B(n48071), .Z(n48069) );
  XOR U48087 ( .A(n48023), .B(n48068), .Z(n48071) );
  AND U48088 ( .A(n48072), .B(n48073), .Z(n48023) );
  XNOR U48089 ( .A(n48020), .B(n48068), .Z(n48070) );
  XNOR U48090 ( .A(n48074), .B(n48075), .Z(n48020) );
  AND U48091 ( .A(n1180), .B(n48076), .Z(n48075) );
  XNOR U48092 ( .A(n48077), .B(n48078), .Z(n48076) );
  XOR U48093 ( .A(n48079), .B(n48080), .Z(n48068) );
  AND U48094 ( .A(n48081), .B(n48082), .Z(n48080) );
  XNOR U48095 ( .A(n48079), .B(n48072), .Z(n48082) );
  IV U48096 ( .A(n48033), .Z(n48072) );
  XOR U48097 ( .A(n48083), .B(n48084), .Z(n48033) );
  XOR U48098 ( .A(n48085), .B(n48073), .Z(n48084) );
  AND U48099 ( .A(n48043), .B(n48086), .Z(n48073) );
  AND U48100 ( .A(n48087), .B(n48088), .Z(n48085) );
  XOR U48101 ( .A(n48089), .B(n48083), .Z(n48087) );
  XNOR U48102 ( .A(n48030), .B(n48079), .Z(n48081) );
  XNOR U48103 ( .A(n48090), .B(n48091), .Z(n48030) );
  AND U48104 ( .A(n1180), .B(n48092), .Z(n48091) );
  XNOR U48105 ( .A(n48093), .B(n48094), .Z(n48092) );
  XOR U48106 ( .A(n48095), .B(n48096), .Z(n48079) );
  AND U48107 ( .A(n48097), .B(n48098), .Z(n48096) );
  XNOR U48108 ( .A(n48095), .B(n48043), .Z(n48098) );
  XOR U48109 ( .A(n48099), .B(n48088), .Z(n48043) );
  XNOR U48110 ( .A(n48100), .B(n48083), .Z(n48088) );
  XOR U48111 ( .A(n48101), .B(n48102), .Z(n48083) );
  AND U48112 ( .A(n48103), .B(n48104), .Z(n48102) );
  XOR U48113 ( .A(n48105), .B(n48101), .Z(n48103) );
  XNOR U48114 ( .A(n48106), .B(n48107), .Z(n48100) );
  AND U48115 ( .A(n48108), .B(n48109), .Z(n48107) );
  XOR U48116 ( .A(n48106), .B(n48110), .Z(n48108) );
  XNOR U48117 ( .A(n48089), .B(n48086), .Z(n48099) );
  AND U48118 ( .A(n48111), .B(n48112), .Z(n48086) );
  XOR U48119 ( .A(n48113), .B(n48114), .Z(n48089) );
  AND U48120 ( .A(n48115), .B(n48116), .Z(n48114) );
  XOR U48121 ( .A(n48113), .B(n48117), .Z(n48115) );
  XNOR U48122 ( .A(n48040), .B(n48095), .Z(n48097) );
  XNOR U48123 ( .A(n48118), .B(n48119), .Z(n48040) );
  AND U48124 ( .A(n1180), .B(n48120), .Z(n48119) );
  XNOR U48125 ( .A(n48121), .B(n48122), .Z(n48120) );
  XOR U48126 ( .A(n48123), .B(n48124), .Z(n48095) );
  AND U48127 ( .A(n48125), .B(n48126), .Z(n48124) );
  XNOR U48128 ( .A(n48123), .B(n48111), .Z(n48126) );
  IV U48129 ( .A(n48053), .Z(n48111) );
  XNOR U48130 ( .A(n48127), .B(n48104), .Z(n48053) );
  XNOR U48131 ( .A(n48128), .B(n48110), .Z(n48104) );
  XOR U48132 ( .A(n48129), .B(n48130), .Z(n48110) );
  AND U48133 ( .A(n48131), .B(n48132), .Z(n48130) );
  XOR U48134 ( .A(n48129), .B(n48133), .Z(n48131) );
  XNOR U48135 ( .A(n48109), .B(n48101), .Z(n48128) );
  XOR U48136 ( .A(n48134), .B(n48135), .Z(n48101) );
  AND U48137 ( .A(n48136), .B(n48137), .Z(n48135) );
  XNOR U48138 ( .A(n48138), .B(n48134), .Z(n48136) );
  XNOR U48139 ( .A(n48139), .B(n48106), .Z(n48109) );
  XOR U48140 ( .A(n48140), .B(n48141), .Z(n48106) );
  AND U48141 ( .A(n48142), .B(n48143), .Z(n48141) );
  XOR U48142 ( .A(n48140), .B(n48144), .Z(n48142) );
  XNOR U48143 ( .A(n48145), .B(n48146), .Z(n48139) );
  AND U48144 ( .A(n48147), .B(n48148), .Z(n48146) );
  XNOR U48145 ( .A(n48145), .B(n48149), .Z(n48147) );
  XNOR U48146 ( .A(n48105), .B(n48112), .Z(n48127) );
  AND U48147 ( .A(n48061), .B(n48150), .Z(n48112) );
  XOR U48148 ( .A(n48117), .B(n48116), .Z(n48105) );
  XNOR U48149 ( .A(n48151), .B(n48113), .Z(n48116) );
  XOR U48150 ( .A(n48152), .B(n48153), .Z(n48113) );
  AND U48151 ( .A(n48154), .B(n48155), .Z(n48153) );
  XOR U48152 ( .A(n48152), .B(n48156), .Z(n48154) );
  XNOR U48153 ( .A(n48157), .B(n48158), .Z(n48151) );
  AND U48154 ( .A(n48159), .B(n48160), .Z(n48158) );
  XOR U48155 ( .A(n48157), .B(n48161), .Z(n48159) );
  XOR U48156 ( .A(n48162), .B(n48163), .Z(n48117) );
  AND U48157 ( .A(n48164), .B(n48165), .Z(n48163) );
  XOR U48158 ( .A(n48162), .B(n48166), .Z(n48164) );
  XNOR U48159 ( .A(n48050), .B(n48123), .Z(n48125) );
  XNOR U48160 ( .A(n48167), .B(n48168), .Z(n48050) );
  AND U48161 ( .A(n1180), .B(n48169), .Z(n48168) );
  XNOR U48162 ( .A(n48170), .B(n48171), .Z(n48169) );
  XOR U48163 ( .A(n48172), .B(n48173), .Z(n48123) );
  AND U48164 ( .A(n48174), .B(n48175), .Z(n48173) );
  XNOR U48165 ( .A(n48172), .B(n48061), .Z(n48175) );
  XOR U48166 ( .A(n48176), .B(n48137), .Z(n48061) );
  XNOR U48167 ( .A(n48177), .B(n48144), .Z(n48137) );
  XOR U48168 ( .A(n48133), .B(n48132), .Z(n48144) );
  XNOR U48169 ( .A(n48178), .B(n48129), .Z(n48132) );
  XOR U48170 ( .A(n48179), .B(n48180), .Z(n48129) );
  AND U48171 ( .A(n48181), .B(n48182), .Z(n48180) );
  XNOR U48172 ( .A(n48183), .B(n48184), .Z(n48181) );
  IV U48173 ( .A(n48179), .Z(n48183) );
  XNOR U48174 ( .A(n48185), .B(n48186), .Z(n48178) );
  NOR U48175 ( .A(n48187), .B(n48188), .Z(n48186) );
  XNOR U48176 ( .A(n48185), .B(n48189), .Z(n48187) );
  XOR U48177 ( .A(n48190), .B(n48191), .Z(n48133) );
  NOR U48178 ( .A(n48192), .B(n48193), .Z(n48191) );
  XNOR U48179 ( .A(n48190), .B(n48194), .Z(n48192) );
  XNOR U48180 ( .A(n48143), .B(n48134), .Z(n48177) );
  XOR U48181 ( .A(n48195), .B(n48196), .Z(n48134) );
  AND U48182 ( .A(n48197), .B(n48198), .Z(n48196) );
  XOR U48183 ( .A(n48195), .B(n48199), .Z(n48197) );
  XOR U48184 ( .A(n48200), .B(n48149), .Z(n48143) );
  XOR U48185 ( .A(n48201), .B(n48202), .Z(n48149) );
  NOR U48186 ( .A(n48203), .B(n48204), .Z(n48202) );
  XOR U48187 ( .A(n48201), .B(n48205), .Z(n48203) );
  XNOR U48188 ( .A(n48148), .B(n48140), .Z(n48200) );
  XOR U48189 ( .A(n48206), .B(n48207), .Z(n48140) );
  AND U48190 ( .A(n48208), .B(n48209), .Z(n48207) );
  XOR U48191 ( .A(n48206), .B(n48210), .Z(n48208) );
  XNOR U48192 ( .A(n48211), .B(n48145), .Z(n48148) );
  XOR U48193 ( .A(n48212), .B(n48213), .Z(n48145) );
  AND U48194 ( .A(n48214), .B(n48215), .Z(n48213) );
  XNOR U48195 ( .A(n48216), .B(n48217), .Z(n48214) );
  IV U48196 ( .A(n48212), .Z(n48216) );
  XNOR U48197 ( .A(n48218), .B(n48219), .Z(n48211) );
  NOR U48198 ( .A(n48220), .B(n48221), .Z(n48219) );
  XNOR U48199 ( .A(n48218), .B(n48222), .Z(n48220) );
  XOR U48200 ( .A(n48138), .B(n48150), .Z(n48176) );
  NOR U48201 ( .A(n48067), .B(n48223), .Z(n48150) );
  XNOR U48202 ( .A(n48156), .B(n48155), .Z(n48138) );
  XNOR U48203 ( .A(n48224), .B(n48161), .Z(n48155) );
  XNOR U48204 ( .A(n48225), .B(n48226), .Z(n48161) );
  NOR U48205 ( .A(n48227), .B(n48228), .Z(n48226) );
  XOR U48206 ( .A(n48225), .B(n48229), .Z(n48227) );
  XNOR U48207 ( .A(n48160), .B(n48152), .Z(n48224) );
  XOR U48208 ( .A(n48230), .B(n48231), .Z(n48152) );
  AND U48209 ( .A(n48232), .B(n48233), .Z(n48231) );
  XOR U48210 ( .A(n48230), .B(n48234), .Z(n48232) );
  XNOR U48211 ( .A(n48235), .B(n48157), .Z(n48160) );
  XOR U48212 ( .A(n48236), .B(n48237), .Z(n48157) );
  AND U48213 ( .A(n48238), .B(n48239), .Z(n48237) );
  XNOR U48214 ( .A(n48240), .B(n48241), .Z(n48238) );
  IV U48215 ( .A(n48236), .Z(n48240) );
  XNOR U48216 ( .A(n48242), .B(n48243), .Z(n48235) );
  NOR U48217 ( .A(n48244), .B(n48245), .Z(n48243) );
  XNOR U48218 ( .A(n48242), .B(n48246), .Z(n48244) );
  XOR U48219 ( .A(n48166), .B(n48165), .Z(n48156) );
  XNOR U48220 ( .A(n48247), .B(n48162), .Z(n48165) );
  XOR U48221 ( .A(n48248), .B(n48249), .Z(n48162) );
  AND U48222 ( .A(n48250), .B(n48251), .Z(n48249) );
  XNOR U48223 ( .A(n48252), .B(n48253), .Z(n48250) );
  IV U48224 ( .A(n48248), .Z(n48252) );
  XNOR U48225 ( .A(n48254), .B(n48255), .Z(n48247) );
  NOR U48226 ( .A(n48256), .B(n48257), .Z(n48255) );
  XNOR U48227 ( .A(n48254), .B(n48258), .Z(n48256) );
  XOR U48228 ( .A(n48259), .B(n48260), .Z(n48166) );
  NOR U48229 ( .A(n48261), .B(n48262), .Z(n48260) );
  XNOR U48230 ( .A(n48259), .B(n48263), .Z(n48261) );
  XNOR U48231 ( .A(n48058), .B(n48172), .Z(n48174) );
  XNOR U48232 ( .A(n48264), .B(n48265), .Z(n48058) );
  AND U48233 ( .A(n1180), .B(n48266), .Z(n48265) );
  XNOR U48234 ( .A(n48267), .B(n48268), .Z(n48266) );
  AND U48235 ( .A(n48064), .B(n48067), .Z(n48172) );
  XOR U48236 ( .A(n48269), .B(n48223), .Z(n48067) );
  XNOR U48237 ( .A(p_input[1760]), .B(p_input[2048]), .Z(n48223) );
  XNOR U48238 ( .A(n48199), .B(n48198), .Z(n48269) );
  XNOR U48239 ( .A(n48270), .B(n48210), .Z(n48198) );
  XOR U48240 ( .A(n48184), .B(n48182), .Z(n48210) );
  XNOR U48241 ( .A(n48271), .B(n48189), .Z(n48182) );
  XOR U48242 ( .A(p_input[1784]), .B(p_input[2072]), .Z(n48189) );
  XOR U48243 ( .A(n48179), .B(n48188), .Z(n48271) );
  XOR U48244 ( .A(n48272), .B(n48185), .Z(n48188) );
  XOR U48245 ( .A(p_input[1782]), .B(p_input[2070]), .Z(n48185) );
  XOR U48246 ( .A(p_input[1783]), .B(n29410), .Z(n48272) );
  XOR U48247 ( .A(p_input[1778]), .B(p_input[2066]), .Z(n48179) );
  XNOR U48248 ( .A(n48194), .B(n48193), .Z(n48184) );
  XOR U48249 ( .A(n48273), .B(n48190), .Z(n48193) );
  XOR U48250 ( .A(p_input[1779]), .B(p_input[2067]), .Z(n48190) );
  XOR U48251 ( .A(p_input[1780]), .B(n29412), .Z(n48273) );
  XOR U48252 ( .A(p_input[1781]), .B(p_input[2069]), .Z(n48194) );
  XOR U48253 ( .A(n48209), .B(n48274), .Z(n48270) );
  IV U48254 ( .A(n48195), .Z(n48274) );
  XOR U48255 ( .A(p_input[1761]), .B(p_input[2049]), .Z(n48195) );
  XNOR U48256 ( .A(n48275), .B(n48217), .Z(n48209) );
  XNOR U48257 ( .A(n48205), .B(n48204), .Z(n48217) );
  XNOR U48258 ( .A(n48276), .B(n48201), .Z(n48204) );
  XNOR U48259 ( .A(p_input[1786]), .B(p_input[2074]), .Z(n48201) );
  XOR U48260 ( .A(p_input[1787]), .B(n29415), .Z(n48276) );
  XOR U48261 ( .A(p_input[1788]), .B(p_input[2076]), .Z(n48205) );
  XOR U48262 ( .A(n48215), .B(n48277), .Z(n48275) );
  IV U48263 ( .A(n48206), .Z(n48277) );
  XOR U48264 ( .A(p_input[1777]), .B(p_input[2065]), .Z(n48206) );
  XNOR U48265 ( .A(n48278), .B(n48222), .Z(n48215) );
  XNOR U48266 ( .A(p_input[1791]), .B(n29418), .Z(n48222) );
  XOR U48267 ( .A(n48212), .B(n48221), .Z(n48278) );
  XOR U48268 ( .A(n48279), .B(n48218), .Z(n48221) );
  XOR U48269 ( .A(p_input[1789]), .B(p_input[2077]), .Z(n48218) );
  XOR U48270 ( .A(p_input[1790]), .B(n29420), .Z(n48279) );
  XOR U48271 ( .A(p_input[1785]), .B(p_input[2073]), .Z(n48212) );
  XOR U48272 ( .A(n48234), .B(n48233), .Z(n48199) );
  XNOR U48273 ( .A(n48280), .B(n48241), .Z(n48233) );
  XNOR U48274 ( .A(n48229), .B(n48228), .Z(n48241) );
  XNOR U48275 ( .A(n48281), .B(n48225), .Z(n48228) );
  XNOR U48276 ( .A(p_input[1771]), .B(p_input[2059]), .Z(n48225) );
  XOR U48277 ( .A(p_input[1772]), .B(n28329), .Z(n48281) );
  XOR U48278 ( .A(p_input[1773]), .B(p_input[2061]), .Z(n48229) );
  XOR U48279 ( .A(n48239), .B(n48282), .Z(n48280) );
  IV U48280 ( .A(n48230), .Z(n48282) );
  XOR U48281 ( .A(p_input[1762]), .B(p_input[2050]), .Z(n48230) );
  XNOR U48282 ( .A(n48283), .B(n48246), .Z(n48239) );
  XNOR U48283 ( .A(p_input[1776]), .B(n28332), .Z(n48246) );
  XOR U48284 ( .A(n48236), .B(n48245), .Z(n48283) );
  XOR U48285 ( .A(n48284), .B(n48242), .Z(n48245) );
  XOR U48286 ( .A(p_input[1774]), .B(p_input[2062]), .Z(n48242) );
  XOR U48287 ( .A(p_input[1775]), .B(n28334), .Z(n48284) );
  XOR U48288 ( .A(p_input[1770]), .B(p_input[2058]), .Z(n48236) );
  XOR U48289 ( .A(n48253), .B(n48251), .Z(n48234) );
  XNOR U48290 ( .A(n48285), .B(n48258), .Z(n48251) );
  XOR U48291 ( .A(p_input[1769]), .B(p_input[2057]), .Z(n48258) );
  XOR U48292 ( .A(n48248), .B(n48257), .Z(n48285) );
  XOR U48293 ( .A(n48286), .B(n48254), .Z(n48257) );
  XOR U48294 ( .A(p_input[1767]), .B(p_input[2055]), .Z(n48254) );
  XOR U48295 ( .A(p_input[1768]), .B(n29427), .Z(n48286) );
  XOR U48296 ( .A(p_input[1763]), .B(p_input[2051]), .Z(n48248) );
  XNOR U48297 ( .A(n48263), .B(n48262), .Z(n48253) );
  XOR U48298 ( .A(n48287), .B(n48259), .Z(n48262) );
  XOR U48299 ( .A(p_input[1764]), .B(p_input[2052]), .Z(n48259) );
  XOR U48300 ( .A(p_input[1765]), .B(n29429), .Z(n48287) );
  XOR U48301 ( .A(p_input[1766]), .B(p_input[2054]), .Z(n48263) );
  XNOR U48302 ( .A(n48288), .B(n48289), .Z(n48064) );
  AND U48303 ( .A(n1180), .B(n48290), .Z(n48289) );
  XNOR U48304 ( .A(n48291), .B(n48292), .Z(n1180) );
  AND U48305 ( .A(n48293), .B(n48294), .Z(n48292) );
  XOR U48306 ( .A(n48078), .B(n48291), .Z(n48294) );
  XNOR U48307 ( .A(n48295), .B(n48291), .Z(n48293) );
  XOR U48308 ( .A(n48296), .B(n48297), .Z(n48291) );
  AND U48309 ( .A(n48298), .B(n48299), .Z(n48297) );
  XOR U48310 ( .A(n48093), .B(n48296), .Z(n48299) );
  XOR U48311 ( .A(n48296), .B(n48094), .Z(n48298) );
  XOR U48312 ( .A(n48300), .B(n48301), .Z(n48296) );
  AND U48313 ( .A(n48302), .B(n48303), .Z(n48301) );
  XOR U48314 ( .A(n48121), .B(n48300), .Z(n48303) );
  XOR U48315 ( .A(n48300), .B(n48122), .Z(n48302) );
  XOR U48316 ( .A(n48304), .B(n48305), .Z(n48300) );
  AND U48317 ( .A(n48306), .B(n48307), .Z(n48305) );
  XOR U48318 ( .A(n48170), .B(n48304), .Z(n48307) );
  XOR U48319 ( .A(n48304), .B(n48171), .Z(n48306) );
  XOR U48320 ( .A(n48308), .B(n48309), .Z(n48304) );
  AND U48321 ( .A(n48310), .B(n48311), .Z(n48309) );
  XOR U48322 ( .A(n48308), .B(n48267), .Z(n48311) );
  XNOR U48323 ( .A(n48312), .B(n48313), .Z(n48014) );
  AND U48324 ( .A(n1184), .B(n48314), .Z(n48313) );
  XNOR U48325 ( .A(n48315), .B(n48316), .Z(n1184) );
  AND U48326 ( .A(n48317), .B(n48318), .Z(n48316) );
  XOR U48327 ( .A(n48315), .B(n48024), .Z(n48318) );
  XNOR U48328 ( .A(n48315), .B(n47974), .Z(n48317) );
  XOR U48329 ( .A(n48319), .B(n48320), .Z(n48315) );
  AND U48330 ( .A(n48321), .B(n48322), .Z(n48320) );
  XNOR U48331 ( .A(n48034), .B(n48319), .Z(n48322) );
  XOR U48332 ( .A(n48319), .B(n47984), .Z(n48321) );
  XOR U48333 ( .A(n48323), .B(n48324), .Z(n48319) );
  AND U48334 ( .A(n48325), .B(n48326), .Z(n48324) );
  XNOR U48335 ( .A(n48044), .B(n48323), .Z(n48326) );
  XOR U48336 ( .A(n48323), .B(n47993), .Z(n48325) );
  XOR U48337 ( .A(n48327), .B(n48328), .Z(n48323) );
  AND U48338 ( .A(n48329), .B(n48330), .Z(n48328) );
  XOR U48339 ( .A(n48327), .B(n48001), .Z(n48329) );
  XOR U48340 ( .A(n48331), .B(n48332), .Z(n47965) );
  AND U48341 ( .A(n1188), .B(n48314), .Z(n48332) );
  XNOR U48342 ( .A(n48312), .B(n48331), .Z(n48314) );
  XNOR U48343 ( .A(n48333), .B(n48334), .Z(n1188) );
  AND U48344 ( .A(n48335), .B(n48336), .Z(n48334) );
  XNOR U48345 ( .A(n48337), .B(n48333), .Z(n48336) );
  IV U48346 ( .A(n48024), .Z(n48337) );
  XOR U48347 ( .A(n48295), .B(n48338), .Z(n48024) );
  AND U48348 ( .A(n1191), .B(n48339), .Z(n48338) );
  XOR U48349 ( .A(n48077), .B(n48074), .Z(n48339) );
  IV U48350 ( .A(n48295), .Z(n48077) );
  XNOR U48351 ( .A(n47974), .B(n48333), .Z(n48335) );
  XOR U48352 ( .A(n48340), .B(n48341), .Z(n47974) );
  AND U48353 ( .A(n1207), .B(n48342), .Z(n48341) );
  XOR U48354 ( .A(n48343), .B(n48344), .Z(n48333) );
  AND U48355 ( .A(n48345), .B(n48346), .Z(n48344) );
  XNOR U48356 ( .A(n48343), .B(n48034), .Z(n48346) );
  XOR U48357 ( .A(n48094), .B(n48347), .Z(n48034) );
  AND U48358 ( .A(n1191), .B(n48348), .Z(n48347) );
  XOR U48359 ( .A(n48090), .B(n48094), .Z(n48348) );
  XNOR U48360 ( .A(n48349), .B(n48343), .Z(n48345) );
  IV U48361 ( .A(n47984), .Z(n48349) );
  XOR U48362 ( .A(n48350), .B(n48351), .Z(n47984) );
  AND U48363 ( .A(n1207), .B(n48352), .Z(n48351) );
  XOR U48364 ( .A(n48353), .B(n48354), .Z(n48343) );
  AND U48365 ( .A(n48355), .B(n48356), .Z(n48354) );
  XNOR U48366 ( .A(n48353), .B(n48044), .Z(n48356) );
  XOR U48367 ( .A(n48122), .B(n48357), .Z(n48044) );
  AND U48368 ( .A(n1191), .B(n48358), .Z(n48357) );
  XOR U48369 ( .A(n48118), .B(n48122), .Z(n48358) );
  XOR U48370 ( .A(n47993), .B(n48353), .Z(n48355) );
  XOR U48371 ( .A(n48359), .B(n48360), .Z(n47993) );
  AND U48372 ( .A(n1207), .B(n48361), .Z(n48360) );
  XOR U48373 ( .A(n48327), .B(n48362), .Z(n48353) );
  AND U48374 ( .A(n48363), .B(n48330), .Z(n48362) );
  XNOR U48375 ( .A(n48054), .B(n48327), .Z(n48330) );
  XOR U48376 ( .A(n48171), .B(n48364), .Z(n48054) );
  AND U48377 ( .A(n1191), .B(n48365), .Z(n48364) );
  XOR U48378 ( .A(n48167), .B(n48171), .Z(n48365) );
  XNOR U48379 ( .A(n48366), .B(n48327), .Z(n48363) );
  IV U48380 ( .A(n48001), .Z(n48366) );
  XOR U48381 ( .A(n48367), .B(n48368), .Z(n48001) );
  AND U48382 ( .A(n1207), .B(n48369), .Z(n48368) );
  XOR U48383 ( .A(n48370), .B(n48371), .Z(n48327) );
  AND U48384 ( .A(n48372), .B(n48373), .Z(n48371) );
  XNOR U48385 ( .A(n48370), .B(n48062), .Z(n48373) );
  XOR U48386 ( .A(n48268), .B(n48374), .Z(n48062) );
  AND U48387 ( .A(n1191), .B(n48375), .Z(n48374) );
  XOR U48388 ( .A(n48264), .B(n48268), .Z(n48375) );
  XNOR U48389 ( .A(n48376), .B(n48370), .Z(n48372) );
  IV U48390 ( .A(n48011), .Z(n48376) );
  XOR U48391 ( .A(n48377), .B(n48378), .Z(n48011) );
  AND U48392 ( .A(n1207), .B(n48379), .Z(n48378) );
  AND U48393 ( .A(n48331), .B(n48312), .Z(n48370) );
  XNOR U48394 ( .A(n48380), .B(n48381), .Z(n48312) );
  AND U48395 ( .A(n1191), .B(n48290), .Z(n48381) );
  XNOR U48396 ( .A(n48288), .B(n48380), .Z(n48290) );
  XNOR U48397 ( .A(n48382), .B(n48383), .Z(n1191) );
  AND U48398 ( .A(n48384), .B(n48385), .Z(n48383) );
  XNOR U48399 ( .A(n48382), .B(n48074), .Z(n48385) );
  IV U48400 ( .A(n48078), .Z(n48074) );
  XOR U48401 ( .A(n48386), .B(n48387), .Z(n48078) );
  AND U48402 ( .A(n1195), .B(n48388), .Z(n48387) );
  XOR U48403 ( .A(n48389), .B(n48386), .Z(n48388) );
  XNOR U48404 ( .A(n48382), .B(n48295), .Z(n48384) );
  XOR U48405 ( .A(n48390), .B(n48391), .Z(n48295) );
  AND U48406 ( .A(n1203), .B(n48342), .Z(n48391) );
  XOR U48407 ( .A(n48340), .B(n48390), .Z(n48342) );
  XOR U48408 ( .A(n48392), .B(n48393), .Z(n48382) );
  AND U48409 ( .A(n48394), .B(n48395), .Z(n48393) );
  XNOR U48410 ( .A(n48392), .B(n48090), .Z(n48395) );
  IV U48411 ( .A(n48093), .Z(n48090) );
  XOR U48412 ( .A(n48396), .B(n48397), .Z(n48093) );
  AND U48413 ( .A(n1195), .B(n48398), .Z(n48397) );
  XOR U48414 ( .A(n48399), .B(n48396), .Z(n48398) );
  XOR U48415 ( .A(n48094), .B(n48392), .Z(n48394) );
  XOR U48416 ( .A(n48400), .B(n48401), .Z(n48094) );
  AND U48417 ( .A(n1203), .B(n48352), .Z(n48401) );
  XOR U48418 ( .A(n48400), .B(n48350), .Z(n48352) );
  XOR U48419 ( .A(n48402), .B(n48403), .Z(n48392) );
  AND U48420 ( .A(n48404), .B(n48405), .Z(n48403) );
  XNOR U48421 ( .A(n48402), .B(n48118), .Z(n48405) );
  IV U48422 ( .A(n48121), .Z(n48118) );
  XOR U48423 ( .A(n48406), .B(n48407), .Z(n48121) );
  AND U48424 ( .A(n1195), .B(n48408), .Z(n48407) );
  XNOR U48425 ( .A(n48409), .B(n48406), .Z(n48408) );
  XOR U48426 ( .A(n48122), .B(n48402), .Z(n48404) );
  XOR U48427 ( .A(n48410), .B(n48411), .Z(n48122) );
  AND U48428 ( .A(n1203), .B(n48361), .Z(n48411) );
  XOR U48429 ( .A(n48410), .B(n48359), .Z(n48361) );
  XOR U48430 ( .A(n48412), .B(n48413), .Z(n48402) );
  AND U48431 ( .A(n48414), .B(n48415), .Z(n48413) );
  XNOR U48432 ( .A(n48412), .B(n48167), .Z(n48415) );
  IV U48433 ( .A(n48170), .Z(n48167) );
  XOR U48434 ( .A(n48416), .B(n48417), .Z(n48170) );
  AND U48435 ( .A(n1195), .B(n48418), .Z(n48417) );
  XOR U48436 ( .A(n48419), .B(n48416), .Z(n48418) );
  XOR U48437 ( .A(n48171), .B(n48412), .Z(n48414) );
  XOR U48438 ( .A(n48420), .B(n48421), .Z(n48171) );
  AND U48439 ( .A(n1203), .B(n48369), .Z(n48421) );
  XOR U48440 ( .A(n48420), .B(n48367), .Z(n48369) );
  XOR U48441 ( .A(n48308), .B(n48422), .Z(n48412) );
  AND U48442 ( .A(n48310), .B(n48423), .Z(n48422) );
  XNOR U48443 ( .A(n48308), .B(n48264), .Z(n48423) );
  IV U48444 ( .A(n48267), .Z(n48264) );
  XOR U48445 ( .A(n48424), .B(n48425), .Z(n48267) );
  AND U48446 ( .A(n1195), .B(n48426), .Z(n48425) );
  XNOR U48447 ( .A(n48427), .B(n48424), .Z(n48426) );
  XOR U48448 ( .A(n48268), .B(n48308), .Z(n48310) );
  XOR U48449 ( .A(n48428), .B(n48429), .Z(n48268) );
  AND U48450 ( .A(n1203), .B(n48379), .Z(n48429) );
  XOR U48451 ( .A(n48428), .B(n48377), .Z(n48379) );
  AND U48452 ( .A(n48380), .B(n48288), .Z(n48308) );
  XNOR U48453 ( .A(n48430), .B(n48431), .Z(n48288) );
  AND U48454 ( .A(n1195), .B(n48432), .Z(n48431) );
  XNOR U48455 ( .A(n48433), .B(n48430), .Z(n48432) );
  XNOR U48456 ( .A(n48434), .B(n48435), .Z(n1195) );
  AND U48457 ( .A(n48436), .B(n48437), .Z(n48435) );
  XOR U48458 ( .A(n48389), .B(n48434), .Z(n48437) );
  AND U48459 ( .A(n48438), .B(n48439), .Z(n48389) );
  XNOR U48460 ( .A(n48386), .B(n48434), .Z(n48436) );
  XNOR U48461 ( .A(n48440), .B(n48441), .Z(n48386) );
  AND U48462 ( .A(n1199), .B(n48442), .Z(n48441) );
  XNOR U48463 ( .A(n48443), .B(n48444), .Z(n48442) );
  XOR U48464 ( .A(n48445), .B(n48446), .Z(n48434) );
  AND U48465 ( .A(n48447), .B(n48448), .Z(n48446) );
  XNOR U48466 ( .A(n48445), .B(n48438), .Z(n48448) );
  IV U48467 ( .A(n48399), .Z(n48438) );
  XOR U48468 ( .A(n48449), .B(n48450), .Z(n48399) );
  XOR U48469 ( .A(n48451), .B(n48439), .Z(n48450) );
  AND U48470 ( .A(n48409), .B(n48452), .Z(n48439) );
  AND U48471 ( .A(n48453), .B(n48454), .Z(n48451) );
  XOR U48472 ( .A(n48455), .B(n48449), .Z(n48453) );
  XNOR U48473 ( .A(n48396), .B(n48445), .Z(n48447) );
  XNOR U48474 ( .A(n48456), .B(n48457), .Z(n48396) );
  AND U48475 ( .A(n1199), .B(n48458), .Z(n48457) );
  XNOR U48476 ( .A(n48459), .B(n48460), .Z(n48458) );
  XOR U48477 ( .A(n48461), .B(n48462), .Z(n48445) );
  AND U48478 ( .A(n48463), .B(n48464), .Z(n48462) );
  XNOR U48479 ( .A(n48461), .B(n48409), .Z(n48464) );
  XOR U48480 ( .A(n48465), .B(n48454), .Z(n48409) );
  XNOR U48481 ( .A(n48466), .B(n48449), .Z(n48454) );
  XOR U48482 ( .A(n48467), .B(n48468), .Z(n48449) );
  AND U48483 ( .A(n48469), .B(n48470), .Z(n48468) );
  XOR U48484 ( .A(n48471), .B(n48467), .Z(n48469) );
  XNOR U48485 ( .A(n48472), .B(n48473), .Z(n48466) );
  AND U48486 ( .A(n48474), .B(n48475), .Z(n48473) );
  XOR U48487 ( .A(n48472), .B(n48476), .Z(n48474) );
  XNOR U48488 ( .A(n48455), .B(n48452), .Z(n48465) );
  AND U48489 ( .A(n48477), .B(n48478), .Z(n48452) );
  XOR U48490 ( .A(n48479), .B(n48480), .Z(n48455) );
  AND U48491 ( .A(n48481), .B(n48482), .Z(n48480) );
  XOR U48492 ( .A(n48479), .B(n48483), .Z(n48481) );
  XNOR U48493 ( .A(n48406), .B(n48461), .Z(n48463) );
  XNOR U48494 ( .A(n48484), .B(n48485), .Z(n48406) );
  AND U48495 ( .A(n1199), .B(n48486), .Z(n48485) );
  XNOR U48496 ( .A(n48487), .B(n48488), .Z(n48486) );
  XOR U48497 ( .A(n48489), .B(n48490), .Z(n48461) );
  AND U48498 ( .A(n48491), .B(n48492), .Z(n48490) );
  XNOR U48499 ( .A(n48489), .B(n48477), .Z(n48492) );
  IV U48500 ( .A(n48419), .Z(n48477) );
  XNOR U48501 ( .A(n48493), .B(n48470), .Z(n48419) );
  XNOR U48502 ( .A(n48494), .B(n48476), .Z(n48470) );
  XOR U48503 ( .A(n48495), .B(n48496), .Z(n48476) );
  AND U48504 ( .A(n48497), .B(n48498), .Z(n48496) );
  XOR U48505 ( .A(n48495), .B(n48499), .Z(n48497) );
  XNOR U48506 ( .A(n48475), .B(n48467), .Z(n48494) );
  XOR U48507 ( .A(n48500), .B(n48501), .Z(n48467) );
  AND U48508 ( .A(n48502), .B(n48503), .Z(n48501) );
  XNOR U48509 ( .A(n48504), .B(n48500), .Z(n48502) );
  XNOR U48510 ( .A(n48505), .B(n48472), .Z(n48475) );
  XOR U48511 ( .A(n48506), .B(n48507), .Z(n48472) );
  AND U48512 ( .A(n48508), .B(n48509), .Z(n48507) );
  XOR U48513 ( .A(n48506), .B(n48510), .Z(n48508) );
  XNOR U48514 ( .A(n48511), .B(n48512), .Z(n48505) );
  AND U48515 ( .A(n48513), .B(n48514), .Z(n48512) );
  XNOR U48516 ( .A(n48511), .B(n48515), .Z(n48513) );
  XNOR U48517 ( .A(n48471), .B(n48478), .Z(n48493) );
  AND U48518 ( .A(n48427), .B(n48516), .Z(n48478) );
  XOR U48519 ( .A(n48483), .B(n48482), .Z(n48471) );
  XNOR U48520 ( .A(n48517), .B(n48479), .Z(n48482) );
  XOR U48521 ( .A(n48518), .B(n48519), .Z(n48479) );
  AND U48522 ( .A(n48520), .B(n48521), .Z(n48519) );
  XOR U48523 ( .A(n48518), .B(n48522), .Z(n48520) );
  XNOR U48524 ( .A(n48523), .B(n48524), .Z(n48517) );
  AND U48525 ( .A(n48525), .B(n48526), .Z(n48524) );
  XOR U48526 ( .A(n48523), .B(n48527), .Z(n48525) );
  XOR U48527 ( .A(n48528), .B(n48529), .Z(n48483) );
  AND U48528 ( .A(n48530), .B(n48531), .Z(n48529) );
  XOR U48529 ( .A(n48528), .B(n48532), .Z(n48530) );
  XNOR U48530 ( .A(n48416), .B(n48489), .Z(n48491) );
  XNOR U48531 ( .A(n48533), .B(n48534), .Z(n48416) );
  AND U48532 ( .A(n1199), .B(n48535), .Z(n48534) );
  XNOR U48533 ( .A(n48536), .B(n48537), .Z(n48535) );
  XOR U48534 ( .A(n48538), .B(n48539), .Z(n48489) );
  AND U48535 ( .A(n48540), .B(n48541), .Z(n48539) );
  XNOR U48536 ( .A(n48538), .B(n48427), .Z(n48541) );
  XOR U48537 ( .A(n48542), .B(n48503), .Z(n48427) );
  XNOR U48538 ( .A(n48543), .B(n48510), .Z(n48503) );
  XOR U48539 ( .A(n48499), .B(n48498), .Z(n48510) );
  XNOR U48540 ( .A(n48544), .B(n48495), .Z(n48498) );
  XOR U48541 ( .A(n48545), .B(n48546), .Z(n48495) );
  AND U48542 ( .A(n48547), .B(n48548), .Z(n48546) );
  XNOR U48543 ( .A(n48549), .B(n48550), .Z(n48547) );
  IV U48544 ( .A(n48545), .Z(n48549) );
  XNOR U48545 ( .A(n48551), .B(n48552), .Z(n48544) );
  NOR U48546 ( .A(n48553), .B(n48554), .Z(n48552) );
  XNOR U48547 ( .A(n48551), .B(n48555), .Z(n48553) );
  XOR U48548 ( .A(n48556), .B(n48557), .Z(n48499) );
  NOR U48549 ( .A(n48558), .B(n48559), .Z(n48557) );
  XNOR U48550 ( .A(n48556), .B(n48560), .Z(n48558) );
  XNOR U48551 ( .A(n48509), .B(n48500), .Z(n48543) );
  XOR U48552 ( .A(n48561), .B(n48562), .Z(n48500) );
  AND U48553 ( .A(n48563), .B(n48564), .Z(n48562) );
  XOR U48554 ( .A(n48561), .B(n48565), .Z(n48563) );
  XOR U48555 ( .A(n48566), .B(n48515), .Z(n48509) );
  XOR U48556 ( .A(n48567), .B(n48568), .Z(n48515) );
  NOR U48557 ( .A(n48569), .B(n48570), .Z(n48568) );
  XOR U48558 ( .A(n48567), .B(n48571), .Z(n48569) );
  XNOR U48559 ( .A(n48514), .B(n48506), .Z(n48566) );
  XOR U48560 ( .A(n48572), .B(n48573), .Z(n48506) );
  AND U48561 ( .A(n48574), .B(n48575), .Z(n48573) );
  XOR U48562 ( .A(n48572), .B(n48576), .Z(n48574) );
  XNOR U48563 ( .A(n48577), .B(n48511), .Z(n48514) );
  XOR U48564 ( .A(n48578), .B(n48579), .Z(n48511) );
  AND U48565 ( .A(n48580), .B(n48581), .Z(n48579) );
  XNOR U48566 ( .A(n48582), .B(n48583), .Z(n48580) );
  IV U48567 ( .A(n48578), .Z(n48582) );
  XNOR U48568 ( .A(n48584), .B(n48585), .Z(n48577) );
  NOR U48569 ( .A(n48586), .B(n48587), .Z(n48585) );
  XNOR U48570 ( .A(n48584), .B(n48588), .Z(n48586) );
  XOR U48571 ( .A(n48504), .B(n48516), .Z(n48542) );
  NOR U48572 ( .A(n48433), .B(n48589), .Z(n48516) );
  XNOR U48573 ( .A(n48522), .B(n48521), .Z(n48504) );
  XNOR U48574 ( .A(n48590), .B(n48527), .Z(n48521) );
  XNOR U48575 ( .A(n48591), .B(n48592), .Z(n48527) );
  NOR U48576 ( .A(n48593), .B(n48594), .Z(n48592) );
  XOR U48577 ( .A(n48591), .B(n48595), .Z(n48593) );
  XNOR U48578 ( .A(n48526), .B(n48518), .Z(n48590) );
  XOR U48579 ( .A(n48596), .B(n48597), .Z(n48518) );
  AND U48580 ( .A(n48598), .B(n48599), .Z(n48597) );
  XOR U48581 ( .A(n48596), .B(n48600), .Z(n48598) );
  XNOR U48582 ( .A(n48601), .B(n48523), .Z(n48526) );
  XOR U48583 ( .A(n48602), .B(n48603), .Z(n48523) );
  AND U48584 ( .A(n48604), .B(n48605), .Z(n48603) );
  XNOR U48585 ( .A(n48606), .B(n48607), .Z(n48604) );
  IV U48586 ( .A(n48602), .Z(n48606) );
  XNOR U48587 ( .A(n48608), .B(n48609), .Z(n48601) );
  NOR U48588 ( .A(n48610), .B(n48611), .Z(n48609) );
  XNOR U48589 ( .A(n48608), .B(n48612), .Z(n48610) );
  XOR U48590 ( .A(n48532), .B(n48531), .Z(n48522) );
  XNOR U48591 ( .A(n48613), .B(n48528), .Z(n48531) );
  XOR U48592 ( .A(n48614), .B(n48615), .Z(n48528) );
  AND U48593 ( .A(n48616), .B(n48617), .Z(n48615) );
  XNOR U48594 ( .A(n48618), .B(n48619), .Z(n48616) );
  IV U48595 ( .A(n48614), .Z(n48618) );
  XNOR U48596 ( .A(n48620), .B(n48621), .Z(n48613) );
  NOR U48597 ( .A(n48622), .B(n48623), .Z(n48621) );
  XNOR U48598 ( .A(n48620), .B(n48624), .Z(n48622) );
  XOR U48599 ( .A(n48625), .B(n48626), .Z(n48532) );
  NOR U48600 ( .A(n48627), .B(n48628), .Z(n48626) );
  XNOR U48601 ( .A(n48625), .B(n48629), .Z(n48627) );
  XNOR U48602 ( .A(n48424), .B(n48538), .Z(n48540) );
  XNOR U48603 ( .A(n48630), .B(n48631), .Z(n48424) );
  AND U48604 ( .A(n1199), .B(n48632), .Z(n48631) );
  XNOR U48605 ( .A(n48633), .B(n48634), .Z(n48632) );
  AND U48606 ( .A(n48430), .B(n48433), .Z(n48538) );
  XOR U48607 ( .A(n48635), .B(n48589), .Z(n48433) );
  XNOR U48608 ( .A(p_input[1792]), .B(p_input[2048]), .Z(n48589) );
  XNOR U48609 ( .A(n48565), .B(n48564), .Z(n48635) );
  XNOR U48610 ( .A(n48636), .B(n48576), .Z(n48564) );
  XOR U48611 ( .A(n48550), .B(n48548), .Z(n48576) );
  XNOR U48612 ( .A(n48637), .B(n48555), .Z(n48548) );
  XOR U48613 ( .A(p_input[1816]), .B(p_input[2072]), .Z(n48555) );
  XOR U48614 ( .A(n48545), .B(n48554), .Z(n48637) );
  XOR U48615 ( .A(n48638), .B(n48551), .Z(n48554) );
  XOR U48616 ( .A(p_input[1814]), .B(p_input[2070]), .Z(n48551) );
  XOR U48617 ( .A(p_input[1815]), .B(n29410), .Z(n48638) );
  XOR U48618 ( .A(p_input[1810]), .B(p_input[2066]), .Z(n48545) );
  XNOR U48619 ( .A(n48560), .B(n48559), .Z(n48550) );
  XOR U48620 ( .A(n48639), .B(n48556), .Z(n48559) );
  XOR U48621 ( .A(p_input[1811]), .B(p_input[2067]), .Z(n48556) );
  XOR U48622 ( .A(p_input[1812]), .B(n29412), .Z(n48639) );
  XOR U48623 ( .A(p_input[1813]), .B(p_input[2069]), .Z(n48560) );
  XOR U48624 ( .A(n48575), .B(n48640), .Z(n48636) );
  IV U48625 ( .A(n48561), .Z(n48640) );
  XOR U48626 ( .A(p_input[1793]), .B(p_input[2049]), .Z(n48561) );
  XNOR U48627 ( .A(n48641), .B(n48583), .Z(n48575) );
  XNOR U48628 ( .A(n48571), .B(n48570), .Z(n48583) );
  XNOR U48629 ( .A(n48642), .B(n48567), .Z(n48570) );
  XNOR U48630 ( .A(p_input[1818]), .B(p_input[2074]), .Z(n48567) );
  XOR U48631 ( .A(p_input[1819]), .B(n29415), .Z(n48642) );
  XOR U48632 ( .A(p_input[1820]), .B(p_input[2076]), .Z(n48571) );
  XOR U48633 ( .A(n48581), .B(n48643), .Z(n48641) );
  IV U48634 ( .A(n48572), .Z(n48643) );
  XOR U48635 ( .A(p_input[1809]), .B(p_input[2065]), .Z(n48572) );
  XNOR U48636 ( .A(n48644), .B(n48588), .Z(n48581) );
  XNOR U48637 ( .A(p_input[1823]), .B(n29418), .Z(n48588) );
  XOR U48638 ( .A(n48578), .B(n48587), .Z(n48644) );
  XOR U48639 ( .A(n48645), .B(n48584), .Z(n48587) );
  XOR U48640 ( .A(p_input[1821]), .B(p_input[2077]), .Z(n48584) );
  XOR U48641 ( .A(p_input[1822]), .B(n29420), .Z(n48645) );
  XOR U48642 ( .A(p_input[1817]), .B(p_input[2073]), .Z(n48578) );
  XOR U48643 ( .A(n48600), .B(n48599), .Z(n48565) );
  XNOR U48644 ( .A(n48646), .B(n48607), .Z(n48599) );
  XNOR U48645 ( .A(n48595), .B(n48594), .Z(n48607) );
  XNOR U48646 ( .A(n48647), .B(n48591), .Z(n48594) );
  XNOR U48647 ( .A(p_input[1803]), .B(p_input[2059]), .Z(n48591) );
  XOR U48648 ( .A(p_input[1804]), .B(n28329), .Z(n48647) );
  XOR U48649 ( .A(p_input[1805]), .B(p_input[2061]), .Z(n48595) );
  XOR U48650 ( .A(n48605), .B(n48648), .Z(n48646) );
  IV U48651 ( .A(n48596), .Z(n48648) );
  XOR U48652 ( .A(p_input[1794]), .B(p_input[2050]), .Z(n48596) );
  XNOR U48653 ( .A(n48649), .B(n48612), .Z(n48605) );
  XNOR U48654 ( .A(p_input[1808]), .B(n28332), .Z(n48612) );
  XOR U48655 ( .A(n48602), .B(n48611), .Z(n48649) );
  XOR U48656 ( .A(n48650), .B(n48608), .Z(n48611) );
  XOR U48657 ( .A(p_input[1806]), .B(p_input[2062]), .Z(n48608) );
  XOR U48658 ( .A(p_input[1807]), .B(n28334), .Z(n48650) );
  XOR U48659 ( .A(p_input[1802]), .B(p_input[2058]), .Z(n48602) );
  XOR U48660 ( .A(n48619), .B(n48617), .Z(n48600) );
  XNOR U48661 ( .A(n48651), .B(n48624), .Z(n48617) );
  XOR U48662 ( .A(p_input[1801]), .B(p_input[2057]), .Z(n48624) );
  XOR U48663 ( .A(n48614), .B(n48623), .Z(n48651) );
  XOR U48664 ( .A(n48652), .B(n48620), .Z(n48623) );
  XOR U48665 ( .A(p_input[1799]), .B(p_input[2055]), .Z(n48620) );
  XOR U48666 ( .A(p_input[1800]), .B(n29427), .Z(n48652) );
  XOR U48667 ( .A(p_input[1795]), .B(p_input[2051]), .Z(n48614) );
  XNOR U48668 ( .A(n48629), .B(n48628), .Z(n48619) );
  XOR U48669 ( .A(n48653), .B(n48625), .Z(n48628) );
  XOR U48670 ( .A(p_input[1796]), .B(p_input[2052]), .Z(n48625) );
  XOR U48671 ( .A(p_input[1797]), .B(n29429), .Z(n48653) );
  XOR U48672 ( .A(p_input[1798]), .B(p_input[2054]), .Z(n48629) );
  XNOR U48673 ( .A(n48654), .B(n48655), .Z(n48430) );
  AND U48674 ( .A(n1199), .B(n48656), .Z(n48655) );
  XNOR U48675 ( .A(n48657), .B(n48658), .Z(n1199) );
  AND U48676 ( .A(n48659), .B(n48660), .Z(n48658) );
  XOR U48677 ( .A(n48444), .B(n48657), .Z(n48660) );
  XNOR U48678 ( .A(n48661), .B(n48657), .Z(n48659) );
  XOR U48679 ( .A(n48662), .B(n48663), .Z(n48657) );
  AND U48680 ( .A(n48664), .B(n48665), .Z(n48663) );
  XOR U48681 ( .A(n48459), .B(n48662), .Z(n48665) );
  XOR U48682 ( .A(n48662), .B(n48460), .Z(n48664) );
  XOR U48683 ( .A(n48666), .B(n48667), .Z(n48662) );
  AND U48684 ( .A(n48668), .B(n48669), .Z(n48667) );
  XOR U48685 ( .A(n48487), .B(n48666), .Z(n48669) );
  XOR U48686 ( .A(n48666), .B(n48488), .Z(n48668) );
  XOR U48687 ( .A(n48670), .B(n48671), .Z(n48666) );
  AND U48688 ( .A(n48672), .B(n48673), .Z(n48671) );
  XOR U48689 ( .A(n48536), .B(n48670), .Z(n48673) );
  XOR U48690 ( .A(n48670), .B(n48537), .Z(n48672) );
  XOR U48691 ( .A(n48674), .B(n48675), .Z(n48670) );
  AND U48692 ( .A(n48676), .B(n48677), .Z(n48675) );
  XOR U48693 ( .A(n48674), .B(n48633), .Z(n48677) );
  XNOR U48694 ( .A(n48678), .B(n48679), .Z(n48380) );
  AND U48695 ( .A(n1203), .B(n48680), .Z(n48679) );
  XNOR U48696 ( .A(n48681), .B(n48682), .Z(n1203) );
  AND U48697 ( .A(n48683), .B(n48684), .Z(n48682) );
  XOR U48698 ( .A(n48681), .B(n48390), .Z(n48684) );
  XNOR U48699 ( .A(n48681), .B(n48340), .Z(n48683) );
  XOR U48700 ( .A(n48685), .B(n48686), .Z(n48681) );
  AND U48701 ( .A(n48687), .B(n48688), .Z(n48686) );
  XNOR U48702 ( .A(n48400), .B(n48685), .Z(n48688) );
  XOR U48703 ( .A(n48685), .B(n48350), .Z(n48687) );
  XOR U48704 ( .A(n48689), .B(n48690), .Z(n48685) );
  AND U48705 ( .A(n48691), .B(n48692), .Z(n48690) );
  XNOR U48706 ( .A(n48410), .B(n48689), .Z(n48692) );
  XOR U48707 ( .A(n48689), .B(n48359), .Z(n48691) );
  XOR U48708 ( .A(n48693), .B(n48694), .Z(n48689) );
  AND U48709 ( .A(n48695), .B(n48696), .Z(n48694) );
  XOR U48710 ( .A(n48693), .B(n48367), .Z(n48695) );
  XOR U48711 ( .A(n48697), .B(n48698), .Z(n48331) );
  AND U48712 ( .A(n1207), .B(n48680), .Z(n48698) );
  XNOR U48713 ( .A(n48678), .B(n48697), .Z(n48680) );
  XNOR U48714 ( .A(n48699), .B(n48700), .Z(n1207) );
  AND U48715 ( .A(n48701), .B(n48702), .Z(n48700) );
  XNOR U48716 ( .A(n48703), .B(n48699), .Z(n48702) );
  IV U48717 ( .A(n48390), .Z(n48703) );
  XOR U48718 ( .A(n48661), .B(n48704), .Z(n48390) );
  AND U48719 ( .A(n1210), .B(n48705), .Z(n48704) );
  XOR U48720 ( .A(n48443), .B(n48440), .Z(n48705) );
  XNOR U48721 ( .A(n48340), .B(n48699), .Z(n48701) );
  XNOR U48722 ( .A(n48706), .B(n48707), .Z(n48340) );
  AND U48723 ( .A(n1226), .B(n48708), .Z(n48707) );
  XNOR U48724 ( .A(n48709), .B(n48710), .Z(n48708) );
  XOR U48725 ( .A(n48711), .B(n48712), .Z(n48699) );
  AND U48726 ( .A(n48713), .B(n48714), .Z(n48712) );
  XNOR U48727 ( .A(n48711), .B(n48400), .Z(n48714) );
  XOR U48728 ( .A(n48460), .B(n48715), .Z(n48400) );
  AND U48729 ( .A(n1210), .B(n48716), .Z(n48715) );
  XOR U48730 ( .A(n48456), .B(n48460), .Z(n48716) );
  XNOR U48731 ( .A(n48717), .B(n48711), .Z(n48713) );
  IV U48732 ( .A(n48350), .Z(n48717) );
  XOR U48733 ( .A(n48718), .B(n48719), .Z(n48350) );
  AND U48734 ( .A(n1226), .B(n48720), .Z(n48719) );
  XOR U48735 ( .A(n48721), .B(n48722), .Z(n48711) );
  AND U48736 ( .A(n48723), .B(n48724), .Z(n48722) );
  XNOR U48737 ( .A(n48721), .B(n48410), .Z(n48724) );
  XOR U48738 ( .A(n48488), .B(n48725), .Z(n48410) );
  AND U48739 ( .A(n1210), .B(n48726), .Z(n48725) );
  XOR U48740 ( .A(n48484), .B(n48488), .Z(n48726) );
  XOR U48741 ( .A(n48359), .B(n48721), .Z(n48723) );
  XOR U48742 ( .A(n48727), .B(n48728), .Z(n48359) );
  AND U48743 ( .A(n1226), .B(n48729), .Z(n48728) );
  XOR U48744 ( .A(n48693), .B(n48730), .Z(n48721) );
  AND U48745 ( .A(n48731), .B(n48696), .Z(n48730) );
  XNOR U48746 ( .A(n48420), .B(n48693), .Z(n48696) );
  XOR U48747 ( .A(n48537), .B(n48732), .Z(n48420) );
  AND U48748 ( .A(n1210), .B(n48733), .Z(n48732) );
  XOR U48749 ( .A(n48533), .B(n48537), .Z(n48733) );
  XNOR U48750 ( .A(n48734), .B(n48693), .Z(n48731) );
  IV U48751 ( .A(n48367), .Z(n48734) );
  XOR U48752 ( .A(n48735), .B(n48736), .Z(n48367) );
  AND U48753 ( .A(n1226), .B(n48737), .Z(n48736) );
  XOR U48754 ( .A(n48738), .B(n48739), .Z(n48693) );
  AND U48755 ( .A(n48740), .B(n48741), .Z(n48739) );
  XNOR U48756 ( .A(n48738), .B(n48428), .Z(n48741) );
  XOR U48757 ( .A(n48634), .B(n48742), .Z(n48428) );
  AND U48758 ( .A(n1210), .B(n48743), .Z(n48742) );
  XOR U48759 ( .A(n48630), .B(n48634), .Z(n48743) );
  XNOR U48760 ( .A(n48744), .B(n48738), .Z(n48740) );
  IV U48761 ( .A(n48377), .Z(n48744) );
  XOR U48762 ( .A(n48745), .B(n48746), .Z(n48377) );
  AND U48763 ( .A(n1226), .B(n48747), .Z(n48746) );
  AND U48764 ( .A(n48697), .B(n48678), .Z(n48738) );
  XNOR U48765 ( .A(n48748), .B(n48749), .Z(n48678) );
  AND U48766 ( .A(n1210), .B(n48656), .Z(n48749) );
  XNOR U48767 ( .A(n48654), .B(n48748), .Z(n48656) );
  XNOR U48768 ( .A(n48750), .B(n48751), .Z(n1210) );
  AND U48769 ( .A(n48752), .B(n48753), .Z(n48751) );
  XNOR U48770 ( .A(n48750), .B(n48440), .Z(n48753) );
  IV U48771 ( .A(n48444), .Z(n48440) );
  XOR U48772 ( .A(n48754), .B(n48755), .Z(n48444) );
  AND U48773 ( .A(n1214), .B(n48756), .Z(n48755) );
  XOR U48774 ( .A(n48757), .B(n48754), .Z(n48756) );
  XNOR U48775 ( .A(n48750), .B(n48661), .Z(n48752) );
  IV U48776 ( .A(n48443), .Z(n48661) );
  XOR U48777 ( .A(n48709), .B(n48758), .Z(n48443) );
  AND U48778 ( .A(n1222), .B(n48759), .Z(n48758) );
  XOR U48779 ( .A(n48709), .B(n48706), .Z(n48759) );
  XOR U48780 ( .A(n48760), .B(n48761), .Z(n48750) );
  AND U48781 ( .A(n48762), .B(n48763), .Z(n48761) );
  XNOR U48782 ( .A(n48760), .B(n48456), .Z(n48763) );
  IV U48783 ( .A(n48459), .Z(n48456) );
  XOR U48784 ( .A(n48764), .B(n48765), .Z(n48459) );
  AND U48785 ( .A(n1214), .B(n48766), .Z(n48765) );
  XOR U48786 ( .A(n48767), .B(n48764), .Z(n48766) );
  XOR U48787 ( .A(n48460), .B(n48760), .Z(n48762) );
  XOR U48788 ( .A(n48768), .B(n48769), .Z(n48460) );
  AND U48789 ( .A(n1222), .B(n48720), .Z(n48769) );
  XOR U48790 ( .A(n48768), .B(n48718), .Z(n48720) );
  XOR U48791 ( .A(n48770), .B(n48771), .Z(n48760) );
  AND U48792 ( .A(n48772), .B(n48773), .Z(n48771) );
  XNOR U48793 ( .A(n48770), .B(n48484), .Z(n48773) );
  IV U48794 ( .A(n48487), .Z(n48484) );
  XOR U48795 ( .A(n48774), .B(n48775), .Z(n48487) );
  AND U48796 ( .A(n1214), .B(n48776), .Z(n48775) );
  XNOR U48797 ( .A(n48777), .B(n48774), .Z(n48776) );
  XOR U48798 ( .A(n48488), .B(n48770), .Z(n48772) );
  XOR U48799 ( .A(n48778), .B(n48779), .Z(n48488) );
  AND U48800 ( .A(n1222), .B(n48729), .Z(n48779) );
  XOR U48801 ( .A(n48778), .B(n48727), .Z(n48729) );
  XOR U48802 ( .A(n48780), .B(n48781), .Z(n48770) );
  AND U48803 ( .A(n48782), .B(n48783), .Z(n48781) );
  XNOR U48804 ( .A(n48780), .B(n48533), .Z(n48783) );
  IV U48805 ( .A(n48536), .Z(n48533) );
  XOR U48806 ( .A(n48784), .B(n48785), .Z(n48536) );
  AND U48807 ( .A(n1214), .B(n48786), .Z(n48785) );
  XOR U48808 ( .A(n48787), .B(n48784), .Z(n48786) );
  XOR U48809 ( .A(n48537), .B(n48780), .Z(n48782) );
  XOR U48810 ( .A(n48788), .B(n48789), .Z(n48537) );
  AND U48811 ( .A(n1222), .B(n48737), .Z(n48789) );
  XOR U48812 ( .A(n48788), .B(n48735), .Z(n48737) );
  XOR U48813 ( .A(n48674), .B(n48790), .Z(n48780) );
  AND U48814 ( .A(n48676), .B(n48791), .Z(n48790) );
  XNOR U48815 ( .A(n48674), .B(n48630), .Z(n48791) );
  IV U48816 ( .A(n48633), .Z(n48630) );
  XOR U48817 ( .A(n48792), .B(n48793), .Z(n48633) );
  AND U48818 ( .A(n1214), .B(n48794), .Z(n48793) );
  XNOR U48819 ( .A(n48795), .B(n48792), .Z(n48794) );
  XOR U48820 ( .A(n48634), .B(n48674), .Z(n48676) );
  XOR U48821 ( .A(n48796), .B(n48797), .Z(n48634) );
  AND U48822 ( .A(n1222), .B(n48747), .Z(n48797) );
  XOR U48823 ( .A(n48796), .B(n48745), .Z(n48747) );
  AND U48824 ( .A(n48748), .B(n48654), .Z(n48674) );
  XNOR U48825 ( .A(n48798), .B(n48799), .Z(n48654) );
  AND U48826 ( .A(n1214), .B(n48800), .Z(n48799) );
  XNOR U48827 ( .A(n48801), .B(n48798), .Z(n48800) );
  XNOR U48828 ( .A(n48802), .B(n48803), .Z(n1214) );
  AND U48829 ( .A(n48804), .B(n48805), .Z(n48803) );
  XOR U48830 ( .A(n48757), .B(n48802), .Z(n48805) );
  AND U48831 ( .A(n48806), .B(n48807), .Z(n48757) );
  XNOR U48832 ( .A(n48754), .B(n48802), .Z(n48804) );
  XNOR U48833 ( .A(n48808), .B(n48809), .Z(n48754) );
  AND U48834 ( .A(n48810), .B(n1218), .Z(n48809) );
  XOR U48835 ( .A(n48811), .B(n48812), .Z(n48802) );
  AND U48836 ( .A(n48813), .B(n48814), .Z(n48812) );
  XNOR U48837 ( .A(n48811), .B(n48806), .Z(n48814) );
  IV U48838 ( .A(n48767), .Z(n48806) );
  XOR U48839 ( .A(n48815), .B(n48816), .Z(n48767) );
  XOR U48840 ( .A(n48817), .B(n48807), .Z(n48816) );
  AND U48841 ( .A(n48777), .B(n48818), .Z(n48807) );
  AND U48842 ( .A(n48819), .B(n48820), .Z(n48817) );
  XOR U48843 ( .A(n48821), .B(n48815), .Z(n48819) );
  XNOR U48844 ( .A(n48764), .B(n48811), .Z(n48813) );
  XNOR U48845 ( .A(n48822), .B(n48823), .Z(n48764) );
  AND U48846 ( .A(n1218), .B(n48824), .Z(n48823) );
  XNOR U48847 ( .A(n48825), .B(n48826), .Z(n48824) );
  XOR U48848 ( .A(n48827), .B(n48828), .Z(n48811) );
  AND U48849 ( .A(n48829), .B(n48830), .Z(n48828) );
  XNOR U48850 ( .A(n48827), .B(n48777), .Z(n48830) );
  XOR U48851 ( .A(n48831), .B(n48820), .Z(n48777) );
  XNOR U48852 ( .A(n48832), .B(n48815), .Z(n48820) );
  XOR U48853 ( .A(n48833), .B(n48834), .Z(n48815) );
  AND U48854 ( .A(n48835), .B(n48836), .Z(n48834) );
  XOR U48855 ( .A(n48837), .B(n48833), .Z(n48835) );
  XNOR U48856 ( .A(n48838), .B(n48839), .Z(n48832) );
  AND U48857 ( .A(n48840), .B(n48841), .Z(n48839) );
  XOR U48858 ( .A(n48838), .B(n48842), .Z(n48840) );
  XNOR U48859 ( .A(n48821), .B(n48818), .Z(n48831) );
  AND U48860 ( .A(n48843), .B(n48844), .Z(n48818) );
  XOR U48861 ( .A(n48845), .B(n48846), .Z(n48821) );
  AND U48862 ( .A(n48847), .B(n48848), .Z(n48846) );
  XOR U48863 ( .A(n48845), .B(n48849), .Z(n48847) );
  XNOR U48864 ( .A(n48774), .B(n48827), .Z(n48829) );
  XNOR U48865 ( .A(n48850), .B(n48851), .Z(n48774) );
  AND U48866 ( .A(n1218), .B(n48852), .Z(n48851) );
  XNOR U48867 ( .A(n48853), .B(n48854), .Z(n48852) );
  XOR U48868 ( .A(n48855), .B(n48856), .Z(n48827) );
  AND U48869 ( .A(n48857), .B(n48858), .Z(n48856) );
  XNOR U48870 ( .A(n48855), .B(n48843), .Z(n48858) );
  IV U48871 ( .A(n48787), .Z(n48843) );
  XNOR U48872 ( .A(n48859), .B(n48836), .Z(n48787) );
  XNOR U48873 ( .A(n48860), .B(n48842), .Z(n48836) );
  XOR U48874 ( .A(n48861), .B(n48862), .Z(n48842) );
  AND U48875 ( .A(n48863), .B(n48864), .Z(n48862) );
  XOR U48876 ( .A(n48861), .B(n48865), .Z(n48863) );
  XNOR U48877 ( .A(n48841), .B(n48833), .Z(n48860) );
  XOR U48878 ( .A(n48866), .B(n48867), .Z(n48833) );
  AND U48879 ( .A(n48868), .B(n48869), .Z(n48867) );
  XNOR U48880 ( .A(n48870), .B(n48866), .Z(n48868) );
  XNOR U48881 ( .A(n48871), .B(n48838), .Z(n48841) );
  XOR U48882 ( .A(n48872), .B(n48873), .Z(n48838) );
  AND U48883 ( .A(n48874), .B(n48875), .Z(n48873) );
  XOR U48884 ( .A(n48872), .B(n48876), .Z(n48874) );
  XNOR U48885 ( .A(n48877), .B(n48878), .Z(n48871) );
  AND U48886 ( .A(n48879), .B(n48880), .Z(n48878) );
  XNOR U48887 ( .A(n48877), .B(n48881), .Z(n48879) );
  XNOR U48888 ( .A(n48837), .B(n48844), .Z(n48859) );
  AND U48889 ( .A(n48795), .B(n48882), .Z(n48844) );
  XOR U48890 ( .A(n48849), .B(n48848), .Z(n48837) );
  XNOR U48891 ( .A(n48883), .B(n48845), .Z(n48848) );
  XOR U48892 ( .A(n48884), .B(n48885), .Z(n48845) );
  AND U48893 ( .A(n48886), .B(n48887), .Z(n48885) );
  XOR U48894 ( .A(n48884), .B(n48888), .Z(n48886) );
  XNOR U48895 ( .A(n48889), .B(n48890), .Z(n48883) );
  AND U48896 ( .A(n48891), .B(n48892), .Z(n48890) );
  XOR U48897 ( .A(n48889), .B(n48893), .Z(n48891) );
  XOR U48898 ( .A(n48894), .B(n48895), .Z(n48849) );
  AND U48899 ( .A(n48896), .B(n48897), .Z(n48895) );
  XOR U48900 ( .A(n48894), .B(n48898), .Z(n48896) );
  XNOR U48901 ( .A(n48784), .B(n48855), .Z(n48857) );
  XNOR U48902 ( .A(n48899), .B(n48900), .Z(n48784) );
  AND U48903 ( .A(n1218), .B(n48901), .Z(n48900) );
  XNOR U48904 ( .A(n48902), .B(n48903), .Z(n48901) );
  XOR U48905 ( .A(n48904), .B(n48905), .Z(n48855) );
  AND U48906 ( .A(n48906), .B(n48907), .Z(n48905) );
  XNOR U48907 ( .A(n48904), .B(n48795), .Z(n48907) );
  XOR U48908 ( .A(n48908), .B(n48869), .Z(n48795) );
  XNOR U48909 ( .A(n48909), .B(n48876), .Z(n48869) );
  XOR U48910 ( .A(n48865), .B(n48864), .Z(n48876) );
  XNOR U48911 ( .A(n48910), .B(n48861), .Z(n48864) );
  XOR U48912 ( .A(n48911), .B(n48912), .Z(n48861) );
  AND U48913 ( .A(n48913), .B(n48914), .Z(n48912) );
  XNOR U48914 ( .A(n48915), .B(n48916), .Z(n48913) );
  IV U48915 ( .A(n48911), .Z(n48915) );
  XNOR U48916 ( .A(n48917), .B(n48918), .Z(n48910) );
  NOR U48917 ( .A(n48919), .B(n48920), .Z(n48918) );
  XNOR U48918 ( .A(n48917), .B(n48921), .Z(n48919) );
  XOR U48919 ( .A(n48922), .B(n48923), .Z(n48865) );
  NOR U48920 ( .A(n48924), .B(n48925), .Z(n48923) );
  XNOR U48921 ( .A(n48922), .B(n48926), .Z(n48924) );
  XNOR U48922 ( .A(n48875), .B(n48866), .Z(n48909) );
  XOR U48923 ( .A(n48927), .B(n48928), .Z(n48866) );
  AND U48924 ( .A(n48929), .B(n48930), .Z(n48928) );
  XOR U48925 ( .A(n48927), .B(n48931), .Z(n48929) );
  XOR U48926 ( .A(n48932), .B(n48881), .Z(n48875) );
  XOR U48927 ( .A(n48933), .B(n48934), .Z(n48881) );
  NOR U48928 ( .A(n48935), .B(n48936), .Z(n48934) );
  XOR U48929 ( .A(n48933), .B(n48937), .Z(n48935) );
  XNOR U48930 ( .A(n48880), .B(n48872), .Z(n48932) );
  XOR U48931 ( .A(n48938), .B(n48939), .Z(n48872) );
  AND U48932 ( .A(n48940), .B(n48941), .Z(n48939) );
  XOR U48933 ( .A(n48938), .B(n48942), .Z(n48940) );
  XNOR U48934 ( .A(n48943), .B(n48877), .Z(n48880) );
  XOR U48935 ( .A(n48944), .B(n48945), .Z(n48877) );
  AND U48936 ( .A(n48946), .B(n48947), .Z(n48945) );
  XNOR U48937 ( .A(n48948), .B(n48949), .Z(n48946) );
  IV U48938 ( .A(n48944), .Z(n48948) );
  XNOR U48939 ( .A(n48950), .B(n48951), .Z(n48943) );
  NOR U48940 ( .A(n48952), .B(n48953), .Z(n48951) );
  XNOR U48941 ( .A(n48950), .B(n48954), .Z(n48952) );
  XOR U48942 ( .A(n48870), .B(n48882), .Z(n48908) );
  NOR U48943 ( .A(n48801), .B(n48955), .Z(n48882) );
  XNOR U48944 ( .A(n48888), .B(n48887), .Z(n48870) );
  XNOR U48945 ( .A(n48956), .B(n48893), .Z(n48887) );
  XNOR U48946 ( .A(n48957), .B(n48958), .Z(n48893) );
  NOR U48947 ( .A(n48959), .B(n48960), .Z(n48958) );
  XOR U48948 ( .A(n48957), .B(n48961), .Z(n48959) );
  XNOR U48949 ( .A(n48892), .B(n48884), .Z(n48956) );
  XOR U48950 ( .A(n48962), .B(n48963), .Z(n48884) );
  AND U48951 ( .A(n48964), .B(n48965), .Z(n48963) );
  XOR U48952 ( .A(n48962), .B(n48966), .Z(n48964) );
  XNOR U48953 ( .A(n48967), .B(n48889), .Z(n48892) );
  XOR U48954 ( .A(n48968), .B(n48969), .Z(n48889) );
  AND U48955 ( .A(n48970), .B(n48971), .Z(n48969) );
  XNOR U48956 ( .A(n48972), .B(n48973), .Z(n48970) );
  IV U48957 ( .A(n48968), .Z(n48972) );
  XNOR U48958 ( .A(n48974), .B(n48975), .Z(n48967) );
  NOR U48959 ( .A(n48976), .B(n48977), .Z(n48975) );
  XNOR U48960 ( .A(n48974), .B(n48978), .Z(n48976) );
  XOR U48961 ( .A(n48898), .B(n48897), .Z(n48888) );
  XNOR U48962 ( .A(n48979), .B(n48894), .Z(n48897) );
  XOR U48963 ( .A(n48980), .B(n48981), .Z(n48894) );
  AND U48964 ( .A(n48982), .B(n48983), .Z(n48981) );
  XNOR U48965 ( .A(n48984), .B(n48985), .Z(n48982) );
  IV U48966 ( .A(n48980), .Z(n48984) );
  XNOR U48967 ( .A(n48986), .B(n48987), .Z(n48979) );
  NOR U48968 ( .A(n48988), .B(n48989), .Z(n48987) );
  XNOR U48969 ( .A(n48986), .B(n48990), .Z(n48988) );
  XOR U48970 ( .A(n48991), .B(n48992), .Z(n48898) );
  NOR U48971 ( .A(n48993), .B(n48994), .Z(n48992) );
  XNOR U48972 ( .A(n48991), .B(n48995), .Z(n48993) );
  XNOR U48973 ( .A(n48792), .B(n48904), .Z(n48906) );
  XNOR U48974 ( .A(n48996), .B(n48997), .Z(n48792) );
  AND U48975 ( .A(n1218), .B(n48998), .Z(n48997) );
  XNOR U48976 ( .A(n48999), .B(n49000), .Z(n48998) );
  AND U48977 ( .A(n48798), .B(n48801), .Z(n48904) );
  XOR U48978 ( .A(n49001), .B(n48955), .Z(n48801) );
  XNOR U48979 ( .A(p_input[1824]), .B(p_input[2048]), .Z(n48955) );
  XNOR U48980 ( .A(n48931), .B(n48930), .Z(n49001) );
  XNOR U48981 ( .A(n49002), .B(n48942), .Z(n48930) );
  XOR U48982 ( .A(n48916), .B(n48914), .Z(n48942) );
  XNOR U48983 ( .A(n49003), .B(n48921), .Z(n48914) );
  XOR U48984 ( .A(p_input[1848]), .B(p_input[2072]), .Z(n48921) );
  XOR U48985 ( .A(n48911), .B(n48920), .Z(n49003) );
  XOR U48986 ( .A(n49004), .B(n48917), .Z(n48920) );
  XOR U48987 ( .A(p_input[1846]), .B(p_input[2070]), .Z(n48917) );
  XOR U48988 ( .A(p_input[1847]), .B(n29410), .Z(n49004) );
  XOR U48989 ( .A(p_input[1842]), .B(p_input[2066]), .Z(n48911) );
  XNOR U48990 ( .A(n48926), .B(n48925), .Z(n48916) );
  XOR U48991 ( .A(n49005), .B(n48922), .Z(n48925) );
  XOR U48992 ( .A(p_input[1843]), .B(p_input[2067]), .Z(n48922) );
  XOR U48993 ( .A(p_input[1844]), .B(n29412), .Z(n49005) );
  XOR U48994 ( .A(p_input[1845]), .B(p_input[2069]), .Z(n48926) );
  XOR U48995 ( .A(n48941), .B(n49006), .Z(n49002) );
  IV U48996 ( .A(n48927), .Z(n49006) );
  XOR U48997 ( .A(p_input[1825]), .B(p_input[2049]), .Z(n48927) );
  XNOR U48998 ( .A(n49007), .B(n48949), .Z(n48941) );
  XNOR U48999 ( .A(n48937), .B(n48936), .Z(n48949) );
  XNOR U49000 ( .A(n49008), .B(n48933), .Z(n48936) );
  XNOR U49001 ( .A(p_input[1850]), .B(p_input[2074]), .Z(n48933) );
  XOR U49002 ( .A(p_input[1851]), .B(n29415), .Z(n49008) );
  XOR U49003 ( .A(p_input[1852]), .B(p_input[2076]), .Z(n48937) );
  XOR U49004 ( .A(n48947), .B(n49009), .Z(n49007) );
  IV U49005 ( .A(n48938), .Z(n49009) );
  XOR U49006 ( .A(p_input[1841]), .B(p_input[2065]), .Z(n48938) );
  XNOR U49007 ( .A(n49010), .B(n48954), .Z(n48947) );
  XNOR U49008 ( .A(p_input[1855]), .B(n29418), .Z(n48954) );
  XOR U49009 ( .A(n48944), .B(n48953), .Z(n49010) );
  XOR U49010 ( .A(n49011), .B(n48950), .Z(n48953) );
  XOR U49011 ( .A(p_input[1853]), .B(p_input[2077]), .Z(n48950) );
  XOR U49012 ( .A(p_input[1854]), .B(n29420), .Z(n49011) );
  XOR U49013 ( .A(p_input[1849]), .B(p_input[2073]), .Z(n48944) );
  XOR U49014 ( .A(n48966), .B(n48965), .Z(n48931) );
  XNOR U49015 ( .A(n49012), .B(n48973), .Z(n48965) );
  XNOR U49016 ( .A(n48961), .B(n48960), .Z(n48973) );
  XNOR U49017 ( .A(n49013), .B(n48957), .Z(n48960) );
  XNOR U49018 ( .A(p_input[1835]), .B(p_input[2059]), .Z(n48957) );
  XOR U49019 ( .A(p_input[1836]), .B(n28329), .Z(n49013) );
  XOR U49020 ( .A(p_input[1837]), .B(p_input[2061]), .Z(n48961) );
  XOR U49021 ( .A(n48971), .B(n49014), .Z(n49012) );
  IV U49022 ( .A(n48962), .Z(n49014) );
  XOR U49023 ( .A(p_input[1826]), .B(p_input[2050]), .Z(n48962) );
  XNOR U49024 ( .A(n49015), .B(n48978), .Z(n48971) );
  XNOR U49025 ( .A(p_input[1840]), .B(n28332), .Z(n48978) );
  XOR U49026 ( .A(n48968), .B(n48977), .Z(n49015) );
  XOR U49027 ( .A(n49016), .B(n48974), .Z(n48977) );
  XOR U49028 ( .A(p_input[1838]), .B(p_input[2062]), .Z(n48974) );
  XOR U49029 ( .A(p_input[1839]), .B(n28334), .Z(n49016) );
  XOR U49030 ( .A(p_input[1834]), .B(p_input[2058]), .Z(n48968) );
  XOR U49031 ( .A(n48985), .B(n48983), .Z(n48966) );
  XNOR U49032 ( .A(n49017), .B(n48990), .Z(n48983) );
  XOR U49033 ( .A(p_input[1833]), .B(p_input[2057]), .Z(n48990) );
  XOR U49034 ( .A(n48980), .B(n48989), .Z(n49017) );
  XOR U49035 ( .A(n49018), .B(n48986), .Z(n48989) );
  XOR U49036 ( .A(p_input[1831]), .B(p_input[2055]), .Z(n48986) );
  XOR U49037 ( .A(p_input[1832]), .B(n29427), .Z(n49018) );
  XOR U49038 ( .A(p_input[1827]), .B(p_input[2051]), .Z(n48980) );
  XNOR U49039 ( .A(n48995), .B(n48994), .Z(n48985) );
  XOR U49040 ( .A(n49019), .B(n48991), .Z(n48994) );
  XOR U49041 ( .A(p_input[1828]), .B(p_input[2052]), .Z(n48991) );
  XOR U49042 ( .A(p_input[1829]), .B(n29429), .Z(n49019) );
  XOR U49043 ( .A(p_input[1830]), .B(p_input[2054]), .Z(n48995) );
  XNOR U49044 ( .A(n49020), .B(n49021), .Z(n48798) );
  AND U49045 ( .A(n1218), .B(n49022), .Z(n49021) );
  XNOR U49046 ( .A(n49023), .B(n49024), .Z(n1218) );
  NOR U49047 ( .A(n49025), .B(n49026), .Z(n49024) );
  XNOR U49048 ( .A(n49027), .B(n49028), .Z(n49026) );
  AND U49049 ( .A(n49027), .B(n48808), .Z(n49025) );
  IV U49050 ( .A(n49023), .Z(n49027) );
  XOR U49051 ( .A(n49029), .B(n49030), .Z(n49023) );
  AND U49052 ( .A(n49031), .B(n49032), .Z(n49030) );
  XOR U49053 ( .A(n48825), .B(n49029), .Z(n49032) );
  XOR U49054 ( .A(n49029), .B(n48826), .Z(n49031) );
  XOR U49055 ( .A(n49033), .B(n49034), .Z(n49029) );
  AND U49056 ( .A(n49035), .B(n49036), .Z(n49034) );
  XOR U49057 ( .A(n48853), .B(n49033), .Z(n49036) );
  XOR U49058 ( .A(n49033), .B(n48854), .Z(n49035) );
  XOR U49059 ( .A(n49037), .B(n49038), .Z(n49033) );
  AND U49060 ( .A(n49039), .B(n49040), .Z(n49038) );
  XOR U49061 ( .A(n48902), .B(n49037), .Z(n49040) );
  XOR U49062 ( .A(n49037), .B(n48903), .Z(n49039) );
  XOR U49063 ( .A(n49041), .B(n49042), .Z(n49037) );
  AND U49064 ( .A(n49043), .B(n49044), .Z(n49042) );
  XOR U49065 ( .A(n49041), .B(n48999), .Z(n49044) );
  XNOR U49066 ( .A(n49045), .B(n49046), .Z(n48748) );
  AND U49067 ( .A(n1222), .B(n49047), .Z(n49046) );
  XNOR U49068 ( .A(n49048), .B(n49049), .Z(n1222) );
  AND U49069 ( .A(n49050), .B(n49051), .Z(n49049) );
  XNOR U49070 ( .A(n49048), .B(n48709), .Z(n49051) );
  XOR U49071 ( .A(n49048), .B(n48706), .Z(n49050) );
  XOR U49072 ( .A(n49052), .B(n49053), .Z(n49048) );
  AND U49073 ( .A(n49054), .B(n49055), .Z(n49053) );
  XNOR U49074 ( .A(n48768), .B(n49052), .Z(n49055) );
  XOR U49075 ( .A(n49052), .B(n48718), .Z(n49054) );
  XOR U49076 ( .A(n49056), .B(n49057), .Z(n49052) );
  AND U49077 ( .A(n49058), .B(n49059), .Z(n49057) );
  XNOR U49078 ( .A(n48778), .B(n49056), .Z(n49059) );
  XOR U49079 ( .A(n49056), .B(n48727), .Z(n49058) );
  XOR U49080 ( .A(n49060), .B(n49061), .Z(n49056) );
  AND U49081 ( .A(n49062), .B(n49063), .Z(n49061) );
  XOR U49082 ( .A(n49060), .B(n48735), .Z(n49062) );
  XOR U49083 ( .A(n49064), .B(n49065), .Z(n48697) );
  AND U49084 ( .A(n1226), .B(n49047), .Z(n49065) );
  XNOR U49085 ( .A(n49045), .B(n49064), .Z(n49047) );
  XNOR U49086 ( .A(n49066), .B(n49067), .Z(n1226) );
  AND U49087 ( .A(n49068), .B(n49069), .Z(n49067) );
  XNOR U49088 ( .A(n48709), .B(n49066), .Z(n49069) );
  XNOR U49089 ( .A(n49028), .B(n49070), .Z(n48709) );
  AND U49090 ( .A(n48810), .B(n1229), .Z(n49070) );
  NOR U49091 ( .A(n49071), .B(n49072), .Z(n48810) );
  XOR U49092 ( .A(n49066), .B(n48706), .Z(n49068) );
  IV U49093 ( .A(n48710), .Z(n48706) );
  AND U49094 ( .A(n49073), .B(n49074), .Z(n48710) );
  XOR U49095 ( .A(n49075), .B(n49076), .Z(n49066) );
  AND U49096 ( .A(n49077), .B(n49078), .Z(n49076) );
  XNOR U49097 ( .A(n49075), .B(n48768), .Z(n49078) );
  XOR U49098 ( .A(n48826), .B(n49079), .Z(n48768) );
  AND U49099 ( .A(n1229), .B(n49080), .Z(n49079) );
  XOR U49100 ( .A(n48822), .B(n48826), .Z(n49080) );
  XNOR U49101 ( .A(n49081), .B(n49075), .Z(n49077) );
  IV U49102 ( .A(n48718), .Z(n49081) );
  XOR U49103 ( .A(n49082), .B(n49083), .Z(n48718) );
  AND U49104 ( .A(n1245), .B(n49084), .Z(n49083) );
  XOR U49105 ( .A(n49085), .B(n49086), .Z(n49075) );
  AND U49106 ( .A(n49087), .B(n49088), .Z(n49086) );
  XNOR U49107 ( .A(n49085), .B(n48778), .Z(n49088) );
  XOR U49108 ( .A(n48854), .B(n49089), .Z(n48778) );
  AND U49109 ( .A(n1229), .B(n49090), .Z(n49089) );
  XOR U49110 ( .A(n48850), .B(n48854), .Z(n49090) );
  XOR U49111 ( .A(n48727), .B(n49085), .Z(n49087) );
  XOR U49112 ( .A(n49091), .B(n49092), .Z(n48727) );
  AND U49113 ( .A(n1245), .B(n49093), .Z(n49092) );
  XOR U49114 ( .A(n49060), .B(n49094), .Z(n49085) );
  AND U49115 ( .A(n49095), .B(n49063), .Z(n49094) );
  XNOR U49116 ( .A(n48788), .B(n49060), .Z(n49063) );
  XOR U49117 ( .A(n48903), .B(n49096), .Z(n48788) );
  AND U49118 ( .A(n1229), .B(n49097), .Z(n49096) );
  XOR U49119 ( .A(n48899), .B(n48903), .Z(n49097) );
  XNOR U49120 ( .A(n49098), .B(n49060), .Z(n49095) );
  IV U49121 ( .A(n48735), .Z(n49098) );
  XOR U49122 ( .A(n49099), .B(n49100), .Z(n48735) );
  AND U49123 ( .A(n1245), .B(n49101), .Z(n49100) );
  XOR U49124 ( .A(n49102), .B(n49103), .Z(n49060) );
  AND U49125 ( .A(n49104), .B(n49105), .Z(n49103) );
  XNOR U49126 ( .A(n49102), .B(n48796), .Z(n49105) );
  XOR U49127 ( .A(n49000), .B(n49106), .Z(n48796) );
  AND U49128 ( .A(n1229), .B(n49107), .Z(n49106) );
  XOR U49129 ( .A(n48996), .B(n49000), .Z(n49107) );
  XNOR U49130 ( .A(n49108), .B(n49102), .Z(n49104) );
  IV U49131 ( .A(n48745), .Z(n49108) );
  XOR U49132 ( .A(n49109), .B(n49110), .Z(n48745) );
  AND U49133 ( .A(n1245), .B(n49111), .Z(n49110) );
  AND U49134 ( .A(n49064), .B(n49045), .Z(n49102) );
  XNOR U49135 ( .A(n49112), .B(n49113), .Z(n49045) );
  AND U49136 ( .A(n1229), .B(n49022), .Z(n49113) );
  XNOR U49137 ( .A(n49020), .B(n49112), .Z(n49022) );
  XNOR U49138 ( .A(n49114), .B(n49115), .Z(n1229) );
  NOR U49139 ( .A(n49116), .B(n49117), .Z(n49115) );
  XNOR U49140 ( .A(n49118), .B(n49028), .Z(n49117) );
  IV U49141 ( .A(n49072), .Z(n49028) );
  NOR U49142 ( .A(n49073), .B(n49074), .Z(n49072) );
  AND U49143 ( .A(n49118), .B(n48808), .Z(n49116) );
  IV U49144 ( .A(n49071), .Z(n48808) );
  AND U49145 ( .A(n49119), .B(n49120), .Z(n49071) );
  IV U49146 ( .A(n49121), .Z(n49119) );
  IV U49147 ( .A(n49114), .Z(n49118) );
  XOR U49148 ( .A(n49122), .B(n49123), .Z(n49114) );
  AND U49149 ( .A(n49124), .B(n49125), .Z(n49123) );
  XNOR U49150 ( .A(n49122), .B(n48822), .Z(n49125) );
  IV U49151 ( .A(n48825), .Z(n48822) );
  XOR U49152 ( .A(n49126), .B(n49127), .Z(n48825) );
  AND U49153 ( .A(n1233), .B(n49128), .Z(n49127) );
  XOR U49154 ( .A(n49129), .B(n49126), .Z(n49128) );
  XOR U49155 ( .A(n48826), .B(n49122), .Z(n49124) );
  XOR U49156 ( .A(n49130), .B(n49131), .Z(n48826) );
  AND U49157 ( .A(n1241), .B(n49084), .Z(n49131) );
  XOR U49158 ( .A(n49130), .B(n49082), .Z(n49084) );
  XOR U49159 ( .A(n49132), .B(n49133), .Z(n49122) );
  AND U49160 ( .A(n49134), .B(n49135), .Z(n49133) );
  XNOR U49161 ( .A(n49132), .B(n48850), .Z(n49135) );
  IV U49162 ( .A(n48853), .Z(n48850) );
  XOR U49163 ( .A(n49136), .B(n49137), .Z(n48853) );
  AND U49164 ( .A(n1233), .B(n49138), .Z(n49137) );
  XNOR U49165 ( .A(n49139), .B(n49136), .Z(n49138) );
  XOR U49166 ( .A(n48854), .B(n49132), .Z(n49134) );
  XOR U49167 ( .A(n49140), .B(n49141), .Z(n48854) );
  AND U49168 ( .A(n1241), .B(n49093), .Z(n49141) );
  XOR U49169 ( .A(n49140), .B(n49091), .Z(n49093) );
  XOR U49170 ( .A(n49142), .B(n49143), .Z(n49132) );
  AND U49171 ( .A(n49144), .B(n49145), .Z(n49143) );
  XNOR U49172 ( .A(n49142), .B(n48899), .Z(n49145) );
  IV U49173 ( .A(n48902), .Z(n48899) );
  XOR U49174 ( .A(n49146), .B(n49147), .Z(n48902) );
  AND U49175 ( .A(n1233), .B(n49148), .Z(n49147) );
  XOR U49176 ( .A(n49149), .B(n49146), .Z(n49148) );
  XOR U49177 ( .A(n48903), .B(n49142), .Z(n49144) );
  XOR U49178 ( .A(n49150), .B(n49151), .Z(n48903) );
  AND U49179 ( .A(n1241), .B(n49101), .Z(n49151) );
  XOR U49180 ( .A(n49150), .B(n49099), .Z(n49101) );
  XOR U49181 ( .A(n49041), .B(n49152), .Z(n49142) );
  AND U49182 ( .A(n49043), .B(n49153), .Z(n49152) );
  XNOR U49183 ( .A(n49041), .B(n48996), .Z(n49153) );
  IV U49184 ( .A(n48999), .Z(n48996) );
  XOR U49185 ( .A(n49154), .B(n49155), .Z(n48999) );
  AND U49186 ( .A(n1233), .B(n49156), .Z(n49155) );
  XNOR U49187 ( .A(n49157), .B(n49154), .Z(n49156) );
  XOR U49188 ( .A(n49000), .B(n49041), .Z(n49043) );
  XOR U49189 ( .A(n49158), .B(n49159), .Z(n49000) );
  AND U49190 ( .A(n1241), .B(n49111), .Z(n49159) );
  XOR U49191 ( .A(n49158), .B(n49109), .Z(n49111) );
  AND U49192 ( .A(n49112), .B(n49020), .Z(n49041) );
  XNOR U49193 ( .A(n49160), .B(n49161), .Z(n49020) );
  AND U49194 ( .A(n1233), .B(n49162), .Z(n49161) );
  XNOR U49195 ( .A(n49163), .B(n49160), .Z(n49162) );
  XNOR U49196 ( .A(n49164), .B(n49165), .Z(n1233) );
  NOR U49197 ( .A(n49166), .B(n49167), .Z(n49165) );
  XNOR U49198 ( .A(n49164), .B(n49121), .Z(n49167) );
  NOR U49199 ( .A(n49168), .B(n49169), .Z(n49121) );
  NOR U49200 ( .A(n49164), .B(n49120), .Z(n49166) );
  AND U49201 ( .A(n49170), .B(n49171), .Z(n49120) );
  XOR U49202 ( .A(n49172), .B(n49173), .Z(n49164) );
  AND U49203 ( .A(n49174), .B(n49175), .Z(n49173) );
  XNOR U49204 ( .A(n49172), .B(n49170), .Z(n49175) );
  IV U49205 ( .A(n49129), .Z(n49170) );
  XOR U49206 ( .A(n49176), .B(n49177), .Z(n49129) );
  XOR U49207 ( .A(n49178), .B(n49171), .Z(n49177) );
  AND U49208 ( .A(n49139), .B(n49179), .Z(n49171) );
  AND U49209 ( .A(n49180), .B(n49181), .Z(n49178) );
  XOR U49210 ( .A(n49182), .B(n49176), .Z(n49180) );
  XNOR U49211 ( .A(n49126), .B(n49172), .Z(n49174) );
  XNOR U49212 ( .A(n49183), .B(n49184), .Z(n49126) );
  AND U49213 ( .A(n1237), .B(n49185), .Z(n49184) );
  XNOR U49214 ( .A(n49186), .B(n49187), .Z(n49185) );
  XOR U49215 ( .A(n49188), .B(n49189), .Z(n49172) );
  AND U49216 ( .A(n49190), .B(n49191), .Z(n49189) );
  XNOR U49217 ( .A(n49188), .B(n49139), .Z(n49191) );
  XOR U49218 ( .A(n49192), .B(n49181), .Z(n49139) );
  XNOR U49219 ( .A(n49193), .B(n49176), .Z(n49181) );
  XOR U49220 ( .A(n49194), .B(n49195), .Z(n49176) );
  AND U49221 ( .A(n49196), .B(n49197), .Z(n49195) );
  XOR U49222 ( .A(n49198), .B(n49194), .Z(n49196) );
  XNOR U49223 ( .A(n49199), .B(n49200), .Z(n49193) );
  AND U49224 ( .A(n49201), .B(n49202), .Z(n49200) );
  XOR U49225 ( .A(n49199), .B(n49203), .Z(n49201) );
  XNOR U49226 ( .A(n49182), .B(n49179), .Z(n49192) );
  AND U49227 ( .A(n49204), .B(n49205), .Z(n49179) );
  XOR U49228 ( .A(n49206), .B(n49207), .Z(n49182) );
  AND U49229 ( .A(n49208), .B(n49209), .Z(n49207) );
  XOR U49230 ( .A(n49206), .B(n49210), .Z(n49208) );
  XNOR U49231 ( .A(n49136), .B(n49188), .Z(n49190) );
  XNOR U49232 ( .A(n49211), .B(n49212), .Z(n49136) );
  AND U49233 ( .A(n1237), .B(n49213), .Z(n49212) );
  XNOR U49234 ( .A(n49214), .B(n49215), .Z(n49213) );
  XOR U49235 ( .A(n49216), .B(n49217), .Z(n49188) );
  AND U49236 ( .A(n49218), .B(n49219), .Z(n49217) );
  XNOR U49237 ( .A(n49216), .B(n49204), .Z(n49219) );
  IV U49238 ( .A(n49149), .Z(n49204) );
  XNOR U49239 ( .A(n49220), .B(n49197), .Z(n49149) );
  XNOR U49240 ( .A(n49221), .B(n49203), .Z(n49197) );
  XOR U49241 ( .A(n49222), .B(n49223), .Z(n49203) );
  AND U49242 ( .A(n49224), .B(n49225), .Z(n49223) );
  XOR U49243 ( .A(n49222), .B(n49226), .Z(n49224) );
  XNOR U49244 ( .A(n49202), .B(n49194), .Z(n49221) );
  XOR U49245 ( .A(n49227), .B(n49228), .Z(n49194) );
  AND U49246 ( .A(n49229), .B(n49230), .Z(n49228) );
  XNOR U49247 ( .A(n49231), .B(n49227), .Z(n49229) );
  XNOR U49248 ( .A(n49232), .B(n49199), .Z(n49202) );
  XOR U49249 ( .A(n49233), .B(n49234), .Z(n49199) );
  AND U49250 ( .A(n49235), .B(n49236), .Z(n49234) );
  XOR U49251 ( .A(n49233), .B(n49237), .Z(n49235) );
  XNOR U49252 ( .A(n49238), .B(n49239), .Z(n49232) );
  AND U49253 ( .A(n49240), .B(n49241), .Z(n49239) );
  XNOR U49254 ( .A(n49238), .B(n49242), .Z(n49240) );
  XNOR U49255 ( .A(n49198), .B(n49205), .Z(n49220) );
  AND U49256 ( .A(n49157), .B(n49243), .Z(n49205) );
  XOR U49257 ( .A(n49210), .B(n49209), .Z(n49198) );
  XNOR U49258 ( .A(n49244), .B(n49206), .Z(n49209) );
  XOR U49259 ( .A(n49245), .B(n49246), .Z(n49206) );
  AND U49260 ( .A(n49247), .B(n49248), .Z(n49246) );
  XOR U49261 ( .A(n49245), .B(n49249), .Z(n49247) );
  XNOR U49262 ( .A(n49250), .B(n49251), .Z(n49244) );
  AND U49263 ( .A(n49252), .B(n49253), .Z(n49251) );
  XOR U49264 ( .A(n49250), .B(n49254), .Z(n49252) );
  XOR U49265 ( .A(n49255), .B(n49256), .Z(n49210) );
  AND U49266 ( .A(n49257), .B(n49258), .Z(n49256) );
  XOR U49267 ( .A(n49255), .B(n49259), .Z(n49257) );
  XNOR U49268 ( .A(n49146), .B(n49216), .Z(n49218) );
  XNOR U49269 ( .A(n49260), .B(n49261), .Z(n49146) );
  AND U49270 ( .A(n1237), .B(n49262), .Z(n49261) );
  XNOR U49271 ( .A(n49263), .B(n49264), .Z(n49262) );
  XOR U49272 ( .A(n49265), .B(n49266), .Z(n49216) );
  AND U49273 ( .A(n49267), .B(n49268), .Z(n49266) );
  XNOR U49274 ( .A(n49265), .B(n49157), .Z(n49268) );
  XOR U49275 ( .A(n49269), .B(n49230), .Z(n49157) );
  XNOR U49276 ( .A(n49270), .B(n49237), .Z(n49230) );
  XOR U49277 ( .A(n49226), .B(n49225), .Z(n49237) );
  XNOR U49278 ( .A(n49271), .B(n49222), .Z(n49225) );
  XOR U49279 ( .A(n49272), .B(n49273), .Z(n49222) );
  AND U49280 ( .A(n49274), .B(n49275), .Z(n49273) );
  XNOR U49281 ( .A(n49276), .B(n49277), .Z(n49274) );
  IV U49282 ( .A(n49272), .Z(n49276) );
  XNOR U49283 ( .A(n49278), .B(n49279), .Z(n49271) );
  NOR U49284 ( .A(n49280), .B(n49281), .Z(n49279) );
  XNOR U49285 ( .A(n49278), .B(n49282), .Z(n49280) );
  XOR U49286 ( .A(n49283), .B(n49284), .Z(n49226) );
  NOR U49287 ( .A(n49285), .B(n49286), .Z(n49284) );
  XNOR U49288 ( .A(n49283), .B(n49287), .Z(n49285) );
  XNOR U49289 ( .A(n49236), .B(n49227), .Z(n49270) );
  XOR U49290 ( .A(n49288), .B(n49289), .Z(n49227) );
  AND U49291 ( .A(n49290), .B(n49291), .Z(n49289) );
  XOR U49292 ( .A(n49288), .B(n49292), .Z(n49290) );
  XOR U49293 ( .A(n49293), .B(n49242), .Z(n49236) );
  XOR U49294 ( .A(n49294), .B(n49295), .Z(n49242) );
  NOR U49295 ( .A(n49296), .B(n49297), .Z(n49295) );
  XOR U49296 ( .A(n49294), .B(n49298), .Z(n49296) );
  XNOR U49297 ( .A(n49241), .B(n49233), .Z(n49293) );
  XOR U49298 ( .A(n49299), .B(n49300), .Z(n49233) );
  AND U49299 ( .A(n49301), .B(n49302), .Z(n49300) );
  XOR U49300 ( .A(n49299), .B(n49303), .Z(n49301) );
  XNOR U49301 ( .A(n49304), .B(n49238), .Z(n49241) );
  XOR U49302 ( .A(n49305), .B(n49306), .Z(n49238) );
  AND U49303 ( .A(n49307), .B(n49308), .Z(n49306) );
  XNOR U49304 ( .A(n49309), .B(n49310), .Z(n49307) );
  IV U49305 ( .A(n49305), .Z(n49309) );
  XNOR U49306 ( .A(n49311), .B(n49312), .Z(n49304) );
  NOR U49307 ( .A(n49313), .B(n49314), .Z(n49312) );
  XNOR U49308 ( .A(n49311), .B(n49315), .Z(n49313) );
  XOR U49309 ( .A(n49231), .B(n49243), .Z(n49269) );
  NOR U49310 ( .A(n49163), .B(n49316), .Z(n49243) );
  XNOR U49311 ( .A(n49249), .B(n49248), .Z(n49231) );
  XNOR U49312 ( .A(n49317), .B(n49254), .Z(n49248) );
  XNOR U49313 ( .A(n49318), .B(n49319), .Z(n49254) );
  NOR U49314 ( .A(n49320), .B(n49321), .Z(n49319) );
  XOR U49315 ( .A(n49318), .B(n49322), .Z(n49320) );
  XNOR U49316 ( .A(n49253), .B(n49245), .Z(n49317) );
  XOR U49317 ( .A(n49323), .B(n49324), .Z(n49245) );
  AND U49318 ( .A(n49325), .B(n49326), .Z(n49324) );
  XOR U49319 ( .A(n49323), .B(n49327), .Z(n49325) );
  XNOR U49320 ( .A(n49328), .B(n49250), .Z(n49253) );
  XOR U49321 ( .A(n49329), .B(n49330), .Z(n49250) );
  AND U49322 ( .A(n49331), .B(n49332), .Z(n49330) );
  XNOR U49323 ( .A(n49333), .B(n49334), .Z(n49331) );
  IV U49324 ( .A(n49329), .Z(n49333) );
  XNOR U49325 ( .A(n49335), .B(n49336), .Z(n49328) );
  NOR U49326 ( .A(n49337), .B(n49338), .Z(n49336) );
  XNOR U49327 ( .A(n49335), .B(n49339), .Z(n49337) );
  XOR U49328 ( .A(n49259), .B(n49258), .Z(n49249) );
  XNOR U49329 ( .A(n49340), .B(n49255), .Z(n49258) );
  XOR U49330 ( .A(n49341), .B(n49342), .Z(n49255) );
  AND U49331 ( .A(n49343), .B(n49344), .Z(n49342) );
  XNOR U49332 ( .A(n49345), .B(n49346), .Z(n49343) );
  IV U49333 ( .A(n49341), .Z(n49345) );
  XNOR U49334 ( .A(n49347), .B(n49348), .Z(n49340) );
  NOR U49335 ( .A(n49349), .B(n49350), .Z(n49348) );
  XNOR U49336 ( .A(n49347), .B(n49351), .Z(n49349) );
  XOR U49337 ( .A(n49352), .B(n49353), .Z(n49259) );
  NOR U49338 ( .A(n49354), .B(n49355), .Z(n49353) );
  XNOR U49339 ( .A(n49352), .B(n49356), .Z(n49354) );
  XNOR U49340 ( .A(n49154), .B(n49265), .Z(n49267) );
  XNOR U49341 ( .A(n49357), .B(n49358), .Z(n49154) );
  AND U49342 ( .A(n1237), .B(n49359), .Z(n49358) );
  XNOR U49343 ( .A(n49360), .B(n49361), .Z(n49359) );
  AND U49344 ( .A(n49160), .B(n49163), .Z(n49265) );
  XOR U49345 ( .A(n49362), .B(n49316), .Z(n49163) );
  XNOR U49346 ( .A(p_input[1856]), .B(p_input[2048]), .Z(n49316) );
  XNOR U49347 ( .A(n49292), .B(n49291), .Z(n49362) );
  XNOR U49348 ( .A(n49363), .B(n49303), .Z(n49291) );
  XOR U49349 ( .A(n49277), .B(n49275), .Z(n49303) );
  XNOR U49350 ( .A(n49364), .B(n49282), .Z(n49275) );
  XOR U49351 ( .A(p_input[1880]), .B(p_input[2072]), .Z(n49282) );
  XOR U49352 ( .A(n49272), .B(n49281), .Z(n49364) );
  XOR U49353 ( .A(n49365), .B(n49278), .Z(n49281) );
  XOR U49354 ( .A(p_input[1878]), .B(p_input[2070]), .Z(n49278) );
  XOR U49355 ( .A(p_input[1879]), .B(n29410), .Z(n49365) );
  XOR U49356 ( .A(p_input[1874]), .B(p_input[2066]), .Z(n49272) );
  XNOR U49357 ( .A(n49287), .B(n49286), .Z(n49277) );
  XOR U49358 ( .A(n49366), .B(n49283), .Z(n49286) );
  XOR U49359 ( .A(p_input[1875]), .B(p_input[2067]), .Z(n49283) );
  XOR U49360 ( .A(p_input[1876]), .B(n29412), .Z(n49366) );
  XOR U49361 ( .A(p_input[1877]), .B(p_input[2069]), .Z(n49287) );
  XOR U49362 ( .A(n49302), .B(n49367), .Z(n49363) );
  IV U49363 ( .A(n49288), .Z(n49367) );
  XOR U49364 ( .A(p_input[1857]), .B(p_input[2049]), .Z(n49288) );
  XNOR U49365 ( .A(n49368), .B(n49310), .Z(n49302) );
  XNOR U49366 ( .A(n49298), .B(n49297), .Z(n49310) );
  XNOR U49367 ( .A(n49369), .B(n49294), .Z(n49297) );
  XNOR U49368 ( .A(p_input[1882]), .B(p_input[2074]), .Z(n49294) );
  XOR U49369 ( .A(p_input[1883]), .B(n29415), .Z(n49369) );
  XOR U49370 ( .A(p_input[1884]), .B(p_input[2076]), .Z(n49298) );
  XOR U49371 ( .A(n49308), .B(n49370), .Z(n49368) );
  IV U49372 ( .A(n49299), .Z(n49370) );
  XOR U49373 ( .A(p_input[1873]), .B(p_input[2065]), .Z(n49299) );
  XNOR U49374 ( .A(n49371), .B(n49315), .Z(n49308) );
  XNOR U49375 ( .A(p_input[1887]), .B(n29418), .Z(n49315) );
  XOR U49376 ( .A(n49305), .B(n49314), .Z(n49371) );
  XOR U49377 ( .A(n49372), .B(n49311), .Z(n49314) );
  XOR U49378 ( .A(p_input[1885]), .B(p_input[2077]), .Z(n49311) );
  XOR U49379 ( .A(p_input[1886]), .B(n29420), .Z(n49372) );
  XOR U49380 ( .A(p_input[1881]), .B(p_input[2073]), .Z(n49305) );
  XOR U49381 ( .A(n49327), .B(n49326), .Z(n49292) );
  XNOR U49382 ( .A(n49373), .B(n49334), .Z(n49326) );
  XNOR U49383 ( .A(n49322), .B(n49321), .Z(n49334) );
  XNOR U49384 ( .A(n49374), .B(n49318), .Z(n49321) );
  XNOR U49385 ( .A(p_input[1867]), .B(p_input[2059]), .Z(n49318) );
  XOR U49386 ( .A(p_input[1868]), .B(n28329), .Z(n49374) );
  XOR U49387 ( .A(p_input[1869]), .B(p_input[2061]), .Z(n49322) );
  XOR U49388 ( .A(n49332), .B(n49375), .Z(n49373) );
  IV U49389 ( .A(n49323), .Z(n49375) );
  XOR U49390 ( .A(p_input[1858]), .B(p_input[2050]), .Z(n49323) );
  XNOR U49391 ( .A(n49376), .B(n49339), .Z(n49332) );
  XNOR U49392 ( .A(p_input[1872]), .B(n28332), .Z(n49339) );
  XOR U49393 ( .A(n49329), .B(n49338), .Z(n49376) );
  XOR U49394 ( .A(n49377), .B(n49335), .Z(n49338) );
  XOR U49395 ( .A(p_input[1870]), .B(p_input[2062]), .Z(n49335) );
  XOR U49396 ( .A(p_input[1871]), .B(n28334), .Z(n49377) );
  XOR U49397 ( .A(p_input[1866]), .B(p_input[2058]), .Z(n49329) );
  XOR U49398 ( .A(n49346), .B(n49344), .Z(n49327) );
  XNOR U49399 ( .A(n49378), .B(n49351), .Z(n49344) );
  XOR U49400 ( .A(p_input[1865]), .B(p_input[2057]), .Z(n49351) );
  XOR U49401 ( .A(n49341), .B(n49350), .Z(n49378) );
  XOR U49402 ( .A(n49379), .B(n49347), .Z(n49350) );
  XOR U49403 ( .A(p_input[1863]), .B(p_input[2055]), .Z(n49347) );
  XOR U49404 ( .A(p_input[1864]), .B(n29427), .Z(n49379) );
  XOR U49405 ( .A(p_input[1859]), .B(p_input[2051]), .Z(n49341) );
  XNOR U49406 ( .A(n49356), .B(n49355), .Z(n49346) );
  XOR U49407 ( .A(n49380), .B(n49352), .Z(n49355) );
  XOR U49408 ( .A(p_input[1860]), .B(p_input[2052]), .Z(n49352) );
  XOR U49409 ( .A(p_input[1861]), .B(n29429), .Z(n49380) );
  XOR U49410 ( .A(p_input[1862]), .B(p_input[2054]), .Z(n49356) );
  XNOR U49411 ( .A(n49381), .B(n49382), .Z(n49160) );
  AND U49412 ( .A(n1237), .B(n49383), .Z(n49382) );
  XNOR U49413 ( .A(n49384), .B(n49385), .Z(n1237) );
  NOR U49414 ( .A(n49386), .B(n49387), .Z(n49385) );
  XNOR U49415 ( .A(n49384), .B(n49388), .Z(n49387) );
  NOR U49416 ( .A(n49384), .B(n49169), .Z(n49386) );
  XOR U49417 ( .A(n49389), .B(n49390), .Z(n49384) );
  AND U49418 ( .A(n49391), .B(n49392), .Z(n49390) );
  XOR U49419 ( .A(n49186), .B(n49389), .Z(n49392) );
  XOR U49420 ( .A(n49389), .B(n49187), .Z(n49391) );
  XOR U49421 ( .A(n49393), .B(n49394), .Z(n49389) );
  AND U49422 ( .A(n49395), .B(n49396), .Z(n49394) );
  XOR U49423 ( .A(n49214), .B(n49393), .Z(n49396) );
  XOR U49424 ( .A(n49393), .B(n49215), .Z(n49395) );
  XOR U49425 ( .A(n49397), .B(n49398), .Z(n49393) );
  AND U49426 ( .A(n49399), .B(n49400), .Z(n49398) );
  XOR U49427 ( .A(n49263), .B(n49397), .Z(n49400) );
  XOR U49428 ( .A(n49397), .B(n49264), .Z(n49399) );
  XOR U49429 ( .A(n49401), .B(n49402), .Z(n49397) );
  AND U49430 ( .A(n49403), .B(n49404), .Z(n49402) );
  XOR U49431 ( .A(n49401), .B(n49360), .Z(n49404) );
  XNOR U49432 ( .A(n49405), .B(n49406), .Z(n49112) );
  AND U49433 ( .A(n1241), .B(n49407), .Z(n49406) );
  XNOR U49434 ( .A(n49408), .B(n49409), .Z(n1241) );
  NOR U49435 ( .A(n49410), .B(n49411), .Z(n49409) );
  XOR U49436 ( .A(n49074), .B(n49408), .Z(n49411) );
  NOR U49437 ( .A(n49408), .B(n49073), .Z(n49410) );
  XOR U49438 ( .A(n49412), .B(n49413), .Z(n49408) );
  AND U49439 ( .A(n49414), .B(n49415), .Z(n49413) );
  XNOR U49440 ( .A(n49130), .B(n49412), .Z(n49415) );
  XOR U49441 ( .A(n49412), .B(n49082), .Z(n49414) );
  XOR U49442 ( .A(n49416), .B(n49417), .Z(n49412) );
  AND U49443 ( .A(n49418), .B(n49419), .Z(n49417) );
  XNOR U49444 ( .A(n49140), .B(n49416), .Z(n49419) );
  XOR U49445 ( .A(n49416), .B(n49091), .Z(n49418) );
  XOR U49446 ( .A(n49420), .B(n49421), .Z(n49416) );
  AND U49447 ( .A(n49422), .B(n49423), .Z(n49421) );
  XOR U49448 ( .A(n49420), .B(n49099), .Z(n49422) );
  XOR U49449 ( .A(n49424), .B(n49425), .Z(n49064) );
  AND U49450 ( .A(n1245), .B(n49407), .Z(n49425) );
  XNOR U49451 ( .A(n49405), .B(n49424), .Z(n49407) );
  XNOR U49452 ( .A(n49426), .B(n49427), .Z(n1245) );
  NOR U49453 ( .A(n49428), .B(n49429), .Z(n49427) );
  XNOR U49454 ( .A(n49074), .B(n49430), .Z(n49429) );
  IV U49455 ( .A(n49426), .Z(n49430) );
  AND U49456 ( .A(n49431), .B(n49432), .Z(n49074) );
  NOR U49457 ( .A(n49426), .B(n49073), .Z(n49428) );
  AND U49458 ( .A(n49169), .B(n49168), .Z(n49073) );
  IV U49459 ( .A(n49388), .Z(n49168) );
  XOR U49460 ( .A(n49433), .B(n49434), .Z(n49426) );
  AND U49461 ( .A(n49435), .B(n49436), .Z(n49434) );
  XNOR U49462 ( .A(n49433), .B(n49130), .Z(n49436) );
  XOR U49463 ( .A(n49187), .B(n49437), .Z(n49130) );
  AND U49464 ( .A(n1248), .B(n49438), .Z(n49437) );
  XOR U49465 ( .A(n49183), .B(n49187), .Z(n49438) );
  XNOR U49466 ( .A(n49439), .B(n49433), .Z(n49435) );
  IV U49467 ( .A(n49082), .Z(n49439) );
  XOR U49468 ( .A(n49440), .B(n49441), .Z(n49082) );
  AND U49469 ( .A(n1264), .B(n49442), .Z(n49441) );
  XOR U49470 ( .A(n49443), .B(n49444), .Z(n49433) );
  AND U49471 ( .A(n49445), .B(n49446), .Z(n49444) );
  XNOR U49472 ( .A(n49443), .B(n49140), .Z(n49446) );
  XOR U49473 ( .A(n49215), .B(n49447), .Z(n49140) );
  AND U49474 ( .A(n1248), .B(n49448), .Z(n49447) );
  XOR U49475 ( .A(n49211), .B(n49215), .Z(n49448) );
  XOR U49476 ( .A(n49091), .B(n49443), .Z(n49445) );
  XOR U49477 ( .A(n49449), .B(n49450), .Z(n49091) );
  AND U49478 ( .A(n1264), .B(n49451), .Z(n49450) );
  XOR U49479 ( .A(n49420), .B(n49452), .Z(n49443) );
  AND U49480 ( .A(n49453), .B(n49423), .Z(n49452) );
  XNOR U49481 ( .A(n49150), .B(n49420), .Z(n49423) );
  XOR U49482 ( .A(n49264), .B(n49454), .Z(n49150) );
  AND U49483 ( .A(n1248), .B(n49455), .Z(n49454) );
  XOR U49484 ( .A(n49260), .B(n49264), .Z(n49455) );
  XNOR U49485 ( .A(n49456), .B(n49420), .Z(n49453) );
  IV U49486 ( .A(n49099), .Z(n49456) );
  XOR U49487 ( .A(n49457), .B(n49458), .Z(n49099) );
  AND U49488 ( .A(n1264), .B(n49459), .Z(n49458) );
  XOR U49489 ( .A(n49460), .B(n49461), .Z(n49420) );
  AND U49490 ( .A(n49462), .B(n49463), .Z(n49461) );
  XNOR U49491 ( .A(n49460), .B(n49158), .Z(n49463) );
  XOR U49492 ( .A(n49361), .B(n49464), .Z(n49158) );
  AND U49493 ( .A(n1248), .B(n49465), .Z(n49464) );
  XOR U49494 ( .A(n49357), .B(n49361), .Z(n49465) );
  XNOR U49495 ( .A(n49466), .B(n49460), .Z(n49462) );
  IV U49496 ( .A(n49109), .Z(n49466) );
  XOR U49497 ( .A(n49467), .B(n49468), .Z(n49109) );
  AND U49498 ( .A(n1264), .B(n49469), .Z(n49468) );
  AND U49499 ( .A(n49424), .B(n49405), .Z(n49460) );
  XNOR U49500 ( .A(n49470), .B(n49471), .Z(n49405) );
  AND U49501 ( .A(n1248), .B(n49383), .Z(n49471) );
  XNOR U49502 ( .A(n49381), .B(n49470), .Z(n49383) );
  XNOR U49503 ( .A(n49472), .B(n49473), .Z(n1248) );
  NOR U49504 ( .A(n49474), .B(n49475), .Z(n49473) );
  XNOR U49505 ( .A(n49472), .B(n49388), .Z(n49475) );
  NOR U49506 ( .A(n49431), .B(n49432), .Z(n49388) );
  NOR U49507 ( .A(n49472), .B(n49169), .Z(n49474) );
  AND U49508 ( .A(n49476), .B(n49477), .Z(n49169) );
  IV U49509 ( .A(n49478), .Z(n49476) );
  XOR U49510 ( .A(n49479), .B(n49480), .Z(n49472) );
  AND U49511 ( .A(n49481), .B(n49482), .Z(n49480) );
  XNOR U49512 ( .A(n49479), .B(n49183), .Z(n49482) );
  IV U49513 ( .A(n49186), .Z(n49183) );
  XOR U49514 ( .A(n49483), .B(n49484), .Z(n49186) );
  AND U49515 ( .A(n1252), .B(n49485), .Z(n49484) );
  XOR U49516 ( .A(n49486), .B(n49483), .Z(n49485) );
  XOR U49517 ( .A(n49187), .B(n49479), .Z(n49481) );
  XOR U49518 ( .A(n49487), .B(n49488), .Z(n49187) );
  AND U49519 ( .A(n1260), .B(n49442), .Z(n49488) );
  XOR U49520 ( .A(n49487), .B(n49440), .Z(n49442) );
  XOR U49521 ( .A(n49489), .B(n49490), .Z(n49479) );
  AND U49522 ( .A(n49491), .B(n49492), .Z(n49490) );
  XNOR U49523 ( .A(n49489), .B(n49211), .Z(n49492) );
  IV U49524 ( .A(n49214), .Z(n49211) );
  XOR U49525 ( .A(n49493), .B(n49494), .Z(n49214) );
  AND U49526 ( .A(n1252), .B(n49495), .Z(n49494) );
  XNOR U49527 ( .A(n49496), .B(n49493), .Z(n49495) );
  XOR U49528 ( .A(n49215), .B(n49489), .Z(n49491) );
  XOR U49529 ( .A(n49497), .B(n49498), .Z(n49215) );
  AND U49530 ( .A(n1260), .B(n49451), .Z(n49498) );
  XOR U49531 ( .A(n49497), .B(n49449), .Z(n49451) );
  XOR U49532 ( .A(n49499), .B(n49500), .Z(n49489) );
  AND U49533 ( .A(n49501), .B(n49502), .Z(n49500) );
  XNOR U49534 ( .A(n49499), .B(n49260), .Z(n49502) );
  IV U49535 ( .A(n49263), .Z(n49260) );
  XOR U49536 ( .A(n49503), .B(n49504), .Z(n49263) );
  AND U49537 ( .A(n1252), .B(n49505), .Z(n49504) );
  XOR U49538 ( .A(n49506), .B(n49503), .Z(n49505) );
  XOR U49539 ( .A(n49264), .B(n49499), .Z(n49501) );
  XOR U49540 ( .A(n49507), .B(n49508), .Z(n49264) );
  AND U49541 ( .A(n1260), .B(n49459), .Z(n49508) );
  XOR U49542 ( .A(n49507), .B(n49457), .Z(n49459) );
  XOR U49543 ( .A(n49401), .B(n49509), .Z(n49499) );
  AND U49544 ( .A(n49403), .B(n49510), .Z(n49509) );
  XNOR U49545 ( .A(n49401), .B(n49357), .Z(n49510) );
  IV U49546 ( .A(n49360), .Z(n49357) );
  XOR U49547 ( .A(n49511), .B(n49512), .Z(n49360) );
  AND U49548 ( .A(n1252), .B(n49513), .Z(n49512) );
  XNOR U49549 ( .A(n49514), .B(n49511), .Z(n49513) );
  XOR U49550 ( .A(n49361), .B(n49401), .Z(n49403) );
  XOR U49551 ( .A(n49515), .B(n49516), .Z(n49361) );
  AND U49552 ( .A(n1260), .B(n49469), .Z(n49516) );
  XOR U49553 ( .A(n49515), .B(n49467), .Z(n49469) );
  AND U49554 ( .A(n49470), .B(n49381), .Z(n49401) );
  XNOR U49555 ( .A(n49517), .B(n49518), .Z(n49381) );
  AND U49556 ( .A(n1252), .B(n49519), .Z(n49518) );
  XNOR U49557 ( .A(n49520), .B(n49517), .Z(n49519) );
  XNOR U49558 ( .A(n49521), .B(n49522), .Z(n1252) );
  NOR U49559 ( .A(n49523), .B(n49524), .Z(n49522) );
  XNOR U49560 ( .A(n49521), .B(n49478), .Z(n49524) );
  NOR U49561 ( .A(n49525), .B(n49526), .Z(n49478) );
  NOR U49562 ( .A(n49521), .B(n49477), .Z(n49523) );
  AND U49563 ( .A(n49527), .B(n49528), .Z(n49477) );
  XOR U49564 ( .A(n49529), .B(n49530), .Z(n49521) );
  AND U49565 ( .A(n49531), .B(n49532), .Z(n49530) );
  XNOR U49566 ( .A(n49529), .B(n49527), .Z(n49532) );
  IV U49567 ( .A(n49486), .Z(n49527) );
  XOR U49568 ( .A(n49533), .B(n49534), .Z(n49486) );
  XOR U49569 ( .A(n49535), .B(n49528), .Z(n49534) );
  AND U49570 ( .A(n49496), .B(n49536), .Z(n49528) );
  AND U49571 ( .A(n49537), .B(n49538), .Z(n49535) );
  XOR U49572 ( .A(n49539), .B(n49533), .Z(n49537) );
  XNOR U49573 ( .A(n49483), .B(n49529), .Z(n49531) );
  XNOR U49574 ( .A(n49540), .B(n49541), .Z(n49483) );
  AND U49575 ( .A(n1256), .B(n49542), .Z(n49541) );
  XNOR U49576 ( .A(n49543), .B(n49544), .Z(n49542) );
  XOR U49577 ( .A(n49545), .B(n49546), .Z(n49529) );
  AND U49578 ( .A(n49547), .B(n49548), .Z(n49546) );
  XNOR U49579 ( .A(n49545), .B(n49496), .Z(n49548) );
  XOR U49580 ( .A(n49549), .B(n49538), .Z(n49496) );
  XNOR U49581 ( .A(n49550), .B(n49533), .Z(n49538) );
  XOR U49582 ( .A(n49551), .B(n49552), .Z(n49533) );
  AND U49583 ( .A(n49553), .B(n49554), .Z(n49552) );
  XOR U49584 ( .A(n49555), .B(n49551), .Z(n49553) );
  XNOR U49585 ( .A(n49556), .B(n49557), .Z(n49550) );
  AND U49586 ( .A(n49558), .B(n49559), .Z(n49557) );
  XOR U49587 ( .A(n49556), .B(n49560), .Z(n49558) );
  XNOR U49588 ( .A(n49539), .B(n49536), .Z(n49549) );
  AND U49589 ( .A(n49561), .B(n49562), .Z(n49536) );
  XOR U49590 ( .A(n49563), .B(n49564), .Z(n49539) );
  AND U49591 ( .A(n49565), .B(n49566), .Z(n49564) );
  XOR U49592 ( .A(n49563), .B(n49567), .Z(n49565) );
  XNOR U49593 ( .A(n49493), .B(n49545), .Z(n49547) );
  XNOR U49594 ( .A(n49568), .B(n49569), .Z(n49493) );
  AND U49595 ( .A(n1256), .B(n49570), .Z(n49569) );
  XNOR U49596 ( .A(n49571), .B(n49572), .Z(n49570) );
  XOR U49597 ( .A(n49573), .B(n49574), .Z(n49545) );
  AND U49598 ( .A(n49575), .B(n49576), .Z(n49574) );
  XNOR U49599 ( .A(n49573), .B(n49561), .Z(n49576) );
  IV U49600 ( .A(n49506), .Z(n49561) );
  XNOR U49601 ( .A(n49577), .B(n49554), .Z(n49506) );
  XNOR U49602 ( .A(n49578), .B(n49560), .Z(n49554) );
  XOR U49603 ( .A(n49579), .B(n49580), .Z(n49560) );
  AND U49604 ( .A(n49581), .B(n49582), .Z(n49580) );
  XOR U49605 ( .A(n49579), .B(n49583), .Z(n49581) );
  XNOR U49606 ( .A(n49559), .B(n49551), .Z(n49578) );
  XOR U49607 ( .A(n49584), .B(n49585), .Z(n49551) );
  AND U49608 ( .A(n49586), .B(n49587), .Z(n49585) );
  XNOR U49609 ( .A(n49588), .B(n49584), .Z(n49586) );
  XNOR U49610 ( .A(n49589), .B(n49556), .Z(n49559) );
  XOR U49611 ( .A(n49590), .B(n49591), .Z(n49556) );
  AND U49612 ( .A(n49592), .B(n49593), .Z(n49591) );
  XOR U49613 ( .A(n49590), .B(n49594), .Z(n49592) );
  XNOR U49614 ( .A(n49595), .B(n49596), .Z(n49589) );
  AND U49615 ( .A(n49597), .B(n49598), .Z(n49596) );
  XNOR U49616 ( .A(n49595), .B(n49599), .Z(n49597) );
  XNOR U49617 ( .A(n49555), .B(n49562), .Z(n49577) );
  AND U49618 ( .A(n49514), .B(n49600), .Z(n49562) );
  XOR U49619 ( .A(n49567), .B(n49566), .Z(n49555) );
  XNOR U49620 ( .A(n49601), .B(n49563), .Z(n49566) );
  XOR U49621 ( .A(n49602), .B(n49603), .Z(n49563) );
  AND U49622 ( .A(n49604), .B(n49605), .Z(n49603) );
  XOR U49623 ( .A(n49602), .B(n49606), .Z(n49604) );
  XNOR U49624 ( .A(n49607), .B(n49608), .Z(n49601) );
  AND U49625 ( .A(n49609), .B(n49610), .Z(n49608) );
  XOR U49626 ( .A(n49607), .B(n49611), .Z(n49609) );
  XOR U49627 ( .A(n49612), .B(n49613), .Z(n49567) );
  AND U49628 ( .A(n49614), .B(n49615), .Z(n49613) );
  XOR U49629 ( .A(n49612), .B(n49616), .Z(n49614) );
  XNOR U49630 ( .A(n49503), .B(n49573), .Z(n49575) );
  XNOR U49631 ( .A(n49617), .B(n49618), .Z(n49503) );
  AND U49632 ( .A(n1256), .B(n49619), .Z(n49618) );
  XNOR U49633 ( .A(n49620), .B(n49621), .Z(n49619) );
  XOR U49634 ( .A(n49622), .B(n49623), .Z(n49573) );
  AND U49635 ( .A(n49624), .B(n49625), .Z(n49623) );
  XNOR U49636 ( .A(n49622), .B(n49514), .Z(n49625) );
  XOR U49637 ( .A(n49626), .B(n49587), .Z(n49514) );
  XNOR U49638 ( .A(n49627), .B(n49594), .Z(n49587) );
  XOR U49639 ( .A(n49583), .B(n49582), .Z(n49594) );
  XNOR U49640 ( .A(n49628), .B(n49579), .Z(n49582) );
  XOR U49641 ( .A(n49629), .B(n49630), .Z(n49579) );
  AND U49642 ( .A(n49631), .B(n49632), .Z(n49630) );
  XNOR U49643 ( .A(n49633), .B(n49634), .Z(n49631) );
  IV U49644 ( .A(n49629), .Z(n49633) );
  XNOR U49645 ( .A(n49635), .B(n49636), .Z(n49628) );
  NOR U49646 ( .A(n49637), .B(n49638), .Z(n49636) );
  XNOR U49647 ( .A(n49635), .B(n49639), .Z(n49637) );
  XOR U49648 ( .A(n49640), .B(n49641), .Z(n49583) );
  NOR U49649 ( .A(n49642), .B(n49643), .Z(n49641) );
  XNOR U49650 ( .A(n49640), .B(n49644), .Z(n49642) );
  XNOR U49651 ( .A(n49593), .B(n49584), .Z(n49627) );
  XOR U49652 ( .A(n49645), .B(n49646), .Z(n49584) );
  AND U49653 ( .A(n49647), .B(n49648), .Z(n49646) );
  XOR U49654 ( .A(n49645), .B(n49649), .Z(n49647) );
  XOR U49655 ( .A(n49650), .B(n49599), .Z(n49593) );
  XOR U49656 ( .A(n49651), .B(n49652), .Z(n49599) );
  NOR U49657 ( .A(n49653), .B(n49654), .Z(n49652) );
  XOR U49658 ( .A(n49651), .B(n49655), .Z(n49653) );
  XNOR U49659 ( .A(n49598), .B(n49590), .Z(n49650) );
  XOR U49660 ( .A(n49656), .B(n49657), .Z(n49590) );
  AND U49661 ( .A(n49658), .B(n49659), .Z(n49657) );
  XOR U49662 ( .A(n49656), .B(n49660), .Z(n49658) );
  XNOR U49663 ( .A(n49661), .B(n49595), .Z(n49598) );
  XOR U49664 ( .A(n49662), .B(n49663), .Z(n49595) );
  AND U49665 ( .A(n49664), .B(n49665), .Z(n49663) );
  XNOR U49666 ( .A(n49666), .B(n49667), .Z(n49664) );
  IV U49667 ( .A(n49662), .Z(n49666) );
  XNOR U49668 ( .A(n49668), .B(n49669), .Z(n49661) );
  NOR U49669 ( .A(n49670), .B(n49671), .Z(n49669) );
  XNOR U49670 ( .A(n49668), .B(n49672), .Z(n49670) );
  XOR U49671 ( .A(n49588), .B(n49600), .Z(n49626) );
  NOR U49672 ( .A(n49520), .B(n49673), .Z(n49600) );
  XNOR U49673 ( .A(n49606), .B(n49605), .Z(n49588) );
  XNOR U49674 ( .A(n49674), .B(n49611), .Z(n49605) );
  XNOR U49675 ( .A(n49675), .B(n49676), .Z(n49611) );
  NOR U49676 ( .A(n49677), .B(n49678), .Z(n49676) );
  XOR U49677 ( .A(n49675), .B(n49679), .Z(n49677) );
  XNOR U49678 ( .A(n49610), .B(n49602), .Z(n49674) );
  XOR U49679 ( .A(n49680), .B(n49681), .Z(n49602) );
  AND U49680 ( .A(n49682), .B(n49683), .Z(n49681) );
  XOR U49681 ( .A(n49680), .B(n49684), .Z(n49682) );
  XNOR U49682 ( .A(n49685), .B(n49607), .Z(n49610) );
  XOR U49683 ( .A(n49686), .B(n49687), .Z(n49607) );
  AND U49684 ( .A(n49688), .B(n49689), .Z(n49687) );
  XNOR U49685 ( .A(n49690), .B(n49691), .Z(n49688) );
  IV U49686 ( .A(n49686), .Z(n49690) );
  XNOR U49687 ( .A(n49692), .B(n49693), .Z(n49685) );
  NOR U49688 ( .A(n49694), .B(n49695), .Z(n49693) );
  XNOR U49689 ( .A(n49692), .B(n49696), .Z(n49694) );
  XOR U49690 ( .A(n49616), .B(n49615), .Z(n49606) );
  XNOR U49691 ( .A(n49697), .B(n49612), .Z(n49615) );
  XOR U49692 ( .A(n49698), .B(n49699), .Z(n49612) );
  AND U49693 ( .A(n49700), .B(n49701), .Z(n49699) );
  XNOR U49694 ( .A(n49702), .B(n49703), .Z(n49700) );
  IV U49695 ( .A(n49698), .Z(n49702) );
  XNOR U49696 ( .A(n49704), .B(n49705), .Z(n49697) );
  NOR U49697 ( .A(n49706), .B(n49707), .Z(n49705) );
  XNOR U49698 ( .A(n49704), .B(n49708), .Z(n49706) );
  XOR U49699 ( .A(n49709), .B(n49710), .Z(n49616) );
  NOR U49700 ( .A(n49711), .B(n49712), .Z(n49710) );
  XNOR U49701 ( .A(n49709), .B(n49713), .Z(n49711) );
  XNOR U49702 ( .A(n49511), .B(n49622), .Z(n49624) );
  XNOR U49703 ( .A(n49714), .B(n49715), .Z(n49511) );
  AND U49704 ( .A(n1256), .B(n49716), .Z(n49715) );
  XNOR U49705 ( .A(n49717), .B(n49718), .Z(n49716) );
  AND U49706 ( .A(n49517), .B(n49520), .Z(n49622) );
  XOR U49707 ( .A(n49719), .B(n49673), .Z(n49520) );
  XNOR U49708 ( .A(p_input[1888]), .B(p_input[2048]), .Z(n49673) );
  XNOR U49709 ( .A(n49649), .B(n49648), .Z(n49719) );
  XNOR U49710 ( .A(n49720), .B(n49660), .Z(n49648) );
  XOR U49711 ( .A(n49634), .B(n49632), .Z(n49660) );
  XNOR U49712 ( .A(n49721), .B(n49639), .Z(n49632) );
  XOR U49713 ( .A(p_input[1912]), .B(p_input[2072]), .Z(n49639) );
  XOR U49714 ( .A(n49629), .B(n49638), .Z(n49721) );
  XOR U49715 ( .A(n49722), .B(n49635), .Z(n49638) );
  XOR U49716 ( .A(p_input[1910]), .B(p_input[2070]), .Z(n49635) );
  XOR U49717 ( .A(p_input[1911]), .B(n29410), .Z(n49722) );
  XOR U49718 ( .A(p_input[1906]), .B(p_input[2066]), .Z(n49629) );
  XNOR U49719 ( .A(n49644), .B(n49643), .Z(n49634) );
  XOR U49720 ( .A(n49723), .B(n49640), .Z(n49643) );
  XOR U49721 ( .A(p_input[1907]), .B(p_input[2067]), .Z(n49640) );
  XOR U49722 ( .A(p_input[1908]), .B(n29412), .Z(n49723) );
  XOR U49723 ( .A(p_input[1909]), .B(p_input[2069]), .Z(n49644) );
  XOR U49724 ( .A(n49659), .B(n49724), .Z(n49720) );
  IV U49725 ( .A(n49645), .Z(n49724) );
  XOR U49726 ( .A(p_input[1889]), .B(p_input[2049]), .Z(n49645) );
  XNOR U49727 ( .A(n49725), .B(n49667), .Z(n49659) );
  XNOR U49728 ( .A(n49655), .B(n49654), .Z(n49667) );
  XNOR U49729 ( .A(n49726), .B(n49651), .Z(n49654) );
  XNOR U49730 ( .A(p_input[1914]), .B(p_input[2074]), .Z(n49651) );
  XOR U49731 ( .A(p_input[1915]), .B(n29415), .Z(n49726) );
  XOR U49732 ( .A(p_input[1916]), .B(p_input[2076]), .Z(n49655) );
  XOR U49733 ( .A(n49665), .B(n49727), .Z(n49725) );
  IV U49734 ( .A(n49656), .Z(n49727) );
  XOR U49735 ( .A(p_input[1905]), .B(p_input[2065]), .Z(n49656) );
  XNOR U49736 ( .A(n49728), .B(n49672), .Z(n49665) );
  XNOR U49737 ( .A(p_input[1919]), .B(n29418), .Z(n49672) );
  XOR U49738 ( .A(n49662), .B(n49671), .Z(n49728) );
  XOR U49739 ( .A(n49729), .B(n49668), .Z(n49671) );
  XOR U49740 ( .A(p_input[1917]), .B(p_input[2077]), .Z(n49668) );
  XOR U49741 ( .A(p_input[1918]), .B(n29420), .Z(n49729) );
  XOR U49742 ( .A(p_input[1913]), .B(p_input[2073]), .Z(n49662) );
  XOR U49743 ( .A(n49684), .B(n49683), .Z(n49649) );
  XNOR U49744 ( .A(n49730), .B(n49691), .Z(n49683) );
  XNOR U49745 ( .A(n49679), .B(n49678), .Z(n49691) );
  XNOR U49746 ( .A(n49731), .B(n49675), .Z(n49678) );
  XNOR U49747 ( .A(p_input[1899]), .B(p_input[2059]), .Z(n49675) );
  XOR U49748 ( .A(p_input[1900]), .B(n28329), .Z(n49731) );
  XOR U49749 ( .A(p_input[1901]), .B(p_input[2061]), .Z(n49679) );
  XOR U49750 ( .A(n49689), .B(n49732), .Z(n49730) );
  IV U49751 ( .A(n49680), .Z(n49732) );
  XOR U49752 ( .A(p_input[1890]), .B(p_input[2050]), .Z(n49680) );
  XNOR U49753 ( .A(n49733), .B(n49696), .Z(n49689) );
  XNOR U49754 ( .A(p_input[1904]), .B(n28332), .Z(n49696) );
  XOR U49755 ( .A(n49686), .B(n49695), .Z(n49733) );
  XOR U49756 ( .A(n49734), .B(n49692), .Z(n49695) );
  XOR U49757 ( .A(p_input[1902]), .B(p_input[2062]), .Z(n49692) );
  XOR U49758 ( .A(p_input[1903]), .B(n28334), .Z(n49734) );
  XOR U49759 ( .A(p_input[1898]), .B(p_input[2058]), .Z(n49686) );
  XOR U49760 ( .A(n49703), .B(n49701), .Z(n49684) );
  XNOR U49761 ( .A(n49735), .B(n49708), .Z(n49701) );
  XOR U49762 ( .A(p_input[1897]), .B(p_input[2057]), .Z(n49708) );
  XOR U49763 ( .A(n49698), .B(n49707), .Z(n49735) );
  XOR U49764 ( .A(n49736), .B(n49704), .Z(n49707) );
  XOR U49765 ( .A(p_input[1895]), .B(p_input[2055]), .Z(n49704) );
  XOR U49766 ( .A(p_input[1896]), .B(n29427), .Z(n49736) );
  XOR U49767 ( .A(p_input[1891]), .B(p_input[2051]), .Z(n49698) );
  XNOR U49768 ( .A(n49713), .B(n49712), .Z(n49703) );
  XOR U49769 ( .A(n49737), .B(n49709), .Z(n49712) );
  XOR U49770 ( .A(p_input[1892]), .B(p_input[2052]), .Z(n49709) );
  XOR U49771 ( .A(p_input[1893]), .B(n29429), .Z(n49737) );
  XOR U49772 ( .A(p_input[1894]), .B(p_input[2054]), .Z(n49713) );
  XNOR U49773 ( .A(n49738), .B(n49739), .Z(n49517) );
  AND U49774 ( .A(n1256), .B(n49740), .Z(n49739) );
  XNOR U49775 ( .A(n49741), .B(n49742), .Z(n1256) );
  NOR U49776 ( .A(n49743), .B(n49744), .Z(n49742) );
  XNOR U49777 ( .A(n49741), .B(n49745), .Z(n49744) );
  NOR U49778 ( .A(n49741), .B(n49526), .Z(n49743) );
  XOR U49779 ( .A(n49746), .B(n49747), .Z(n49741) );
  AND U49780 ( .A(n49748), .B(n49749), .Z(n49747) );
  XOR U49781 ( .A(n49543), .B(n49746), .Z(n49749) );
  XOR U49782 ( .A(n49746), .B(n49544), .Z(n49748) );
  XOR U49783 ( .A(n49750), .B(n49751), .Z(n49746) );
  AND U49784 ( .A(n49752), .B(n49753), .Z(n49751) );
  XOR U49785 ( .A(n49571), .B(n49750), .Z(n49753) );
  XOR U49786 ( .A(n49750), .B(n49572), .Z(n49752) );
  XOR U49787 ( .A(n49754), .B(n49755), .Z(n49750) );
  AND U49788 ( .A(n49756), .B(n49757), .Z(n49755) );
  XOR U49789 ( .A(n49620), .B(n49754), .Z(n49757) );
  XOR U49790 ( .A(n49754), .B(n49621), .Z(n49756) );
  XOR U49791 ( .A(n49758), .B(n49759), .Z(n49754) );
  AND U49792 ( .A(n49760), .B(n49761), .Z(n49759) );
  XOR U49793 ( .A(n49758), .B(n49717), .Z(n49761) );
  XNOR U49794 ( .A(n49762), .B(n49763), .Z(n49470) );
  AND U49795 ( .A(n1260), .B(n49764), .Z(n49763) );
  XNOR U49796 ( .A(n49765), .B(n49766), .Z(n1260) );
  NOR U49797 ( .A(n49767), .B(n49768), .Z(n49766) );
  XOR U49798 ( .A(n49432), .B(n49765), .Z(n49768) );
  NOR U49799 ( .A(n49765), .B(n49431), .Z(n49767) );
  XOR U49800 ( .A(n49769), .B(n49770), .Z(n49765) );
  AND U49801 ( .A(n49771), .B(n49772), .Z(n49770) );
  XNOR U49802 ( .A(n49487), .B(n49769), .Z(n49772) );
  XOR U49803 ( .A(n49769), .B(n49440), .Z(n49771) );
  XOR U49804 ( .A(n49773), .B(n49774), .Z(n49769) );
  AND U49805 ( .A(n49775), .B(n49776), .Z(n49774) );
  XNOR U49806 ( .A(n49497), .B(n49773), .Z(n49776) );
  XOR U49807 ( .A(n49773), .B(n49449), .Z(n49775) );
  XOR U49808 ( .A(n49777), .B(n49778), .Z(n49773) );
  AND U49809 ( .A(n49779), .B(n49780), .Z(n49778) );
  XOR U49810 ( .A(n49777), .B(n49457), .Z(n49779) );
  XOR U49811 ( .A(n49781), .B(n49782), .Z(n49424) );
  AND U49812 ( .A(n1264), .B(n49764), .Z(n49782) );
  XNOR U49813 ( .A(n49762), .B(n49781), .Z(n49764) );
  XNOR U49814 ( .A(n49783), .B(n49784), .Z(n1264) );
  NOR U49815 ( .A(n49785), .B(n49786), .Z(n49784) );
  XNOR U49816 ( .A(n49432), .B(n49787), .Z(n49786) );
  IV U49817 ( .A(n49783), .Z(n49787) );
  AND U49818 ( .A(n49788), .B(n49789), .Z(n49432) );
  NOR U49819 ( .A(n49783), .B(n49431), .Z(n49785) );
  AND U49820 ( .A(n49526), .B(n49525), .Z(n49431) );
  IV U49821 ( .A(n49745), .Z(n49525) );
  XOR U49822 ( .A(n49790), .B(n49791), .Z(n49783) );
  AND U49823 ( .A(n49792), .B(n49793), .Z(n49791) );
  XNOR U49824 ( .A(n49790), .B(n49487), .Z(n49793) );
  XOR U49825 ( .A(n49544), .B(n49794), .Z(n49487) );
  AND U49826 ( .A(n1267), .B(n49795), .Z(n49794) );
  XOR U49827 ( .A(n49540), .B(n49544), .Z(n49795) );
  XNOR U49828 ( .A(n49796), .B(n49790), .Z(n49792) );
  IV U49829 ( .A(n49440), .Z(n49796) );
  XOR U49830 ( .A(n49797), .B(n49798), .Z(n49440) );
  AND U49831 ( .A(n1282), .B(n49799), .Z(n49798) );
  XOR U49832 ( .A(n49800), .B(n49801), .Z(n49790) );
  AND U49833 ( .A(n49802), .B(n49803), .Z(n49801) );
  XNOR U49834 ( .A(n49800), .B(n49497), .Z(n49803) );
  XOR U49835 ( .A(n49572), .B(n49804), .Z(n49497) );
  AND U49836 ( .A(n1267), .B(n49805), .Z(n49804) );
  XOR U49837 ( .A(n49568), .B(n49572), .Z(n49805) );
  XOR U49838 ( .A(n49449), .B(n49800), .Z(n49802) );
  XOR U49839 ( .A(n49806), .B(n49807), .Z(n49449) );
  AND U49840 ( .A(n1282), .B(n49808), .Z(n49807) );
  XOR U49841 ( .A(n49777), .B(n49809), .Z(n49800) );
  AND U49842 ( .A(n49810), .B(n49780), .Z(n49809) );
  XNOR U49843 ( .A(n49507), .B(n49777), .Z(n49780) );
  XOR U49844 ( .A(n49621), .B(n49811), .Z(n49507) );
  AND U49845 ( .A(n1267), .B(n49812), .Z(n49811) );
  XOR U49846 ( .A(n49617), .B(n49621), .Z(n49812) );
  XNOR U49847 ( .A(n49813), .B(n49777), .Z(n49810) );
  IV U49848 ( .A(n49457), .Z(n49813) );
  XOR U49849 ( .A(n49814), .B(n49815), .Z(n49457) );
  AND U49850 ( .A(n1282), .B(n49816), .Z(n49815) );
  XOR U49851 ( .A(n49817), .B(n49818), .Z(n49777) );
  AND U49852 ( .A(n49819), .B(n49820), .Z(n49818) );
  XNOR U49853 ( .A(n49817), .B(n49515), .Z(n49820) );
  XOR U49854 ( .A(n49718), .B(n49821), .Z(n49515) );
  AND U49855 ( .A(n1267), .B(n49822), .Z(n49821) );
  XOR U49856 ( .A(n49714), .B(n49718), .Z(n49822) );
  XNOR U49857 ( .A(n49823), .B(n49817), .Z(n49819) );
  IV U49858 ( .A(n49467), .Z(n49823) );
  XOR U49859 ( .A(n49824), .B(n49825), .Z(n49467) );
  AND U49860 ( .A(n1282), .B(n49826), .Z(n49825) );
  AND U49861 ( .A(n49781), .B(n49762), .Z(n49817) );
  XNOR U49862 ( .A(n49827), .B(n49828), .Z(n49762) );
  AND U49863 ( .A(n1267), .B(n49740), .Z(n49828) );
  XNOR U49864 ( .A(n49738), .B(n49827), .Z(n49740) );
  XNOR U49865 ( .A(n49829), .B(n49830), .Z(n1267) );
  NOR U49866 ( .A(n49831), .B(n49832), .Z(n49830) );
  XNOR U49867 ( .A(n49829), .B(n49745), .Z(n49832) );
  NOR U49868 ( .A(n49788), .B(n49789), .Z(n49745) );
  NOR U49869 ( .A(n49829), .B(n49526), .Z(n49831) );
  AND U49870 ( .A(n49833), .B(n49834), .Z(n49526) );
  IV U49871 ( .A(n49835), .Z(n49833) );
  XOR U49872 ( .A(n49836), .B(n49837), .Z(n49829) );
  AND U49873 ( .A(n49838), .B(n49839), .Z(n49837) );
  XNOR U49874 ( .A(n49836), .B(n49540), .Z(n49839) );
  IV U49875 ( .A(n49543), .Z(n49540) );
  XOR U49876 ( .A(n49840), .B(n49841), .Z(n49543) );
  AND U49877 ( .A(n1271), .B(n49842), .Z(n49841) );
  XOR U49878 ( .A(n49843), .B(n49840), .Z(n49842) );
  XOR U49879 ( .A(n49544), .B(n49836), .Z(n49838) );
  XOR U49880 ( .A(n49844), .B(n49845), .Z(n49544) );
  AND U49881 ( .A(n1278), .B(n49799), .Z(n49845) );
  XOR U49882 ( .A(n49844), .B(n49797), .Z(n49799) );
  XOR U49883 ( .A(n49846), .B(n49847), .Z(n49836) );
  AND U49884 ( .A(n49848), .B(n49849), .Z(n49847) );
  XNOR U49885 ( .A(n49846), .B(n49568), .Z(n49849) );
  IV U49886 ( .A(n49571), .Z(n49568) );
  XOR U49887 ( .A(n49850), .B(n49851), .Z(n49571) );
  AND U49888 ( .A(n1271), .B(n49852), .Z(n49851) );
  XNOR U49889 ( .A(n49853), .B(n49850), .Z(n49852) );
  XOR U49890 ( .A(n49572), .B(n49846), .Z(n49848) );
  XOR U49891 ( .A(n49854), .B(n49855), .Z(n49572) );
  AND U49892 ( .A(n1278), .B(n49808), .Z(n49855) );
  XOR U49893 ( .A(n49854), .B(n49806), .Z(n49808) );
  XOR U49894 ( .A(n49856), .B(n49857), .Z(n49846) );
  AND U49895 ( .A(n49858), .B(n49859), .Z(n49857) );
  XNOR U49896 ( .A(n49856), .B(n49617), .Z(n49859) );
  IV U49897 ( .A(n49620), .Z(n49617) );
  XOR U49898 ( .A(n49860), .B(n49861), .Z(n49620) );
  AND U49899 ( .A(n1271), .B(n49862), .Z(n49861) );
  XOR U49900 ( .A(n49863), .B(n49860), .Z(n49862) );
  XOR U49901 ( .A(n49621), .B(n49856), .Z(n49858) );
  XOR U49902 ( .A(n49864), .B(n49865), .Z(n49621) );
  AND U49903 ( .A(n1278), .B(n49816), .Z(n49865) );
  XOR U49904 ( .A(n49864), .B(n49814), .Z(n49816) );
  XOR U49905 ( .A(n49758), .B(n49866), .Z(n49856) );
  AND U49906 ( .A(n49760), .B(n49867), .Z(n49866) );
  XNOR U49907 ( .A(n49758), .B(n49714), .Z(n49867) );
  IV U49908 ( .A(n49717), .Z(n49714) );
  XOR U49909 ( .A(n49868), .B(n49869), .Z(n49717) );
  AND U49910 ( .A(n1271), .B(n49870), .Z(n49869) );
  XNOR U49911 ( .A(n49871), .B(n49868), .Z(n49870) );
  XOR U49912 ( .A(n49718), .B(n49758), .Z(n49760) );
  XOR U49913 ( .A(n49872), .B(n49873), .Z(n49718) );
  AND U49914 ( .A(n1278), .B(n49826), .Z(n49873) );
  XOR U49915 ( .A(n49872), .B(n49824), .Z(n49826) );
  AND U49916 ( .A(n49827), .B(n49738), .Z(n49758) );
  XNOR U49917 ( .A(n49874), .B(n49875), .Z(n49738) );
  AND U49918 ( .A(n1271), .B(n49876), .Z(n49875) );
  XNOR U49919 ( .A(n49877), .B(n49874), .Z(n49876) );
  XNOR U49920 ( .A(n49878), .B(n49879), .Z(n1271) );
  NOR U49921 ( .A(n49880), .B(n49881), .Z(n49879) );
  XNOR U49922 ( .A(n49878), .B(n49835), .Z(n49881) );
  NOR U49923 ( .A(n49882), .B(n49883), .Z(n49835) );
  NOR U49924 ( .A(n49878), .B(n49834), .Z(n49880) );
  AND U49925 ( .A(n49884), .B(n49885), .Z(n49834) );
  XOR U49926 ( .A(n49886), .B(n49887), .Z(n49878) );
  AND U49927 ( .A(n49888), .B(n49889), .Z(n49887) );
  XNOR U49928 ( .A(n49886), .B(n49884), .Z(n49889) );
  IV U49929 ( .A(n49843), .Z(n49884) );
  XOR U49930 ( .A(n49890), .B(n49891), .Z(n49843) );
  XOR U49931 ( .A(n49892), .B(n49885), .Z(n49891) );
  AND U49932 ( .A(n49853), .B(n49893), .Z(n49885) );
  AND U49933 ( .A(n49894), .B(n49895), .Z(n49892) );
  XOR U49934 ( .A(n49896), .B(n49890), .Z(n49894) );
  XNOR U49935 ( .A(n49840), .B(n49886), .Z(n49888) );
  XNOR U49936 ( .A(n49897), .B(n49898), .Z(n49840) );
  AND U49937 ( .A(n1274), .B(n49899), .Z(n49898) );
  XOR U49938 ( .A(n49900), .B(n49901), .Z(n49886) );
  AND U49939 ( .A(n49902), .B(n49903), .Z(n49901) );
  XNOR U49940 ( .A(n49900), .B(n49853), .Z(n49903) );
  XOR U49941 ( .A(n49904), .B(n49895), .Z(n49853) );
  XNOR U49942 ( .A(n49905), .B(n49890), .Z(n49895) );
  XOR U49943 ( .A(n49906), .B(n49907), .Z(n49890) );
  AND U49944 ( .A(n49908), .B(n49909), .Z(n49907) );
  XOR U49945 ( .A(n49910), .B(n49906), .Z(n49908) );
  XNOR U49946 ( .A(n49911), .B(n49912), .Z(n49905) );
  AND U49947 ( .A(n49913), .B(n49914), .Z(n49912) );
  XOR U49948 ( .A(n49911), .B(n49915), .Z(n49913) );
  XNOR U49949 ( .A(n49896), .B(n49893), .Z(n49904) );
  AND U49950 ( .A(n49916), .B(n49917), .Z(n49893) );
  XOR U49951 ( .A(n49918), .B(n49919), .Z(n49896) );
  AND U49952 ( .A(n49920), .B(n49921), .Z(n49919) );
  XOR U49953 ( .A(n49918), .B(n49922), .Z(n49920) );
  XNOR U49954 ( .A(n49850), .B(n49900), .Z(n49902) );
  XNOR U49955 ( .A(n49923), .B(n49924), .Z(n49850) );
  AND U49956 ( .A(n1274), .B(n49925), .Z(n49924) );
  XOR U49957 ( .A(n49926), .B(n49927), .Z(n49900) );
  AND U49958 ( .A(n49928), .B(n49929), .Z(n49927) );
  XNOR U49959 ( .A(n49926), .B(n49916), .Z(n49929) );
  IV U49960 ( .A(n49863), .Z(n49916) );
  XNOR U49961 ( .A(n49930), .B(n49909), .Z(n49863) );
  XNOR U49962 ( .A(n49931), .B(n49915), .Z(n49909) );
  XOR U49963 ( .A(n49932), .B(n49933), .Z(n49915) );
  AND U49964 ( .A(n49934), .B(n49935), .Z(n49933) );
  XOR U49965 ( .A(n49932), .B(n49936), .Z(n49934) );
  XNOR U49966 ( .A(n49914), .B(n49906), .Z(n49931) );
  XOR U49967 ( .A(n49937), .B(n49938), .Z(n49906) );
  AND U49968 ( .A(n49939), .B(n49940), .Z(n49938) );
  XNOR U49969 ( .A(n49941), .B(n49937), .Z(n49939) );
  XNOR U49970 ( .A(n49942), .B(n49911), .Z(n49914) );
  XOR U49971 ( .A(n49943), .B(n49944), .Z(n49911) );
  AND U49972 ( .A(n49945), .B(n49946), .Z(n49944) );
  XOR U49973 ( .A(n49943), .B(n49947), .Z(n49945) );
  XNOR U49974 ( .A(n49948), .B(n49949), .Z(n49942) );
  AND U49975 ( .A(n49950), .B(n49951), .Z(n49949) );
  XNOR U49976 ( .A(n49948), .B(n49952), .Z(n49950) );
  XNOR U49977 ( .A(n49910), .B(n49917), .Z(n49930) );
  AND U49978 ( .A(n49871), .B(n49953), .Z(n49917) );
  XOR U49979 ( .A(n49922), .B(n49921), .Z(n49910) );
  XNOR U49980 ( .A(n49954), .B(n49918), .Z(n49921) );
  XOR U49981 ( .A(n49955), .B(n49956), .Z(n49918) );
  AND U49982 ( .A(n49957), .B(n49958), .Z(n49956) );
  XOR U49983 ( .A(n49955), .B(n49959), .Z(n49957) );
  XNOR U49984 ( .A(n49960), .B(n49961), .Z(n49954) );
  AND U49985 ( .A(n49962), .B(n49963), .Z(n49961) );
  XOR U49986 ( .A(n49960), .B(n49964), .Z(n49962) );
  XOR U49987 ( .A(n49965), .B(n49966), .Z(n49922) );
  AND U49988 ( .A(n49967), .B(n49968), .Z(n49966) );
  XOR U49989 ( .A(n49965), .B(n49969), .Z(n49967) );
  XNOR U49990 ( .A(n49860), .B(n49926), .Z(n49928) );
  XNOR U49991 ( .A(n49970), .B(n49971), .Z(n49860) );
  AND U49992 ( .A(n1274), .B(n49972), .Z(n49971) );
  XNOR U49993 ( .A(n49973), .B(n49974), .Z(n49972) );
  XOR U49994 ( .A(n49975), .B(n49976), .Z(n49926) );
  AND U49995 ( .A(n49977), .B(n49978), .Z(n49976) );
  XNOR U49996 ( .A(n49975), .B(n49871), .Z(n49978) );
  XOR U49997 ( .A(n49979), .B(n49940), .Z(n49871) );
  XNOR U49998 ( .A(n49980), .B(n49947), .Z(n49940) );
  XOR U49999 ( .A(n49936), .B(n49935), .Z(n49947) );
  XNOR U50000 ( .A(n49981), .B(n49932), .Z(n49935) );
  XOR U50001 ( .A(n49982), .B(n49983), .Z(n49932) );
  AND U50002 ( .A(n49984), .B(n49985), .Z(n49983) );
  XNOR U50003 ( .A(n49986), .B(n49987), .Z(n49984) );
  IV U50004 ( .A(n49982), .Z(n49986) );
  XNOR U50005 ( .A(n49988), .B(n49989), .Z(n49981) );
  NOR U50006 ( .A(n49990), .B(n49991), .Z(n49989) );
  XNOR U50007 ( .A(n49988), .B(n49992), .Z(n49990) );
  XOR U50008 ( .A(n49993), .B(n49994), .Z(n49936) );
  NOR U50009 ( .A(n49995), .B(n49996), .Z(n49994) );
  XNOR U50010 ( .A(n49993), .B(n49997), .Z(n49995) );
  XNOR U50011 ( .A(n49946), .B(n49937), .Z(n49980) );
  XOR U50012 ( .A(n49998), .B(n49999), .Z(n49937) );
  AND U50013 ( .A(n50000), .B(n50001), .Z(n49999) );
  XOR U50014 ( .A(n49998), .B(n50002), .Z(n50000) );
  XOR U50015 ( .A(n50003), .B(n49952), .Z(n49946) );
  XOR U50016 ( .A(n50004), .B(n50005), .Z(n49952) );
  NOR U50017 ( .A(n50006), .B(n50007), .Z(n50005) );
  XOR U50018 ( .A(n50004), .B(n50008), .Z(n50006) );
  XNOR U50019 ( .A(n49951), .B(n49943), .Z(n50003) );
  XOR U50020 ( .A(n50009), .B(n50010), .Z(n49943) );
  AND U50021 ( .A(n50011), .B(n50012), .Z(n50010) );
  XOR U50022 ( .A(n50009), .B(n50013), .Z(n50011) );
  XNOR U50023 ( .A(n50014), .B(n49948), .Z(n49951) );
  XOR U50024 ( .A(n50015), .B(n50016), .Z(n49948) );
  AND U50025 ( .A(n50017), .B(n50018), .Z(n50016) );
  XNOR U50026 ( .A(n50019), .B(n50020), .Z(n50017) );
  IV U50027 ( .A(n50015), .Z(n50019) );
  XNOR U50028 ( .A(n50021), .B(n50022), .Z(n50014) );
  NOR U50029 ( .A(n50023), .B(n50024), .Z(n50022) );
  XNOR U50030 ( .A(n50021), .B(n50025), .Z(n50023) );
  XOR U50031 ( .A(n49941), .B(n49953), .Z(n49979) );
  NOR U50032 ( .A(n49877), .B(n50026), .Z(n49953) );
  XNOR U50033 ( .A(n49959), .B(n49958), .Z(n49941) );
  XNOR U50034 ( .A(n50027), .B(n49964), .Z(n49958) );
  XNOR U50035 ( .A(n50028), .B(n50029), .Z(n49964) );
  NOR U50036 ( .A(n50030), .B(n50031), .Z(n50029) );
  XOR U50037 ( .A(n50028), .B(n50032), .Z(n50030) );
  XNOR U50038 ( .A(n49963), .B(n49955), .Z(n50027) );
  XOR U50039 ( .A(n50033), .B(n50034), .Z(n49955) );
  AND U50040 ( .A(n50035), .B(n50036), .Z(n50034) );
  XOR U50041 ( .A(n50033), .B(n50037), .Z(n50035) );
  XNOR U50042 ( .A(n50038), .B(n49960), .Z(n49963) );
  XOR U50043 ( .A(n50039), .B(n50040), .Z(n49960) );
  AND U50044 ( .A(n50041), .B(n50042), .Z(n50040) );
  XNOR U50045 ( .A(n50043), .B(n50044), .Z(n50041) );
  IV U50046 ( .A(n50039), .Z(n50043) );
  XNOR U50047 ( .A(n50045), .B(n50046), .Z(n50038) );
  NOR U50048 ( .A(n50047), .B(n50048), .Z(n50046) );
  XNOR U50049 ( .A(n50045), .B(n50049), .Z(n50047) );
  XOR U50050 ( .A(n49969), .B(n49968), .Z(n49959) );
  XNOR U50051 ( .A(n50050), .B(n49965), .Z(n49968) );
  XOR U50052 ( .A(n50051), .B(n50052), .Z(n49965) );
  AND U50053 ( .A(n50053), .B(n50054), .Z(n50052) );
  XNOR U50054 ( .A(n50055), .B(n50056), .Z(n50053) );
  IV U50055 ( .A(n50051), .Z(n50055) );
  XNOR U50056 ( .A(n50057), .B(n50058), .Z(n50050) );
  NOR U50057 ( .A(n50059), .B(n50060), .Z(n50058) );
  XNOR U50058 ( .A(n50057), .B(n50061), .Z(n50059) );
  XOR U50059 ( .A(n50062), .B(n50063), .Z(n49969) );
  NOR U50060 ( .A(n50064), .B(n50065), .Z(n50063) );
  XNOR U50061 ( .A(n50062), .B(n50066), .Z(n50064) );
  XNOR U50062 ( .A(n49868), .B(n49975), .Z(n49977) );
  XNOR U50063 ( .A(n50067), .B(n50068), .Z(n49868) );
  AND U50064 ( .A(n1274), .B(n50069), .Z(n50068) );
  AND U50065 ( .A(n49874), .B(n49877), .Z(n49975) );
  XOR U50066 ( .A(n50070), .B(n50026), .Z(n49877) );
  XNOR U50067 ( .A(p_input[1920]), .B(p_input[2048]), .Z(n50026) );
  XNOR U50068 ( .A(n50002), .B(n50001), .Z(n50070) );
  XNOR U50069 ( .A(n50071), .B(n50013), .Z(n50001) );
  XOR U50070 ( .A(n49987), .B(n49985), .Z(n50013) );
  XNOR U50071 ( .A(n50072), .B(n49992), .Z(n49985) );
  XOR U50072 ( .A(p_input[1944]), .B(p_input[2072]), .Z(n49992) );
  XOR U50073 ( .A(n49982), .B(n49991), .Z(n50072) );
  XOR U50074 ( .A(n50073), .B(n49988), .Z(n49991) );
  XOR U50075 ( .A(p_input[1942]), .B(p_input[2070]), .Z(n49988) );
  XOR U50076 ( .A(p_input[1943]), .B(n29410), .Z(n50073) );
  XOR U50077 ( .A(p_input[1938]), .B(p_input[2066]), .Z(n49982) );
  XNOR U50078 ( .A(n49997), .B(n49996), .Z(n49987) );
  XOR U50079 ( .A(n50074), .B(n49993), .Z(n49996) );
  XOR U50080 ( .A(p_input[1939]), .B(p_input[2067]), .Z(n49993) );
  XOR U50081 ( .A(p_input[1940]), .B(n29412), .Z(n50074) );
  XOR U50082 ( .A(p_input[1941]), .B(p_input[2069]), .Z(n49997) );
  XOR U50083 ( .A(n50012), .B(n50075), .Z(n50071) );
  IV U50084 ( .A(n49998), .Z(n50075) );
  XOR U50085 ( .A(p_input[1921]), .B(p_input[2049]), .Z(n49998) );
  XNOR U50086 ( .A(n50076), .B(n50020), .Z(n50012) );
  XNOR U50087 ( .A(n50008), .B(n50007), .Z(n50020) );
  XNOR U50088 ( .A(n50077), .B(n50004), .Z(n50007) );
  XNOR U50089 ( .A(p_input[1946]), .B(p_input[2074]), .Z(n50004) );
  XOR U50090 ( .A(p_input[1947]), .B(n29415), .Z(n50077) );
  XOR U50091 ( .A(p_input[1948]), .B(p_input[2076]), .Z(n50008) );
  XOR U50092 ( .A(n50018), .B(n50078), .Z(n50076) );
  IV U50093 ( .A(n50009), .Z(n50078) );
  XOR U50094 ( .A(p_input[1937]), .B(p_input[2065]), .Z(n50009) );
  XNOR U50095 ( .A(n50079), .B(n50025), .Z(n50018) );
  XNOR U50096 ( .A(p_input[1951]), .B(n29418), .Z(n50025) );
  IV U50097 ( .A(p_input[2079]), .Z(n29418) );
  XOR U50098 ( .A(n50015), .B(n50024), .Z(n50079) );
  XOR U50099 ( .A(n50080), .B(n50021), .Z(n50024) );
  XOR U50100 ( .A(p_input[1949]), .B(p_input[2077]), .Z(n50021) );
  XOR U50101 ( .A(p_input[1950]), .B(n29420), .Z(n50080) );
  XOR U50102 ( .A(p_input[1945]), .B(p_input[2073]), .Z(n50015) );
  XOR U50103 ( .A(n50037), .B(n50036), .Z(n50002) );
  XNOR U50104 ( .A(n50081), .B(n50044), .Z(n50036) );
  XNOR U50105 ( .A(n50032), .B(n50031), .Z(n50044) );
  XNOR U50106 ( .A(n50082), .B(n50028), .Z(n50031) );
  XNOR U50107 ( .A(p_input[1931]), .B(p_input[2059]), .Z(n50028) );
  XOR U50108 ( .A(p_input[1932]), .B(n28329), .Z(n50082) );
  XOR U50109 ( .A(p_input[1933]), .B(p_input[2061]), .Z(n50032) );
  XOR U50110 ( .A(n50042), .B(n50083), .Z(n50081) );
  IV U50111 ( .A(n50033), .Z(n50083) );
  XOR U50112 ( .A(p_input[1922]), .B(p_input[2050]), .Z(n50033) );
  XNOR U50113 ( .A(n50084), .B(n50049), .Z(n50042) );
  XNOR U50114 ( .A(p_input[1936]), .B(n28332), .Z(n50049) );
  IV U50115 ( .A(p_input[2064]), .Z(n28332) );
  XOR U50116 ( .A(n50039), .B(n50048), .Z(n50084) );
  XOR U50117 ( .A(n50085), .B(n50045), .Z(n50048) );
  XOR U50118 ( .A(p_input[1934]), .B(p_input[2062]), .Z(n50045) );
  XOR U50119 ( .A(p_input[1935]), .B(n28334), .Z(n50085) );
  XOR U50120 ( .A(p_input[1930]), .B(p_input[2058]), .Z(n50039) );
  XOR U50121 ( .A(n50056), .B(n50054), .Z(n50037) );
  XNOR U50122 ( .A(n50086), .B(n50061), .Z(n50054) );
  XOR U50123 ( .A(p_input[1929]), .B(p_input[2057]), .Z(n50061) );
  XOR U50124 ( .A(n50051), .B(n50060), .Z(n50086) );
  XOR U50125 ( .A(n50087), .B(n50057), .Z(n50060) );
  XOR U50126 ( .A(p_input[1927]), .B(p_input[2055]), .Z(n50057) );
  XOR U50127 ( .A(p_input[1928]), .B(n29427), .Z(n50087) );
  XOR U50128 ( .A(p_input[1923]), .B(p_input[2051]), .Z(n50051) );
  XNOR U50129 ( .A(n50066), .B(n50065), .Z(n50056) );
  XOR U50130 ( .A(n50088), .B(n50062), .Z(n50065) );
  XOR U50131 ( .A(p_input[1924]), .B(p_input[2052]), .Z(n50062) );
  XOR U50132 ( .A(p_input[1925]), .B(n29429), .Z(n50088) );
  XOR U50133 ( .A(p_input[1926]), .B(p_input[2054]), .Z(n50066) );
  XNOR U50134 ( .A(n50089), .B(n50090), .Z(n49874) );
  AND U50135 ( .A(n1274), .B(n50091), .Z(n50090) );
  XNOR U50136 ( .A(n50092), .B(n50093), .Z(n1274) );
  NOR U50137 ( .A(n50094), .B(n50095), .Z(n50093) );
  XOR U50138 ( .A(n50092), .B(n49882), .Z(n50095) );
  XNOR U50139 ( .A(n50096), .B(n50097), .Z(n49827) );
  AND U50140 ( .A(n1278), .B(n50098), .Z(n50097) );
  XNOR U50141 ( .A(n50099), .B(n50100), .Z(n1278) );
  NOR U50142 ( .A(n50101), .B(n50102), .Z(n50100) );
  XOR U50143 ( .A(n49789), .B(n50099), .Z(n50102) );
  NOR U50144 ( .A(n50099), .B(n49788), .Z(n50101) );
  XOR U50145 ( .A(n50103), .B(n50104), .Z(n50099) );
  AND U50146 ( .A(n50105), .B(n50106), .Z(n50104) );
  XNOR U50147 ( .A(n49844), .B(n50103), .Z(n50106) );
  XOR U50148 ( .A(n50103), .B(n49797), .Z(n50105) );
  XOR U50149 ( .A(n50107), .B(n50108), .Z(n50103) );
  AND U50150 ( .A(n50109), .B(n50110), .Z(n50108) );
  XNOR U50151 ( .A(n49854), .B(n50107), .Z(n50110) );
  XOR U50152 ( .A(n50107), .B(n49806), .Z(n50109) );
  XOR U50153 ( .A(n50111), .B(n50112), .Z(n50107) );
  AND U50154 ( .A(n50113), .B(n50114), .Z(n50112) );
  XOR U50155 ( .A(n50111), .B(n49814), .Z(n50113) );
  XOR U50156 ( .A(n50115), .B(n50116), .Z(n49781) );
  AND U50157 ( .A(n1282), .B(n50098), .Z(n50116) );
  XNOR U50158 ( .A(n50096), .B(n50115), .Z(n50098) );
  XNOR U50159 ( .A(n50117), .B(n50118), .Z(n1282) );
  NOR U50160 ( .A(n50119), .B(n50120), .Z(n50118) );
  XNOR U50161 ( .A(n49789), .B(n50121), .Z(n50120) );
  IV U50162 ( .A(n50117), .Z(n50121) );
  AND U50163 ( .A(n50122), .B(n50123), .Z(n49789) );
  NOR U50164 ( .A(n50117), .B(n49788), .Z(n50119) );
  AND U50165 ( .A(n49882), .B(n49883), .Z(n49788) );
  IV U50166 ( .A(n50124), .Z(n49882) );
  XOR U50167 ( .A(n50125), .B(n50126), .Z(n50117) );
  AND U50168 ( .A(n50127), .B(n50128), .Z(n50126) );
  XNOR U50169 ( .A(n50125), .B(n49844), .Z(n50128) );
  XOR U50170 ( .A(n50129), .B(n50130), .Z(n49844) );
  AND U50171 ( .A(n1285), .B(n49899), .Z(n50130) );
  XOR U50172 ( .A(n49897), .B(n50129), .Z(n49899) );
  XNOR U50173 ( .A(n50131), .B(n50125), .Z(n50127) );
  IV U50174 ( .A(n49797), .Z(n50131) );
  XOR U50175 ( .A(n50132), .B(n50133), .Z(n49797) );
  AND U50176 ( .A(n1290), .B(n50134), .Z(n50133) );
  XOR U50177 ( .A(n50135), .B(n50136), .Z(n50125) );
  AND U50178 ( .A(n50137), .B(n50138), .Z(n50136) );
  XNOR U50179 ( .A(n50135), .B(n49854), .Z(n50138) );
  XOR U50180 ( .A(n50139), .B(n50140), .Z(n49854) );
  AND U50181 ( .A(n1285), .B(n49925), .Z(n50140) );
  XOR U50182 ( .A(n49923), .B(n50139), .Z(n49925) );
  XOR U50183 ( .A(n49806), .B(n50135), .Z(n50137) );
  XOR U50184 ( .A(n50141), .B(n50142), .Z(n49806) );
  AND U50185 ( .A(n1290), .B(n50143), .Z(n50142) );
  XOR U50186 ( .A(n50111), .B(n50144), .Z(n50135) );
  AND U50187 ( .A(n50145), .B(n50114), .Z(n50144) );
  XNOR U50188 ( .A(n49864), .B(n50111), .Z(n50114) );
  XOR U50189 ( .A(n49974), .B(n50146), .Z(n49864) );
  AND U50190 ( .A(n1285), .B(n50147), .Z(n50146) );
  XOR U50191 ( .A(n49970), .B(n49974), .Z(n50147) );
  XNOR U50192 ( .A(n50148), .B(n50111), .Z(n50145) );
  IV U50193 ( .A(n49814), .Z(n50148) );
  XOR U50194 ( .A(n50149), .B(n50150), .Z(n49814) );
  AND U50195 ( .A(n1290), .B(n50151), .Z(n50150) );
  XOR U50196 ( .A(n50152), .B(n50153), .Z(n50111) );
  AND U50197 ( .A(n50154), .B(n50155), .Z(n50153) );
  XNOR U50198 ( .A(n50152), .B(n49872), .Z(n50155) );
  XNOR U50199 ( .A(n50156), .B(n50157), .Z(n49872) );
  AND U50200 ( .A(n1285), .B(n50069), .Z(n50157) );
  XOR U50201 ( .A(n50067), .B(n50158), .Z(n50069) );
  IV U50202 ( .A(n50156), .Z(n50158) );
  XNOR U50203 ( .A(n50159), .B(n50152), .Z(n50154) );
  IV U50204 ( .A(n49824), .Z(n50159) );
  XOR U50205 ( .A(n50160), .B(n50161), .Z(n49824) );
  AND U50206 ( .A(n1290), .B(n50162), .Z(n50161) );
  AND U50207 ( .A(n50115), .B(n50096), .Z(n50152) );
  XNOR U50208 ( .A(n50163), .B(n50164), .Z(n50096) );
  AND U50209 ( .A(n1285), .B(n50091), .Z(n50164) );
  XOR U50210 ( .A(n50165), .B(n50163), .Z(n50091) );
  XNOR U50211 ( .A(n50092), .B(n50166), .Z(n1285) );
  NOR U50212 ( .A(n50094), .B(n50167), .Z(n50166) );
  XNOR U50213 ( .A(n50092), .B(n50124), .Z(n50167) );
  NOR U50214 ( .A(n50122), .B(n50123), .Z(n50124) );
  NOR U50215 ( .A(n50092), .B(n49883), .Z(n50094) );
  AND U50216 ( .A(n49897), .B(n50168), .Z(n49883) );
  XOR U50217 ( .A(n50169), .B(n50170), .Z(n50092) );
  AND U50218 ( .A(n50171), .B(n50172), .Z(n50170) );
  XNOR U50219 ( .A(n49897), .B(n50169), .Z(n50172) );
  XNOR U50220 ( .A(n50173), .B(n50174), .Z(n49897) );
  XOR U50221 ( .A(n50175), .B(n50168), .Z(n50174) );
  AND U50222 ( .A(n49923), .B(n50176), .Z(n50168) );
  AND U50223 ( .A(n50177), .B(n50178), .Z(n50175) );
  XOR U50224 ( .A(n50179), .B(n50173), .Z(n50177) );
  XOR U50225 ( .A(n50169), .B(n50129), .Z(n50171) );
  XOR U50226 ( .A(n50180), .B(n50181), .Z(n50129) );
  AND U50227 ( .A(n1287), .B(n50134), .Z(n50181) );
  XOR U50228 ( .A(n50180), .B(n50132), .Z(n50134) );
  XOR U50229 ( .A(n50182), .B(n50183), .Z(n50169) );
  AND U50230 ( .A(n50184), .B(n50185), .Z(n50183) );
  XNOR U50231 ( .A(n49923), .B(n50182), .Z(n50185) );
  XOR U50232 ( .A(n50186), .B(n50178), .Z(n49923) );
  XNOR U50233 ( .A(n50187), .B(n50173), .Z(n50178) );
  XOR U50234 ( .A(n50188), .B(n50189), .Z(n50173) );
  AND U50235 ( .A(n50190), .B(n50191), .Z(n50189) );
  XOR U50236 ( .A(n50192), .B(n50188), .Z(n50190) );
  XNOR U50237 ( .A(n50193), .B(n50194), .Z(n50187) );
  AND U50238 ( .A(n50195), .B(n50196), .Z(n50194) );
  XOR U50239 ( .A(n50193), .B(n50197), .Z(n50195) );
  XNOR U50240 ( .A(n50179), .B(n50176), .Z(n50186) );
  AND U50241 ( .A(n49970), .B(n50198), .Z(n50176) );
  XOR U50242 ( .A(n50199), .B(n50200), .Z(n50179) );
  AND U50243 ( .A(n50201), .B(n50202), .Z(n50200) );
  XOR U50244 ( .A(n50199), .B(n50203), .Z(n50201) );
  XOR U50245 ( .A(n50182), .B(n50139), .Z(n50184) );
  XOR U50246 ( .A(n50204), .B(n50205), .Z(n50139) );
  AND U50247 ( .A(n1287), .B(n50143), .Z(n50205) );
  XOR U50248 ( .A(n50204), .B(n50141), .Z(n50143) );
  XOR U50249 ( .A(n50206), .B(n50207), .Z(n50182) );
  AND U50250 ( .A(n50208), .B(n50209), .Z(n50207) );
  XNOR U50251 ( .A(n49970), .B(n50206), .Z(n50209) );
  IV U50252 ( .A(n49973), .Z(n49970) );
  XNOR U50253 ( .A(n50210), .B(n50191), .Z(n49973) );
  XNOR U50254 ( .A(n50211), .B(n50197), .Z(n50191) );
  XOR U50255 ( .A(n50212), .B(n50213), .Z(n50197) );
  AND U50256 ( .A(n50214), .B(n50215), .Z(n50213) );
  XOR U50257 ( .A(n50212), .B(n50216), .Z(n50214) );
  XNOR U50258 ( .A(n50196), .B(n50188), .Z(n50211) );
  XOR U50259 ( .A(n50217), .B(n50218), .Z(n50188) );
  AND U50260 ( .A(n50219), .B(n50220), .Z(n50218) );
  XNOR U50261 ( .A(n50221), .B(n50217), .Z(n50219) );
  XNOR U50262 ( .A(n50222), .B(n50193), .Z(n50196) );
  XOR U50263 ( .A(n50223), .B(n50224), .Z(n50193) );
  AND U50264 ( .A(n50225), .B(n50226), .Z(n50224) );
  XOR U50265 ( .A(n50223), .B(n50227), .Z(n50225) );
  XNOR U50266 ( .A(n50228), .B(n50229), .Z(n50222) );
  AND U50267 ( .A(n50230), .B(n50231), .Z(n50229) );
  XNOR U50268 ( .A(n50228), .B(n50232), .Z(n50230) );
  XNOR U50269 ( .A(n50192), .B(n50198), .Z(n50210) );
  AND U50270 ( .A(n50067), .B(n50233), .Z(n50198) );
  XOR U50271 ( .A(n50203), .B(n50202), .Z(n50192) );
  XNOR U50272 ( .A(n50234), .B(n50199), .Z(n50202) );
  XOR U50273 ( .A(n50235), .B(n50236), .Z(n50199) );
  AND U50274 ( .A(n50237), .B(n50238), .Z(n50236) );
  XOR U50275 ( .A(n50235), .B(n50239), .Z(n50237) );
  XNOR U50276 ( .A(n50240), .B(n50241), .Z(n50234) );
  AND U50277 ( .A(n50242), .B(n50243), .Z(n50241) );
  XOR U50278 ( .A(n50240), .B(n50244), .Z(n50242) );
  XOR U50279 ( .A(n50245), .B(n50246), .Z(n50203) );
  AND U50280 ( .A(n50247), .B(n50248), .Z(n50246) );
  XOR U50281 ( .A(n50245), .B(n50249), .Z(n50247) );
  XOR U50282 ( .A(n50206), .B(n49974), .Z(n50208) );
  XOR U50283 ( .A(n50250), .B(n50251), .Z(n49974) );
  AND U50284 ( .A(n1287), .B(n50151), .Z(n50251) );
  XOR U50285 ( .A(n50250), .B(n50149), .Z(n50151) );
  XOR U50286 ( .A(n50252), .B(n50253), .Z(n50206) );
  AND U50287 ( .A(n50254), .B(n50255), .Z(n50253) );
  XNOR U50288 ( .A(n50252), .B(n50067), .Z(n50255) );
  XOR U50289 ( .A(n50256), .B(n50220), .Z(n50067) );
  XNOR U50290 ( .A(n50257), .B(n50227), .Z(n50220) );
  XOR U50291 ( .A(n50216), .B(n50215), .Z(n50227) );
  XNOR U50292 ( .A(n50258), .B(n50212), .Z(n50215) );
  XOR U50293 ( .A(n50259), .B(n50260), .Z(n50212) );
  AND U50294 ( .A(n50261), .B(n50262), .Z(n50260) );
  XOR U50295 ( .A(n50259), .B(n50263), .Z(n50261) );
  XNOR U50296 ( .A(n50264), .B(n50265), .Z(n50258) );
  NOR U50297 ( .A(n50266), .B(n50267), .Z(n50265) );
  XNOR U50298 ( .A(n50264), .B(n50268), .Z(n50266) );
  XOR U50299 ( .A(n50269), .B(n50270), .Z(n50216) );
  NOR U50300 ( .A(n50271), .B(n50272), .Z(n50270) );
  XNOR U50301 ( .A(n50269), .B(n50273), .Z(n50271) );
  XNOR U50302 ( .A(n50226), .B(n50217), .Z(n50257) );
  XOR U50303 ( .A(n50274), .B(n50275), .Z(n50217) );
  NOR U50304 ( .A(n50276), .B(n50277), .Z(n50275) );
  XNOR U50305 ( .A(n50274), .B(n50278), .Z(n50276) );
  XOR U50306 ( .A(n50279), .B(n50232), .Z(n50226) );
  XNOR U50307 ( .A(n50280), .B(n50281), .Z(n50232) );
  NOR U50308 ( .A(n50282), .B(n50283), .Z(n50281) );
  XNOR U50309 ( .A(n50280), .B(n50284), .Z(n50282) );
  XNOR U50310 ( .A(n50231), .B(n50223), .Z(n50279) );
  XOR U50311 ( .A(n50285), .B(n50286), .Z(n50223) );
  AND U50312 ( .A(n50287), .B(n50288), .Z(n50286) );
  XOR U50313 ( .A(n50285), .B(n50289), .Z(n50287) );
  XNOR U50314 ( .A(n50290), .B(n50228), .Z(n50231) );
  XOR U50315 ( .A(n50291), .B(n50292), .Z(n50228) );
  AND U50316 ( .A(n50293), .B(n50294), .Z(n50292) );
  XOR U50317 ( .A(n50291), .B(n50295), .Z(n50293) );
  XNOR U50318 ( .A(n50296), .B(n50297), .Z(n50290) );
  NOR U50319 ( .A(n50298), .B(n50299), .Z(n50297) );
  XOR U50320 ( .A(n50296), .B(n50300), .Z(n50298) );
  XOR U50321 ( .A(n50221), .B(n50233), .Z(n50256) );
  AND U50322 ( .A(n50165), .B(n50301), .Z(n50233) );
  IV U50323 ( .A(n50089), .Z(n50165) );
  XNOR U50324 ( .A(n50239), .B(n50238), .Z(n50221) );
  XNOR U50325 ( .A(n50302), .B(n50244), .Z(n50238) );
  XOR U50326 ( .A(n50303), .B(n50304), .Z(n50244) );
  NOR U50327 ( .A(n50305), .B(n50306), .Z(n50304) );
  XNOR U50328 ( .A(n50303), .B(n50307), .Z(n50305) );
  XNOR U50329 ( .A(n50243), .B(n50235), .Z(n50302) );
  XOR U50330 ( .A(n50308), .B(n50309), .Z(n50235) );
  AND U50331 ( .A(n50310), .B(n50311), .Z(n50309) );
  XNOR U50332 ( .A(n50308), .B(n50312), .Z(n50310) );
  XNOR U50333 ( .A(n50313), .B(n50240), .Z(n50243) );
  XOR U50334 ( .A(n50314), .B(n50315), .Z(n50240) );
  AND U50335 ( .A(n50316), .B(n50317), .Z(n50315) );
  XOR U50336 ( .A(n50314), .B(n50318), .Z(n50316) );
  XNOR U50337 ( .A(n50319), .B(n50320), .Z(n50313) );
  NOR U50338 ( .A(n50321), .B(n50322), .Z(n50320) );
  XOR U50339 ( .A(n50319), .B(n50323), .Z(n50321) );
  XOR U50340 ( .A(n50249), .B(n50248), .Z(n50239) );
  XNOR U50341 ( .A(n50324), .B(n50245), .Z(n50248) );
  XOR U50342 ( .A(n50325), .B(n50326), .Z(n50245) );
  AND U50343 ( .A(n50327), .B(n50328), .Z(n50326) );
  XOR U50344 ( .A(n50325), .B(n50329), .Z(n50327) );
  XNOR U50345 ( .A(n50330), .B(n50331), .Z(n50324) );
  NOR U50346 ( .A(n50332), .B(n50333), .Z(n50331) );
  XNOR U50347 ( .A(n50330), .B(n50334), .Z(n50332) );
  XOR U50348 ( .A(n50335), .B(n50336), .Z(n50249) );
  NOR U50349 ( .A(n50337), .B(n50338), .Z(n50336) );
  XNOR U50350 ( .A(n50335), .B(n50339), .Z(n50337) );
  XNOR U50351 ( .A(n50156), .B(n50252), .Z(n50254) );
  XNOR U50352 ( .A(n50340), .B(n50341), .Z(n50156) );
  AND U50353 ( .A(n1287), .B(n50162), .Z(n50341) );
  XOR U50354 ( .A(n50340), .B(n50160), .Z(n50162) );
  AND U50355 ( .A(n50163), .B(n50089), .Z(n50252) );
  XNOR U50356 ( .A(n50342), .B(n50301), .Z(n50089) );
  XOR U50357 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(
        p_input[2048]), .Z(n50301) );
  XOR U50358 ( .A(n50278), .B(n50277), .Z(n50342) );
  XOR U50359 ( .A(n50343), .B(n50289), .Z(n50277) );
  XOR U50360 ( .A(n50263), .B(n50262), .Z(n50289) );
  XNOR U50361 ( .A(n50344), .B(n50268), .Z(n50262) );
  XOR U50362 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][24] ), .B(
        p_input[2072]), .Z(n50268) );
  XOR U50363 ( .A(n50259), .B(n50267), .Z(n50344) );
  XOR U50364 ( .A(n50345), .B(n50264), .Z(n50267) );
  XOR U50365 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][22] ), .B(
        p_input[2070]), .Z(n50264) );
  XOR U50366 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][23] ), .B(n29410), 
        .Z(n50345) );
  XNOR U50367 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][18] ), .B(n28684), 
        .Z(n50259) );
  XNOR U50368 ( .A(n50273), .B(n50272), .Z(n50263) );
  XOR U50369 ( .A(n50346), .B(n50269), .Z(n50272) );
  XOR U50370 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][19] ), .B(
        p_input[2067]), .Z(n50269) );
  XOR U50371 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][20] ), .B(n29412), 
        .Z(n50346) );
  XOR U50372 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][21] ), .B(
        p_input[2069]), .Z(n50273) );
  XNOR U50373 ( .A(n50288), .B(n50274), .Z(n50343) );
  XNOR U50374 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n28686), 
        .Z(n50274) );
  XNOR U50375 ( .A(n50347), .B(n50295), .Z(n50288) );
  XNOR U50376 ( .A(n50284), .B(n50283), .Z(n50295) );
  XOR U50377 ( .A(n50348), .B(n50280), .Z(n50283) );
  XNOR U50378 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][26] ), .B(n28322), 
        .Z(n50280) );
  XOR U50379 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][27] ), .B(n29415), 
        .Z(n50348) );
  XOR U50380 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][28] ), .B(
        p_input[2076]), .Z(n50284) );
  XNOR U50381 ( .A(n50294), .B(n50285), .Z(n50347) );
  XNOR U50382 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][17] ), .B(n28689), 
        .Z(n50285) );
  XOR U50383 ( .A(n50349), .B(n50300), .Z(n50294) );
  XNOR U50384 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][31] ), .B(
        p_input[2079]), .Z(n50300) );
  XOR U50385 ( .A(n50291), .B(n50299), .Z(n50349) );
  XOR U50386 ( .A(n50350), .B(n50296), .Z(n50299) );
  XOR U50387 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][29] ), .B(
        p_input[2077]), .Z(n50296) );
  XOR U50388 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][30] ), .B(n29420), 
        .Z(n50350) );
  XNOR U50389 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][25] ), .B(n28326), 
        .Z(n50291) );
  XNOR U50390 ( .A(n50312), .B(n50311), .Z(n50278) );
  XNOR U50391 ( .A(n50351), .B(n50318), .Z(n50311) );
  XNOR U50392 ( .A(n50307), .B(n50306), .Z(n50318) );
  XOR U50393 ( .A(n50352), .B(n50303), .Z(n50306) );
  XNOR U50394 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n28694), 
        .Z(n50303) );
  XOR U50395 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n28329), 
        .Z(n50352) );
  XOR U50396 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(
        p_input[2061]), .Z(n50307) );
  XNOR U50397 ( .A(n50317), .B(n50308), .Z(n50351) );
  XNOR U50398 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n28330), 
        .Z(n50308) );
  XOR U50399 ( .A(n50353), .B(n50323), .Z(n50317) );
  XNOR U50400 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][16] ), .B(
        p_input[2064]), .Z(n50323) );
  XOR U50401 ( .A(n50314), .B(n50322), .Z(n50353) );
  XOR U50402 ( .A(n50354), .B(n50319), .Z(n50322) );
  XOR U50403 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(
        p_input[2062]), .Z(n50319) );
  XOR U50404 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n28334), 
        .Z(n50354) );
  XNOR U50405 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n28697), 
        .Z(n50314) );
  XNOR U50406 ( .A(n50329), .B(n50328), .Z(n50312) );
  XNOR U50407 ( .A(n50355), .B(n50334), .Z(n50328) );
  XOR U50408 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(
        p_input[2057]), .Z(n50334) );
  XOR U50409 ( .A(n50325), .B(n50333), .Z(n50355) );
  XOR U50410 ( .A(n50356), .B(n50330), .Z(n50333) );
  XOR U50411 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(
        p_input[2055]), .Z(n50330) );
  XOR U50412 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n29427), 
        .Z(n50356) );
  XNOR U50413 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(n28337), 
        .Z(n50325) );
  XNOR U50414 ( .A(n50339), .B(n50338), .Z(n50329) );
  XOR U50415 ( .A(n50357), .B(n50335), .Z(n50338) );
  XOR U50416 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(
        p_input[2052]), .Z(n50335) );
  XOR U50417 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n29429), 
        .Z(n50357) );
  XOR U50418 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(
        p_input[2054]), .Z(n50339) );
  XNOR U50419 ( .A(n50358), .B(n50359), .Z(n50163) );
  AND U50420 ( .A(n1287), .B(n50360), .Z(n50359) );
  XNOR U50421 ( .A(n50361), .B(n50362), .Z(n1287) );
  NOR U50422 ( .A(n50363), .B(n50364), .Z(n50362) );
  XOR U50423 ( .A(n50123), .B(n50361), .Z(n50364) );
  NOR U50424 ( .A(n50361), .B(n50122), .Z(n50363) );
  XOR U50425 ( .A(n50365), .B(n50366), .Z(n50361) );
  AND U50426 ( .A(n50367), .B(n50368), .Z(n50366) );
  XNOR U50427 ( .A(n50180), .B(n50365), .Z(n50368) );
  XOR U50428 ( .A(n50365), .B(n50132), .Z(n50367) );
  XOR U50429 ( .A(n50369), .B(n50370), .Z(n50365) );
  AND U50430 ( .A(n50371), .B(n50372), .Z(n50370) );
  XNOR U50431 ( .A(n50204), .B(n50369), .Z(n50372) );
  XOR U50432 ( .A(n50369), .B(n50141), .Z(n50371) );
  XOR U50433 ( .A(n50373), .B(n50374), .Z(n50369) );
  AND U50434 ( .A(n50375), .B(n50376), .Z(n50374) );
  XOR U50435 ( .A(n50373), .B(n50149), .Z(n50375) );
  XOR U50436 ( .A(n50377), .B(n50378), .Z(n50115) );
  AND U50437 ( .A(n1290), .B(n50360), .Z(n50378) );
  XOR U50438 ( .A(n50379), .B(n50377), .Z(n50360) );
  XNOR U50439 ( .A(n50380), .B(n50381), .Z(n1290) );
  NOR U50440 ( .A(n50382), .B(n50383), .Z(n50381) );
  XNOR U50441 ( .A(n50123), .B(n50384), .Z(n50383) );
  IV U50442 ( .A(n50380), .Z(n50384) );
  AND U50443 ( .A(n50132), .B(n50385), .Z(n50123) );
  NOR U50444 ( .A(n50380), .B(n50122), .Z(n50382) );
  AND U50445 ( .A(n50180), .B(n50386), .Z(n50122) );
  XOR U50446 ( .A(n50387), .B(n50388), .Z(n50380) );
  AND U50447 ( .A(n50389), .B(n50390), .Z(n50388) );
  XNOR U50448 ( .A(n50387), .B(n50180), .Z(n50390) );
  XNOR U50449 ( .A(n50391), .B(n50392), .Z(n50180) );
  XOR U50450 ( .A(n50393), .B(n50386), .Z(n50392) );
  AND U50451 ( .A(n50204), .B(n50394), .Z(n50386) );
  AND U50452 ( .A(n50395), .B(n50396), .Z(n50393) );
  XOR U50453 ( .A(n50397), .B(n50391), .Z(n50395) );
  XNOR U50454 ( .A(n50398), .B(n50387), .Z(n50389) );
  IV U50455 ( .A(n50132), .Z(n50398) );
  XNOR U50456 ( .A(n50399), .B(n50400), .Z(n50132) );
  XOR U50457 ( .A(n50401), .B(n50385), .Z(n50400) );
  AND U50458 ( .A(n50141), .B(n50402), .Z(n50385) );
  AND U50459 ( .A(n50403), .B(n50404), .Z(n50401) );
  XNOR U50460 ( .A(n50399), .B(n50405), .Z(n50403) );
  XOR U50461 ( .A(n50406), .B(n50407), .Z(n50387) );
  AND U50462 ( .A(n50408), .B(n50409), .Z(n50407) );
  XNOR U50463 ( .A(n50406), .B(n50204), .Z(n50409) );
  XOR U50464 ( .A(n50410), .B(n50396), .Z(n50204) );
  XNOR U50465 ( .A(n50411), .B(n50391), .Z(n50396) );
  XOR U50466 ( .A(n50412), .B(n50413), .Z(n50391) );
  AND U50467 ( .A(n50414), .B(n50415), .Z(n50413) );
  XOR U50468 ( .A(n50416), .B(n50412), .Z(n50414) );
  XNOR U50469 ( .A(n50417), .B(n50418), .Z(n50411) );
  AND U50470 ( .A(n50419), .B(n50420), .Z(n50418) );
  XOR U50471 ( .A(n50417), .B(n50421), .Z(n50419) );
  XNOR U50472 ( .A(n50397), .B(n50394), .Z(n50410) );
  AND U50473 ( .A(n50250), .B(n50422), .Z(n50394) );
  XOR U50474 ( .A(n50423), .B(n50424), .Z(n50397) );
  AND U50475 ( .A(n50425), .B(n50426), .Z(n50424) );
  XOR U50476 ( .A(n50423), .B(n50427), .Z(n50425) );
  XOR U50477 ( .A(n50141), .B(n50406), .Z(n50408) );
  XNOR U50478 ( .A(n50428), .B(n50405), .Z(n50141) );
  XNOR U50479 ( .A(n50429), .B(n50430), .Z(n50405) );
  AND U50480 ( .A(n50431), .B(n50432), .Z(n50430) );
  XOR U50481 ( .A(n50429), .B(n50433), .Z(n50431) );
  XNOR U50482 ( .A(n50404), .B(n50402), .Z(n50428) );
  AND U50483 ( .A(n50149), .B(n50434), .Z(n50402) );
  XNOR U50484 ( .A(n50435), .B(n50399), .Z(n50404) );
  XOR U50485 ( .A(n50436), .B(n50437), .Z(n50399) );
  AND U50486 ( .A(n50438), .B(n50439), .Z(n50437) );
  XOR U50487 ( .A(n50436), .B(n50440), .Z(n50438) );
  XNOR U50488 ( .A(n50441), .B(n50442), .Z(n50435) );
  AND U50489 ( .A(n50443), .B(n50444), .Z(n50442) );
  XNOR U50490 ( .A(n50441), .B(n50445), .Z(n50443) );
  XOR U50491 ( .A(n50373), .B(n50446), .Z(n50406) );
  AND U50492 ( .A(n50447), .B(n50376), .Z(n50446) );
  XNOR U50493 ( .A(n50250), .B(n50373), .Z(n50376) );
  XOR U50494 ( .A(n50448), .B(n50415), .Z(n50250) );
  XNOR U50495 ( .A(n50449), .B(n50421), .Z(n50415) );
  XOR U50496 ( .A(n50450), .B(n50451), .Z(n50421) );
  AND U50497 ( .A(n50452), .B(n50453), .Z(n50451) );
  XOR U50498 ( .A(n50450), .B(n50454), .Z(n50452) );
  XNOR U50499 ( .A(n50420), .B(n50412), .Z(n50449) );
  XOR U50500 ( .A(n50455), .B(n50456), .Z(n50412) );
  AND U50501 ( .A(n50457), .B(n50458), .Z(n50456) );
  XNOR U50502 ( .A(n50459), .B(n50455), .Z(n50457) );
  XNOR U50503 ( .A(n50460), .B(n50417), .Z(n50420) );
  XOR U50504 ( .A(n50461), .B(n50462), .Z(n50417) );
  AND U50505 ( .A(n50463), .B(n50464), .Z(n50462) );
  XOR U50506 ( .A(n50461), .B(n50465), .Z(n50463) );
  XNOR U50507 ( .A(n50466), .B(n50467), .Z(n50460) );
  AND U50508 ( .A(n50468), .B(n50469), .Z(n50467) );
  XNOR U50509 ( .A(n50466), .B(n50470), .Z(n50468) );
  XNOR U50510 ( .A(n50416), .B(n50422), .Z(n50448) );
  AND U50511 ( .A(n50340), .B(n50471), .Z(n50422) );
  XOR U50512 ( .A(n50427), .B(n50426), .Z(n50416) );
  XNOR U50513 ( .A(n50472), .B(n50423), .Z(n50426) );
  XOR U50514 ( .A(n50473), .B(n50474), .Z(n50423) );
  AND U50515 ( .A(n50475), .B(n50476), .Z(n50474) );
  XOR U50516 ( .A(n50473), .B(n50477), .Z(n50475) );
  XNOR U50517 ( .A(n50478), .B(n50479), .Z(n50472) );
  AND U50518 ( .A(n50480), .B(n50481), .Z(n50479) );
  XOR U50519 ( .A(n50478), .B(n50482), .Z(n50480) );
  XOR U50520 ( .A(n50483), .B(n50484), .Z(n50427) );
  AND U50521 ( .A(n50485), .B(n50486), .Z(n50484) );
  XOR U50522 ( .A(n50483), .B(n50487), .Z(n50485) );
  XNOR U50523 ( .A(n50488), .B(n50373), .Z(n50447) );
  IV U50524 ( .A(n50149), .Z(n50488) );
  XOR U50525 ( .A(n50489), .B(n50440), .Z(n50149) );
  XOR U50526 ( .A(n50433), .B(n50432), .Z(n50440) );
  XNOR U50527 ( .A(n50490), .B(n50429), .Z(n50432) );
  XOR U50528 ( .A(n50491), .B(n50492), .Z(n50429) );
  AND U50529 ( .A(n50493), .B(n50494), .Z(n50492) );
  XOR U50530 ( .A(n50491), .B(n50495), .Z(n50493) );
  XNOR U50531 ( .A(n50496), .B(n50497), .Z(n50490) );
  AND U50532 ( .A(n50498), .B(n50499), .Z(n50497) );
  XOR U50533 ( .A(n50496), .B(n50500), .Z(n50498) );
  XOR U50534 ( .A(n50501), .B(n50502), .Z(n50433) );
  AND U50535 ( .A(n50503), .B(n50504), .Z(n50502) );
  XOR U50536 ( .A(n50501), .B(n50505), .Z(n50503) );
  XNOR U50537 ( .A(n50439), .B(n50434), .Z(n50489) );
  AND U50538 ( .A(n50160), .B(n50506), .Z(n50434) );
  XOR U50539 ( .A(n50507), .B(n50445), .Z(n50439) );
  XNOR U50540 ( .A(n50508), .B(n50509), .Z(n50445) );
  AND U50541 ( .A(n50510), .B(n50511), .Z(n50509) );
  XOR U50542 ( .A(n50508), .B(n50512), .Z(n50510) );
  XNOR U50543 ( .A(n50444), .B(n50436), .Z(n50507) );
  XOR U50544 ( .A(n50513), .B(n50514), .Z(n50436) );
  AND U50545 ( .A(n50515), .B(n50516), .Z(n50514) );
  XOR U50546 ( .A(n50513), .B(n50517), .Z(n50515) );
  XNOR U50547 ( .A(n50518), .B(n50441), .Z(n50444) );
  XOR U50548 ( .A(n50519), .B(n50520), .Z(n50441) );
  AND U50549 ( .A(n50521), .B(n50522), .Z(n50520) );
  XOR U50550 ( .A(n50519), .B(n50523), .Z(n50521) );
  XNOR U50551 ( .A(n50524), .B(n50525), .Z(n50518) );
  AND U50552 ( .A(n50526), .B(n50527), .Z(n50525) );
  XNOR U50553 ( .A(n50524), .B(n50528), .Z(n50526) );
  XOR U50554 ( .A(n50529), .B(n50530), .Z(n50373) );
  AND U50555 ( .A(n50531), .B(n50532), .Z(n50530) );
  XNOR U50556 ( .A(n50529), .B(n50340), .Z(n50532) );
  XOR U50557 ( .A(n50533), .B(n50458), .Z(n50340) );
  XNOR U50558 ( .A(n50534), .B(n50465), .Z(n50458) );
  XOR U50559 ( .A(n50454), .B(n50453), .Z(n50465) );
  XNOR U50560 ( .A(n50535), .B(n50450), .Z(n50453) );
  XOR U50561 ( .A(n50536), .B(n50537), .Z(n50450) );
  AND U50562 ( .A(n50538), .B(n50539), .Z(n50537) );
  XOR U50563 ( .A(n50536), .B(n50540), .Z(n50538) );
  XNOR U50564 ( .A(n50541), .B(n50542), .Z(n50535) );
  NOR U50565 ( .A(n50543), .B(n50544), .Z(n50542) );
  XNOR U50566 ( .A(n50541), .B(n50545), .Z(n50543) );
  XOR U50567 ( .A(n50546), .B(n50547), .Z(n50454) );
  NOR U50568 ( .A(n50548), .B(n50549), .Z(n50547) );
  XNOR U50569 ( .A(n50546), .B(n50550), .Z(n50548) );
  XNOR U50570 ( .A(n50464), .B(n50455), .Z(n50534) );
  XOR U50571 ( .A(n50551), .B(n50552), .Z(n50455) );
  NOR U50572 ( .A(n50553), .B(n50554), .Z(n50552) );
  XNOR U50573 ( .A(n50551), .B(n50555), .Z(n50553) );
  XOR U50574 ( .A(n50556), .B(n50470), .Z(n50464) );
  XNOR U50575 ( .A(n50557), .B(n50558), .Z(n50470) );
  NOR U50576 ( .A(n50559), .B(n50560), .Z(n50558) );
  XNOR U50577 ( .A(n50557), .B(n50561), .Z(n50559) );
  XNOR U50578 ( .A(n50469), .B(n50461), .Z(n50556) );
  XOR U50579 ( .A(n50562), .B(n50563), .Z(n50461) );
  AND U50580 ( .A(n50564), .B(n50565), .Z(n50563) );
  XOR U50581 ( .A(n50562), .B(n50566), .Z(n50564) );
  XNOR U50582 ( .A(n50567), .B(n50466), .Z(n50469) );
  XOR U50583 ( .A(n50568), .B(n50569), .Z(n50466) );
  AND U50584 ( .A(n50570), .B(n50571), .Z(n50569) );
  XOR U50585 ( .A(n50568), .B(n50572), .Z(n50570) );
  XNOR U50586 ( .A(n50573), .B(n50574), .Z(n50567) );
  NOR U50587 ( .A(n50575), .B(n50576), .Z(n50574) );
  XOR U50588 ( .A(n50573), .B(n50577), .Z(n50575) );
  XOR U50589 ( .A(n50459), .B(n50471), .Z(n50533) );
  AND U50590 ( .A(n50379), .B(n50578), .Z(n50471) );
  IV U50591 ( .A(n50358), .Z(n50379) );
  XNOR U50592 ( .A(n50477), .B(n50476), .Z(n50459) );
  XNOR U50593 ( .A(n50579), .B(n50482), .Z(n50476) );
  XOR U50594 ( .A(n50580), .B(n50581), .Z(n50482) );
  NOR U50595 ( .A(n50582), .B(n50583), .Z(n50581) );
  XNOR U50596 ( .A(n50580), .B(n50584), .Z(n50582) );
  XNOR U50597 ( .A(n50481), .B(n50473), .Z(n50579) );
  XOR U50598 ( .A(n50585), .B(n50586), .Z(n50473) );
  AND U50599 ( .A(n50587), .B(n50588), .Z(n50586) );
  XNOR U50600 ( .A(n50585), .B(n50589), .Z(n50587) );
  XNOR U50601 ( .A(n50590), .B(n50478), .Z(n50481) );
  XOR U50602 ( .A(n50591), .B(n50592), .Z(n50478) );
  AND U50603 ( .A(n50593), .B(n50594), .Z(n50592) );
  XOR U50604 ( .A(n50591), .B(n50595), .Z(n50593) );
  XNOR U50605 ( .A(n50596), .B(n50597), .Z(n50590) );
  NOR U50606 ( .A(n50598), .B(n50599), .Z(n50597) );
  XOR U50607 ( .A(n50596), .B(n50600), .Z(n50598) );
  XOR U50608 ( .A(n50487), .B(n50486), .Z(n50477) );
  XNOR U50609 ( .A(n50601), .B(n50483), .Z(n50486) );
  XOR U50610 ( .A(n50602), .B(n50603), .Z(n50483) );
  AND U50611 ( .A(n50604), .B(n50605), .Z(n50603) );
  XOR U50612 ( .A(n50602), .B(n50606), .Z(n50604) );
  XNOR U50613 ( .A(n50607), .B(n50608), .Z(n50601) );
  NOR U50614 ( .A(n50609), .B(n50610), .Z(n50608) );
  XNOR U50615 ( .A(n50607), .B(n50611), .Z(n50609) );
  XOR U50616 ( .A(n50612), .B(n50613), .Z(n50487) );
  NOR U50617 ( .A(n50614), .B(n50615), .Z(n50613) );
  XNOR U50618 ( .A(n50612), .B(n50616), .Z(n50614) );
  XNOR U50619 ( .A(n50617), .B(n50529), .Z(n50531) );
  IV U50620 ( .A(n50160), .Z(n50617) );
  XOR U50621 ( .A(n50618), .B(n50517), .Z(n50160) );
  XOR U50622 ( .A(n50495), .B(n50494), .Z(n50517) );
  XNOR U50623 ( .A(n50619), .B(n50500), .Z(n50494) );
  XOR U50624 ( .A(n50620), .B(n50621), .Z(n50500) );
  NOR U50625 ( .A(n50622), .B(n50623), .Z(n50621) );
  XNOR U50626 ( .A(n50620), .B(n50624), .Z(n50622) );
  XNOR U50627 ( .A(n50499), .B(n50491), .Z(n50619) );
  XOR U50628 ( .A(n50625), .B(n50626), .Z(n50491) );
  AND U50629 ( .A(n50627), .B(n50628), .Z(n50626) );
  XNOR U50630 ( .A(n50625), .B(n50629), .Z(n50627) );
  XNOR U50631 ( .A(n50630), .B(n50496), .Z(n50499) );
  XOR U50632 ( .A(n50631), .B(n50632), .Z(n50496) );
  AND U50633 ( .A(n50633), .B(n50634), .Z(n50632) );
  XOR U50634 ( .A(n50631), .B(n50635), .Z(n50633) );
  XNOR U50635 ( .A(n50636), .B(n50637), .Z(n50630) );
  NOR U50636 ( .A(n50638), .B(n50639), .Z(n50637) );
  XOR U50637 ( .A(n50636), .B(n50640), .Z(n50638) );
  XOR U50638 ( .A(n50505), .B(n50504), .Z(n50495) );
  XNOR U50639 ( .A(n50641), .B(n50501), .Z(n50504) );
  XOR U50640 ( .A(n50642), .B(n50643), .Z(n50501) );
  AND U50641 ( .A(n50644), .B(n50645), .Z(n50643) );
  XOR U50642 ( .A(n50642), .B(n50646), .Z(n50644) );
  XNOR U50643 ( .A(n50647), .B(n50648), .Z(n50641) );
  NOR U50644 ( .A(n50649), .B(n50650), .Z(n50648) );
  XNOR U50645 ( .A(n50647), .B(n50651), .Z(n50649) );
  XOR U50646 ( .A(n50652), .B(n50653), .Z(n50505) );
  NOR U50647 ( .A(n50654), .B(n50655), .Z(n50653) );
  XNOR U50648 ( .A(n50652), .B(n50656), .Z(n50654) );
  XNOR U50649 ( .A(n50516), .B(n50506), .Z(n50618) );
  AND U50650 ( .A(n50377), .B(n50657), .Z(n50506) );
  XNOR U50651 ( .A(n50658), .B(n50523), .Z(n50516) );
  XOR U50652 ( .A(n50512), .B(n50511), .Z(n50523) );
  XNOR U50653 ( .A(n50659), .B(n50508), .Z(n50511) );
  XOR U50654 ( .A(n50660), .B(n50661), .Z(n50508) );
  AND U50655 ( .A(n50662), .B(n50663), .Z(n50661) );
  XOR U50656 ( .A(n50660), .B(n50664), .Z(n50662) );
  XNOR U50657 ( .A(n50665), .B(n50666), .Z(n50659) );
  NOR U50658 ( .A(n50667), .B(n50668), .Z(n50666) );
  XNOR U50659 ( .A(n50665), .B(n50669), .Z(n50667) );
  XOR U50660 ( .A(n50670), .B(n50671), .Z(n50512) );
  NOR U50661 ( .A(n50672), .B(n50673), .Z(n50671) );
  XNOR U50662 ( .A(n50670), .B(n50674), .Z(n50672) );
  XNOR U50663 ( .A(n50522), .B(n50513), .Z(n50658) );
  XOR U50664 ( .A(n50675), .B(n50676), .Z(n50513) );
  NOR U50665 ( .A(n50677), .B(n50678), .Z(n50676) );
  XNOR U50666 ( .A(n50675), .B(n50679), .Z(n50677) );
  XOR U50667 ( .A(n50680), .B(n50528), .Z(n50522) );
  XNOR U50668 ( .A(n50681), .B(n50682), .Z(n50528) );
  NOR U50669 ( .A(n50683), .B(n50684), .Z(n50682) );
  XNOR U50670 ( .A(n50681), .B(n50685), .Z(n50683) );
  XNOR U50671 ( .A(n50527), .B(n50519), .Z(n50680) );
  XOR U50672 ( .A(n50686), .B(n50687), .Z(n50519) );
  AND U50673 ( .A(n50688), .B(n50689), .Z(n50687) );
  XOR U50674 ( .A(n50686), .B(n50690), .Z(n50688) );
  XNOR U50675 ( .A(n50691), .B(n50524), .Z(n50527) );
  XOR U50676 ( .A(n50692), .B(n50693), .Z(n50524) );
  AND U50677 ( .A(n50694), .B(n50695), .Z(n50693) );
  XOR U50678 ( .A(n50692), .B(n50696), .Z(n50694) );
  XNOR U50679 ( .A(n50697), .B(n50698), .Z(n50691) );
  NOR U50680 ( .A(n50699), .B(n50700), .Z(n50698) );
  XOR U50681 ( .A(n50697), .B(n50701), .Z(n50699) );
  AND U50682 ( .A(n50377), .B(n50358), .Z(n50529) );
  XNOR U50683 ( .A(n50702), .B(n50578), .Z(n50358) );
  XOR U50684 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(
        p_input[2048]), .Z(n50578) );
  XOR U50685 ( .A(n50555), .B(n50554), .Z(n50702) );
  XOR U50686 ( .A(n50703), .B(n50566), .Z(n50554) );
  XOR U50687 ( .A(n50540), .B(n50539), .Z(n50566) );
  XNOR U50688 ( .A(n50704), .B(n50545), .Z(n50539) );
  XOR U50689 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .B(
        p_input[2072]), .Z(n50545) );
  XOR U50690 ( .A(n50536), .B(n50544), .Z(n50704) );
  XOR U50691 ( .A(n50705), .B(n50541), .Z(n50544) );
  XOR U50692 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .B(
        p_input[2070]), .Z(n50541) );
  XOR U50693 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .B(n29410), 
        .Z(n50705) );
  XNOR U50694 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .B(n28684), 
        .Z(n50536) );
  XNOR U50695 ( .A(n50550), .B(n50549), .Z(n50540) );
  XOR U50696 ( .A(n50706), .B(n50546), .Z(n50549) );
  XOR U50697 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .B(
        p_input[2067]), .Z(n50546) );
  XOR U50698 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .B(n29412), 
        .Z(n50706) );
  XOR U50699 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .B(
        p_input[2069]), .Z(n50550) );
  XNOR U50700 ( .A(n50565), .B(n50551), .Z(n50703) );
  XNOR U50701 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(n28686), 
        .Z(n50551) );
  XNOR U50702 ( .A(n50707), .B(n50572), .Z(n50565) );
  XNOR U50703 ( .A(n50561), .B(n50560), .Z(n50572) );
  XOR U50704 ( .A(n50708), .B(n50557), .Z(n50560) );
  XNOR U50705 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .B(n28322), 
        .Z(n50557) );
  XOR U50706 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .B(n29415), 
        .Z(n50708) );
  XOR U50707 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .B(
        p_input[2076]), .Z(n50561) );
  XNOR U50708 ( .A(n50571), .B(n50562), .Z(n50707) );
  XNOR U50709 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .B(n28689), 
        .Z(n50562) );
  XOR U50710 ( .A(n50709), .B(n50577), .Z(n50571) );
  XNOR U50711 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .B(
        p_input[2079]), .Z(n50577) );
  XOR U50712 ( .A(n50568), .B(n50576), .Z(n50709) );
  XOR U50713 ( .A(n50710), .B(n50573), .Z(n50576) );
  XOR U50714 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .B(
        p_input[2077]), .Z(n50573) );
  XOR U50715 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .B(n29420), 
        .Z(n50710) );
  XNOR U50716 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .B(n28326), 
        .Z(n50568) );
  XNOR U50717 ( .A(n50589), .B(n50588), .Z(n50555) );
  XNOR U50718 ( .A(n50711), .B(n50595), .Z(n50588) );
  XNOR U50719 ( .A(n50584), .B(n50583), .Z(n50595) );
  XOR U50720 ( .A(n50712), .B(n50580), .Z(n50583) );
  XNOR U50721 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n28694), 
        .Z(n50580) );
  XOR U50722 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(n28329), 
        .Z(n50712) );
  XOR U50723 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(
        p_input[2061]), .Z(n50584) );
  XNOR U50724 ( .A(n50594), .B(n50585), .Z(n50711) );
  XNOR U50725 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .B(n28330), 
        .Z(n50585) );
  XOR U50726 ( .A(n50713), .B(n50600), .Z(n50594) );
  XNOR U50727 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .B(
        p_input[2064]), .Z(n50600) );
  XOR U50728 ( .A(n50591), .B(n50599), .Z(n50713) );
  XOR U50729 ( .A(n50714), .B(n50596), .Z(n50599) );
  XOR U50730 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(
        p_input[2062]), .Z(n50596) );
  XOR U50731 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(n28334), 
        .Z(n50714) );
  XNOR U50732 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(n28697), 
        .Z(n50591) );
  XNOR U50733 ( .A(n50606), .B(n50605), .Z(n50589) );
  XNOR U50734 ( .A(n50715), .B(n50611), .Z(n50605) );
  XNOR U50735 ( .A(n1292), .B(p_input[2057]), .Z(n50611) );
  IV U50736 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .Z(n1292) );
  XOR U50737 ( .A(n50602), .B(n50610), .Z(n50715) );
  XOR U50738 ( .A(n50716), .B(n50607), .Z(n50610) );
  XNOR U50739 ( .A(n3020), .B(p_input[2055]), .Z(n50607) );
  IV U50740 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .Z(n3020) );
  XOR U50741 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .B(n29427), 
        .Z(n50716) );
  XNOR U50742 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .B(n28337), 
        .Z(n50602) );
  XNOR U50743 ( .A(n50616), .B(n50615), .Z(n50606) );
  XOR U50744 ( .A(n50717), .B(n50612), .Z(n50615) );
  XOR U50745 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(
        p_input[2052]), .Z(n50612) );
  XOR U50746 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(n29429), 
        .Z(n50717) );
  XOR U50747 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .B(
        p_input[2054]), .Z(n50616) );
  XOR U50748 ( .A(n50718), .B(n50679), .Z(n50377) );
  XNOR U50749 ( .A(n50629), .B(n50628), .Z(n50679) );
  XNOR U50750 ( .A(n50719), .B(n50635), .Z(n50628) );
  XNOR U50751 ( .A(n50624), .B(n50623), .Z(n50635) );
  XOR U50752 ( .A(n50720), .B(n50620), .Z(n50623) );
  XNOR U50753 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n28694), .Z(n50620) );
  IV U50754 ( .A(p_input[2059]), .Z(n28694) );
  XOR U50755 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n28329), .Z(n50720) );
  IV U50756 ( .A(p_input[2060]), .Z(n28329) );
  XOR U50757 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[2061]), .Z(
        n50624) );
  XNOR U50758 ( .A(n50634), .B(n50625), .Z(n50719) );
  XNOR U50759 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n28330), .Z(n50625) );
  IV U50760 ( .A(p_input[2050]), .Z(n28330) );
  XOR U50761 ( .A(n50721), .B(n50640), .Z(n50634) );
  XNOR U50762 ( .A(\knn_comb_/min_val_out[0][16] ), .B(p_input[2064]), .Z(
        n50640) );
  XOR U50763 ( .A(n50631), .B(n50639), .Z(n50721) );
  XOR U50764 ( .A(n50722), .B(n50636), .Z(n50639) );
  XOR U50765 ( .A(\knn_comb_/min_val_out[0][14] ), .B(p_input[2062]), .Z(
        n50636) );
  XOR U50766 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n28334), .Z(n50722) );
  IV U50767 ( .A(p_input[2063]), .Z(n28334) );
  XNOR U50768 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n28697), .Z(n50631) );
  IV U50769 ( .A(p_input[2058]), .Z(n28697) );
  XNOR U50770 ( .A(n50646), .B(n50645), .Z(n50629) );
  XNOR U50771 ( .A(n50723), .B(n50651), .Z(n50645) );
  XNOR U50772 ( .A(n1291), .B(p_input[2057]), .Z(n50651) );
  IV U50773 ( .A(\knn_comb_/min_val_out[0][9] ), .Z(n1291) );
  XOR U50774 ( .A(n50642), .B(n50650), .Z(n50723) );
  XOR U50775 ( .A(n50724), .B(n50647), .Z(n50650) );
  XNOR U50776 ( .A(n3019), .B(p_input[2055]), .Z(n50647) );
  IV U50777 ( .A(\knn_comb_/min_val_out[0][7] ), .Z(n3019) );
  XOR U50778 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n29427), .Z(n50724) );
  IV U50779 ( .A(p_input[2056]), .Z(n29427) );
  XNOR U50780 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n28337), .Z(n50642) );
  IV U50781 ( .A(p_input[2051]), .Z(n28337) );
  XNOR U50782 ( .A(n50656), .B(n50655), .Z(n50646) );
  XOR U50783 ( .A(n50725), .B(n50652), .Z(n50655) );
  XOR U50784 ( .A(\knn_comb_/min_val_out[0][4] ), .B(p_input[2052]), .Z(n50652) );
  XOR U50785 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n29429), .Z(n50725) );
  IV U50786 ( .A(p_input[2053]), .Z(n29429) );
  XOR U50787 ( .A(\knn_comb_/min_val_out[0][6] ), .B(p_input[2054]), .Z(n50656) );
  XOR U50788 ( .A(n50678), .B(n50657), .Z(n50718) );
  XOR U50789 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[2048]), .Z(n50657) );
  XOR U50790 ( .A(n50726), .B(n50690), .Z(n50678) );
  XOR U50791 ( .A(n50664), .B(n50663), .Z(n50690) );
  XNOR U50792 ( .A(n50727), .B(n50669), .Z(n50663) );
  XOR U50793 ( .A(\knn_comb_/min_val_out[0][24] ), .B(p_input[2072]), .Z(
        n50669) );
  XOR U50794 ( .A(n50660), .B(n50668), .Z(n50727) );
  XOR U50795 ( .A(n50728), .B(n50665), .Z(n50668) );
  XOR U50796 ( .A(\knn_comb_/min_val_out[0][22] ), .B(p_input[2070]), .Z(
        n50665) );
  XOR U50797 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n29410), .Z(n50728) );
  IV U50798 ( .A(p_input[2071]), .Z(n29410) );
  XNOR U50799 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n28684), .Z(n50660) );
  IV U50800 ( .A(p_input[2066]), .Z(n28684) );
  XNOR U50801 ( .A(n50674), .B(n50673), .Z(n50664) );
  XOR U50802 ( .A(n50729), .B(n50670), .Z(n50673) );
  XOR U50803 ( .A(\knn_comb_/min_val_out[0][19] ), .B(p_input[2067]), .Z(
        n50670) );
  XOR U50804 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n29412), .Z(n50729) );
  IV U50805 ( .A(p_input[2068]), .Z(n29412) );
  XOR U50806 ( .A(\knn_comb_/min_val_out[0][21] ), .B(p_input[2069]), .Z(
        n50674) );
  XNOR U50807 ( .A(n50689), .B(n50675), .Z(n50726) );
  XNOR U50808 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n28686), .Z(n50675) );
  IV U50809 ( .A(p_input[2049]), .Z(n28686) );
  XNOR U50810 ( .A(n50730), .B(n50696), .Z(n50689) );
  XNOR U50811 ( .A(n50685), .B(n50684), .Z(n50696) );
  XOR U50812 ( .A(n50731), .B(n50681), .Z(n50684) );
  XNOR U50813 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n28322), .Z(n50681) );
  IV U50814 ( .A(p_input[2074]), .Z(n28322) );
  XOR U50815 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n29415), .Z(n50731) );
  IV U50816 ( .A(p_input[2075]), .Z(n29415) );
  XOR U50817 ( .A(\knn_comb_/min_val_out[0][28] ), .B(p_input[2076]), .Z(
        n50685) );
  XNOR U50818 ( .A(n50695), .B(n50686), .Z(n50730) );
  XNOR U50819 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n28689), .Z(n50686) );
  IV U50820 ( .A(p_input[2065]), .Z(n28689) );
  XOR U50821 ( .A(n50732), .B(n50701), .Z(n50695) );
  XNOR U50822 ( .A(\knn_comb_/min_val_out[0][31] ), .B(p_input[2079]), .Z(
        n50701) );
  XOR U50823 ( .A(n50692), .B(n50700), .Z(n50732) );
  XOR U50824 ( .A(n50733), .B(n50697), .Z(n50700) );
  XOR U50825 ( .A(\knn_comb_/min_val_out[0][29] ), .B(p_input[2077]), .Z(
        n50697) );
  XOR U50826 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n29420), .Z(n50733) );
  IV U50827 ( .A(p_input[2078]), .Z(n29420) );
  XNOR U50828 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n28326), .Z(n50692) );
  IV U50829 ( .A(p_input[2073]), .Z(n28326) );
endmodule

