
module knn_comb_BMR_W32_K1_N16 ( p_input, o );
  input [543:0] p_input;
  output [31:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/min_val_out[0][16] , \knn_comb_/min_val_out[0][17] ,
         \knn_comb_/min_val_out[0][18] , \knn_comb_/min_val_out[0][19] ,
         \knn_comb_/min_val_out[0][20] , \knn_comb_/min_val_out[0][21] ,
         \knn_comb_/min_val_out[0][22] , \knn_comb_/min_val_out[0][23] ,
         \knn_comb_/min_val_out[0][24] , \knn_comb_/min_val_out[0][25] ,
         \knn_comb_/min_val_out[0][26] , \knn_comb_/min_val_out[0][27] ,
         \knn_comb_/min_val_out[0][28] , \knn_comb_/min_val_out[0][29] ,
         \knn_comb_/min_val_out[0][30] , \knn_comb_/min_val_out[0][31] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860;
  assign \knn_comb_/min_val_out[0][0]  = p_input[480];
  assign \knn_comb_/min_val_out[0][1]  = p_input[481];
  assign \knn_comb_/min_val_out[0][2]  = p_input[482];
  assign \knn_comb_/min_val_out[0][3]  = p_input[483];
  assign \knn_comb_/min_val_out[0][4]  = p_input[484];
  assign \knn_comb_/min_val_out[0][5]  = p_input[485];
  assign \knn_comb_/min_val_out[0][6]  = p_input[486];
  assign \knn_comb_/min_val_out[0][7]  = p_input[487];
  assign \knn_comb_/min_val_out[0][8]  = p_input[488];
  assign \knn_comb_/min_val_out[0][9]  = p_input[489];
  assign \knn_comb_/min_val_out[0][10]  = p_input[490];
  assign \knn_comb_/min_val_out[0][11]  = p_input[491];
  assign \knn_comb_/min_val_out[0][12]  = p_input[492];
  assign \knn_comb_/min_val_out[0][13]  = p_input[493];
  assign \knn_comb_/min_val_out[0][14]  = p_input[494];
  assign \knn_comb_/min_val_out[0][15]  = p_input[495];
  assign \knn_comb_/min_val_out[0][16]  = p_input[496];
  assign \knn_comb_/min_val_out[0][17]  = p_input[497];
  assign \knn_comb_/min_val_out[0][18]  = p_input[498];
  assign \knn_comb_/min_val_out[0][19]  = p_input[499];
  assign \knn_comb_/min_val_out[0][20]  = p_input[500];
  assign \knn_comb_/min_val_out[0][21]  = p_input[501];
  assign \knn_comb_/min_val_out[0][22]  = p_input[502];
  assign \knn_comb_/min_val_out[0][23]  = p_input[503];
  assign \knn_comb_/min_val_out[0][24]  = p_input[504];
  assign \knn_comb_/min_val_out[0][25]  = p_input[505];
  assign \knn_comb_/min_val_out[0][26]  = p_input[506];
  assign \knn_comb_/min_val_out[0][27]  = p_input[507];
  assign \knn_comb_/min_val_out[0][28]  = p_input[508];
  assign \knn_comb_/min_val_out[0][29]  = p_input[509];
  assign \knn_comb_/min_val_out[0][30]  = p_input[510];
  assign \knn_comb_/min_val_out[0][31]  = p_input[511];

  XNOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(n3), .B(n4), .Z(n1) );
  XNOR U3 ( .A(p_input[9]), .B(n2), .Z(n4) );
  XOR U4 ( .A(n5), .B(n6), .Z(n2) );
  AND U5 ( .A(n7), .B(n8), .Z(n6) );
  XNOR U6 ( .A(p_input[41]), .B(n5), .Z(n8) );
  XOR U7 ( .A(n9), .B(n10), .Z(n5) );
  AND U8 ( .A(n11), .B(n12), .Z(n10) );
  XNOR U9 ( .A(p_input[73]), .B(n9), .Z(n12) );
  XOR U10 ( .A(n13), .B(n14), .Z(n9) );
  AND U11 ( .A(n15), .B(n16), .Z(n14) );
  XNOR U12 ( .A(p_input[105]), .B(n13), .Z(n16) );
  XOR U13 ( .A(n17), .B(n18), .Z(n13) );
  AND U14 ( .A(n19), .B(n20), .Z(n18) );
  XNOR U15 ( .A(p_input[137]), .B(n17), .Z(n20) );
  XOR U16 ( .A(n21), .B(n22), .Z(n17) );
  AND U17 ( .A(n23), .B(n24), .Z(n22) );
  XNOR U18 ( .A(p_input[169]), .B(n21), .Z(n24) );
  XOR U19 ( .A(n25), .B(n26), .Z(n21) );
  AND U20 ( .A(n27), .B(n28), .Z(n26) );
  XNOR U21 ( .A(p_input[201]), .B(n25), .Z(n28) );
  XOR U22 ( .A(n29), .B(n30), .Z(n25) );
  AND U23 ( .A(n31), .B(n32), .Z(n30) );
  XNOR U24 ( .A(p_input[233]), .B(n29), .Z(n32) );
  XOR U25 ( .A(n33), .B(n34), .Z(n29) );
  AND U26 ( .A(n35), .B(n36), .Z(n34) );
  XNOR U27 ( .A(p_input[265]), .B(n33), .Z(n36) );
  XOR U28 ( .A(n37), .B(n38), .Z(n33) );
  AND U29 ( .A(n39), .B(n40), .Z(n38) );
  XNOR U30 ( .A(p_input[297]), .B(n37), .Z(n40) );
  XOR U31 ( .A(n41), .B(n42), .Z(n37) );
  AND U32 ( .A(n43), .B(n44), .Z(n42) );
  XNOR U33 ( .A(p_input[329]), .B(n41), .Z(n44) );
  XOR U34 ( .A(n45), .B(n46), .Z(n41) );
  AND U35 ( .A(n47), .B(n48), .Z(n46) );
  XNOR U36 ( .A(p_input[361]), .B(n45), .Z(n48) );
  XOR U37 ( .A(n49), .B(n50), .Z(n45) );
  AND U38 ( .A(n51), .B(n52), .Z(n50) );
  XNOR U39 ( .A(p_input[393]), .B(n49), .Z(n52) );
  XNOR U40 ( .A(n53), .B(n54), .Z(n49) );
  AND U41 ( .A(n55), .B(n56), .Z(n54) );
  XOR U42 ( .A(p_input[425]), .B(n53), .Z(n56) );
  XOR U43 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n57), .Z(n53) );
  AND U44 ( .A(n58), .B(n59), .Z(n57) );
  XOR U45 ( .A(p_input[457]), .B(\knn_comb_/min_val_out[0][9] ), .Z(n59) );
  XNOR U46 ( .A(n60), .B(n61), .Z(o[8]) );
  AND U47 ( .A(n3), .B(n62), .Z(n60) );
  XNOR U48 ( .A(p_input[8]), .B(n61), .Z(n62) );
  XOR U49 ( .A(n63), .B(n64), .Z(n61) );
  AND U50 ( .A(n7), .B(n65), .Z(n64) );
  XNOR U51 ( .A(p_input[40]), .B(n63), .Z(n65) );
  XOR U52 ( .A(n66), .B(n67), .Z(n63) );
  AND U53 ( .A(n11), .B(n68), .Z(n67) );
  XNOR U54 ( .A(p_input[72]), .B(n66), .Z(n68) );
  XOR U55 ( .A(n69), .B(n70), .Z(n66) );
  AND U56 ( .A(n15), .B(n71), .Z(n70) );
  XNOR U57 ( .A(p_input[104]), .B(n69), .Z(n71) );
  XOR U58 ( .A(n72), .B(n73), .Z(n69) );
  AND U59 ( .A(n19), .B(n74), .Z(n73) );
  XNOR U60 ( .A(p_input[136]), .B(n72), .Z(n74) );
  XOR U61 ( .A(n75), .B(n76), .Z(n72) );
  AND U62 ( .A(n23), .B(n77), .Z(n76) );
  XNOR U63 ( .A(p_input[168]), .B(n75), .Z(n77) );
  XOR U64 ( .A(n78), .B(n79), .Z(n75) );
  AND U65 ( .A(n27), .B(n80), .Z(n79) );
  XNOR U66 ( .A(p_input[200]), .B(n78), .Z(n80) );
  XOR U67 ( .A(n81), .B(n82), .Z(n78) );
  AND U68 ( .A(n31), .B(n83), .Z(n82) );
  XNOR U69 ( .A(p_input[232]), .B(n81), .Z(n83) );
  XOR U70 ( .A(n84), .B(n85), .Z(n81) );
  AND U71 ( .A(n35), .B(n86), .Z(n85) );
  XNOR U72 ( .A(p_input[264]), .B(n84), .Z(n86) );
  XOR U73 ( .A(n87), .B(n88), .Z(n84) );
  AND U74 ( .A(n39), .B(n89), .Z(n88) );
  XNOR U75 ( .A(p_input[296]), .B(n87), .Z(n89) );
  XOR U76 ( .A(n90), .B(n91), .Z(n87) );
  AND U77 ( .A(n43), .B(n92), .Z(n91) );
  XNOR U78 ( .A(p_input[328]), .B(n90), .Z(n92) );
  XOR U79 ( .A(n93), .B(n94), .Z(n90) );
  AND U80 ( .A(n47), .B(n95), .Z(n94) );
  XNOR U81 ( .A(p_input[360]), .B(n93), .Z(n95) );
  XOR U82 ( .A(n96), .B(n97), .Z(n93) );
  AND U83 ( .A(n51), .B(n98), .Z(n97) );
  XNOR U84 ( .A(p_input[392]), .B(n96), .Z(n98) );
  XNOR U85 ( .A(n99), .B(n100), .Z(n96) );
  AND U86 ( .A(n55), .B(n101), .Z(n100) );
  XOR U87 ( .A(p_input[424]), .B(n99), .Z(n101) );
  XOR U88 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n102), .Z(n99) );
  AND U89 ( .A(n58), .B(n103), .Z(n102) );
  XOR U90 ( .A(p_input[456]), .B(\knn_comb_/min_val_out[0][8] ), .Z(n103) );
  XNOR U91 ( .A(n104), .B(n105), .Z(o[7]) );
  AND U92 ( .A(n3), .B(n106), .Z(n104) );
  XNOR U93 ( .A(p_input[7]), .B(n105), .Z(n106) );
  XOR U94 ( .A(n107), .B(n108), .Z(n105) );
  AND U95 ( .A(n7), .B(n109), .Z(n108) );
  XNOR U96 ( .A(p_input[39]), .B(n107), .Z(n109) );
  XOR U97 ( .A(n110), .B(n111), .Z(n107) );
  AND U98 ( .A(n11), .B(n112), .Z(n111) );
  XNOR U99 ( .A(p_input[71]), .B(n110), .Z(n112) );
  XOR U100 ( .A(n113), .B(n114), .Z(n110) );
  AND U101 ( .A(n15), .B(n115), .Z(n114) );
  XNOR U102 ( .A(p_input[103]), .B(n113), .Z(n115) );
  XOR U103 ( .A(n116), .B(n117), .Z(n113) );
  AND U104 ( .A(n19), .B(n118), .Z(n117) );
  XNOR U105 ( .A(p_input[135]), .B(n116), .Z(n118) );
  XOR U106 ( .A(n119), .B(n120), .Z(n116) );
  AND U107 ( .A(n23), .B(n121), .Z(n120) );
  XNOR U108 ( .A(p_input[167]), .B(n119), .Z(n121) );
  XOR U109 ( .A(n122), .B(n123), .Z(n119) );
  AND U110 ( .A(n27), .B(n124), .Z(n123) );
  XNOR U111 ( .A(p_input[199]), .B(n122), .Z(n124) );
  XOR U112 ( .A(n125), .B(n126), .Z(n122) );
  AND U113 ( .A(n31), .B(n127), .Z(n126) );
  XNOR U114 ( .A(p_input[231]), .B(n125), .Z(n127) );
  XOR U115 ( .A(n128), .B(n129), .Z(n125) );
  AND U116 ( .A(n35), .B(n130), .Z(n129) );
  XNOR U117 ( .A(p_input[263]), .B(n128), .Z(n130) );
  XOR U118 ( .A(n131), .B(n132), .Z(n128) );
  AND U119 ( .A(n39), .B(n133), .Z(n132) );
  XNOR U120 ( .A(p_input[295]), .B(n131), .Z(n133) );
  XOR U121 ( .A(n134), .B(n135), .Z(n131) );
  AND U122 ( .A(n43), .B(n136), .Z(n135) );
  XNOR U123 ( .A(p_input[327]), .B(n134), .Z(n136) );
  XOR U124 ( .A(n137), .B(n138), .Z(n134) );
  AND U125 ( .A(n47), .B(n139), .Z(n138) );
  XNOR U126 ( .A(p_input[359]), .B(n137), .Z(n139) );
  XOR U127 ( .A(n140), .B(n141), .Z(n137) );
  AND U128 ( .A(n51), .B(n142), .Z(n141) );
  XNOR U129 ( .A(p_input[391]), .B(n140), .Z(n142) );
  XNOR U130 ( .A(n143), .B(n144), .Z(n140) );
  AND U131 ( .A(n55), .B(n145), .Z(n144) );
  XOR U132 ( .A(p_input[423]), .B(n143), .Z(n145) );
  XOR U133 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n146), .Z(n143) );
  AND U134 ( .A(n58), .B(n147), .Z(n146) );
  XOR U135 ( .A(p_input[455]), .B(\knn_comb_/min_val_out[0][7] ), .Z(n147) );
  XNOR U136 ( .A(n148), .B(n149), .Z(o[6]) );
  AND U137 ( .A(n3), .B(n150), .Z(n148) );
  XNOR U138 ( .A(p_input[6]), .B(n149), .Z(n150) );
  XOR U139 ( .A(n151), .B(n152), .Z(n149) );
  AND U140 ( .A(n7), .B(n153), .Z(n152) );
  XNOR U141 ( .A(p_input[38]), .B(n151), .Z(n153) );
  XOR U142 ( .A(n154), .B(n155), .Z(n151) );
  AND U143 ( .A(n11), .B(n156), .Z(n155) );
  XNOR U144 ( .A(p_input[70]), .B(n154), .Z(n156) );
  XOR U145 ( .A(n157), .B(n158), .Z(n154) );
  AND U146 ( .A(n15), .B(n159), .Z(n158) );
  XNOR U147 ( .A(p_input[102]), .B(n157), .Z(n159) );
  XOR U148 ( .A(n160), .B(n161), .Z(n157) );
  AND U149 ( .A(n19), .B(n162), .Z(n161) );
  XNOR U150 ( .A(p_input[134]), .B(n160), .Z(n162) );
  XOR U151 ( .A(n163), .B(n164), .Z(n160) );
  AND U152 ( .A(n23), .B(n165), .Z(n164) );
  XNOR U153 ( .A(p_input[166]), .B(n163), .Z(n165) );
  XOR U154 ( .A(n166), .B(n167), .Z(n163) );
  AND U155 ( .A(n27), .B(n168), .Z(n167) );
  XNOR U156 ( .A(p_input[198]), .B(n166), .Z(n168) );
  XOR U157 ( .A(n169), .B(n170), .Z(n166) );
  AND U158 ( .A(n31), .B(n171), .Z(n170) );
  XNOR U159 ( .A(p_input[230]), .B(n169), .Z(n171) );
  XOR U160 ( .A(n172), .B(n173), .Z(n169) );
  AND U161 ( .A(n35), .B(n174), .Z(n173) );
  XNOR U162 ( .A(p_input[262]), .B(n172), .Z(n174) );
  XOR U163 ( .A(n175), .B(n176), .Z(n172) );
  AND U164 ( .A(n39), .B(n177), .Z(n176) );
  XNOR U165 ( .A(p_input[294]), .B(n175), .Z(n177) );
  XOR U166 ( .A(n178), .B(n179), .Z(n175) );
  AND U167 ( .A(n43), .B(n180), .Z(n179) );
  XNOR U168 ( .A(p_input[326]), .B(n178), .Z(n180) );
  XOR U169 ( .A(n181), .B(n182), .Z(n178) );
  AND U170 ( .A(n47), .B(n183), .Z(n182) );
  XNOR U171 ( .A(p_input[358]), .B(n181), .Z(n183) );
  XOR U172 ( .A(n184), .B(n185), .Z(n181) );
  AND U173 ( .A(n51), .B(n186), .Z(n185) );
  XNOR U174 ( .A(p_input[390]), .B(n184), .Z(n186) );
  XNOR U175 ( .A(n187), .B(n188), .Z(n184) );
  AND U176 ( .A(n55), .B(n189), .Z(n188) );
  XOR U177 ( .A(p_input[422]), .B(n187), .Z(n189) );
  XOR U178 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n190), .Z(n187) );
  AND U179 ( .A(n58), .B(n191), .Z(n190) );
  XOR U180 ( .A(p_input[454]), .B(\knn_comb_/min_val_out[0][6] ), .Z(n191) );
  XNOR U181 ( .A(n192), .B(n193), .Z(o[5]) );
  AND U182 ( .A(n3), .B(n194), .Z(n192) );
  XNOR U183 ( .A(p_input[5]), .B(n193), .Z(n194) );
  XOR U184 ( .A(n195), .B(n196), .Z(n193) );
  AND U185 ( .A(n7), .B(n197), .Z(n196) );
  XNOR U186 ( .A(p_input[37]), .B(n195), .Z(n197) );
  XOR U187 ( .A(n198), .B(n199), .Z(n195) );
  AND U188 ( .A(n11), .B(n200), .Z(n199) );
  XNOR U189 ( .A(p_input[69]), .B(n198), .Z(n200) );
  XOR U190 ( .A(n201), .B(n202), .Z(n198) );
  AND U191 ( .A(n15), .B(n203), .Z(n202) );
  XNOR U192 ( .A(p_input[101]), .B(n201), .Z(n203) );
  XOR U193 ( .A(n204), .B(n205), .Z(n201) );
  AND U194 ( .A(n19), .B(n206), .Z(n205) );
  XNOR U195 ( .A(p_input[133]), .B(n204), .Z(n206) );
  XOR U196 ( .A(n207), .B(n208), .Z(n204) );
  AND U197 ( .A(n23), .B(n209), .Z(n208) );
  XNOR U198 ( .A(p_input[165]), .B(n207), .Z(n209) );
  XOR U199 ( .A(n210), .B(n211), .Z(n207) );
  AND U200 ( .A(n27), .B(n212), .Z(n211) );
  XNOR U201 ( .A(p_input[197]), .B(n210), .Z(n212) );
  XOR U202 ( .A(n213), .B(n214), .Z(n210) );
  AND U203 ( .A(n31), .B(n215), .Z(n214) );
  XNOR U204 ( .A(p_input[229]), .B(n213), .Z(n215) );
  XOR U205 ( .A(n216), .B(n217), .Z(n213) );
  AND U206 ( .A(n35), .B(n218), .Z(n217) );
  XNOR U207 ( .A(p_input[261]), .B(n216), .Z(n218) );
  XOR U208 ( .A(n219), .B(n220), .Z(n216) );
  AND U209 ( .A(n39), .B(n221), .Z(n220) );
  XNOR U210 ( .A(p_input[293]), .B(n219), .Z(n221) );
  XOR U211 ( .A(n222), .B(n223), .Z(n219) );
  AND U212 ( .A(n43), .B(n224), .Z(n223) );
  XNOR U213 ( .A(p_input[325]), .B(n222), .Z(n224) );
  XOR U214 ( .A(n225), .B(n226), .Z(n222) );
  AND U215 ( .A(n47), .B(n227), .Z(n226) );
  XNOR U216 ( .A(p_input[357]), .B(n225), .Z(n227) );
  XOR U217 ( .A(n228), .B(n229), .Z(n225) );
  AND U218 ( .A(n51), .B(n230), .Z(n229) );
  XNOR U219 ( .A(p_input[389]), .B(n228), .Z(n230) );
  XNOR U220 ( .A(n231), .B(n232), .Z(n228) );
  AND U221 ( .A(n55), .B(n233), .Z(n232) );
  XOR U222 ( .A(p_input[421]), .B(n231), .Z(n233) );
  XOR U223 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n234), .Z(n231) );
  AND U224 ( .A(n58), .B(n235), .Z(n234) );
  XOR U225 ( .A(p_input[453]), .B(\knn_comb_/min_val_out[0][5] ), .Z(n235) );
  XNOR U226 ( .A(n236), .B(n237), .Z(o[4]) );
  AND U227 ( .A(n3), .B(n238), .Z(n236) );
  XNOR U228 ( .A(p_input[4]), .B(n237), .Z(n238) );
  XOR U229 ( .A(n239), .B(n240), .Z(n237) );
  AND U230 ( .A(n7), .B(n241), .Z(n240) );
  XNOR U231 ( .A(p_input[36]), .B(n239), .Z(n241) );
  XOR U232 ( .A(n242), .B(n243), .Z(n239) );
  AND U233 ( .A(n11), .B(n244), .Z(n243) );
  XNOR U234 ( .A(p_input[68]), .B(n242), .Z(n244) );
  XOR U235 ( .A(n245), .B(n246), .Z(n242) );
  AND U236 ( .A(n15), .B(n247), .Z(n246) );
  XNOR U237 ( .A(p_input[100]), .B(n245), .Z(n247) );
  XOR U238 ( .A(n248), .B(n249), .Z(n245) );
  AND U239 ( .A(n19), .B(n250), .Z(n249) );
  XNOR U240 ( .A(p_input[132]), .B(n248), .Z(n250) );
  XOR U241 ( .A(n251), .B(n252), .Z(n248) );
  AND U242 ( .A(n23), .B(n253), .Z(n252) );
  XNOR U243 ( .A(p_input[164]), .B(n251), .Z(n253) );
  XOR U244 ( .A(n254), .B(n255), .Z(n251) );
  AND U245 ( .A(n27), .B(n256), .Z(n255) );
  XNOR U246 ( .A(p_input[196]), .B(n254), .Z(n256) );
  XOR U247 ( .A(n257), .B(n258), .Z(n254) );
  AND U248 ( .A(n31), .B(n259), .Z(n258) );
  XNOR U249 ( .A(p_input[228]), .B(n257), .Z(n259) );
  XOR U250 ( .A(n260), .B(n261), .Z(n257) );
  AND U251 ( .A(n35), .B(n262), .Z(n261) );
  XNOR U252 ( .A(p_input[260]), .B(n260), .Z(n262) );
  XOR U253 ( .A(n263), .B(n264), .Z(n260) );
  AND U254 ( .A(n39), .B(n265), .Z(n264) );
  XNOR U255 ( .A(p_input[292]), .B(n263), .Z(n265) );
  XOR U256 ( .A(n266), .B(n267), .Z(n263) );
  AND U257 ( .A(n43), .B(n268), .Z(n267) );
  XNOR U258 ( .A(p_input[324]), .B(n266), .Z(n268) );
  XOR U259 ( .A(n269), .B(n270), .Z(n266) );
  AND U260 ( .A(n47), .B(n271), .Z(n270) );
  XNOR U261 ( .A(p_input[356]), .B(n269), .Z(n271) );
  XOR U262 ( .A(n272), .B(n273), .Z(n269) );
  AND U263 ( .A(n51), .B(n274), .Z(n273) );
  XNOR U264 ( .A(p_input[388]), .B(n272), .Z(n274) );
  XNOR U265 ( .A(n275), .B(n276), .Z(n272) );
  AND U266 ( .A(n55), .B(n277), .Z(n276) );
  XOR U267 ( .A(p_input[420]), .B(n275), .Z(n277) );
  XOR U268 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n278), .Z(n275) );
  AND U269 ( .A(n58), .B(n279), .Z(n278) );
  XOR U270 ( .A(p_input[452]), .B(\knn_comb_/min_val_out[0][4] ), .Z(n279) );
  XNOR U271 ( .A(n280), .B(n281), .Z(o[3]) );
  AND U272 ( .A(n3), .B(n282), .Z(n280) );
  XNOR U273 ( .A(p_input[3]), .B(n281), .Z(n282) );
  XOR U274 ( .A(n283), .B(n284), .Z(n281) );
  AND U275 ( .A(n7), .B(n285), .Z(n284) );
  XNOR U276 ( .A(p_input[35]), .B(n283), .Z(n285) );
  XOR U277 ( .A(n286), .B(n287), .Z(n283) );
  AND U278 ( .A(n11), .B(n288), .Z(n287) );
  XNOR U279 ( .A(p_input[67]), .B(n286), .Z(n288) );
  XOR U280 ( .A(n289), .B(n290), .Z(n286) );
  AND U281 ( .A(n15), .B(n291), .Z(n290) );
  XNOR U282 ( .A(p_input[99]), .B(n289), .Z(n291) );
  XOR U283 ( .A(n292), .B(n293), .Z(n289) );
  AND U284 ( .A(n19), .B(n294), .Z(n293) );
  XNOR U285 ( .A(p_input[131]), .B(n292), .Z(n294) );
  XOR U286 ( .A(n295), .B(n296), .Z(n292) );
  AND U287 ( .A(n23), .B(n297), .Z(n296) );
  XNOR U288 ( .A(p_input[163]), .B(n295), .Z(n297) );
  XOR U289 ( .A(n298), .B(n299), .Z(n295) );
  AND U290 ( .A(n27), .B(n300), .Z(n299) );
  XNOR U291 ( .A(p_input[195]), .B(n298), .Z(n300) );
  XOR U292 ( .A(n301), .B(n302), .Z(n298) );
  AND U293 ( .A(n31), .B(n303), .Z(n302) );
  XNOR U294 ( .A(p_input[227]), .B(n301), .Z(n303) );
  XOR U295 ( .A(n304), .B(n305), .Z(n301) );
  AND U296 ( .A(n35), .B(n306), .Z(n305) );
  XNOR U297 ( .A(p_input[259]), .B(n304), .Z(n306) );
  XOR U298 ( .A(n307), .B(n308), .Z(n304) );
  AND U299 ( .A(n39), .B(n309), .Z(n308) );
  XNOR U300 ( .A(p_input[291]), .B(n307), .Z(n309) );
  XOR U301 ( .A(n310), .B(n311), .Z(n307) );
  AND U302 ( .A(n43), .B(n312), .Z(n311) );
  XNOR U303 ( .A(p_input[323]), .B(n310), .Z(n312) );
  XOR U304 ( .A(n313), .B(n314), .Z(n310) );
  AND U305 ( .A(n47), .B(n315), .Z(n314) );
  XNOR U306 ( .A(p_input[355]), .B(n313), .Z(n315) );
  XOR U307 ( .A(n316), .B(n317), .Z(n313) );
  AND U308 ( .A(n51), .B(n318), .Z(n317) );
  XNOR U309 ( .A(p_input[387]), .B(n316), .Z(n318) );
  XNOR U310 ( .A(n319), .B(n320), .Z(n316) );
  AND U311 ( .A(n55), .B(n321), .Z(n320) );
  XOR U312 ( .A(p_input[419]), .B(n319), .Z(n321) );
  XOR U313 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n322), .Z(n319) );
  AND U314 ( .A(n58), .B(n323), .Z(n322) );
  XOR U315 ( .A(p_input[451]), .B(\knn_comb_/min_val_out[0][3] ), .Z(n323) );
  XNOR U316 ( .A(n324), .B(n325), .Z(o[31]) );
  AND U317 ( .A(n3), .B(n326), .Z(n324) );
  XNOR U318 ( .A(p_input[31]), .B(n325), .Z(n326) );
  XOR U319 ( .A(n327), .B(n328), .Z(n325) );
  AND U320 ( .A(n7), .B(n329), .Z(n328) );
  XNOR U321 ( .A(p_input[63]), .B(n327), .Z(n329) );
  XOR U322 ( .A(n330), .B(n331), .Z(n327) );
  AND U323 ( .A(n11), .B(n332), .Z(n331) );
  XNOR U324 ( .A(p_input[95]), .B(n330), .Z(n332) );
  XOR U325 ( .A(n333), .B(n334), .Z(n330) );
  AND U326 ( .A(n15), .B(n335), .Z(n334) );
  XNOR U327 ( .A(p_input[127]), .B(n333), .Z(n335) );
  XOR U328 ( .A(n336), .B(n337), .Z(n333) );
  AND U329 ( .A(n19), .B(n338), .Z(n337) );
  XNOR U330 ( .A(p_input[159]), .B(n336), .Z(n338) );
  XOR U331 ( .A(n339), .B(n340), .Z(n336) );
  AND U332 ( .A(n23), .B(n341), .Z(n340) );
  XNOR U333 ( .A(p_input[191]), .B(n339), .Z(n341) );
  XOR U334 ( .A(n342), .B(n343), .Z(n339) );
  AND U335 ( .A(n27), .B(n344), .Z(n343) );
  XNOR U336 ( .A(p_input[223]), .B(n342), .Z(n344) );
  XOR U337 ( .A(n345), .B(n346), .Z(n342) );
  AND U338 ( .A(n31), .B(n347), .Z(n346) );
  XNOR U339 ( .A(p_input[255]), .B(n345), .Z(n347) );
  XOR U340 ( .A(n348), .B(n349), .Z(n345) );
  AND U341 ( .A(n35), .B(n350), .Z(n349) );
  XNOR U342 ( .A(p_input[287]), .B(n348), .Z(n350) );
  XOR U343 ( .A(n351), .B(n352), .Z(n348) );
  AND U344 ( .A(n39), .B(n353), .Z(n352) );
  XNOR U345 ( .A(p_input[319]), .B(n351), .Z(n353) );
  XOR U346 ( .A(n354), .B(n355), .Z(n351) );
  AND U347 ( .A(n43), .B(n356), .Z(n355) );
  XNOR U348 ( .A(p_input[351]), .B(n354), .Z(n356) );
  XOR U349 ( .A(n357), .B(n358), .Z(n354) );
  AND U350 ( .A(n47), .B(n359), .Z(n358) );
  XNOR U351 ( .A(p_input[383]), .B(n357), .Z(n359) );
  XOR U352 ( .A(n360), .B(n361), .Z(n357) );
  AND U353 ( .A(n51), .B(n362), .Z(n361) );
  XNOR U354 ( .A(p_input[415]), .B(n360), .Z(n362) );
  XNOR U355 ( .A(n363), .B(n364), .Z(n360) );
  AND U356 ( .A(n55), .B(n365), .Z(n364) );
  XOR U357 ( .A(p_input[447]), .B(n363), .Z(n365) );
  XOR U358 ( .A(\knn_comb_/min_val_out[0][31] ), .B(n366), .Z(n363) );
  AND U359 ( .A(n58), .B(n367), .Z(n366) );
  XOR U360 ( .A(p_input[479]), .B(\knn_comb_/min_val_out[0][31] ), .Z(n367) );
  XNOR U361 ( .A(n368), .B(n369), .Z(o[30]) );
  AND U362 ( .A(n3), .B(n370), .Z(n368) );
  XNOR U363 ( .A(p_input[30]), .B(n369), .Z(n370) );
  XOR U364 ( .A(n371), .B(n372), .Z(n369) );
  AND U365 ( .A(n7), .B(n373), .Z(n372) );
  XNOR U366 ( .A(p_input[62]), .B(n371), .Z(n373) );
  XOR U367 ( .A(n374), .B(n375), .Z(n371) );
  AND U368 ( .A(n11), .B(n376), .Z(n375) );
  XNOR U369 ( .A(p_input[94]), .B(n374), .Z(n376) );
  XOR U370 ( .A(n377), .B(n378), .Z(n374) );
  AND U371 ( .A(n15), .B(n379), .Z(n378) );
  XNOR U372 ( .A(p_input[126]), .B(n377), .Z(n379) );
  XOR U373 ( .A(n380), .B(n381), .Z(n377) );
  AND U374 ( .A(n19), .B(n382), .Z(n381) );
  XNOR U375 ( .A(p_input[158]), .B(n380), .Z(n382) );
  XOR U376 ( .A(n383), .B(n384), .Z(n380) );
  AND U377 ( .A(n23), .B(n385), .Z(n384) );
  XNOR U378 ( .A(p_input[190]), .B(n383), .Z(n385) );
  XOR U379 ( .A(n386), .B(n387), .Z(n383) );
  AND U380 ( .A(n27), .B(n388), .Z(n387) );
  XNOR U381 ( .A(p_input[222]), .B(n386), .Z(n388) );
  XOR U382 ( .A(n389), .B(n390), .Z(n386) );
  AND U383 ( .A(n31), .B(n391), .Z(n390) );
  XNOR U384 ( .A(p_input[254]), .B(n389), .Z(n391) );
  XOR U385 ( .A(n392), .B(n393), .Z(n389) );
  AND U386 ( .A(n35), .B(n394), .Z(n393) );
  XNOR U387 ( .A(p_input[286]), .B(n392), .Z(n394) );
  XOR U388 ( .A(n395), .B(n396), .Z(n392) );
  AND U389 ( .A(n39), .B(n397), .Z(n396) );
  XNOR U390 ( .A(p_input[318]), .B(n395), .Z(n397) );
  XOR U391 ( .A(n398), .B(n399), .Z(n395) );
  AND U392 ( .A(n43), .B(n400), .Z(n399) );
  XNOR U393 ( .A(p_input[350]), .B(n398), .Z(n400) );
  XOR U394 ( .A(n401), .B(n402), .Z(n398) );
  AND U395 ( .A(n47), .B(n403), .Z(n402) );
  XNOR U396 ( .A(p_input[382]), .B(n401), .Z(n403) );
  XOR U397 ( .A(n404), .B(n405), .Z(n401) );
  AND U398 ( .A(n51), .B(n406), .Z(n405) );
  XNOR U399 ( .A(p_input[414]), .B(n404), .Z(n406) );
  XNOR U400 ( .A(n407), .B(n408), .Z(n404) );
  AND U401 ( .A(n55), .B(n409), .Z(n408) );
  XOR U402 ( .A(p_input[446]), .B(n407), .Z(n409) );
  XOR U403 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n410), .Z(n407) );
  AND U404 ( .A(n58), .B(n411), .Z(n410) );
  XOR U405 ( .A(p_input[478]), .B(\knn_comb_/min_val_out[0][30] ), .Z(n411) );
  XNOR U406 ( .A(n412), .B(n413), .Z(o[2]) );
  AND U407 ( .A(n3), .B(n414), .Z(n412) );
  XNOR U408 ( .A(p_input[2]), .B(n413), .Z(n414) );
  XOR U409 ( .A(n415), .B(n416), .Z(n413) );
  AND U410 ( .A(n7), .B(n417), .Z(n416) );
  XNOR U411 ( .A(p_input[34]), .B(n415), .Z(n417) );
  XOR U412 ( .A(n418), .B(n419), .Z(n415) );
  AND U413 ( .A(n11), .B(n420), .Z(n419) );
  XNOR U414 ( .A(p_input[66]), .B(n418), .Z(n420) );
  XOR U415 ( .A(n421), .B(n422), .Z(n418) );
  AND U416 ( .A(n15), .B(n423), .Z(n422) );
  XNOR U417 ( .A(p_input[98]), .B(n421), .Z(n423) );
  XOR U418 ( .A(n424), .B(n425), .Z(n421) );
  AND U419 ( .A(n19), .B(n426), .Z(n425) );
  XNOR U420 ( .A(p_input[130]), .B(n424), .Z(n426) );
  XOR U421 ( .A(n427), .B(n428), .Z(n424) );
  AND U422 ( .A(n23), .B(n429), .Z(n428) );
  XNOR U423 ( .A(p_input[162]), .B(n427), .Z(n429) );
  XOR U424 ( .A(n430), .B(n431), .Z(n427) );
  AND U425 ( .A(n27), .B(n432), .Z(n431) );
  XNOR U426 ( .A(p_input[194]), .B(n430), .Z(n432) );
  XOR U427 ( .A(n433), .B(n434), .Z(n430) );
  AND U428 ( .A(n31), .B(n435), .Z(n434) );
  XNOR U429 ( .A(p_input[226]), .B(n433), .Z(n435) );
  XOR U430 ( .A(n436), .B(n437), .Z(n433) );
  AND U431 ( .A(n35), .B(n438), .Z(n437) );
  XNOR U432 ( .A(p_input[258]), .B(n436), .Z(n438) );
  XOR U433 ( .A(n439), .B(n440), .Z(n436) );
  AND U434 ( .A(n39), .B(n441), .Z(n440) );
  XNOR U435 ( .A(p_input[290]), .B(n439), .Z(n441) );
  XOR U436 ( .A(n442), .B(n443), .Z(n439) );
  AND U437 ( .A(n43), .B(n444), .Z(n443) );
  XNOR U438 ( .A(p_input[322]), .B(n442), .Z(n444) );
  XOR U439 ( .A(n445), .B(n446), .Z(n442) );
  AND U440 ( .A(n47), .B(n447), .Z(n446) );
  XNOR U441 ( .A(p_input[354]), .B(n445), .Z(n447) );
  XOR U442 ( .A(n448), .B(n449), .Z(n445) );
  AND U443 ( .A(n51), .B(n450), .Z(n449) );
  XNOR U444 ( .A(p_input[386]), .B(n448), .Z(n450) );
  XNOR U445 ( .A(n451), .B(n452), .Z(n448) );
  AND U446 ( .A(n55), .B(n453), .Z(n452) );
  XOR U447 ( .A(p_input[418]), .B(n451), .Z(n453) );
  XOR U448 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n454), .Z(n451) );
  AND U449 ( .A(n58), .B(n455), .Z(n454) );
  XOR U450 ( .A(p_input[450]), .B(\knn_comb_/min_val_out[0][2] ), .Z(n455) );
  XNOR U451 ( .A(n456), .B(n457), .Z(o[29]) );
  AND U452 ( .A(n3), .B(n458), .Z(n456) );
  XNOR U453 ( .A(p_input[29]), .B(n457), .Z(n458) );
  XOR U454 ( .A(n459), .B(n460), .Z(n457) );
  AND U455 ( .A(n7), .B(n461), .Z(n460) );
  XNOR U456 ( .A(p_input[61]), .B(n459), .Z(n461) );
  XOR U457 ( .A(n462), .B(n463), .Z(n459) );
  AND U458 ( .A(n11), .B(n464), .Z(n463) );
  XNOR U459 ( .A(p_input[93]), .B(n462), .Z(n464) );
  XOR U460 ( .A(n465), .B(n466), .Z(n462) );
  AND U461 ( .A(n15), .B(n467), .Z(n466) );
  XNOR U462 ( .A(p_input[125]), .B(n465), .Z(n467) );
  XOR U463 ( .A(n468), .B(n469), .Z(n465) );
  AND U464 ( .A(n19), .B(n470), .Z(n469) );
  XNOR U465 ( .A(p_input[157]), .B(n468), .Z(n470) );
  XOR U466 ( .A(n471), .B(n472), .Z(n468) );
  AND U467 ( .A(n23), .B(n473), .Z(n472) );
  XNOR U468 ( .A(p_input[189]), .B(n471), .Z(n473) );
  XOR U469 ( .A(n474), .B(n475), .Z(n471) );
  AND U470 ( .A(n27), .B(n476), .Z(n475) );
  XNOR U471 ( .A(p_input[221]), .B(n474), .Z(n476) );
  XOR U472 ( .A(n477), .B(n478), .Z(n474) );
  AND U473 ( .A(n31), .B(n479), .Z(n478) );
  XNOR U474 ( .A(p_input[253]), .B(n477), .Z(n479) );
  XOR U475 ( .A(n480), .B(n481), .Z(n477) );
  AND U476 ( .A(n35), .B(n482), .Z(n481) );
  XNOR U477 ( .A(p_input[285]), .B(n480), .Z(n482) );
  XOR U478 ( .A(n483), .B(n484), .Z(n480) );
  AND U479 ( .A(n39), .B(n485), .Z(n484) );
  XNOR U480 ( .A(p_input[317]), .B(n483), .Z(n485) );
  XOR U481 ( .A(n486), .B(n487), .Z(n483) );
  AND U482 ( .A(n43), .B(n488), .Z(n487) );
  XNOR U483 ( .A(p_input[349]), .B(n486), .Z(n488) );
  XOR U484 ( .A(n489), .B(n490), .Z(n486) );
  AND U485 ( .A(n47), .B(n491), .Z(n490) );
  XNOR U486 ( .A(p_input[381]), .B(n489), .Z(n491) );
  XOR U487 ( .A(n492), .B(n493), .Z(n489) );
  AND U488 ( .A(n51), .B(n494), .Z(n493) );
  XNOR U489 ( .A(p_input[413]), .B(n492), .Z(n494) );
  XNOR U490 ( .A(n495), .B(n496), .Z(n492) );
  AND U491 ( .A(n55), .B(n497), .Z(n496) );
  XOR U492 ( .A(p_input[445]), .B(n495), .Z(n497) );
  XOR U493 ( .A(\knn_comb_/min_val_out[0][29] ), .B(n498), .Z(n495) );
  AND U494 ( .A(n58), .B(n499), .Z(n498) );
  XOR U495 ( .A(p_input[477]), .B(\knn_comb_/min_val_out[0][29] ), .Z(n499) );
  XNOR U496 ( .A(n500), .B(n501), .Z(o[28]) );
  AND U497 ( .A(n3), .B(n502), .Z(n500) );
  XNOR U498 ( .A(p_input[28]), .B(n501), .Z(n502) );
  XOR U499 ( .A(n503), .B(n504), .Z(n501) );
  AND U500 ( .A(n7), .B(n505), .Z(n504) );
  XNOR U501 ( .A(p_input[60]), .B(n503), .Z(n505) );
  XOR U502 ( .A(n506), .B(n507), .Z(n503) );
  AND U503 ( .A(n11), .B(n508), .Z(n507) );
  XNOR U504 ( .A(p_input[92]), .B(n506), .Z(n508) );
  XOR U505 ( .A(n509), .B(n510), .Z(n506) );
  AND U506 ( .A(n15), .B(n511), .Z(n510) );
  XNOR U507 ( .A(p_input[124]), .B(n509), .Z(n511) );
  XOR U508 ( .A(n512), .B(n513), .Z(n509) );
  AND U509 ( .A(n19), .B(n514), .Z(n513) );
  XNOR U510 ( .A(p_input[156]), .B(n512), .Z(n514) );
  XOR U511 ( .A(n515), .B(n516), .Z(n512) );
  AND U512 ( .A(n23), .B(n517), .Z(n516) );
  XNOR U513 ( .A(p_input[188]), .B(n515), .Z(n517) );
  XOR U514 ( .A(n518), .B(n519), .Z(n515) );
  AND U515 ( .A(n27), .B(n520), .Z(n519) );
  XNOR U516 ( .A(p_input[220]), .B(n518), .Z(n520) );
  XOR U517 ( .A(n521), .B(n522), .Z(n518) );
  AND U518 ( .A(n31), .B(n523), .Z(n522) );
  XNOR U519 ( .A(p_input[252]), .B(n521), .Z(n523) );
  XOR U520 ( .A(n524), .B(n525), .Z(n521) );
  AND U521 ( .A(n35), .B(n526), .Z(n525) );
  XNOR U522 ( .A(p_input[284]), .B(n524), .Z(n526) );
  XOR U523 ( .A(n527), .B(n528), .Z(n524) );
  AND U524 ( .A(n39), .B(n529), .Z(n528) );
  XNOR U525 ( .A(p_input[316]), .B(n527), .Z(n529) );
  XOR U526 ( .A(n530), .B(n531), .Z(n527) );
  AND U527 ( .A(n43), .B(n532), .Z(n531) );
  XNOR U528 ( .A(p_input[348]), .B(n530), .Z(n532) );
  XOR U529 ( .A(n533), .B(n534), .Z(n530) );
  AND U530 ( .A(n47), .B(n535), .Z(n534) );
  XNOR U531 ( .A(p_input[380]), .B(n533), .Z(n535) );
  XOR U532 ( .A(n536), .B(n537), .Z(n533) );
  AND U533 ( .A(n51), .B(n538), .Z(n537) );
  XNOR U534 ( .A(p_input[412]), .B(n536), .Z(n538) );
  XNOR U535 ( .A(n539), .B(n540), .Z(n536) );
  AND U536 ( .A(n55), .B(n541), .Z(n540) );
  XOR U537 ( .A(p_input[444]), .B(n539), .Z(n541) );
  XOR U538 ( .A(\knn_comb_/min_val_out[0][28] ), .B(n542), .Z(n539) );
  AND U539 ( .A(n58), .B(n543), .Z(n542) );
  XOR U540 ( .A(p_input[476]), .B(\knn_comb_/min_val_out[0][28] ), .Z(n543) );
  XNOR U541 ( .A(n544), .B(n545), .Z(o[27]) );
  AND U542 ( .A(n3), .B(n546), .Z(n544) );
  XNOR U543 ( .A(p_input[27]), .B(n545), .Z(n546) );
  XOR U544 ( .A(n547), .B(n548), .Z(n545) );
  AND U545 ( .A(n7), .B(n549), .Z(n548) );
  XNOR U546 ( .A(p_input[59]), .B(n547), .Z(n549) );
  XOR U547 ( .A(n550), .B(n551), .Z(n547) );
  AND U548 ( .A(n11), .B(n552), .Z(n551) );
  XNOR U549 ( .A(p_input[91]), .B(n550), .Z(n552) );
  XOR U550 ( .A(n553), .B(n554), .Z(n550) );
  AND U551 ( .A(n15), .B(n555), .Z(n554) );
  XNOR U552 ( .A(p_input[123]), .B(n553), .Z(n555) );
  XOR U553 ( .A(n556), .B(n557), .Z(n553) );
  AND U554 ( .A(n19), .B(n558), .Z(n557) );
  XNOR U555 ( .A(p_input[155]), .B(n556), .Z(n558) );
  XOR U556 ( .A(n559), .B(n560), .Z(n556) );
  AND U557 ( .A(n23), .B(n561), .Z(n560) );
  XNOR U558 ( .A(p_input[187]), .B(n559), .Z(n561) );
  XOR U559 ( .A(n562), .B(n563), .Z(n559) );
  AND U560 ( .A(n27), .B(n564), .Z(n563) );
  XNOR U561 ( .A(p_input[219]), .B(n562), .Z(n564) );
  XOR U562 ( .A(n565), .B(n566), .Z(n562) );
  AND U563 ( .A(n31), .B(n567), .Z(n566) );
  XNOR U564 ( .A(p_input[251]), .B(n565), .Z(n567) );
  XOR U565 ( .A(n568), .B(n569), .Z(n565) );
  AND U566 ( .A(n35), .B(n570), .Z(n569) );
  XNOR U567 ( .A(p_input[283]), .B(n568), .Z(n570) );
  XOR U568 ( .A(n571), .B(n572), .Z(n568) );
  AND U569 ( .A(n39), .B(n573), .Z(n572) );
  XNOR U570 ( .A(p_input[315]), .B(n571), .Z(n573) );
  XOR U571 ( .A(n574), .B(n575), .Z(n571) );
  AND U572 ( .A(n43), .B(n576), .Z(n575) );
  XNOR U573 ( .A(p_input[347]), .B(n574), .Z(n576) );
  XOR U574 ( .A(n577), .B(n578), .Z(n574) );
  AND U575 ( .A(n47), .B(n579), .Z(n578) );
  XNOR U576 ( .A(p_input[379]), .B(n577), .Z(n579) );
  XOR U577 ( .A(n580), .B(n581), .Z(n577) );
  AND U578 ( .A(n51), .B(n582), .Z(n581) );
  XNOR U579 ( .A(p_input[411]), .B(n580), .Z(n582) );
  XNOR U580 ( .A(n583), .B(n584), .Z(n580) );
  AND U581 ( .A(n55), .B(n585), .Z(n584) );
  XOR U582 ( .A(p_input[443]), .B(n583), .Z(n585) );
  XOR U583 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n586), .Z(n583) );
  AND U584 ( .A(n58), .B(n587), .Z(n586) );
  XOR U585 ( .A(p_input[475]), .B(\knn_comb_/min_val_out[0][27] ), .Z(n587) );
  XNOR U586 ( .A(n588), .B(n589), .Z(o[26]) );
  AND U587 ( .A(n3), .B(n590), .Z(n588) );
  XNOR U588 ( .A(p_input[26]), .B(n589), .Z(n590) );
  XOR U589 ( .A(n591), .B(n592), .Z(n589) );
  AND U590 ( .A(n7), .B(n593), .Z(n592) );
  XNOR U591 ( .A(p_input[58]), .B(n591), .Z(n593) );
  XOR U592 ( .A(n594), .B(n595), .Z(n591) );
  AND U593 ( .A(n11), .B(n596), .Z(n595) );
  XNOR U594 ( .A(p_input[90]), .B(n594), .Z(n596) );
  XOR U595 ( .A(n597), .B(n598), .Z(n594) );
  AND U596 ( .A(n15), .B(n599), .Z(n598) );
  XNOR U597 ( .A(p_input[122]), .B(n597), .Z(n599) );
  XOR U598 ( .A(n600), .B(n601), .Z(n597) );
  AND U599 ( .A(n19), .B(n602), .Z(n601) );
  XNOR U600 ( .A(p_input[154]), .B(n600), .Z(n602) );
  XOR U601 ( .A(n603), .B(n604), .Z(n600) );
  AND U602 ( .A(n23), .B(n605), .Z(n604) );
  XNOR U603 ( .A(p_input[186]), .B(n603), .Z(n605) );
  XOR U604 ( .A(n606), .B(n607), .Z(n603) );
  AND U605 ( .A(n27), .B(n608), .Z(n607) );
  XNOR U606 ( .A(p_input[218]), .B(n606), .Z(n608) );
  XOR U607 ( .A(n609), .B(n610), .Z(n606) );
  AND U608 ( .A(n31), .B(n611), .Z(n610) );
  XNOR U609 ( .A(p_input[250]), .B(n609), .Z(n611) );
  XOR U610 ( .A(n612), .B(n613), .Z(n609) );
  AND U611 ( .A(n35), .B(n614), .Z(n613) );
  XNOR U612 ( .A(p_input[282]), .B(n612), .Z(n614) );
  XOR U613 ( .A(n615), .B(n616), .Z(n612) );
  AND U614 ( .A(n39), .B(n617), .Z(n616) );
  XNOR U615 ( .A(p_input[314]), .B(n615), .Z(n617) );
  XOR U616 ( .A(n618), .B(n619), .Z(n615) );
  AND U617 ( .A(n43), .B(n620), .Z(n619) );
  XNOR U618 ( .A(p_input[346]), .B(n618), .Z(n620) );
  XOR U619 ( .A(n621), .B(n622), .Z(n618) );
  AND U620 ( .A(n47), .B(n623), .Z(n622) );
  XNOR U621 ( .A(p_input[378]), .B(n621), .Z(n623) );
  XOR U622 ( .A(n624), .B(n625), .Z(n621) );
  AND U623 ( .A(n51), .B(n626), .Z(n625) );
  XNOR U624 ( .A(p_input[410]), .B(n624), .Z(n626) );
  XNOR U625 ( .A(n627), .B(n628), .Z(n624) );
  AND U626 ( .A(n55), .B(n629), .Z(n628) );
  XOR U627 ( .A(p_input[442]), .B(n627), .Z(n629) );
  XOR U628 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n630), .Z(n627) );
  AND U629 ( .A(n58), .B(n631), .Z(n630) );
  XOR U630 ( .A(p_input[474]), .B(\knn_comb_/min_val_out[0][26] ), .Z(n631) );
  XNOR U631 ( .A(n632), .B(n633), .Z(o[25]) );
  AND U632 ( .A(n3), .B(n634), .Z(n632) );
  XNOR U633 ( .A(p_input[25]), .B(n633), .Z(n634) );
  XOR U634 ( .A(n635), .B(n636), .Z(n633) );
  AND U635 ( .A(n7), .B(n637), .Z(n636) );
  XNOR U636 ( .A(p_input[57]), .B(n635), .Z(n637) );
  XOR U637 ( .A(n638), .B(n639), .Z(n635) );
  AND U638 ( .A(n11), .B(n640), .Z(n639) );
  XNOR U639 ( .A(p_input[89]), .B(n638), .Z(n640) );
  XOR U640 ( .A(n641), .B(n642), .Z(n638) );
  AND U641 ( .A(n15), .B(n643), .Z(n642) );
  XNOR U642 ( .A(p_input[121]), .B(n641), .Z(n643) );
  XOR U643 ( .A(n644), .B(n645), .Z(n641) );
  AND U644 ( .A(n19), .B(n646), .Z(n645) );
  XNOR U645 ( .A(p_input[153]), .B(n644), .Z(n646) );
  XOR U646 ( .A(n647), .B(n648), .Z(n644) );
  AND U647 ( .A(n23), .B(n649), .Z(n648) );
  XNOR U648 ( .A(p_input[185]), .B(n647), .Z(n649) );
  XOR U649 ( .A(n650), .B(n651), .Z(n647) );
  AND U650 ( .A(n27), .B(n652), .Z(n651) );
  XNOR U651 ( .A(p_input[217]), .B(n650), .Z(n652) );
  XOR U652 ( .A(n653), .B(n654), .Z(n650) );
  AND U653 ( .A(n31), .B(n655), .Z(n654) );
  XNOR U654 ( .A(p_input[249]), .B(n653), .Z(n655) );
  XOR U655 ( .A(n656), .B(n657), .Z(n653) );
  AND U656 ( .A(n35), .B(n658), .Z(n657) );
  XNOR U657 ( .A(p_input[281]), .B(n656), .Z(n658) );
  XOR U658 ( .A(n659), .B(n660), .Z(n656) );
  AND U659 ( .A(n39), .B(n661), .Z(n660) );
  XNOR U660 ( .A(p_input[313]), .B(n659), .Z(n661) );
  XOR U661 ( .A(n662), .B(n663), .Z(n659) );
  AND U662 ( .A(n43), .B(n664), .Z(n663) );
  XNOR U663 ( .A(p_input[345]), .B(n662), .Z(n664) );
  XOR U664 ( .A(n665), .B(n666), .Z(n662) );
  AND U665 ( .A(n47), .B(n667), .Z(n666) );
  XNOR U666 ( .A(p_input[377]), .B(n665), .Z(n667) );
  XOR U667 ( .A(n668), .B(n669), .Z(n665) );
  AND U668 ( .A(n51), .B(n670), .Z(n669) );
  XNOR U669 ( .A(p_input[409]), .B(n668), .Z(n670) );
  XNOR U670 ( .A(n671), .B(n672), .Z(n668) );
  AND U671 ( .A(n55), .B(n673), .Z(n672) );
  XOR U672 ( .A(p_input[441]), .B(n671), .Z(n673) );
  XOR U673 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n674), .Z(n671) );
  AND U674 ( .A(n58), .B(n675), .Z(n674) );
  XOR U675 ( .A(p_input[473]), .B(\knn_comb_/min_val_out[0][25] ), .Z(n675) );
  XNOR U676 ( .A(n676), .B(n677), .Z(o[24]) );
  AND U677 ( .A(n3), .B(n678), .Z(n676) );
  XNOR U678 ( .A(p_input[24]), .B(n677), .Z(n678) );
  XOR U679 ( .A(n679), .B(n680), .Z(n677) );
  AND U680 ( .A(n7), .B(n681), .Z(n680) );
  XNOR U681 ( .A(p_input[56]), .B(n679), .Z(n681) );
  XOR U682 ( .A(n682), .B(n683), .Z(n679) );
  AND U683 ( .A(n11), .B(n684), .Z(n683) );
  XNOR U684 ( .A(p_input[88]), .B(n682), .Z(n684) );
  XOR U685 ( .A(n685), .B(n686), .Z(n682) );
  AND U686 ( .A(n15), .B(n687), .Z(n686) );
  XNOR U687 ( .A(p_input[120]), .B(n685), .Z(n687) );
  XOR U688 ( .A(n688), .B(n689), .Z(n685) );
  AND U689 ( .A(n19), .B(n690), .Z(n689) );
  XNOR U690 ( .A(p_input[152]), .B(n688), .Z(n690) );
  XOR U691 ( .A(n691), .B(n692), .Z(n688) );
  AND U692 ( .A(n23), .B(n693), .Z(n692) );
  XNOR U693 ( .A(p_input[184]), .B(n691), .Z(n693) );
  XOR U694 ( .A(n694), .B(n695), .Z(n691) );
  AND U695 ( .A(n27), .B(n696), .Z(n695) );
  XNOR U696 ( .A(p_input[216]), .B(n694), .Z(n696) );
  XOR U697 ( .A(n697), .B(n698), .Z(n694) );
  AND U698 ( .A(n31), .B(n699), .Z(n698) );
  XNOR U699 ( .A(p_input[248]), .B(n697), .Z(n699) );
  XOR U700 ( .A(n700), .B(n701), .Z(n697) );
  AND U701 ( .A(n35), .B(n702), .Z(n701) );
  XNOR U702 ( .A(p_input[280]), .B(n700), .Z(n702) );
  XOR U703 ( .A(n703), .B(n704), .Z(n700) );
  AND U704 ( .A(n39), .B(n705), .Z(n704) );
  XNOR U705 ( .A(p_input[312]), .B(n703), .Z(n705) );
  XOR U706 ( .A(n706), .B(n707), .Z(n703) );
  AND U707 ( .A(n43), .B(n708), .Z(n707) );
  XNOR U708 ( .A(p_input[344]), .B(n706), .Z(n708) );
  XOR U709 ( .A(n709), .B(n710), .Z(n706) );
  AND U710 ( .A(n47), .B(n711), .Z(n710) );
  XNOR U711 ( .A(p_input[376]), .B(n709), .Z(n711) );
  XOR U712 ( .A(n712), .B(n713), .Z(n709) );
  AND U713 ( .A(n51), .B(n714), .Z(n713) );
  XNOR U714 ( .A(p_input[408]), .B(n712), .Z(n714) );
  XNOR U715 ( .A(n715), .B(n716), .Z(n712) );
  AND U716 ( .A(n55), .B(n717), .Z(n716) );
  XOR U717 ( .A(p_input[440]), .B(n715), .Z(n717) );
  XOR U718 ( .A(\knn_comb_/min_val_out[0][24] ), .B(n718), .Z(n715) );
  AND U719 ( .A(n58), .B(n719), .Z(n718) );
  XOR U720 ( .A(p_input[472]), .B(\knn_comb_/min_val_out[0][24] ), .Z(n719) );
  XNOR U721 ( .A(n720), .B(n721), .Z(o[23]) );
  AND U722 ( .A(n3), .B(n722), .Z(n720) );
  XNOR U723 ( .A(p_input[23]), .B(n721), .Z(n722) );
  XOR U724 ( .A(n723), .B(n724), .Z(n721) );
  AND U725 ( .A(n7), .B(n725), .Z(n724) );
  XNOR U726 ( .A(p_input[55]), .B(n723), .Z(n725) );
  XOR U727 ( .A(n726), .B(n727), .Z(n723) );
  AND U728 ( .A(n11), .B(n728), .Z(n727) );
  XNOR U729 ( .A(p_input[87]), .B(n726), .Z(n728) );
  XOR U730 ( .A(n729), .B(n730), .Z(n726) );
  AND U731 ( .A(n15), .B(n731), .Z(n730) );
  XNOR U732 ( .A(p_input[119]), .B(n729), .Z(n731) );
  XOR U733 ( .A(n732), .B(n733), .Z(n729) );
  AND U734 ( .A(n19), .B(n734), .Z(n733) );
  XNOR U735 ( .A(p_input[151]), .B(n732), .Z(n734) );
  XOR U736 ( .A(n735), .B(n736), .Z(n732) );
  AND U737 ( .A(n23), .B(n737), .Z(n736) );
  XNOR U738 ( .A(p_input[183]), .B(n735), .Z(n737) );
  XOR U739 ( .A(n738), .B(n739), .Z(n735) );
  AND U740 ( .A(n27), .B(n740), .Z(n739) );
  XNOR U741 ( .A(p_input[215]), .B(n738), .Z(n740) );
  XOR U742 ( .A(n741), .B(n742), .Z(n738) );
  AND U743 ( .A(n31), .B(n743), .Z(n742) );
  XNOR U744 ( .A(p_input[247]), .B(n741), .Z(n743) );
  XOR U745 ( .A(n744), .B(n745), .Z(n741) );
  AND U746 ( .A(n35), .B(n746), .Z(n745) );
  XNOR U747 ( .A(p_input[279]), .B(n744), .Z(n746) );
  XOR U748 ( .A(n747), .B(n748), .Z(n744) );
  AND U749 ( .A(n39), .B(n749), .Z(n748) );
  XNOR U750 ( .A(p_input[311]), .B(n747), .Z(n749) );
  XOR U751 ( .A(n750), .B(n751), .Z(n747) );
  AND U752 ( .A(n43), .B(n752), .Z(n751) );
  XNOR U753 ( .A(p_input[343]), .B(n750), .Z(n752) );
  XOR U754 ( .A(n753), .B(n754), .Z(n750) );
  AND U755 ( .A(n47), .B(n755), .Z(n754) );
  XNOR U756 ( .A(p_input[375]), .B(n753), .Z(n755) );
  XOR U757 ( .A(n756), .B(n757), .Z(n753) );
  AND U758 ( .A(n51), .B(n758), .Z(n757) );
  XNOR U759 ( .A(p_input[407]), .B(n756), .Z(n758) );
  XNOR U760 ( .A(n759), .B(n760), .Z(n756) );
  AND U761 ( .A(n55), .B(n761), .Z(n760) );
  XOR U762 ( .A(p_input[439]), .B(n759), .Z(n761) );
  XOR U763 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n762), .Z(n759) );
  AND U764 ( .A(n58), .B(n763), .Z(n762) );
  XOR U765 ( .A(p_input[471]), .B(\knn_comb_/min_val_out[0][23] ), .Z(n763) );
  XNOR U766 ( .A(n764), .B(n765), .Z(o[22]) );
  AND U767 ( .A(n3), .B(n766), .Z(n764) );
  XNOR U768 ( .A(p_input[22]), .B(n765), .Z(n766) );
  XOR U769 ( .A(n767), .B(n768), .Z(n765) );
  AND U770 ( .A(n7), .B(n769), .Z(n768) );
  XNOR U771 ( .A(p_input[54]), .B(n767), .Z(n769) );
  XOR U772 ( .A(n770), .B(n771), .Z(n767) );
  AND U773 ( .A(n11), .B(n772), .Z(n771) );
  XNOR U774 ( .A(p_input[86]), .B(n770), .Z(n772) );
  XOR U775 ( .A(n773), .B(n774), .Z(n770) );
  AND U776 ( .A(n15), .B(n775), .Z(n774) );
  XNOR U777 ( .A(p_input[118]), .B(n773), .Z(n775) );
  XOR U778 ( .A(n776), .B(n777), .Z(n773) );
  AND U779 ( .A(n19), .B(n778), .Z(n777) );
  XNOR U780 ( .A(p_input[150]), .B(n776), .Z(n778) );
  XOR U781 ( .A(n779), .B(n780), .Z(n776) );
  AND U782 ( .A(n23), .B(n781), .Z(n780) );
  XNOR U783 ( .A(p_input[182]), .B(n779), .Z(n781) );
  XOR U784 ( .A(n782), .B(n783), .Z(n779) );
  AND U785 ( .A(n27), .B(n784), .Z(n783) );
  XNOR U786 ( .A(p_input[214]), .B(n782), .Z(n784) );
  XOR U787 ( .A(n785), .B(n786), .Z(n782) );
  AND U788 ( .A(n31), .B(n787), .Z(n786) );
  XNOR U789 ( .A(p_input[246]), .B(n785), .Z(n787) );
  XOR U790 ( .A(n788), .B(n789), .Z(n785) );
  AND U791 ( .A(n35), .B(n790), .Z(n789) );
  XNOR U792 ( .A(p_input[278]), .B(n788), .Z(n790) );
  XOR U793 ( .A(n791), .B(n792), .Z(n788) );
  AND U794 ( .A(n39), .B(n793), .Z(n792) );
  XNOR U795 ( .A(p_input[310]), .B(n791), .Z(n793) );
  XOR U796 ( .A(n794), .B(n795), .Z(n791) );
  AND U797 ( .A(n43), .B(n796), .Z(n795) );
  XNOR U798 ( .A(p_input[342]), .B(n794), .Z(n796) );
  XOR U799 ( .A(n797), .B(n798), .Z(n794) );
  AND U800 ( .A(n47), .B(n799), .Z(n798) );
  XNOR U801 ( .A(p_input[374]), .B(n797), .Z(n799) );
  XOR U802 ( .A(n800), .B(n801), .Z(n797) );
  AND U803 ( .A(n51), .B(n802), .Z(n801) );
  XNOR U804 ( .A(p_input[406]), .B(n800), .Z(n802) );
  XNOR U805 ( .A(n803), .B(n804), .Z(n800) );
  AND U806 ( .A(n55), .B(n805), .Z(n804) );
  XOR U807 ( .A(p_input[438]), .B(n803), .Z(n805) );
  XOR U808 ( .A(\knn_comb_/min_val_out[0][22] ), .B(n806), .Z(n803) );
  AND U809 ( .A(n58), .B(n807), .Z(n806) );
  XOR U810 ( .A(p_input[470]), .B(\knn_comb_/min_val_out[0][22] ), .Z(n807) );
  XNOR U811 ( .A(n808), .B(n809), .Z(o[21]) );
  AND U812 ( .A(n3), .B(n810), .Z(n808) );
  XNOR U813 ( .A(p_input[21]), .B(n809), .Z(n810) );
  XOR U814 ( .A(n811), .B(n812), .Z(n809) );
  AND U815 ( .A(n7), .B(n813), .Z(n812) );
  XNOR U816 ( .A(p_input[53]), .B(n811), .Z(n813) );
  XOR U817 ( .A(n814), .B(n815), .Z(n811) );
  AND U818 ( .A(n11), .B(n816), .Z(n815) );
  XNOR U819 ( .A(p_input[85]), .B(n814), .Z(n816) );
  XOR U820 ( .A(n817), .B(n818), .Z(n814) );
  AND U821 ( .A(n15), .B(n819), .Z(n818) );
  XNOR U822 ( .A(p_input[117]), .B(n817), .Z(n819) );
  XOR U823 ( .A(n820), .B(n821), .Z(n817) );
  AND U824 ( .A(n19), .B(n822), .Z(n821) );
  XNOR U825 ( .A(p_input[149]), .B(n820), .Z(n822) );
  XOR U826 ( .A(n823), .B(n824), .Z(n820) );
  AND U827 ( .A(n23), .B(n825), .Z(n824) );
  XNOR U828 ( .A(p_input[181]), .B(n823), .Z(n825) );
  XOR U829 ( .A(n826), .B(n827), .Z(n823) );
  AND U830 ( .A(n27), .B(n828), .Z(n827) );
  XNOR U831 ( .A(p_input[213]), .B(n826), .Z(n828) );
  XOR U832 ( .A(n829), .B(n830), .Z(n826) );
  AND U833 ( .A(n31), .B(n831), .Z(n830) );
  XNOR U834 ( .A(p_input[245]), .B(n829), .Z(n831) );
  XOR U835 ( .A(n832), .B(n833), .Z(n829) );
  AND U836 ( .A(n35), .B(n834), .Z(n833) );
  XNOR U837 ( .A(p_input[277]), .B(n832), .Z(n834) );
  XOR U838 ( .A(n835), .B(n836), .Z(n832) );
  AND U839 ( .A(n39), .B(n837), .Z(n836) );
  XNOR U840 ( .A(p_input[309]), .B(n835), .Z(n837) );
  XOR U841 ( .A(n838), .B(n839), .Z(n835) );
  AND U842 ( .A(n43), .B(n840), .Z(n839) );
  XNOR U843 ( .A(p_input[341]), .B(n838), .Z(n840) );
  XOR U844 ( .A(n841), .B(n842), .Z(n838) );
  AND U845 ( .A(n47), .B(n843), .Z(n842) );
  XNOR U846 ( .A(p_input[373]), .B(n841), .Z(n843) );
  XOR U847 ( .A(n844), .B(n845), .Z(n841) );
  AND U848 ( .A(n51), .B(n846), .Z(n845) );
  XNOR U849 ( .A(p_input[405]), .B(n844), .Z(n846) );
  XNOR U850 ( .A(n847), .B(n848), .Z(n844) );
  AND U851 ( .A(n55), .B(n849), .Z(n848) );
  XOR U852 ( .A(p_input[437]), .B(n847), .Z(n849) );
  XOR U853 ( .A(\knn_comb_/min_val_out[0][21] ), .B(n850), .Z(n847) );
  AND U854 ( .A(n58), .B(n851), .Z(n850) );
  XOR U855 ( .A(p_input[469]), .B(\knn_comb_/min_val_out[0][21] ), .Z(n851) );
  XNOR U856 ( .A(n852), .B(n853), .Z(o[20]) );
  AND U857 ( .A(n3), .B(n854), .Z(n852) );
  XNOR U858 ( .A(p_input[20]), .B(n853), .Z(n854) );
  XOR U859 ( .A(n855), .B(n856), .Z(n853) );
  AND U860 ( .A(n7), .B(n857), .Z(n856) );
  XNOR U861 ( .A(p_input[52]), .B(n855), .Z(n857) );
  XOR U862 ( .A(n858), .B(n859), .Z(n855) );
  AND U863 ( .A(n11), .B(n860), .Z(n859) );
  XNOR U864 ( .A(p_input[84]), .B(n858), .Z(n860) );
  XOR U865 ( .A(n861), .B(n862), .Z(n858) );
  AND U866 ( .A(n15), .B(n863), .Z(n862) );
  XNOR U867 ( .A(p_input[116]), .B(n861), .Z(n863) );
  XOR U868 ( .A(n864), .B(n865), .Z(n861) );
  AND U869 ( .A(n19), .B(n866), .Z(n865) );
  XNOR U870 ( .A(p_input[148]), .B(n864), .Z(n866) );
  XOR U871 ( .A(n867), .B(n868), .Z(n864) );
  AND U872 ( .A(n23), .B(n869), .Z(n868) );
  XNOR U873 ( .A(p_input[180]), .B(n867), .Z(n869) );
  XOR U874 ( .A(n870), .B(n871), .Z(n867) );
  AND U875 ( .A(n27), .B(n872), .Z(n871) );
  XNOR U876 ( .A(p_input[212]), .B(n870), .Z(n872) );
  XOR U877 ( .A(n873), .B(n874), .Z(n870) );
  AND U878 ( .A(n31), .B(n875), .Z(n874) );
  XNOR U879 ( .A(p_input[244]), .B(n873), .Z(n875) );
  XOR U880 ( .A(n876), .B(n877), .Z(n873) );
  AND U881 ( .A(n35), .B(n878), .Z(n877) );
  XNOR U882 ( .A(p_input[276]), .B(n876), .Z(n878) );
  XOR U883 ( .A(n879), .B(n880), .Z(n876) );
  AND U884 ( .A(n39), .B(n881), .Z(n880) );
  XNOR U885 ( .A(p_input[308]), .B(n879), .Z(n881) );
  XOR U886 ( .A(n882), .B(n883), .Z(n879) );
  AND U887 ( .A(n43), .B(n884), .Z(n883) );
  XNOR U888 ( .A(p_input[340]), .B(n882), .Z(n884) );
  XOR U889 ( .A(n885), .B(n886), .Z(n882) );
  AND U890 ( .A(n47), .B(n887), .Z(n886) );
  XNOR U891 ( .A(p_input[372]), .B(n885), .Z(n887) );
  XOR U892 ( .A(n888), .B(n889), .Z(n885) );
  AND U893 ( .A(n51), .B(n890), .Z(n889) );
  XNOR U894 ( .A(p_input[404]), .B(n888), .Z(n890) );
  XNOR U895 ( .A(n891), .B(n892), .Z(n888) );
  AND U896 ( .A(n55), .B(n893), .Z(n892) );
  XOR U897 ( .A(p_input[436]), .B(n891), .Z(n893) );
  XOR U898 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n894), .Z(n891) );
  AND U899 ( .A(n58), .B(n895), .Z(n894) );
  XOR U900 ( .A(p_input[468]), .B(\knn_comb_/min_val_out[0][20] ), .Z(n895) );
  XNOR U901 ( .A(n896), .B(n897), .Z(o[1]) );
  AND U902 ( .A(n3), .B(n898), .Z(n896) );
  XNOR U903 ( .A(p_input[1]), .B(n897), .Z(n898) );
  XOR U904 ( .A(n899), .B(n900), .Z(n897) );
  AND U905 ( .A(n7), .B(n901), .Z(n900) );
  XNOR U906 ( .A(p_input[33]), .B(n899), .Z(n901) );
  XOR U907 ( .A(n902), .B(n903), .Z(n899) );
  AND U908 ( .A(n11), .B(n904), .Z(n903) );
  XNOR U909 ( .A(p_input[65]), .B(n902), .Z(n904) );
  XOR U910 ( .A(n905), .B(n906), .Z(n902) );
  AND U911 ( .A(n15), .B(n907), .Z(n906) );
  XNOR U912 ( .A(p_input[97]), .B(n905), .Z(n907) );
  XOR U913 ( .A(n908), .B(n909), .Z(n905) );
  AND U914 ( .A(n19), .B(n910), .Z(n909) );
  XNOR U915 ( .A(p_input[129]), .B(n908), .Z(n910) );
  XOR U916 ( .A(n911), .B(n912), .Z(n908) );
  AND U917 ( .A(n23), .B(n913), .Z(n912) );
  XNOR U918 ( .A(p_input[161]), .B(n911), .Z(n913) );
  XOR U919 ( .A(n914), .B(n915), .Z(n911) );
  AND U920 ( .A(n27), .B(n916), .Z(n915) );
  XNOR U921 ( .A(p_input[193]), .B(n914), .Z(n916) );
  XOR U922 ( .A(n917), .B(n918), .Z(n914) );
  AND U923 ( .A(n31), .B(n919), .Z(n918) );
  XNOR U924 ( .A(p_input[225]), .B(n917), .Z(n919) );
  XOR U925 ( .A(n920), .B(n921), .Z(n917) );
  AND U926 ( .A(n35), .B(n922), .Z(n921) );
  XNOR U927 ( .A(p_input[257]), .B(n920), .Z(n922) );
  XOR U928 ( .A(n923), .B(n924), .Z(n920) );
  AND U929 ( .A(n39), .B(n925), .Z(n924) );
  XNOR U930 ( .A(p_input[289]), .B(n923), .Z(n925) );
  XOR U931 ( .A(n926), .B(n927), .Z(n923) );
  AND U932 ( .A(n43), .B(n928), .Z(n927) );
  XNOR U933 ( .A(p_input[321]), .B(n926), .Z(n928) );
  XOR U934 ( .A(n929), .B(n930), .Z(n926) );
  AND U935 ( .A(n47), .B(n931), .Z(n930) );
  XNOR U936 ( .A(p_input[353]), .B(n929), .Z(n931) );
  XOR U937 ( .A(n932), .B(n933), .Z(n929) );
  AND U938 ( .A(n51), .B(n934), .Z(n933) );
  XNOR U939 ( .A(p_input[385]), .B(n932), .Z(n934) );
  XNOR U940 ( .A(n935), .B(n936), .Z(n932) );
  AND U941 ( .A(n55), .B(n937), .Z(n936) );
  XOR U942 ( .A(p_input[417]), .B(n935), .Z(n937) );
  XOR U943 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n938), .Z(n935) );
  AND U944 ( .A(n58), .B(n939), .Z(n938) );
  XOR U945 ( .A(p_input[449]), .B(\knn_comb_/min_val_out[0][1] ), .Z(n939) );
  XNOR U946 ( .A(n940), .B(n941), .Z(o[19]) );
  AND U947 ( .A(n3), .B(n942), .Z(n940) );
  XNOR U948 ( .A(p_input[19]), .B(n941), .Z(n942) );
  XOR U949 ( .A(n943), .B(n944), .Z(n941) );
  AND U950 ( .A(n7), .B(n945), .Z(n944) );
  XNOR U951 ( .A(p_input[51]), .B(n943), .Z(n945) );
  XOR U952 ( .A(n946), .B(n947), .Z(n943) );
  AND U953 ( .A(n11), .B(n948), .Z(n947) );
  XNOR U954 ( .A(p_input[83]), .B(n946), .Z(n948) );
  XOR U955 ( .A(n949), .B(n950), .Z(n946) );
  AND U956 ( .A(n15), .B(n951), .Z(n950) );
  XNOR U957 ( .A(p_input[115]), .B(n949), .Z(n951) );
  XOR U958 ( .A(n952), .B(n953), .Z(n949) );
  AND U959 ( .A(n19), .B(n954), .Z(n953) );
  XNOR U960 ( .A(p_input[147]), .B(n952), .Z(n954) );
  XOR U961 ( .A(n955), .B(n956), .Z(n952) );
  AND U962 ( .A(n23), .B(n957), .Z(n956) );
  XNOR U963 ( .A(p_input[179]), .B(n955), .Z(n957) );
  XOR U964 ( .A(n958), .B(n959), .Z(n955) );
  AND U965 ( .A(n27), .B(n960), .Z(n959) );
  XNOR U966 ( .A(p_input[211]), .B(n958), .Z(n960) );
  XOR U967 ( .A(n961), .B(n962), .Z(n958) );
  AND U968 ( .A(n31), .B(n963), .Z(n962) );
  XNOR U969 ( .A(p_input[243]), .B(n961), .Z(n963) );
  XOR U970 ( .A(n964), .B(n965), .Z(n961) );
  AND U971 ( .A(n35), .B(n966), .Z(n965) );
  XNOR U972 ( .A(p_input[275]), .B(n964), .Z(n966) );
  XOR U973 ( .A(n967), .B(n968), .Z(n964) );
  AND U974 ( .A(n39), .B(n969), .Z(n968) );
  XNOR U975 ( .A(p_input[307]), .B(n967), .Z(n969) );
  XOR U976 ( .A(n970), .B(n971), .Z(n967) );
  AND U977 ( .A(n43), .B(n972), .Z(n971) );
  XNOR U978 ( .A(p_input[339]), .B(n970), .Z(n972) );
  XOR U979 ( .A(n973), .B(n974), .Z(n970) );
  AND U980 ( .A(n47), .B(n975), .Z(n974) );
  XNOR U981 ( .A(p_input[371]), .B(n973), .Z(n975) );
  XOR U982 ( .A(n976), .B(n977), .Z(n973) );
  AND U983 ( .A(n51), .B(n978), .Z(n977) );
  XNOR U984 ( .A(p_input[403]), .B(n976), .Z(n978) );
  XNOR U985 ( .A(n979), .B(n980), .Z(n976) );
  AND U986 ( .A(n55), .B(n981), .Z(n980) );
  XOR U987 ( .A(p_input[435]), .B(n979), .Z(n981) );
  XOR U988 ( .A(\knn_comb_/min_val_out[0][19] ), .B(n982), .Z(n979) );
  AND U989 ( .A(n58), .B(n983), .Z(n982) );
  XOR U990 ( .A(p_input[467]), .B(\knn_comb_/min_val_out[0][19] ), .Z(n983) );
  XNOR U991 ( .A(n984), .B(n985), .Z(o[18]) );
  AND U992 ( .A(n3), .B(n986), .Z(n984) );
  XNOR U993 ( .A(p_input[18]), .B(n985), .Z(n986) );
  XOR U994 ( .A(n987), .B(n988), .Z(n985) );
  AND U995 ( .A(n7), .B(n989), .Z(n988) );
  XNOR U996 ( .A(p_input[50]), .B(n987), .Z(n989) );
  XOR U997 ( .A(n990), .B(n991), .Z(n987) );
  AND U998 ( .A(n11), .B(n992), .Z(n991) );
  XNOR U999 ( .A(p_input[82]), .B(n990), .Z(n992) );
  XOR U1000 ( .A(n993), .B(n994), .Z(n990) );
  AND U1001 ( .A(n15), .B(n995), .Z(n994) );
  XNOR U1002 ( .A(p_input[114]), .B(n993), .Z(n995) );
  XOR U1003 ( .A(n996), .B(n997), .Z(n993) );
  AND U1004 ( .A(n19), .B(n998), .Z(n997) );
  XNOR U1005 ( .A(p_input[146]), .B(n996), .Z(n998) );
  XOR U1006 ( .A(n999), .B(n1000), .Z(n996) );
  AND U1007 ( .A(n23), .B(n1001), .Z(n1000) );
  XNOR U1008 ( .A(p_input[178]), .B(n999), .Z(n1001) );
  XOR U1009 ( .A(n1002), .B(n1003), .Z(n999) );
  AND U1010 ( .A(n27), .B(n1004), .Z(n1003) );
  XNOR U1011 ( .A(p_input[210]), .B(n1002), .Z(n1004) );
  XOR U1012 ( .A(n1005), .B(n1006), .Z(n1002) );
  AND U1013 ( .A(n31), .B(n1007), .Z(n1006) );
  XNOR U1014 ( .A(p_input[242]), .B(n1005), .Z(n1007) );
  XOR U1015 ( .A(n1008), .B(n1009), .Z(n1005) );
  AND U1016 ( .A(n35), .B(n1010), .Z(n1009) );
  XNOR U1017 ( .A(p_input[274]), .B(n1008), .Z(n1010) );
  XOR U1018 ( .A(n1011), .B(n1012), .Z(n1008) );
  AND U1019 ( .A(n39), .B(n1013), .Z(n1012) );
  XNOR U1020 ( .A(p_input[306]), .B(n1011), .Z(n1013) );
  XOR U1021 ( .A(n1014), .B(n1015), .Z(n1011) );
  AND U1022 ( .A(n43), .B(n1016), .Z(n1015) );
  XNOR U1023 ( .A(p_input[338]), .B(n1014), .Z(n1016) );
  XOR U1024 ( .A(n1017), .B(n1018), .Z(n1014) );
  AND U1025 ( .A(n47), .B(n1019), .Z(n1018) );
  XNOR U1026 ( .A(p_input[370]), .B(n1017), .Z(n1019) );
  XOR U1027 ( .A(n1020), .B(n1021), .Z(n1017) );
  AND U1028 ( .A(n51), .B(n1022), .Z(n1021) );
  XNOR U1029 ( .A(p_input[402]), .B(n1020), .Z(n1022) );
  XNOR U1030 ( .A(n1023), .B(n1024), .Z(n1020) );
  AND U1031 ( .A(n55), .B(n1025), .Z(n1024) );
  XOR U1032 ( .A(p_input[434]), .B(n1023), .Z(n1025) );
  XOR U1033 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n1026), .Z(n1023) );
  AND U1034 ( .A(n58), .B(n1027), .Z(n1026) );
  XOR U1035 ( .A(p_input[466]), .B(\knn_comb_/min_val_out[0][18] ), .Z(n1027)
         );
  XNOR U1036 ( .A(n1028), .B(n1029), .Z(o[17]) );
  AND U1037 ( .A(n3), .B(n1030), .Z(n1028) );
  XNOR U1038 ( .A(p_input[17]), .B(n1029), .Z(n1030) );
  XOR U1039 ( .A(n1031), .B(n1032), .Z(n1029) );
  AND U1040 ( .A(n7), .B(n1033), .Z(n1032) );
  XNOR U1041 ( .A(p_input[49]), .B(n1031), .Z(n1033) );
  XOR U1042 ( .A(n1034), .B(n1035), .Z(n1031) );
  AND U1043 ( .A(n11), .B(n1036), .Z(n1035) );
  XNOR U1044 ( .A(p_input[81]), .B(n1034), .Z(n1036) );
  XOR U1045 ( .A(n1037), .B(n1038), .Z(n1034) );
  AND U1046 ( .A(n15), .B(n1039), .Z(n1038) );
  XNOR U1047 ( .A(p_input[113]), .B(n1037), .Z(n1039) );
  XOR U1048 ( .A(n1040), .B(n1041), .Z(n1037) );
  AND U1049 ( .A(n19), .B(n1042), .Z(n1041) );
  XNOR U1050 ( .A(p_input[145]), .B(n1040), .Z(n1042) );
  XOR U1051 ( .A(n1043), .B(n1044), .Z(n1040) );
  AND U1052 ( .A(n23), .B(n1045), .Z(n1044) );
  XNOR U1053 ( .A(p_input[177]), .B(n1043), .Z(n1045) );
  XOR U1054 ( .A(n1046), .B(n1047), .Z(n1043) );
  AND U1055 ( .A(n27), .B(n1048), .Z(n1047) );
  XNOR U1056 ( .A(p_input[209]), .B(n1046), .Z(n1048) );
  XOR U1057 ( .A(n1049), .B(n1050), .Z(n1046) );
  AND U1058 ( .A(n31), .B(n1051), .Z(n1050) );
  XNOR U1059 ( .A(p_input[241]), .B(n1049), .Z(n1051) );
  XOR U1060 ( .A(n1052), .B(n1053), .Z(n1049) );
  AND U1061 ( .A(n35), .B(n1054), .Z(n1053) );
  XNOR U1062 ( .A(p_input[273]), .B(n1052), .Z(n1054) );
  XOR U1063 ( .A(n1055), .B(n1056), .Z(n1052) );
  AND U1064 ( .A(n39), .B(n1057), .Z(n1056) );
  XNOR U1065 ( .A(p_input[305]), .B(n1055), .Z(n1057) );
  XOR U1066 ( .A(n1058), .B(n1059), .Z(n1055) );
  AND U1067 ( .A(n43), .B(n1060), .Z(n1059) );
  XNOR U1068 ( .A(p_input[337]), .B(n1058), .Z(n1060) );
  XOR U1069 ( .A(n1061), .B(n1062), .Z(n1058) );
  AND U1070 ( .A(n47), .B(n1063), .Z(n1062) );
  XNOR U1071 ( .A(p_input[369]), .B(n1061), .Z(n1063) );
  XOR U1072 ( .A(n1064), .B(n1065), .Z(n1061) );
  AND U1073 ( .A(n51), .B(n1066), .Z(n1065) );
  XNOR U1074 ( .A(p_input[401]), .B(n1064), .Z(n1066) );
  XNOR U1075 ( .A(n1067), .B(n1068), .Z(n1064) );
  AND U1076 ( .A(n55), .B(n1069), .Z(n1068) );
  XOR U1077 ( .A(p_input[433]), .B(n1067), .Z(n1069) );
  XOR U1078 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n1070), .Z(n1067) );
  AND U1079 ( .A(n58), .B(n1071), .Z(n1070) );
  XOR U1080 ( .A(p_input[465]), .B(\knn_comb_/min_val_out[0][17] ), .Z(n1071)
         );
  XNOR U1081 ( .A(n1072), .B(n1073), .Z(o[16]) );
  AND U1082 ( .A(n3), .B(n1074), .Z(n1072) );
  XNOR U1083 ( .A(p_input[16]), .B(n1073), .Z(n1074) );
  XOR U1084 ( .A(n1075), .B(n1076), .Z(n1073) );
  AND U1085 ( .A(n7), .B(n1077), .Z(n1076) );
  XNOR U1086 ( .A(p_input[48]), .B(n1075), .Z(n1077) );
  XOR U1087 ( .A(n1078), .B(n1079), .Z(n1075) );
  AND U1088 ( .A(n11), .B(n1080), .Z(n1079) );
  XNOR U1089 ( .A(p_input[80]), .B(n1078), .Z(n1080) );
  XOR U1090 ( .A(n1081), .B(n1082), .Z(n1078) );
  AND U1091 ( .A(n15), .B(n1083), .Z(n1082) );
  XNOR U1092 ( .A(p_input[112]), .B(n1081), .Z(n1083) );
  XOR U1093 ( .A(n1084), .B(n1085), .Z(n1081) );
  AND U1094 ( .A(n19), .B(n1086), .Z(n1085) );
  XNOR U1095 ( .A(p_input[144]), .B(n1084), .Z(n1086) );
  XOR U1096 ( .A(n1087), .B(n1088), .Z(n1084) );
  AND U1097 ( .A(n23), .B(n1089), .Z(n1088) );
  XNOR U1098 ( .A(p_input[176]), .B(n1087), .Z(n1089) );
  XOR U1099 ( .A(n1090), .B(n1091), .Z(n1087) );
  AND U1100 ( .A(n27), .B(n1092), .Z(n1091) );
  XNOR U1101 ( .A(p_input[208]), .B(n1090), .Z(n1092) );
  XOR U1102 ( .A(n1093), .B(n1094), .Z(n1090) );
  AND U1103 ( .A(n31), .B(n1095), .Z(n1094) );
  XNOR U1104 ( .A(p_input[240]), .B(n1093), .Z(n1095) );
  XOR U1105 ( .A(n1096), .B(n1097), .Z(n1093) );
  AND U1106 ( .A(n35), .B(n1098), .Z(n1097) );
  XNOR U1107 ( .A(p_input[272]), .B(n1096), .Z(n1098) );
  XOR U1108 ( .A(n1099), .B(n1100), .Z(n1096) );
  AND U1109 ( .A(n39), .B(n1101), .Z(n1100) );
  XNOR U1110 ( .A(p_input[304]), .B(n1099), .Z(n1101) );
  XOR U1111 ( .A(n1102), .B(n1103), .Z(n1099) );
  AND U1112 ( .A(n43), .B(n1104), .Z(n1103) );
  XNOR U1113 ( .A(p_input[336]), .B(n1102), .Z(n1104) );
  XOR U1114 ( .A(n1105), .B(n1106), .Z(n1102) );
  AND U1115 ( .A(n47), .B(n1107), .Z(n1106) );
  XNOR U1116 ( .A(p_input[368]), .B(n1105), .Z(n1107) );
  XOR U1117 ( .A(n1108), .B(n1109), .Z(n1105) );
  AND U1118 ( .A(n51), .B(n1110), .Z(n1109) );
  XNOR U1119 ( .A(p_input[400]), .B(n1108), .Z(n1110) );
  XNOR U1120 ( .A(n1111), .B(n1112), .Z(n1108) );
  AND U1121 ( .A(n55), .B(n1113), .Z(n1112) );
  XOR U1122 ( .A(p_input[432]), .B(n1111), .Z(n1113) );
  XOR U1123 ( .A(\knn_comb_/min_val_out[0][16] ), .B(n1114), .Z(n1111) );
  AND U1124 ( .A(n58), .B(n1115), .Z(n1114) );
  XOR U1125 ( .A(p_input[464]), .B(\knn_comb_/min_val_out[0][16] ), .Z(n1115)
         );
  XNOR U1126 ( .A(n1116), .B(n1117), .Z(o[15]) );
  AND U1127 ( .A(n3), .B(n1118), .Z(n1116) );
  XNOR U1128 ( .A(p_input[15]), .B(n1117), .Z(n1118) );
  XOR U1129 ( .A(n1119), .B(n1120), .Z(n1117) );
  AND U1130 ( .A(n7), .B(n1121), .Z(n1120) );
  XNOR U1131 ( .A(p_input[47]), .B(n1119), .Z(n1121) );
  XOR U1132 ( .A(n1122), .B(n1123), .Z(n1119) );
  AND U1133 ( .A(n11), .B(n1124), .Z(n1123) );
  XNOR U1134 ( .A(p_input[79]), .B(n1122), .Z(n1124) );
  XOR U1135 ( .A(n1125), .B(n1126), .Z(n1122) );
  AND U1136 ( .A(n15), .B(n1127), .Z(n1126) );
  XNOR U1137 ( .A(p_input[111]), .B(n1125), .Z(n1127) );
  XOR U1138 ( .A(n1128), .B(n1129), .Z(n1125) );
  AND U1139 ( .A(n19), .B(n1130), .Z(n1129) );
  XNOR U1140 ( .A(p_input[143]), .B(n1128), .Z(n1130) );
  XOR U1141 ( .A(n1131), .B(n1132), .Z(n1128) );
  AND U1142 ( .A(n23), .B(n1133), .Z(n1132) );
  XNOR U1143 ( .A(p_input[175]), .B(n1131), .Z(n1133) );
  XOR U1144 ( .A(n1134), .B(n1135), .Z(n1131) );
  AND U1145 ( .A(n27), .B(n1136), .Z(n1135) );
  XNOR U1146 ( .A(p_input[207]), .B(n1134), .Z(n1136) );
  XOR U1147 ( .A(n1137), .B(n1138), .Z(n1134) );
  AND U1148 ( .A(n31), .B(n1139), .Z(n1138) );
  XNOR U1149 ( .A(p_input[239]), .B(n1137), .Z(n1139) );
  XOR U1150 ( .A(n1140), .B(n1141), .Z(n1137) );
  AND U1151 ( .A(n35), .B(n1142), .Z(n1141) );
  XNOR U1152 ( .A(p_input[271]), .B(n1140), .Z(n1142) );
  XOR U1153 ( .A(n1143), .B(n1144), .Z(n1140) );
  AND U1154 ( .A(n39), .B(n1145), .Z(n1144) );
  XNOR U1155 ( .A(p_input[303]), .B(n1143), .Z(n1145) );
  XOR U1156 ( .A(n1146), .B(n1147), .Z(n1143) );
  AND U1157 ( .A(n43), .B(n1148), .Z(n1147) );
  XNOR U1158 ( .A(p_input[335]), .B(n1146), .Z(n1148) );
  XOR U1159 ( .A(n1149), .B(n1150), .Z(n1146) );
  AND U1160 ( .A(n47), .B(n1151), .Z(n1150) );
  XNOR U1161 ( .A(p_input[367]), .B(n1149), .Z(n1151) );
  XOR U1162 ( .A(n1152), .B(n1153), .Z(n1149) );
  AND U1163 ( .A(n51), .B(n1154), .Z(n1153) );
  XNOR U1164 ( .A(p_input[399]), .B(n1152), .Z(n1154) );
  XNOR U1165 ( .A(n1155), .B(n1156), .Z(n1152) );
  AND U1166 ( .A(n55), .B(n1157), .Z(n1156) );
  XOR U1167 ( .A(p_input[431]), .B(n1155), .Z(n1157) );
  XOR U1168 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n1158), .Z(n1155) );
  AND U1169 ( .A(n58), .B(n1159), .Z(n1158) );
  XOR U1170 ( .A(p_input[463]), .B(\knn_comb_/min_val_out[0][15] ), .Z(n1159)
         );
  XNOR U1171 ( .A(n1160), .B(n1161), .Z(o[14]) );
  AND U1172 ( .A(n3), .B(n1162), .Z(n1160) );
  XNOR U1173 ( .A(p_input[14]), .B(n1161), .Z(n1162) );
  XOR U1174 ( .A(n1163), .B(n1164), .Z(n1161) );
  AND U1175 ( .A(n7), .B(n1165), .Z(n1164) );
  XNOR U1176 ( .A(p_input[46]), .B(n1163), .Z(n1165) );
  XOR U1177 ( .A(n1166), .B(n1167), .Z(n1163) );
  AND U1178 ( .A(n11), .B(n1168), .Z(n1167) );
  XNOR U1179 ( .A(p_input[78]), .B(n1166), .Z(n1168) );
  XOR U1180 ( .A(n1169), .B(n1170), .Z(n1166) );
  AND U1181 ( .A(n15), .B(n1171), .Z(n1170) );
  XNOR U1182 ( .A(p_input[110]), .B(n1169), .Z(n1171) );
  XOR U1183 ( .A(n1172), .B(n1173), .Z(n1169) );
  AND U1184 ( .A(n19), .B(n1174), .Z(n1173) );
  XNOR U1185 ( .A(p_input[142]), .B(n1172), .Z(n1174) );
  XOR U1186 ( .A(n1175), .B(n1176), .Z(n1172) );
  AND U1187 ( .A(n23), .B(n1177), .Z(n1176) );
  XNOR U1188 ( .A(p_input[174]), .B(n1175), .Z(n1177) );
  XOR U1189 ( .A(n1178), .B(n1179), .Z(n1175) );
  AND U1190 ( .A(n27), .B(n1180), .Z(n1179) );
  XNOR U1191 ( .A(p_input[206]), .B(n1178), .Z(n1180) );
  XOR U1192 ( .A(n1181), .B(n1182), .Z(n1178) );
  AND U1193 ( .A(n31), .B(n1183), .Z(n1182) );
  XNOR U1194 ( .A(p_input[238]), .B(n1181), .Z(n1183) );
  XOR U1195 ( .A(n1184), .B(n1185), .Z(n1181) );
  AND U1196 ( .A(n35), .B(n1186), .Z(n1185) );
  XNOR U1197 ( .A(p_input[270]), .B(n1184), .Z(n1186) );
  XOR U1198 ( .A(n1187), .B(n1188), .Z(n1184) );
  AND U1199 ( .A(n39), .B(n1189), .Z(n1188) );
  XNOR U1200 ( .A(p_input[302]), .B(n1187), .Z(n1189) );
  XOR U1201 ( .A(n1190), .B(n1191), .Z(n1187) );
  AND U1202 ( .A(n43), .B(n1192), .Z(n1191) );
  XNOR U1203 ( .A(p_input[334]), .B(n1190), .Z(n1192) );
  XOR U1204 ( .A(n1193), .B(n1194), .Z(n1190) );
  AND U1205 ( .A(n47), .B(n1195), .Z(n1194) );
  XNOR U1206 ( .A(p_input[366]), .B(n1193), .Z(n1195) );
  XOR U1207 ( .A(n1196), .B(n1197), .Z(n1193) );
  AND U1208 ( .A(n51), .B(n1198), .Z(n1197) );
  XNOR U1209 ( .A(p_input[398]), .B(n1196), .Z(n1198) );
  XNOR U1210 ( .A(n1199), .B(n1200), .Z(n1196) );
  AND U1211 ( .A(n55), .B(n1201), .Z(n1200) );
  XOR U1212 ( .A(p_input[430]), .B(n1199), .Z(n1201) );
  XOR U1213 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n1202), .Z(n1199) );
  AND U1214 ( .A(n58), .B(n1203), .Z(n1202) );
  XOR U1215 ( .A(p_input[462]), .B(\knn_comb_/min_val_out[0][14] ), .Z(n1203)
         );
  XNOR U1216 ( .A(n1204), .B(n1205), .Z(o[13]) );
  AND U1217 ( .A(n3), .B(n1206), .Z(n1204) );
  XNOR U1218 ( .A(p_input[13]), .B(n1205), .Z(n1206) );
  XOR U1219 ( .A(n1207), .B(n1208), .Z(n1205) );
  AND U1220 ( .A(n7), .B(n1209), .Z(n1208) );
  XNOR U1221 ( .A(p_input[45]), .B(n1207), .Z(n1209) );
  XOR U1222 ( .A(n1210), .B(n1211), .Z(n1207) );
  AND U1223 ( .A(n11), .B(n1212), .Z(n1211) );
  XNOR U1224 ( .A(p_input[77]), .B(n1210), .Z(n1212) );
  XOR U1225 ( .A(n1213), .B(n1214), .Z(n1210) );
  AND U1226 ( .A(n15), .B(n1215), .Z(n1214) );
  XNOR U1227 ( .A(p_input[109]), .B(n1213), .Z(n1215) );
  XOR U1228 ( .A(n1216), .B(n1217), .Z(n1213) );
  AND U1229 ( .A(n19), .B(n1218), .Z(n1217) );
  XNOR U1230 ( .A(p_input[141]), .B(n1216), .Z(n1218) );
  XOR U1231 ( .A(n1219), .B(n1220), .Z(n1216) );
  AND U1232 ( .A(n23), .B(n1221), .Z(n1220) );
  XNOR U1233 ( .A(p_input[173]), .B(n1219), .Z(n1221) );
  XOR U1234 ( .A(n1222), .B(n1223), .Z(n1219) );
  AND U1235 ( .A(n27), .B(n1224), .Z(n1223) );
  XNOR U1236 ( .A(p_input[205]), .B(n1222), .Z(n1224) );
  XOR U1237 ( .A(n1225), .B(n1226), .Z(n1222) );
  AND U1238 ( .A(n31), .B(n1227), .Z(n1226) );
  XNOR U1239 ( .A(p_input[237]), .B(n1225), .Z(n1227) );
  XOR U1240 ( .A(n1228), .B(n1229), .Z(n1225) );
  AND U1241 ( .A(n35), .B(n1230), .Z(n1229) );
  XNOR U1242 ( .A(p_input[269]), .B(n1228), .Z(n1230) );
  XOR U1243 ( .A(n1231), .B(n1232), .Z(n1228) );
  AND U1244 ( .A(n39), .B(n1233), .Z(n1232) );
  XNOR U1245 ( .A(p_input[301]), .B(n1231), .Z(n1233) );
  XOR U1246 ( .A(n1234), .B(n1235), .Z(n1231) );
  AND U1247 ( .A(n43), .B(n1236), .Z(n1235) );
  XNOR U1248 ( .A(p_input[333]), .B(n1234), .Z(n1236) );
  XOR U1249 ( .A(n1237), .B(n1238), .Z(n1234) );
  AND U1250 ( .A(n47), .B(n1239), .Z(n1238) );
  XNOR U1251 ( .A(p_input[365]), .B(n1237), .Z(n1239) );
  XOR U1252 ( .A(n1240), .B(n1241), .Z(n1237) );
  AND U1253 ( .A(n51), .B(n1242), .Z(n1241) );
  XNOR U1254 ( .A(p_input[397]), .B(n1240), .Z(n1242) );
  XNOR U1255 ( .A(n1243), .B(n1244), .Z(n1240) );
  AND U1256 ( .A(n55), .B(n1245), .Z(n1244) );
  XOR U1257 ( .A(p_input[429]), .B(n1243), .Z(n1245) );
  XOR U1258 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n1246), .Z(n1243) );
  AND U1259 ( .A(n58), .B(n1247), .Z(n1246) );
  XOR U1260 ( .A(p_input[461]), .B(\knn_comb_/min_val_out[0][13] ), .Z(n1247)
         );
  XNOR U1261 ( .A(n1248), .B(n1249), .Z(o[12]) );
  AND U1262 ( .A(n3), .B(n1250), .Z(n1248) );
  XNOR U1263 ( .A(p_input[12]), .B(n1249), .Z(n1250) );
  XOR U1264 ( .A(n1251), .B(n1252), .Z(n1249) );
  AND U1265 ( .A(n7), .B(n1253), .Z(n1252) );
  XNOR U1266 ( .A(p_input[44]), .B(n1251), .Z(n1253) );
  XOR U1267 ( .A(n1254), .B(n1255), .Z(n1251) );
  AND U1268 ( .A(n11), .B(n1256), .Z(n1255) );
  XNOR U1269 ( .A(p_input[76]), .B(n1254), .Z(n1256) );
  XOR U1270 ( .A(n1257), .B(n1258), .Z(n1254) );
  AND U1271 ( .A(n15), .B(n1259), .Z(n1258) );
  XNOR U1272 ( .A(p_input[108]), .B(n1257), .Z(n1259) );
  XOR U1273 ( .A(n1260), .B(n1261), .Z(n1257) );
  AND U1274 ( .A(n19), .B(n1262), .Z(n1261) );
  XNOR U1275 ( .A(p_input[140]), .B(n1260), .Z(n1262) );
  XOR U1276 ( .A(n1263), .B(n1264), .Z(n1260) );
  AND U1277 ( .A(n23), .B(n1265), .Z(n1264) );
  XNOR U1278 ( .A(p_input[172]), .B(n1263), .Z(n1265) );
  XOR U1279 ( .A(n1266), .B(n1267), .Z(n1263) );
  AND U1280 ( .A(n27), .B(n1268), .Z(n1267) );
  XNOR U1281 ( .A(p_input[204]), .B(n1266), .Z(n1268) );
  XOR U1282 ( .A(n1269), .B(n1270), .Z(n1266) );
  AND U1283 ( .A(n31), .B(n1271), .Z(n1270) );
  XNOR U1284 ( .A(p_input[236]), .B(n1269), .Z(n1271) );
  XOR U1285 ( .A(n1272), .B(n1273), .Z(n1269) );
  AND U1286 ( .A(n35), .B(n1274), .Z(n1273) );
  XNOR U1287 ( .A(p_input[268]), .B(n1272), .Z(n1274) );
  XOR U1288 ( .A(n1275), .B(n1276), .Z(n1272) );
  AND U1289 ( .A(n39), .B(n1277), .Z(n1276) );
  XNOR U1290 ( .A(p_input[300]), .B(n1275), .Z(n1277) );
  XOR U1291 ( .A(n1278), .B(n1279), .Z(n1275) );
  AND U1292 ( .A(n43), .B(n1280), .Z(n1279) );
  XNOR U1293 ( .A(p_input[332]), .B(n1278), .Z(n1280) );
  XOR U1294 ( .A(n1281), .B(n1282), .Z(n1278) );
  AND U1295 ( .A(n47), .B(n1283), .Z(n1282) );
  XNOR U1296 ( .A(p_input[364]), .B(n1281), .Z(n1283) );
  XOR U1297 ( .A(n1284), .B(n1285), .Z(n1281) );
  AND U1298 ( .A(n51), .B(n1286), .Z(n1285) );
  XNOR U1299 ( .A(p_input[396]), .B(n1284), .Z(n1286) );
  XNOR U1300 ( .A(n1287), .B(n1288), .Z(n1284) );
  AND U1301 ( .A(n55), .B(n1289), .Z(n1288) );
  XOR U1302 ( .A(p_input[428]), .B(n1287), .Z(n1289) );
  XOR U1303 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n1290), .Z(n1287) );
  AND U1304 ( .A(n58), .B(n1291), .Z(n1290) );
  XOR U1305 ( .A(p_input[460]), .B(\knn_comb_/min_val_out[0][12] ), .Z(n1291)
         );
  XNOR U1306 ( .A(n1292), .B(n1293), .Z(o[11]) );
  AND U1307 ( .A(n3), .B(n1294), .Z(n1292) );
  XNOR U1308 ( .A(p_input[11]), .B(n1293), .Z(n1294) );
  XOR U1309 ( .A(n1295), .B(n1296), .Z(n1293) );
  AND U1310 ( .A(n7), .B(n1297), .Z(n1296) );
  XNOR U1311 ( .A(p_input[43]), .B(n1295), .Z(n1297) );
  XOR U1312 ( .A(n1298), .B(n1299), .Z(n1295) );
  AND U1313 ( .A(n11), .B(n1300), .Z(n1299) );
  XNOR U1314 ( .A(p_input[75]), .B(n1298), .Z(n1300) );
  XOR U1315 ( .A(n1301), .B(n1302), .Z(n1298) );
  AND U1316 ( .A(n15), .B(n1303), .Z(n1302) );
  XNOR U1317 ( .A(p_input[107]), .B(n1301), .Z(n1303) );
  XOR U1318 ( .A(n1304), .B(n1305), .Z(n1301) );
  AND U1319 ( .A(n19), .B(n1306), .Z(n1305) );
  XNOR U1320 ( .A(p_input[139]), .B(n1304), .Z(n1306) );
  XOR U1321 ( .A(n1307), .B(n1308), .Z(n1304) );
  AND U1322 ( .A(n23), .B(n1309), .Z(n1308) );
  XNOR U1323 ( .A(p_input[171]), .B(n1307), .Z(n1309) );
  XOR U1324 ( .A(n1310), .B(n1311), .Z(n1307) );
  AND U1325 ( .A(n27), .B(n1312), .Z(n1311) );
  XNOR U1326 ( .A(p_input[203]), .B(n1310), .Z(n1312) );
  XOR U1327 ( .A(n1313), .B(n1314), .Z(n1310) );
  AND U1328 ( .A(n31), .B(n1315), .Z(n1314) );
  XNOR U1329 ( .A(p_input[235]), .B(n1313), .Z(n1315) );
  XOR U1330 ( .A(n1316), .B(n1317), .Z(n1313) );
  AND U1331 ( .A(n35), .B(n1318), .Z(n1317) );
  XNOR U1332 ( .A(p_input[267]), .B(n1316), .Z(n1318) );
  XOR U1333 ( .A(n1319), .B(n1320), .Z(n1316) );
  AND U1334 ( .A(n39), .B(n1321), .Z(n1320) );
  XNOR U1335 ( .A(p_input[299]), .B(n1319), .Z(n1321) );
  XOR U1336 ( .A(n1322), .B(n1323), .Z(n1319) );
  AND U1337 ( .A(n43), .B(n1324), .Z(n1323) );
  XNOR U1338 ( .A(p_input[331]), .B(n1322), .Z(n1324) );
  XOR U1339 ( .A(n1325), .B(n1326), .Z(n1322) );
  AND U1340 ( .A(n47), .B(n1327), .Z(n1326) );
  XNOR U1341 ( .A(p_input[363]), .B(n1325), .Z(n1327) );
  XOR U1342 ( .A(n1328), .B(n1329), .Z(n1325) );
  AND U1343 ( .A(n51), .B(n1330), .Z(n1329) );
  XNOR U1344 ( .A(p_input[395]), .B(n1328), .Z(n1330) );
  XNOR U1345 ( .A(n1331), .B(n1332), .Z(n1328) );
  AND U1346 ( .A(n55), .B(n1333), .Z(n1332) );
  XOR U1347 ( .A(p_input[427]), .B(n1331), .Z(n1333) );
  XOR U1348 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n1334), .Z(n1331) );
  AND U1349 ( .A(n58), .B(n1335), .Z(n1334) );
  XOR U1350 ( .A(p_input[459]), .B(\knn_comb_/min_val_out[0][11] ), .Z(n1335)
         );
  XNOR U1351 ( .A(n1336), .B(n1337), .Z(o[10]) );
  AND U1352 ( .A(n3), .B(n1338), .Z(n1336) );
  XNOR U1353 ( .A(p_input[10]), .B(n1337), .Z(n1338) );
  XOR U1354 ( .A(n1339), .B(n1340), .Z(n1337) );
  AND U1355 ( .A(n7), .B(n1341), .Z(n1340) );
  XNOR U1356 ( .A(p_input[42]), .B(n1339), .Z(n1341) );
  XOR U1357 ( .A(n1342), .B(n1343), .Z(n1339) );
  AND U1358 ( .A(n11), .B(n1344), .Z(n1343) );
  XNOR U1359 ( .A(p_input[74]), .B(n1342), .Z(n1344) );
  XOR U1360 ( .A(n1345), .B(n1346), .Z(n1342) );
  AND U1361 ( .A(n15), .B(n1347), .Z(n1346) );
  XNOR U1362 ( .A(p_input[106]), .B(n1345), .Z(n1347) );
  XOR U1363 ( .A(n1348), .B(n1349), .Z(n1345) );
  AND U1364 ( .A(n19), .B(n1350), .Z(n1349) );
  XNOR U1365 ( .A(p_input[138]), .B(n1348), .Z(n1350) );
  XOR U1366 ( .A(n1351), .B(n1352), .Z(n1348) );
  AND U1367 ( .A(n23), .B(n1353), .Z(n1352) );
  XNOR U1368 ( .A(p_input[170]), .B(n1351), .Z(n1353) );
  XOR U1369 ( .A(n1354), .B(n1355), .Z(n1351) );
  AND U1370 ( .A(n27), .B(n1356), .Z(n1355) );
  XNOR U1371 ( .A(p_input[202]), .B(n1354), .Z(n1356) );
  XOR U1372 ( .A(n1357), .B(n1358), .Z(n1354) );
  AND U1373 ( .A(n31), .B(n1359), .Z(n1358) );
  XNOR U1374 ( .A(p_input[234]), .B(n1357), .Z(n1359) );
  XOR U1375 ( .A(n1360), .B(n1361), .Z(n1357) );
  AND U1376 ( .A(n35), .B(n1362), .Z(n1361) );
  XNOR U1377 ( .A(p_input[266]), .B(n1360), .Z(n1362) );
  XOR U1378 ( .A(n1363), .B(n1364), .Z(n1360) );
  AND U1379 ( .A(n39), .B(n1365), .Z(n1364) );
  XNOR U1380 ( .A(p_input[298]), .B(n1363), .Z(n1365) );
  XOR U1381 ( .A(n1366), .B(n1367), .Z(n1363) );
  AND U1382 ( .A(n43), .B(n1368), .Z(n1367) );
  XNOR U1383 ( .A(p_input[330]), .B(n1366), .Z(n1368) );
  XOR U1384 ( .A(n1369), .B(n1370), .Z(n1366) );
  AND U1385 ( .A(n47), .B(n1371), .Z(n1370) );
  XNOR U1386 ( .A(p_input[362]), .B(n1369), .Z(n1371) );
  XOR U1387 ( .A(n1372), .B(n1373), .Z(n1369) );
  AND U1388 ( .A(n51), .B(n1374), .Z(n1373) );
  XNOR U1389 ( .A(p_input[394]), .B(n1372), .Z(n1374) );
  XNOR U1390 ( .A(n1375), .B(n1376), .Z(n1372) );
  AND U1391 ( .A(n55), .B(n1377), .Z(n1376) );
  XOR U1392 ( .A(p_input[426]), .B(n1375), .Z(n1377) );
  XOR U1393 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n1378), .Z(n1375) );
  AND U1394 ( .A(n58), .B(n1379), .Z(n1378) );
  XOR U1395 ( .A(p_input[458]), .B(\knn_comb_/min_val_out[0][10] ), .Z(n1379)
         );
  XNOR U1396 ( .A(n1380), .B(n1381), .Z(o[0]) );
  AND U1397 ( .A(n3), .B(n1382), .Z(n1380) );
  XNOR U1398 ( .A(p_input[0]), .B(n1381), .Z(n1382) );
  XOR U1399 ( .A(n1383), .B(n1384), .Z(n1381) );
  AND U1400 ( .A(n7), .B(n1385), .Z(n1384) );
  XNOR U1401 ( .A(p_input[32]), .B(n1383), .Z(n1385) );
  XOR U1402 ( .A(n1386), .B(n1387), .Z(n1383) );
  AND U1403 ( .A(n11), .B(n1388), .Z(n1387) );
  XNOR U1404 ( .A(p_input[64]), .B(n1386), .Z(n1388) );
  XOR U1405 ( .A(n1389), .B(n1390), .Z(n1386) );
  AND U1406 ( .A(n15), .B(n1391), .Z(n1390) );
  XNOR U1407 ( .A(p_input[96]), .B(n1389), .Z(n1391) );
  XOR U1408 ( .A(n1392), .B(n1393), .Z(n1389) );
  AND U1409 ( .A(n19), .B(n1394), .Z(n1393) );
  XNOR U1410 ( .A(p_input[128]), .B(n1392), .Z(n1394) );
  XOR U1411 ( .A(n1395), .B(n1396), .Z(n1392) );
  AND U1412 ( .A(n23), .B(n1397), .Z(n1396) );
  XNOR U1413 ( .A(p_input[160]), .B(n1395), .Z(n1397) );
  XOR U1414 ( .A(n1398), .B(n1399), .Z(n1395) );
  AND U1415 ( .A(n27), .B(n1400), .Z(n1399) );
  XNOR U1416 ( .A(p_input[192]), .B(n1398), .Z(n1400) );
  XOR U1417 ( .A(n1401), .B(n1402), .Z(n1398) );
  AND U1418 ( .A(n31), .B(n1403), .Z(n1402) );
  XNOR U1419 ( .A(p_input[224]), .B(n1401), .Z(n1403) );
  XOR U1420 ( .A(n1404), .B(n1405), .Z(n1401) );
  AND U1421 ( .A(n35), .B(n1406), .Z(n1405) );
  XNOR U1422 ( .A(p_input[256]), .B(n1404), .Z(n1406) );
  XOR U1423 ( .A(n1407), .B(n1408), .Z(n1404) );
  AND U1424 ( .A(n39), .B(n1409), .Z(n1408) );
  XNOR U1425 ( .A(p_input[288]), .B(n1407), .Z(n1409) );
  XOR U1426 ( .A(n1410), .B(n1411), .Z(n1407) );
  AND U1427 ( .A(n43), .B(n1412), .Z(n1411) );
  XNOR U1428 ( .A(p_input[320]), .B(n1410), .Z(n1412) );
  XOR U1429 ( .A(n1413), .B(n1414), .Z(n1410) );
  AND U1430 ( .A(n47), .B(n1415), .Z(n1414) );
  XNOR U1431 ( .A(p_input[352]), .B(n1413), .Z(n1415) );
  XOR U1432 ( .A(n1416), .B(n1417), .Z(n1413) );
  AND U1433 ( .A(n51), .B(n1418), .Z(n1417) );
  XNOR U1434 ( .A(p_input[384]), .B(n1416), .Z(n1418) );
  XNOR U1435 ( .A(n1419), .B(n1420), .Z(n1416) );
  AND U1436 ( .A(n55), .B(n1421), .Z(n1420) );
  XOR U1437 ( .A(p_input[416]), .B(n1419), .Z(n1421) );
  XOR U1438 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n1422), .Z(n1419) );
  AND U1439 ( .A(n58), .B(n1423), .Z(n1422) );
  XOR U1440 ( .A(p_input[448]), .B(\knn_comb_/min_val_out[0][0] ), .Z(n1423)
         );
  XNOR U1441 ( .A(n1424), .B(n1425), .Z(n3) );
  AND U1442 ( .A(n1426), .B(n1427), .Z(n1425) );
  XOR U1443 ( .A(n1428), .B(n1424), .Z(n1427) );
  AND U1444 ( .A(n1429), .B(n1430), .Z(n1428) );
  XOR U1445 ( .A(n1431), .B(n1424), .Z(n1426) );
  XNOR U1446 ( .A(n1432), .B(n1433), .Z(n1431) );
  AND U1447 ( .A(n7), .B(n1434), .Z(n1433) );
  XOR U1448 ( .A(n1435), .B(n1432), .Z(n1434) );
  XOR U1449 ( .A(n1436), .B(n1437), .Z(n1424) );
  AND U1450 ( .A(n1438), .B(n1439), .Z(n1437) );
  XNOR U1451 ( .A(n1436), .B(n1429), .Z(n1439) );
  XNOR U1452 ( .A(n1440), .B(n1441), .Z(n1429) );
  XOR U1453 ( .A(n1442), .B(n1430), .Z(n1441) );
  AND U1454 ( .A(n1443), .B(n1444), .Z(n1430) );
  AND U1455 ( .A(n1445), .B(n1446), .Z(n1442) );
  XOR U1456 ( .A(n1447), .B(n1440), .Z(n1445) );
  XOR U1457 ( .A(n1448), .B(n1436), .Z(n1438) );
  XNOR U1458 ( .A(n1449), .B(n1450), .Z(n1448) );
  AND U1459 ( .A(n7), .B(n1451), .Z(n1450) );
  XOR U1460 ( .A(n1452), .B(n1449), .Z(n1451) );
  XOR U1461 ( .A(n1453), .B(n1454), .Z(n1436) );
  AND U1462 ( .A(n1455), .B(n1456), .Z(n1454) );
  XNOR U1463 ( .A(n1453), .B(n1443), .Z(n1456) );
  XOR U1464 ( .A(n1457), .B(n1446), .Z(n1443) );
  XNOR U1465 ( .A(n1458), .B(n1440), .Z(n1446) );
  XOR U1466 ( .A(n1459), .B(n1460), .Z(n1440) );
  AND U1467 ( .A(n1461), .B(n1462), .Z(n1460) );
  XOR U1468 ( .A(n1463), .B(n1459), .Z(n1461) );
  XNOR U1469 ( .A(n1464), .B(n1465), .Z(n1458) );
  AND U1470 ( .A(n1466), .B(n1467), .Z(n1465) );
  XOR U1471 ( .A(n1464), .B(n1468), .Z(n1466) );
  XNOR U1472 ( .A(n1447), .B(n1444), .Z(n1457) );
  AND U1473 ( .A(n1469), .B(n1470), .Z(n1444) );
  XOR U1474 ( .A(n1471), .B(n1472), .Z(n1447) );
  AND U1475 ( .A(n1473), .B(n1474), .Z(n1472) );
  XOR U1476 ( .A(n1471), .B(n1475), .Z(n1473) );
  XOR U1477 ( .A(n1476), .B(n1453), .Z(n1455) );
  XNOR U1478 ( .A(n1477), .B(n1478), .Z(n1476) );
  AND U1479 ( .A(n7), .B(n1479), .Z(n1478) );
  XNOR U1480 ( .A(n1480), .B(n1477), .Z(n1479) );
  XOR U1481 ( .A(n1481), .B(n1482), .Z(n1453) );
  AND U1482 ( .A(n1483), .B(n1484), .Z(n1482) );
  XNOR U1483 ( .A(n1481), .B(n1469), .Z(n1484) );
  XOR U1484 ( .A(n1485), .B(n1462), .Z(n1469) );
  XNOR U1485 ( .A(n1486), .B(n1468), .Z(n1462) );
  XOR U1486 ( .A(n1487), .B(n1488), .Z(n1468) );
  AND U1487 ( .A(n1489), .B(n1490), .Z(n1488) );
  XOR U1488 ( .A(n1487), .B(n1491), .Z(n1489) );
  XNOR U1489 ( .A(n1467), .B(n1459), .Z(n1486) );
  XOR U1490 ( .A(n1492), .B(n1493), .Z(n1459) );
  AND U1491 ( .A(n1494), .B(n1495), .Z(n1493) );
  XNOR U1492 ( .A(n1496), .B(n1492), .Z(n1494) );
  XNOR U1493 ( .A(n1497), .B(n1464), .Z(n1467) );
  XOR U1494 ( .A(n1498), .B(n1499), .Z(n1464) );
  AND U1495 ( .A(n1500), .B(n1501), .Z(n1499) );
  XOR U1496 ( .A(n1498), .B(n1502), .Z(n1500) );
  XNOR U1497 ( .A(n1503), .B(n1504), .Z(n1497) );
  AND U1498 ( .A(n1505), .B(n1506), .Z(n1504) );
  XNOR U1499 ( .A(n1503), .B(n1507), .Z(n1505) );
  XNOR U1500 ( .A(n1463), .B(n1470), .Z(n1485) );
  AND U1501 ( .A(n1508), .B(n1509), .Z(n1470) );
  XOR U1502 ( .A(n1475), .B(n1474), .Z(n1463) );
  XNOR U1503 ( .A(n1510), .B(n1471), .Z(n1474) );
  XOR U1504 ( .A(n1511), .B(n1512), .Z(n1471) );
  AND U1505 ( .A(n1513), .B(n1514), .Z(n1512) );
  XOR U1506 ( .A(n1511), .B(n1515), .Z(n1513) );
  XNOR U1507 ( .A(n1516), .B(n1517), .Z(n1510) );
  AND U1508 ( .A(n1518), .B(n1519), .Z(n1517) );
  XOR U1509 ( .A(n1516), .B(n1520), .Z(n1518) );
  XOR U1510 ( .A(n1521), .B(n1522), .Z(n1475) );
  AND U1511 ( .A(n1523), .B(n1524), .Z(n1522) );
  XOR U1512 ( .A(n1521), .B(n1525), .Z(n1523) );
  XOR U1513 ( .A(n1526), .B(n1481), .Z(n1483) );
  XNOR U1514 ( .A(n1527), .B(n1528), .Z(n1526) );
  AND U1515 ( .A(n7), .B(n1529), .Z(n1528) );
  XOR U1516 ( .A(n1530), .B(n1527), .Z(n1529) );
  XOR U1517 ( .A(n1531), .B(n1532), .Z(n1481) );
  AND U1518 ( .A(n1533), .B(n1534), .Z(n1532) );
  XNOR U1519 ( .A(n1531), .B(n1508), .Z(n1534) );
  XOR U1520 ( .A(n1535), .B(n1495), .Z(n1508) );
  XNOR U1521 ( .A(n1536), .B(n1502), .Z(n1495) );
  XOR U1522 ( .A(n1491), .B(n1490), .Z(n1502) );
  XNOR U1523 ( .A(n1537), .B(n1487), .Z(n1490) );
  XOR U1524 ( .A(n1538), .B(n1539), .Z(n1487) );
  AND U1525 ( .A(n1540), .B(n1541), .Z(n1539) );
  XNOR U1526 ( .A(n1542), .B(n1543), .Z(n1540) );
  IV U1527 ( .A(n1538), .Z(n1542) );
  XNOR U1528 ( .A(n1544), .B(n1545), .Z(n1537) );
  NOR U1529 ( .A(n1546), .B(n1547), .Z(n1545) );
  XNOR U1530 ( .A(n1544), .B(n1548), .Z(n1546) );
  XOR U1531 ( .A(n1549), .B(n1550), .Z(n1491) );
  NOR U1532 ( .A(n1551), .B(n1552), .Z(n1550) );
  XNOR U1533 ( .A(n1549), .B(n1553), .Z(n1551) );
  XNOR U1534 ( .A(n1501), .B(n1492), .Z(n1536) );
  XOR U1535 ( .A(n1554), .B(n1555), .Z(n1492) );
  AND U1536 ( .A(n1556), .B(n1557), .Z(n1555) );
  XOR U1537 ( .A(n1554), .B(n1558), .Z(n1556) );
  XOR U1538 ( .A(n1559), .B(n1507), .Z(n1501) );
  XOR U1539 ( .A(n1560), .B(n1561), .Z(n1507) );
  NOR U1540 ( .A(n1562), .B(n1563), .Z(n1561) );
  XOR U1541 ( .A(n1560), .B(n1564), .Z(n1562) );
  XNOR U1542 ( .A(n1506), .B(n1498), .Z(n1559) );
  XOR U1543 ( .A(n1565), .B(n1566), .Z(n1498) );
  AND U1544 ( .A(n1567), .B(n1568), .Z(n1566) );
  XOR U1545 ( .A(n1565), .B(n1569), .Z(n1567) );
  XNOR U1546 ( .A(n1570), .B(n1503), .Z(n1506) );
  XOR U1547 ( .A(n1571), .B(n1572), .Z(n1503) );
  AND U1548 ( .A(n1573), .B(n1574), .Z(n1572) );
  XNOR U1549 ( .A(n1575), .B(n1576), .Z(n1573) );
  IV U1550 ( .A(n1571), .Z(n1575) );
  XNOR U1551 ( .A(n1577), .B(n1578), .Z(n1570) );
  NOR U1552 ( .A(n1579), .B(n1580), .Z(n1578) );
  XNOR U1553 ( .A(n1577), .B(n1581), .Z(n1579) );
  XOR U1554 ( .A(n1496), .B(n1509), .Z(n1535) );
  NOR U1555 ( .A(n1582), .B(n1583), .Z(n1509) );
  XNOR U1556 ( .A(n1515), .B(n1514), .Z(n1496) );
  XNOR U1557 ( .A(n1584), .B(n1520), .Z(n1514) );
  XNOR U1558 ( .A(n1585), .B(n1586), .Z(n1520) );
  NOR U1559 ( .A(n1587), .B(n1588), .Z(n1586) );
  XOR U1560 ( .A(n1585), .B(n1589), .Z(n1587) );
  XNOR U1561 ( .A(n1519), .B(n1511), .Z(n1584) );
  XOR U1562 ( .A(n1590), .B(n1591), .Z(n1511) );
  AND U1563 ( .A(n1592), .B(n1593), .Z(n1591) );
  XNOR U1564 ( .A(n1590), .B(n1594), .Z(n1592) );
  XNOR U1565 ( .A(n1595), .B(n1516), .Z(n1519) );
  XOR U1566 ( .A(n1596), .B(n1597), .Z(n1516) );
  AND U1567 ( .A(n1598), .B(n1599), .Z(n1597) );
  XNOR U1568 ( .A(n1600), .B(n1601), .Z(n1598) );
  IV U1569 ( .A(n1596), .Z(n1600) );
  XNOR U1570 ( .A(n1602), .B(n1603), .Z(n1595) );
  NOR U1571 ( .A(n1604), .B(n1605), .Z(n1603) );
  XNOR U1572 ( .A(n1602), .B(n1606), .Z(n1604) );
  XOR U1573 ( .A(n1525), .B(n1524), .Z(n1515) );
  XNOR U1574 ( .A(n1607), .B(n1521), .Z(n1524) );
  XOR U1575 ( .A(n1608), .B(n1609), .Z(n1521) );
  AND U1576 ( .A(n1610), .B(n1611), .Z(n1609) );
  XNOR U1577 ( .A(n1612), .B(n1613), .Z(n1610) );
  IV U1578 ( .A(n1608), .Z(n1612) );
  XNOR U1579 ( .A(n1614), .B(n1615), .Z(n1607) );
  NOR U1580 ( .A(n1616), .B(n1617), .Z(n1615) );
  XNOR U1581 ( .A(n1614), .B(n1618), .Z(n1616) );
  XOR U1582 ( .A(n1619), .B(n1620), .Z(n1525) );
  NOR U1583 ( .A(n1621), .B(n1622), .Z(n1620) );
  XNOR U1584 ( .A(n1619), .B(n1623), .Z(n1621) );
  XNOR U1585 ( .A(n1624), .B(n1625), .Z(n1533) );
  XOR U1586 ( .A(n1531), .B(n1626), .Z(n1625) );
  AND U1587 ( .A(n7), .B(n1627), .Z(n1626) );
  XNOR U1588 ( .A(n1628), .B(n1624), .Z(n1627) );
  AND U1589 ( .A(n1629), .B(n1582), .Z(n1531) );
  XOR U1590 ( .A(n1630), .B(n1583), .Z(n1582) );
  XNOR U1591 ( .A(p_input[0]), .B(p_input[512]), .Z(n1583) );
  XNOR U1592 ( .A(n1558), .B(n1557), .Z(n1630) );
  XNOR U1593 ( .A(n1631), .B(n1569), .Z(n1557) );
  XOR U1594 ( .A(n1543), .B(n1541), .Z(n1569) );
  XNOR U1595 ( .A(n1632), .B(n1548), .Z(n1541) );
  XOR U1596 ( .A(p_input[24]), .B(p_input[536]), .Z(n1548) );
  XOR U1597 ( .A(n1538), .B(n1547), .Z(n1632) );
  XOR U1598 ( .A(n1633), .B(n1544), .Z(n1547) );
  XOR U1599 ( .A(p_input[22]), .B(p_input[534]), .Z(n1544) );
  XOR U1600 ( .A(p_input[23]), .B(n1634), .Z(n1633) );
  XOR U1601 ( .A(p_input[18]), .B(p_input[530]), .Z(n1538) );
  XNOR U1602 ( .A(n1553), .B(n1552), .Z(n1543) );
  XOR U1603 ( .A(n1635), .B(n1549), .Z(n1552) );
  XOR U1604 ( .A(p_input[19]), .B(p_input[531]), .Z(n1549) );
  XOR U1605 ( .A(p_input[20]), .B(n1636), .Z(n1635) );
  XOR U1606 ( .A(p_input[21]), .B(p_input[533]), .Z(n1553) );
  XOR U1607 ( .A(n1568), .B(n1637), .Z(n1631) );
  IV U1608 ( .A(n1554), .Z(n1637) );
  XOR U1609 ( .A(p_input[1]), .B(p_input[513]), .Z(n1554) );
  XNOR U1610 ( .A(n1638), .B(n1576), .Z(n1568) );
  XNOR U1611 ( .A(n1564), .B(n1563), .Z(n1576) );
  XNOR U1612 ( .A(n1639), .B(n1560), .Z(n1563) );
  XNOR U1613 ( .A(p_input[26]), .B(p_input[538]), .Z(n1560) );
  XOR U1614 ( .A(p_input[27]), .B(n1640), .Z(n1639) );
  XOR U1615 ( .A(p_input[28]), .B(p_input[540]), .Z(n1564) );
  XOR U1616 ( .A(n1574), .B(n1641), .Z(n1638) );
  IV U1617 ( .A(n1565), .Z(n1641) );
  XOR U1618 ( .A(p_input[17]), .B(p_input[529]), .Z(n1565) );
  XNOR U1619 ( .A(n1642), .B(n1581), .Z(n1574) );
  XNOR U1620 ( .A(p_input[31]), .B(n1643), .Z(n1581) );
  XOR U1621 ( .A(n1571), .B(n1580), .Z(n1642) );
  XOR U1622 ( .A(n1644), .B(n1577), .Z(n1580) );
  XOR U1623 ( .A(p_input[29]), .B(p_input[541]), .Z(n1577) );
  XOR U1624 ( .A(p_input[30]), .B(n1645), .Z(n1644) );
  XOR U1625 ( .A(p_input[25]), .B(p_input[537]), .Z(n1571) );
  XNOR U1626 ( .A(n1594), .B(n1593), .Z(n1558) );
  XNOR U1627 ( .A(n1646), .B(n1601), .Z(n1593) );
  XNOR U1628 ( .A(n1589), .B(n1588), .Z(n1601) );
  XNOR U1629 ( .A(n1647), .B(n1585), .Z(n1588) );
  XNOR U1630 ( .A(p_input[11]), .B(p_input[523]), .Z(n1585) );
  XOR U1631 ( .A(p_input[12]), .B(n1648), .Z(n1647) );
  XOR U1632 ( .A(p_input[13]), .B(p_input[525]), .Z(n1589) );
  XOR U1633 ( .A(n1599), .B(n1649), .Z(n1646) );
  IV U1634 ( .A(n1590), .Z(n1649) );
  XOR U1635 ( .A(p_input[2]), .B(p_input[514]), .Z(n1590) );
  XNOR U1636 ( .A(n1650), .B(n1606), .Z(n1599) );
  XNOR U1637 ( .A(p_input[16]), .B(n1651), .Z(n1606) );
  XOR U1638 ( .A(n1596), .B(n1605), .Z(n1650) );
  XOR U1639 ( .A(n1652), .B(n1602), .Z(n1605) );
  XOR U1640 ( .A(p_input[14]), .B(p_input[526]), .Z(n1602) );
  XOR U1641 ( .A(p_input[15]), .B(n1653), .Z(n1652) );
  XOR U1642 ( .A(p_input[10]), .B(p_input[522]), .Z(n1596) );
  XNOR U1643 ( .A(n1613), .B(n1611), .Z(n1594) );
  XNOR U1644 ( .A(n1654), .B(n1618), .Z(n1611) );
  XOR U1645 ( .A(p_input[521]), .B(p_input[9]), .Z(n1618) );
  XOR U1646 ( .A(n1608), .B(n1617), .Z(n1654) );
  XOR U1647 ( .A(n1655), .B(n1614), .Z(n1617) );
  XOR U1648 ( .A(p_input[519]), .B(p_input[7]), .Z(n1614) );
  XNOR U1649 ( .A(p_input[520]), .B(p_input[8]), .Z(n1655) );
  XOR U1650 ( .A(p_input[3]), .B(p_input[515]), .Z(n1608) );
  XNOR U1651 ( .A(n1623), .B(n1622), .Z(n1613) );
  XOR U1652 ( .A(n1656), .B(n1619), .Z(n1622) );
  XOR U1653 ( .A(p_input[4]), .B(p_input[516]), .Z(n1619) );
  XNOR U1654 ( .A(p_input[517]), .B(p_input[5]), .Z(n1656) );
  XOR U1655 ( .A(p_input[518]), .B(p_input[6]), .Z(n1623) );
  XNOR U1656 ( .A(n1657), .B(n1658), .Z(n1629) );
  AND U1657 ( .A(n7), .B(n1659), .Z(n1658) );
  XNOR U1658 ( .A(n1660), .B(n1661), .Z(n1659) );
  XNOR U1659 ( .A(n1662), .B(n1663), .Z(n7) );
  AND U1660 ( .A(n1664), .B(n1665), .Z(n1663) );
  XOR U1661 ( .A(n1435), .B(n1662), .Z(n1665) );
  AND U1662 ( .A(n1666), .B(n1667), .Z(n1435) );
  XNOR U1663 ( .A(n1432), .B(n1662), .Z(n1664) );
  XOR U1664 ( .A(n1668), .B(n1669), .Z(n1432) );
  AND U1665 ( .A(n11), .B(n1670), .Z(n1669) );
  XOR U1666 ( .A(n1671), .B(n1668), .Z(n1670) );
  XOR U1667 ( .A(n1672), .B(n1673), .Z(n1662) );
  AND U1668 ( .A(n1674), .B(n1675), .Z(n1673) );
  XNOR U1669 ( .A(n1672), .B(n1666), .Z(n1675) );
  IV U1670 ( .A(n1452), .Z(n1666) );
  XOR U1671 ( .A(n1676), .B(n1677), .Z(n1452) );
  XOR U1672 ( .A(n1678), .B(n1667), .Z(n1677) );
  AND U1673 ( .A(n1480), .B(n1679), .Z(n1667) );
  AND U1674 ( .A(n1680), .B(n1681), .Z(n1678) );
  XOR U1675 ( .A(n1682), .B(n1676), .Z(n1680) );
  XNOR U1676 ( .A(n1449), .B(n1672), .Z(n1674) );
  XOR U1677 ( .A(n1683), .B(n1684), .Z(n1449) );
  AND U1678 ( .A(n11), .B(n1685), .Z(n1684) );
  XOR U1679 ( .A(n1686), .B(n1683), .Z(n1685) );
  XOR U1680 ( .A(n1687), .B(n1688), .Z(n1672) );
  AND U1681 ( .A(n1689), .B(n1690), .Z(n1688) );
  XNOR U1682 ( .A(n1687), .B(n1480), .Z(n1690) );
  XOR U1683 ( .A(n1691), .B(n1681), .Z(n1480) );
  XNOR U1684 ( .A(n1692), .B(n1676), .Z(n1681) );
  XOR U1685 ( .A(n1693), .B(n1694), .Z(n1676) );
  AND U1686 ( .A(n1695), .B(n1696), .Z(n1694) );
  XOR U1687 ( .A(n1697), .B(n1693), .Z(n1695) );
  XNOR U1688 ( .A(n1698), .B(n1699), .Z(n1692) );
  AND U1689 ( .A(n1700), .B(n1701), .Z(n1699) );
  XOR U1690 ( .A(n1698), .B(n1702), .Z(n1700) );
  XNOR U1691 ( .A(n1682), .B(n1679), .Z(n1691) );
  AND U1692 ( .A(n1703), .B(n1704), .Z(n1679) );
  XOR U1693 ( .A(n1705), .B(n1706), .Z(n1682) );
  AND U1694 ( .A(n1707), .B(n1708), .Z(n1706) );
  XOR U1695 ( .A(n1705), .B(n1709), .Z(n1707) );
  XNOR U1696 ( .A(n1477), .B(n1687), .Z(n1689) );
  XOR U1697 ( .A(n1710), .B(n1711), .Z(n1477) );
  AND U1698 ( .A(n11), .B(n1712), .Z(n1711) );
  XNOR U1699 ( .A(n1713), .B(n1710), .Z(n1712) );
  XOR U1700 ( .A(n1714), .B(n1715), .Z(n1687) );
  AND U1701 ( .A(n1716), .B(n1717), .Z(n1715) );
  XNOR U1702 ( .A(n1714), .B(n1703), .Z(n1717) );
  IV U1703 ( .A(n1530), .Z(n1703) );
  XNOR U1704 ( .A(n1718), .B(n1696), .Z(n1530) );
  XNOR U1705 ( .A(n1719), .B(n1702), .Z(n1696) );
  XOR U1706 ( .A(n1720), .B(n1721), .Z(n1702) );
  AND U1707 ( .A(n1722), .B(n1723), .Z(n1721) );
  XOR U1708 ( .A(n1720), .B(n1724), .Z(n1722) );
  XNOR U1709 ( .A(n1701), .B(n1693), .Z(n1719) );
  XOR U1710 ( .A(n1725), .B(n1726), .Z(n1693) );
  AND U1711 ( .A(n1727), .B(n1728), .Z(n1726) );
  XNOR U1712 ( .A(n1729), .B(n1725), .Z(n1727) );
  XNOR U1713 ( .A(n1730), .B(n1698), .Z(n1701) );
  XOR U1714 ( .A(n1731), .B(n1732), .Z(n1698) );
  AND U1715 ( .A(n1733), .B(n1734), .Z(n1732) );
  XOR U1716 ( .A(n1731), .B(n1735), .Z(n1733) );
  XNOR U1717 ( .A(n1736), .B(n1737), .Z(n1730) );
  AND U1718 ( .A(n1738), .B(n1739), .Z(n1737) );
  XNOR U1719 ( .A(n1736), .B(n1740), .Z(n1738) );
  XNOR U1720 ( .A(n1697), .B(n1704), .Z(n1718) );
  AND U1721 ( .A(n1628), .B(n1741), .Z(n1704) );
  XOR U1722 ( .A(n1709), .B(n1708), .Z(n1697) );
  XNOR U1723 ( .A(n1742), .B(n1705), .Z(n1708) );
  XOR U1724 ( .A(n1743), .B(n1744), .Z(n1705) );
  AND U1725 ( .A(n1745), .B(n1746), .Z(n1744) );
  XOR U1726 ( .A(n1743), .B(n1747), .Z(n1745) );
  XNOR U1727 ( .A(n1748), .B(n1749), .Z(n1742) );
  AND U1728 ( .A(n1750), .B(n1751), .Z(n1749) );
  XOR U1729 ( .A(n1748), .B(n1752), .Z(n1750) );
  XOR U1730 ( .A(n1753), .B(n1754), .Z(n1709) );
  AND U1731 ( .A(n1755), .B(n1756), .Z(n1754) );
  XOR U1732 ( .A(n1753), .B(n1757), .Z(n1755) );
  XNOR U1733 ( .A(n1527), .B(n1714), .Z(n1716) );
  XOR U1734 ( .A(n1758), .B(n1759), .Z(n1527) );
  AND U1735 ( .A(n11), .B(n1760), .Z(n1759) );
  XOR U1736 ( .A(n1761), .B(n1758), .Z(n1760) );
  XOR U1737 ( .A(n1762), .B(n1763), .Z(n1714) );
  AND U1738 ( .A(n1764), .B(n1765), .Z(n1763) );
  XNOR U1739 ( .A(n1762), .B(n1628), .Z(n1765) );
  XOR U1740 ( .A(n1766), .B(n1728), .Z(n1628) );
  XNOR U1741 ( .A(n1767), .B(n1735), .Z(n1728) );
  XOR U1742 ( .A(n1724), .B(n1723), .Z(n1735) );
  XNOR U1743 ( .A(n1768), .B(n1720), .Z(n1723) );
  XOR U1744 ( .A(n1769), .B(n1770), .Z(n1720) );
  AND U1745 ( .A(n1771), .B(n1772), .Z(n1770) );
  XNOR U1746 ( .A(n1773), .B(n1774), .Z(n1771) );
  IV U1747 ( .A(n1769), .Z(n1773) );
  XNOR U1748 ( .A(n1775), .B(n1776), .Z(n1768) );
  NOR U1749 ( .A(n1777), .B(n1778), .Z(n1776) );
  XNOR U1750 ( .A(n1775), .B(n1779), .Z(n1777) );
  XOR U1751 ( .A(n1780), .B(n1781), .Z(n1724) );
  NOR U1752 ( .A(n1782), .B(n1783), .Z(n1781) );
  XNOR U1753 ( .A(n1780), .B(n1784), .Z(n1782) );
  XNOR U1754 ( .A(n1734), .B(n1725), .Z(n1767) );
  XOR U1755 ( .A(n1785), .B(n1786), .Z(n1725) );
  NOR U1756 ( .A(n1787), .B(n1788), .Z(n1786) );
  XOR U1757 ( .A(n1789), .B(n1790), .Z(n1787) );
  XOR U1758 ( .A(n1791), .B(n1740), .Z(n1734) );
  XNOR U1759 ( .A(n1792), .B(n1793), .Z(n1740) );
  NOR U1760 ( .A(n1794), .B(n1795), .Z(n1793) );
  XNOR U1761 ( .A(n1792), .B(n1796), .Z(n1794) );
  XNOR U1762 ( .A(n1739), .B(n1731), .Z(n1791) );
  XOR U1763 ( .A(n1797), .B(n1798), .Z(n1731) );
  AND U1764 ( .A(n1799), .B(n1800), .Z(n1798) );
  XOR U1765 ( .A(n1797), .B(n1801), .Z(n1799) );
  XNOR U1766 ( .A(n1802), .B(n1736), .Z(n1739) );
  XOR U1767 ( .A(n1803), .B(n1804), .Z(n1736) );
  AND U1768 ( .A(n1805), .B(n1806), .Z(n1804) );
  XOR U1769 ( .A(n1803), .B(n1807), .Z(n1805) );
  XNOR U1770 ( .A(n1808), .B(n1809), .Z(n1802) );
  NOR U1771 ( .A(n1810), .B(n1811), .Z(n1809) );
  XOR U1772 ( .A(n1808), .B(n1812), .Z(n1810) );
  XOR U1773 ( .A(n1729), .B(n1741), .Z(n1766) );
  NOR U1774 ( .A(n1660), .B(n1813), .Z(n1741) );
  XNOR U1775 ( .A(n1747), .B(n1746), .Z(n1729) );
  XNOR U1776 ( .A(n1814), .B(n1752), .Z(n1746) );
  XNOR U1777 ( .A(n1815), .B(n1816), .Z(n1752) );
  NOR U1778 ( .A(n1817), .B(n1818), .Z(n1816) );
  XOR U1779 ( .A(n1815), .B(n1819), .Z(n1817) );
  XNOR U1780 ( .A(n1751), .B(n1743), .Z(n1814) );
  XOR U1781 ( .A(n1820), .B(n1821), .Z(n1743) );
  AND U1782 ( .A(n1822), .B(n1823), .Z(n1821) );
  XOR U1783 ( .A(n1820), .B(n1824), .Z(n1822) );
  XNOR U1784 ( .A(n1825), .B(n1748), .Z(n1751) );
  XOR U1785 ( .A(n1826), .B(n1827), .Z(n1748) );
  AND U1786 ( .A(n1828), .B(n1829), .Z(n1827) );
  XNOR U1787 ( .A(n1830), .B(n1831), .Z(n1828) );
  IV U1788 ( .A(n1826), .Z(n1830) );
  XNOR U1789 ( .A(n1832), .B(n1833), .Z(n1825) );
  NOR U1790 ( .A(n1834), .B(n1835), .Z(n1833) );
  XNOR U1791 ( .A(n1832), .B(n1836), .Z(n1834) );
  XOR U1792 ( .A(n1757), .B(n1756), .Z(n1747) );
  XNOR U1793 ( .A(n1837), .B(n1753), .Z(n1756) );
  XOR U1794 ( .A(n1838), .B(n1839), .Z(n1753) );
  AND U1795 ( .A(n1840), .B(n1841), .Z(n1839) );
  XNOR U1796 ( .A(n1842), .B(n1843), .Z(n1840) );
  IV U1797 ( .A(n1838), .Z(n1842) );
  XNOR U1798 ( .A(n1844), .B(n1845), .Z(n1837) );
  NOR U1799 ( .A(n1846), .B(n1847), .Z(n1845) );
  XNOR U1800 ( .A(n1844), .B(n1848), .Z(n1846) );
  XOR U1801 ( .A(n1849), .B(n1850), .Z(n1757) );
  NOR U1802 ( .A(n1851), .B(n1852), .Z(n1850) );
  XNOR U1803 ( .A(n1849), .B(n1853), .Z(n1851) );
  XNOR U1804 ( .A(n1624), .B(n1762), .Z(n1764) );
  XOR U1805 ( .A(n1854), .B(n1855), .Z(n1624) );
  AND U1806 ( .A(n11), .B(n1856), .Z(n1855) );
  XNOR U1807 ( .A(n1857), .B(n1854), .Z(n1856) );
  AND U1808 ( .A(n1661), .B(n1660), .Z(n1762) );
  XOR U1809 ( .A(n1858), .B(n1813), .Z(n1660) );
  XNOR U1810 ( .A(p_input[32]), .B(p_input[512]), .Z(n1813) );
  XOR U1811 ( .A(n1790), .B(n1788), .Z(n1858) );
  XOR U1812 ( .A(n1859), .B(n1801), .Z(n1788) );
  XOR U1813 ( .A(n1774), .B(n1772), .Z(n1801) );
  XNOR U1814 ( .A(n1860), .B(n1779), .Z(n1772) );
  XOR U1815 ( .A(p_input[536]), .B(p_input[56]), .Z(n1779) );
  XOR U1816 ( .A(n1769), .B(n1778), .Z(n1860) );
  XOR U1817 ( .A(n1861), .B(n1775), .Z(n1778) );
  XOR U1818 ( .A(p_input[534]), .B(p_input[54]), .Z(n1775) );
  XNOR U1819 ( .A(p_input[535]), .B(p_input[55]), .Z(n1861) );
  XOR U1820 ( .A(p_input[50]), .B(p_input[530]), .Z(n1769) );
  XNOR U1821 ( .A(n1784), .B(n1783), .Z(n1774) );
  XOR U1822 ( .A(n1862), .B(n1780), .Z(n1783) );
  XOR U1823 ( .A(p_input[51]), .B(p_input[531]), .Z(n1780) );
  XOR U1824 ( .A(p_input[52]), .B(n1636), .Z(n1862) );
  XOR U1825 ( .A(p_input[533]), .B(p_input[53]), .Z(n1784) );
  XOR U1826 ( .A(n1800), .B(n1789), .Z(n1859) );
  IV U1827 ( .A(n1785), .Z(n1789) );
  XOR U1828 ( .A(p_input[33]), .B(p_input[513]), .Z(n1785) );
  XNOR U1829 ( .A(n1863), .B(n1807), .Z(n1800) );
  XNOR U1830 ( .A(n1796), .B(n1795), .Z(n1807) );
  XOR U1831 ( .A(n1864), .B(n1792), .Z(n1795) );
  XNOR U1832 ( .A(n1865), .B(p_input[58]), .Z(n1792) );
  XNOR U1833 ( .A(p_input[539]), .B(p_input[59]), .Z(n1864) );
  XOR U1834 ( .A(p_input[540]), .B(p_input[60]), .Z(n1796) );
  XOR U1835 ( .A(n1806), .B(n1866), .Z(n1863) );
  IV U1836 ( .A(n1797), .Z(n1866) );
  XOR U1837 ( .A(p_input[49]), .B(p_input[529]), .Z(n1797) );
  XOR U1838 ( .A(n1867), .B(n1812), .Z(n1806) );
  XNOR U1839 ( .A(p_input[543]), .B(p_input[63]), .Z(n1812) );
  XOR U1840 ( .A(n1803), .B(n1811), .Z(n1867) );
  XOR U1841 ( .A(n1868), .B(n1808), .Z(n1811) );
  XOR U1842 ( .A(p_input[541]), .B(p_input[61]), .Z(n1808) );
  XNOR U1843 ( .A(p_input[542]), .B(p_input[62]), .Z(n1868) );
  XNOR U1844 ( .A(n1869), .B(p_input[57]), .Z(n1803) );
  XOR U1845 ( .A(n1824), .B(n1823), .Z(n1790) );
  XNOR U1846 ( .A(n1870), .B(n1831), .Z(n1823) );
  XNOR U1847 ( .A(n1819), .B(n1818), .Z(n1831) );
  XNOR U1848 ( .A(n1871), .B(n1815), .Z(n1818) );
  XNOR U1849 ( .A(p_input[43]), .B(p_input[523]), .Z(n1815) );
  XOR U1850 ( .A(p_input[44]), .B(n1648), .Z(n1871) );
  XOR U1851 ( .A(p_input[45]), .B(p_input[525]), .Z(n1819) );
  XOR U1852 ( .A(n1829), .B(n1872), .Z(n1870) );
  IV U1853 ( .A(n1820), .Z(n1872) );
  XOR U1854 ( .A(p_input[34]), .B(p_input[514]), .Z(n1820) );
  XNOR U1855 ( .A(n1873), .B(n1836), .Z(n1829) );
  XNOR U1856 ( .A(p_input[48]), .B(n1651), .Z(n1836) );
  XOR U1857 ( .A(n1826), .B(n1835), .Z(n1873) );
  XOR U1858 ( .A(n1874), .B(n1832), .Z(n1835) );
  XOR U1859 ( .A(p_input[46]), .B(p_input[526]), .Z(n1832) );
  XOR U1860 ( .A(p_input[47]), .B(n1653), .Z(n1874) );
  XOR U1861 ( .A(p_input[42]), .B(p_input[522]), .Z(n1826) );
  XOR U1862 ( .A(n1843), .B(n1841), .Z(n1824) );
  XNOR U1863 ( .A(n1875), .B(n1848), .Z(n1841) );
  XOR U1864 ( .A(p_input[41]), .B(p_input[521]), .Z(n1848) );
  XOR U1865 ( .A(n1838), .B(n1847), .Z(n1875) );
  XOR U1866 ( .A(n1876), .B(n1844), .Z(n1847) );
  XOR U1867 ( .A(p_input[39]), .B(p_input[519]), .Z(n1844) );
  XOR U1868 ( .A(p_input[40]), .B(n1877), .Z(n1876) );
  XOR U1869 ( .A(p_input[35]), .B(p_input[515]), .Z(n1838) );
  XNOR U1870 ( .A(n1853), .B(n1852), .Z(n1843) );
  XOR U1871 ( .A(n1878), .B(n1849), .Z(n1852) );
  XOR U1872 ( .A(p_input[36]), .B(p_input[516]), .Z(n1849) );
  XOR U1873 ( .A(p_input[37]), .B(n1879), .Z(n1878) );
  XOR U1874 ( .A(p_input[38]), .B(p_input[518]), .Z(n1853) );
  IV U1875 ( .A(n1657), .Z(n1661) );
  XNOR U1876 ( .A(n1880), .B(n1881), .Z(n1657) );
  AND U1877 ( .A(n11), .B(n1882), .Z(n1881) );
  XNOR U1878 ( .A(n1883), .B(n1880), .Z(n1882) );
  XNOR U1879 ( .A(n1884), .B(n1885), .Z(n11) );
  AND U1880 ( .A(n1886), .B(n1887), .Z(n1885) );
  XOR U1881 ( .A(n1671), .B(n1884), .Z(n1887) );
  AND U1882 ( .A(n1888), .B(n1889), .Z(n1671) );
  XNOR U1883 ( .A(n1668), .B(n1884), .Z(n1886) );
  XOR U1884 ( .A(n1890), .B(n1891), .Z(n1668) );
  AND U1885 ( .A(n15), .B(n1892), .Z(n1891) );
  XOR U1886 ( .A(n1893), .B(n1890), .Z(n1892) );
  XOR U1887 ( .A(n1894), .B(n1895), .Z(n1884) );
  AND U1888 ( .A(n1896), .B(n1897), .Z(n1895) );
  XNOR U1889 ( .A(n1894), .B(n1888), .Z(n1897) );
  IV U1890 ( .A(n1686), .Z(n1888) );
  XOR U1891 ( .A(n1898), .B(n1899), .Z(n1686) );
  XOR U1892 ( .A(n1900), .B(n1889), .Z(n1899) );
  AND U1893 ( .A(n1713), .B(n1901), .Z(n1889) );
  AND U1894 ( .A(n1902), .B(n1903), .Z(n1900) );
  XOR U1895 ( .A(n1904), .B(n1898), .Z(n1902) );
  XNOR U1896 ( .A(n1683), .B(n1894), .Z(n1896) );
  XOR U1897 ( .A(n1905), .B(n1906), .Z(n1683) );
  AND U1898 ( .A(n15), .B(n1907), .Z(n1906) );
  XOR U1899 ( .A(n1908), .B(n1905), .Z(n1907) );
  XOR U1900 ( .A(n1909), .B(n1910), .Z(n1894) );
  AND U1901 ( .A(n1911), .B(n1912), .Z(n1910) );
  XNOR U1902 ( .A(n1909), .B(n1713), .Z(n1912) );
  XOR U1903 ( .A(n1913), .B(n1903), .Z(n1713) );
  XNOR U1904 ( .A(n1914), .B(n1898), .Z(n1903) );
  XOR U1905 ( .A(n1915), .B(n1916), .Z(n1898) );
  AND U1906 ( .A(n1917), .B(n1918), .Z(n1916) );
  XOR U1907 ( .A(n1919), .B(n1915), .Z(n1917) );
  XNOR U1908 ( .A(n1920), .B(n1921), .Z(n1914) );
  AND U1909 ( .A(n1922), .B(n1923), .Z(n1921) );
  XOR U1910 ( .A(n1920), .B(n1924), .Z(n1922) );
  XNOR U1911 ( .A(n1904), .B(n1901), .Z(n1913) );
  AND U1912 ( .A(n1925), .B(n1926), .Z(n1901) );
  XOR U1913 ( .A(n1927), .B(n1928), .Z(n1904) );
  AND U1914 ( .A(n1929), .B(n1930), .Z(n1928) );
  XOR U1915 ( .A(n1927), .B(n1931), .Z(n1929) );
  XNOR U1916 ( .A(n1710), .B(n1909), .Z(n1911) );
  XOR U1917 ( .A(n1932), .B(n1933), .Z(n1710) );
  AND U1918 ( .A(n15), .B(n1934), .Z(n1933) );
  XNOR U1919 ( .A(n1935), .B(n1932), .Z(n1934) );
  XOR U1920 ( .A(n1936), .B(n1937), .Z(n1909) );
  AND U1921 ( .A(n1938), .B(n1939), .Z(n1937) );
  XNOR U1922 ( .A(n1936), .B(n1925), .Z(n1939) );
  IV U1923 ( .A(n1761), .Z(n1925) );
  XNOR U1924 ( .A(n1940), .B(n1918), .Z(n1761) );
  XNOR U1925 ( .A(n1941), .B(n1924), .Z(n1918) );
  XOR U1926 ( .A(n1942), .B(n1943), .Z(n1924) );
  AND U1927 ( .A(n1944), .B(n1945), .Z(n1943) );
  XOR U1928 ( .A(n1942), .B(n1946), .Z(n1944) );
  XNOR U1929 ( .A(n1923), .B(n1915), .Z(n1941) );
  XOR U1930 ( .A(n1947), .B(n1948), .Z(n1915) );
  AND U1931 ( .A(n1949), .B(n1950), .Z(n1948) );
  XNOR U1932 ( .A(n1951), .B(n1947), .Z(n1949) );
  XNOR U1933 ( .A(n1952), .B(n1920), .Z(n1923) );
  XOR U1934 ( .A(n1953), .B(n1954), .Z(n1920) );
  AND U1935 ( .A(n1955), .B(n1956), .Z(n1954) );
  XOR U1936 ( .A(n1953), .B(n1957), .Z(n1955) );
  XNOR U1937 ( .A(n1958), .B(n1959), .Z(n1952) );
  AND U1938 ( .A(n1960), .B(n1961), .Z(n1959) );
  XNOR U1939 ( .A(n1958), .B(n1962), .Z(n1960) );
  XNOR U1940 ( .A(n1919), .B(n1926), .Z(n1940) );
  AND U1941 ( .A(n1857), .B(n1963), .Z(n1926) );
  XOR U1942 ( .A(n1931), .B(n1930), .Z(n1919) );
  XNOR U1943 ( .A(n1964), .B(n1927), .Z(n1930) );
  XOR U1944 ( .A(n1965), .B(n1966), .Z(n1927) );
  AND U1945 ( .A(n1967), .B(n1968), .Z(n1966) );
  XOR U1946 ( .A(n1965), .B(n1969), .Z(n1967) );
  XNOR U1947 ( .A(n1970), .B(n1971), .Z(n1964) );
  AND U1948 ( .A(n1972), .B(n1973), .Z(n1971) );
  XOR U1949 ( .A(n1970), .B(n1974), .Z(n1972) );
  XOR U1950 ( .A(n1975), .B(n1976), .Z(n1931) );
  AND U1951 ( .A(n1977), .B(n1978), .Z(n1976) );
  XOR U1952 ( .A(n1975), .B(n1979), .Z(n1977) );
  XNOR U1953 ( .A(n1758), .B(n1936), .Z(n1938) );
  XOR U1954 ( .A(n1980), .B(n1981), .Z(n1758) );
  AND U1955 ( .A(n15), .B(n1982), .Z(n1981) );
  XOR U1956 ( .A(n1983), .B(n1980), .Z(n1982) );
  XOR U1957 ( .A(n1984), .B(n1985), .Z(n1936) );
  AND U1958 ( .A(n1986), .B(n1987), .Z(n1985) );
  XNOR U1959 ( .A(n1984), .B(n1857), .Z(n1987) );
  XOR U1960 ( .A(n1988), .B(n1950), .Z(n1857) );
  XNOR U1961 ( .A(n1989), .B(n1957), .Z(n1950) );
  XOR U1962 ( .A(n1946), .B(n1945), .Z(n1957) );
  XNOR U1963 ( .A(n1990), .B(n1942), .Z(n1945) );
  XOR U1964 ( .A(n1991), .B(n1992), .Z(n1942) );
  AND U1965 ( .A(n1993), .B(n1994), .Z(n1992) );
  XOR U1966 ( .A(n1991), .B(n1995), .Z(n1993) );
  XNOR U1967 ( .A(n1996), .B(n1997), .Z(n1990) );
  NOR U1968 ( .A(n1998), .B(n1999), .Z(n1997) );
  XNOR U1969 ( .A(n1996), .B(n2000), .Z(n1998) );
  XOR U1970 ( .A(n2001), .B(n2002), .Z(n1946) );
  NOR U1971 ( .A(n2003), .B(n2004), .Z(n2002) );
  XNOR U1972 ( .A(n2001), .B(n2005), .Z(n2003) );
  XNOR U1973 ( .A(n1956), .B(n1947), .Z(n1989) );
  XOR U1974 ( .A(n2006), .B(n2007), .Z(n1947) );
  NOR U1975 ( .A(n2008), .B(n2009), .Z(n2007) );
  XNOR U1976 ( .A(n2006), .B(n2010), .Z(n2008) );
  XOR U1977 ( .A(n2011), .B(n1962), .Z(n1956) );
  XNOR U1978 ( .A(n2012), .B(n2013), .Z(n1962) );
  NOR U1979 ( .A(n2014), .B(n2015), .Z(n2013) );
  XNOR U1980 ( .A(n2012), .B(n2016), .Z(n2014) );
  XNOR U1981 ( .A(n1961), .B(n1953), .Z(n2011) );
  XOR U1982 ( .A(n2017), .B(n2018), .Z(n1953) );
  AND U1983 ( .A(n2019), .B(n2020), .Z(n2018) );
  XOR U1984 ( .A(n2017), .B(n2021), .Z(n2019) );
  XNOR U1985 ( .A(n2022), .B(n1958), .Z(n1961) );
  XOR U1986 ( .A(n2023), .B(n2024), .Z(n1958) );
  AND U1987 ( .A(n2025), .B(n2026), .Z(n2024) );
  XOR U1988 ( .A(n2023), .B(n2027), .Z(n2025) );
  XNOR U1989 ( .A(n2028), .B(n2029), .Z(n2022) );
  NOR U1990 ( .A(n2030), .B(n2031), .Z(n2029) );
  XOR U1991 ( .A(n2028), .B(n2032), .Z(n2030) );
  XOR U1992 ( .A(n1951), .B(n1963), .Z(n1988) );
  NOR U1993 ( .A(n1883), .B(n2033), .Z(n1963) );
  XNOR U1994 ( .A(n1969), .B(n1968), .Z(n1951) );
  XNOR U1995 ( .A(n2034), .B(n1974), .Z(n1968) );
  XOR U1996 ( .A(n2035), .B(n2036), .Z(n1974) );
  NOR U1997 ( .A(n2037), .B(n2038), .Z(n2036) );
  XNOR U1998 ( .A(n2035), .B(n2039), .Z(n2037) );
  XNOR U1999 ( .A(n1973), .B(n1965), .Z(n2034) );
  XOR U2000 ( .A(n2040), .B(n2041), .Z(n1965) );
  AND U2001 ( .A(n2042), .B(n2043), .Z(n2041) );
  XNOR U2002 ( .A(n2040), .B(n2044), .Z(n2042) );
  XNOR U2003 ( .A(n2045), .B(n1970), .Z(n1973) );
  XOR U2004 ( .A(n2046), .B(n2047), .Z(n1970) );
  AND U2005 ( .A(n2048), .B(n2049), .Z(n2047) );
  XOR U2006 ( .A(n2046), .B(n2050), .Z(n2048) );
  XNOR U2007 ( .A(n2051), .B(n2052), .Z(n2045) );
  NOR U2008 ( .A(n2053), .B(n2054), .Z(n2052) );
  XOR U2009 ( .A(n2051), .B(n2055), .Z(n2053) );
  XOR U2010 ( .A(n1979), .B(n1978), .Z(n1969) );
  XNOR U2011 ( .A(n2056), .B(n1975), .Z(n1978) );
  XOR U2012 ( .A(n2057), .B(n2058), .Z(n1975) );
  AND U2013 ( .A(n2059), .B(n2060), .Z(n2058) );
  XOR U2014 ( .A(n2057), .B(n2061), .Z(n2059) );
  XNOR U2015 ( .A(n2062), .B(n2063), .Z(n2056) );
  NOR U2016 ( .A(n2064), .B(n2065), .Z(n2063) );
  XNOR U2017 ( .A(n2062), .B(n2066), .Z(n2064) );
  XOR U2018 ( .A(n2067), .B(n2068), .Z(n1979) );
  NOR U2019 ( .A(n2069), .B(n2070), .Z(n2068) );
  XNOR U2020 ( .A(n2067), .B(n2071), .Z(n2069) );
  XNOR U2021 ( .A(n1854), .B(n1984), .Z(n1986) );
  XOR U2022 ( .A(n2072), .B(n2073), .Z(n1854) );
  AND U2023 ( .A(n15), .B(n2074), .Z(n2073) );
  XNOR U2024 ( .A(n2075), .B(n2072), .Z(n2074) );
  AND U2025 ( .A(n1880), .B(n1883), .Z(n1984) );
  XOR U2026 ( .A(n2076), .B(n2033), .Z(n1883) );
  XNOR U2027 ( .A(p_input[512]), .B(p_input[64]), .Z(n2033) );
  XOR U2028 ( .A(n2010), .B(n2009), .Z(n2076) );
  XOR U2029 ( .A(n2077), .B(n2021), .Z(n2009) );
  XOR U2030 ( .A(n1995), .B(n1994), .Z(n2021) );
  XNOR U2031 ( .A(n2078), .B(n2000), .Z(n1994) );
  XOR U2032 ( .A(p_input[536]), .B(p_input[88]), .Z(n2000) );
  XOR U2033 ( .A(n1991), .B(n1999), .Z(n2078) );
  XOR U2034 ( .A(n2079), .B(n1996), .Z(n1999) );
  XOR U2035 ( .A(p_input[534]), .B(p_input[86]), .Z(n1996) );
  XNOR U2036 ( .A(p_input[535]), .B(p_input[87]), .Z(n2079) );
  XNOR U2037 ( .A(n2080), .B(p_input[82]), .Z(n1991) );
  XNOR U2038 ( .A(n2005), .B(n2004), .Z(n1995) );
  XOR U2039 ( .A(n2081), .B(n2001), .Z(n2004) );
  XOR U2040 ( .A(p_input[531]), .B(p_input[83]), .Z(n2001) );
  XNOR U2041 ( .A(p_input[532]), .B(p_input[84]), .Z(n2081) );
  XOR U2042 ( .A(p_input[533]), .B(p_input[85]), .Z(n2005) );
  XNOR U2043 ( .A(n2020), .B(n2006), .Z(n2077) );
  XNOR U2044 ( .A(n2082), .B(p_input[65]), .Z(n2006) );
  XNOR U2045 ( .A(n2083), .B(n2027), .Z(n2020) );
  XNOR U2046 ( .A(n2016), .B(n2015), .Z(n2027) );
  XOR U2047 ( .A(n2084), .B(n2012), .Z(n2015) );
  XNOR U2048 ( .A(n1865), .B(p_input[90]), .Z(n2012) );
  XNOR U2049 ( .A(p_input[539]), .B(p_input[91]), .Z(n2084) );
  XOR U2050 ( .A(p_input[540]), .B(p_input[92]), .Z(n2016) );
  XNOR U2051 ( .A(n2026), .B(n2017), .Z(n2083) );
  XNOR U2052 ( .A(n2085), .B(p_input[81]), .Z(n2017) );
  XOR U2053 ( .A(n2086), .B(n2032), .Z(n2026) );
  XNOR U2054 ( .A(p_input[543]), .B(p_input[95]), .Z(n2032) );
  XOR U2055 ( .A(n2023), .B(n2031), .Z(n2086) );
  XOR U2056 ( .A(n2087), .B(n2028), .Z(n2031) );
  XOR U2057 ( .A(p_input[541]), .B(p_input[93]), .Z(n2028) );
  XNOR U2058 ( .A(p_input[542]), .B(p_input[94]), .Z(n2087) );
  XNOR U2059 ( .A(n1869), .B(p_input[89]), .Z(n2023) );
  XNOR U2060 ( .A(n2044), .B(n2043), .Z(n2010) );
  XNOR U2061 ( .A(n2088), .B(n2050), .Z(n2043) );
  XNOR U2062 ( .A(n2039), .B(n2038), .Z(n2050) );
  XOR U2063 ( .A(n2089), .B(n2035), .Z(n2038) );
  XNOR U2064 ( .A(n2090), .B(p_input[75]), .Z(n2035) );
  XNOR U2065 ( .A(p_input[524]), .B(p_input[76]), .Z(n2089) );
  XOR U2066 ( .A(p_input[525]), .B(p_input[77]), .Z(n2039) );
  XNOR U2067 ( .A(n2049), .B(n2040), .Z(n2088) );
  XNOR U2068 ( .A(n2091), .B(p_input[66]), .Z(n2040) );
  XOR U2069 ( .A(n2092), .B(n2055), .Z(n2049) );
  XNOR U2070 ( .A(p_input[528]), .B(p_input[80]), .Z(n2055) );
  XOR U2071 ( .A(n2046), .B(n2054), .Z(n2092) );
  XOR U2072 ( .A(n2093), .B(n2051), .Z(n2054) );
  XOR U2073 ( .A(p_input[526]), .B(p_input[78]), .Z(n2051) );
  XNOR U2074 ( .A(p_input[527]), .B(p_input[79]), .Z(n2093) );
  XNOR U2075 ( .A(n2094), .B(p_input[74]), .Z(n2046) );
  XNOR U2076 ( .A(n2061), .B(n2060), .Z(n2044) );
  XNOR U2077 ( .A(n2095), .B(n2066), .Z(n2060) );
  XOR U2078 ( .A(p_input[521]), .B(p_input[73]), .Z(n2066) );
  XOR U2079 ( .A(n2057), .B(n2065), .Z(n2095) );
  XOR U2080 ( .A(n2096), .B(n2062), .Z(n2065) );
  XOR U2081 ( .A(p_input[519]), .B(p_input[71]), .Z(n2062) );
  XNOR U2082 ( .A(p_input[520]), .B(p_input[72]), .Z(n2096) );
  XNOR U2083 ( .A(n2097), .B(p_input[67]), .Z(n2057) );
  XNOR U2084 ( .A(n2071), .B(n2070), .Z(n2061) );
  XOR U2085 ( .A(n2098), .B(n2067), .Z(n2070) );
  XOR U2086 ( .A(p_input[516]), .B(p_input[68]), .Z(n2067) );
  XNOR U2087 ( .A(p_input[517]), .B(p_input[69]), .Z(n2098) );
  XOR U2088 ( .A(p_input[518]), .B(p_input[70]), .Z(n2071) );
  XOR U2089 ( .A(n2099), .B(n2100), .Z(n1880) );
  AND U2090 ( .A(n15), .B(n2101), .Z(n2100) );
  XNOR U2091 ( .A(n2102), .B(n2099), .Z(n2101) );
  XNOR U2092 ( .A(n2103), .B(n2104), .Z(n15) );
  AND U2093 ( .A(n2105), .B(n2106), .Z(n2104) );
  XOR U2094 ( .A(n1893), .B(n2103), .Z(n2106) );
  AND U2095 ( .A(n2107), .B(n2108), .Z(n1893) );
  XNOR U2096 ( .A(n1890), .B(n2103), .Z(n2105) );
  XOR U2097 ( .A(n2109), .B(n2110), .Z(n1890) );
  AND U2098 ( .A(n19), .B(n2111), .Z(n2110) );
  XOR U2099 ( .A(n2112), .B(n2109), .Z(n2111) );
  XOR U2100 ( .A(n2113), .B(n2114), .Z(n2103) );
  AND U2101 ( .A(n2115), .B(n2116), .Z(n2114) );
  XNOR U2102 ( .A(n2113), .B(n2107), .Z(n2116) );
  IV U2103 ( .A(n1908), .Z(n2107) );
  XOR U2104 ( .A(n2117), .B(n2118), .Z(n1908) );
  XOR U2105 ( .A(n2119), .B(n2108), .Z(n2118) );
  AND U2106 ( .A(n1935), .B(n2120), .Z(n2108) );
  AND U2107 ( .A(n2121), .B(n2122), .Z(n2119) );
  XOR U2108 ( .A(n2123), .B(n2117), .Z(n2121) );
  XNOR U2109 ( .A(n1905), .B(n2113), .Z(n2115) );
  XOR U2110 ( .A(n2124), .B(n2125), .Z(n1905) );
  AND U2111 ( .A(n19), .B(n2126), .Z(n2125) );
  XOR U2112 ( .A(n2127), .B(n2124), .Z(n2126) );
  XOR U2113 ( .A(n2128), .B(n2129), .Z(n2113) );
  AND U2114 ( .A(n2130), .B(n2131), .Z(n2129) );
  XNOR U2115 ( .A(n2128), .B(n1935), .Z(n2131) );
  XOR U2116 ( .A(n2132), .B(n2122), .Z(n1935) );
  XNOR U2117 ( .A(n2133), .B(n2117), .Z(n2122) );
  XOR U2118 ( .A(n2134), .B(n2135), .Z(n2117) );
  AND U2119 ( .A(n2136), .B(n2137), .Z(n2135) );
  XOR U2120 ( .A(n2138), .B(n2134), .Z(n2136) );
  XNOR U2121 ( .A(n2139), .B(n2140), .Z(n2133) );
  AND U2122 ( .A(n2141), .B(n2142), .Z(n2140) );
  XOR U2123 ( .A(n2139), .B(n2143), .Z(n2141) );
  XNOR U2124 ( .A(n2123), .B(n2120), .Z(n2132) );
  AND U2125 ( .A(n2144), .B(n2145), .Z(n2120) );
  XOR U2126 ( .A(n2146), .B(n2147), .Z(n2123) );
  AND U2127 ( .A(n2148), .B(n2149), .Z(n2147) );
  XOR U2128 ( .A(n2146), .B(n2150), .Z(n2148) );
  XNOR U2129 ( .A(n1932), .B(n2128), .Z(n2130) );
  XOR U2130 ( .A(n2151), .B(n2152), .Z(n1932) );
  AND U2131 ( .A(n19), .B(n2153), .Z(n2152) );
  XNOR U2132 ( .A(n2154), .B(n2151), .Z(n2153) );
  XOR U2133 ( .A(n2155), .B(n2156), .Z(n2128) );
  AND U2134 ( .A(n2157), .B(n2158), .Z(n2156) );
  XNOR U2135 ( .A(n2155), .B(n2144), .Z(n2158) );
  IV U2136 ( .A(n1983), .Z(n2144) );
  XNOR U2137 ( .A(n2159), .B(n2137), .Z(n1983) );
  XNOR U2138 ( .A(n2160), .B(n2143), .Z(n2137) );
  XOR U2139 ( .A(n2161), .B(n2162), .Z(n2143) );
  AND U2140 ( .A(n2163), .B(n2164), .Z(n2162) );
  XOR U2141 ( .A(n2161), .B(n2165), .Z(n2163) );
  XNOR U2142 ( .A(n2142), .B(n2134), .Z(n2160) );
  XOR U2143 ( .A(n2166), .B(n2167), .Z(n2134) );
  AND U2144 ( .A(n2168), .B(n2169), .Z(n2167) );
  XNOR U2145 ( .A(n2170), .B(n2166), .Z(n2168) );
  XNOR U2146 ( .A(n2171), .B(n2139), .Z(n2142) );
  XOR U2147 ( .A(n2172), .B(n2173), .Z(n2139) );
  AND U2148 ( .A(n2174), .B(n2175), .Z(n2173) );
  XOR U2149 ( .A(n2172), .B(n2176), .Z(n2174) );
  XNOR U2150 ( .A(n2177), .B(n2178), .Z(n2171) );
  AND U2151 ( .A(n2179), .B(n2180), .Z(n2178) );
  XNOR U2152 ( .A(n2177), .B(n2181), .Z(n2179) );
  XNOR U2153 ( .A(n2138), .B(n2145), .Z(n2159) );
  AND U2154 ( .A(n2075), .B(n2182), .Z(n2145) );
  XOR U2155 ( .A(n2150), .B(n2149), .Z(n2138) );
  XNOR U2156 ( .A(n2183), .B(n2146), .Z(n2149) );
  XOR U2157 ( .A(n2184), .B(n2185), .Z(n2146) );
  AND U2158 ( .A(n2186), .B(n2187), .Z(n2185) );
  XOR U2159 ( .A(n2184), .B(n2188), .Z(n2186) );
  XNOR U2160 ( .A(n2189), .B(n2190), .Z(n2183) );
  AND U2161 ( .A(n2191), .B(n2192), .Z(n2190) );
  XOR U2162 ( .A(n2189), .B(n2193), .Z(n2191) );
  XOR U2163 ( .A(n2194), .B(n2195), .Z(n2150) );
  AND U2164 ( .A(n2196), .B(n2197), .Z(n2195) );
  XOR U2165 ( .A(n2194), .B(n2198), .Z(n2196) );
  XNOR U2166 ( .A(n1980), .B(n2155), .Z(n2157) );
  XOR U2167 ( .A(n2199), .B(n2200), .Z(n1980) );
  AND U2168 ( .A(n19), .B(n2201), .Z(n2200) );
  XOR U2169 ( .A(n2202), .B(n2199), .Z(n2201) );
  XOR U2170 ( .A(n2203), .B(n2204), .Z(n2155) );
  AND U2171 ( .A(n2205), .B(n2206), .Z(n2204) );
  XNOR U2172 ( .A(n2203), .B(n2075), .Z(n2206) );
  XOR U2173 ( .A(n2207), .B(n2169), .Z(n2075) );
  XNOR U2174 ( .A(n2208), .B(n2176), .Z(n2169) );
  XOR U2175 ( .A(n2165), .B(n2164), .Z(n2176) );
  XNOR U2176 ( .A(n2209), .B(n2161), .Z(n2164) );
  XOR U2177 ( .A(n2210), .B(n2211), .Z(n2161) );
  AND U2178 ( .A(n2212), .B(n2213), .Z(n2211) );
  XNOR U2179 ( .A(n2214), .B(n2215), .Z(n2212) );
  IV U2180 ( .A(n2210), .Z(n2214) );
  XNOR U2181 ( .A(n2216), .B(n2217), .Z(n2209) );
  NOR U2182 ( .A(n2218), .B(n2219), .Z(n2217) );
  XNOR U2183 ( .A(n2216), .B(n2220), .Z(n2218) );
  XOR U2184 ( .A(n2221), .B(n2222), .Z(n2165) );
  NOR U2185 ( .A(n2223), .B(n2224), .Z(n2222) );
  XNOR U2186 ( .A(n2221), .B(n2225), .Z(n2223) );
  XNOR U2187 ( .A(n2175), .B(n2166), .Z(n2208) );
  XOR U2188 ( .A(n2226), .B(n2227), .Z(n2166) );
  AND U2189 ( .A(n2228), .B(n2229), .Z(n2227) );
  XOR U2190 ( .A(n2226), .B(n2230), .Z(n2228) );
  XOR U2191 ( .A(n2231), .B(n2181), .Z(n2175) );
  XOR U2192 ( .A(n2232), .B(n2233), .Z(n2181) );
  NOR U2193 ( .A(n2234), .B(n2235), .Z(n2233) );
  XOR U2194 ( .A(n2232), .B(n2236), .Z(n2234) );
  XNOR U2195 ( .A(n2180), .B(n2172), .Z(n2231) );
  XOR U2196 ( .A(n2237), .B(n2238), .Z(n2172) );
  AND U2197 ( .A(n2239), .B(n2240), .Z(n2238) );
  XOR U2198 ( .A(n2237), .B(n2241), .Z(n2239) );
  XNOR U2199 ( .A(n2242), .B(n2177), .Z(n2180) );
  XOR U2200 ( .A(n2243), .B(n2244), .Z(n2177) );
  AND U2201 ( .A(n2245), .B(n2246), .Z(n2244) );
  XNOR U2202 ( .A(n2247), .B(n2248), .Z(n2245) );
  IV U2203 ( .A(n2243), .Z(n2247) );
  XNOR U2204 ( .A(n2249), .B(n2250), .Z(n2242) );
  NOR U2205 ( .A(n2251), .B(n2252), .Z(n2250) );
  XNOR U2206 ( .A(n2249), .B(n2253), .Z(n2251) );
  XOR U2207 ( .A(n2170), .B(n2182), .Z(n2207) );
  NOR U2208 ( .A(n2102), .B(n2254), .Z(n2182) );
  XNOR U2209 ( .A(n2188), .B(n2187), .Z(n2170) );
  XNOR U2210 ( .A(n2255), .B(n2193), .Z(n2187) );
  XNOR U2211 ( .A(n2256), .B(n2257), .Z(n2193) );
  NOR U2212 ( .A(n2258), .B(n2259), .Z(n2257) );
  XOR U2213 ( .A(n2256), .B(n2260), .Z(n2258) );
  XNOR U2214 ( .A(n2192), .B(n2184), .Z(n2255) );
  XOR U2215 ( .A(n2261), .B(n2262), .Z(n2184) );
  AND U2216 ( .A(n2263), .B(n2264), .Z(n2262) );
  XOR U2217 ( .A(n2261), .B(n2265), .Z(n2263) );
  XNOR U2218 ( .A(n2266), .B(n2189), .Z(n2192) );
  XOR U2219 ( .A(n2267), .B(n2268), .Z(n2189) );
  AND U2220 ( .A(n2269), .B(n2270), .Z(n2268) );
  XNOR U2221 ( .A(n2271), .B(n2272), .Z(n2269) );
  IV U2222 ( .A(n2267), .Z(n2271) );
  XNOR U2223 ( .A(n2273), .B(n2274), .Z(n2266) );
  NOR U2224 ( .A(n2275), .B(n2276), .Z(n2274) );
  XNOR U2225 ( .A(n2273), .B(n2277), .Z(n2275) );
  XOR U2226 ( .A(n2198), .B(n2197), .Z(n2188) );
  XNOR U2227 ( .A(n2278), .B(n2194), .Z(n2197) );
  XOR U2228 ( .A(n2279), .B(n2280), .Z(n2194) );
  AND U2229 ( .A(n2281), .B(n2282), .Z(n2280) );
  XOR U2230 ( .A(n2279), .B(n2283), .Z(n2281) );
  XNOR U2231 ( .A(n2284), .B(n2285), .Z(n2278) );
  NOR U2232 ( .A(n2286), .B(n2287), .Z(n2285) );
  XNOR U2233 ( .A(n2284), .B(n2288), .Z(n2286) );
  XOR U2234 ( .A(n2289), .B(n2290), .Z(n2198) );
  NOR U2235 ( .A(n2291), .B(n2292), .Z(n2290) );
  XNOR U2236 ( .A(n2289), .B(n2293), .Z(n2291) );
  XNOR U2237 ( .A(n2072), .B(n2203), .Z(n2205) );
  XOR U2238 ( .A(n2294), .B(n2295), .Z(n2072) );
  AND U2239 ( .A(n19), .B(n2296), .Z(n2295) );
  XNOR U2240 ( .A(n2297), .B(n2294), .Z(n2296) );
  AND U2241 ( .A(n2099), .B(n2102), .Z(n2203) );
  XOR U2242 ( .A(n2298), .B(n2254), .Z(n2102) );
  XNOR U2243 ( .A(p_input[512]), .B(p_input[96]), .Z(n2254) );
  XNOR U2244 ( .A(n2230), .B(n2229), .Z(n2298) );
  XNOR U2245 ( .A(n2299), .B(n2241), .Z(n2229) );
  XOR U2246 ( .A(n2215), .B(n2213), .Z(n2241) );
  XNOR U2247 ( .A(n2300), .B(n2220), .Z(n2213) );
  XOR U2248 ( .A(p_input[120]), .B(p_input[536]), .Z(n2220) );
  XOR U2249 ( .A(n2210), .B(n2219), .Z(n2300) );
  XOR U2250 ( .A(n2301), .B(n2216), .Z(n2219) );
  XOR U2251 ( .A(p_input[118]), .B(p_input[534]), .Z(n2216) );
  XOR U2252 ( .A(p_input[119]), .B(n1634), .Z(n2301) );
  XOR U2253 ( .A(p_input[114]), .B(p_input[530]), .Z(n2210) );
  XNOR U2254 ( .A(n2225), .B(n2224), .Z(n2215) );
  XOR U2255 ( .A(n2302), .B(n2221), .Z(n2224) );
  XOR U2256 ( .A(p_input[115]), .B(p_input[531]), .Z(n2221) );
  XOR U2257 ( .A(p_input[116]), .B(n1636), .Z(n2302) );
  XOR U2258 ( .A(p_input[117]), .B(p_input[533]), .Z(n2225) );
  XNOR U2259 ( .A(n2240), .B(n2226), .Z(n2299) );
  XNOR U2260 ( .A(n2082), .B(p_input[97]), .Z(n2226) );
  XNOR U2261 ( .A(n2303), .B(n2248), .Z(n2240) );
  XNOR U2262 ( .A(n2236), .B(n2235), .Z(n2248) );
  XNOR U2263 ( .A(n2304), .B(n2232), .Z(n2235) );
  XNOR U2264 ( .A(p_input[122]), .B(p_input[538]), .Z(n2232) );
  XOR U2265 ( .A(p_input[123]), .B(n1640), .Z(n2304) );
  XOR U2266 ( .A(p_input[124]), .B(p_input[540]), .Z(n2236) );
  XOR U2267 ( .A(n2246), .B(n2305), .Z(n2303) );
  IV U2268 ( .A(n2237), .Z(n2305) );
  XOR U2269 ( .A(p_input[113]), .B(p_input[529]), .Z(n2237) );
  XNOR U2270 ( .A(n2306), .B(n2253), .Z(n2246) );
  XNOR U2271 ( .A(p_input[127]), .B(n1643), .Z(n2253) );
  XOR U2272 ( .A(n2243), .B(n2252), .Z(n2306) );
  XOR U2273 ( .A(n2307), .B(n2249), .Z(n2252) );
  XOR U2274 ( .A(p_input[125]), .B(p_input[541]), .Z(n2249) );
  XOR U2275 ( .A(p_input[126]), .B(n1645), .Z(n2307) );
  XOR U2276 ( .A(p_input[121]), .B(p_input[537]), .Z(n2243) );
  XOR U2277 ( .A(n2265), .B(n2264), .Z(n2230) );
  XNOR U2278 ( .A(n2308), .B(n2272), .Z(n2264) );
  XNOR U2279 ( .A(n2260), .B(n2259), .Z(n2272) );
  XNOR U2280 ( .A(n2309), .B(n2256), .Z(n2259) );
  XNOR U2281 ( .A(p_input[107]), .B(p_input[523]), .Z(n2256) );
  XOR U2282 ( .A(p_input[108]), .B(n1648), .Z(n2309) );
  XOR U2283 ( .A(p_input[109]), .B(p_input[525]), .Z(n2260) );
  XNOR U2284 ( .A(n2270), .B(n2261), .Z(n2308) );
  XNOR U2285 ( .A(n2091), .B(p_input[98]), .Z(n2261) );
  XNOR U2286 ( .A(n2310), .B(n2277), .Z(n2270) );
  XNOR U2287 ( .A(p_input[112]), .B(n1651), .Z(n2277) );
  XOR U2288 ( .A(n2267), .B(n2276), .Z(n2310) );
  XOR U2289 ( .A(n2311), .B(n2273), .Z(n2276) );
  XOR U2290 ( .A(p_input[110]), .B(p_input[526]), .Z(n2273) );
  XOR U2291 ( .A(p_input[111]), .B(n1653), .Z(n2311) );
  XOR U2292 ( .A(p_input[106]), .B(p_input[522]), .Z(n2267) );
  XOR U2293 ( .A(n2283), .B(n2282), .Z(n2265) );
  XNOR U2294 ( .A(n2312), .B(n2288), .Z(n2282) );
  XOR U2295 ( .A(p_input[105]), .B(p_input[521]), .Z(n2288) );
  XOR U2296 ( .A(n2279), .B(n2287), .Z(n2312) );
  XOR U2297 ( .A(n2313), .B(n2284), .Z(n2287) );
  XOR U2298 ( .A(p_input[103]), .B(p_input[519]), .Z(n2284) );
  XOR U2299 ( .A(p_input[104]), .B(n1877), .Z(n2313) );
  XNOR U2300 ( .A(n2097), .B(p_input[99]), .Z(n2279) );
  XNOR U2301 ( .A(n2293), .B(n2292), .Z(n2283) );
  XOR U2302 ( .A(n2314), .B(n2289), .Z(n2292) );
  XOR U2303 ( .A(p_input[100]), .B(p_input[516]), .Z(n2289) );
  XOR U2304 ( .A(p_input[101]), .B(n1879), .Z(n2314) );
  XOR U2305 ( .A(p_input[102]), .B(p_input[518]), .Z(n2293) );
  XOR U2306 ( .A(n2315), .B(n2316), .Z(n2099) );
  AND U2307 ( .A(n19), .B(n2317), .Z(n2316) );
  XNOR U2308 ( .A(n2318), .B(n2315), .Z(n2317) );
  XNOR U2309 ( .A(n2319), .B(n2320), .Z(n19) );
  AND U2310 ( .A(n2321), .B(n2322), .Z(n2320) );
  XOR U2311 ( .A(n2112), .B(n2319), .Z(n2322) );
  AND U2312 ( .A(n2323), .B(n2324), .Z(n2112) );
  XNOR U2313 ( .A(n2109), .B(n2319), .Z(n2321) );
  XOR U2314 ( .A(n2325), .B(n2326), .Z(n2109) );
  AND U2315 ( .A(n23), .B(n2327), .Z(n2326) );
  XOR U2316 ( .A(n2328), .B(n2325), .Z(n2327) );
  XOR U2317 ( .A(n2329), .B(n2330), .Z(n2319) );
  AND U2318 ( .A(n2331), .B(n2332), .Z(n2330) );
  XNOR U2319 ( .A(n2329), .B(n2323), .Z(n2332) );
  IV U2320 ( .A(n2127), .Z(n2323) );
  XOR U2321 ( .A(n2333), .B(n2334), .Z(n2127) );
  XOR U2322 ( .A(n2335), .B(n2324), .Z(n2334) );
  AND U2323 ( .A(n2154), .B(n2336), .Z(n2324) );
  AND U2324 ( .A(n2337), .B(n2338), .Z(n2335) );
  XOR U2325 ( .A(n2339), .B(n2333), .Z(n2337) );
  XNOR U2326 ( .A(n2124), .B(n2329), .Z(n2331) );
  XOR U2327 ( .A(n2340), .B(n2341), .Z(n2124) );
  AND U2328 ( .A(n23), .B(n2342), .Z(n2341) );
  XOR U2329 ( .A(n2343), .B(n2340), .Z(n2342) );
  XOR U2330 ( .A(n2344), .B(n2345), .Z(n2329) );
  AND U2331 ( .A(n2346), .B(n2347), .Z(n2345) );
  XNOR U2332 ( .A(n2344), .B(n2154), .Z(n2347) );
  XOR U2333 ( .A(n2348), .B(n2338), .Z(n2154) );
  XNOR U2334 ( .A(n2349), .B(n2333), .Z(n2338) );
  XOR U2335 ( .A(n2350), .B(n2351), .Z(n2333) );
  AND U2336 ( .A(n2352), .B(n2353), .Z(n2351) );
  XOR U2337 ( .A(n2354), .B(n2350), .Z(n2352) );
  XNOR U2338 ( .A(n2355), .B(n2356), .Z(n2349) );
  AND U2339 ( .A(n2357), .B(n2358), .Z(n2356) );
  XOR U2340 ( .A(n2355), .B(n2359), .Z(n2357) );
  XNOR U2341 ( .A(n2339), .B(n2336), .Z(n2348) );
  AND U2342 ( .A(n2360), .B(n2361), .Z(n2336) );
  XOR U2343 ( .A(n2362), .B(n2363), .Z(n2339) );
  AND U2344 ( .A(n2364), .B(n2365), .Z(n2363) );
  XOR U2345 ( .A(n2362), .B(n2366), .Z(n2364) );
  XNOR U2346 ( .A(n2151), .B(n2344), .Z(n2346) );
  XOR U2347 ( .A(n2367), .B(n2368), .Z(n2151) );
  AND U2348 ( .A(n23), .B(n2369), .Z(n2368) );
  XNOR U2349 ( .A(n2370), .B(n2367), .Z(n2369) );
  XOR U2350 ( .A(n2371), .B(n2372), .Z(n2344) );
  AND U2351 ( .A(n2373), .B(n2374), .Z(n2372) );
  XNOR U2352 ( .A(n2371), .B(n2360), .Z(n2374) );
  IV U2353 ( .A(n2202), .Z(n2360) );
  XNOR U2354 ( .A(n2375), .B(n2353), .Z(n2202) );
  XNOR U2355 ( .A(n2376), .B(n2359), .Z(n2353) );
  XOR U2356 ( .A(n2377), .B(n2378), .Z(n2359) );
  AND U2357 ( .A(n2379), .B(n2380), .Z(n2378) );
  XOR U2358 ( .A(n2377), .B(n2381), .Z(n2379) );
  XNOR U2359 ( .A(n2358), .B(n2350), .Z(n2376) );
  XOR U2360 ( .A(n2382), .B(n2383), .Z(n2350) );
  AND U2361 ( .A(n2384), .B(n2385), .Z(n2383) );
  XNOR U2362 ( .A(n2386), .B(n2382), .Z(n2384) );
  XNOR U2363 ( .A(n2387), .B(n2355), .Z(n2358) );
  XOR U2364 ( .A(n2388), .B(n2389), .Z(n2355) );
  AND U2365 ( .A(n2390), .B(n2391), .Z(n2389) );
  XOR U2366 ( .A(n2388), .B(n2392), .Z(n2390) );
  XNOR U2367 ( .A(n2393), .B(n2394), .Z(n2387) );
  AND U2368 ( .A(n2395), .B(n2396), .Z(n2394) );
  XNOR U2369 ( .A(n2393), .B(n2397), .Z(n2395) );
  XNOR U2370 ( .A(n2354), .B(n2361), .Z(n2375) );
  AND U2371 ( .A(n2297), .B(n2398), .Z(n2361) );
  XOR U2372 ( .A(n2366), .B(n2365), .Z(n2354) );
  XNOR U2373 ( .A(n2399), .B(n2362), .Z(n2365) );
  XOR U2374 ( .A(n2400), .B(n2401), .Z(n2362) );
  AND U2375 ( .A(n2402), .B(n2403), .Z(n2401) );
  XOR U2376 ( .A(n2400), .B(n2404), .Z(n2402) );
  XNOR U2377 ( .A(n2405), .B(n2406), .Z(n2399) );
  AND U2378 ( .A(n2407), .B(n2408), .Z(n2406) );
  XOR U2379 ( .A(n2405), .B(n2409), .Z(n2407) );
  XOR U2380 ( .A(n2410), .B(n2411), .Z(n2366) );
  AND U2381 ( .A(n2412), .B(n2413), .Z(n2411) );
  XOR U2382 ( .A(n2410), .B(n2414), .Z(n2412) );
  XNOR U2383 ( .A(n2199), .B(n2371), .Z(n2373) );
  XOR U2384 ( .A(n2415), .B(n2416), .Z(n2199) );
  AND U2385 ( .A(n23), .B(n2417), .Z(n2416) );
  XOR U2386 ( .A(n2418), .B(n2415), .Z(n2417) );
  XOR U2387 ( .A(n2419), .B(n2420), .Z(n2371) );
  AND U2388 ( .A(n2421), .B(n2422), .Z(n2420) );
  XNOR U2389 ( .A(n2419), .B(n2297), .Z(n2422) );
  XOR U2390 ( .A(n2423), .B(n2385), .Z(n2297) );
  XNOR U2391 ( .A(n2424), .B(n2392), .Z(n2385) );
  XOR U2392 ( .A(n2381), .B(n2380), .Z(n2392) );
  XNOR U2393 ( .A(n2425), .B(n2377), .Z(n2380) );
  XOR U2394 ( .A(n2426), .B(n2427), .Z(n2377) );
  AND U2395 ( .A(n2428), .B(n2429), .Z(n2427) );
  XNOR U2396 ( .A(n2430), .B(n2431), .Z(n2428) );
  IV U2397 ( .A(n2426), .Z(n2430) );
  XNOR U2398 ( .A(n2432), .B(n2433), .Z(n2425) );
  NOR U2399 ( .A(n2434), .B(n2435), .Z(n2433) );
  XNOR U2400 ( .A(n2432), .B(n2436), .Z(n2434) );
  XOR U2401 ( .A(n2437), .B(n2438), .Z(n2381) );
  NOR U2402 ( .A(n2439), .B(n2440), .Z(n2438) );
  XNOR U2403 ( .A(n2437), .B(n2441), .Z(n2439) );
  XNOR U2404 ( .A(n2391), .B(n2382), .Z(n2424) );
  XOR U2405 ( .A(n2442), .B(n2443), .Z(n2382) );
  AND U2406 ( .A(n2444), .B(n2445), .Z(n2443) );
  XOR U2407 ( .A(n2442), .B(n2446), .Z(n2444) );
  XOR U2408 ( .A(n2447), .B(n2397), .Z(n2391) );
  XOR U2409 ( .A(n2448), .B(n2449), .Z(n2397) );
  NOR U2410 ( .A(n2450), .B(n2451), .Z(n2449) );
  XOR U2411 ( .A(n2448), .B(n2452), .Z(n2450) );
  XNOR U2412 ( .A(n2396), .B(n2388), .Z(n2447) );
  XOR U2413 ( .A(n2453), .B(n2454), .Z(n2388) );
  AND U2414 ( .A(n2455), .B(n2456), .Z(n2454) );
  XOR U2415 ( .A(n2453), .B(n2457), .Z(n2455) );
  XNOR U2416 ( .A(n2458), .B(n2393), .Z(n2396) );
  XOR U2417 ( .A(n2459), .B(n2460), .Z(n2393) );
  AND U2418 ( .A(n2461), .B(n2462), .Z(n2460) );
  XNOR U2419 ( .A(n2463), .B(n2464), .Z(n2461) );
  IV U2420 ( .A(n2459), .Z(n2463) );
  XNOR U2421 ( .A(n2465), .B(n2466), .Z(n2458) );
  NOR U2422 ( .A(n2467), .B(n2468), .Z(n2466) );
  XNOR U2423 ( .A(n2465), .B(n2469), .Z(n2467) );
  XOR U2424 ( .A(n2386), .B(n2398), .Z(n2423) );
  NOR U2425 ( .A(n2318), .B(n2470), .Z(n2398) );
  XNOR U2426 ( .A(n2404), .B(n2403), .Z(n2386) );
  XNOR U2427 ( .A(n2471), .B(n2409), .Z(n2403) );
  XNOR U2428 ( .A(n2472), .B(n2473), .Z(n2409) );
  NOR U2429 ( .A(n2474), .B(n2475), .Z(n2473) );
  XOR U2430 ( .A(n2472), .B(n2476), .Z(n2474) );
  XNOR U2431 ( .A(n2408), .B(n2400), .Z(n2471) );
  XOR U2432 ( .A(n2477), .B(n2478), .Z(n2400) );
  AND U2433 ( .A(n2479), .B(n2480), .Z(n2478) );
  XOR U2434 ( .A(n2477), .B(n2481), .Z(n2479) );
  XNOR U2435 ( .A(n2482), .B(n2405), .Z(n2408) );
  XOR U2436 ( .A(n2483), .B(n2484), .Z(n2405) );
  AND U2437 ( .A(n2485), .B(n2486), .Z(n2484) );
  XNOR U2438 ( .A(n2487), .B(n2488), .Z(n2485) );
  IV U2439 ( .A(n2483), .Z(n2487) );
  XNOR U2440 ( .A(n2489), .B(n2490), .Z(n2482) );
  NOR U2441 ( .A(n2491), .B(n2492), .Z(n2490) );
  XNOR U2442 ( .A(n2489), .B(n2493), .Z(n2491) );
  XOR U2443 ( .A(n2414), .B(n2413), .Z(n2404) );
  XNOR U2444 ( .A(n2494), .B(n2410), .Z(n2413) );
  XOR U2445 ( .A(n2495), .B(n2496), .Z(n2410) );
  AND U2446 ( .A(n2497), .B(n2498), .Z(n2496) );
  XNOR U2447 ( .A(n2499), .B(n2500), .Z(n2497) );
  IV U2448 ( .A(n2495), .Z(n2499) );
  XNOR U2449 ( .A(n2501), .B(n2502), .Z(n2494) );
  NOR U2450 ( .A(n2503), .B(n2504), .Z(n2502) );
  XNOR U2451 ( .A(n2501), .B(n2505), .Z(n2503) );
  XOR U2452 ( .A(n2506), .B(n2507), .Z(n2414) );
  NOR U2453 ( .A(n2508), .B(n2509), .Z(n2507) );
  XNOR U2454 ( .A(n2506), .B(n2510), .Z(n2508) );
  XNOR U2455 ( .A(n2294), .B(n2419), .Z(n2421) );
  XOR U2456 ( .A(n2511), .B(n2512), .Z(n2294) );
  AND U2457 ( .A(n23), .B(n2513), .Z(n2512) );
  XNOR U2458 ( .A(n2514), .B(n2511), .Z(n2513) );
  AND U2459 ( .A(n2315), .B(n2318), .Z(n2419) );
  XOR U2460 ( .A(n2515), .B(n2470), .Z(n2318) );
  XNOR U2461 ( .A(p_input[128]), .B(p_input[512]), .Z(n2470) );
  XNOR U2462 ( .A(n2446), .B(n2445), .Z(n2515) );
  XNOR U2463 ( .A(n2516), .B(n2457), .Z(n2445) );
  XOR U2464 ( .A(n2431), .B(n2429), .Z(n2457) );
  XNOR U2465 ( .A(n2517), .B(n2436), .Z(n2429) );
  XOR U2466 ( .A(p_input[152]), .B(p_input[536]), .Z(n2436) );
  XOR U2467 ( .A(n2426), .B(n2435), .Z(n2517) );
  XOR U2468 ( .A(n2518), .B(n2432), .Z(n2435) );
  XOR U2469 ( .A(p_input[150]), .B(p_input[534]), .Z(n2432) );
  XOR U2470 ( .A(p_input[151]), .B(n1634), .Z(n2518) );
  XOR U2471 ( .A(p_input[146]), .B(p_input[530]), .Z(n2426) );
  XNOR U2472 ( .A(n2441), .B(n2440), .Z(n2431) );
  XOR U2473 ( .A(n2519), .B(n2437), .Z(n2440) );
  XOR U2474 ( .A(p_input[147]), .B(p_input[531]), .Z(n2437) );
  XOR U2475 ( .A(p_input[148]), .B(n1636), .Z(n2519) );
  XOR U2476 ( .A(p_input[149]), .B(p_input[533]), .Z(n2441) );
  XOR U2477 ( .A(n2456), .B(n2520), .Z(n2516) );
  IV U2478 ( .A(n2442), .Z(n2520) );
  XOR U2479 ( .A(p_input[129]), .B(p_input[513]), .Z(n2442) );
  XNOR U2480 ( .A(n2521), .B(n2464), .Z(n2456) );
  XNOR U2481 ( .A(n2452), .B(n2451), .Z(n2464) );
  XNOR U2482 ( .A(n2522), .B(n2448), .Z(n2451) );
  XNOR U2483 ( .A(p_input[154]), .B(p_input[538]), .Z(n2448) );
  XOR U2484 ( .A(p_input[155]), .B(n1640), .Z(n2522) );
  XOR U2485 ( .A(p_input[156]), .B(p_input[540]), .Z(n2452) );
  XOR U2486 ( .A(n2462), .B(n2523), .Z(n2521) );
  IV U2487 ( .A(n2453), .Z(n2523) );
  XOR U2488 ( .A(p_input[145]), .B(p_input[529]), .Z(n2453) );
  XNOR U2489 ( .A(n2524), .B(n2469), .Z(n2462) );
  XNOR U2490 ( .A(p_input[159]), .B(n1643), .Z(n2469) );
  XOR U2491 ( .A(n2459), .B(n2468), .Z(n2524) );
  XOR U2492 ( .A(n2525), .B(n2465), .Z(n2468) );
  XOR U2493 ( .A(p_input[157]), .B(p_input[541]), .Z(n2465) );
  XOR U2494 ( .A(p_input[158]), .B(n1645), .Z(n2525) );
  XOR U2495 ( .A(p_input[153]), .B(p_input[537]), .Z(n2459) );
  XOR U2496 ( .A(n2481), .B(n2480), .Z(n2446) );
  XNOR U2497 ( .A(n2526), .B(n2488), .Z(n2480) );
  XNOR U2498 ( .A(n2476), .B(n2475), .Z(n2488) );
  XNOR U2499 ( .A(n2527), .B(n2472), .Z(n2475) );
  XNOR U2500 ( .A(p_input[139]), .B(p_input[523]), .Z(n2472) );
  XOR U2501 ( .A(p_input[140]), .B(n1648), .Z(n2527) );
  XOR U2502 ( .A(p_input[141]), .B(p_input[525]), .Z(n2476) );
  XOR U2503 ( .A(n2486), .B(n2528), .Z(n2526) );
  IV U2504 ( .A(n2477), .Z(n2528) );
  XOR U2505 ( .A(p_input[130]), .B(p_input[514]), .Z(n2477) );
  XNOR U2506 ( .A(n2529), .B(n2493), .Z(n2486) );
  XNOR U2507 ( .A(p_input[144]), .B(n1651), .Z(n2493) );
  XOR U2508 ( .A(n2483), .B(n2492), .Z(n2529) );
  XOR U2509 ( .A(n2530), .B(n2489), .Z(n2492) );
  XOR U2510 ( .A(p_input[142]), .B(p_input[526]), .Z(n2489) );
  XOR U2511 ( .A(p_input[143]), .B(n1653), .Z(n2530) );
  XOR U2512 ( .A(p_input[138]), .B(p_input[522]), .Z(n2483) );
  XOR U2513 ( .A(n2500), .B(n2498), .Z(n2481) );
  XNOR U2514 ( .A(n2531), .B(n2505), .Z(n2498) );
  XOR U2515 ( .A(p_input[137]), .B(p_input[521]), .Z(n2505) );
  XOR U2516 ( .A(n2495), .B(n2504), .Z(n2531) );
  XOR U2517 ( .A(n2532), .B(n2501), .Z(n2504) );
  XOR U2518 ( .A(p_input[135]), .B(p_input[519]), .Z(n2501) );
  XOR U2519 ( .A(p_input[136]), .B(n1877), .Z(n2532) );
  XOR U2520 ( .A(p_input[131]), .B(p_input[515]), .Z(n2495) );
  XNOR U2521 ( .A(n2510), .B(n2509), .Z(n2500) );
  XOR U2522 ( .A(n2533), .B(n2506), .Z(n2509) );
  XOR U2523 ( .A(p_input[132]), .B(p_input[516]), .Z(n2506) );
  XOR U2524 ( .A(p_input[133]), .B(n1879), .Z(n2533) );
  XOR U2525 ( .A(p_input[134]), .B(p_input[518]), .Z(n2510) );
  XOR U2526 ( .A(n2534), .B(n2535), .Z(n2315) );
  AND U2527 ( .A(n23), .B(n2536), .Z(n2535) );
  XNOR U2528 ( .A(n2537), .B(n2534), .Z(n2536) );
  XNOR U2529 ( .A(n2538), .B(n2539), .Z(n23) );
  AND U2530 ( .A(n2540), .B(n2541), .Z(n2539) );
  XOR U2531 ( .A(n2328), .B(n2538), .Z(n2541) );
  AND U2532 ( .A(n2542), .B(n2543), .Z(n2328) );
  XNOR U2533 ( .A(n2325), .B(n2538), .Z(n2540) );
  XNOR U2534 ( .A(n2544), .B(n2545), .Z(n2325) );
  AND U2535 ( .A(n27), .B(n2546), .Z(n2545) );
  XNOR U2536 ( .A(n2547), .B(n2544), .Z(n2546) );
  XOR U2537 ( .A(n2548), .B(n2549), .Z(n2538) );
  AND U2538 ( .A(n2550), .B(n2551), .Z(n2549) );
  XNOR U2539 ( .A(n2548), .B(n2542), .Z(n2551) );
  IV U2540 ( .A(n2343), .Z(n2542) );
  XOR U2541 ( .A(n2552), .B(n2553), .Z(n2343) );
  XOR U2542 ( .A(n2554), .B(n2543), .Z(n2553) );
  AND U2543 ( .A(n2370), .B(n2555), .Z(n2543) );
  AND U2544 ( .A(n2556), .B(n2557), .Z(n2554) );
  XOR U2545 ( .A(n2558), .B(n2552), .Z(n2556) );
  XNOR U2546 ( .A(n2340), .B(n2548), .Z(n2550) );
  XOR U2547 ( .A(n2559), .B(n2560), .Z(n2340) );
  AND U2548 ( .A(n27), .B(n2561), .Z(n2560) );
  XOR U2549 ( .A(n2562), .B(n2559), .Z(n2561) );
  XOR U2550 ( .A(n2563), .B(n2564), .Z(n2548) );
  AND U2551 ( .A(n2565), .B(n2566), .Z(n2564) );
  XNOR U2552 ( .A(n2563), .B(n2370), .Z(n2566) );
  XOR U2553 ( .A(n2567), .B(n2557), .Z(n2370) );
  XNOR U2554 ( .A(n2568), .B(n2552), .Z(n2557) );
  XOR U2555 ( .A(n2569), .B(n2570), .Z(n2552) );
  AND U2556 ( .A(n2571), .B(n2572), .Z(n2570) );
  XOR U2557 ( .A(n2573), .B(n2569), .Z(n2571) );
  XNOR U2558 ( .A(n2574), .B(n2575), .Z(n2568) );
  AND U2559 ( .A(n2576), .B(n2577), .Z(n2575) );
  XOR U2560 ( .A(n2574), .B(n2578), .Z(n2576) );
  XNOR U2561 ( .A(n2558), .B(n2555), .Z(n2567) );
  AND U2562 ( .A(n2579), .B(n2580), .Z(n2555) );
  XOR U2563 ( .A(n2581), .B(n2582), .Z(n2558) );
  AND U2564 ( .A(n2583), .B(n2584), .Z(n2582) );
  XOR U2565 ( .A(n2581), .B(n2585), .Z(n2583) );
  XNOR U2566 ( .A(n2367), .B(n2563), .Z(n2565) );
  XOR U2567 ( .A(n2586), .B(n2587), .Z(n2367) );
  AND U2568 ( .A(n27), .B(n2588), .Z(n2587) );
  XNOR U2569 ( .A(n2589), .B(n2586), .Z(n2588) );
  XOR U2570 ( .A(n2590), .B(n2591), .Z(n2563) );
  AND U2571 ( .A(n2592), .B(n2593), .Z(n2591) );
  XNOR U2572 ( .A(n2590), .B(n2579), .Z(n2593) );
  IV U2573 ( .A(n2418), .Z(n2579) );
  XNOR U2574 ( .A(n2594), .B(n2572), .Z(n2418) );
  XNOR U2575 ( .A(n2595), .B(n2578), .Z(n2572) );
  XOR U2576 ( .A(n2596), .B(n2597), .Z(n2578) );
  AND U2577 ( .A(n2598), .B(n2599), .Z(n2597) );
  XOR U2578 ( .A(n2596), .B(n2600), .Z(n2598) );
  XNOR U2579 ( .A(n2577), .B(n2569), .Z(n2595) );
  XOR U2580 ( .A(n2601), .B(n2602), .Z(n2569) );
  AND U2581 ( .A(n2603), .B(n2604), .Z(n2602) );
  XNOR U2582 ( .A(n2605), .B(n2601), .Z(n2603) );
  XNOR U2583 ( .A(n2606), .B(n2574), .Z(n2577) );
  XOR U2584 ( .A(n2607), .B(n2608), .Z(n2574) );
  AND U2585 ( .A(n2609), .B(n2610), .Z(n2608) );
  XOR U2586 ( .A(n2607), .B(n2611), .Z(n2609) );
  XNOR U2587 ( .A(n2612), .B(n2613), .Z(n2606) );
  AND U2588 ( .A(n2614), .B(n2615), .Z(n2613) );
  XNOR U2589 ( .A(n2612), .B(n2616), .Z(n2614) );
  XNOR U2590 ( .A(n2573), .B(n2580), .Z(n2594) );
  AND U2591 ( .A(n2514), .B(n2617), .Z(n2580) );
  XOR U2592 ( .A(n2585), .B(n2584), .Z(n2573) );
  XNOR U2593 ( .A(n2618), .B(n2581), .Z(n2584) );
  XOR U2594 ( .A(n2619), .B(n2620), .Z(n2581) );
  AND U2595 ( .A(n2621), .B(n2622), .Z(n2620) );
  XOR U2596 ( .A(n2619), .B(n2623), .Z(n2621) );
  XNOR U2597 ( .A(n2624), .B(n2625), .Z(n2618) );
  AND U2598 ( .A(n2626), .B(n2627), .Z(n2625) );
  XOR U2599 ( .A(n2624), .B(n2628), .Z(n2626) );
  XOR U2600 ( .A(n2629), .B(n2630), .Z(n2585) );
  AND U2601 ( .A(n2631), .B(n2632), .Z(n2630) );
  XOR U2602 ( .A(n2629), .B(n2633), .Z(n2631) );
  XNOR U2603 ( .A(n2415), .B(n2590), .Z(n2592) );
  XOR U2604 ( .A(n2634), .B(n2635), .Z(n2415) );
  AND U2605 ( .A(n27), .B(n2636), .Z(n2635) );
  XOR U2606 ( .A(n2637), .B(n2634), .Z(n2636) );
  XOR U2607 ( .A(n2638), .B(n2639), .Z(n2590) );
  AND U2608 ( .A(n2640), .B(n2641), .Z(n2639) );
  XNOR U2609 ( .A(n2638), .B(n2514), .Z(n2641) );
  XOR U2610 ( .A(n2642), .B(n2604), .Z(n2514) );
  XNOR U2611 ( .A(n2643), .B(n2611), .Z(n2604) );
  XOR U2612 ( .A(n2600), .B(n2599), .Z(n2611) );
  XNOR U2613 ( .A(n2644), .B(n2596), .Z(n2599) );
  XOR U2614 ( .A(n2645), .B(n2646), .Z(n2596) );
  AND U2615 ( .A(n2647), .B(n2648), .Z(n2646) );
  XNOR U2616 ( .A(n2649), .B(n2650), .Z(n2647) );
  IV U2617 ( .A(n2645), .Z(n2649) );
  XNOR U2618 ( .A(n2651), .B(n2652), .Z(n2644) );
  NOR U2619 ( .A(n2653), .B(n2654), .Z(n2652) );
  XNOR U2620 ( .A(n2651), .B(n2655), .Z(n2653) );
  XOR U2621 ( .A(n2656), .B(n2657), .Z(n2600) );
  NOR U2622 ( .A(n2658), .B(n2659), .Z(n2657) );
  XNOR U2623 ( .A(n2656), .B(n2660), .Z(n2658) );
  XNOR U2624 ( .A(n2610), .B(n2601), .Z(n2643) );
  XOR U2625 ( .A(n2661), .B(n2662), .Z(n2601) );
  AND U2626 ( .A(n2663), .B(n2664), .Z(n2662) );
  XOR U2627 ( .A(n2661), .B(n2665), .Z(n2663) );
  XOR U2628 ( .A(n2666), .B(n2616), .Z(n2610) );
  XOR U2629 ( .A(n2667), .B(n2668), .Z(n2616) );
  NOR U2630 ( .A(n2669), .B(n2670), .Z(n2668) );
  XOR U2631 ( .A(n2667), .B(n2671), .Z(n2669) );
  XNOR U2632 ( .A(n2615), .B(n2607), .Z(n2666) );
  XOR U2633 ( .A(n2672), .B(n2673), .Z(n2607) );
  AND U2634 ( .A(n2674), .B(n2675), .Z(n2673) );
  XOR U2635 ( .A(n2672), .B(n2676), .Z(n2674) );
  XNOR U2636 ( .A(n2677), .B(n2612), .Z(n2615) );
  XOR U2637 ( .A(n2678), .B(n2679), .Z(n2612) );
  AND U2638 ( .A(n2680), .B(n2681), .Z(n2679) );
  XNOR U2639 ( .A(n2682), .B(n2683), .Z(n2680) );
  IV U2640 ( .A(n2678), .Z(n2682) );
  XNOR U2641 ( .A(n2684), .B(n2685), .Z(n2677) );
  NOR U2642 ( .A(n2686), .B(n2687), .Z(n2685) );
  XNOR U2643 ( .A(n2684), .B(n2688), .Z(n2686) );
  XOR U2644 ( .A(n2605), .B(n2617), .Z(n2642) );
  NOR U2645 ( .A(n2537), .B(n2689), .Z(n2617) );
  XNOR U2646 ( .A(n2623), .B(n2622), .Z(n2605) );
  XNOR U2647 ( .A(n2690), .B(n2628), .Z(n2622) );
  XNOR U2648 ( .A(n2691), .B(n2692), .Z(n2628) );
  NOR U2649 ( .A(n2693), .B(n2694), .Z(n2692) );
  XOR U2650 ( .A(n2691), .B(n2695), .Z(n2693) );
  XNOR U2651 ( .A(n2627), .B(n2619), .Z(n2690) );
  XOR U2652 ( .A(n2696), .B(n2697), .Z(n2619) );
  AND U2653 ( .A(n2698), .B(n2699), .Z(n2697) );
  XOR U2654 ( .A(n2696), .B(n2700), .Z(n2698) );
  XNOR U2655 ( .A(n2701), .B(n2624), .Z(n2627) );
  XOR U2656 ( .A(n2702), .B(n2703), .Z(n2624) );
  AND U2657 ( .A(n2704), .B(n2705), .Z(n2703) );
  XNOR U2658 ( .A(n2706), .B(n2707), .Z(n2704) );
  IV U2659 ( .A(n2702), .Z(n2706) );
  XNOR U2660 ( .A(n2708), .B(n2709), .Z(n2701) );
  NOR U2661 ( .A(n2710), .B(n2711), .Z(n2709) );
  XNOR U2662 ( .A(n2708), .B(n2712), .Z(n2710) );
  XOR U2663 ( .A(n2633), .B(n2632), .Z(n2623) );
  XNOR U2664 ( .A(n2713), .B(n2629), .Z(n2632) );
  XOR U2665 ( .A(n2714), .B(n2715), .Z(n2629) );
  AND U2666 ( .A(n2716), .B(n2717), .Z(n2715) );
  XNOR U2667 ( .A(n2718), .B(n2719), .Z(n2716) );
  IV U2668 ( .A(n2714), .Z(n2718) );
  XNOR U2669 ( .A(n2720), .B(n2721), .Z(n2713) );
  NOR U2670 ( .A(n2722), .B(n2723), .Z(n2721) );
  XNOR U2671 ( .A(n2720), .B(n2724), .Z(n2722) );
  XOR U2672 ( .A(n2725), .B(n2726), .Z(n2633) );
  NOR U2673 ( .A(n2727), .B(n2728), .Z(n2726) );
  XNOR U2674 ( .A(n2725), .B(n2729), .Z(n2727) );
  XNOR U2675 ( .A(n2511), .B(n2638), .Z(n2640) );
  XOR U2676 ( .A(n2730), .B(n2731), .Z(n2511) );
  AND U2677 ( .A(n27), .B(n2732), .Z(n2731) );
  XNOR U2678 ( .A(n2733), .B(n2730), .Z(n2732) );
  AND U2679 ( .A(n2534), .B(n2537), .Z(n2638) );
  XOR U2680 ( .A(n2734), .B(n2689), .Z(n2537) );
  XNOR U2681 ( .A(p_input[160]), .B(p_input[512]), .Z(n2689) );
  XNOR U2682 ( .A(n2665), .B(n2664), .Z(n2734) );
  XNOR U2683 ( .A(n2735), .B(n2676), .Z(n2664) );
  XOR U2684 ( .A(n2650), .B(n2648), .Z(n2676) );
  XNOR U2685 ( .A(n2736), .B(n2655), .Z(n2648) );
  XOR U2686 ( .A(p_input[184]), .B(p_input[536]), .Z(n2655) );
  XOR U2687 ( .A(n2645), .B(n2654), .Z(n2736) );
  XOR U2688 ( .A(n2737), .B(n2651), .Z(n2654) );
  XOR U2689 ( .A(p_input[182]), .B(p_input[534]), .Z(n2651) );
  XOR U2690 ( .A(p_input[183]), .B(n1634), .Z(n2737) );
  XOR U2691 ( .A(p_input[178]), .B(p_input[530]), .Z(n2645) );
  XNOR U2692 ( .A(n2660), .B(n2659), .Z(n2650) );
  XOR U2693 ( .A(n2738), .B(n2656), .Z(n2659) );
  XOR U2694 ( .A(p_input[179]), .B(p_input[531]), .Z(n2656) );
  XOR U2695 ( .A(p_input[180]), .B(n1636), .Z(n2738) );
  XOR U2696 ( .A(p_input[181]), .B(p_input[533]), .Z(n2660) );
  XOR U2697 ( .A(n2675), .B(n2739), .Z(n2735) );
  IV U2698 ( .A(n2661), .Z(n2739) );
  XOR U2699 ( .A(p_input[161]), .B(p_input[513]), .Z(n2661) );
  XNOR U2700 ( .A(n2740), .B(n2683), .Z(n2675) );
  XNOR U2701 ( .A(n2671), .B(n2670), .Z(n2683) );
  XNOR U2702 ( .A(n2741), .B(n2667), .Z(n2670) );
  XNOR U2703 ( .A(p_input[186]), .B(p_input[538]), .Z(n2667) );
  XOR U2704 ( .A(p_input[187]), .B(n1640), .Z(n2741) );
  XOR U2705 ( .A(p_input[188]), .B(p_input[540]), .Z(n2671) );
  XOR U2706 ( .A(n2681), .B(n2742), .Z(n2740) );
  IV U2707 ( .A(n2672), .Z(n2742) );
  XOR U2708 ( .A(p_input[177]), .B(p_input[529]), .Z(n2672) );
  XNOR U2709 ( .A(n2743), .B(n2688), .Z(n2681) );
  XNOR U2710 ( .A(p_input[191]), .B(n1643), .Z(n2688) );
  XOR U2711 ( .A(n2678), .B(n2687), .Z(n2743) );
  XOR U2712 ( .A(n2744), .B(n2684), .Z(n2687) );
  XOR U2713 ( .A(p_input[189]), .B(p_input[541]), .Z(n2684) );
  XOR U2714 ( .A(p_input[190]), .B(n1645), .Z(n2744) );
  XOR U2715 ( .A(p_input[185]), .B(p_input[537]), .Z(n2678) );
  XOR U2716 ( .A(n2700), .B(n2699), .Z(n2665) );
  XNOR U2717 ( .A(n2745), .B(n2707), .Z(n2699) );
  XNOR U2718 ( .A(n2695), .B(n2694), .Z(n2707) );
  XNOR U2719 ( .A(n2746), .B(n2691), .Z(n2694) );
  XNOR U2720 ( .A(p_input[171]), .B(p_input[523]), .Z(n2691) );
  XOR U2721 ( .A(p_input[172]), .B(n1648), .Z(n2746) );
  XOR U2722 ( .A(p_input[173]), .B(p_input[525]), .Z(n2695) );
  XOR U2723 ( .A(n2705), .B(n2747), .Z(n2745) );
  IV U2724 ( .A(n2696), .Z(n2747) );
  XOR U2725 ( .A(p_input[162]), .B(p_input[514]), .Z(n2696) );
  XNOR U2726 ( .A(n2748), .B(n2712), .Z(n2705) );
  XNOR U2727 ( .A(p_input[176]), .B(n1651), .Z(n2712) );
  XOR U2728 ( .A(n2702), .B(n2711), .Z(n2748) );
  XOR U2729 ( .A(n2749), .B(n2708), .Z(n2711) );
  XOR U2730 ( .A(p_input[174]), .B(p_input[526]), .Z(n2708) );
  XOR U2731 ( .A(p_input[175]), .B(n1653), .Z(n2749) );
  XOR U2732 ( .A(p_input[170]), .B(p_input[522]), .Z(n2702) );
  XOR U2733 ( .A(n2719), .B(n2717), .Z(n2700) );
  XNOR U2734 ( .A(n2750), .B(n2724), .Z(n2717) );
  XOR U2735 ( .A(p_input[169]), .B(p_input[521]), .Z(n2724) );
  XOR U2736 ( .A(n2714), .B(n2723), .Z(n2750) );
  XOR U2737 ( .A(n2751), .B(n2720), .Z(n2723) );
  XOR U2738 ( .A(p_input[167]), .B(p_input[519]), .Z(n2720) );
  XOR U2739 ( .A(p_input[168]), .B(n1877), .Z(n2751) );
  XOR U2740 ( .A(p_input[163]), .B(p_input[515]), .Z(n2714) );
  XNOR U2741 ( .A(n2729), .B(n2728), .Z(n2719) );
  XOR U2742 ( .A(n2752), .B(n2725), .Z(n2728) );
  XOR U2743 ( .A(p_input[164]), .B(p_input[516]), .Z(n2725) );
  XOR U2744 ( .A(p_input[165]), .B(n1879), .Z(n2752) );
  XOR U2745 ( .A(p_input[166]), .B(p_input[518]), .Z(n2729) );
  XOR U2746 ( .A(n2753), .B(n2754), .Z(n2534) );
  AND U2747 ( .A(n27), .B(n2755), .Z(n2754) );
  XNOR U2748 ( .A(n2756), .B(n2753), .Z(n2755) );
  XNOR U2749 ( .A(n2757), .B(n2758), .Z(n27) );
  AND U2750 ( .A(n2759), .B(n2760), .Z(n2758) );
  XOR U2751 ( .A(n2547), .B(n2757), .Z(n2760) );
  AND U2752 ( .A(n2761), .B(n2762), .Z(n2547) );
  XNOR U2753 ( .A(n2763), .B(n2757), .Z(n2759) );
  IV U2754 ( .A(n2544), .Z(n2763) );
  XNOR U2755 ( .A(n2764), .B(n2765), .Z(n2544) );
  AND U2756 ( .A(n2766), .B(n31), .Z(n2765) );
  AND U2757 ( .A(n2764), .B(n2767), .Z(n2766) );
  IV U2758 ( .A(n2768), .Z(n2767) );
  XOR U2759 ( .A(n2769), .B(n2770), .Z(n2757) );
  AND U2760 ( .A(n2771), .B(n2772), .Z(n2770) );
  XNOR U2761 ( .A(n2769), .B(n2761), .Z(n2772) );
  IV U2762 ( .A(n2562), .Z(n2761) );
  XOR U2763 ( .A(n2773), .B(n2774), .Z(n2562) );
  XOR U2764 ( .A(n2775), .B(n2762), .Z(n2774) );
  AND U2765 ( .A(n2589), .B(n2776), .Z(n2762) );
  AND U2766 ( .A(n2777), .B(n2778), .Z(n2775) );
  XOR U2767 ( .A(n2779), .B(n2773), .Z(n2777) );
  XNOR U2768 ( .A(n2559), .B(n2769), .Z(n2771) );
  XOR U2769 ( .A(n2780), .B(n2781), .Z(n2559) );
  AND U2770 ( .A(n31), .B(n2782), .Z(n2781) );
  XOR U2771 ( .A(n2783), .B(n2780), .Z(n2782) );
  XOR U2772 ( .A(n2784), .B(n2785), .Z(n2769) );
  AND U2773 ( .A(n2786), .B(n2787), .Z(n2785) );
  XNOR U2774 ( .A(n2784), .B(n2589), .Z(n2787) );
  XOR U2775 ( .A(n2788), .B(n2778), .Z(n2589) );
  XNOR U2776 ( .A(n2789), .B(n2773), .Z(n2778) );
  XOR U2777 ( .A(n2790), .B(n2791), .Z(n2773) );
  AND U2778 ( .A(n2792), .B(n2793), .Z(n2791) );
  XOR U2779 ( .A(n2794), .B(n2790), .Z(n2792) );
  XNOR U2780 ( .A(n2795), .B(n2796), .Z(n2789) );
  AND U2781 ( .A(n2797), .B(n2798), .Z(n2796) );
  XOR U2782 ( .A(n2795), .B(n2799), .Z(n2797) );
  XNOR U2783 ( .A(n2779), .B(n2776), .Z(n2788) );
  AND U2784 ( .A(n2800), .B(n2801), .Z(n2776) );
  XOR U2785 ( .A(n2802), .B(n2803), .Z(n2779) );
  AND U2786 ( .A(n2804), .B(n2805), .Z(n2803) );
  XOR U2787 ( .A(n2802), .B(n2806), .Z(n2804) );
  XNOR U2788 ( .A(n2586), .B(n2784), .Z(n2786) );
  XOR U2789 ( .A(n2807), .B(n2808), .Z(n2586) );
  AND U2790 ( .A(n31), .B(n2809), .Z(n2808) );
  XNOR U2791 ( .A(n2810), .B(n2807), .Z(n2809) );
  XOR U2792 ( .A(n2811), .B(n2812), .Z(n2784) );
  AND U2793 ( .A(n2813), .B(n2814), .Z(n2812) );
  XNOR U2794 ( .A(n2811), .B(n2800), .Z(n2814) );
  IV U2795 ( .A(n2637), .Z(n2800) );
  XNOR U2796 ( .A(n2815), .B(n2793), .Z(n2637) );
  XNOR U2797 ( .A(n2816), .B(n2799), .Z(n2793) );
  XOR U2798 ( .A(n2817), .B(n2818), .Z(n2799) );
  AND U2799 ( .A(n2819), .B(n2820), .Z(n2818) );
  XOR U2800 ( .A(n2817), .B(n2821), .Z(n2819) );
  XNOR U2801 ( .A(n2798), .B(n2790), .Z(n2816) );
  XOR U2802 ( .A(n2822), .B(n2823), .Z(n2790) );
  AND U2803 ( .A(n2824), .B(n2825), .Z(n2823) );
  XNOR U2804 ( .A(n2826), .B(n2822), .Z(n2824) );
  XNOR U2805 ( .A(n2827), .B(n2795), .Z(n2798) );
  XOR U2806 ( .A(n2828), .B(n2829), .Z(n2795) );
  AND U2807 ( .A(n2830), .B(n2831), .Z(n2829) );
  XOR U2808 ( .A(n2828), .B(n2832), .Z(n2830) );
  XNOR U2809 ( .A(n2833), .B(n2834), .Z(n2827) );
  AND U2810 ( .A(n2835), .B(n2836), .Z(n2834) );
  XNOR U2811 ( .A(n2833), .B(n2837), .Z(n2835) );
  XNOR U2812 ( .A(n2794), .B(n2801), .Z(n2815) );
  AND U2813 ( .A(n2733), .B(n2838), .Z(n2801) );
  XOR U2814 ( .A(n2806), .B(n2805), .Z(n2794) );
  XNOR U2815 ( .A(n2839), .B(n2802), .Z(n2805) );
  XOR U2816 ( .A(n2840), .B(n2841), .Z(n2802) );
  AND U2817 ( .A(n2842), .B(n2843), .Z(n2841) );
  XOR U2818 ( .A(n2840), .B(n2844), .Z(n2842) );
  XNOR U2819 ( .A(n2845), .B(n2846), .Z(n2839) );
  AND U2820 ( .A(n2847), .B(n2848), .Z(n2846) );
  XOR U2821 ( .A(n2845), .B(n2849), .Z(n2847) );
  XOR U2822 ( .A(n2850), .B(n2851), .Z(n2806) );
  AND U2823 ( .A(n2852), .B(n2853), .Z(n2851) );
  XOR U2824 ( .A(n2850), .B(n2854), .Z(n2852) );
  XNOR U2825 ( .A(n2634), .B(n2811), .Z(n2813) );
  XOR U2826 ( .A(n2855), .B(n2856), .Z(n2634) );
  AND U2827 ( .A(n31), .B(n2857), .Z(n2856) );
  XOR U2828 ( .A(n2858), .B(n2855), .Z(n2857) );
  XOR U2829 ( .A(n2859), .B(n2860), .Z(n2811) );
  AND U2830 ( .A(n2861), .B(n2862), .Z(n2860) );
  XNOR U2831 ( .A(n2859), .B(n2733), .Z(n2862) );
  XOR U2832 ( .A(n2863), .B(n2825), .Z(n2733) );
  XNOR U2833 ( .A(n2864), .B(n2832), .Z(n2825) );
  XOR U2834 ( .A(n2821), .B(n2820), .Z(n2832) );
  XNOR U2835 ( .A(n2865), .B(n2817), .Z(n2820) );
  XOR U2836 ( .A(n2866), .B(n2867), .Z(n2817) );
  AND U2837 ( .A(n2868), .B(n2869), .Z(n2867) );
  XNOR U2838 ( .A(n2870), .B(n2871), .Z(n2868) );
  IV U2839 ( .A(n2866), .Z(n2870) );
  XNOR U2840 ( .A(n2872), .B(n2873), .Z(n2865) );
  NOR U2841 ( .A(n2874), .B(n2875), .Z(n2873) );
  XNOR U2842 ( .A(n2872), .B(n2876), .Z(n2874) );
  XOR U2843 ( .A(n2877), .B(n2878), .Z(n2821) );
  NOR U2844 ( .A(n2879), .B(n2880), .Z(n2878) );
  XNOR U2845 ( .A(n2877), .B(n2881), .Z(n2879) );
  XNOR U2846 ( .A(n2831), .B(n2822), .Z(n2864) );
  XOR U2847 ( .A(n2882), .B(n2883), .Z(n2822) );
  AND U2848 ( .A(n2884), .B(n2885), .Z(n2883) );
  XOR U2849 ( .A(n2882), .B(n2886), .Z(n2884) );
  XOR U2850 ( .A(n2887), .B(n2837), .Z(n2831) );
  XOR U2851 ( .A(n2888), .B(n2889), .Z(n2837) );
  NOR U2852 ( .A(n2890), .B(n2891), .Z(n2889) );
  XOR U2853 ( .A(n2888), .B(n2892), .Z(n2890) );
  XNOR U2854 ( .A(n2836), .B(n2828), .Z(n2887) );
  XOR U2855 ( .A(n2893), .B(n2894), .Z(n2828) );
  AND U2856 ( .A(n2895), .B(n2896), .Z(n2894) );
  XOR U2857 ( .A(n2893), .B(n2897), .Z(n2895) );
  XNOR U2858 ( .A(n2898), .B(n2833), .Z(n2836) );
  XOR U2859 ( .A(n2899), .B(n2900), .Z(n2833) );
  AND U2860 ( .A(n2901), .B(n2902), .Z(n2900) );
  XNOR U2861 ( .A(n2903), .B(n2904), .Z(n2901) );
  IV U2862 ( .A(n2899), .Z(n2903) );
  XNOR U2863 ( .A(n2905), .B(n2906), .Z(n2898) );
  NOR U2864 ( .A(n2907), .B(n2908), .Z(n2906) );
  XNOR U2865 ( .A(n2905), .B(n2909), .Z(n2907) );
  XOR U2866 ( .A(n2826), .B(n2838), .Z(n2863) );
  NOR U2867 ( .A(n2756), .B(n2910), .Z(n2838) );
  XNOR U2868 ( .A(n2844), .B(n2843), .Z(n2826) );
  XNOR U2869 ( .A(n2911), .B(n2849), .Z(n2843) );
  XNOR U2870 ( .A(n2912), .B(n2913), .Z(n2849) );
  NOR U2871 ( .A(n2914), .B(n2915), .Z(n2913) );
  XOR U2872 ( .A(n2912), .B(n2916), .Z(n2914) );
  XNOR U2873 ( .A(n2848), .B(n2840), .Z(n2911) );
  XOR U2874 ( .A(n2917), .B(n2918), .Z(n2840) );
  AND U2875 ( .A(n2919), .B(n2920), .Z(n2918) );
  XOR U2876 ( .A(n2917), .B(n2921), .Z(n2919) );
  XNOR U2877 ( .A(n2922), .B(n2845), .Z(n2848) );
  XOR U2878 ( .A(n2923), .B(n2924), .Z(n2845) );
  AND U2879 ( .A(n2925), .B(n2926), .Z(n2924) );
  XNOR U2880 ( .A(n2927), .B(n2928), .Z(n2925) );
  IV U2881 ( .A(n2923), .Z(n2927) );
  XNOR U2882 ( .A(n2929), .B(n2930), .Z(n2922) );
  NOR U2883 ( .A(n2931), .B(n2932), .Z(n2930) );
  XNOR U2884 ( .A(n2929), .B(n2933), .Z(n2931) );
  XOR U2885 ( .A(n2854), .B(n2853), .Z(n2844) );
  XNOR U2886 ( .A(n2934), .B(n2850), .Z(n2853) );
  XOR U2887 ( .A(n2935), .B(n2936), .Z(n2850) );
  AND U2888 ( .A(n2937), .B(n2938), .Z(n2936) );
  XNOR U2889 ( .A(n2939), .B(n2940), .Z(n2937) );
  IV U2890 ( .A(n2935), .Z(n2939) );
  XNOR U2891 ( .A(n2941), .B(n2942), .Z(n2934) );
  NOR U2892 ( .A(n2943), .B(n2944), .Z(n2942) );
  XNOR U2893 ( .A(n2941), .B(n2945), .Z(n2943) );
  XOR U2894 ( .A(n2946), .B(n2947), .Z(n2854) );
  NOR U2895 ( .A(n2948), .B(n2949), .Z(n2947) );
  XNOR U2896 ( .A(n2946), .B(n2950), .Z(n2948) );
  XNOR U2897 ( .A(n2730), .B(n2859), .Z(n2861) );
  XOR U2898 ( .A(n2951), .B(n2952), .Z(n2730) );
  AND U2899 ( .A(n31), .B(n2953), .Z(n2952) );
  XNOR U2900 ( .A(n2954), .B(n2951), .Z(n2953) );
  AND U2901 ( .A(n2753), .B(n2756), .Z(n2859) );
  XOR U2902 ( .A(n2955), .B(n2910), .Z(n2756) );
  XNOR U2903 ( .A(p_input[192]), .B(p_input[512]), .Z(n2910) );
  XNOR U2904 ( .A(n2886), .B(n2885), .Z(n2955) );
  XNOR U2905 ( .A(n2956), .B(n2897), .Z(n2885) );
  XOR U2906 ( .A(n2871), .B(n2869), .Z(n2897) );
  XNOR U2907 ( .A(n2957), .B(n2876), .Z(n2869) );
  XOR U2908 ( .A(p_input[216]), .B(p_input[536]), .Z(n2876) );
  XOR U2909 ( .A(n2866), .B(n2875), .Z(n2957) );
  XOR U2910 ( .A(n2958), .B(n2872), .Z(n2875) );
  XOR U2911 ( .A(p_input[214]), .B(p_input[534]), .Z(n2872) );
  XOR U2912 ( .A(p_input[215]), .B(n1634), .Z(n2958) );
  XOR U2913 ( .A(p_input[210]), .B(p_input[530]), .Z(n2866) );
  XNOR U2914 ( .A(n2881), .B(n2880), .Z(n2871) );
  XOR U2915 ( .A(n2959), .B(n2877), .Z(n2880) );
  XOR U2916 ( .A(p_input[211]), .B(p_input[531]), .Z(n2877) );
  XOR U2917 ( .A(p_input[212]), .B(n1636), .Z(n2959) );
  XOR U2918 ( .A(p_input[213]), .B(p_input[533]), .Z(n2881) );
  XOR U2919 ( .A(n2896), .B(n2960), .Z(n2956) );
  IV U2920 ( .A(n2882), .Z(n2960) );
  XOR U2921 ( .A(p_input[193]), .B(p_input[513]), .Z(n2882) );
  XNOR U2922 ( .A(n2961), .B(n2904), .Z(n2896) );
  XNOR U2923 ( .A(n2892), .B(n2891), .Z(n2904) );
  XNOR U2924 ( .A(n2962), .B(n2888), .Z(n2891) );
  XNOR U2925 ( .A(p_input[218]), .B(p_input[538]), .Z(n2888) );
  XOR U2926 ( .A(p_input[219]), .B(n1640), .Z(n2962) );
  XOR U2927 ( .A(p_input[220]), .B(p_input[540]), .Z(n2892) );
  XOR U2928 ( .A(n2902), .B(n2963), .Z(n2961) );
  IV U2929 ( .A(n2893), .Z(n2963) );
  XOR U2930 ( .A(p_input[209]), .B(p_input[529]), .Z(n2893) );
  XNOR U2931 ( .A(n2964), .B(n2909), .Z(n2902) );
  XNOR U2932 ( .A(p_input[223]), .B(n1643), .Z(n2909) );
  XOR U2933 ( .A(n2899), .B(n2908), .Z(n2964) );
  XOR U2934 ( .A(n2965), .B(n2905), .Z(n2908) );
  XOR U2935 ( .A(p_input[221]), .B(p_input[541]), .Z(n2905) );
  XOR U2936 ( .A(p_input[222]), .B(n1645), .Z(n2965) );
  XOR U2937 ( .A(p_input[217]), .B(p_input[537]), .Z(n2899) );
  XOR U2938 ( .A(n2921), .B(n2920), .Z(n2886) );
  XNOR U2939 ( .A(n2966), .B(n2928), .Z(n2920) );
  XNOR U2940 ( .A(n2916), .B(n2915), .Z(n2928) );
  XNOR U2941 ( .A(n2967), .B(n2912), .Z(n2915) );
  XNOR U2942 ( .A(p_input[203]), .B(p_input[523]), .Z(n2912) );
  XOR U2943 ( .A(p_input[204]), .B(n1648), .Z(n2967) );
  XOR U2944 ( .A(p_input[205]), .B(p_input[525]), .Z(n2916) );
  XOR U2945 ( .A(n2926), .B(n2968), .Z(n2966) );
  IV U2946 ( .A(n2917), .Z(n2968) );
  XOR U2947 ( .A(p_input[194]), .B(p_input[514]), .Z(n2917) );
  XNOR U2948 ( .A(n2969), .B(n2933), .Z(n2926) );
  XNOR U2949 ( .A(p_input[208]), .B(n1651), .Z(n2933) );
  XOR U2950 ( .A(n2923), .B(n2932), .Z(n2969) );
  XOR U2951 ( .A(n2970), .B(n2929), .Z(n2932) );
  XOR U2952 ( .A(p_input[206]), .B(p_input[526]), .Z(n2929) );
  XOR U2953 ( .A(p_input[207]), .B(n1653), .Z(n2970) );
  XOR U2954 ( .A(p_input[202]), .B(p_input[522]), .Z(n2923) );
  XOR U2955 ( .A(n2940), .B(n2938), .Z(n2921) );
  XNOR U2956 ( .A(n2971), .B(n2945), .Z(n2938) );
  XOR U2957 ( .A(p_input[201]), .B(p_input[521]), .Z(n2945) );
  XOR U2958 ( .A(n2935), .B(n2944), .Z(n2971) );
  XOR U2959 ( .A(n2972), .B(n2941), .Z(n2944) );
  XOR U2960 ( .A(p_input[199]), .B(p_input[519]), .Z(n2941) );
  XOR U2961 ( .A(p_input[200]), .B(n1877), .Z(n2972) );
  XOR U2962 ( .A(p_input[195]), .B(p_input[515]), .Z(n2935) );
  XNOR U2963 ( .A(n2950), .B(n2949), .Z(n2940) );
  XOR U2964 ( .A(n2973), .B(n2946), .Z(n2949) );
  XOR U2965 ( .A(p_input[196]), .B(p_input[516]), .Z(n2946) );
  XOR U2966 ( .A(p_input[197]), .B(n1879), .Z(n2973) );
  XOR U2967 ( .A(p_input[198]), .B(p_input[518]), .Z(n2950) );
  XOR U2968 ( .A(n2974), .B(n2975), .Z(n2753) );
  AND U2969 ( .A(n31), .B(n2976), .Z(n2975) );
  XNOR U2970 ( .A(n2977), .B(n2974), .Z(n2976) );
  XNOR U2971 ( .A(n2978), .B(n2979), .Z(n31) );
  NOR U2972 ( .A(n2980), .B(n2981), .Z(n2979) );
  XOR U2973 ( .A(n2764), .B(n2978), .Z(n2981) );
  AND U2974 ( .A(n2982), .B(n2983), .Z(n2764) );
  NOR U2975 ( .A(n2978), .B(n2768), .Z(n2980) );
  AND U2976 ( .A(n2984), .B(n2985), .Z(n2768) );
  XOR U2977 ( .A(n2986), .B(n2987), .Z(n2978) );
  AND U2978 ( .A(n2988), .B(n2989), .Z(n2987) );
  XNOR U2979 ( .A(n2986), .B(n2984), .Z(n2989) );
  IV U2980 ( .A(n2783), .Z(n2984) );
  XOR U2981 ( .A(n2990), .B(n2991), .Z(n2783) );
  XOR U2982 ( .A(n2992), .B(n2985), .Z(n2991) );
  AND U2983 ( .A(n2810), .B(n2993), .Z(n2985) );
  AND U2984 ( .A(n2994), .B(n2995), .Z(n2992) );
  XOR U2985 ( .A(n2996), .B(n2990), .Z(n2994) );
  XNOR U2986 ( .A(n2780), .B(n2986), .Z(n2988) );
  XOR U2987 ( .A(n2997), .B(n2998), .Z(n2780) );
  AND U2988 ( .A(n35), .B(n2999), .Z(n2998) );
  XOR U2989 ( .A(n3000), .B(n2997), .Z(n2999) );
  XOR U2990 ( .A(n3001), .B(n3002), .Z(n2986) );
  AND U2991 ( .A(n3003), .B(n3004), .Z(n3002) );
  XNOR U2992 ( .A(n3001), .B(n2810), .Z(n3004) );
  XOR U2993 ( .A(n3005), .B(n2995), .Z(n2810) );
  XNOR U2994 ( .A(n3006), .B(n2990), .Z(n2995) );
  XOR U2995 ( .A(n3007), .B(n3008), .Z(n2990) );
  AND U2996 ( .A(n3009), .B(n3010), .Z(n3008) );
  XOR U2997 ( .A(n3011), .B(n3007), .Z(n3009) );
  XNOR U2998 ( .A(n3012), .B(n3013), .Z(n3006) );
  AND U2999 ( .A(n3014), .B(n3015), .Z(n3013) );
  XOR U3000 ( .A(n3012), .B(n3016), .Z(n3014) );
  XNOR U3001 ( .A(n2996), .B(n2993), .Z(n3005) );
  AND U3002 ( .A(n3017), .B(n3018), .Z(n2993) );
  XOR U3003 ( .A(n3019), .B(n3020), .Z(n2996) );
  AND U3004 ( .A(n3021), .B(n3022), .Z(n3020) );
  XOR U3005 ( .A(n3019), .B(n3023), .Z(n3021) );
  XNOR U3006 ( .A(n2807), .B(n3001), .Z(n3003) );
  XOR U3007 ( .A(n3024), .B(n3025), .Z(n2807) );
  AND U3008 ( .A(n35), .B(n3026), .Z(n3025) );
  XNOR U3009 ( .A(n3027), .B(n3024), .Z(n3026) );
  XOR U3010 ( .A(n3028), .B(n3029), .Z(n3001) );
  AND U3011 ( .A(n3030), .B(n3031), .Z(n3029) );
  XNOR U3012 ( .A(n3028), .B(n3017), .Z(n3031) );
  IV U3013 ( .A(n2858), .Z(n3017) );
  XNOR U3014 ( .A(n3032), .B(n3010), .Z(n2858) );
  XNOR U3015 ( .A(n3033), .B(n3016), .Z(n3010) );
  XOR U3016 ( .A(n3034), .B(n3035), .Z(n3016) );
  AND U3017 ( .A(n3036), .B(n3037), .Z(n3035) );
  XOR U3018 ( .A(n3034), .B(n3038), .Z(n3036) );
  XNOR U3019 ( .A(n3015), .B(n3007), .Z(n3033) );
  XOR U3020 ( .A(n3039), .B(n3040), .Z(n3007) );
  AND U3021 ( .A(n3041), .B(n3042), .Z(n3040) );
  XNOR U3022 ( .A(n3043), .B(n3039), .Z(n3041) );
  XNOR U3023 ( .A(n3044), .B(n3012), .Z(n3015) );
  XOR U3024 ( .A(n3045), .B(n3046), .Z(n3012) );
  AND U3025 ( .A(n3047), .B(n3048), .Z(n3046) );
  XOR U3026 ( .A(n3045), .B(n3049), .Z(n3047) );
  XNOR U3027 ( .A(n3050), .B(n3051), .Z(n3044) );
  AND U3028 ( .A(n3052), .B(n3053), .Z(n3051) );
  XNOR U3029 ( .A(n3050), .B(n3054), .Z(n3052) );
  XNOR U3030 ( .A(n3011), .B(n3018), .Z(n3032) );
  AND U3031 ( .A(n2954), .B(n3055), .Z(n3018) );
  XOR U3032 ( .A(n3023), .B(n3022), .Z(n3011) );
  XNOR U3033 ( .A(n3056), .B(n3019), .Z(n3022) );
  XOR U3034 ( .A(n3057), .B(n3058), .Z(n3019) );
  AND U3035 ( .A(n3059), .B(n3060), .Z(n3058) );
  XOR U3036 ( .A(n3057), .B(n3061), .Z(n3059) );
  XNOR U3037 ( .A(n3062), .B(n3063), .Z(n3056) );
  AND U3038 ( .A(n3064), .B(n3065), .Z(n3063) );
  XOR U3039 ( .A(n3062), .B(n3066), .Z(n3064) );
  XOR U3040 ( .A(n3067), .B(n3068), .Z(n3023) );
  AND U3041 ( .A(n3069), .B(n3070), .Z(n3068) );
  XOR U3042 ( .A(n3067), .B(n3071), .Z(n3069) );
  XNOR U3043 ( .A(n2855), .B(n3028), .Z(n3030) );
  XOR U3044 ( .A(n3072), .B(n3073), .Z(n2855) );
  AND U3045 ( .A(n35), .B(n3074), .Z(n3073) );
  XOR U3046 ( .A(n3075), .B(n3072), .Z(n3074) );
  XOR U3047 ( .A(n3076), .B(n3077), .Z(n3028) );
  AND U3048 ( .A(n3078), .B(n3079), .Z(n3077) );
  XNOR U3049 ( .A(n3076), .B(n2954), .Z(n3079) );
  XOR U3050 ( .A(n3080), .B(n3042), .Z(n2954) );
  XNOR U3051 ( .A(n3081), .B(n3049), .Z(n3042) );
  XOR U3052 ( .A(n3038), .B(n3037), .Z(n3049) );
  XNOR U3053 ( .A(n3082), .B(n3034), .Z(n3037) );
  XOR U3054 ( .A(n3083), .B(n3084), .Z(n3034) );
  AND U3055 ( .A(n3085), .B(n3086), .Z(n3084) );
  XNOR U3056 ( .A(n3087), .B(n3088), .Z(n3085) );
  IV U3057 ( .A(n3083), .Z(n3087) );
  XNOR U3058 ( .A(n3089), .B(n3090), .Z(n3082) );
  NOR U3059 ( .A(n3091), .B(n3092), .Z(n3090) );
  XNOR U3060 ( .A(n3089), .B(n3093), .Z(n3091) );
  XOR U3061 ( .A(n3094), .B(n3095), .Z(n3038) );
  NOR U3062 ( .A(n3096), .B(n3097), .Z(n3095) );
  XNOR U3063 ( .A(n3094), .B(n3098), .Z(n3096) );
  XNOR U3064 ( .A(n3048), .B(n3039), .Z(n3081) );
  XOR U3065 ( .A(n3099), .B(n3100), .Z(n3039) );
  AND U3066 ( .A(n3101), .B(n3102), .Z(n3100) );
  XOR U3067 ( .A(n3099), .B(n3103), .Z(n3101) );
  XOR U3068 ( .A(n3104), .B(n3054), .Z(n3048) );
  XOR U3069 ( .A(n3105), .B(n3106), .Z(n3054) );
  NOR U3070 ( .A(n3107), .B(n3108), .Z(n3106) );
  XOR U3071 ( .A(n3105), .B(n3109), .Z(n3107) );
  XNOR U3072 ( .A(n3053), .B(n3045), .Z(n3104) );
  XOR U3073 ( .A(n3110), .B(n3111), .Z(n3045) );
  AND U3074 ( .A(n3112), .B(n3113), .Z(n3111) );
  XOR U3075 ( .A(n3110), .B(n3114), .Z(n3112) );
  XNOR U3076 ( .A(n3115), .B(n3050), .Z(n3053) );
  XOR U3077 ( .A(n3116), .B(n3117), .Z(n3050) );
  AND U3078 ( .A(n3118), .B(n3119), .Z(n3117) );
  XNOR U3079 ( .A(n3120), .B(n3121), .Z(n3118) );
  IV U3080 ( .A(n3116), .Z(n3120) );
  XNOR U3081 ( .A(n3122), .B(n3123), .Z(n3115) );
  NOR U3082 ( .A(n3124), .B(n3125), .Z(n3123) );
  XNOR U3083 ( .A(n3122), .B(n3126), .Z(n3124) );
  XOR U3084 ( .A(n3043), .B(n3055), .Z(n3080) );
  NOR U3085 ( .A(n2977), .B(n3127), .Z(n3055) );
  XNOR U3086 ( .A(n3061), .B(n3060), .Z(n3043) );
  XNOR U3087 ( .A(n3128), .B(n3066), .Z(n3060) );
  XNOR U3088 ( .A(n3129), .B(n3130), .Z(n3066) );
  NOR U3089 ( .A(n3131), .B(n3132), .Z(n3130) );
  XOR U3090 ( .A(n3129), .B(n3133), .Z(n3131) );
  XNOR U3091 ( .A(n3065), .B(n3057), .Z(n3128) );
  XOR U3092 ( .A(n3134), .B(n3135), .Z(n3057) );
  AND U3093 ( .A(n3136), .B(n3137), .Z(n3135) );
  XOR U3094 ( .A(n3134), .B(n3138), .Z(n3136) );
  XNOR U3095 ( .A(n3139), .B(n3062), .Z(n3065) );
  XOR U3096 ( .A(n3140), .B(n3141), .Z(n3062) );
  AND U3097 ( .A(n3142), .B(n3143), .Z(n3141) );
  XNOR U3098 ( .A(n3144), .B(n3145), .Z(n3142) );
  IV U3099 ( .A(n3140), .Z(n3144) );
  XNOR U3100 ( .A(n3146), .B(n3147), .Z(n3139) );
  NOR U3101 ( .A(n3148), .B(n3149), .Z(n3147) );
  XNOR U3102 ( .A(n3146), .B(n3150), .Z(n3148) );
  XOR U3103 ( .A(n3071), .B(n3070), .Z(n3061) );
  XNOR U3104 ( .A(n3151), .B(n3067), .Z(n3070) );
  XOR U3105 ( .A(n3152), .B(n3153), .Z(n3067) );
  AND U3106 ( .A(n3154), .B(n3155), .Z(n3153) );
  XNOR U3107 ( .A(n3156), .B(n3157), .Z(n3154) );
  IV U3108 ( .A(n3152), .Z(n3156) );
  XNOR U3109 ( .A(n3158), .B(n3159), .Z(n3151) );
  NOR U3110 ( .A(n3160), .B(n3161), .Z(n3159) );
  XNOR U3111 ( .A(n3158), .B(n3162), .Z(n3160) );
  XOR U3112 ( .A(n3163), .B(n3164), .Z(n3071) );
  NOR U3113 ( .A(n3165), .B(n3166), .Z(n3164) );
  XNOR U3114 ( .A(n3163), .B(n3167), .Z(n3165) );
  XNOR U3115 ( .A(n2951), .B(n3076), .Z(n3078) );
  XOR U3116 ( .A(n3168), .B(n3169), .Z(n2951) );
  AND U3117 ( .A(n35), .B(n3170), .Z(n3169) );
  XNOR U3118 ( .A(n3171), .B(n3168), .Z(n3170) );
  AND U3119 ( .A(n2974), .B(n2977), .Z(n3076) );
  XOR U3120 ( .A(n3172), .B(n3127), .Z(n2977) );
  XNOR U3121 ( .A(p_input[224]), .B(p_input[512]), .Z(n3127) );
  XNOR U3122 ( .A(n3103), .B(n3102), .Z(n3172) );
  XNOR U3123 ( .A(n3173), .B(n3114), .Z(n3102) );
  XOR U3124 ( .A(n3088), .B(n3086), .Z(n3114) );
  XNOR U3125 ( .A(n3174), .B(n3093), .Z(n3086) );
  XOR U3126 ( .A(p_input[248]), .B(p_input[536]), .Z(n3093) );
  XOR U3127 ( .A(n3083), .B(n3092), .Z(n3174) );
  XOR U3128 ( .A(n3175), .B(n3089), .Z(n3092) );
  XOR U3129 ( .A(p_input[246]), .B(p_input[534]), .Z(n3089) );
  XOR U3130 ( .A(p_input[247]), .B(n1634), .Z(n3175) );
  XOR U3131 ( .A(p_input[242]), .B(p_input[530]), .Z(n3083) );
  XNOR U3132 ( .A(n3098), .B(n3097), .Z(n3088) );
  XOR U3133 ( .A(n3176), .B(n3094), .Z(n3097) );
  XOR U3134 ( .A(p_input[243]), .B(p_input[531]), .Z(n3094) );
  XOR U3135 ( .A(p_input[244]), .B(n1636), .Z(n3176) );
  XOR U3136 ( .A(p_input[245]), .B(p_input[533]), .Z(n3098) );
  XOR U3137 ( .A(n3113), .B(n3177), .Z(n3173) );
  IV U3138 ( .A(n3099), .Z(n3177) );
  XOR U3139 ( .A(p_input[225]), .B(p_input[513]), .Z(n3099) );
  XNOR U3140 ( .A(n3178), .B(n3121), .Z(n3113) );
  XNOR U3141 ( .A(n3109), .B(n3108), .Z(n3121) );
  XNOR U3142 ( .A(n3179), .B(n3105), .Z(n3108) );
  XNOR U3143 ( .A(p_input[250]), .B(p_input[538]), .Z(n3105) );
  XOR U3144 ( .A(p_input[251]), .B(n1640), .Z(n3179) );
  XOR U3145 ( .A(p_input[252]), .B(p_input[540]), .Z(n3109) );
  XOR U3146 ( .A(n3119), .B(n3180), .Z(n3178) );
  IV U3147 ( .A(n3110), .Z(n3180) );
  XOR U3148 ( .A(p_input[241]), .B(p_input[529]), .Z(n3110) );
  XNOR U3149 ( .A(n3181), .B(n3126), .Z(n3119) );
  XNOR U3150 ( .A(p_input[255]), .B(n1643), .Z(n3126) );
  XOR U3151 ( .A(n3116), .B(n3125), .Z(n3181) );
  XOR U3152 ( .A(n3182), .B(n3122), .Z(n3125) );
  XOR U3153 ( .A(p_input[253]), .B(p_input[541]), .Z(n3122) );
  XOR U3154 ( .A(p_input[254]), .B(n1645), .Z(n3182) );
  XOR U3155 ( .A(p_input[249]), .B(p_input[537]), .Z(n3116) );
  XOR U3156 ( .A(n3138), .B(n3137), .Z(n3103) );
  XNOR U3157 ( .A(n3183), .B(n3145), .Z(n3137) );
  XNOR U3158 ( .A(n3133), .B(n3132), .Z(n3145) );
  XNOR U3159 ( .A(n3184), .B(n3129), .Z(n3132) );
  XNOR U3160 ( .A(p_input[235]), .B(p_input[523]), .Z(n3129) );
  XOR U3161 ( .A(p_input[236]), .B(n1648), .Z(n3184) );
  XOR U3162 ( .A(p_input[237]), .B(p_input[525]), .Z(n3133) );
  XOR U3163 ( .A(n3143), .B(n3185), .Z(n3183) );
  IV U3164 ( .A(n3134), .Z(n3185) );
  XOR U3165 ( .A(p_input[226]), .B(p_input[514]), .Z(n3134) );
  XNOR U3166 ( .A(n3186), .B(n3150), .Z(n3143) );
  XNOR U3167 ( .A(p_input[240]), .B(n1651), .Z(n3150) );
  XOR U3168 ( .A(n3140), .B(n3149), .Z(n3186) );
  XOR U3169 ( .A(n3187), .B(n3146), .Z(n3149) );
  XOR U3170 ( .A(p_input[238]), .B(p_input[526]), .Z(n3146) );
  XOR U3171 ( .A(p_input[239]), .B(n1653), .Z(n3187) );
  XOR U3172 ( .A(p_input[234]), .B(p_input[522]), .Z(n3140) );
  XOR U3173 ( .A(n3157), .B(n3155), .Z(n3138) );
  XNOR U3174 ( .A(n3188), .B(n3162), .Z(n3155) );
  XOR U3175 ( .A(p_input[233]), .B(p_input[521]), .Z(n3162) );
  XOR U3176 ( .A(n3152), .B(n3161), .Z(n3188) );
  XOR U3177 ( .A(n3189), .B(n3158), .Z(n3161) );
  XOR U3178 ( .A(p_input[231]), .B(p_input[519]), .Z(n3158) );
  XOR U3179 ( .A(p_input[232]), .B(n1877), .Z(n3189) );
  XOR U3180 ( .A(p_input[227]), .B(p_input[515]), .Z(n3152) );
  XNOR U3181 ( .A(n3167), .B(n3166), .Z(n3157) );
  XOR U3182 ( .A(n3190), .B(n3163), .Z(n3166) );
  XOR U3183 ( .A(p_input[228]), .B(p_input[516]), .Z(n3163) );
  XOR U3184 ( .A(p_input[229]), .B(n1879), .Z(n3190) );
  XOR U3185 ( .A(p_input[230]), .B(p_input[518]), .Z(n3167) );
  XOR U3186 ( .A(n3191), .B(n3192), .Z(n2974) );
  AND U3187 ( .A(n35), .B(n3193), .Z(n3192) );
  XNOR U3188 ( .A(n3194), .B(n3191), .Z(n3193) );
  XNOR U3189 ( .A(n3195), .B(n3196), .Z(n35) );
  NOR U3190 ( .A(n3197), .B(n3198), .Z(n3196) );
  XOR U3191 ( .A(n2983), .B(n3195), .Z(n3198) );
  AND U3192 ( .A(n3199), .B(n3200), .Z(n2983) );
  NOR U3193 ( .A(n3195), .B(n2982), .Z(n3197) );
  AND U3194 ( .A(n3201), .B(n3202), .Z(n2982) );
  XOR U3195 ( .A(n3203), .B(n3204), .Z(n3195) );
  AND U3196 ( .A(n3205), .B(n3206), .Z(n3204) );
  XNOR U3197 ( .A(n3203), .B(n3201), .Z(n3206) );
  IV U3198 ( .A(n3000), .Z(n3201) );
  XOR U3199 ( .A(n3207), .B(n3208), .Z(n3000) );
  XOR U3200 ( .A(n3209), .B(n3202), .Z(n3208) );
  AND U3201 ( .A(n3027), .B(n3210), .Z(n3202) );
  AND U3202 ( .A(n3211), .B(n3212), .Z(n3209) );
  XOR U3203 ( .A(n3213), .B(n3207), .Z(n3211) );
  XNOR U3204 ( .A(n2997), .B(n3203), .Z(n3205) );
  XOR U3205 ( .A(n3214), .B(n3215), .Z(n2997) );
  AND U3206 ( .A(n39), .B(n3216), .Z(n3215) );
  XOR U3207 ( .A(n3217), .B(n3214), .Z(n3216) );
  XOR U3208 ( .A(n3218), .B(n3219), .Z(n3203) );
  AND U3209 ( .A(n3220), .B(n3221), .Z(n3219) );
  XNOR U3210 ( .A(n3218), .B(n3027), .Z(n3221) );
  XOR U3211 ( .A(n3222), .B(n3212), .Z(n3027) );
  XNOR U3212 ( .A(n3223), .B(n3207), .Z(n3212) );
  XOR U3213 ( .A(n3224), .B(n3225), .Z(n3207) );
  AND U3214 ( .A(n3226), .B(n3227), .Z(n3225) );
  XOR U3215 ( .A(n3228), .B(n3224), .Z(n3226) );
  XNOR U3216 ( .A(n3229), .B(n3230), .Z(n3223) );
  AND U3217 ( .A(n3231), .B(n3232), .Z(n3230) );
  XOR U3218 ( .A(n3229), .B(n3233), .Z(n3231) );
  XNOR U3219 ( .A(n3213), .B(n3210), .Z(n3222) );
  AND U3220 ( .A(n3234), .B(n3235), .Z(n3210) );
  XOR U3221 ( .A(n3236), .B(n3237), .Z(n3213) );
  AND U3222 ( .A(n3238), .B(n3239), .Z(n3237) );
  XOR U3223 ( .A(n3236), .B(n3240), .Z(n3238) );
  XNOR U3224 ( .A(n3024), .B(n3218), .Z(n3220) );
  XOR U3225 ( .A(n3241), .B(n3242), .Z(n3024) );
  AND U3226 ( .A(n39), .B(n3243), .Z(n3242) );
  XNOR U3227 ( .A(n3244), .B(n3241), .Z(n3243) );
  XOR U3228 ( .A(n3245), .B(n3246), .Z(n3218) );
  AND U3229 ( .A(n3247), .B(n3248), .Z(n3246) );
  XNOR U3230 ( .A(n3245), .B(n3234), .Z(n3248) );
  IV U3231 ( .A(n3075), .Z(n3234) );
  XNOR U3232 ( .A(n3249), .B(n3227), .Z(n3075) );
  XNOR U3233 ( .A(n3250), .B(n3233), .Z(n3227) );
  XOR U3234 ( .A(n3251), .B(n3252), .Z(n3233) );
  AND U3235 ( .A(n3253), .B(n3254), .Z(n3252) );
  XOR U3236 ( .A(n3251), .B(n3255), .Z(n3253) );
  XNOR U3237 ( .A(n3232), .B(n3224), .Z(n3250) );
  XOR U3238 ( .A(n3256), .B(n3257), .Z(n3224) );
  AND U3239 ( .A(n3258), .B(n3259), .Z(n3257) );
  XNOR U3240 ( .A(n3260), .B(n3256), .Z(n3258) );
  XNOR U3241 ( .A(n3261), .B(n3229), .Z(n3232) );
  XOR U3242 ( .A(n3262), .B(n3263), .Z(n3229) );
  AND U3243 ( .A(n3264), .B(n3265), .Z(n3263) );
  XOR U3244 ( .A(n3262), .B(n3266), .Z(n3264) );
  XNOR U3245 ( .A(n3267), .B(n3268), .Z(n3261) );
  AND U3246 ( .A(n3269), .B(n3270), .Z(n3268) );
  XNOR U3247 ( .A(n3267), .B(n3271), .Z(n3269) );
  XNOR U3248 ( .A(n3228), .B(n3235), .Z(n3249) );
  AND U3249 ( .A(n3171), .B(n3272), .Z(n3235) );
  XOR U3250 ( .A(n3240), .B(n3239), .Z(n3228) );
  XNOR U3251 ( .A(n3273), .B(n3236), .Z(n3239) );
  XOR U3252 ( .A(n3274), .B(n3275), .Z(n3236) );
  AND U3253 ( .A(n3276), .B(n3277), .Z(n3275) );
  XOR U3254 ( .A(n3274), .B(n3278), .Z(n3276) );
  XNOR U3255 ( .A(n3279), .B(n3280), .Z(n3273) );
  AND U3256 ( .A(n3281), .B(n3282), .Z(n3280) );
  XOR U3257 ( .A(n3279), .B(n3283), .Z(n3281) );
  XOR U3258 ( .A(n3284), .B(n3285), .Z(n3240) );
  AND U3259 ( .A(n3286), .B(n3287), .Z(n3285) );
  XOR U3260 ( .A(n3284), .B(n3288), .Z(n3286) );
  XNOR U3261 ( .A(n3072), .B(n3245), .Z(n3247) );
  XOR U3262 ( .A(n3289), .B(n3290), .Z(n3072) );
  AND U3263 ( .A(n39), .B(n3291), .Z(n3290) );
  XOR U3264 ( .A(n3292), .B(n3289), .Z(n3291) );
  XOR U3265 ( .A(n3293), .B(n3294), .Z(n3245) );
  AND U3266 ( .A(n3295), .B(n3296), .Z(n3294) );
  XNOR U3267 ( .A(n3293), .B(n3171), .Z(n3296) );
  XOR U3268 ( .A(n3297), .B(n3259), .Z(n3171) );
  XNOR U3269 ( .A(n3298), .B(n3266), .Z(n3259) );
  XOR U3270 ( .A(n3255), .B(n3254), .Z(n3266) );
  XNOR U3271 ( .A(n3299), .B(n3251), .Z(n3254) );
  XOR U3272 ( .A(n3300), .B(n3301), .Z(n3251) );
  AND U3273 ( .A(n3302), .B(n3303), .Z(n3301) );
  XNOR U3274 ( .A(n3304), .B(n3305), .Z(n3302) );
  IV U3275 ( .A(n3300), .Z(n3304) );
  XNOR U3276 ( .A(n3306), .B(n3307), .Z(n3299) );
  NOR U3277 ( .A(n3308), .B(n3309), .Z(n3307) );
  XNOR U3278 ( .A(n3306), .B(n3310), .Z(n3308) );
  XOR U3279 ( .A(n3311), .B(n3312), .Z(n3255) );
  NOR U3280 ( .A(n3313), .B(n3314), .Z(n3312) );
  XNOR U3281 ( .A(n3311), .B(n3315), .Z(n3313) );
  XNOR U3282 ( .A(n3265), .B(n3256), .Z(n3298) );
  XOR U3283 ( .A(n3316), .B(n3317), .Z(n3256) );
  AND U3284 ( .A(n3318), .B(n3319), .Z(n3317) );
  XOR U3285 ( .A(n3316), .B(n3320), .Z(n3318) );
  XOR U3286 ( .A(n3321), .B(n3271), .Z(n3265) );
  XOR U3287 ( .A(n3322), .B(n3323), .Z(n3271) );
  NOR U3288 ( .A(n3324), .B(n3325), .Z(n3323) );
  XOR U3289 ( .A(n3322), .B(n3326), .Z(n3324) );
  XNOR U3290 ( .A(n3270), .B(n3262), .Z(n3321) );
  XOR U3291 ( .A(n3327), .B(n3328), .Z(n3262) );
  AND U3292 ( .A(n3329), .B(n3330), .Z(n3328) );
  XOR U3293 ( .A(n3327), .B(n3331), .Z(n3329) );
  XNOR U3294 ( .A(n3332), .B(n3267), .Z(n3270) );
  XOR U3295 ( .A(n3333), .B(n3334), .Z(n3267) );
  AND U3296 ( .A(n3335), .B(n3336), .Z(n3334) );
  XNOR U3297 ( .A(n3337), .B(n3338), .Z(n3335) );
  IV U3298 ( .A(n3333), .Z(n3337) );
  XNOR U3299 ( .A(n3339), .B(n3340), .Z(n3332) );
  NOR U3300 ( .A(n3341), .B(n3342), .Z(n3340) );
  XNOR U3301 ( .A(n3339), .B(n3343), .Z(n3341) );
  XOR U3302 ( .A(n3260), .B(n3272), .Z(n3297) );
  NOR U3303 ( .A(n3194), .B(n3344), .Z(n3272) );
  XNOR U3304 ( .A(n3278), .B(n3277), .Z(n3260) );
  XNOR U3305 ( .A(n3345), .B(n3283), .Z(n3277) );
  XNOR U3306 ( .A(n3346), .B(n3347), .Z(n3283) );
  NOR U3307 ( .A(n3348), .B(n3349), .Z(n3347) );
  XOR U3308 ( .A(n3346), .B(n3350), .Z(n3348) );
  XNOR U3309 ( .A(n3282), .B(n3274), .Z(n3345) );
  XOR U3310 ( .A(n3351), .B(n3352), .Z(n3274) );
  AND U3311 ( .A(n3353), .B(n3354), .Z(n3352) );
  XOR U3312 ( .A(n3351), .B(n3355), .Z(n3353) );
  XNOR U3313 ( .A(n3356), .B(n3279), .Z(n3282) );
  XOR U3314 ( .A(n3357), .B(n3358), .Z(n3279) );
  AND U3315 ( .A(n3359), .B(n3360), .Z(n3358) );
  XNOR U3316 ( .A(n3361), .B(n3362), .Z(n3359) );
  IV U3317 ( .A(n3357), .Z(n3361) );
  XNOR U3318 ( .A(n3363), .B(n3364), .Z(n3356) );
  NOR U3319 ( .A(n3365), .B(n3366), .Z(n3364) );
  XNOR U3320 ( .A(n3363), .B(n3367), .Z(n3365) );
  XOR U3321 ( .A(n3288), .B(n3287), .Z(n3278) );
  XNOR U3322 ( .A(n3368), .B(n3284), .Z(n3287) );
  XOR U3323 ( .A(n3369), .B(n3370), .Z(n3284) );
  AND U3324 ( .A(n3371), .B(n3372), .Z(n3370) );
  XNOR U3325 ( .A(n3373), .B(n3374), .Z(n3371) );
  IV U3326 ( .A(n3369), .Z(n3373) );
  XNOR U3327 ( .A(n3375), .B(n3376), .Z(n3368) );
  NOR U3328 ( .A(n3377), .B(n3378), .Z(n3376) );
  XNOR U3329 ( .A(n3375), .B(n3379), .Z(n3377) );
  XOR U3330 ( .A(n3380), .B(n3381), .Z(n3288) );
  NOR U3331 ( .A(n3382), .B(n3383), .Z(n3381) );
  XNOR U3332 ( .A(n3380), .B(n3384), .Z(n3382) );
  XNOR U3333 ( .A(n3168), .B(n3293), .Z(n3295) );
  XOR U3334 ( .A(n3385), .B(n3386), .Z(n3168) );
  AND U3335 ( .A(n39), .B(n3387), .Z(n3386) );
  XNOR U3336 ( .A(n3388), .B(n3385), .Z(n3387) );
  AND U3337 ( .A(n3191), .B(n3194), .Z(n3293) );
  XOR U3338 ( .A(n3389), .B(n3344), .Z(n3194) );
  XNOR U3339 ( .A(p_input[256]), .B(p_input[512]), .Z(n3344) );
  XNOR U3340 ( .A(n3320), .B(n3319), .Z(n3389) );
  XNOR U3341 ( .A(n3390), .B(n3331), .Z(n3319) );
  XOR U3342 ( .A(n3305), .B(n3303), .Z(n3331) );
  XNOR U3343 ( .A(n3391), .B(n3310), .Z(n3303) );
  XOR U3344 ( .A(p_input[280]), .B(p_input[536]), .Z(n3310) );
  XOR U3345 ( .A(n3300), .B(n3309), .Z(n3391) );
  XOR U3346 ( .A(n3392), .B(n3306), .Z(n3309) );
  XOR U3347 ( .A(p_input[278]), .B(p_input[534]), .Z(n3306) );
  XOR U3348 ( .A(p_input[279]), .B(n1634), .Z(n3392) );
  XOR U3349 ( .A(p_input[274]), .B(p_input[530]), .Z(n3300) );
  XNOR U3350 ( .A(n3315), .B(n3314), .Z(n3305) );
  XOR U3351 ( .A(n3393), .B(n3311), .Z(n3314) );
  XOR U3352 ( .A(p_input[275]), .B(p_input[531]), .Z(n3311) );
  XOR U3353 ( .A(p_input[276]), .B(n1636), .Z(n3393) );
  XOR U3354 ( .A(p_input[277]), .B(p_input[533]), .Z(n3315) );
  XOR U3355 ( .A(n3330), .B(n3394), .Z(n3390) );
  IV U3356 ( .A(n3316), .Z(n3394) );
  XOR U3357 ( .A(p_input[257]), .B(p_input[513]), .Z(n3316) );
  XNOR U3358 ( .A(n3395), .B(n3338), .Z(n3330) );
  XNOR U3359 ( .A(n3326), .B(n3325), .Z(n3338) );
  XNOR U3360 ( .A(n3396), .B(n3322), .Z(n3325) );
  XNOR U3361 ( .A(p_input[282]), .B(p_input[538]), .Z(n3322) );
  XOR U3362 ( .A(p_input[283]), .B(n1640), .Z(n3396) );
  XOR U3363 ( .A(p_input[284]), .B(p_input[540]), .Z(n3326) );
  XOR U3364 ( .A(n3336), .B(n3397), .Z(n3395) );
  IV U3365 ( .A(n3327), .Z(n3397) );
  XOR U3366 ( .A(p_input[273]), .B(p_input[529]), .Z(n3327) );
  XNOR U3367 ( .A(n3398), .B(n3343), .Z(n3336) );
  XNOR U3368 ( .A(p_input[287]), .B(n1643), .Z(n3343) );
  XOR U3369 ( .A(n3333), .B(n3342), .Z(n3398) );
  XOR U3370 ( .A(n3399), .B(n3339), .Z(n3342) );
  XOR U3371 ( .A(p_input[285]), .B(p_input[541]), .Z(n3339) );
  XOR U3372 ( .A(p_input[286]), .B(n1645), .Z(n3399) );
  XOR U3373 ( .A(p_input[281]), .B(p_input[537]), .Z(n3333) );
  XOR U3374 ( .A(n3355), .B(n3354), .Z(n3320) );
  XNOR U3375 ( .A(n3400), .B(n3362), .Z(n3354) );
  XNOR U3376 ( .A(n3350), .B(n3349), .Z(n3362) );
  XNOR U3377 ( .A(n3401), .B(n3346), .Z(n3349) );
  XNOR U3378 ( .A(p_input[267]), .B(p_input[523]), .Z(n3346) );
  XOR U3379 ( .A(p_input[268]), .B(n1648), .Z(n3401) );
  XOR U3380 ( .A(p_input[269]), .B(p_input[525]), .Z(n3350) );
  XOR U3381 ( .A(n3360), .B(n3402), .Z(n3400) );
  IV U3382 ( .A(n3351), .Z(n3402) );
  XOR U3383 ( .A(p_input[258]), .B(p_input[514]), .Z(n3351) );
  XNOR U3384 ( .A(n3403), .B(n3367), .Z(n3360) );
  XNOR U3385 ( .A(p_input[272]), .B(n1651), .Z(n3367) );
  XOR U3386 ( .A(n3357), .B(n3366), .Z(n3403) );
  XOR U3387 ( .A(n3404), .B(n3363), .Z(n3366) );
  XOR U3388 ( .A(p_input[270]), .B(p_input[526]), .Z(n3363) );
  XOR U3389 ( .A(p_input[271]), .B(n1653), .Z(n3404) );
  XOR U3390 ( .A(p_input[266]), .B(p_input[522]), .Z(n3357) );
  XOR U3391 ( .A(n3374), .B(n3372), .Z(n3355) );
  XNOR U3392 ( .A(n3405), .B(n3379), .Z(n3372) );
  XOR U3393 ( .A(p_input[265]), .B(p_input[521]), .Z(n3379) );
  XOR U3394 ( .A(n3369), .B(n3378), .Z(n3405) );
  XOR U3395 ( .A(n3406), .B(n3375), .Z(n3378) );
  XOR U3396 ( .A(p_input[263]), .B(p_input[519]), .Z(n3375) );
  XOR U3397 ( .A(p_input[264]), .B(n1877), .Z(n3406) );
  XOR U3398 ( .A(p_input[259]), .B(p_input[515]), .Z(n3369) );
  XNOR U3399 ( .A(n3384), .B(n3383), .Z(n3374) );
  XOR U3400 ( .A(n3407), .B(n3380), .Z(n3383) );
  XOR U3401 ( .A(p_input[260]), .B(p_input[516]), .Z(n3380) );
  XOR U3402 ( .A(p_input[261]), .B(n1879), .Z(n3407) );
  XOR U3403 ( .A(p_input[262]), .B(p_input[518]), .Z(n3384) );
  XOR U3404 ( .A(n3408), .B(n3409), .Z(n3191) );
  AND U3405 ( .A(n39), .B(n3410), .Z(n3409) );
  XNOR U3406 ( .A(n3411), .B(n3408), .Z(n3410) );
  XNOR U3407 ( .A(n3412), .B(n3413), .Z(n39) );
  NOR U3408 ( .A(n3414), .B(n3415), .Z(n3413) );
  XOR U3409 ( .A(n3200), .B(n3412), .Z(n3415) );
  AND U3410 ( .A(n3416), .B(n3417), .Z(n3200) );
  NOR U3411 ( .A(n3412), .B(n3199), .Z(n3414) );
  AND U3412 ( .A(n3418), .B(n3419), .Z(n3199) );
  XOR U3413 ( .A(n3420), .B(n3421), .Z(n3412) );
  AND U3414 ( .A(n3422), .B(n3423), .Z(n3421) );
  XNOR U3415 ( .A(n3420), .B(n3418), .Z(n3423) );
  IV U3416 ( .A(n3217), .Z(n3418) );
  XOR U3417 ( .A(n3424), .B(n3425), .Z(n3217) );
  XOR U3418 ( .A(n3426), .B(n3419), .Z(n3425) );
  AND U3419 ( .A(n3244), .B(n3427), .Z(n3419) );
  AND U3420 ( .A(n3428), .B(n3429), .Z(n3426) );
  XOR U3421 ( .A(n3430), .B(n3424), .Z(n3428) );
  XNOR U3422 ( .A(n3214), .B(n3420), .Z(n3422) );
  XOR U3423 ( .A(n3431), .B(n3432), .Z(n3214) );
  AND U3424 ( .A(n43), .B(n3433), .Z(n3432) );
  XOR U3425 ( .A(n3434), .B(n3431), .Z(n3433) );
  XOR U3426 ( .A(n3435), .B(n3436), .Z(n3420) );
  AND U3427 ( .A(n3437), .B(n3438), .Z(n3436) );
  XNOR U3428 ( .A(n3435), .B(n3244), .Z(n3438) );
  XOR U3429 ( .A(n3439), .B(n3429), .Z(n3244) );
  XNOR U3430 ( .A(n3440), .B(n3424), .Z(n3429) );
  XOR U3431 ( .A(n3441), .B(n3442), .Z(n3424) );
  AND U3432 ( .A(n3443), .B(n3444), .Z(n3442) );
  XOR U3433 ( .A(n3445), .B(n3441), .Z(n3443) );
  XNOR U3434 ( .A(n3446), .B(n3447), .Z(n3440) );
  AND U3435 ( .A(n3448), .B(n3449), .Z(n3447) );
  XOR U3436 ( .A(n3446), .B(n3450), .Z(n3448) );
  XNOR U3437 ( .A(n3430), .B(n3427), .Z(n3439) );
  AND U3438 ( .A(n3451), .B(n3452), .Z(n3427) );
  XOR U3439 ( .A(n3453), .B(n3454), .Z(n3430) );
  AND U3440 ( .A(n3455), .B(n3456), .Z(n3454) );
  XOR U3441 ( .A(n3453), .B(n3457), .Z(n3455) );
  XNOR U3442 ( .A(n3241), .B(n3435), .Z(n3437) );
  XOR U3443 ( .A(n3458), .B(n3459), .Z(n3241) );
  AND U3444 ( .A(n43), .B(n3460), .Z(n3459) );
  XNOR U3445 ( .A(n3461), .B(n3458), .Z(n3460) );
  XOR U3446 ( .A(n3462), .B(n3463), .Z(n3435) );
  AND U3447 ( .A(n3464), .B(n3465), .Z(n3463) );
  XNOR U3448 ( .A(n3462), .B(n3451), .Z(n3465) );
  IV U3449 ( .A(n3292), .Z(n3451) );
  XNOR U3450 ( .A(n3466), .B(n3444), .Z(n3292) );
  XNOR U3451 ( .A(n3467), .B(n3450), .Z(n3444) );
  XOR U3452 ( .A(n3468), .B(n3469), .Z(n3450) );
  AND U3453 ( .A(n3470), .B(n3471), .Z(n3469) );
  XOR U3454 ( .A(n3468), .B(n3472), .Z(n3470) );
  XNOR U3455 ( .A(n3449), .B(n3441), .Z(n3467) );
  XOR U3456 ( .A(n3473), .B(n3474), .Z(n3441) );
  AND U3457 ( .A(n3475), .B(n3476), .Z(n3474) );
  XNOR U3458 ( .A(n3477), .B(n3473), .Z(n3475) );
  XNOR U3459 ( .A(n3478), .B(n3446), .Z(n3449) );
  XOR U3460 ( .A(n3479), .B(n3480), .Z(n3446) );
  AND U3461 ( .A(n3481), .B(n3482), .Z(n3480) );
  XOR U3462 ( .A(n3479), .B(n3483), .Z(n3481) );
  XNOR U3463 ( .A(n3484), .B(n3485), .Z(n3478) );
  AND U3464 ( .A(n3486), .B(n3487), .Z(n3485) );
  XNOR U3465 ( .A(n3484), .B(n3488), .Z(n3486) );
  XNOR U3466 ( .A(n3445), .B(n3452), .Z(n3466) );
  AND U3467 ( .A(n3388), .B(n3489), .Z(n3452) );
  XOR U3468 ( .A(n3457), .B(n3456), .Z(n3445) );
  XNOR U3469 ( .A(n3490), .B(n3453), .Z(n3456) );
  XOR U3470 ( .A(n3491), .B(n3492), .Z(n3453) );
  AND U3471 ( .A(n3493), .B(n3494), .Z(n3492) );
  XOR U3472 ( .A(n3491), .B(n3495), .Z(n3493) );
  XNOR U3473 ( .A(n3496), .B(n3497), .Z(n3490) );
  AND U3474 ( .A(n3498), .B(n3499), .Z(n3497) );
  XOR U3475 ( .A(n3496), .B(n3500), .Z(n3498) );
  XOR U3476 ( .A(n3501), .B(n3502), .Z(n3457) );
  AND U3477 ( .A(n3503), .B(n3504), .Z(n3502) );
  XOR U3478 ( .A(n3501), .B(n3505), .Z(n3503) );
  XNOR U3479 ( .A(n3289), .B(n3462), .Z(n3464) );
  XOR U3480 ( .A(n3506), .B(n3507), .Z(n3289) );
  AND U3481 ( .A(n43), .B(n3508), .Z(n3507) );
  XOR U3482 ( .A(n3509), .B(n3506), .Z(n3508) );
  XOR U3483 ( .A(n3510), .B(n3511), .Z(n3462) );
  AND U3484 ( .A(n3512), .B(n3513), .Z(n3511) );
  XNOR U3485 ( .A(n3510), .B(n3388), .Z(n3513) );
  XOR U3486 ( .A(n3514), .B(n3476), .Z(n3388) );
  XNOR U3487 ( .A(n3515), .B(n3483), .Z(n3476) );
  XOR U3488 ( .A(n3472), .B(n3471), .Z(n3483) );
  XNOR U3489 ( .A(n3516), .B(n3468), .Z(n3471) );
  XOR U3490 ( .A(n3517), .B(n3518), .Z(n3468) );
  AND U3491 ( .A(n3519), .B(n3520), .Z(n3518) );
  XNOR U3492 ( .A(n3521), .B(n3522), .Z(n3519) );
  IV U3493 ( .A(n3517), .Z(n3521) );
  XNOR U3494 ( .A(n3523), .B(n3524), .Z(n3516) );
  NOR U3495 ( .A(n3525), .B(n3526), .Z(n3524) );
  XNOR U3496 ( .A(n3523), .B(n3527), .Z(n3525) );
  XOR U3497 ( .A(n3528), .B(n3529), .Z(n3472) );
  NOR U3498 ( .A(n3530), .B(n3531), .Z(n3529) );
  XNOR U3499 ( .A(n3528), .B(n3532), .Z(n3530) );
  XNOR U3500 ( .A(n3482), .B(n3473), .Z(n3515) );
  XOR U3501 ( .A(n3533), .B(n3534), .Z(n3473) );
  AND U3502 ( .A(n3535), .B(n3536), .Z(n3534) );
  XOR U3503 ( .A(n3533), .B(n3537), .Z(n3535) );
  XOR U3504 ( .A(n3538), .B(n3488), .Z(n3482) );
  XOR U3505 ( .A(n3539), .B(n3540), .Z(n3488) );
  NOR U3506 ( .A(n3541), .B(n3542), .Z(n3540) );
  XOR U3507 ( .A(n3539), .B(n3543), .Z(n3541) );
  XNOR U3508 ( .A(n3487), .B(n3479), .Z(n3538) );
  XOR U3509 ( .A(n3544), .B(n3545), .Z(n3479) );
  AND U3510 ( .A(n3546), .B(n3547), .Z(n3545) );
  XOR U3511 ( .A(n3544), .B(n3548), .Z(n3546) );
  XNOR U3512 ( .A(n3549), .B(n3484), .Z(n3487) );
  XOR U3513 ( .A(n3550), .B(n3551), .Z(n3484) );
  AND U3514 ( .A(n3552), .B(n3553), .Z(n3551) );
  XNOR U3515 ( .A(n3554), .B(n3555), .Z(n3552) );
  IV U3516 ( .A(n3550), .Z(n3554) );
  XNOR U3517 ( .A(n3556), .B(n3557), .Z(n3549) );
  NOR U3518 ( .A(n3558), .B(n3559), .Z(n3557) );
  XNOR U3519 ( .A(n3556), .B(n3560), .Z(n3558) );
  XOR U3520 ( .A(n3477), .B(n3489), .Z(n3514) );
  NOR U3521 ( .A(n3411), .B(n3561), .Z(n3489) );
  XNOR U3522 ( .A(n3495), .B(n3494), .Z(n3477) );
  XNOR U3523 ( .A(n3562), .B(n3500), .Z(n3494) );
  XNOR U3524 ( .A(n3563), .B(n3564), .Z(n3500) );
  NOR U3525 ( .A(n3565), .B(n3566), .Z(n3564) );
  XOR U3526 ( .A(n3563), .B(n3567), .Z(n3565) );
  XNOR U3527 ( .A(n3499), .B(n3491), .Z(n3562) );
  XOR U3528 ( .A(n3568), .B(n3569), .Z(n3491) );
  AND U3529 ( .A(n3570), .B(n3571), .Z(n3569) );
  XOR U3530 ( .A(n3568), .B(n3572), .Z(n3570) );
  XNOR U3531 ( .A(n3573), .B(n3496), .Z(n3499) );
  XOR U3532 ( .A(n3574), .B(n3575), .Z(n3496) );
  AND U3533 ( .A(n3576), .B(n3577), .Z(n3575) );
  XNOR U3534 ( .A(n3578), .B(n3579), .Z(n3576) );
  IV U3535 ( .A(n3574), .Z(n3578) );
  XNOR U3536 ( .A(n3580), .B(n3581), .Z(n3573) );
  NOR U3537 ( .A(n3582), .B(n3583), .Z(n3581) );
  XNOR U3538 ( .A(n3580), .B(n3584), .Z(n3582) );
  XOR U3539 ( .A(n3505), .B(n3504), .Z(n3495) );
  XNOR U3540 ( .A(n3585), .B(n3501), .Z(n3504) );
  XOR U3541 ( .A(n3586), .B(n3587), .Z(n3501) );
  AND U3542 ( .A(n3588), .B(n3589), .Z(n3587) );
  XNOR U3543 ( .A(n3590), .B(n3591), .Z(n3588) );
  IV U3544 ( .A(n3586), .Z(n3590) );
  XNOR U3545 ( .A(n3592), .B(n3593), .Z(n3585) );
  NOR U3546 ( .A(n3594), .B(n3595), .Z(n3593) );
  XNOR U3547 ( .A(n3592), .B(n3596), .Z(n3594) );
  XOR U3548 ( .A(n3597), .B(n3598), .Z(n3505) );
  NOR U3549 ( .A(n3599), .B(n3600), .Z(n3598) );
  XNOR U3550 ( .A(n3597), .B(n3601), .Z(n3599) );
  XNOR U3551 ( .A(n3385), .B(n3510), .Z(n3512) );
  XOR U3552 ( .A(n3602), .B(n3603), .Z(n3385) );
  AND U3553 ( .A(n43), .B(n3604), .Z(n3603) );
  XNOR U3554 ( .A(n3605), .B(n3602), .Z(n3604) );
  AND U3555 ( .A(n3408), .B(n3411), .Z(n3510) );
  XOR U3556 ( .A(n3606), .B(n3561), .Z(n3411) );
  XNOR U3557 ( .A(p_input[288]), .B(p_input[512]), .Z(n3561) );
  XNOR U3558 ( .A(n3537), .B(n3536), .Z(n3606) );
  XNOR U3559 ( .A(n3607), .B(n3548), .Z(n3536) );
  XOR U3560 ( .A(n3522), .B(n3520), .Z(n3548) );
  XNOR U3561 ( .A(n3608), .B(n3527), .Z(n3520) );
  XOR U3562 ( .A(p_input[312]), .B(p_input[536]), .Z(n3527) );
  XOR U3563 ( .A(n3517), .B(n3526), .Z(n3608) );
  XOR U3564 ( .A(n3609), .B(n3523), .Z(n3526) );
  XOR U3565 ( .A(p_input[310]), .B(p_input[534]), .Z(n3523) );
  XOR U3566 ( .A(p_input[311]), .B(n1634), .Z(n3609) );
  XOR U3567 ( .A(p_input[306]), .B(p_input[530]), .Z(n3517) );
  XNOR U3568 ( .A(n3532), .B(n3531), .Z(n3522) );
  XOR U3569 ( .A(n3610), .B(n3528), .Z(n3531) );
  XOR U3570 ( .A(p_input[307]), .B(p_input[531]), .Z(n3528) );
  XOR U3571 ( .A(p_input[308]), .B(n1636), .Z(n3610) );
  XOR U3572 ( .A(p_input[309]), .B(p_input[533]), .Z(n3532) );
  XOR U3573 ( .A(n3547), .B(n3611), .Z(n3607) );
  IV U3574 ( .A(n3533), .Z(n3611) );
  XOR U3575 ( .A(p_input[289]), .B(p_input[513]), .Z(n3533) );
  XNOR U3576 ( .A(n3612), .B(n3555), .Z(n3547) );
  XNOR U3577 ( .A(n3543), .B(n3542), .Z(n3555) );
  XNOR U3578 ( .A(n3613), .B(n3539), .Z(n3542) );
  XNOR U3579 ( .A(p_input[314]), .B(p_input[538]), .Z(n3539) );
  XOR U3580 ( .A(p_input[315]), .B(n1640), .Z(n3613) );
  XOR U3581 ( .A(p_input[316]), .B(p_input[540]), .Z(n3543) );
  XOR U3582 ( .A(n3553), .B(n3614), .Z(n3612) );
  IV U3583 ( .A(n3544), .Z(n3614) );
  XOR U3584 ( .A(p_input[305]), .B(p_input[529]), .Z(n3544) );
  XNOR U3585 ( .A(n3615), .B(n3560), .Z(n3553) );
  XNOR U3586 ( .A(p_input[319]), .B(n1643), .Z(n3560) );
  XOR U3587 ( .A(n3550), .B(n3559), .Z(n3615) );
  XOR U3588 ( .A(n3616), .B(n3556), .Z(n3559) );
  XOR U3589 ( .A(p_input[317]), .B(p_input[541]), .Z(n3556) );
  XOR U3590 ( .A(p_input[318]), .B(n1645), .Z(n3616) );
  XOR U3591 ( .A(p_input[313]), .B(p_input[537]), .Z(n3550) );
  XOR U3592 ( .A(n3572), .B(n3571), .Z(n3537) );
  XNOR U3593 ( .A(n3617), .B(n3579), .Z(n3571) );
  XNOR U3594 ( .A(n3567), .B(n3566), .Z(n3579) );
  XNOR U3595 ( .A(n3618), .B(n3563), .Z(n3566) );
  XNOR U3596 ( .A(p_input[299]), .B(p_input[523]), .Z(n3563) );
  XOR U3597 ( .A(p_input[300]), .B(n1648), .Z(n3618) );
  XOR U3598 ( .A(p_input[301]), .B(p_input[525]), .Z(n3567) );
  XOR U3599 ( .A(n3577), .B(n3619), .Z(n3617) );
  IV U3600 ( .A(n3568), .Z(n3619) );
  XOR U3601 ( .A(p_input[290]), .B(p_input[514]), .Z(n3568) );
  XNOR U3602 ( .A(n3620), .B(n3584), .Z(n3577) );
  XNOR U3603 ( .A(p_input[304]), .B(n1651), .Z(n3584) );
  XOR U3604 ( .A(n3574), .B(n3583), .Z(n3620) );
  XOR U3605 ( .A(n3621), .B(n3580), .Z(n3583) );
  XOR U3606 ( .A(p_input[302]), .B(p_input[526]), .Z(n3580) );
  XOR U3607 ( .A(p_input[303]), .B(n1653), .Z(n3621) );
  XOR U3608 ( .A(p_input[298]), .B(p_input[522]), .Z(n3574) );
  XOR U3609 ( .A(n3591), .B(n3589), .Z(n3572) );
  XNOR U3610 ( .A(n3622), .B(n3596), .Z(n3589) );
  XOR U3611 ( .A(p_input[297]), .B(p_input[521]), .Z(n3596) );
  XOR U3612 ( .A(n3586), .B(n3595), .Z(n3622) );
  XOR U3613 ( .A(n3623), .B(n3592), .Z(n3595) );
  XOR U3614 ( .A(p_input[295]), .B(p_input[519]), .Z(n3592) );
  XOR U3615 ( .A(p_input[296]), .B(n1877), .Z(n3623) );
  XOR U3616 ( .A(p_input[291]), .B(p_input[515]), .Z(n3586) );
  XNOR U3617 ( .A(n3601), .B(n3600), .Z(n3591) );
  XOR U3618 ( .A(n3624), .B(n3597), .Z(n3600) );
  XOR U3619 ( .A(p_input[292]), .B(p_input[516]), .Z(n3597) );
  XOR U3620 ( .A(p_input[293]), .B(n1879), .Z(n3624) );
  XOR U3621 ( .A(p_input[294]), .B(p_input[518]), .Z(n3601) );
  XOR U3622 ( .A(n3625), .B(n3626), .Z(n3408) );
  AND U3623 ( .A(n43), .B(n3627), .Z(n3626) );
  XNOR U3624 ( .A(n3628), .B(n3625), .Z(n3627) );
  XNOR U3625 ( .A(n3629), .B(n3630), .Z(n43) );
  NOR U3626 ( .A(n3631), .B(n3632), .Z(n3630) );
  XOR U3627 ( .A(n3417), .B(n3629), .Z(n3632) );
  AND U3628 ( .A(n3633), .B(n3634), .Z(n3417) );
  NOR U3629 ( .A(n3629), .B(n3416), .Z(n3631) );
  AND U3630 ( .A(n3635), .B(n3636), .Z(n3416) );
  XOR U3631 ( .A(n3637), .B(n3638), .Z(n3629) );
  AND U3632 ( .A(n3639), .B(n3640), .Z(n3638) );
  XNOR U3633 ( .A(n3637), .B(n3635), .Z(n3640) );
  IV U3634 ( .A(n3434), .Z(n3635) );
  XOR U3635 ( .A(n3641), .B(n3642), .Z(n3434) );
  XOR U3636 ( .A(n3643), .B(n3636), .Z(n3642) );
  AND U3637 ( .A(n3461), .B(n3644), .Z(n3636) );
  AND U3638 ( .A(n3645), .B(n3646), .Z(n3643) );
  XOR U3639 ( .A(n3647), .B(n3641), .Z(n3645) );
  XNOR U3640 ( .A(n3431), .B(n3637), .Z(n3639) );
  XOR U3641 ( .A(n3648), .B(n3649), .Z(n3431) );
  AND U3642 ( .A(n47), .B(n3650), .Z(n3649) );
  XOR U3643 ( .A(n3651), .B(n3648), .Z(n3650) );
  XOR U3644 ( .A(n3652), .B(n3653), .Z(n3637) );
  AND U3645 ( .A(n3654), .B(n3655), .Z(n3653) );
  XNOR U3646 ( .A(n3652), .B(n3461), .Z(n3655) );
  XOR U3647 ( .A(n3656), .B(n3646), .Z(n3461) );
  XNOR U3648 ( .A(n3657), .B(n3641), .Z(n3646) );
  XOR U3649 ( .A(n3658), .B(n3659), .Z(n3641) );
  AND U3650 ( .A(n3660), .B(n3661), .Z(n3659) );
  XOR U3651 ( .A(n3662), .B(n3658), .Z(n3660) );
  XNOR U3652 ( .A(n3663), .B(n3664), .Z(n3657) );
  AND U3653 ( .A(n3665), .B(n3666), .Z(n3664) );
  XOR U3654 ( .A(n3663), .B(n3667), .Z(n3665) );
  XNOR U3655 ( .A(n3647), .B(n3644), .Z(n3656) );
  AND U3656 ( .A(n3668), .B(n3669), .Z(n3644) );
  XOR U3657 ( .A(n3670), .B(n3671), .Z(n3647) );
  AND U3658 ( .A(n3672), .B(n3673), .Z(n3671) );
  XOR U3659 ( .A(n3670), .B(n3674), .Z(n3672) );
  XNOR U3660 ( .A(n3458), .B(n3652), .Z(n3654) );
  XOR U3661 ( .A(n3675), .B(n3676), .Z(n3458) );
  AND U3662 ( .A(n47), .B(n3677), .Z(n3676) );
  XNOR U3663 ( .A(n3678), .B(n3675), .Z(n3677) );
  XOR U3664 ( .A(n3679), .B(n3680), .Z(n3652) );
  AND U3665 ( .A(n3681), .B(n3682), .Z(n3680) );
  XNOR U3666 ( .A(n3679), .B(n3668), .Z(n3682) );
  IV U3667 ( .A(n3509), .Z(n3668) );
  XNOR U3668 ( .A(n3683), .B(n3661), .Z(n3509) );
  XNOR U3669 ( .A(n3684), .B(n3667), .Z(n3661) );
  XOR U3670 ( .A(n3685), .B(n3686), .Z(n3667) );
  AND U3671 ( .A(n3687), .B(n3688), .Z(n3686) );
  XOR U3672 ( .A(n3685), .B(n3689), .Z(n3687) );
  XNOR U3673 ( .A(n3666), .B(n3658), .Z(n3684) );
  XOR U3674 ( .A(n3690), .B(n3691), .Z(n3658) );
  AND U3675 ( .A(n3692), .B(n3693), .Z(n3691) );
  XNOR U3676 ( .A(n3694), .B(n3690), .Z(n3692) );
  XNOR U3677 ( .A(n3695), .B(n3663), .Z(n3666) );
  XOR U3678 ( .A(n3696), .B(n3697), .Z(n3663) );
  AND U3679 ( .A(n3698), .B(n3699), .Z(n3697) );
  XOR U3680 ( .A(n3696), .B(n3700), .Z(n3698) );
  XNOR U3681 ( .A(n3701), .B(n3702), .Z(n3695) );
  AND U3682 ( .A(n3703), .B(n3704), .Z(n3702) );
  XNOR U3683 ( .A(n3701), .B(n3705), .Z(n3703) );
  XNOR U3684 ( .A(n3662), .B(n3669), .Z(n3683) );
  AND U3685 ( .A(n3605), .B(n3706), .Z(n3669) );
  XOR U3686 ( .A(n3674), .B(n3673), .Z(n3662) );
  XNOR U3687 ( .A(n3707), .B(n3670), .Z(n3673) );
  XOR U3688 ( .A(n3708), .B(n3709), .Z(n3670) );
  AND U3689 ( .A(n3710), .B(n3711), .Z(n3709) );
  XOR U3690 ( .A(n3708), .B(n3712), .Z(n3710) );
  XNOR U3691 ( .A(n3713), .B(n3714), .Z(n3707) );
  AND U3692 ( .A(n3715), .B(n3716), .Z(n3714) );
  XOR U3693 ( .A(n3713), .B(n3717), .Z(n3715) );
  XOR U3694 ( .A(n3718), .B(n3719), .Z(n3674) );
  AND U3695 ( .A(n3720), .B(n3721), .Z(n3719) );
  XOR U3696 ( .A(n3718), .B(n3722), .Z(n3720) );
  XNOR U3697 ( .A(n3506), .B(n3679), .Z(n3681) );
  XOR U3698 ( .A(n3723), .B(n3724), .Z(n3506) );
  AND U3699 ( .A(n47), .B(n3725), .Z(n3724) );
  XOR U3700 ( .A(n3726), .B(n3723), .Z(n3725) );
  XOR U3701 ( .A(n3727), .B(n3728), .Z(n3679) );
  AND U3702 ( .A(n3729), .B(n3730), .Z(n3728) );
  XNOR U3703 ( .A(n3727), .B(n3605), .Z(n3730) );
  XOR U3704 ( .A(n3731), .B(n3693), .Z(n3605) );
  XNOR U3705 ( .A(n3732), .B(n3700), .Z(n3693) );
  XOR U3706 ( .A(n3689), .B(n3688), .Z(n3700) );
  XNOR U3707 ( .A(n3733), .B(n3685), .Z(n3688) );
  XOR U3708 ( .A(n3734), .B(n3735), .Z(n3685) );
  AND U3709 ( .A(n3736), .B(n3737), .Z(n3735) );
  XNOR U3710 ( .A(n3738), .B(n3739), .Z(n3736) );
  IV U3711 ( .A(n3734), .Z(n3738) );
  XNOR U3712 ( .A(n3740), .B(n3741), .Z(n3733) );
  NOR U3713 ( .A(n3742), .B(n3743), .Z(n3741) );
  XNOR U3714 ( .A(n3740), .B(n3744), .Z(n3742) );
  XOR U3715 ( .A(n3745), .B(n3746), .Z(n3689) );
  NOR U3716 ( .A(n3747), .B(n3748), .Z(n3746) );
  XNOR U3717 ( .A(n3745), .B(n3749), .Z(n3747) );
  XNOR U3718 ( .A(n3699), .B(n3690), .Z(n3732) );
  XOR U3719 ( .A(n3750), .B(n3751), .Z(n3690) );
  AND U3720 ( .A(n3752), .B(n3753), .Z(n3751) );
  XOR U3721 ( .A(n3750), .B(n3754), .Z(n3752) );
  XOR U3722 ( .A(n3755), .B(n3705), .Z(n3699) );
  XOR U3723 ( .A(n3756), .B(n3757), .Z(n3705) );
  NOR U3724 ( .A(n3758), .B(n3759), .Z(n3757) );
  XOR U3725 ( .A(n3756), .B(n3760), .Z(n3758) );
  XNOR U3726 ( .A(n3704), .B(n3696), .Z(n3755) );
  XOR U3727 ( .A(n3761), .B(n3762), .Z(n3696) );
  AND U3728 ( .A(n3763), .B(n3764), .Z(n3762) );
  XOR U3729 ( .A(n3761), .B(n3765), .Z(n3763) );
  XNOR U3730 ( .A(n3766), .B(n3701), .Z(n3704) );
  XOR U3731 ( .A(n3767), .B(n3768), .Z(n3701) );
  AND U3732 ( .A(n3769), .B(n3770), .Z(n3768) );
  XNOR U3733 ( .A(n3771), .B(n3772), .Z(n3769) );
  IV U3734 ( .A(n3767), .Z(n3771) );
  XNOR U3735 ( .A(n3773), .B(n3774), .Z(n3766) );
  NOR U3736 ( .A(n3775), .B(n3776), .Z(n3774) );
  XNOR U3737 ( .A(n3773), .B(n3777), .Z(n3775) );
  XOR U3738 ( .A(n3694), .B(n3706), .Z(n3731) );
  NOR U3739 ( .A(n3628), .B(n3778), .Z(n3706) );
  XNOR U3740 ( .A(n3712), .B(n3711), .Z(n3694) );
  XNOR U3741 ( .A(n3779), .B(n3717), .Z(n3711) );
  XNOR U3742 ( .A(n3780), .B(n3781), .Z(n3717) );
  NOR U3743 ( .A(n3782), .B(n3783), .Z(n3781) );
  XOR U3744 ( .A(n3780), .B(n3784), .Z(n3782) );
  XNOR U3745 ( .A(n3716), .B(n3708), .Z(n3779) );
  XOR U3746 ( .A(n3785), .B(n3786), .Z(n3708) );
  AND U3747 ( .A(n3787), .B(n3788), .Z(n3786) );
  XOR U3748 ( .A(n3785), .B(n3789), .Z(n3787) );
  XNOR U3749 ( .A(n3790), .B(n3713), .Z(n3716) );
  XOR U3750 ( .A(n3791), .B(n3792), .Z(n3713) );
  AND U3751 ( .A(n3793), .B(n3794), .Z(n3792) );
  XNOR U3752 ( .A(n3795), .B(n3796), .Z(n3793) );
  IV U3753 ( .A(n3791), .Z(n3795) );
  XNOR U3754 ( .A(n3797), .B(n3798), .Z(n3790) );
  NOR U3755 ( .A(n3799), .B(n3800), .Z(n3798) );
  XNOR U3756 ( .A(n3797), .B(n3801), .Z(n3799) );
  XOR U3757 ( .A(n3722), .B(n3721), .Z(n3712) );
  XNOR U3758 ( .A(n3802), .B(n3718), .Z(n3721) );
  XOR U3759 ( .A(n3803), .B(n3804), .Z(n3718) );
  AND U3760 ( .A(n3805), .B(n3806), .Z(n3804) );
  XNOR U3761 ( .A(n3807), .B(n3808), .Z(n3805) );
  IV U3762 ( .A(n3803), .Z(n3807) );
  XNOR U3763 ( .A(n3809), .B(n3810), .Z(n3802) );
  NOR U3764 ( .A(n3811), .B(n3812), .Z(n3810) );
  XNOR U3765 ( .A(n3809), .B(n3813), .Z(n3811) );
  XOR U3766 ( .A(n3814), .B(n3815), .Z(n3722) );
  NOR U3767 ( .A(n3816), .B(n3817), .Z(n3815) );
  XNOR U3768 ( .A(n3814), .B(n3818), .Z(n3816) );
  XNOR U3769 ( .A(n3602), .B(n3727), .Z(n3729) );
  XOR U3770 ( .A(n3819), .B(n3820), .Z(n3602) );
  AND U3771 ( .A(n47), .B(n3821), .Z(n3820) );
  XNOR U3772 ( .A(n3822), .B(n3819), .Z(n3821) );
  AND U3773 ( .A(n3625), .B(n3628), .Z(n3727) );
  XOR U3774 ( .A(n3823), .B(n3778), .Z(n3628) );
  XNOR U3775 ( .A(p_input[320]), .B(p_input[512]), .Z(n3778) );
  XNOR U3776 ( .A(n3754), .B(n3753), .Z(n3823) );
  XNOR U3777 ( .A(n3824), .B(n3765), .Z(n3753) );
  XOR U3778 ( .A(n3739), .B(n3737), .Z(n3765) );
  XNOR U3779 ( .A(n3825), .B(n3744), .Z(n3737) );
  XOR U3780 ( .A(p_input[344]), .B(p_input[536]), .Z(n3744) );
  XOR U3781 ( .A(n3734), .B(n3743), .Z(n3825) );
  XOR U3782 ( .A(n3826), .B(n3740), .Z(n3743) );
  XOR U3783 ( .A(p_input[342]), .B(p_input[534]), .Z(n3740) );
  XOR U3784 ( .A(p_input[343]), .B(n1634), .Z(n3826) );
  XOR U3785 ( .A(p_input[338]), .B(p_input[530]), .Z(n3734) );
  XNOR U3786 ( .A(n3749), .B(n3748), .Z(n3739) );
  XOR U3787 ( .A(n3827), .B(n3745), .Z(n3748) );
  XOR U3788 ( .A(p_input[339]), .B(p_input[531]), .Z(n3745) );
  XOR U3789 ( .A(p_input[340]), .B(n1636), .Z(n3827) );
  XOR U3790 ( .A(p_input[341]), .B(p_input[533]), .Z(n3749) );
  XOR U3791 ( .A(n3764), .B(n3828), .Z(n3824) );
  IV U3792 ( .A(n3750), .Z(n3828) );
  XOR U3793 ( .A(p_input[321]), .B(p_input[513]), .Z(n3750) );
  XNOR U3794 ( .A(n3829), .B(n3772), .Z(n3764) );
  XNOR U3795 ( .A(n3760), .B(n3759), .Z(n3772) );
  XNOR U3796 ( .A(n3830), .B(n3756), .Z(n3759) );
  XNOR U3797 ( .A(p_input[346]), .B(p_input[538]), .Z(n3756) );
  XOR U3798 ( .A(p_input[347]), .B(n1640), .Z(n3830) );
  XOR U3799 ( .A(p_input[348]), .B(p_input[540]), .Z(n3760) );
  XOR U3800 ( .A(n3770), .B(n3831), .Z(n3829) );
  IV U3801 ( .A(n3761), .Z(n3831) );
  XOR U3802 ( .A(p_input[337]), .B(p_input[529]), .Z(n3761) );
  XNOR U3803 ( .A(n3832), .B(n3777), .Z(n3770) );
  XNOR U3804 ( .A(p_input[351]), .B(n1643), .Z(n3777) );
  XOR U3805 ( .A(n3767), .B(n3776), .Z(n3832) );
  XOR U3806 ( .A(n3833), .B(n3773), .Z(n3776) );
  XOR U3807 ( .A(p_input[349]), .B(p_input[541]), .Z(n3773) );
  XOR U3808 ( .A(p_input[350]), .B(n1645), .Z(n3833) );
  XOR U3809 ( .A(p_input[345]), .B(p_input[537]), .Z(n3767) );
  XOR U3810 ( .A(n3789), .B(n3788), .Z(n3754) );
  XNOR U3811 ( .A(n3834), .B(n3796), .Z(n3788) );
  XNOR U3812 ( .A(n3784), .B(n3783), .Z(n3796) );
  XNOR U3813 ( .A(n3835), .B(n3780), .Z(n3783) );
  XNOR U3814 ( .A(p_input[331]), .B(p_input[523]), .Z(n3780) );
  XOR U3815 ( .A(p_input[332]), .B(n1648), .Z(n3835) );
  XOR U3816 ( .A(p_input[333]), .B(p_input[525]), .Z(n3784) );
  XOR U3817 ( .A(n3794), .B(n3836), .Z(n3834) );
  IV U3818 ( .A(n3785), .Z(n3836) );
  XOR U3819 ( .A(p_input[322]), .B(p_input[514]), .Z(n3785) );
  XNOR U3820 ( .A(n3837), .B(n3801), .Z(n3794) );
  XNOR U3821 ( .A(p_input[336]), .B(n1651), .Z(n3801) );
  XOR U3822 ( .A(n3791), .B(n3800), .Z(n3837) );
  XOR U3823 ( .A(n3838), .B(n3797), .Z(n3800) );
  XOR U3824 ( .A(p_input[334]), .B(p_input[526]), .Z(n3797) );
  XOR U3825 ( .A(p_input[335]), .B(n1653), .Z(n3838) );
  XOR U3826 ( .A(p_input[330]), .B(p_input[522]), .Z(n3791) );
  XOR U3827 ( .A(n3808), .B(n3806), .Z(n3789) );
  XNOR U3828 ( .A(n3839), .B(n3813), .Z(n3806) );
  XOR U3829 ( .A(p_input[329]), .B(p_input[521]), .Z(n3813) );
  XOR U3830 ( .A(n3803), .B(n3812), .Z(n3839) );
  XOR U3831 ( .A(n3840), .B(n3809), .Z(n3812) );
  XOR U3832 ( .A(p_input[327]), .B(p_input[519]), .Z(n3809) );
  XOR U3833 ( .A(p_input[328]), .B(n1877), .Z(n3840) );
  XOR U3834 ( .A(p_input[323]), .B(p_input[515]), .Z(n3803) );
  XNOR U3835 ( .A(n3818), .B(n3817), .Z(n3808) );
  XOR U3836 ( .A(n3841), .B(n3814), .Z(n3817) );
  XOR U3837 ( .A(p_input[324]), .B(p_input[516]), .Z(n3814) );
  XOR U3838 ( .A(p_input[325]), .B(n1879), .Z(n3841) );
  XOR U3839 ( .A(p_input[326]), .B(p_input[518]), .Z(n3818) );
  XOR U3840 ( .A(n3842), .B(n3843), .Z(n3625) );
  AND U3841 ( .A(n47), .B(n3844), .Z(n3843) );
  XNOR U3842 ( .A(n3845), .B(n3842), .Z(n3844) );
  XNOR U3843 ( .A(n3846), .B(n3847), .Z(n47) );
  NOR U3844 ( .A(n3848), .B(n3849), .Z(n3847) );
  XOR U3845 ( .A(n3634), .B(n3846), .Z(n3849) );
  AND U3846 ( .A(n3850), .B(n3851), .Z(n3634) );
  NOR U3847 ( .A(n3846), .B(n3633), .Z(n3848) );
  AND U3848 ( .A(n3852), .B(n3853), .Z(n3633) );
  XOR U3849 ( .A(n3854), .B(n3855), .Z(n3846) );
  AND U3850 ( .A(n3856), .B(n3857), .Z(n3855) );
  XNOR U3851 ( .A(n3854), .B(n3852), .Z(n3857) );
  IV U3852 ( .A(n3651), .Z(n3852) );
  XOR U3853 ( .A(n3858), .B(n3859), .Z(n3651) );
  XOR U3854 ( .A(n3860), .B(n3853), .Z(n3859) );
  AND U3855 ( .A(n3678), .B(n3861), .Z(n3853) );
  AND U3856 ( .A(n3862), .B(n3863), .Z(n3860) );
  XOR U3857 ( .A(n3864), .B(n3858), .Z(n3862) );
  XNOR U3858 ( .A(n3648), .B(n3854), .Z(n3856) );
  XOR U3859 ( .A(n3865), .B(n3866), .Z(n3648) );
  AND U3860 ( .A(n51), .B(n3867), .Z(n3866) );
  XOR U3861 ( .A(n3868), .B(n3865), .Z(n3867) );
  XOR U3862 ( .A(n3869), .B(n3870), .Z(n3854) );
  AND U3863 ( .A(n3871), .B(n3872), .Z(n3870) );
  XNOR U3864 ( .A(n3869), .B(n3678), .Z(n3872) );
  XOR U3865 ( .A(n3873), .B(n3863), .Z(n3678) );
  XNOR U3866 ( .A(n3874), .B(n3858), .Z(n3863) );
  XOR U3867 ( .A(n3875), .B(n3876), .Z(n3858) );
  AND U3868 ( .A(n3877), .B(n3878), .Z(n3876) );
  XOR U3869 ( .A(n3879), .B(n3875), .Z(n3877) );
  XNOR U3870 ( .A(n3880), .B(n3881), .Z(n3874) );
  AND U3871 ( .A(n3882), .B(n3883), .Z(n3881) );
  XOR U3872 ( .A(n3880), .B(n3884), .Z(n3882) );
  XNOR U3873 ( .A(n3864), .B(n3861), .Z(n3873) );
  AND U3874 ( .A(n3885), .B(n3886), .Z(n3861) );
  XOR U3875 ( .A(n3887), .B(n3888), .Z(n3864) );
  AND U3876 ( .A(n3889), .B(n3890), .Z(n3888) );
  XOR U3877 ( .A(n3887), .B(n3891), .Z(n3889) );
  XNOR U3878 ( .A(n3675), .B(n3869), .Z(n3871) );
  XOR U3879 ( .A(n3892), .B(n3893), .Z(n3675) );
  AND U3880 ( .A(n51), .B(n3894), .Z(n3893) );
  XNOR U3881 ( .A(n3895), .B(n3892), .Z(n3894) );
  XOR U3882 ( .A(n3896), .B(n3897), .Z(n3869) );
  AND U3883 ( .A(n3898), .B(n3899), .Z(n3897) );
  XNOR U3884 ( .A(n3896), .B(n3885), .Z(n3899) );
  IV U3885 ( .A(n3726), .Z(n3885) );
  XNOR U3886 ( .A(n3900), .B(n3878), .Z(n3726) );
  XNOR U3887 ( .A(n3901), .B(n3884), .Z(n3878) );
  XOR U3888 ( .A(n3902), .B(n3903), .Z(n3884) );
  AND U3889 ( .A(n3904), .B(n3905), .Z(n3903) );
  XOR U3890 ( .A(n3902), .B(n3906), .Z(n3904) );
  XNOR U3891 ( .A(n3883), .B(n3875), .Z(n3901) );
  XOR U3892 ( .A(n3907), .B(n3908), .Z(n3875) );
  AND U3893 ( .A(n3909), .B(n3910), .Z(n3908) );
  XNOR U3894 ( .A(n3911), .B(n3907), .Z(n3909) );
  XNOR U3895 ( .A(n3912), .B(n3880), .Z(n3883) );
  XOR U3896 ( .A(n3913), .B(n3914), .Z(n3880) );
  AND U3897 ( .A(n3915), .B(n3916), .Z(n3914) );
  XOR U3898 ( .A(n3913), .B(n3917), .Z(n3915) );
  XNOR U3899 ( .A(n3918), .B(n3919), .Z(n3912) );
  AND U3900 ( .A(n3920), .B(n3921), .Z(n3919) );
  XNOR U3901 ( .A(n3918), .B(n3922), .Z(n3920) );
  XNOR U3902 ( .A(n3879), .B(n3886), .Z(n3900) );
  AND U3903 ( .A(n3822), .B(n3923), .Z(n3886) );
  XOR U3904 ( .A(n3891), .B(n3890), .Z(n3879) );
  XNOR U3905 ( .A(n3924), .B(n3887), .Z(n3890) );
  XOR U3906 ( .A(n3925), .B(n3926), .Z(n3887) );
  AND U3907 ( .A(n3927), .B(n3928), .Z(n3926) );
  XOR U3908 ( .A(n3925), .B(n3929), .Z(n3927) );
  XNOR U3909 ( .A(n3930), .B(n3931), .Z(n3924) );
  AND U3910 ( .A(n3932), .B(n3933), .Z(n3931) );
  XOR U3911 ( .A(n3930), .B(n3934), .Z(n3932) );
  XOR U3912 ( .A(n3935), .B(n3936), .Z(n3891) );
  AND U3913 ( .A(n3937), .B(n3938), .Z(n3936) );
  XOR U3914 ( .A(n3935), .B(n3939), .Z(n3937) );
  XNOR U3915 ( .A(n3723), .B(n3896), .Z(n3898) );
  XOR U3916 ( .A(n3940), .B(n3941), .Z(n3723) );
  AND U3917 ( .A(n51), .B(n3942), .Z(n3941) );
  XOR U3918 ( .A(n3943), .B(n3940), .Z(n3942) );
  XOR U3919 ( .A(n3944), .B(n3945), .Z(n3896) );
  AND U3920 ( .A(n3946), .B(n3947), .Z(n3945) );
  XNOR U3921 ( .A(n3944), .B(n3822), .Z(n3947) );
  XOR U3922 ( .A(n3948), .B(n3910), .Z(n3822) );
  XNOR U3923 ( .A(n3949), .B(n3917), .Z(n3910) );
  XOR U3924 ( .A(n3906), .B(n3905), .Z(n3917) );
  XNOR U3925 ( .A(n3950), .B(n3902), .Z(n3905) );
  XOR U3926 ( .A(n3951), .B(n3952), .Z(n3902) );
  AND U3927 ( .A(n3953), .B(n3954), .Z(n3952) );
  XNOR U3928 ( .A(n3955), .B(n3956), .Z(n3953) );
  IV U3929 ( .A(n3951), .Z(n3955) );
  XNOR U3930 ( .A(n3957), .B(n3958), .Z(n3950) );
  NOR U3931 ( .A(n3959), .B(n3960), .Z(n3958) );
  XNOR U3932 ( .A(n3957), .B(n3961), .Z(n3959) );
  XOR U3933 ( .A(n3962), .B(n3963), .Z(n3906) );
  NOR U3934 ( .A(n3964), .B(n3965), .Z(n3963) );
  XNOR U3935 ( .A(n3962), .B(n3966), .Z(n3964) );
  XNOR U3936 ( .A(n3916), .B(n3907), .Z(n3949) );
  XOR U3937 ( .A(n3967), .B(n3968), .Z(n3907) );
  AND U3938 ( .A(n3969), .B(n3970), .Z(n3968) );
  XOR U3939 ( .A(n3967), .B(n3971), .Z(n3969) );
  XOR U3940 ( .A(n3972), .B(n3922), .Z(n3916) );
  XOR U3941 ( .A(n3973), .B(n3974), .Z(n3922) );
  NOR U3942 ( .A(n3975), .B(n3976), .Z(n3974) );
  XOR U3943 ( .A(n3973), .B(n3977), .Z(n3975) );
  XNOR U3944 ( .A(n3921), .B(n3913), .Z(n3972) );
  XOR U3945 ( .A(n3978), .B(n3979), .Z(n3913) );
  AND U3946 ( .A(n3980), .B(n3981), .Z(n3979) );
  XOR U3947 ( .A(n3978), .B(n3982), .Z(n3980) );
  XNOR U3948 ( .A(n3983), .B(n3918), .Z(n3921) );
  XOR U3949 ( .A(n3984), .B(n3985), .Z(n3918) );
  AND U3950 ( .A(n3986), .B(n3987), .Z(n3985) );
  XNOR U3951 ( .A(n3988), .B(n3989), .Z(n3986) );
  IV U3952 ( .A(n3984), .Z(n3988) );
  XNOR U3953 ( .A(n3990), .B(n3991), .Z(n3983) );
  NOR U3954 ( .A(n3992), .B(n3993), .Z(n3991) );
  XNOR U3955 ( .A(n3990), .B(n3994), .Z(n3992) );
  XOR U3956 ( .A(n3911), .B(n3923), .Z(n3948) );
  NOR U3957 ( .A(n3845), .B(n3995), .Z(n3923) );
  XNOR U3958 ( .A(n3929), .B(n3928), .Z(n3911) );
  XNOR U3959 ( .A(n3996), .B(n3934), .Z(n3928) );
  XNOR U3960 ( .A(n3997), .B(n3998), .Z(n3934) );
  NOR U3961 ( .A(n3999), .B(n4000), .Z(n3998) );
  XOR U3962 ( .A(n3997), .B(n4001), .Z(n3999) );
  XNOR U3963 ( .A(n3933), .B(n3925), .Z(n3996) );
  XOR U3964 ( .A(n4002), .B(n4003), .Z(n3925) );
  AND U3965 ( .A(n4004), .B(n4005), .Z(n4003) );
  XOR U3966 ( .A(n4002), .B(n4006), .Z(n4004) );
  XNOR U3967 ( .A(n4007), .B(n3930), .Z(n3933) );
  XOR U3968 ( .A(n4008), .B(n4009), .Z(n3930) );
  AND U3969 ( .A(n4010), .B(n4011), .Z(n4009) );
  XNOR U3970 ( .A(n4012), .B(n4013), .Z(n4010) );
  IV U3971 ( .A(n4008), .Z(n4012) );
  XNOR U3972 ( .A(n4014), .B(n4015), .Z(n4007) );
  NOR U3973 ( .A(n4016), .B(n4017), .Z(n4015) );
  XNOR U3974 ( .A(n4014), .B(n4018), .Z(n4016) );
  XOR U3975 ( .A(n3939), .B(n3938), .Z(n3929) );
  XNOR U3976 ( .A(n4019), .B(n3935), .Z(n3938) );
  XOR U3977 ( .A(n4020), .B(n4021), .Z(n3935) );
  AND U3978 ( .A(n4022), .B(n4023), .Z(n4021) );
  XNOR U3979 ( .A(n4024), .B(n4025), .Z(n4022) );
  IV U3980 ( .A(n4020), .Z(n4024) );
  XNOR U3981 ( .A(n4026), .B(n4027), .Z(n4019) );
  NOR U3982 ( .A(n4028), .B(n4029), .Z(n4027) );
  XNOR U3983 ( .A(n4026), .B(n4030), .Z(n4028) );
  XOR U3984 ( .A(n4031), .B(n4032), .Z(n3939) );
  NOR U3985 ( .A(n4033), .B(n4034), .Z(n4032) );
  XNOR U3986 ( .A(n4031), .B(n4035), .Z(n4033) );
  XNOR U3987 ( .A(n3819), .B(n3944), .Z(n3946) );
  XOR U3988 ( .A(n4036), .B(n4037), .Z(n3819) );
  AND U3989 ( .A(n51), .B(n4038), .Z(n4037) );
  XNOR U3990 ( .A(n4039), .B(n4036), .Z(n4038) );
  AND U3991 ( .A(n3842), .B(n3845), .Z(n3944) );
  XOR U3992 ( .A(n4040), .B(n3995), .Z(n3845) );
  XNOR U3993 ( .A(p_input[352]), .B(p_input[512]), .Z(n3995) );
  XNOR U3994 ( .A(n3971), .B(n3970), .Z(n4040) );
  XNOR U3995 ( .A(n4041), .B(n3982), .Z(n3970) );
  XOR U3996 ( .A(n3956), .B(n3954), .Z(n3982) );
  XNOR U3997 ( .A(n4042), .B(n3961), .Z(n3954) );
  XOR U3998 ( .A(p_input[376]), .B(p_input[536]), .Z(n3961) );
  XOR U3999 ( .A(n3951), .B(n3960), .Z(n4042) );
  XOR U4000 ( .A(n4043), .B(n3957), .Z(n3960) );
  XOR U4001 ( .A(p_input[374]), .B(p_input[534]), .Z(n3957) );
  XOR U4002 ( .A(p_input[375]), .B(n1634), .Z(n4043) );
  XOR U4003 ( .A(p_input[370]), .B(p_input[530]), .Z(n3951) );
  XNOR U4004 ( .A(n3966), .B(n3965), .Z(n3956) );
  XOR U4005 ( .A(n4044), .B(n3962), .Z(n3965) );
  XOR U4006 ( .A(p_input[371]), .B(p_input[531]), .Z(n3962) );
  XOR U4007 ( .A(p_input[372]), .B(n1636), .Z(n4044) );
  XOR U4008 ( .A(p_input[373]), .B(p_input[533]), .Z(n3966) );
  XOR U4009 ( .A(n3981), .B(n4045), .Z(n4041) );
  IV U4010 ( .A(n3967), .Z(n4045) );
  XOR U4011 ( .A(p_input[353]), .B(p_input[513]), .Z(n3967) );
  XNOR U4012 ( .A(n4046), .B(n3989), .Z(n3981) );
  XNOR U4013 ( .A(n3977), .B(n3976), .Z(n3989) );
  XNOR U4014 ( .A(n4047), .B(n3973), .Z(n3976) );
  XNOR U4015 ( .A(p_input[378]), .B(p_input[538]), .Z(n3973) );
  XOR U4016 ( .A(p_input[379]), .B(n1640), .Z(n4047) );
  XOR U4017 ( .A(p_input[380]), .B(p_input[540]), .Z(n3977) );
  XOR U4018 ( .A(n3987), .B(n4048), .Z(n4046) );
  IV U4019 ( .A(n3978), .Z(n4048) );
  XOR U4020 ( .A(p_input[369]), .B(p_input[529]), .Z(n3978) );
  XNOR U4021 ( .A(n4049), .B(n3994), .Z(n3987) );
  XNOR U4022 ( .A(p_input[383]), .B(n1643), .Z(n3994) );
  XOR U4023 ( .A(n3984), .B(n3993), .Z(n4049) );
  XOR U4024 ( .A(n4050), .B(n3990), .Z(n3993) );
  XOR U4025 ( .A(p_input[381]), .B(p_input[541]), .Z(n3990) );
  XOR U4026 ( .A(p_input[382]), .B(n1645), .Z(n4050) );
  XOR U4027 ( .A(p_input[377]), .B(p_input[537]), .Z(n3984) );
  XOR U4028 ( .A(n4006), .B(n4005), .Z(n3971) );
  XNOR U4029 ( .A(n4051), .B(n4013), .Z(n4005) );
  XNOR U4030 ( .A(n4001), .B(n4000), .Z(n4013) );
  XNOR U4031 ( .A(n4052), .B(n3997), .Z(n4000) );
  XNOR U4032 ( .A(p_input[363]), .B(p_input[523]), .Z(n3997) );
  XOR U4033 ( .A(p_input[364]), .B(n1648), .Z(n4052) );
  XOR U4034 ( .A(p_input[365]), .B(p_input[525]), .Z(n4001) );
  XOR U4035 ( .A(n4011), .B(n4053), .Z(n4051) );
  IV U4036 ( .A(n4002), .Z(n4053) );
  XOR U4037 ( .A(p_input[354]), .B(p_input[514]), .Z(n4002) );
  XNOR U4038 ( .A(n4054), .B(n4018), .Z(n4011) );
  XNOR U4039 ( .A(p_input[368]), .B(n1651), .Z(n4018) );
  XOR U4040 ( .A(n4008), .B(n4017), .Z(n4054) );
  XOR U4041 ( .A(n4055), .B(n4014), .Z(n4017) );
  XOR U4042 ( .A(p_input[366]), .B(p_input[526]), .Z(n4014) );
  XOR U4043 ( .A(p_input[367]), .B(n1653), .Z(n4055) );
  XOR U4044 ( .A(p_input[362]), .B(p_input[522]), .Z(n4008) );
  XOR U4045 ( .A(n4025), .B(n4023), .Z(n4006) );
  XNOR U4046 ( .A(n4056), .B(n4030), .Z(n4023) );
  XOR U4047 ( .A(p_input[361]), .B(p_input[521]), .Z(n4030) );
  XOR U4048 ( .A(n4020), .B(n4029), .Z(n4056) );
  XOR U4049 ( .A(n4057), .B(n4026), .Z(n4029) );
  XOR U4050 ( .A(p_input[359]), .B(p_input[519]), .Z(n4026) );
  XOR U4051 ( .A(p_input[360]), .B(n1877), .Z(n4057) );
  XOR U4052 ( .A(p_input[355]), .B(p_input[515]), .Z(n4020) );
  XNOR U4053 ( .A(n4035), .B(n4034), .Z(n4025) );
  XOR U4054 ( .A(n4058), .B(n4031), .Z(n4034) );
  XOR U4055 ( .A(p_input[356]), .B(p_input[516]), .Z(n4031) );
  XOR U4056 ( .A(p_input[357]), .B(n1879), .Z(n4058) );
  XOR U4057 ( .A(p_input[358]), .B(p_input[518]), .Z(n4035) );
  XOR U4058 ( .A(n4059), .B(n4060), .Z(n3842) );
  AND U4059 ( .A(n51), .B(n4061), .Z(n4060) );
  XNOR U4060 ( .A(n4062), .B(n4059), .Z(n4061) );
  XNOR U4061 ( .A(n4063), .B(n4064), .Z(n51) );
  NOR U4062 ( .A(n4065), .B(n4066), .Z(n4064) );
  XOR U4063 ( .A(n3851), .B(n4063), .Z(n4066) );
  AND U4064 ( .A(n4067), .B(n4068), .Z(n3851) );
  NOR U4065 ( .A(n4063), .B(n3850), .Z(n4065) );
  AND U4066 ( .A(n4069), .B(n4070), .Z(n3850) );
  XOR U4067 ( .A(n4071), .B(n4072), .Z(n4063) );
  AND U4068 ( .A(n4073), .B(n4074), .Z(n4072) );
  XNOR U4069 ( .A(n4071), .B(n4069), .Z(n4074) );
  IV U4070 ( .A(n3868), .Z(n4069) );
  XOR U4071 ( .A(n4075), .B(n4076), .Z(n3868) );
  XOR U4072 ( .A(n4077), .B(n4070), .Z(n4076) );
  AND U4073 ( .A(n3895), .B(n4078), .Z(n4070) );
  AND U4074 ( .A(n4079), .B(n4080), .Z(n4077) );
  XOR U4075 ( .A(n4081), .B(n4075), .Z(n4079) );
  XNOR U4076 ( .A(n3865), .B(n4071), .Z(n4073) );
  XOR U4077 ( .A(n4082), .B(n4083), .Z(n3865) );
  AND U4078 ( .A(n55), .B(n4084), .Z(n4083) );
  XOR U4079 ( .A(n4085), .B(n4082), .Z(n4084) );
  XOR U4080 ( .A(n4086), .B(n4087), .Z(n4071) );
  AND U4081 ( .A(n4088), .B(n4089), .Z(n4087) );
  XNOR U4082 ( .A(n4086), .B(n3895), .Z(n4089) );
  XOR U4083 ( .A(n4090), .B(n4080), .Z(n3895) );
  XNOR U4084 ( .A(n4091), .B(n4075), .Z(n4080) );
  XOR U4085 ( .A(n4092), .B(n4093), .Z(n4075) );
  AND U4086 ( .A(n4094), .B(n4095), .Z(n4093) );
  XOR U4087 ( .A(n4096), .B(n4092), .Z(n4094) );
  XNOR U4088 ( .A(n4097), .B(n4098), .Z(n4091) );
  AND U4089 ( .A(n4099), .B(n4100), .Z(n4098) );
  XOR U4090 ( .A(n4097), .B(n4101), .Z(n4099) );
  XNOR U4091 ( .A(n4081), .B(n4078), .Z(n4090) );
  AND U4092 ( .A(n4102), .B(n4103), .Z(n4078) );
  XOR U4093 ( .A(n4104), .B(n4105), .Z(n4081) );
  AND U4094 ( .A(n4106), .B(n4107), .Z(n4105) );
  XOR U4095 ( .A(n4104), .B(n4108), .Z(n4106) );
  XNOR U4096 ( .A(n3892), .B(n4086), .Z(n4088) );
  XOR U4097 ( .A(n4109), .B(n4110), .Z(n3892) );
  AND U4098 ( .A(n55), .B(n4111), .Z(n4110) );
  XNOR U4099 ( .A(n4112), .B(n4109), .Z(n4111) );
  XOR U4100 ( .A(n4113), .B(n4114), .Z(n4086) );
  AND U4101 ( .A(n4115), .B(n4116), .Z(n4114) );
  XNOR U4102 ( .A(n4113), .B(n4102), .Z(n4116) );
  IV U4103 ( .A(n3943), .Z(n4102) );
  XNOR U4104 ( .A(n4117), .B(n4095), .Z(n3943) );
  XNOR U4105 ( .A(n4118), .B(n4101), .Z(n4095) );
  XOR U4106 ( .A(n4119), .B(n4120), .Z(n4101) );
  AND U4107 ( .A(n4121), .B(n4122), .Z(n4120) );
  XOR U4108 ( .A(n4119), .B(n4123), .Z(n4121) );
  XNOR U4109 ( .A(n4100), .B(n4092), .Z(n4118) );
  XOR U4110 ( .A(n4124), .B(n4125), .Z(n4092) );
  AND U4111 ( .A(n4126), .B(n4127), .Z(n4125) );
  XNOR U4112 ( .A(n4128), .B(n4124), .Z(n4126) );
  XNOR U4113 ( .A(n4129), .B(n4097), .Z(n4100) );
  XOR U4114 ( .A(n4130), .B(n4131), .Z(n4097) );
  AND U4115 ( .A(n4132), .B(n4133), .Z(n4131) );
  XOR U4116 ( .A(n4130), .B(n4134), .Z(n4132) );
  XNOR U4117 ( .A(n4135), .B(n4136), .Z(n4129) );
  AND U4118 ( .A(n4137), .B(n4138), .Z(n4136) );
  XNOR U4119 ( .A(n4135), .B(n4139), .Z(n4137) );
  XNOR U4120 ( .A(n4096), .B(n4103), .Z(n4117) );
  AND U4121 ( .A(n4039), .B(n4140), .Z(n4103) );
  XOR U4122 ( .A(n4108), .B(n4107), .Z(n4096) );
  XNOR U4123 ( .A(n4141), .B(n4104), .Z(n4107) );
  XOR U4124 ( .A(n4142), .B(n4143), .Z(n4104) );
  AND U4125 ( .A(n4144), .B(n4145), .Z(n4143) );
  XOR U4126 ( .A(n4142), .B(n4146), .Z(n4144) );
  XNOR U4127 ( .A(n4147), .B(n4148), .Z(n4141) );
  AND U4128 ( .A(n4149), .B(n4150), .Z(n4148) );
  XOR U4129 ( .A(n4147), .B(n4151), .Z(n4149) );
  XOR U4130 ( .A(n4152), .B(n4153), .Z(n4108) );
  AND U4131 ( .A(n4154), .B(n4155), .Z(n4153) );
  XOR U4132 ( .A(n4152), .B(n4156), .Z(n4154) );
  XNOR U4133 ( .A(n3940), .B(n4113), .Z(n4115) );
  XOR U4134 ( .A(n4157), .B(n4158), .Z(n3940) );
  AND U4135 ( .A(n55), .B(n4159), .Z(n4158) );
  XOR U4136 ( .A(n4160), .B(n4157), .Z(n4159) );
  XOR U4137 ( .A(n4161), .B(n4162), .Z(n4113) );
  AND U4138 ( .A(n4163), .B(n4164), .Z(n4162) );
  XNOR U4139 ( .A(n4161), .B(n4039), .Z(n4164) );
  XOR U4140 ( .A(n4165), .B(n4127), .Z(n4039) );
  XNOR U4141 ( .A(n4166), .B(n4134), .Z(n4127) );
  XOR U4142 ( .A(n4123), .B(n4122), .Z(n4134) );
  XNOR U4143 ( .A(n4167), .B(n4119), .Z(n4122) );
  XOR U4144 ( .A(n4168), .B(n4169), .Z(n4119) );
  AND U4145 ( .A(n4170), .B(n4171), .Z(n4169) );
  XNOR U4146 ( .A(n4172), .B(n4173), .Z(n4170) );
  IV U4147 ( .A(n4168), .Z(n4172) );
  XNOR U4148 ( .A(n4174), .B(n4175), .Z(n4167) );
  NOR U4149 ( .A(n4176), .B(n4177), .Z(n4175) );
  XNOR U4150 ( .A(n4174), .B(n4178), .Z(n4176) );
  XOR U4151 ( .A(n4179), .B(n4180), .Z(n4123) );
  NOR U4152 ( .A(n4181), .B(n4182), .Z(n4180) );
  XNOR U4153 ( .A(n4179), .B(n4183), .Z(n4181) );
  XNOR U4154 ( .A(n4133), .B(n4124), .Z(n4166) );
  XOR U4155 ( .A(n4184), .B(n4185), .Z(n4124) );
  AND U4156 ( .A(n4186), .B(n4187), .Z(n4185) );
  XOR U4157 ( .A(n4184), .B(n4188), .Z(n4186) );
  XOR U4158 ( .A(n4189), .B(n4139), .Z(n4133) );
  XOR U4159 ( .A(n4190), .B(n4191), .Z(n4139) );
  NOR U4160 ( .A(n4192), .B(n4193), .Z(n4191) );
  XOR U4161 ( .A(n4190), .B(n4194), .Z(n4192) );
  XNOR U4162 ( .A(n4138), .B(n4130), .Z(n4189) );
  XOR U4163 ( .A(n4195), .B(n4196), .Z(n4130) );
  AND U4164 ( .A(n4197), .B(n4198), .Z(n4196) );
  XOR U4165 ( .A(n4195), .B(n4199), .Z(n4197) );
  XNOR U4166 ( .A(n4200), .B(n4135), .Z(n4138) );
  XOR U4167 ( .A(n4201), .B(n4202), .Z(n4135) );
  AND U4168 ( .A(n4203), .B(n4204), .Z(n4202) );
  XNOR U4169 ( .A(n4205), .B(n4206), .Z(n4203) );
  IV U4170 ( .A(n4201), .Z(n4205) );
  XNOR U4171 ( .A(n4207), .B(n4208), .Z(n4200) );
  NOR U4172 ( .A(n4209), .B(n4210), .Z(n4208) );
  XNOR U4173 ( .A(n4207), .B(n4211), .Z(n4209) );
  XOR U4174 ( .A(n4128), .B(n4140), .Z(n4165) );
  NOR U4175 ( .A(n4062), .B(n4212), .Z(n4140) );
  XNOR U4176 ( .A(n4146), .B(n4145), .Z(n4128) );
  XNOR U4177 ( .A(n4213), .B(n4151), .Z(n4145) );
  XNOR U4178 ( .A(n4214), .B(n4215), .Z(n4151) );
  NOR U4179 ( .A(n4216), .B(n4217), .Z(n4215) );
  XOR U4180 ( .A(n4214), .B(n4218), .Z(n4216) );
  XNOR U4181 ( .A(n4150), .B(n4142), .Z(n4213) );
  XOR U4182 ( .A(n4219), .B(n4220), .Z(n4142) );
  AND U4183 ( .A(n4221), .B(n4222), .Z(n4220) );
  XOR U4184 ( .A(n4219), .B(n4223), .Z(n4221) );
  XNOR U4185 ( .A(n4224), .B(n4147), .Z(n4150) );
  XOR U4186 ( .A(n4225), .B(n4226), .Z(n4147) );
  AND U4187 ( .A(n4227), .B(n4228), .Z(n4226) );
  XNOR U4188 ( .A(n4229), .B(n4230), .Z(n4227) );
  IV U4189 ( .A(n4225), .Z(n4229) );
  XNOR U4190 ( .A(n4231), .B(n4232), .Z(n4224) );
  NOR U4191 ( .A(n4233), .B(n4234), .Z(n4232) );
  XNOR U4192 ( .A(n4231), .B(n4235), .Z(n4233) );
  XOR U4193 ( .A(n4156), .B(n4155), .Z(n4146) );
  XNOR U4194 ( .A(n4236), .B(n4152), .Z(n4155) );
  XOR U4195 ( .A(n4237), .B(n4238), .Z(n4152) );
  AND U4196 ( .A(n4239), .B(n4240), .Z(n4238) );
  XNOR U4197 ( .A(n4241), .B(n4242), .Z(n4239) );
  IV U4198 ( .A(n4237), .Z(n4241) );
  XNOR U4199 ( .A(n4243), .B(n4244), .Z(n4236) );
  NOR U4200 ( .A(n4245), .B(n4246), .Z(n4244) );
  XNOR U4201 ( .A(n4243), .B(n4247), .Z(n4245) );
  XOR U4202 ( .A(n4248), .B(n4249), .Z(n4156) );
  NOR U4203 ( .A(n4250), .B(n4251), .Z(n4249) );
  XNOR U4204 ( .A(n4248), .B(n4252), .Z(n4250) );
  XNOR U4205 ( .A(n4036), .B(n4161), .Z(n4163) );
  XOR U4206 ( .A(n4253), .B(n4254), .Z(n4036) );
  AND U4207 ( .A(n55), .B(n4255), .Z(n4254) );
  XNOR U4208 ( .A(n4256), .B(n4253), .Z(n4255) );
  AND U4209 ( .A(n4059), .B(n4062), .Z(n4161) );
  XOR U4210 ( .A(n4257), .B(n4212), .Z(n4062) );
  XNOR U4211 ( .A(p_input[384]), .B(p_input[512]), .Z(n4212) );
  XNOR U4212 ( .A(n4188), .B(n4187), .Z(n4257) );
  XNOR U4213 ( .A(n4258), .B(n4199), .Z(n4187) );
  XOR U4214 ( .A(n4173), .B(n4171), .Z(n4199) );
  XNOR U4215 ( .A(n4259), .B(n4178), .Z(n4171) );
  XOR U4216 ( .A(p_input[408]), .B(p_input[536]), .Z(n4178) );
  XOR U4217 ( .A(n4168), .B(n4177), .Z(n4259) );
  XOR U4218 ( .A(n4260), .B(n4174), .Z(n4177) );
  XOR U4219 ( .A(p_input[406]), .B(p_input[534]), .Z(n4174) );
  XOR U4220 ( .A(p_input[407]), .B(n1634), .Z(n4260) );
  XOR U4221 ( .A(p_input[402]), .B(p_input[530]), .Z(n4168) );
  XNOR U4222 ( .A(n4183), .B(n4182), .Z(n4173) );
  XOR U4223 ( .A(n4261), .B(n4179), .Z(n4182) );
  XOR U4224 ( .A(p_input[403]), .B(p_input[531]), .Z(n4179) );
  XOR U4225 ( .A(p_input[404]), .B(n1636), .Z(n4261) );
  XOR U4226 ( .A(p_input[405]), .B(p_input[533]), .Z(n4183) );
  XOR U4227 ( .A(n4198), .B(n4262), .Z(n4258) );
  IV U4228 ( .A(n4184), .Z(n4262) );
  XOR U4229 ( .A(p_input[385]), .B(p_input[513]), .Z(n4184) );
  XNOR U4230 ( .A(n4263), .B(n4206), .Z(n4198) );
  XNOR U4231 ( .A(n4194), .B(n4193), .Z(n4206) );
  XNOR U4232 ( .A(n4264), .B(n4190), .Z(n4193) );
  XNOR U4233 ( .A(p_input[410]), .B(p_input[538]), .Z(n4190) );
  XOR U4234 ( .A(p_input[411]), .B(n1640), .Z(n4264) );
  XOR U4235 ( .A(p_input[412]), .B(p_input[540]), .Z(n4194) );
  XOR U4236 ( .A(n4204), .B(n4265), .Z(n4263) );
  IV U4237 ( .A(n4195), .Z(n4265) );
  XOR U4238 ( .A(p_input[401]), .B(p_input[529]), .Z(n4195) );
  XNOR U4239 ( .A(n4266), .B(n4211), .Z(n4204) );
  XNOR U4240 ( .A(p_input[415]), .B(n1643), .Z(n4211) );
  XOR U4241 ( .A(n4201), .B(n4210), .Z(n4266) );
  XOR U4242 ( .A(n4267), .B(n4207), .Z(n4210) );
  XOR U4243 ( .A(p_input[413]), .B(p_input[541]), .Z(n4207) );
  XOR U4244 ( .A(p_input[414]), .B(n1645), .Z(n4267) );
  XOR U4245 ( .A(p_input[409]), .B(p_input[537]), .Z(n4201) );
  XOR U4246 ( .A(n4223), .B(n4222), .Z(n4188) );
  XNOR U4247 ( .A(n4268), .B(n4230), .Z(n4222) );
  XNOR U4248 ( .A(n4218), .B(n4217), .Z(n4230) );
  XNOR U4249 ( .A(n4269), .B(n4214), .Z(n4217) );
  XNOR U4250 ( .A(p_input[395]), .B(p_input[523]), .Z(n4214) );
  XOR U4251 ( .A(p_input[396]), .B(n1648), .Z(n4269) );
  XOR U4252 ( .A(p_input[397]), .B(p_input[525]), .Z(n4218) );
  XOR U4253 ( .A(n4228), .B(n4270), .Z(n4268) );
  IV U4254 ( .A(n4219), .Z(n4270) );
  XOR U4255 ( .A(p_input[386]), .B(p_input[514]), .Z(n4219) );
  XNOR U4256 ( .A(n4271), .B(n4235), .Z(n4228) );
  XNOR U4257 ( .A(p_input[400]), .B(n1651), .Z(n4235) );
  XOR U4258 ( .A(n4225), .B(n4234), .Z(n4271) );
  XOR U4259 ( .A(n4272), .B(n4231), .Z(n4234) );
  XOR U4260 ( .A(p_input[398]), .B(p_input[526]), .Z(n4231) );
  XOR U4261 ( .A(p_input[399]), .B(n1653), .Z(n4272) );
  XOR U4262 ( .A(p_input[394]), .B(p_input[522]), .Z(n4225) );
  XOR U4263 ( .A(n4242), .B(n4240), .Z(n4223) );
  XNOR U4264 ( .A(n4273), .B(n4247), .Z(n4240) );
  XOR U4265 ( .A(p_input[393]), .B(p_input[521]), .Z(n4247) );
  XOR U4266 ( .A(n4237), .B(n4246), .Z(n4273) );
  XOR U4267 ( .A(n4274), .B(n4243), .Z(n4246) );
  XOR U4268 ( .A(p_input[391]), .B(p_input[519]), .Z(n4243) );
  XOR U4269 ( .A(p_input[392]), .B(n1877), .Z(n4274) );
  XOR U4270 ( .A(p_input[387]), .B(p_input[515]), .Z(n4237) );
  XNOR U4271 ( .A(n4252), .B(n4251), .Z(n4242) );
  XOR U4272 ( .A(n4275), .B(n4248), .Z(n4251) );
  XOR U4273 ( .A(p_input[388]), .B(p_input[516]), .Z(n4248) );
  XOR U4274 ( .A(p_input[389]), .B(n1879), .Z(n4275) );
  XOR U4275 ( .A(p_input[390]), .B(p_input[518]), .Z(n4252) );
  XOR U4276 ( .A(n4276), .B(n4277), .Z(n4059) );
  AND U4277 ( .A(n55), .B(n4278), .Z(n4277) );
  XNOR U4278 ( .A(n4279), .B(n4276), .Z(n4278) );
  XNOR U4279 ( .A(n4280), .B(n4281), .Z(n55) );
  NOR U4280 ( .A(n4282), .B(n4283), .Z(n4281) );
  XOR U4281 ( .A(n4068), .B(n4280), .Z(n4283) );
  AND U4282 ( .A(n4284), .B(n4285), .Z(n4068) );
  NOR U4283 ( .A(n4280), .B(n4067), .Z(n4282) );
  AND U4284 ( .A(n4286), .B(n4287), .Z(n4067) );
  XOR U4285 ( .A(n4288), .B(n4289), .Z(n4280) );
  AND U4286 ( .A(n4290), .B(n4291), .Z(n4289) );
  XNOR U4287 ( .A(n4288), .B(n4286), .Z(n4291) );
  IV U4288 ( .A(n4085), .Z(n4286) );
  XOR U4289 ( .A(n4292), .B(n4293), .Z(n4085) );
  XOR U4290 ( .A(n4294), .B(n4287), .Z(n4293) );
  AND U4291 ( .A(n4112), .B(n4295), .Z(n4287) );
  AND U4292 ( .A(n4296), .B(n4297), .Z(n4294) );
  XOR U4293 ( .A(n4298), .B(n4292), .Z(n4296) );
  XNOR U4294 ( .A(n4082), .B(n4288), .Z(n4290) );
  XNOR U4295 ( .A(n4299), .B(n4300), .Z(n4082) );
  AND U4296 ( .A(n58), .B(n4301), .Z(n4300) );
  XNOR U4297 ( .A(n4302), .B(n4299), .Z(n4301) );
  XOR U4298 ( .A(n4303), .B(n4304), .Z(n4288) );
  AND U4299 ( .A(n4305), .B(n4306), .Z(n4304) );
  XNOR U4300 ( .A(n4303), .B(n4112), .Z(n4306) );
  XOR U4301 ( .A(n4307), .B(n4297), .Z(n4112) );
  XNOR U4302 ( .A(n4308), .B(n4292), .Z(n4297) );
  XOR U4303 ( .A(n4309), .B(n4310), .Z(n4292) );
  AND U4304 ( .A(n4311), .B(n4312), .Z(n4310) );
  XOR U4305 ( .A(n4313), .B(n4309), .Z(n4311) );
  XNOR U4306 ( .A(n4314), .B(n4315), .Z(n4308) );
  AND U4307 ( .A(n4316), .B(n4317), .Z(n4315) );
  XOR U4308 ( .A(n4314), .B(n4318), .Z(n4316) );
  XNOR U4309 ( .A(n4298), .B(n4295), .Z(n4307) );
  AND U4310 ( .A(n4319), .B(n4320), .Z(n4295) );
  XOR U4311 ( .A(n4321), .B(n4322), .Z(n4298) );
  AND U4312 ( .A(n4323), .B(n4324), .Z(n4322) );
  XOR U4313 ( .A(n4321), .B(n4325), .Z(n4323) );
  XNOR U4314 ( .A(n4109), .B(n4303), .Z(n4305) );
  XNOR U4315 ( .A(n4326), .B(n4327), .Z(n4109) );
  AND U4316 ( .A(n58), .B(n4328), .Z(n4327) );
  XOR U4317 ( .A(n4329), .B(n4326), .Z(n4328) );
  XOR U4318 ( .A(n4330), .B(n4331), .Z(n4303) );
  AND U4319 ( .A(n4332), .B(n4333), .Z(n4331) );
  XNOR U4320 ( .A(n4330), .B(n4319), .Z(n4333) );
  IV U4321 ( .A(n4160), .Z(n4319) );
  XNOR U4322 ( .A(n4334), .B(n4312), .Z(n4160) );
  XNOR U4323 ( .A(n4335), .B(n4318), .Z(n4312) );
  XOR U4324 ( .A(n4336), .B(n4337), .Z(n4318) );
  AND U4325 ( .A(n4338), .B(n4339), .Z(n4337) );
  XOR U4326 ( .A(n4336), .B(n4340), .Z(n4338) );
  XNOR U4327 ( .A(n4317), .B(n4309), .Z(n4335) );
  XOR U4328 ( .A(n4341), .B(n4342), .Z(n4309) );
  AND U4329 ( .A(n4343), .B(n4344), .Z(n4342) );
  XNOR U4330 ( .A(n4345), .B(n4341), .Z(n4343) );
  XNOR U4331 ( .A(n4346), .B(n4314), .Z(n4317) );
  XOR U4332 ( .A(n4347), .B(n4348), .Z(n4314) );
  AND U4333 ( .A(n4349), .B(n4350), .Z(n4348) );
  XOR U4334 ( .A(n4347), .B(n4351), .Z(n4349) );
  XNOR U4335 ( .A(n4352), .B(n4353), .Z(n4346) );
  AND U4336 ( .A(n4354), .B(n4355), .Z(n4353) );
  XNOR U4337 ( .A(n4352), .B(n4356), .Z(n4354) );
  XNOR U4338 ( .A(n4313), .B(n4320), .Z(n4334) );
  AND U4339 ( .A(n4256), .B(n4357), .Z(n4320) );
  XOR U4340 ( .A(n4325), .B(n4324), .Z(n4313) );
  XNOR U4341 ( .A(n4358), .B(n4321), .Z(n4324) );
  XOR U4342 ( .A(n4359), .B(n4360), .Z(n4321) );
  AND U4343 ( .A(n4361), .B(n4362), .Z(n4360) );
  XOR U4344 ( .A(n4359), .B(n4363), .Z(n4361) );
  XNOR U4345 ( .A(n4364), .B(n4365), .Z(n4358) );
  AND U4346 ( .A(n4366), .B(n4367), .Z(n4365) );
  XOR U4347 ( .A(n4364), .B(n4368), .Z(n4366) );
  XOR U4348 ( .A(n4369), .B(n4370), .Z(n4325) );
  AND U4349 ( .A(n4371), .B(n4372), .Z(n4370) );
  XOR U4350 ( .A(n4369), .B(n4373), .Z(n4371) );
  XNOR U4351 ( .A(n4157), .B(n4330), .Z(n4332) );
  XNOR U4352 ( .A(n4374), .B(n4375), .Z(n4157) );
  AND U4353 ( .A(n58), .B(n4376), .Z(n4375) );
  XNOR U4354 ( .A(n4377), .B(n4374), .Z(n4376) );
  XOR U4355 ( .A(n4378), .B(n4379), .Z(n4330) );
  AND U4356 ( .A(n4380), .B(n4381), .Z(n4379) );
  XNOR U4357 ( .A(n4378), .B(n4256), .Z(n4381) );
  XOR U4358 ( .A(n4382), .B(n4344), .Z(n4256) );
  XNOR U4359 ( .A(n4383), .B(n4351), .Z(n4344) );
  XOR U4360 ( .A(n4340), .B(n4339), .Z(n4351) );
  XNOR U4361 ( .A(n4384), .B(n4336), .Z(n4339) );
  XOR U4362 ( .A(n4385), .B(n4386), .Z(n4336) );
  AND U4363 ( .A(n4387), .B(n4388), .Z(n4386) );
  XNOR U4364 ( .A(n4389), .B(n4390), .Z(n4387) );
  IV U4365 ( .A(n4385), .Z(n4389) );
  XNOR U4366 ( .A(n4391), .B(n4392), .Z(n4384) );
  NOR U4367 ( .A(n4393), .B(n4394), .Z(n4392) );
  XNOR U4368 ( .A(n4391), .B(n4395), .Z(n4393) );
  XOR U4369 ( .A(n4396), .B(n4397), .Z(n4340) );
  NOR U4370 ( .A(n4398), .B(n4399), .Z(n4397) );
  XNOR U4371 ( .A(n4396), .B(n4400), .Z(n4398) );
  XNOR U4372 ( .A(n4350), .B(n4341), .Z(n4383) );
  XOR U4373 ( .A(n4401), .B(n4402), .Z(n4341) );
  AND U4374 ( .A(n4403), .B(n4404), .Z(n4402) );
  XOR U4375 ( .A(n4401), .B(n4405), .Z(n4403) );
  XOR U4376 ( .A(n4406), .B(n4356), .Z(n4350) );
  XOR U4377 ( .A(n4407), .B(n4408), .Z(n4356) );
  NOR U4378 ( .A(n4409), .B(n4410), .Z(n4408) );
  XOR U4379 ( .A(n4407), .B(n4411), .Z(n4409) );
  XNOR U4380 ( .A(n4355), .B(n4347), .Z(n4406) );
  XOR U4381 ( .A(n4412), .B(n4413), .Z(n4347) );
  AND U4382 ( .A(n4414), .B(n4415), .Z(n4413) );
  XOR U4383 ( .A(n4412), .B(n4416), .Z(n4414) );
  XNOR U4384 ( .A(n4417), .B(n4352), .Z(n4355) );
  XOR U4385 ( .A(n4418), .B(n4419), .Z(n4352) );
  AND U4386 ( .A(n4420), .B(n4421), .Z(n4419) );
  XNOR U4387 ( .A(n4422), .B(n4423), .Z(n4420) );
  IV U4388 ( .A(n4418), .Z(n4422) );
  XNOR U4389 ( .A(n4424), .B(n4425), .Z(n4417) );
  NOR U4390 ( .A(n4426), .B(n4427), .Z(n4425) );
  XNOR U4391 ( .A(n4424), .B(n4428), .Z(n4426) );
  XOR U4392 ( .A(n4345), .B(n4357), .Z(n4382) );
  NOR U4393 ( .A(n4279), .B(n4429), .Z(n4357) );
  XNOR U4394 ( .A(n4363), .B(n4362), .Z(n4345) );
  XNOR U4395 ( .A(n4430), .B(n4368), .Z(n4362) );
  XNOR U4396 ( .A(n4431), .B(n4432), .Z(n4368) );
  NOR U4397 ( .A(n4433), .B(n4434), .Z(n4432) );
  XOR U4398 ( .A(n4431), .B(n4435), .Z(n4433) );
  XNOR U4399 ( .A(n4367), .B(n4359), .Z(n4430) );
  XOR U4400 ( .A(n4436), .B(n4437), .Z(n4359) );
  AND U4401 ( .A(n4438), .B(n4439), .Z(n4437) );
  XOR U4402 ( .A(n4436), .B(n4440), .Z(n4438) );
  XNOR U4403 ( .A(n4441), .B(n4364), .Z(n4367) );
  XOR U4404 ( .A(n4442), .B(n4443), .Z(n4364) );
  AND U4405 ( .A(n4444), .B(n4445), .Z(n4443) );
  XNOR U4406 ( .A(n4446), .B(n4447), .Z(n4444) );
  IV U4407 ( .A(n4442), .Z(n4446) );
  XNOR U4408 ( .A(n4448), .B(n4449), .Z(n4441) );
  NOR U4409 ( .A(n4450), .B(n4451), .Z(n4449) );
  XNOR U4410 ( .A(n4448), .B(n4452), .Z(n4450) );
  XOR U4411 ( .A(n4373), .B(n4372), .Z(n4363) );
  XNOR U4412 ( .A(n4453), .B(n4369), .Z(n4372) );
  XOR U4413 ( .A(n4454), .B(n4455), .Z(n4369) );
  AND U4414 ( .A(n4456), .B(n4457), .Z(n4455) );
  XNOR U4415 ( .A(n4458), .B(n4459), .Z(n4456) );
  IV U4416 ( .A(n4454), .Z(n4458) );
  XNOR U4417 ( .A(n4460), .B(n4461), .Z(n4453) );
  NOR U4418 ( .A(n4462), .B(n4463), .Z(n4461) );
  XNOR U4419 ( .A(n4460), .B(n4464), .Z(n4462) );
  XOR U4420 ( .A(n4465), .B(n4466), .Z(n4373) );
  NOR U4421 ( .A(n4467), .B(n4468), .Z(n4466) );
  XNOR U4422 ( .A(n4465), .B(n4469), .Z(n4467) );
  XNOR U4423 ( .A(n4253), .B(n4378), .Z(n4380) );
  XNOR U4424 ( .A(n4470), .B(n4471), .Z(n4253) );
  AND U4425 ( .A(n58), .B(n4472), .Z(n4471) );
  XOR U4426 ( .A(n4473), .B(n4470), .Z(n4472) );
  AND U4427 ( .A(n4276), .B(n4279), .Z(n4378) );
  XOR U4428 ( .A(n4474), .B(n4429), .Z(n4279) );
  XNOR U4429 ( .A(p_input[416]), .B(p_input[512]), .Z(n4429) );
  XNOR U4430 ( .A(n4405), .B(n4404), .Z(n4474) );
  XNOR U4431 ( .A(n4475), .B(n4416), .Z(n4404) );
  XOR U4432 ( .A(n4390), .B(n4388), .Z(n4416) );
  XNOR U4433 ( .A(n4476), .B(n4395), .Z(n4388) );
  XOR U4434 ( .A(p_input[440]), .B(p_input[536]), .Z(n4395) );
  XOR U4435 ( .A(n4385), .B(n4394), .Z(n4476) );
  XOR U4436 ( .A(n4477), .B(n4391), .Z(n4394) );
  XOR U4437 ( .A(p_input[438]), .B(p_input[534]), .Z(n4391) );
  XOR U4438 ( .A(p_input[439]), .B(n1634), .Z(n4477) );
  XOR U4439 ( .A(p_input[434]), .B(p_input[530]), .Z(n4385) );
  XNOR U4440 ( .A(n4400), .B(n4399), .Z(n4390) );
  XOR U4441 ( .A(n4478), .B(n4396), .Z(n4399) );
  XOR U4442 ( .A(p_input[435]), .B(p_input[531]), .Z(n4396) );
  XOR U4443 ( .A(p_input[436]), .B(n1636), .Z(n4478) );
  XOR U4444 ( .A(p_input[437]), .B(p_input[533]), .Z(n4400) );
  XOR U4445 ( .A(n4415), .B(n4479), .Z(n4475) );
  IV U4446 ( .A(n4401), .Z(n4479) );
  XOR U4447 ( .A(p_input[417]), .B(p_input[513]), .Z(n4401) );
  XNOR U4448 ( .A(n4480), .B(n4423), .Z(n4415) );
  XNOR U4449 ( .A(n4411), .B(n4410), .Z(n4423) );
  XNOR U4450 ( .A(n4481), .B(n4407), .Z(n4410) );
  XNOR U4451 ( .A(p_input[442]), .B(p_input[538]), .Z(n4407) );
  XOR U4452 ( .A(p_input[443]), .B(n1640), .Z(n4481) );
  XOR U4453 ( .A(p_input[444]), .B(p_input[540]), .Z(n4411) );
  XOR U4454 ( .A(n4421), .B(n4482), .Z(n4480) );
  IV U4455 ( .A(n4412), .Z(n4482) );
  XOR U4456 ( .A(p_input[433]), .B(p_input[529]), .Z(n4412) );
  XNOR U4457 ( .A(n4483), .B(n4428), .Z(n4421) );
  XNOR U4458 ( .A(p_input[447]), .B(n1643), .Z(n4428) );
  XOR U4459 ( .A(n4418), .B(n4427), .Z(n4483) );
  XOR U4460 ( .A(n4484), .B(n4424), .Z(n4427) );
  XOR U4461 ( .A(p_input[445]), .B(p_input[541]), .Z(n4424) );
  XOR U4462 ( .A(p_input[446]), .B(n1645), .Z(n4484) );
  XOR U4463 ( .A(p_input[441]), .B(p_input[537]), .Z(n4418) );
  XOR U4464 ( .A(n4440), .B(n4439), .Z(n4405) );
  XNOR U4465 ( .A(n4485), .B(n4447), .Z(n4439) );
  XNOR U4466 ( .A(n4435), .B(n4434), .Z(n4447) );
  XNOR U4467 ( .A(n4486), .B(n4431), .Z(n4434) );
  XNOR U4468 ( .A(p_input[427]), .B(p_input[523]), .Z(n4431) );
  XOR U4469 ( .A(p_input[428]), .B(n1648), .Z(n4486) );
  XOR U4470 ( .A(p_input[429]), .B(p_input[525]), .Z(n4435) );
  XOR U4471 ( .A(n4445), .B(n4487), .Z(n4485) );
  IV U4472 ( .A(n4436), .Z(n4487) );
  XOR U4473 ( .A(p_input[418]), .B(p_input[514]), .Z(n4436) );
  XNOR U4474 ( .A(n4488), .B(n4452), .Z(n4445) );
  XNOR U4475 ( .A(p_input[432]), .B(n1651), .Z(n4452) );
  XOR U4476 ( .A(n4442), .B(n4451), .Z(n4488) );
  XOR U4477 ( .A(n4489), .B(n4448), .Z(n4451) );
  XOR U4478 ( .A(p_input[430]), .B(p_input[526]), .Z(n4448) );
  XOR U4479 ( .A(p_input[431]), .B(n1653), .Z(n4489) );
  XOR U4480 ( .A(p_input[426]), .B(p_input[522]), .Z(n4442) );
  XOR U4481 ( .A(n4459), .B(n4457), .Z(n4440) );
  XNOR U4482 ( .A(n4490), .B(n4464), .Z(n4457) );
  XOR U4483 ( .A(p_input[425]), .B(p_input[521]), .Z(n4464) );
  XOR U4484 ( .A(n4454), .B(n4463), .Z(n4490) );
  XOR U4485 ( .A(n4491), .B(n4460), .Z(n4463) );
  XOR U4486 ( .A(p_input[423]), .B(p_input[519]), .Z(n4460) );
  XOR U4487 ( .A(p_input[424]), .B(n1877), .Z(n4491) );
  XOR U4488 ( .A(p_input[419]), .B(p_input[515]), .Z(n4454) );
  XNOR U4489 ( .A(n4469), .B(n4468), .Z(n4459) );
  XOR U4490 ( .A(n4492), .B(n4465), .Z(n4468) );
  XOR U4491 ( .A(p_input[420]), .B(p_input[516]), .Z(n4465) );
  XOR U4492 ( .A(p_input[421]), .B(n1879), .Z(n4492) );
  XOR U4493 ( .A(p_input[422]), .B(p_input[518]), .Z(n4469) );
  XOR U4494 ( .A(n4493), .B(n4494), .Z(n4276) );
  AND U4495 ( .A(n58), .B(n4495), .Z(n4494) );
  XNOR U4496 ( .A(n4496), .B(n4493), .Z(n4495) );
  XNOR U4497 ( .A(n4497), .B(n4498), .Z(n58) );
  NOR U4498 ( .A(n4499), .B(n4500), .Z(n4498) );
  XOR U4499 ( .A(n4285), .B(n4497), .Z(n4500) );
  AND U4500 ( .A(n4299), .B(n4501), .Z(n4285) );
  NOR U4501 ( .A(n4497), .B(n4284), .Z(n4499) );
  AND U4502 ( .A(n4502), .B(n4503), .Z(n4284) );
  XOR U4503 ( .A(n4504), .B(n4505), .Z(n4497) );
  AND U4504 ( .A(n4506), .B(n4507), .Z(n4505) );
  XNOR U4505 ( .A(n4504), .B(n4502), .Z(n4507) );
  IV U4506 ( .A(n4302), .Z(n4502) );
  XOR U4507 ( .A(n4508), .B(n4509), .Z(n4302) );
  XOR U4508 ( .A(n4510), .B(n4503), .Z(n4509) );
  AND U4509 ( .A(n4329), .B(n4511), .Z(n4503) );
  AND U4510 ( .A(n4512), .B(n4513), .Z(n4510) );
  XOR U4511 ( .A(n4514), .B(n4508), .Z(n4512) );
  XNOR U4512 ( .A(n4515), .B(n4504), .Z(n4506) );
  IV U4513 ( .A(n4299), .Z(n4515) );
  XNOR U4514 ( .A(n4516), .B(n4517), .Z(n4299) );
  XOR U4515 ( .A(n4518), .B(n4501), .Z(n4517) );
  AND U4516 ( .A(n4326), .B(n4519), .Z(n4501) );
  AND U4517 ( .A(n4520), .B(n4521), .Z(n4518) );
  XNOR U4518 ( .A(n4516), .B(n4522), .Z(n4520) );
  XOR U4519 ( .A(n4523), .B(n4524), .Z(n4504) );
  AND U4520 ( .A(n4525), .B(n4526), .Z(n4524) );
  XNOR U4521 ( .A(n4523), .B(n4329), .Z(n4526) );
  XOR U4522 ( .A(n4527), .B(n4513), .Z(n4329) );
  XNOR U4523 ( .A(n4528), .B(n4508), .Z(n4513) );
  XOR U4524 ( .A(n4529), .B(n4530), .Z(n4508) );
  AND U4525 ( .A(n4531), .B(n4532), .Z(n4530) );
  XOR U4526 ( .A(n4533), .B(n4529), .Z(n4531) );
  XNOR U4527 ( .A(n4534), .B(n4535), .Z(n4528) );
  AND U4528 ( .A(n4536), .B(n4537), .Z(n4535) );
  XOR U4529 ( .A(n4534), .B(n4538), .Z(n4536) );
  XNOR U4530 ( .A(n4514), .B(n4511), .Z(n4527) );
  AND U4531 ( .A(n4539), .B(n4540), .Z(n4511) );
  XOR U4532 ( .A(n4541), .B(n4542), .Z(n4514) );
  AND U4533 ( .A(n4543), .B(n4544), .Z(n4542) );
  XOR U4534 ( .A(n4541), .B(n4545), .Z(n4543) );
  XOR U4535 ( .A(n4326), .B(n4523), .Z(n4525) );
  XNOR U4536 ( .A(n4546), .B(n4522), .Z(n4326) );
  XNOR U4537 ( .A(n4547), .B(n4548), .Z(n4522) );
  AND U4538 ( .A(n4549), .B(n4550), .Z(n4548) );
  XOR U4539 ( .A(n4547), .B(n4551), .Z(n4549) );
  XNOR U4540 ( .A(n4521), .B(n4519), .Z(n4546) );
  AND U4541 ( .A(n4374), .B(n4552), .Z(n4519) );
  XNOR U4542 ( .A(n4553), .B(n4516), .Z(n4521) );
  XOR U4543 ( .A(n4554), .B(n4555), .Z(n4516) );
  AND U4544 ( .A(n4556), .B(n4557), .Z(n4555) );
  XOR U4545 ( .A(n4554), .B(n4558), .Z(n4556) );
  XNOR U4546 ( .A(n4559), .B(n4560), .Z(n4553) );
  AND U4547 ( .A(n4561), .B(n4562), .Z(n4560) );
  XNOR U4548 ( .A(n4559), .B(n4563), .Z(n4561) );
  XOR U4549 ( .A(n4564), .B(n4565), .Z(n4523) );
  AND U4550 ( .A(n4566), .B(n4567), .Z(n4565) );
  XNOR U4551 ( .A(n4564), .B(n4539), .Z(n4567) );
  IV U4552 ( .A(n4377), .Z(n4539) );
  XNOR U4553 ( .A(n4568), .B(n4532), .Z(n4377) );
  XNOR U4554 ( .A(n4569), .B(n4538), .Z(n4532) );
  XOR U4555 ( .A(n4570), .B(n4571), .Z(n4538) );
  AND U4556 ( .A(n4572), .B(n4573), .Z(n4571) );
  XOR U4557 ( .A(n4570), .B(n4574), .Z(n4572) );
  XNOR U4558 ( .A(n4537), .B(n4529), .Z(n4569) );
  XOR U4559 ( .A(n4575), .B(n4576), .Z(n4529) );
  AND U4560 ( .A(n4577), .B(n4578), .Z(n4576) );
  XNOR U4561 ( .A(n4579), .B(n4575), .Z(n4577) );
  XNOR U4562 ( .A(n4580), .B(n4534), .Z(n4537) );
  XOR U4563 ( .A(n4581), .B(n4582), .Z(n4534) );
  AND U4564 ( .A(n4583), .B(n4584), .Z(n4582) );
  XOR U4565 ( .A(n4581), .B(n4585), .Z(n4583) );
  XNOR U4566 ( .A(n4586), .B(n4587), .Z(n4580) );
  AND U4567 ( .A(n4588), .B(n4589), .Z(n4587) );
  XNOR U4568 ( .A(n4586), .B(n4590), .Z(n4588) );
  XNOR U4569 ( .A(n4533), .B(n4540), .Z(n4568) );
  AND U4570 ( .A(n4473), .B(n4591), .Z(n4540) );
  XOR U4571 ( .A(n4545), .B(n4544), .Z(n4533) );
  XNOR U4572 ( .A(n4592), .B(n4541), .Z(n4544) );
  XOR U4573 ( .A(n4593), .B(n4594), .Z(n4541) );
  AND U4574 ( .A(n4595), .B(n4596), .Z(n4594) );
  XOR U4575 ( .A(n4593), .B(n4597), .Z(n4595) );
  XNOR U4576 ( .A(n4598), .B(n4599), .Z(n4592) );
  AND U4577 ( .A(n4600), .B(n4601), .Z(n4599) );
  XOR U4578 ( .A(n4598), .B(n4602), .Z(n4600) );
  XOR U4579 ( .A(n4603), .B(n4604), .Z(n4545) );
  AND U4580 ( .A(n4605), .B(n4606), .Z(n4604) );
  XOR U4581 ( .A(n4603), .B(n4607), .Z(n4605) );
  XNOR U4582 ( .A(n4608), .B(n4564), .Z(n4566) );
  IV U4583 ( .A(n4374), .Z(n4608) );
  XOR U4584 ( .A(n4609), .B(n4558), .Z(n4374) );
  XOR U4585 ( .A(n4551), .B(n4550), .Z(n4558) );
  XNOR U4586 ( .A(n4610), .B(n4547), .Z(n4550) );
  XOR U4587 ( .A(n4611), .B(n4612), .Z(n4547) );
  AND U4588 ( .A(n4613), .B(n4614), .Z(n4612) );
  XOR U4589 ( .A(n4611), .B(n4615), .Z(n4613) );
  XNOR U4590 ( .A(n4616), .B(n4617), .Z(n4610) );
  AND U4591 ( .A(n4618), .B(n4619), .Z(n4617) );
  XOR U4592 ( .A(n4616), .B(n4620), .Z(n4618) );
  XOR U4593 ( .A(n4621), .B(n4622), .Z(n4551) );
  AND U4594 ( .A(n4623), .B(n4624), .Z(n4622) );
  XOR U4595 ( .A(n4621), .B(n4625), .Z(n4623) );
  XNOR U4596 ( .A(n4557), .B(n4552), .Z(n4609) );
  AND U4597 ( .A(n4470), .B(n4626), .Z(n4552) );
  XOR U4598 ( .A(n4627), .B(n4563), .Z(n4557) );
  XNOR U4599 ( .A(n4628), .B(n4629), .Z(n4563) );
  AND U4600 ( .A(n4630), .B(n4631), .Z(n4629) );
  XOR U4601 ( .A(n4628), .B(n4632), .Z(n4630) );
  XNOR U4602 ( .A(n4562), .B(n4554), .Z(n4627) );
  XOR U4603 ( .A(n4633), .B(n4634), .Z(n4554) );
  AND U4604 ( .A(n4635), .B(n4636), .Z(n4634) );
  XOR U4605 ( .A(n4633), .B(n4637), .Z(n4635) );
  XNOR U4606 ( .A(n4638), .B(n4559), .Z(n4562) );
  XOR U4607 ( .A(n4639), .B(n4640), .Z(n4559) );
  AND U4608 ( .A(n4641), .B(n4642), .Z(n4640) );
  XOR U4609 ( .A(n4639), .B(n4643), .Z(n4641) );
  XNOR U4610 ( .A(n4644), .B(n4645), .Z(n4638) );
  AND U4611 ( .A(n4646), .B(n4647), .Z(n4645) );
  XNOR U4612 ( .A(n4644), .B(n4648), .Z(n4646) );
  XOR U4613 ( .A(n4649), .B(n4650), .Z(n4564) );
  AND U4614 ( .A(n4651), .B(n4652), .Z(n4650) );
  XNOR U4615 ( .A(n4649), .B(n4473), .Z(n4652) );
  XOR U4616 ( .A(n4653), .B(n4578), .Z(n4473) );
  XNOR U4617 ( .A(n4654), .B(n4585), .Z(n4578) );
  XOR U4618 ( .A(n4574), .B(n4573), .Z(n4585) );
  XNOR U4619 ( .A(n4655), .B(n4570), .Z(n4573) );
  XOR U4620 ( .A(n4656), .B(n4657), .Z(n4570) );
  AND U4621 ( .A(n4658), .B(n4659), .Z(n4657) );
  XNOR U4622 ( .A(n4660), .B(n4661), .Z(n4658) );
  IV U4623 ( .A(n4656), .Z(n4660) );
  XNOR U4624 ( .A(n4662), .B(n4663), .Z(n4655) );
  NOR U4625 ( .A(n4664), .B(n4665), .Z(n4663) );
  XNOR U4626 ( .A(n4662), .B(n4666), .Z(n4664) );
  XOR U4627 ( .A(n4667), .B(n4668), .Z(n4574) );
  NOR U4628 ( .A(n4669), .B(n4670), .Z(n4668) );
  XNOR U4629 ( .A(n4667), .B(n4671), .Z(n4669) );
  XNOR U4630 ( .A(n4584), .B(n4575), .Z(n4654) );
  XOR U4631 ( .A(n4672), .B(n4673), .Z(n4575) );
  AND U4632 ( .A(n4674), .B(n4675), .Z(n4673) );
  XOR U4633 ( .A(n4672), .B(n4676), .Z(n4674) );
  XOR U4634 ( .A(n4677), .B(n4590), .Z(n4584) );
  XOR U4635 ( .A(n4678), .B(n4679), .Z(n4590) );
  NOR U4636 ( .A(n4680), .B(n4681), .Z(n4679) );
  XOR U4637 ( .A(n4678), .B(n4682), .Z(n4680) );
  XNOR U4638 ( .A(n4589), .B(n4581), .Z(n4677) );
  XOR U4639 ( .A(n4683), .B(n4684), .Z(n4581) );
  AND U4640 ( .A(n4685), .B(n4686), .Z(n4684) );
  XOR U4641 ( .A(n4683), .B(n4687), .Z(n4685) );
  XNOR U4642 ( .A(n4688), .B(n4586), .Z(n4589) );
  XOR U4643 ( .A(n4689), .B(n4690), .Z(n4586) );
  AND U4644 ( .A(n4691), .B(n4692), .Z(n4690) );
  XNOR U4645 ( .A(n4693), .B(n4694), .Z(n4691) );
  IV U4646 ( .A(n4689), .Z(n4693) );
  XNOR U4647 ( .A(n4695), .B(n4696), .Z(n4688) );
  NOR U4648 ( .A(n4697), .B(n4698), .Z(n4696) );
  XNOR U4649 ( .A(n4695), .B(n4699), .Z(n4697) );
  XOR U4650 ( .A(n4579), .B(n4591), .Z(n4653) );
  NOR U4651 ( .A(n4496), .B(n4700), .Z(n4591) );
  XNOR U4652 ( .A(n4597), .B(n4596), .Z(n4579) );
  XNOR U4653 ( .A(n4701), .B(n4602), .Z(n4596) );
  XNOR U4654 ( .A(n4702), .B(n4703), .Z(n4602) );
  NOR U4655 ( .A(n4704), .B(n4705), .Z(n4703) );
  XOR U4656 ( .A(n4702), .B(n4706), .Z(n4704) );
  XNOR U4657 ( .A(n4601), .B(n4593), .Z(n4701) );
  XOR U4658 ( .A(n4707), .B(n4708), .Z(n4593) );
  AND U4659 ( .A(n4709), .B(n4710), .Z(n4708) );
  XOR U4660 ( .A(n4707), .B(n4711), .Z(n4709) );
  XNOR U4661 ( .A(n4712), .B(n4598), .Z(n4601) );
  XOR U4662 ( .A(n4713), .B(n4714), .Z(n4598) );
  AND U4663 ( .A(n4715), .B(n4716), .Z(n4714) );
  XNOR U4664 ( .A(n4717), .B(n4718), .Z(n4715) );
  IV U4665 ( .A(n4713), .Z(n4717) );
  XNOR U4666 ( .A(n4719), .B(n4720), .Z(n4712) );
  NOR U4667 ( .A(n4721), .B(n4722), .Z(n4720) );
  XNOR U4668 ( .A(n4719), .B(n4723), .Z(n4721) );
  XOR U4669 ( .A(n4607), .B(n4606), .Z(n4597) );
  XNOR U4670 ( .A(n4724), .B(n4603), .Z(n4606) );
  XOR U4671 ( .A(n4725), .B(n4726), .Z(n4603) );
  AND U4672 ( .A(n4727), .B(n4728), .Z(n4726) );
  XNOR U4673 ( .A(n4729), .B(n4730), .Z(n4727) );
  IV U4674 ( .A(n4725), .Z(n4729) );
  XNOR U4675 ( .A(n4731), .B(n4732), .Z(n4724) );
  NOR U4676 ( .A(n4733), .B(n4734), .Z(n4732) );
  XNOR U4677 ( .A(n4731), .B(n4735), .Z(n4733) );
  XOR U4678 ( .A(n4736), .B(n4737), .Z(n4607) );
  NOR U4679 ( .A(n4738), .B(n4739), .Z(n4737) );
  XNOR U4680 ( .A(n4736), .B(n4740), .Z(n4738) );
  XNOR U4681 ( .A(n4741), .B(n4649), .Z(n4651) );
  IV U4682 ( .A(n4470), .Z(n4741) );
  XOR U4683 ( .A(n4742), .B(n4637), .Z(n4470) );
  XOR U4684 ( .A(n4615), .B(n4614), .Z(n4637) );
  XNOR U4685 ( .A(n4743), .B(n4620), .Z(n4614) );
  XOR U4686 ( .A(n4744), .B(n4745), .Z(n4620) );
  NOR U4687 ( .A(n4746), .B(n4747), .Z(n4745) );
  XNOR U4688 ( .A(n4744), .B(n4748), .Z(n4746) );
  XNOR U4689 ( .A(n4619), .B(n4611), .Z(n4743) );
  XOR U4690 ( .A(n4749), .B(n4750), .Z(n4611) );
  AND U4691 ( .A(n4751), .B(n4752), .Z(n4750) );
  XNOR U4692 ( .A(n4749), .B(n4753), .Z(n4751) );
  XNOR U4693 ( .A(n4754), .B(n4616), .Z(n4619) );
  XOR U4694 ( .A(n4755), .B(n4756), .Z(n4616) );
  AND U4695 ( .A(n4757), .B(n4758), .Z(n4756) );
  XOR U4696 ( .A(n4755), .B(n4759), .Z(n4757) );
  XNOR U4697 ( .A(n4760), .B(n4761), .Z(n4754) );
  NOR U4698 ( .A(n4762), .B(n4763), .Z(n4761) );
  XOR U4699 ( .A(n4760), .B(n4764), .Z(n4762) );
  XOR U4700 ( .A(n4625), .B(n4624), .Z(n4615) );
  XNOR U4701 ( .A(n4765), .B(n4621), .Z(n4624) );
  XOR U4702 ( .A(n4766), .B(n4767), .Z(n4621) );
  AND U4703 ( .A(n4768), .B(n4769), .Z(n4767) );
  XOR U4704 ( .A(n4766), .B(n4770), .Z(n4768) );
  XNOR U4705 ( .A(n4771), .B(n4772), .Z(n4765) );
  NOR U4706 ( .A(n4773), .B(n4774), .Z(n4772) );
  XNOR U4707 ( .A(n4771), .B(n4775), .Z(n4773) );
  XOR U4708 ( .A(n4776), .B(n4777), .Z(n4625) );
  NOR U4709 ( .A(n4778), .B(n4779), .Z(n4777) );
  XNOR U4710 ( .A(n4776), .B(n4780), .Z(n4778) );
  XNOR U4711 ( .A(n4636), .B(n4626), .Z(n4742) );
  AND U4712 ( .A(n4493), .B(n4781), .Z(n4626) );
  XNOR U4713 ( .A(n4782), .B(n4643), .Z(n4636) );
  XOR U4714 ( .A(n4632), .B(n4631), .Z(n4643) );
  XNOR U4715 ( .A(n4783), .B(n4628), .Z(n4631) );
  XOR U4716 ( .A(n4784), .B(n4785), .Z(n4628) );
  AND U4717 ( .A(n4786), .B(n4787), .Z(n4785) );
  XOR U4718 ( .A(n4784), .B(n4788), .Z(n4786) );
  XNOR U4719 ( .A(n4789), .B(n4790), .Z(n4783) );
  NOR U4720 ( .A(n4791), .B(n4792), .Z(n4790) );
  XNOR U4721 ( .A(n4789), .B(n4793), .Z(n4791) );
  XOR U4722 ( .A(n4794), .B(n4795), .Z(n4632) );
  NOR U4723 ( .A(n4796), .B(n4797), .Z(n4795) );
  XNOR U4724 ( .A(n4794), .B(n4798), .Z(n4796) );
  XNOR U4725 ( .A(n4642), .B(n4633), .Z(n4782) );
  XOR U4726 ( .A(n4799), .B(n4800), .Z(n4633) );
  NOR U4727 ( .A(n4801), .B(n4802), .Z(n4800) );
  XNOR U4728 ( .A(n4799), .B(n4803), .Z(n4801) );
  XOR U4729 ( .A(n4804), .B(n4648), .Z(n4642) );
  XNOR U4730 ( .A(n4805), .B(n4806), .Z(n4648) );
  NOR U4731 ( .A(n4807), .B(n4808), .Z(n4806) );
  XNOR U4732 ( .A(n4805), .B(n4809), .Z(n4807) );
  XNOR U4733 ( .A(n4647), .B(n4639), .Z(n4804) );
  XOR U4734 ( .A(n4810), .B(n4811), .Z(n4639) );
  AND U4735 ( .A(n4812), .B(n4813), .Z(n4811) );
  XOR U4736 ( .A(n4810), .B(n4814), .Z(n4812) );
  XNOR U4737 ( .A(n4815), .B(n4644), .Z(n4647) );
  XOR U4738 ( .A(n4816), .B(n4817), .Z(n4644) );
  AND U4739 ( .A(n4818), .B(n4819), .Z(n4817) );
  XOR U4740 ( .A(n4816), .B(n4820), .Z(n4818) );
  XNOR U4741 ( .A(n4821), .B(n4822), .Z(n4815) );
  NOR U4742 ( .A(n4823), .B(n4824), .Z(n4822) );
  XOR U4743 ( .A(n4821), .B(n4825), .Z(n4823) );
  AND U4744 ( .A(n4493), .B(n4496), .Z(n4649) );
  XOR U4745 ( .A(n4826), .B(n4700), .Z(n4496) );
  XNOR U4746 ( .A(p_input[448]), .B(p_input[512]), .Z(n4700) );
  XNOR U4747 ( .A(n4676), .B(n4675), .Z(n4826) );
  XNOR U4748 ( .A(n4827), .B(n4687), .Z(n4675) );
  XOR U4749 ( .A(n4661), .B(n4659), .Z(n4687) );
  XNOR U4750 ( .A(n4828), .B(n4666), .Z(n4659) );
  XOR U4751 ( .A(p_input[472]), .B(p_input[536]), .Z(n4666) );
  XOR U4752 ( .A(n4656), .B(n4665), .Z(n4828) );
  XOR U4753 ( .A(n4829), .B(n4662), .Z(n4665) );
  XOR U4754 ( .A(p_input[470]), .B(p_input[534]), .Z(n4662) );
  XOR U4755 ( .A(p_input[471]), .B(n1634), .Z(n4829) );
  XOR U4756 ( .A(p_input[466]), .B(p_input[530]), .Z(n4656) );
  XNOR U4757 ( .A(n4671), .B(n4670), .Z(n4661) );
  XOR U4758 ( .A(n4830), .B(n4667), .Z(n4670) );
  XOR U4759 ( .A(p_input[467]), .B(p_input[531]), .Z(n4667) );
  XOR U4760 ( .A(p_input[468]), .B(n1636), .Z(n4830) );
  XOR U4761 ( .A(p_input[469]), .B(p_input[533]), .Z(n4671) );
  XOR U4762 ( .A(n4686), .B(n4831), .Z(n4827) );
  IV U4763 ( .A(n4672), .Z(n4831) );
  XOR U4764 ( .A(p_input[449]), .B(p_input[513]), .Z(n4672) );
  XNOR U4765 ( .A(n4832), .B(n4694), .Z(n4686) );
  XNOR U4766 ( .A(n4682), .B(n4681), .Z(n4694) );
  XNOR U4767 ( .A(n4833), .B(n4678), .Z(n4681) );
  XNOR U4768 ( .A(p_input[474]), .B(p_input[538]), .Z(n4678) );
  XOR U4769 ( .A(p_input[475]), .B(n1640), .Z(n4833) );
  XOR U4770 ( .A(p_input[476]), .B(p_input[540]), .Z(n4682) );
  XOR U4771 ( .A(n4692), .B(n4834), .Z(n4832) );
  IV U4772 ( .A(n4683), .Z(n4834) );
  XOR U4773 ( .A(p_input[465]), .B(p_input[529]), .Z(n4683) );
  XNOR U4774 ( .A(n4835), .B(n4699), .Z(n4692) );
  XNOR U4775 ( .A(p_input[479]), .B(n1643), .Z(n4699) );
  IV U4776 ( .A(p_input[543]), .Z(n1643) );
  XOR U4777 ( .A(n4689), .B(n4698), .Z(n4835) );
  XOR U4778 ( .A(n4836), .B(n4695), .Z(n4698) );
  XOR U4779 ( .A(p_input[477]), .B(p_input[541]), .Z(n4695) );
  XOR U4780 ( .A(p_input[478]), .B(n1645), .Z(n4836) );
  XOR U4781 ( .A(p_input[473]), .B(p_input[537]), .Z(n4689) );
  XOR U4782 ( .A(n4711), .B(n4710), .Z(n4676) );
  XNOR U4783 ( .A(n4837), .B(n4718), .Z(n4710) );
  XNOR U4784 ( .A(n4706), .B(n4705), .Z(n4718) );
  XNOR U4785 ( .A(n4838), .B(n4702), .Z(n4705) );
  XNOR U4786 ( .A(p_input[459]), .B(p_input[523]), .Z(n4702) );
  XOR U4787 ( .A(p_input[460]), .B(n1648), .Z(n4838) );
  XOR U4788 ( .A(p_input[461]), .B(p_input[525]), .Z(n4706) );
  XOR U4789 ( .A(n4716), .B(n4839), .Z(n4837) );
  IV U4790 ( .A(n4707), .Z(n4839) );
  XOR U4791 ( .A(p_input[450]), .B(p_input[514]), .Z(n4707) );
  XNOR U4792 ( .A(n4840), .B(n4723), .Z(n4716) );
  XNOR U4793 ( .A(p_input[464]), .B(n1651), .Z(n4723) );
  IV U4794 ( .A(p_input[528]), .Z(n1651) );
  XOR U4795 ( .A(n4713), .B(n4722), .Z(n4840) );
  XOR U4796 ( .A(n4841), .B(n4719), .Z(n4722) );
  XOR U4797 ( .A(p_input[462]), .B(p_input[526]), .Z(n4719) );
  XOR U4798 ( .A(p_input[463]), .B(n1653), .Z(n4841) );
  XOR U4799 ( .A(p_input[458]), .B(p_input[522]), .Z(n4713) );
  XOR U4800 ( .A(n4730), .B(n4728), .Z(n4711) );
  XNOR U4801 ( .A(n4842), .B(n4735), .Z(n4728) );
  XOR U4802 ( .A(p_input[457]), .B(p_input[521]), .Z(n4735) );
  XOR U4803 ( .A(n4725), .B(n4734), .Z(n4842) );
  XOR U4804 ( .A(n4843), .B(n4731), .Z(n4734) );
  XOR U4805 ( .A(p_input[455]), .B(p_input[519]), .Z(n4731) );
  XOR U4806 ( .A(p_input[456]), .B(n1877), .Z(n4843) );
  XOR U4807 ( .A(p_input[451]), .B(p_input[515]), .Z(n4725) );
  XNOR U4808 ( .A(n4740), .B(n4739), .Z(n4730) );
  XOR U4809 ( .A(n4844), .B(n4736), .Z(n4739) );
  XOR U4810 ( .A(p_input[452]), .B(p_input[516]), .Z(n4736) );
  XOR U4811 ( .A(p_input[453]), .B(n1879), .Z(n4844) );
  XOR U4812 ( .A(p_input[454]), .B(p_input[518]), .Z(n4740) );
  XOR U4813 ( .A(n4845), .B(n4803), .Z(n4493) );
  XNOR U4814 ( .A(n4753), .B(n4752), .Z(n4803) );
  XNOR U4815 ( .A(n4846), .B(n4759), .Z(n4752) );
  XNOR U4816 ( .A(n4748), .B(n4747), .Z(n4759) );
  XOR U4817 ( .A(n4847), .B(n4744), .Z(n4747) );
  XNOR U4818 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n2090), .Z(n4744) );
  IV U4819 ( .A(p_input[523]), .Z(n2090) );
  XOR U4820 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n1648), .Z(n4847) );
  IV U4821 ( .A(p_input[524]), .Z(n1648) );
  XOR U4822 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[525]), .Z(n4748)
         );
  XNOR U4823 ( .A(n4758), .B(n4749), .Z(n4846) );
  XNOR U4824 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n2091), .Z(n4749) );
  IV U4825 ( .A(p_input[514]), .Z(n2091) );
  XOR U4826 ( .A(n4848), .B(n4764), .Z(n4758) );
  XNOR U4827 ( .A(\knn_comb_/min_val_out[0][16] ), .B(p_input[528]), .Z(n4764)
         );
  XOR U4828 ( .A(n4755), .B(n4763), .Z(n4848) );
  XOR U4829 ( .A(n4849), .B(n4760), .Z(n4763) );
  XOR U4830 ( .A(\knn_comb_/min_val_out[0][14] ), .B(p_input[526]), .Z(n4760)
         );
  XOR U4831 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n1653), .Z(n4849) );
  IV U4832 ( .A(p_input[527]), .Z(n1653) );
  XNOR U4833 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n2094), .Z(n4755) );
  IV U4834 ( .A(p_input[522]), .Z(n2094) );
  XNOR U4835 ( .A(n4770), .B(n4769), .Z(n4753) );
  XNOR U4836 ( .A(n4850), .B(n4775), .Z(n4769) );
  XOR U4837 ( .A(\knn_comb_/min_val_out[0][9] ), .B(p_input[521]), .Z(n4775)
         );
  XOR U4838 ( .A(n4766), .B(n4774), .Z(n4850) );
  XOR U4839 ( .A(n4851), .B(n4771), .Z(n4774) );
  XOR U4840 ( .A(\knn_comb_/min_val_out[0][7] ), .B(p_input[519]), .Z(n4771)
         );
  XOR U4841 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n1877), .Z(n4851) );
  IV U4842 ( .A(p_input[520]), .Z(n1877) );
  XNOR U4843 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n2097), .Z(n4766) );
  IV U4844 ( .A(p_input[515]), .Z(n2097) );
  XNOR U4845 ( .A(n4780), .B(n4779), .Z(n4770) );
  XOR U4846 ( .A(n4852), .B(n4776), .Z(n4779) );
  XOR U4847 ( .A(\knn_comb_/min_val_out[0][4] ), .B(p_input[516]), .Z(n4776)
         );
  XOR U4848 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n1879), .Z(n4852) );
  IV U4849 ( .A(p_input[517]), .Z(n1879) );
  XOR U4850 ( .A(\knn_comb_/min_val_out[0][6] ), .B(p_input[518]), .Z(n4780)
         );
  XOR U4851 ( .A(n4802), .B(n4781), .Z(n4845) );
  XOR U4852 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[512]), .Z(n4781)
         );
  XOR U4853 ( .A(n4853), .B(n4814), .Z(n4802) );
  XOR U4854 ( .A(n4788), .B(n4787), .Z(n4814) );
  XNOR U4855 ( .A(n4854), .B(n4793), .Z(n4787) );
  XOR U4856 ( .A(\knn_comb_/min_val_out[0][24] ), .B(p_input[536]), .Z(n4793)
         );
  XOR U4857 ( .A(n4784), .B(n4792), .Z(n4854) );
  XOR U4858 ( .A(n4855), .B(n4789), .Z(n4792) );
  XOR U4859 ( .A(\knn_comb_/min_val_out[0][22] ), .B(p_input[534]), .Z(n4789)
         );
  XOR U4860 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n1634), .Z(n4855) );
  IV U4861 ( .A(p_input[535]), .Z(n1634) );
  XNOR U4862 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n2080), .Z(n4784) );
  IV U4863 ( .A(p_input[530]), .Z(n2080) );
  XNOR U4864 ( .A(n4798), .B(n4797), .Z(n4788) );
  XOR U4865 ( .A(n4856), .B(n4794), .Z(n4797) );
  XOR U4866 ( .A(\knn_comb_/min_val_out[0][19] ), .B(p_input[531]), .Z(n4794)
         );
  XOR U4867 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n1636), .Z(n4856) );
  IV U4868 ( .A(p_input[532]), .Z(n1636) );
  XOR U4869 ( .A(\knn_comb_/min_val_out[0][21] ), .B(p_input[533]), .Z(n4798)
         );
  XNOR U4870 ( .A(n4813), .B(n4799), .Z(n4853) );
  XNOR U4871 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n2082), .Z(n4799) );
  IV U4872 ( .A(p_input[513]), .Z(n2082) );
  XNOR U4873 ( .A(n4857), .B(n4820), .Z(n4813) );
  XNOR U4874 ( .A(n4809), .B(n4808), .Z(n4820) );
  XOR U4875 ( .A(n4858), .B(n4805), .Z(n4808) );
  XNOR U4876 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n1865), .Z(n4805) );
  IV U4877 ( .A(p_input[538]), .Z(n1865) );
  XOR U4878 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n1640), .Z(n4858) );
  IV U4879 ( .A(p_input[539]), .Z(n1640) );
  XOR U4880 ( .A(\knn_comb_/min_val_out[0][28] ), .B(p_input[540]), .Z(n4809)
         );
  XNOR U4881 ( .A(n4819), .B(n4810), .Z(n4857) );
  XNOR U4882 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n2085), .Z(n4810) );
  IV U4883 ( .A(p_input[529]), .Z(n2085) );
  XOR U4884 ( .A(n4859), .B(n4825), .Z(n4819) );
  XNOR U4885 ( .A(\knn_comb_/min_val_out[0][31] ), .B(p_input[543]), .Z(n4825)
         );
  XOR U4886 ( .A(n4816), .B(n4824), .Z(n4859) );
  XOR U4887 ( .A(n4860), .B(n4821), .Z(n4824) );
  XOR U4888 ( .A(\knn_comb_/min_val_out[0][29] ), .B(p_input[541]), .Z(n4821)
         );
  XOR U4889 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n1645), .Z(n4860) );
  IV U4890 ( .A(p_input[542]), .Z(n1645) );
  XNOR U4891 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n1869), .Z(n4816) );
  IV U4892 ( .A(p_input[537]), .Z(n1869) );
endmodule

