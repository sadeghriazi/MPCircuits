
module psi_BMR_b100_n10 ( p_input, o );
  input [999:0] p_input;
  output [99:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800;

  AND U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(n3), .B(n4), .Z(n2) );
  AND U3 ( .A(n5), .B(p_input[309]), .Z(n4) );
  AND U4 ( .A(p_input[209]), .B(p_input[109]), .Z(n5) );
  AND U5 ( .A(p_input[509]), .B(p_input[409]), .Z(n3) );
  AND U6 ( .A(n6), .B(n7), .Z(n1) );
  AND U7 ( .A(n8), .B(p_input[809]), .Z(n7) );
  AND U8 ( .A(p_input[709]), .B(p_input[609]), .Z(n8) );
  AND U9 ( .A(p_input[9]), .B(p_input[909]), .Z(n6) );
  AND U10 ( .A(n9), .B(n10), .Z(o[99]) );
  AND U11 ( .A(n11), .B(n12), .Z(n10) );
  AND U12 ( .A(n13), .B(p_input[399]), .Z(n12) );
  AND U13 ( .A(p_input[299]), .B(p_input[199]), .Z(n13) );
  AND U14 ( .A(p_input[599]), .B(p_input[499]), .Z(n11) );
  AND U15 ( .A(n14), .B(n15), .Z(n9) );
  AND U16 ( .A(n16), .B(p_input[899]), .Z(n15) );
  AND U17 ( .A(p_input[799]), .B(p_input[699]), .Z(n16) );
  AND U18 ( .A(p_input[99]), .B(p_input[999]), .Z(n14) );
  AND U19 ( .A(n17), .B(n18), .Z(o[98]) );
  AND U20 ( .A(n19), .B(n20), .Z(n18) );
  AND U21 ( .A(n21), .B(p_input[398]), .Z(n20) );
  AND U22 ( .A(p_input[298]), .B(p_input[198]), .Z(n21) );
  AND U23 ( .A(p_input[598]), .B(p_input[498]), .Z(n19) );
  AND U24 ( .A(n22), .B(n23), .Z(n17) );
  AND U25 ( .A(n24), .B(p_input[898]), .Z(n23) );
  AND U26 ( .A(p_input[798]), .B(p_input[698]), .Z(n24) );
  AND U27 ( .A(p_input[998]), .B(p_input[98]), .Z(n22) );
  AND U28 ( .A(n25), .B(n26), .Z(o[97]) );
  AND U29 ( .A(n27), .B(n28), .Z(n26) );
  AND U30 ( .A(n29), .B(p_input[397]), .Z(n28) );
  AND U31 ( .A(p_input[297]), .B(p_input[197]), .Z(n29) );
  AND U32 ( .A(p_input[597]), .B(p_input[497]), .Z(n27) );
  AND U33 ( .A(n30), .B(n31), .Z(n25) );
  AND U34 ( .A(n32), .B(p_input[897]), .Z(n31) );
  AND U35 ( .A(p_input[797]), .B(p_input[697]), .Z(n32) );
  AND U36 ( .A(p_input[997]), .B(p_input[97]), .Z(n30) );
  AND U37 ( .A(n33), .B(n34), .Z(o[96]) );
  AND U38 ( .A(n35), .B(n36), .Z(n34) );
  AND U39 ( .A(n37), .B(p_input[396]), .Z(n36) );
  AND U40 ( .A(p_input[296]), .B(p_input[196]), .Z(n37) );
  AND U41 ( .A(p_input[596]), .B(p_input[496]), .Z(n35) );
  AND U42 ( .A(n38), .B(n39), .Z(n33) );
  AND U43 ( .A(n40), .B(p_input[896]), .Z(n39) );
  AND U44 ( .A(p_input[796]), .B(p_input[696]), .Z(n40) );
  AND U45 ( .A(p_input[996]), .B(p_input[96]), .Z(n38) );
  AND U46 ( .A(n41), .B(n42), .Z(o[95]) );
  AND U47 ( .A(n43), .B(n44), .Z(n42) );
  AND U48 ( .A(n45), .B(p_input[395]), .Z(n44) );
  AND U49 ( .A(p_input[295]), .B(p_input[195]), .Z(n45) );
  AND U50 ( .A(p_input[595]), .B(p_input[495]), .Z(n43) );
  AND U51 ( .A(n46), .B(n47), .Z(n41) );
  AND U52 ( .A(n48), .B(p_input[895]), .Z(n47) );
  AND U53 ( .A(p_input[795]), .B(p_input[695]), .Z(n48) );
  AND U54 ( .A(p_input[995]), .B(p_input[95]), .Z(n46) );
  AND U55 ( .A(n49), .B(n50), .Z(o[94]) );
  AND U56 ( .A(n51), .B(n52), .Z(n50) );
  AND U57 ( .A(n53), .B(p_input[394]), .Z(n52) );
  AND U58 ( .A(p_input[294]), .B(p_input[194]), .Z(n53) );
  AND U59 ( .A(p_input[594]), .B(p_input[494]), .Z(n51) );
  AND U60 ( .A(n54), .B(n55), .Z(n49) );
  AND U61 ( .A(n56), .B(p_input[894]), .Z(n55) );
  AND U62 ( .A(p_input[794]), .B(p_input[694]), .Z(n56) );
  AND U63 ( .A(p_input[994]), .B(p_input[94]), .Z(n54) );
  AND U64 ( .A(n57), .B(n58), .Z(o[93]) );
  AND U65 ( .A(n59), .B(n60), .Z(n58) );
  AND U66 ( .A(n61), .B(p_input[393]), .Z(n60) );
  AND U67 ( .A(p_input[293]), .B(p_input[193]), .Z(n61) );
  AND U68 ( .A(p_input[593]), .B(p_input[493]), .Z(n59) );
  AND U69 ( .A(n62), .B(n63), .Z(n57) );
  AND U70 ( .A(n64), .B(p_input[893]), .Z(n63) );
  AND U71 ( .A(p_input[793]), .B(p_input[693]), .Z(n64) );
  AND U72 ( .A(p_input[993]), .B(p_input[93]), .Z(n62) );
  AND U73 ( .A(n65), .B(n66), .Z(o[92]) );
  AND U74 ( .A(n67), .B(n68), .Z(n66) );
  AND U75 ( .A(n69), .B(p_input[392]), .Z(n68) );
  AND U76 ( .A(p_input[292]), .B(p_input[192]), .Z(n69) );
  AND U77 ( .A(p_input[592]), .B(p_input[492]), .Z(n67) );
  AND U78 ( .A(n70), .B(n71), .Z(n65) );
  AND U79 ( .A(n72), .B(p_input[892]), .Z(n71) );
  AND U80 ( .A(p_input[792]), .B(p_input[692]), .Z(n72) );
  AND U81 ( .A(p_input[992]), .B(p_input[92]), .Z(n70) );
  AND U82 ( .A(n73), .B(n74), .Z(o[91]) );
  AND U83 ( .A(n75), .B(n76), .Z(n74) );
  AND U84 ( .A(n77), .B(p_input[391]), .Z(n76) );
  AND U85 ( .A(p_input[291]), .B(p_input[191]), .Z(n77) );
  AND U86 ( .A(p_input[591]), .B(p_input[491]), .Z(n75) );
  AND U87 ( .A(n78), .B(n79), .Z(n73) );
  AND U88 ( .A(n80), .B(p_input[891]), .Z(n79) );
  AND U89 ( .A(p_input[791]), .B(p_input[691]), .Z(n80) );
  AND U90 ( .A(p_input[991]), .B(p_input[91]), .Z(n78) );
  AND U91 ( .A(n81), .B(n82), .Z(o[90]) );
  AND U92 ( .A(n83), .B(n84), .Z(n82) );
  AND U93 ( .A(n85), .B(p_input[390]), .Z(n84) );
  AND U94 ( .A(p_input[290]), .B(p_input[190]), .Z(n85) );
  AND U95 ( .A(p_input[590]), .B(p_input[490]), .Z(n83) );
  AND U96 ( .A(n86), .B(n87), .Z(n81) );
  AND U97 ( .A(n88), .B(p_input[890]), .Z(n87) );
  AND U98 ( .A(p_input[790]), .B(p_input[690]), .Z(n88) );
  AND U99 ( .A(p_input[990]), .B(p_input[90]), .Z(n86) );
  AND U100 ( .A(n89), .B(n90), .Z(o[8]) );
  AND U101 ( .A(n91), .B(n92), .Z(n90) );
  AND U102 ( .A(n93), .B(p_input[308]), .Z(n92) );
  AND U103 ( .A(p_input[208]), .B(p_input[108]), .Z(n93) );
  AND U104 ( .A(p_input[508]), .B(p_input[408]), .Z(n91) );
  AND U105 ( .A(n94), .B(n95), .Z(n89) );
  AND U106 ( .A(n96), .B(p_input[808]), .Z(n95) );
  AND U107 ( .A(p_input[708]), .B(p_input[608]), .Z(n96) );
  AND U108 ( .A(p_input[908]), .B(p_input[8]), .Z(n94) );
  AND U109 ( .A(n97), .B(n98), .Z(o[89]) );
  AND U110 ( .A(n99), .B(n100), .Z(n98) );
  AND U111 ( .A(n101), .B(p_input[389]), .Z(n100) );
  AND U112 ( .A(p_input[289]), .B(p_input[189]), .Z(n101) );
  AND U113 ( .A(p_input[589]), .B(p_input[489]), .Z(n99) );
  AND U114 ( .A(n102), .B(n103), .Z(n97) );
  AND U115 ( .A(n104), .B(p_input[889]), .Z(n103) );
  AND U116 ( .A(p_input[789]), .B(p_input[689]), .Z(n104) );
  AND U117 ( .A(p_input[989]), .B(p_input[89]), .Z(n102) );
  AND U118 ( .A(n105), .B(n106), .Z(o[88]) );
  AND U119 ( .A(n107), .B(n108), .Z(n106) );
  AND U120 ( .A(n109), .B(p_input[388]), .Z(n108) );
  AND U121 ( .A(p_input[288]), .B(p_input[188]), .Z(n109) );
  AND U122 ( .A(p_input[588]), .B(p_input[488]), .Z(n107) );
  AND U123 ( .A(n110), .B(n111), .Z(n105) );
  AND U124 ( .A(n112), .B(p_input[888]), .Z(n111) );
  AND U125 ( .A(p_input[788]), .B(p_input[688]), .Z(n112) );
  AND U126 ( .A(p_input[988]), .B(p_input[88]), .Z(n110) );
  AND U127 ( .A(n113), .B(n114), .Z(o[87]) );
  AND U128 ( .A(n115), .B(n116), .Z(n114) );
  AND U129 ( .A(n117), .B(p_input[387]), .Z(n116) );
  AND U130 ( .A(p_input[287]), .B(p_input[187]), .Z(n117) );
  AND U131 ( .A(p_input[587]), .B(p_input[487]), .Z(n115) );
  AND U132 ( .A(n118), .B(n119), .Z(n113) );
  AND U133 ( .A(n120), .B(p_input[87]), .Z(n119) );
  AND U134 ( .A(p_input[787]), .B(p_input[687]), .Z(n120) );
  AND U135 ( .A(p_input[987]), .B(p_input[887]), .Z(n118) );
  AND U136 ( .A(n121), .B(n122), .Z(o[86]) );
  AND U137 ( .A(n123), .B(n124), .Z(n122) );
  AND U138 ( .A(n125), .B(p_input[386]), .Z(n124) );
  AND U139 ( .A(p_input[286]), .B(p_input[186]), .Z(n125) );
  AND U140 ( .A(p_input[586]), .B(p_input[486]), .Z(n123) );
  AND U141 ( .A(n126), .B(n127), .Z(n121) );
  AND U142 ( .A(n128), .B(p_input[86]), .Z(n127) );
  AND U143 ( .A(p_input[786]), .B(p_input[686]), .Z(n128) );
  AND U144 ( .A(p_input[986]), .B(p_input[886]), .Z(n126) );
  AND U145 ( .A(n129), .B(n130), .Z(o[85]) );
  AND U146 ( .A(n131), .B(n132), .Z(n130) );
  AND U147 ( .A(n133), .B(p_input[385]), .Z(n132) );
  AND U148 ( .A(p_input[285]), .B(p_input[185]), .Z(n133) );
  AND U149 ( .A(p_input[585]), .B(p_input[485]), .Z(n131) );
  AND U150 ( .A(n134), .B(n135), .Z(n129) );
  AND U151 ( .A(n136), .B(p_input[85]), .Z(n135) );
  AND U152 ( .A(p_input[785]), .B(p_input[685]), .Z(n136) );
  AND U153 ( .A(p_input[985]), .B(p_input[885]), .Z(n134) );
  AND U154 ( .A(n137), .B(n138), .Z(o[84]) );
  AND U155 ( .A(n139), .B(n140), .Z(n138) );
  AND U156 ( .A(n141), .B(p_input[384]), .Z(n140) );
  AND U157 ( .A(p_input[284]), .B(p_input[184]), .Z(n141) );
  AND U158 ( .A(p_input[584]), .B(p_input[484]), .Z(n139) );
  AND U159 ( .A(n142), .B(n143), .Z(n137) );
  AND U160 ( .A(n144), .B(p_input[84]), .Z(n143) );
  AND U161 ( .A(p_input[784]), .B(p_input[684]), .Z(n144) );
  AND U162 ( .A(p_input[984]), .B(p_input[884]), .Z(n142) );
  AND U163 ( .A(n145), .B(n146), .Z(o[83]) );
  AND U164 ( .A(n147), .B(n148), .Z(n146) );
  AND U165 ( .A(n149), .B(p_input[383]), .Z(n148) );
  AND U166 ( .A(p_input[283]), .B(p_input[183]), .Z(n149) );
  AND U167 ( .A(p_input[583]), .B(p_input[483]), .Z(n147) );
  AND U168 ( .A(n150), .B(n151), .Z(n145) );
  AND U169 ( .A(n152), .B(p_input[83]), .Z(n151) );
  AND U170 ( .A(p_input[783]), .B(p_input[683]), .Z(n152) );
  AND U171 ( .A(p_input[983]), .B(p_input[883]), .Z(n150) );
  AND U172 ( .A(n153), .B(n154), .Z(o[82]) );
  AND U173 ( .A(n155), .B(n156), .Z(n154) );
  AND U174 ( .A(n157), .B(p_input[382]), .Z(n156) );
  AND U175 ( .A(p_input[282]), .B(p_input[182]), .Z(n157) );
  AND U176 ( .A(p_input[582]), .B(p_input[482]), .Z(n155) );
  AND U177 ( .A(n158), .B(n159), .Z(n153) );
  AND U178 ( .A(n160), .B(p_input[82]), .Z(n159) );
  AND U179 ( .A(p_input[782]), .B(p_input[682]), .Z(n160) );
  AND U180 ( .A(p_input[982]), .B(p_input[882]), .Z(n158) );
  AND U181 ( .A(n161), .B(n162), .Z(o[81]) );
  AND U182 ( .A(n163), .B(n164), .Z(n162) );
  AND U183 ( .A(n165), .B(p_input[381]), .Z(n164) );
  AND U184 ( .A(p_input[281]), .B(p_input[181]), .Z(n165) );
  AND U185 ( .A(p_input[581]), .B(p_input[481]), .Z(n163) );
  AND U186 ( .A(n166), .B(n167), .Z(n161) );
  AND U187 ( .A(n168), .B(p_input[81]), .Z(n167) );
  AND U188 ( .A(p_input[781]), .B(p_input[681]), .Z(n168) );
  AND U189 ( .A(p_input[981]), .B(p_input[881]), .Z(n166) );
  AND U190 ( .A(n169), .B(n170), .Z(o[80]) );
  AND U191 ( .A(n171), .B(n172), .Z(n170) );
  AND U192 ( .A(n173), .B(p_input[380]), .Z(n172) );
  AND U193 ( .A(p_input[280]), .B(p_input[180]), .Z(n173) );
  AND U194 ( .A(p_input[580]), .B(p_input[480]), .Z(n171) );
  AND U195 ( .A(n174), .B(n175), .Z(n169) );
  AND U196 ( .A(n176), .B(p_input[80]), .Z(n175) );
  AND U197 ( .A(p_input[780]), .B(p_input[680]), .Z(n176) );
  AND U198 ( .A(p_input[980]), .B(p_input[880]), .Z(n174) );
  AND U199 ( .A(n177), .B(n178), .Z(o[7]) );
  AND U200 ( .A(n179), .B(n180), .Z(n178) );
  AND U201 ( .A(n181), .B(p_input[307]), .Z(n180) );
  AND U202 ( .A(p_input[207]), .B(p_input[107]), .Z(n181) );
  AND U203 ( .A(p_input[507]), .B(p_input[407]), .Z(n179) );
  AND U204 ( .A(n182), .B(n183), .Z(n177) );
  AND U205 ( .A(n184), .B(p_input[7]), .Z(n183) );
  AND U206 ( .A(p_input[707]), .B(p_input[607]), .Z(n184) );
  AND U207 ( .A(p_input[907]), .B(p_input[807]), .Z(n182) );
  AND U208 ( .A(n185), .B(n186), .Z(o[79]) );
  AND U209 ( .A(n187), .B(n188), .Z(n186) );
  AND U210 ( .A(n189), .B(p_input[379]), .Z(n188) );
  AND U211 ( .A(p_input[279]), .B(p_input[179]), .Z(n189) );
  AND U212 ( .A(p_input[579]), .B(p_input[479]), .Z(n187) );
  AND U213 ( .A(n190), .B(n191), .Z(n185) );
  AND U214 ( .A(n192), .B(p_input[79]), .Z(n191) );
  AND U215 ( .A(p_input[779]), .B(p_input[679]), .Z(n192) );
  AND U216 ( .A(p_input[979]), .B(p_input[879]), .Z(n190) );
  AND U217 ( .A(n193), .B(n194), .Z(o[78]) );
  AND U218 ( .A(n195), .B(n196), .Z(n194) );
  AND U219 ( .A(n197), .B(p_input[378]), .Z(n196) );
  AND U220 ( .A(p_input[278]), .B(p_input[178]), .Z(n197) );
  AND U221 ( .A(p_input[578]), .B(p_input[478]), .Z(n195) );
  AND U222 ( .A(n198), .B(n199), .Z(n193) );
  AND U223 ( .A(n200), .B(p_input[78]), .Z(n199) );
  AND U224 ( .A(p_input[778]), .B(p_input[678]), .Z(n200) );
  AND U225 ( .A(p_input[978]), .B(p_input[878]), .Z(n198) );
  AND U226 ( .A(n201), .B(n202), .Z(o[77]) );
  AND U227 ( .A(n203), .B(n204), .Z(n202) );
  AND U228 ( .A(n205), .B(p_input[377]), .Z(n204) );
  AND U229 ( .A(p_input[277]), .B(p_input[177]), .Z(n205) );
  AND U230 ( .A(p_input[577]), .B(p_input[477]), .Z(n203) );
  AND U231 ( .A(n206), .B(n207), .Z(n201) );
  AND U232 ( .A(n208), .B(p_input[77]), .Z(n207) );
  AND U233 ( .A(p_input[777]), .B(p_input[677]), .Z(n208) );
  AND U234 ( .A(p_input[977]), .B(p_input[877]), .Z(n206) );
  AND U235 ( .A(n209), .B(n210), .Z(o[76]) );
  AND U236 ( .A(n211), .B(n212), .Z(n210) );
  AND U237 ( .A(n213), .B(p_input[376]), .Z(n212) );
  AND U238 ( .A(p_input[276]), .B(p_input[176]), .Z(n213) );
  AND U239 ( .A(p_input[576]), .B(p_input[476]), .Z(n211) );
  AND U240 ( .A(n214), .B(n215), .Z(n209) );
  AND U241 ( .A(n216), .B(p_input[776]), .Z(n215) );
  AND U242 ( .A(p_input[76]), .B(p_input[676]), .Z(n216) );
  AND U243 ( .A(p_input[976]), .B(p_input[876]), .Z(n214) );
  AND U244 ( .A(n217), .B(n218), .Z(o[75]) );
  AND U245 ( .A(n219), .B(n220), .Z(n218) );
  AND U246 ( .A(n221), .B(p_input[375]), .Z(n220) );
  AND U247 ( .A(p_input[275]), .B(p_input[175]), .Z(n221) );
  AND U248 ( .A(p_input[575]), .B(p_input[475]), .Z(n219) );
  AND U249 ( .A(n222), .B(n223), .Z(n217) );
  AND U250 ( .A(n224), .B(p_input[775]), .Z(n223) );
  AND U251 ( .A(p_input[75]), .B(p_input[675]), .Z(n224) );
  AND U252 ( .A(p_input[975]), .B(p_input[875]), .Z(n222) );
  AND U253 ( .A(n225), .B(n226), .Z(o[74]) );
  AND U254 ( .A(n227), .B(n228), .Z(n226) );
  AND U255 ( .A(n229), .B(p_input[374]), .Z(n228) );
  AND U256 ( .A(p_input[274]), .B(p_input[174]), .Z(n229) );
  AND U257 ( .A(p_input[574]), .B(p_input[474]), .Z(n227) );
  AND U258 ( .A(n230), .B(n231), .Z(n225) );
  AND U259 ( .A(n232), .B(p_input[774]), .Z(n231) );
  AND U260 ( .A(p_input[74]), .B(p_input[674]), .Z(n232) );
  AND U261 ( .A(p_input[974]), .B(p_input[874]), .Z(n230) );
  AND U262 ( .A(n233), .B(n234), .Z(o[73]) );
  AND U263 ( .A(n235), .B(n236), .Z(n234) );
  AND U264 ( .A(n237), .B(p_input[373]), .Z(n236) );
  AND U265 ( .A(p_input[273]), .B(p_input[173]), .Z(n237) );
  AND U266 ( .A(p_input[573]), .B(p_input[473]), .Z(n235) );
  AND U267 ( .A(n238), .B(n239), .Z(n233) );
  AND U268 ( .A(n240), .B(p_input[773]), .Z(n239) );
  AND U269 ( .A(p_input[73]), .B(p_input[673]), .Z(n240) );
  AND U270 ( .A(p_input[973]), .B(p_input[873]), .Z(n238) );
  AND U271 ( .A(n241), .B(n242), .Z(o[72]) );
  AND U272 ( .A(n243), .B(n244), .Z(n242) );
  AND U273 ( .A(n245), .B(p_input[372]), .Z(n244) );
  AND U274 ( .A(p_input[272]), .B(p_input[172]), .Z(n245) );
  AND U275 ( .A(p_input[572]), .B(p_input[472]), .Z(n243) );
  AND U276 ( .A(n246), .B(n247), .Z(n241) );
  AND U277 ( .A(n248), .B(p_input[772]), .Z(n247) );
  AND U278 ( .A(p_input[72]), .B(p_input[672]), .Z(n248) );
  AND U279 ( .A(p_input[972]), .B(p_input[872]), .Z(n246) );
  AND U280 ( .A(n249), .B(n250), .Z(o[71]) );
  AND U281 ( .A(n251), .B(n252), .Z(n250) );
  AND U282 ( .A(n253), .B(p_input[371]), .Z(n252) );
  AND U283 ( .A(p_input[271]), .B(p_input[171]), .Z(n253) );
  AND U284 ( .A(p_input[571]), .B(p_input[471]), .Z(n251) );
  AND U285 ( .A(n254), .B(n255), .Z(n249) );
  AND U286 ( .A(n256), .B(p_input[771]), .Z(n255) );
  AND U287 ( .A(p_input[71]), .B(p_input[671]), .Z(n256) );
  AND U288 ( .A(p_input[971]), .B(p_input[871]), .Z(n254) );
  AND U289 ( .A(n257), .B(n258), .Z(o[70]) );
  AND U290 ( .A(n259), .B(n260), .Z(n258) );
  AND U291 ( .A(n261), .B(p_input[370]), .Z(n260) );
  AND U292 ( .A(p_input[270]), .B(p_input[170]), .Z(n261) );
  AND U293 ( .A(p_input[570]), .B(p_input[470]), .Z(n259) );
  AND U294 ( .A(n262), .B(n263), .Z(n257) );
  AND U295 ( .A(n264), .B(p_input[770]), .Z(n263) );
  AND U296 ( .A(p_input[70]), .B(p_input[670]), .Z(n264) );
  AND U297 ( .A(p_input[970]), .B(p_input[870]), .Z(n262) );
  AND U298 ( .A(n265), .B(n266), .Z(o[6]) );
  AND U299 ( .A(n267), .B(n268), .Z(n266) );
  AND U300 ( .A(n269), .B(p_input[306]), .Z(n268) );
  AND U301 ( .A(p_input[206]), .B(p_input[106]), .Z(n269) );
  AND U302 ( .A(p_input[506]), .B(p_input[406]), .Z(n267) );
  AND U303 ( .A(n270), .B(n271), .Z(n265) );
  AND U304 ( .A(n272), .B(p_input[706]), .Z(n271) );
  AND U305 ( .A(p_input[6]), .B(p_input[606]), .Z(n272) );
  AND U306 ( .A(p_input[906]), .B(p_input[806]), .Z(n270) );
  AND U307 ( .A(n273), .B(n274), .Z(o[69]) );
  AND U308 ( .A(n275), .B(n276), .Z(n274) );
  AND U309 ( .A(n277), .B(p_input[369]), .Z(n276) );
  AND U310 ( .A(p_input[269]), .B(p_input[169]), .Z(n277) );
  AND U311 ( .A(p_input[569]), .B(p_input[469]), .Z(n275) );
  AND U312 ( .A(n278), .B(n279), .Z(n273) );
  AND U313 ( .A(n280), .B(p_input[769]), .Z(n279) );
  AND U314 ( .A(p_input[69]), .B(p_input[669]), .Z(n280) );
  AND U315 ( .A(p_input[969]), .B(p_input[869]), .Z(n278) );
  AND U316 ( .A(n281), .B(n282), .Z(o[68]) );
  AND U317 ( .A(n283), .B(n284), .Z(n282) );
  AND U318 ( .A(n285), .B(p_input[368]), .Z(n284) );
  AND U319 ( .A(p_input[268]), .B(p_input[168]), .Z(n285) );
  AND U320 ( .A(p_input[568]), .B(p_input[468]), .Z(n283) );
  AND U321 ( .A(n286), .B(n287), .Z(n281) );
  AND U322 ( .A(n288), .B(p_input[768]), .Z(n287) );
  AND U323 ( .A(p_input[68]), .B(p_input[668]), .Z(n288) );
  AND U324 ( .A(p_input[968]), .B(p_input[868]), .Z(n286) );
  AND U325 ( .A(n289), .B(n290), .Z(o[67]) );
  AND U326 ( .A(n291), .B(n292), .Z(n290) );
  AND U327 ( .A(n293), .B(p_input[367]), .Z(n292) );
  AND U328 ( .A(p_input[267]), .B(p_input[167]), .Z(n293) );
  AND U329 ( .A(p_input[567]), .B(p_input[467]), .Z(n291) );
  AND U330 ( .A(n294), .B(n295), .Z(n289) );
  AND U331 ( .A(n296), .B(p_input[767]), .Z(n295) );
  AND U332 ( .A(p_input[67]), .B(p_input[667]), .Z(n296) );
  AND U333 ( .A(p_input[967]), .B(p_input[867]), .Z(n294) );
  AND U334 ( .A(n297), .B(n298), .Z(o[66]) );
  AND U335 ( .A(n299), .B(n300), .Z(n298) );
  AND U336 ( .A(n301), .B(p_input[366]), .Z(n300) );
  AND U337 ( .A(p_input[266]), .B(p_input[166]), .Z(n301) );
  AND U338 ( .A(p_input[566]), .B(p_input[466]), .Z(n299) );
  AND U339 ( .A(n302), .B(n303), .Z(n297) );
  AND U340 ( .A(n304), .B(p_input[766]), .Z(n303) );
  AND U341 ( .A(p_input[66]), .B(p_input[666]), .Z(n304) );
  AND U342 ( .A(p_input[966]), .B(p_input[866]), .Z(n302) );
  AND U343 ( .A(n305), .B(n306), .Z(o[65]) );
  AND U344 ( .A(n307), .B(n308), .Z(n306) );
  AND U345 ( .A(n309), .B(p_input[365]), .Z(n308) );
  AND U346 ( .A(p_input[265]), .B(p_input[165]), .Z(n309) );
  AND U347 ( .A(p_input[565]), .B(p_input[465]), .Z(n307) );
  AND U348 ( .A(n310), .B(n311), .Z(n305) );
  AND U349 ( .A(n312), .B(p_input[765]), .Z(n311) );
  AND U350 ( .A(p_input[665]), .B(p_input[65]), .Z(n312) );
  AND U351 ( .A(p_input[965]), .B(p_input[865]), .Z(n310) );
  AND U352 ( .A(n313), .B(n314), .Z(o[64]) );
  AND U353 ( .A(n315), .B(n316), .Z(n314) );
  AND U354 ( .A(n317), .B(p_input[364]), .Z(n316) );
  AND U355 ( .A(p_input[264]), .B(p_input[164]), .Z(n317) );
  AND U356 ( .A(p_input[564]), .B(p_input[464]), .Z(n315) );
  AND U357 ( .A(n318), .B(n319), .Z(n313) );
  AND U358 ( .A(n320), .B(p_input[764]), .Z(n319) );
  AND U359 ( .A(p_input[664]), .B(p_input[64]), .Z(n320) );
  AND U360 ( .A(p_input[964]), .B(p_input[864]), .Z(n318) );
  AND U361 ( .A(n321), .B(n322), .Z(o[63]) );
  AND U362 ( .A(n323), .B(n324), .Z(n322) );
  AND U363 ( .A(n325), .B(p_input[363]), .Z(n324) );
  AND U364 ( .A(p_input[263]), .B(p_input[163]), .Z(n325) );
  AND U365 ( .A(p_input[563]), .B(p_input[463]), .Z(n323) );
  AND U366 ( .A(n326), .B(n327), .Z(n321) );
  AND U367 ( .A(n328), .B(p_input[763]), .Z(n327) );
  AND U368 ( .A(p_input[663]), .B(p_input[63]), .Z(n328) );
  AND U369 ( .A(p_input[963]), .B(p_input[863]), .Z(n326) );
  AND U370 ( .A(n329), .B(n330), .Z(o[62]) );
  AND U371 ( .A(n331), .B(n332), .Z(n330) );
  AND U372 ( .A(n333), .B(p_input[362]), .Z(n332) );
  AND U373 ( .A(p_input[262]), .B(p_input[162]), .Z(n333) );
  AND U374 ( .A(p_input[562]), .B(p_input[462]), .Z(n331) );
  AND U375 ( .A(n334), .B(n335), .Z(n329) );
  AND U376 ( .A(n336), .B(p_input[762]), .Z(n335) );
  AND U377 ( .A(p_input[662]), .B(p_input[62]), .Z(n336) );
  AND U378 ( .A(p_input[962]), .B(p_input[862]), .Z(n334) );
  AND U379 ( .A(n337), .B(n338), .Z(o[61]) );
  AND U380 ( .A(n339), .B(n340), .Z(n338) );
  AND U381 ( .A(n341), .B(p_input[361]), .Z(n340) );
  AND U382 ( .A(p_input[261]), .B(p_input[161]), .Z(n341) );
  AND U383 ( .A(p_input[561]), .B(p_input[461]), .Z(n339) );
  AND U384 ( .A(n342), .B(n343), .Z(n337) );
  AND U385 ( .A(n344), .B(p_input[761]), .Z(n343) );
  AND U386 ( .A(p_input[661]), .B(p_input[61]), .Z(n344) );
  AND U387 ( .A(p_input[961]), .B(p_input[861]), .Z(n342) );
  AND U388 ( .A(n345), .B(n346), .Z(o[60]) );
  AND U389 ( .A(n347), .B(n348), .Z(n346) );
  AND U390 ( .A(n349), .B(p_input[360]), .Z(n348) );
  AND U391 ( .A(p_input[260]), .B(p_input[160]), .Z(n349) );
  AND U392 ( .A(p_input[560]), .B(p_input[460]), .Z(n347) );
  AND U393 ( .A(n350), .B(n351), .Z(n345) );
  AND U394 ( .A(n352), .B(p_input[760]), .Z(n351) );
  AND U395 ( .A(p_input[660]), .B(p_input[60]), .Z(n352) );
  AND U396 ( .A(p_input[960]), .B(p_input[860]), .Z(n350) );
  AND U397 ( .A(n353), .B(n354), .Z(o[5]) );
  AND U398 ( .A(n355), .B(n356), .Z(n354) );
  AND U399 ( .A(n357), .B(p_input[305]), .Z(n356) );
  AND U400 ( .A(p_input[205]), .B(p_input[105]), .Z(n357) );
  AND U401 ( .A(p_input[505]), .B(p_input[405]), .Z(n355) );
  AND U402 ( .A(n358), .B(n359), .Z(n353) );
  AND U403 ( .A(n360), .B(p_input[705]), .Z(n359) );
  AND U404 ( .A(p_input[605]), .B(p_input[5]), .Z(n360) );
  AND U405 ( .A(p_input[905]), .B(p_input[805]), .Z(n358) );
  AND U406 ( .A(n361), .B(n362), .Z(o[59]) );
  AND U407 ( .A(n363), .B(n364), .Z(n362) );
  AND U408 ( .A(n365), .B(p_input[359]), .Z(n364) );
  AND U409 ( .A(p_input[259]), .B(p_input[159]), .Z(n365) );
  AND U410 ( .A(p_input[559]), .B(p_input[459]), .Z(n363) );
  AND U411 ( .A(n366), .B(n367), .Z(n361) );
  AND U412 ( .A(n368), .B(p_input[759]), .Z(n367) );
  AND U413 ( .A(p_input[659]), .B(p_input[59]), .Z(n368) );
  AND U414 ( .A(p_input[959]), .B(p_input[859]), .Z(n366) );
  AND U415 ( .A(n369), .B(n370), .Z(o[58]) );
  AND U416 ( .A(n371), .B(n372), .Z(n370) );
  AND U417 ( .A(n373), .B(p_input[358]), .Z(n372) );
  AND U418 ( .A(p_input[258]), .B(p_input[158]), .Z(n373) );
  AND U419 ( .A(p_input[558]), .B(p_input[458]), .Z(n371) );
  AND U420 ( .A(n374), .B(n375), .Z(n369) );
  AND U421 ( .A(n376), .B(p_input[758]), .Z(n375) );
  AND U422 ( .A(p_input[658]), .B(p_input[58]), .Z(n376) );
  AND U423 ( .A(p_input[958]), .B(p_input[858]), .Z(n374) );
  AND U424 ( .A(n377), .B(n378), .Z(o[57]) );
  AND U425 ( .A(n379), .B(n380), .Z(n378) );
  AND U426 ( .A(n381), .B(p_input[357]), .Z(n380) );
  AND U427 ( .A(p_input[257]), .B(p_input[157]), .Z(n381) );
  AND U428 ( .A(p_input[557]), .B(p_input[457]), .Z(n379) );
  AND U429 ( .A(n382), .B(n383), .Z(n377) );
  AND U430 ( .A(n384), .B(p_input[757]), .Z(n383) );
  AND U431 ( .A(p_input[657]), .B(p_input[57]), .Z(n384) );
  AND U432 ( .A(p_input[957]), .B(p_input[857]), .Z(n382) );
  AND U433 ( .A(n385), .B(n386), .Z(o[56]) );
  AND U434 ( .A(n387), .B(n388), .Z(n386) );
  AND U435 ( .A(n389), .B(p_input[356]), .Z(n388) );
  AND U436 ( .A(p_input[256]), .B(p_input[156]), .Z(n389) );
  AND U437 ( .A(p_input[556]), .B(p_input[456]), .Z(n387) );
  AND U438 ( .A(n390), .B(n391), .Z(n385) );
  AND U439 ( .A(n392), .B(p_input[756]), .Z(n391) );
  AND U440 ( .A(p_input[656]), .B(p_input[56]), .Z(n392) );
  AND U441 ( .A(p_input[956]), .B(p_input[856]), .Z(n390) );
  AND U442 ( .A(n393), .B(n394), .Z(o[55]) );
  AND U443 ( .A(n395), .B(n396), .Z(n394) );
  AND U444 ( .A(n397), .B(p_input[355]), .Z(n396) );
  AND U445 ( .A(p_input[255]), .B(p_input[155]), .Z(n397) );
  AND U446 ( .A(p_input[555]), .B(p_input[455]), .Z(n395) );
  AND U447 ( .A(n398), .B(n399), .Z(n393) );
  AND U448 ( .A(n400), .B(p_input[755]), .Z(n399) );
  AND U449 ( .A(p_input[655]), .B(p_input[55]), .Z(n400) );
  AND U450 ( .A(p_input[955]), .B(p_input[855]), .Z(n398) );
  AND U451 ( .A(n401), .B(n402), .Z(o[54]) );
  AND U452 ( .A(n403), .B(n404), .Z(n402) );
  AND U453 ( .A(n405), .B(p_input[354]), .Z(n404) );
  AND U454 ( .A(p_input[254]), .B(p_input[154]), .Z(n405) );
  AND U455 ( .A(p_input[54]), .B(p_input[454]), .Z(n403) );
  AND U456 ( .A(n406), .B(n407), .Z(n401) );
  AND U457 ( .A(n408), .B(p_input[754]), .Z(n407) );
  AND U458 ( .A(p_input[654]), .B(p_input[554]), .Z(n408) );
  AND U459 ( .A(p_input[954]), .B(p_input[854]), .Z(n406) );
  AND U460 ( .A(n409), .B(n410), .Z(o[53]) );
  AND U461 ( .A(n411), .B(n412), .Z(n410) );
  AND U462 ( .A(n413), .B(p_input[353]), .Z(n412) );
  AND U463 ( .A(p_input[253]), .B(p_input[153]), .Z(n413) );
  AND U464 ( .A(p_input[53]), .B(p_input[453]), .Z(n411) );
  AND U465 ( .A(n414), .B(n415), .Z(n409) );
  AND U466 ( .A(n416), .B(p_input[753]), .Z(n415) );
  AND U467 ( .A(p_input[653]), .B(p_input[553]), .Z(n416) );
  AND U468 ( .A(p_input[953]), .B(p_input[853]), .Z(n414) );
  AND U469 ( .A(n417), .B(n418), .Z(o[52]) );
  AND U470 ( .A(n419), .B(n420), .Z(n418) );
  AND U471 ( .A(n421), .B(p_input[352]), .Z(n420) );
  AND U472 ( .A(p_input[252]), .B(p_input[152]), .Z(n421) );
  AND U473 ( .A(p_input[52]), .B(p_input[452]), .Z(n419) );
  AND U474 ( .A(n422), .B(n423), .Z(n417) );
  AND U475 ( .A(n424), .B(p_input[752]), .Z(n423) );
  AND U476 ( .A(p_input[652]), .B(p_input[552]), .Z(n424) );
  AND U477 ( .A(p_input[952]), .B(p_input[852]), .Z(n422) );
  AND U478 ( .A(n425), .B(n426), .Z(o[51]) );
  AND U479 ( .A(n427), .B(n428), .Z(n426) );
  AND U480 ( .A(n429), .B(p_input[351]), .Z(n428) );
  AND U481 ( .A(p_input[251]), .B(p_input[151]), .Z(n429) );
  AND U482 ( .A(p_input[51]), .B(p_input[451]), .Z(n427) );
  AND U483 ( .A(n430), .B(n431), .Z(n425) );
  AND U484 ( .A(n432), .B(p_input[751]), .Z(n431) );
  AND U485 ( .A(p_input[651]), .B(p_input[551]), .Z(n432) );
  AND U486 ( .A(p_input[951]), .B(p_input[851]), .Z(n430) );
  AND U487 ( .A(n433), .B(n434), .Z(o[50]) );
  AND U488 ( .A(n435), .B(n436), .Z(n434) );
  AND U489 ( .A(n437), .B(p_input[350]), .Z(n436) );
  AND U490 ( .A(p_input[250]), .B(p_input[150]), .Z(n437) );
  AND U491 ( .A(p_input[50]), .B(p_input[450]), .Z(n435) );
  AND U492 ( .A(n438), .B(n439), .Z(n433) );
  AND U493 ( .A(n440), .B(p_input[750]), .Z(n439) );
  AND U494 ( .A(p_input[650]), .B(p_input[550]), .Z(n440) );
  AND U495 ( .A(p_input[950]), .B(p_input[850]), .Z(n438) );
  AND U496 ( .A(n441), .B(n442), .Z(o[4]) );
  AND U497 ( .A(n443), .B(n444), .Z(n442) );
  AND U498 ( .A(n445), .B(p_input[304]), .Z(n444) );
  AND U499 ( .A(p_input[204]), .B(p_input[104]), .Z(n445) );
  AND U500 ( .A(p_input[4]), .B(p_input[404]), .Z(n443) );
  AND U501 ( .A(n446), .B(n447), .Z(n441) );
  AND U502 ( .A(n448), .B(p_input[704]), .Z(n447) );
  AND U503 ( .A(p_input[604]), .B(p_input[504]), .Z(n448) );
  AND U504 ( .A(p_input[904]), .B(p_input[804]), .Z(n446) );
  AND U505 ( .A(n449), .B(n450), .Z(o[49]) );
  AND U506 ( .A(n451), .B(n452), .Z(n450) );
  AND U507 ( .A(n453), .B(p_input[349]), .Z(n452) );
  AND U508 ( .A(p_input[249]), .B(p_input[149]), .Z(n453) );
  AND U509 ( .A(p_input[49]), .B(p_input[449]), .Z(n451) );
  AND U510 ( .A(n454), .B(n455), .Z(n449) );
  AND U511 ( .A(n456), .B(p_input[749]), .Z(n455) );
  AND U512 ( .A(p_input[649]), .B(p_input[549]), .Z(n456) );
  AND U513 ( .A(p_input[949]), .B(p_input[849]), .Z(n454) );
  AND U514 ( .A(n457), .B(n458), .Z(o[48]) );
  AND U515 ( .A(n459), .B(n460), .Z(n458) );
  AND U516 ( .A(n461), .B(p_input[348]), .Z(n460) );
  AND U517 ( .A(p_input[248]), .B(p_input[148]), .Z(n461) );
  AND U518 ( .A(p_input[48]), .B(p_input[448]), .Z(n459) );
  AND U519 ( .A(n462), .B(n463), .Z(n457) );
  AND U520 ( .A(n464), .B(p_input[748]), .Z(n463) );
  AND U521 ( .A(p_input[648]), .B(p_input[548]), .Z(n464) );
  AND U522 ( .A(p_input[948]), .B(p_input[848]), .Z(n462) );
  AND U523 ( .A(n465), .B(n466), .Z(o[47]) );
  AND U524 ( .A(n467), .B(n468), .Z(n466) );
  AND U525 ( .A(n469), .B(p_input[347]), .Z(n468) );
  AND U526 ( .A(p_input[247]), .B(p_input[147]), .Z(n469) );
  AND U527 ( .A(p_input[47]), .B(p_input[447]), .Z(n467) );
  AND U528 ( .A(n470), .B(n471), .Z(n465) );
  AND U529 ( .A(n472), .B(p_input[747]), .Z(n471) );
  AND U530 ( .A(p_input[647]), .B(p_input[547]), .Z(n472) );
  AND U531 ( .A(p_input[947]), .B(p_input[847]), .Z(n470) );
  AND U532 ( .A(n473), .B(n474), .Z(o[46]) );
  AND U533 ( .A(n475), .B(n476), .Z(n474) );
  AND U534 ( .A(n477), .B(p_input[346]), .Z(n476) );
  AND U535 ( .A(p_input[246]), .B(p_input[146]), .Z(n477) );
  AND U536 ( .A(p_input[46]), .B(p_input[446]), .Z(n475) );
  AND U537 ( .A(n478), .B(n479), .Z(n473) );
  AND U538 ( .A(n480), .B(p_input[746]), .Z(n479) );
  AND U539 ( .A(p_input[646]), .B(p_input[546]), .Z(n480) );
  AND U540 ( .A(p_input[946]), .B(p_input[846]), .Z(n478) );
  AND U541 ( .A(n481), .B(n482), .Z(o[45]) );
  AND U542 ( .A(n483), .B(n484), .Z(n482) );
  AND U543 ( .A(n485), .B(p_input[345]), .Z(n484) );
  AND U544 ( .A(p_input[245]), .B(p_input[145]), .Z(n485) );
  AND U545 ( .A(p_input[45]), .B(p_input[445]), .Z(n483) );
  AND U546 ( .A(n486), .B(n487), .Z(n481) );
  AND U547 ( .A(n488), .B(p_input[745]), .Z(n487) );
  AND U548 ( .A(p_input[645]), .B(p_input[545]), .Z(n488) );
  AND U549 ( .A(p_input[945]), .B(p_input[845]), .Z(n486) );
  AND U550 ( .A(n489), .B(n490), .Z(o[44]) );
  AND U551 ( .A(n491), .B(n492), .Z(n490) );
  AND U552 ( .A(n493), .B(p_input[344]), .Z(n492) );
  AND U553 ( .A(p_input[244]), .B(p_input[144]), .Z(n493) );
  AND U554 ( .A(p_input[44]), .B(p_input[444]), .Z(n491) );
  AND U555 ( .A(n494), .B(n495), .Z(n489) );
  AND U556 ( .A(n496), .B(p_input[744]), .Z(n495) );
  AND U557 ( .A(p_input[644]), .B(p_input[544]), .Z(n496) );
  AND U558 ( .A(p_input[944]), .B(p_input[844]), .Z(n494) );
  AND U559 ( .A(n497), .B(n498), .Z(o[43]) );
  AND U560 ( .A(n499), .B(n500), .Z(n498) );
  AND U561 ( .A(n501), .B(p_input[343]), .Z(n500) );
  AND U562 ( .A(p_input[243]), .B(p_input[143]), .Z(n501) );
  AND U563 ( .A(p_input[443]), .B(p_input[43]), .Z(n499) );
  AND U564 ( .A(n502), .B(n503), .Z(n497) );
  AND U565 ( .A(n504), .B(p_input[743]), .Z(n503) );
  AND U566 ( .A(p_input[643]), .B(p_input[543]), .Z(n504) );
  AND U567 ( .A(p_input[943]), .B(p_input[843]), .Z(n502) );
  AND U568 ( .A(n505), .B(n506), .Z(o[42]) );
  AND U569 ( .A(n507), .B(n508), .Z(n506) );
  AND U570 ( .A(n509), .B(p_input[342]), .Z(n508) );
  AND U571 ( .A(p_input[242]), .B(p_input[142]), .Z(n509) );
  AND U572 ( .A(p_input[442]), .B(p_input[42]), .Z(n507) );
  AND U573 ( .A(n510), .B(n511), .Z(n505) );
  AND U574 ( .A(n512), .B(p_input[742]), .Z(n511) );
  AND U575 ( .A(p_input[642]), .B(p_input[542]), .Z(n512) );
  AND U576 ( .A(p_input[942]), .B(p_input[842]), .Z(n510) );
  AND U577 ( .A(n513), .B(n514), .Z(o[41]) );
  AND U578 ( .A(n515), .B(n516), .Z(n514) );
  AND U579 ( .A(n517), .B(p_input[341]), .Z(n516) );
  AND U580 ( .A(p_input[241]), .B(p_input[141]), .Z(n517) );
  AND U581 ( .A(p_input[441]), .B(p_input[41]), .Z(n515) );
  AND U582 ( .A(n518), .B(n519), .Z(n513) );
  AND U583 ( .A(n520), .B(p_input[741]), .Z(n519) );
  AND U584 ( .A(p_input[641]), .B(p_input[541]), .Z(n520) );
  AND U585 ( .A(p_input[941]), .B(p_input[841]), .Z(n518) );
  AND U586 ( .A(n521), .B(n522), .Z(o[40]) );
  AND U587 ( .A(n523), .B(n524), .Z(n522) );
  AND U588 ( .A(n525), .B(p_input[340]), .Z(n524) );
  AND U589 ( .A(p_input[240]), .B(p_input[140]), .Z(n525) );
  AND U590 ( .A(p_input[440]), .B(p_input[40]), .Z(n523) );
  AND U591 ( .A(n526), .B(n527), .Z(n521) );
  AND U592 ( .A(n528), .B(p_input[740]), .Z(n527) );
  AND U593 ( .A(p_input[640]), .B(p_input[540]), .Z(n528) );
  AND U594 ( .A(p_input[940]), .B(p_input[840]), .Z(n526) );
  AND U595 ( .A(n529), .B(n530), .Z(o[3]) );
  AND U596 ( .A(n531), .B(n532), .Z(n530) );
  AND U597 ( .A(n533), .B(p_input[303]), .Z(n532) );
  AND U598 ( .A(p_input[203]), .B(p_input[103]), .Z(n533) );
  AND U599 ( .A(p_input[403]), .B(p_input[3]), .Z(n531) );
  AND U600 ( .A(n534), .B(n535), .Z(n529) );
  AND U601 ( .A(n536), .B(p_input[703]), .Z(n535) );
  AND U602 ( .A(p_input[603]), .B(p_input[503]), .Z(n536) );
  AND U603 ( .A(p_input[903]), .B(p_input[803]), .Z(n534) );
  AND U604 ( .A(n537), .B(n538), .Z(o[39]) );
  AND U605 ( .A(n539), .B(n540), .Z(n538) );
  AND U606 ( .A(n541), .B(p_input[339]), .Z(n540) );
  AND U607 ( .A(p_input[239]), .B(p_input[139]), .Z(n541) );
  AND U608 ( .A(p_input[439]), .B(p_input[39]), .Z(n539) );
  AND U609 ( .A(n542), .B(n543), .Z(n537) );
  AND U610 ( .A(n544), .B(p_input[739]), .Z(n543) );
  AND U611 ( .A(p_input[639]), .B(p_input[539]), .Z(n544) );
  AND U612 ( .A(p_input[939]), .B(p_input[839]), .Z(n542) );
  AND U613 ( .A(n545), .B(n546), .Z(o[38]) );
  AND U614 ( .A(n547), .B(n548), .Z(n546) );
  AND U615 ( .A(n549), .B(p_input[338]), .Z(n548) );
  AND U616 ( .A(p_input[238]), .B(p_input[138]), .Z(n549) );
  AND U617 ( .A(p_input[438]), .B(p_input[38]), .Z(n547) );
  AND U618 ( .A(n550), .B(n551), .Z(n545) );
  AND U619 ( .A(n552), .B(p_input[738]), .Z(n551) );
  AND U620 ( .A(p_input[638]), .B(p_input[538]), .Z(n552) );
  AND U621 ( .A(p_input[938]), .B(p_input[838]), .Z(n550) );
  AND U622 ( .A(n553), .B(n554), .Z(o[37]) );
  AND U623 ( .A(n555), .B(n556), .Z(n554) );
  AND U624 ( .A(n557), .B(p_input[337]), .Z(n556) );
  AND U625 ( .A(p_input[237]), .B(p_input[137]), .Z(n557) );
  AND U626 ( .A(p_input[437]), .B(p_input[37]), .Z(n555) );
  AND U627 ( .A(n558), .B(n559), .Z(n553) );
  AND U628 ( .A(n560), .B(p_input[737]), .Z(n559) );
  AND U629 ( .A(p_input[637]), .B(p_input[537]), .Z(n560) );
  AND U630 ( .A(p_input[937]), .B(p_input[837]), .Z(n558) );
  AND U631 ( .A(n561), .B(n562), .Z(o[36]) );
  AND U632 ( .A(n563), .B(n564), .Z(n562) );
  AND U633 ( .A(n565), .B(p_input[336]), .Z(n564) );
  AND U634 ( .A(p_input[236]), .B(p_input[136]), .Z(n565) );
  AND U635 ( .A(p_input[436]), .B(p_input[36]), .Z(n563) );
  AND U636 ( .A(n566), .B(n567), .Z(n561) );
  AND U637 ( .A(n568), .B(p_input[736]), .Z(n567) );
  AND U638 ( .A(p_input[636]), .B(p_input[536]), .Z(n568) );
  AND U639 ( .A(p_input[936]), .B(p_input[836]), .Z(n566) );
  AND U640 ( .A(n569), .B(n570), .Z(o[35]) );
  AND U641 ( .A(n571), .B(n572), .Z(n570) );
  AND U642 ( .A(n573), .B(p_input[335]), .Z(n572) );
  AND U643 ( .A(p_input[235]), .B(p_input[135]), .Z(n573) );
  AND U644 ( .A(p_input[435]), .B(p_input[35]), .Z(n571) );
  AND U645 ( .A(n574), .B(n575), .Z(n569) );
  AND U646 ( .A(n576), .B(p_input[735]), .Z(n575) );
  AND U647 ( .A(p_input[635]), .B(p_input[535]), .Z(n576) );
  AND U648 ( .A(p_input[935]), .B(p_input[835]), .Z(n574) );
  AND U649 ( .A(n577), .B(n578), .Z(o[34]) );
  AND U650 ( .A(n579), .B(n580), .Z(n578) );
  AND U651 ( .A(n581), .B(p_input[334]), .Z(n580) );
  AND U652 ( .A(p_input[234]), .B(p_input[134]), .Z(n581) );
  AND U653 ( .A(p_input[434]), .B(p_input[34]), .Z(n579) );
  AND U654 ( .A(n582), .B(n583), .Z(n577) );
  AND U655 ( .A(n584), .B(p_input[734]), .Z(n583) );
  AND U656 ( .A(p_input[634]), .B(p_input[534]), .Z(n584) );
  AND U657 ( .A(p_input[934]), .B(p_input[834]), .Z(n582) );
  AND U658 ( .A(n585), .B(n586), .Z(o[33]) );
  AND U659 ( .A(n587), .B(n588), .Z(n586) );
  AND U660 ( .A(n589), .B(p_input[333]), .Z(n588) );
  AND U661 ( .A(p_input[233]), .B(p_input[133]), .Z(n589) );
  AND U662 ( .A(p_input[433]), .B(p_input[33]), .Z(n587) );
  AND U663 ( .A(n590), .B(n591), .Z(n585) );
  AND U664 ( .A(n592), .B(p_input[733]), .Z(n591) );
  AND U665 ( .A(p_input[633]), .B(p_input[533]), .Z(n592) );
  AND U666 ( .A(p_input[933]), .B(p_input[833]), .Z(n590) );
  AND U667 ( .A(n593), .B(n594), .Z(o[32]) );
  AND U668 ( .A(n595), .B(n596), .Z(n594) );
  AND U669 ( .A(n597), .B(p_input[32]), .Z(n596) );
  AND U670 ( .A(p_input[232]), .B(p_input[132]), .Z(n597) );
  AND U671 ( .A(p_input[432]), .B(p_input[332]), .Z(n595) );
  AND U672 ( .A(n598), .B(n599), .Z(n593) );
  AND U673 ( .A(n600), .B(p_input[732]), .Z(n599) );
  AND U674 ( .A(p_input[632]), .B(p_input[532]), .Z(n600) );
  AND U675 ( .A(p_input[932]), .B(p_input[832]), .Z(n598) );
  AND U676 ( .A(n601), .B(n602), .Z(o[31]) );
  AND U677 ( .A(n603), .B(n604), .Z(n602) );
  AND U678 ( .A(n605), .B(p_input[31]), .Z(n604) );
  AND U679 ( .A(p_input[231]), .B(p_input[131]), .Z(n605) );
  AND U680 ( .A(p_input[431]), .B(p_input[331]), .Z(n603) );
  AND U681 ( .A(n606), .B(n607), .Z(n601) );
  AND U682 ( .A(n608), .B(p_input[731]), .Z(n607) );
  AND U683 ( .A(p_input[631]), .B(p_input[531]), .Z(n608) );
  AND U684 ( .A(p_input[931]), .B(p_input[831]), .Z(n606) );
  AND U685 ( .A(n609), .B(n610), .Z(o[30]) );
  AND U686 ( .A(n611), .B(n612), .Z(n610) );
  AND U687 ( .A(n613), .B(p_input[30]), .Z(n612) );
  AND U688 ( .A(p_input[230]), .B(p_input[130]), .Z(n613) );
  AND U689 ( .A(p_input[430]), .B(p_input[330]), .Z(n611) );
  AND U690 ( .A(n614), .B(n615), .Z(n609) );
  AND U691 ( .A(n616), .B(p_input[730]), .Z(n615) );
  AND U692 ( .A(p_input[630]), .B(p_input[530]), .Z(n616) );
  AND U693 ( .A(p_input[930]), .B(p_input[830]), .Z(n614) );
  AND U694 ( .A(n617), .B(n618), .Z(o[2]) );
  AND U695 ( .A(n619), .B(n620), .Z(n618) );
  AND U696 ( .A(n621), .B(p_input[2]), .Z(n620) );
  AND U697 ( .A(p_input[202]), .B(p_input[102]), .Z(n621) );
  AND U698 ( .A(p_input[402]), .B(p_input[302]), .Z(n619) );
  AND U699 ( .A(n622), .B(n623), .Z(n617) );
  AND U700 ( .A(n624), .B(p_input[702]), .Z(n623) );
  AND U701 ( .A(p_input[602]), .B(p_input[502]), .Z(n624) );
  AND U702 ( .A(p_input[902]), .B(p_input[802]), .Z(n622) );
  AND U703 ( .A(n625), .B(n626), .Z(o[29]) );
  AND U704 ( .A(n627), .B(n628), .Z(n626) );
  AND U705 ( .A(n629), .B(p_input[29]), .Z(n628) );
  AND U706 ( .A(p_input[229]), .B(p_input[129]), .Z(n629) );
  AND U707 ( .A(p_input[429]), .B(p_input[329]), .Z(n627) );
  AND U708 ( .A(n630), .B(n631), .Z(n625) );
  AND U709 ( .A(n632), .B(p_input[729]), .Z(n631) );
  AND U710 ( .A(p_input[629]), .B(p_input[529]), .Z(n632) );
  AND U711 ( .A(p_input[929]), .B(p_input[829]), .Z(n630) );
  AND U712 ( .A(n633), .B(n634), .Z(o[28]) );
  AND U713 ( .A(n635), .B(n636), .Z(n634) );
  AND U714 ( .A(n637), .B(p_input[28]), .Z(n636) );
  AND U715 ( .A(p_input[228]), .B(p_input[128]), .Z(n637) );
  AND U716 ( .A(p_input[428]), .B(p_input[328]), .Z(n635) );
  AND U717 ( .A(n638), .B(n639), .Z(n633) );
  AND U718 ( .A(n640), .B(p_input[728]), .Z(n639) );
  AND U719 ( .A(p_input[628]), .B(p_input[528]), .Z(n640) );
  AND U720 ( .A(p_input[928]), .B(p_input[828]), .Z(n638) );
  AND U721 ( .A(n641), .B(n642), .Z(o[27]) );
  AND U722 ( .A(n643), .B(n644), .Z(n642) );
  AND U723 ( .A(n645), .B(p_input[27]), .Z(n644) );
  AND U724 ( .A(p_input[227]), .B(p_input[127]), .Z(n645) );
  AND U725 ( .A(p_input[427]), .B(p_input[327]), .Z(n643) );
  AND U726 ( .A(n646), .B(n647), .Z(n641) );
  AND U727 ( .A(n648), .B(p_input[727]), .Z(n647) );
  AND U728 ( .A(p_input[627]), .B(p_input[527]), .Z(n648) );
  AND U729 ( .A(p_input[927]), .B(p_input[827]), .Z(n646) );
  AND U730 ( .A(n649), .B(n650), .Z(o[26]) );
  AND U731 ( .A(n651), .B(n652), .Z(n650) );
  AND U732 ( .A(n653), .B(p_input[26]), .Z(n652) );
  AND U733 ( .A(p_input[226]), .B(p_input[126]), .Z(n653) );
  AND U734 ( .A(p_input[426]), .B(p_input[326]), .Z(n651) );
  AND U735 ( .A(n654), .B(n655), .Z(n649) );
  AND U736 ( .A(n656), .B(p_input[726]), .Z(n655) );
  AND U737 ( .A(p_input[626]), .B(p_input[526]), .Z(n656) );
  AND U738 ( .A(p_input[926]), .B(p_input[826]), .Z(n654) );
  AND U739 ( .A(n657), .B(n658), .Z(o[25]) );
  AND U740 ( .A(n659), .B(n660), .Z(n658) );
  AND U741 ( .A(n661), .B(p_input[25]), .Z(n660) );
  AND U742 ( .A(p_input[225]), .B(p_input[125]), .Z(n661) );
  AND U743 ( .A(p_input[425]), .B(p_input[325]), .Z(n659) );
  AND U744 ( .A(n662), .B(n663), .Z(n657) );
  AND U745 ( .A(n664), .B(p_input[725]), .Z(n663) );
  AND U746 ( .A(p_input[625]), .B(p_input[525]), .Z(n664) );
  AND U747 ( .A(p_input[925]), .B(p_input[825]), .Z(n662) );
  AND U748 ( .A(n665), .B(n666), .Z(o[24]) );
  AND U749 ( .A(n667), .B(n668), .Z(n666) );
  AND U750 ( .A(n669), .B(p_input[24]), .Z(n668) );
  AND U751 ( .A(p_input[224]), .B(p_input[124]), .Z(n669) );
  AND U752 ( .A(p_input[424]), .B(p_input[324]), .Z(n667) );
  AND U753 ( .A(n670), .B(n671), .Z(n665) );
  AND U754 ( .A(n672), .B(p_input[724]), .Z(n671) );
  AND U755 ( .A(p_input[624]), .B(p_input[524]), .Z(n672) );
  AND U756 ( .A(p_input[924]), .B(p_input[824]), .Z(n670) );
  AND U757 ( .A(n673), .B(n674), .Z(o[23]) );
  AND U758 ( .A(n675), .B(n676), .Z(n674) );
  AND U759 ( .A(n677), .B(p_input[23]), .Z(n676) );
  AND U760 ( .A(p_input[223]), .B(p_input[123]), .Z(n677) );
  AND U761 ( .A(p_input[423]), .B(p_input[323]), .Z(n675) );
  AND U762 ( .A(n678), .B(n679), .Z(n673) );
  AND U763 ( .A(n680), .B(p_input[723]), .Z(n679) );
  AND U764 ( .A(p_input[623]), .B(p_input[523]), .Z(n680) );
  AND U765 ( .A(p_input[923]), .B(p_input[823]), .Z(n678) );
  AND U766 ( .A(n681), .B(n682), .Z(o[22]) );
  AND U767 ( .A(n683), .B(n684), .Z(n682) );
  AND U768 ( .A(n685), .B(p_input[22]), .Z(n684) );
  AND U769 ( .A(p_input[222]), .B(p_input[122]), .Z(n685) );
  AND U770 ( .A(p_input[422]), .B(p_input[322]), .Z(n683) );
  AND U771 ( .A(n686), .B(n687), .Z(n681) );
  AND U772 ( .A(n688), .B(p_input[722]), .Z(n687) );
  AND U773 ( .A(p_input[622]), .B(p_input[522]), .Z(n688) );
  AND U774 ( .A(p_input[922]), .B(p_input[822]), .Z(n686) );
  AND U775 ( .A(n689), .B(n690), .Z(o[21]) );
  AND U776 ( .A(n691), .B(n692), .Z(n690) );
  AND U777 ( .A(n693), .B(p_input[221]), .Z(n692) );
  AND U778 ( .A(p_input[21]), .B(p_input[121]), .Z(n693) );
  AND U779 ( .A(p_input[421]), .B(p_input[321]), .Z(n691) );
  AND U780 ( .A(n694), .B(n695), .Z(n689) );
  AND U781 ( .A(n696), .B(p_input[721]), .Z(n695) );
  AND U782 ( .A(p_input[621]), .B(p_input[521]), .Z(n696) );
  AND U783 ( .A(p_input[921]), .B(p_input[821]), .Z(n694) );
  AND U784 ( .A(n697), .B(n698), .Z(o[20]) );
  AND U785 ( .A(n699), .B(n700), .Z(n698) );
  AND U786 ( .A(n701), .B(p_input[220]), .Z(n700) );
  AND U787 ( .A(p_input[20]), .B(p_input[120]), .Z(n701) );
  AND U788 ( .A(p_input[420]), .B(p_input[320]), .Z(n699) );
  AND U789 ( .A(n702), .B(n703), .Z(n697) );
  AND U790 ( .A(n704), .B(p_input[720]), .Z(n703) );
  AND U791 ( .A(p_input[620]), .B(p_input[520]), .Z(n704) );
  AND U792 ( .A(p_input[920]), .B(p_input[820]), .Z(n702) );
  AND U793 ( .A(n705), .B(n706), .Z(o[1]) );
  AND U794 ( .A(n707), .B(n708), .Z(n706) );
  AND U795 ( .A(n709), .B(p_input[201]), .Z(n708) );
  AND U796 ( .A(p_input[1]), .B(p_input[101]), .Z(n709) );
  AND U797 ( .A(p_input[401]), .B(p_input[301]), .Z(n707) );
  AND U798 ( .A(n710), .B(n711), .Z(n705) );
  AND U799 ( .A(n712), .B(p_input[701]), .Z(n711) );
  AND U800 ( .A(p_input[601]), .B(p_input[501]), .Z(n712) );
  AND U801 ( .A(p_input[901]), .B(p_input[801]), .Z(n710) );
  AND U802 ( .A(n713), .B(n714), .Z(o[19]) );
  AND U803 ( .A(n715), .B(n716), .Z(n714) );
  AND U804 ( .A(n717), .B(p_input[219]), .Z(n716) );
  AND U805 ( .A(p_input[19]), .B(p_input[119]), .Z(n717) );
  AND U806 ( .A(p_input[419]), .B(p_input[319]), .Z(n715) );
  AND U807 ( .A(n718), .B(n719), .Z(n713) );
  AND U808 ( .A(n720), .B(p_input[719]), .Z(n719) );
  AND U809 ( .A(p_input[619]), .B(p_input[519]), .Z(n720) );
  AND U810 ( .A(p_input[919]), .B(p_input[819]), .Z(n718) );
  AND U811 ( .A(n721), .B(n722), .Z(o[18]) );
  AND U812 ( .A(n723), .B(n724), .Z(n722) );
  AND U813 ( .A(n725), .B(p_input[218]), .Z(n724) );
  AND U814 ( .A(p_input[18]), .B(p_input[118]), .Z(n725) );
  AND U815 ( .A(p_input[418]), .B(p_input[318]), .Z(n723) );
  AND U816 ( .A(n726), .B(n727), .Z(n721) );
  AND U817 ( .A(n728), .B(p_input[718]), .Z(n727) );
  AND U818 ( .A(p_input[618]), .B(p_input[518]), .Z(n728) );
  AND U819 ( .A(p_input[918]), .B(p_input[818]), .Z(n726) );
  AND U820 ( .A(n729), .B(n730), .Z(o[17]) );
  AND U821 ( .A(n731), .B(n732), .Z(n730) );
  AND U822 ( .A(n733), .B(p_input[217]), .Z(n732) );
  AND U823 ( .A(p_input[17]), .B(p_input[117]), .Z(n733) );
  AND U824 ( .A(p_input[417]), .B(p_input[317]), .Z(n731) );
  AND U825 ( .A(n734), .B(n735), .Z(n729) );
  AND U826 ( .A(n736), .B(p_input[717]), .Z(n735) );
  AND U827 ( .A(p_input[617]), .B(p_input[517]), .Z(n736) );
  AND U828 ( .A(p_input[917]), .B(p_input[817]), .Z(n734) );
  AND U829 ( .A(n737), .B(n738), .Z(o[16]) );
  AND U830 ( .A(n739), .B(n740), .Z(n738) );
  AND U831 ( .A(n741), .B(p_input[216]), .Z(n740) );
  AND U832 ( .A(p_input[16]), .B(p_input[116]), .Z(n741) );
  AND U833 ( .A(p_input[416]), .B(p_input[316]), .Z(n739) );
  AND U834 ( .A(n742), .B(n743), .Z(n737) );
  AND U835 ( .A(n744), .B(p_input[716]), .Z(n743) );
  AND U836 ( .A(p_input[616]), .B(p_input[516]), .Z(n744) );
  AND U837 ( .A(p_input[916]), .B(p_input[816]), .Z(n742) );
  AND U838 ( .A(n745), .B(n746), .Z(o[15]) );
  AND U839 ( .A(n747), .B(n748), .Z(n746) );
  AND U840 ( .A(n749), .B(p_input[215]), .Z(n748) );
  AND U841 ( .A(p_input[15]), .B(p_input[115]), .Z(n749) );
  AND U842 ( .A(p_input[415]), .B(p_input[315]), .Z(n747) );
  AND U843 ( .A(n750), .B(n751), .Z(n745) );
  AND U844 ( .A(n752), .B(p_input[715]), .Z(n751) );
  AND U845 ( .A(p_input[615]), .B(p_input[515]), .Z(n752) );
  AND U846 ( .A(p_input[915]), .B(p_input[815]), .Z(n750) );
  AND U847 ( .A(n753), .B(n754), .Z(o[14]) );
  AND U848 ( .A(n755), .B(n756), .Z(n754) );
  AND U849 ( .A(n757), .B(p_input[214]), .Z(n756) );
  AND U850 ( .A(p_input[14]), .B(p_input[114]), .Z(n757) );
  AND U851 ( .A(p_input[414]), .B(p_input[314]), .Z(n755) );
  AND U852 ( .A(n758), .B(n759), .Z(n753) );
  AND U853 ( .A(n760), .B(p_input[714]), .Z(n759) );
  AND U854 ( .A(p_input[614]), .B(p_input[514]), .Z(n760) );
  AND U855 ( .A(p_input[914]), .B(p_input[814]), .Z(n758) );
  AND U856 ( .A(n761), .B(n762), .Z(o[13]) );
  AND U857 ( .A(n763), .B(n764), .Z(n762) );
  AND U858 ( .A(n765), .B(p_input[213]), .Z(n764) );
  AND U859 ( .A(p_input[13]), .B(p_input[113]), .Z(n765) );
  AND U860 ( .A(p_input[413]), .B(p_input[313]), .Z(n763) );
  AND U861 ( .A(n766), .B(n767), .Z(n761) );
  AND U862 ( .A(n768), .B(p_input[713]), .Z(n767) );
  AND U863 ( .A(p_input[613]), .B(p_input[513]), .Z(n768) );
  AND U864 ( .A(p_input[913]), .B(p_input[813]), .Z(n766) );
  AND U865 ( .A(n769), .B(n770), .Z(o[12]) );
  AND U866 ( .A(n771), .B(n772), .Z(n770) );
  AND U867 ( .A(n773), .B(p_input[212]), .Z(n772) );
  AND U868 ( .A(p_input[12]), .B(p_input[112]), .Z(n773) );
  AND U869 ( .A(p_input[412]), .B(p_input[312]), .Z(n771) );
  AND U870 ( .A(n774), .B(n775), .Z(n769) );
  AND U871 ( .A(n776), .B(p_input[712]), .Z(n775) );
  AND U872 ( .A(p_input[612]), .B(p_input[512]), .Z(n776) );
  AND U873 ( .A(p_input[912]), .B(p_input[812]), .Z(n774) );
  AND U874 ( .A(n777), .B(n778), .Z(o[11]) );
  AND U875 ( .A(n779), .B(n780), .Z(n778) );
  AND U876 ( .A(n781), .B(p_input[211]), .Z(n780) );
  AND U877 ( .A(p_input[11]), .B(p_input[111]), .Z(n781) );
  AND U878 ( .A(p_input[411]), .B(p_input[311]), .Z(n779) );
  AND U879 ( .A(n782), .B(n783), .Z(n777) );
  AND U880 ( .A(n784), .B(p_input[711]), .Z(n783) );
  AND U881 ( .A(p_input[611]), .B(p_input[511]), .Z(n784) );
  AND U882 ( .A(p_input[911]), .B(p_input[811]), .Z(n782) );
  AND U883 ( .A(n785), .B(n786), .Z(o[10]) );
  AND U884 ( .A(n787), .B(n788), .Z(n786) );
  AND U885 ( .A(n789), .B(p_input[210]), .Z(n788) );
  AND U886 ( .A(p_input[110]), .B(p_input[10]), .Z(n789) );
  AND U887 ( .A(p_input[410]), .B(p_input[310]), .Z(n787) );
  AND U888 ( .A(n790), .B(n791), .Z(n785) );
  AND U889 ( .A(n792), .B(p_input[710]), .Z(n791) );
  AND U890 ( .A(p_input[610]), .B(p_input[510]), .Z(n792) );
  AND U891 ( .A(p_input[910]), .B(p_input[810]), .Z(n790) );
  AND U892 ( .A(n793), .B(n794), .Z(o[0]) );
  AND U893 ( .A(n795), .B(n796), .Z(n794) );
  AND U894 ( .A(n797), .B(p_input[200]), .Z(n796) );
  AND U895 ( .A(p_input[100]), .B(p_input[0]), .Z(n797) );
  AND U896 ( .A(p_input[400]), .B(p_input[300]), .Z(n795) );
  AND U897 ( .A(n798), .B(n799), .Z(n793) );
  AND U898 ( .A(n800), .B(p_input[700]), .Z(n799) );
  AND U899 ( .A(p_input[600]), .B(p_input[500]), .Z(n800) );
  AND U900 ( .A(p_input[900]), .B(p_input[800]), .Z(n798) );
endmodule

