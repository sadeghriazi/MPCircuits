
module knn_comb_BMR_W16_K1_N4 ( p_input, o );
  input [79:0] p_input;
  output [15:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529;
  assign \knn_comb_/min_val_out[0][0]  = p_input[48];
  assign \knn_comb_/min_val_out[0][1]  = p_input[49];
  assign \knn_comb_/min_val_out[0][2]  = p_input[50];
  assign \knn_comb_/min_val_out[0][3]  = p_input[51];
  assign \knn_comb_/min_val_out[0][4]  = p_input[52];
  assign \knn_comb_/min_val_out[0][5]  = p_input[53];
  assign \knn_comb_/min_val_out[0][6]  = p_input[54];
  assign \knn_comb_/min_val_out[0][7]  = p_input[55];
  assign \knn_comb_/min_val_out[0][8]  = p_input[56];
  assign \knn_comb_/min_val_out[0][9]  = p_input[57];
  assign \knn_comb_/min_val_out[0][10]  = p_input[58];
  assign \knn_comb_/min_val_out[0][11]  = p_input[59];
  assign \knn_comb_/min_val_out[0][12]  = p_input[60];
  assign \knn_comb_/min_val_out[0][13]  = p_input[61];
  assign \knn_comb_/min_val_out[0][14]  = p_input[62];
  assign \knn_comb_/min_val_out[0][15]  = p_input[63];

  XNOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(n3), .B(n4), .Z(n1) );
  XNOR U3 ( .A(p_input[9]), .B(n2), .Z(n4) );
  XOR U4 ( .A(n5), .B(n6), .Z(n2) );
  AND U5 ( .A(n7), .B(n8), .Z(n6) );
  XNOR U6 ( .A(p_input[25]), .B(n5), .Z(n8) );
  XNOR U7 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n9), .Z(n5) );
  AND U8 ( .A(n10), .B(n11), .Z(n9) );
  XOR U9 ( .A(p_input[41]), .B(\knn_comb_/min_val_out[0][9] ), .Z(n11) );
  XNOR U10 ( .A(n12), .B(n13), .Z(o[8]) );
  AND U11 ( .A(n3), .B(n14), .Z(n12) );
  XNOR U12 ( .A(p_input[8]), .B(n13), .Z(n14) );
  XOR U13 ( .A(n15), .B(n16), .Z(n13) );
  AND U14 ( .A(n7), .B(n17), .Z(n16) );
  XNOR U15 ( .A(p_input[24]), .B(n15), .Z(n17) );
  XNOR U16 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n18), .Z(n15) );
  AND U17 ( .A(n10), .B(n19), .Z(n18) );
  XOR U18 ( .A(p_input[40]), .B(\knn_comb_/min_val_out[0][8] ), .Z(n19) );
  XNOR U19 ( .A(n20), .B(n21), .Z(o[7]) );
  AND U20 ( .A(n3), .B(n22), .Z(n20) );
  XNOR U21 ( .A(p_input[7]), .B(n21), .Z(n22) );
  XOR U22 ( .A(n23), .B(n24), .Z(n21) );
  AND U23 ( .A(n7), .B(n25), .Z(n24) );
  XNOR U24 ( .A(p_input[23]), .B(n23), .Z(n25) );
  XNOR U25 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n26), .Z(n23) );
  AND U26 ( .A(n10), .B(n27), .Z(n26) );
  XNOR U27 ( .A(p_input[39]), .B(n28), .Z(n27) );
  IV U28 ( .A(\knn_comb_/min_val_out[0][7] ), .Z(n28) );
  XNOR U29 ( .A(n29), .B(n30), .Z(o[6]) );
  AND U30 ( .A(n3), .B(n31), .Z(n29) );
  XNOR U31 ( .A(p_input[6]), .B(n30), .Z(n31) );
  XOR U32 ( .A(n32), .B(n33), .Z(n30) );
  AND U33 ( .A(n7), .B(n34), .Z(n33) );
  XNOR U34 ( .A(p_input[22]), .B(n32), .Z(n34) );
  XNOR U35 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n35), .Z(n32) );
  AND U36 ( .A(n10), .B(n36), .Z(n35) );
  XOR U37 ( .A(p_input[38]), .B(\knn_comb_/min_val_out[0][6] ), .Z(n36) );
  XNOR U38 ( .A(n37), .B(n38), .Z(o[5]) );
  AND U39 ( .A(n3), .B(n39), .Z(n37) );
  XNOR U40 ( .A(p_input[5]), .B(n38), .Z(n39) );
  XOR U41 ( .A(n40), .B(n41), .Z(n38) );
  AND U42 ( .A(n7), .B(n42), .Z(n41) );
  XNOR U43 ( .A(p_input[21]), .B(n40), .Z(n42) );
  XNOR U44 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n43), .Z(n40) );
  AND U45 ( .A(n10), .B(n44), .Z(n43) );
  XOR U46 ( .A(p_input[37]), .B(\knn_comb_/min_val_out[0][5] ), .Z(n44) );
  XNOR U47 ( .A(n45), .B(n46), .Z(o[4]) );
  AND U48 ( .A(n3), .B(n47), .Z(n45) );
  XNOR U49 ( .A(p_input[4]), .B(n46), .Z(n47) );
  XOR U50 ( .A(n48), .B(n49), .Z(n46) );
  AND U51 ( .A(n7), .B(n50), .Z(n49) );
  XNOR U52 ( .A(p_input[20]), .B(n48), .Z(n50) );
  XNOR U53 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n51), .Z(n48) );
  AND U54 ( .A(n10), .B(n52), .Z(n51) );
  XNOR U55 ( .A(p_input[36]), .B(n53), .Z(n52) );
  IV U56 ( .A(\knn_comb_/min_val_out[0][4] ), .Z(n53) );
  XNOR U57 ( .A(n54), .B(n55), .Z(o[3]) );
  AND U58 ( .A(n3), .B(n56), .Z(n54) );
  XNOR U59 ( .A(p_input[3]), .B(n55), .Z(n56) );
  XOR U60 ( .A(n57), .B(n58), .Z(n55) );
  AND U61 ( .A(n7), .B(n59), .Z(n58) );
  XNOR U62 ( .A(p_input[19]), .B(n57), .Z(n59) );
  XNOR U63 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n60), .Z(n57) );
  AND U64 ( .A(n10), .B(n61), .Z(n60) );
  XOR U65 ( .A(p_input[35]), .B(\knn_comb_/min_val_out[0][3] ), .Z(n61) );
  XNOR U66 ( .A(n62), .B(n63), .Z(o[2]) );
  AND U67 ( .A(n3), .B(n64), .Z(n62) );
  XNOR U68 ( .A(p_input[2]), .B(n63), .Z(n64) );
  XOR U69 ( .A(n65), .B(n66), .Z(n63) );
  AND U70 ( .A(n7), .B(n67), .Z(n66) );
  XNOR U71 ( .A(p_input[18]), .B(n65), .Z(n67) );
  XNOR U72 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n68), .Z(n65) );
  AND U73 ( .A(n10), .B(n69), .Z(n68) );
  XOR U74 ( .A(p_input[34]), .B(\knn_comb_/min_val_out[0][2] ), .Z(n69) );
  XNOR U75 ( .A(n70), .B(n71), .Z(o[1]) );
  AND U76 ( .A(n3), .B(n72), .Z(n70) );
  XNOR U77 ( .A(p_input[1]), .B(n71), .Z(n72) );
  XOR U78 ( .A(n73), .B(n74), .Z(n71) );
  AND U79 ( .A(n7), .B(n75), .Z(n74) );
  XNOR U80 ( .A(p_input[17]), .B(n73), .Z(n75) );
  XNOR U81 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n76), .Z(n73) );
  AND U82 ( .A(n10), .B(n77), .Z(n76) );
  XOR U83 ( .A(p_input[33]), .B(\knn_comb_/min_val_out[0][1] ), .Z(n77) );
  XNOR U84 ( .A(n78), .B(n79), .Z(o[15]) );
  AND U85 ( .A(n3), .B(n80), .Z(n78) );
  XNOR U86 ( .A(p_input[15]), .B(n79), .Z(n80) );
  XOR U87 ( .A(n81), .B(n82), .Z(n79) );
  AND U88 ( .A(n7), .B(n83), .Z(n82) );
  XNOR U89 ( .A(p_input[31]), .B(n81), .Z(n83) );
  XNOR U90 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n84), .Z(n81) );
  AND U91 ( .A(n10), .B(n85), .Z(n84) );
  XOR U92 ( .A(p_input[47]), .B(\knn_comb_/min_val_out[0][15] ), .Z(n85) );
  XNOR U93 ( .A(n86), .B(n87), .Z(o[14]) );
  AND U94 ( .A(n3), .B(n88), .Z(n86) );
  XNOR U95 ( .A(p_input[14]), .B(n87), .Z(n88) );
  XOR U96 ( .A(n89), .B(n90), .Z(n87) );
  AND U97 ( .A(n7), .B(n91), .Z(n90) );
  XNOR U98 ( .A(p_input[30]), .B(n89), .Z(n91) );
  XNOR U99 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n92), .Z(n89) );
  AND U100 ( .A(n10), .B(n93), .Z(n92) );
  XNOR U101 ( .A(p_input[46]), .B(n94), .Z(n93) );
  IV U102 ( .A(\knn_comb_/min_val_out[0][14] ), .Z(n94) );
  XNOR U103 ( .A(n95), .B(n96), .Z(o[13]) );
  AND U104 ( .A(n3), .B(n97), .Z(n95) );
  XNOR U105 ( .A(p_input[13]), .B(n96), .Z(n97) );
  XOR U106 ( .A(n98), .B(n99), .Z(n96) );
  AND U107 ( .A(n7), .B(n100), .Z(n99) );
  XNOR U108 ( .A(p_input[29]), .B(n98), .Z(n100) );
  XNOR U109 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n101), .Z(n98) );
  AND U110 ( .A(n10), .B(n102), .Z(n101) );
  XOR U111 ( .A(p_input[45]), .B(\knn_comb_/min_val_out[0][13] ), .Z(n102) );
  XNOR U112 ( .A(n103), .B(n104), .Z(o[12]) );
  AND U113 ( .A(n3), .B(n105), .Z(n103) );
  XNOR U114 ( .A(p_input[12]), .B(n104), .Z(n105) );
  XOR U115 ( .A(n106), .B(n107), .Z(n104) );
  AND U116 ( .A(n7), .B(n108), .Z(n107) );
  XNOR U117 ( .A(p_input[28]), .B(n106), .Z(n108) );
  XNOR U118 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n109), .Z(n106) );
  AND U119 ( .A(n10), .B(n110), .Z(n109) );
  XOR U120 ( .A(p_input[44]), .B(\knn_comb_/min_val_out[0][12] ), .Z(n110) );
  XNOR U121 ( .A(n111), .B(n112), .Z(o[11]) );
  AND U122 ( .A(n3), .B(n113), .Z(n111) );
  XNOR U123 ( .A(p_input[11]), .B(n112), .Z(n113) );
  XOR U124 ( .A(n114), .B(n115), .Z(n112) );
  AND U125 ( .A(n7), .B(n116), .Z(n115) );
  XNOR U126 ( .A(p_input[27]), .B(n114), .Z(n116) );
  XNOR U127 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n117), .Z(n114) );
  AND U128 ( .A(n10), .B(n118), .Z(n117) );
  XNOR U129 ( .A(p_input[43]), .B(n119), .Z(n118) );
  IV U130 ( .A(\knn_comb_/min_val_out[0][11] ), .Z(n119) );
  XNOR U131 ( .A(n120), .B(n121), .Z(o[10]) );
  AND U132 ( .A(n3), .B(n122), .Z(n120) );
  XNOR U133 ( .A(p_input[10]), .B(n121), .Z(n122) );
  XOR U134 ( .A(n123), .B(n124), .Z(n121) );
  AND U135 ( .A(n7), .B(n125), .Z(n124) );
  XNOR U136 ( .A(p_input[26]), .B(n123), .Z(n125) );
  XNOR U137 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n126), .Z(n123) );
  AND U138 ( .A(n10), .B(n127), .Z(n126) );
  XOR U139 ( .A(p_input[42]), .B(\knn_comb_/min_val_out[0][10] ), .Z(n127) );
  XNOR U140 ( .A(n128), .B(n129), .Z(o[0]) );
  AND U141 ( .A(n3), .B(n130), .Z(n128) );
  XNOR U142 ( .A(p_input[0]), .B(n129), .Z(n130) );
  XOR U143 ( .A(n131), .B(n132), .Z(n129) );
  AND U144 ( .A(n7), .B(n133), .Z(n132) );
  XNOR U145 ( .A(p_input[16]), .B(n131), .Z(n133) );
  XNOR U146 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n134), .Z(n131) );
  AND U147 ( .A(n10), .B(n135), .Z(n134) );
  XOR U148 ( .A(p_input[32]), .B(\knn_comb_/min_val_out[0][0] ), .Z(n135) );
  XOR U149 ( .A(n136), .B(n137), .Z(n3) );
  MUX U150 ( .IN0(n138), .IN1(n139), .SEL(n137), .F(n136) );
  XOR U151 ( .A(n140), .B(n141), .Z(n137) );
  AND U152 ( .A(n142), .B(n143), .Z(n141) );
  XOR U153 ( .A(n140), .B(n144), .Z(n143) );
  XNOR U154 ( .A(n145), .B(n140), .Z(n142) );
  XOR U155 ( .A(n146), .B(n147), .Z(n145) );
  AND U156 ( .A(n7), .B(n148), .Z(n147) );
  XOR U157 ( .A(n149), .B(n146), .Z(n148) );
  XOR U158 ( .A(n150), .B(n151), .Z(n140) );
  AND U159 ( .A(n152), .B(n153), .Z(n151) );
  XOR U160 ( .A(n150), .B(n154), .Z(n153) );
  XNOR U161 ( .A(n155), .B(n150), .Z(n152) );
  XOR U162 ( .A(n156), .B(n157), .Z(n155) );
  AND U163 ( .A(n7), .B(n158), .Z(n157) );
  XOR U164 ( .A(n159), .B(n156), .Z(n158) );
  XOR U165 ( .A(n160), .B(n161), .Z(n150) );
  AND U166 ( .A(n162), .B(n163), .Z(n161) );
  XNOR U167 ( .A(n164), .B(n165), .Z(n163) );
  XOR U168 ( .A(n166), .B(n167), .Z(n162) );
  XNOR U169 ( .A(n160), .B(n168), .Z(n167) );
  AND U170 ( .A(n7), .B(n169), .Z(n168) );
  XOR U171 ( .A(n170), .B(n166), .Z(n169) );
  IV U172 ( .A(n164), .Z(n160) );
  AND U173 ( .A(n171), .B(n172), .Z(n164) );
  XNOR U174 ( .A(n173), .B(n174), .Z(n171) );
  AND U175 ( .A(n7), .B(n175), .Z(n174) );
  XOR U176 ( .A(n176), .B(n177), .Z(n175) );
  IV U177 ( .A(n173), .Z(n177) );
  XOR U178 ( .A(n178), .B(n179), .Z(n7) );
  MUX U179 ( .IN0(n180), .IN1(n181), .SEL(n178), .F(n179) );
  XOR U180 ( .A(n182), .B(n183), .Z(n178) );
  AND U181 ( .A(n184), .B(n185), .Z(n183) );
  XOR U182 ( .A(n182), .B(n149), .Z(n185) );
  XNOR U183 ( .A(n146), .B(n182), .Z(n184) );
  XOR U184 ( .A(n186), .B(n187), .Z(n146) );
  AND U185 ( .A(n10), .B(n188), .Z(n187) );
  XOR U186 ( .A(n189), .B(n186), .Z(n188) );
  XOR U187 ( .A(n190), .B(n191), .Z(n182) );
  AND U188 ( .A(n192), .B(n193), .Z(n191) );
  XOR U189 ( .A(n190), .B(n159), .Z(n193) );
  XNOR U190 ( .A(n156), .B(n190), .Z(n192) );
  XOR U191 ( .A(n194), .B(n195), .Z(n156) );
  AND U192 ( .A(n10), .B(n196), .Z(n195) );
  XOR U193 ( .A(n197), .B(n194), .Z(n196) );
  XOR U194 ( .A(n198), .B(n199), .Z(n190) );
  AND U195 ( .A(n200), .B(n201), .Z(n199) );
  XNOR U196 ( .A(n202), .B(n170), .Z(n201) );
  XNOR U197 ( .A(n166), .B(n198), .Z(n200) );
  XOR U198 ( .A(n203), .B(n204), .Z(n166) );
  AND U199 ( .A(n10), .B(n205), .Z(n204) );
  XOR U200 ( .A(n206), .B(n203), .Z(n205) );
  IV U201 ( .A(n202), .Z(n198) );
  NOR U202 ( .A(n173), .B(n176), .Z(n202) );
  XOR U203 ( .A(n207), .B(n208), .Z(n173) );
  AND U204 ( .A(n10), .B(n209), .Z(n208) );
  XNOR U205 ( .A(n210), .B(n207), .Z(n209) );
  XOR U206 ( .A(n211), .B(n212), .Z(n10) );
  MUX U207 ( .IN0(n213), .IN1(n214), .SEL(n211), .F(n212) );
  XOR U208 ( .A(n215), .B(n216), .Z(n211) );
  AND U209 ( .A(n217), .B(n218), .Z(n216) );
  XOR U210 ( .A(n215), .B(n189), .Z(n218) );
  XOR U211 ( .A(n219), .B(n215), .Z(n217) );
  IV U212 ( .A(n186), .Z(n219) );
  XOR U213 ( .A(n220), .B(n221), .Z(n215) );
  AND U214 ( .A(n222), .B(n223), .Z(n221) );
  XOR U215 ( .A(n220), .B(n197), .Z(n223) );
  XNOR U216 ( .A(n194), .B(n220), .Z(n222) );
  XOR U217 ( .A(n224), .B(n225), .Z(n220) );
  AND U218 ( .A(n226), .B(n227), .Z(n225) );
  XNOR U219 ( .A(n228), .B(n206), .Z(n227) );
  XNOR U220 ( .A(n203), .B(n224), .Z(n226) );
  IV U221 ( .A(n228), .Z(n224) );
  NOR U222 ( .A(n207), .B(n210), .Z(n228) );
  AND U223 ( .A(n144), .B(n229), .Z(n139) );
  XOR U224 ( .A(n230), .B(n231), .Z(n144) );
  XOR U225 ( .A(n232), .B(n229), .Z(n231) );
  AND U226 ( .A(n154), .B(n233), .Z(n229) );
  XNOR U227 ( .A(n234), .B(n235), .Z(n154) );
  XOR U228 ( .A(n236), .B(n233), .Z(n234) );
  AND U229 ( .A(n165), .B(n237), .Z(n233) );
  XNOR U230 ( .A(n238), .B(n239), .Z(n165) );
  XOR U231 ( .A(n240), .B(n237), .Z(n238) );
  NOR U232 ( .A(n172), .B(n241), .Z(n237) );
  XOR U233 ( .A(n242), .B(n241), .Z(n172) );
  XNOR U234 ( .A(p_input[0]), .B(p_input[64]), .Z(n241) );
  XOR U235 ( .A(n243), .B(n244), .Z(n242) );
  NOR U236 ( .A(n245), .B(n235), .Z(n232) );
  XNOR U237 ( .A(n246), .B(n230), .Z(n235) );
  XOR U238 ( .A(n247), .B(n248), .Z(n246) );
  AND U239 ( .A(n249), .B(n250), .Z(n248) );
  XOR U240 ( .A(n247), .B(n251), .Z(n249) );
  XNOR U241 ( .A(n236), .B(n230), .Z(n245) );
  XOR U242 ( .A(n252), .B(n253), .Z(n236) );
  AND U243 ( .A(n254), .B(n255), .Z(n253) );
  XOR U244 ( .A(n252), .B(n256), .Z(n254) );
  XOR U245 ( .A(n257), .B(n258), .Z(n230) );
  NOR U246 ( .A(n259), .B(n239), .Z(n258) );
  XNOR U247 ( .A(n260), .B(n251), .Z(n239) );
  XOR U248 ( .A(n261), .B(n262), .Z(n251) );
  AND U249 ( .A(n263), .B(n264), .Z(n262) );
  XOR U250 ( .A(n261), .B(n265), .Z(n263) );
  XOR U251 ( .A(n250), .B(n257), .Z(n260) );
  XOR U252 ( .A(n266), .B(n247), .Z(n250) );
  XOR U253 ( .A(n267), .B(n268), .Z(n247) );
  AND U254 ( .A(n269), .B(n270), .Z(n268) );
  XOR U255 ( .A(n267), .B(n271), .Z(n269) );
  XOR U256 ( .A(n272), .B(n273), .Z(n266) );
  AND U257 ( .A(n274), .B(n275), .Z(n273) );
  XOR U258 ( .A(n272), .B(n276), .Z(n274) );
  XNOR U259 ( .A(n240), .B(n257), .Z(n259) );
  XOR U260 ( .A(n256), .B(n255), .Z(n240) );
  XOR U261 ( .A(n277), .B(n252), .Z(n255) );
  XOR U262 ( .A(n278), .B(n279), .Z(n252) );
  AND U263 ( .A(n280), .B(n281), .Z(n279) );
  XOR U264 ( .A(n278), .B(n282), .Z(n280) );
  XOR U265 ( .A(n283), .B(n284), .Z(n277) );
  AND U266 ( .A(n285), .B(n286), .Z(n284) );
  XOR U267 ( .A(n283), .B(n287), .Z(n285) );
  XNOR U268 ( .A(n288), .B(n289), .Z(n256) );
  AND U269 ( .A(n290), .B(n291), .Z(n289) );
  XNOR U270 ( .A(n288), .B(n292), .Z(n290) );
  XNOR U271 ( .A(n293), .B(n294), .Z(n257) );
  AND U272 ( .A(n295), .B(n244), .Z(n294) );
  XOR U273 ( .A(n296), .B(n271), .Z(n244) );
  XOR U274 ( .A(n265), .B(n264), .Z(n271) );
  XOR U275 ( .A(n297), .B(n261), .Z(n264) );
  XNOR U276 ( .A(p_input[10]), .B(p_input[74]), .Z(n261) );
  XNOR U277 ( .A(p_input[11]), .B(p_input[75]), .Z(n297) );
  XNOR U278 ( .A(p_input[12]), .B(p_input[76]), .Z(n265) );
  XNOR U279 ( .A(n270), .B(n293), .Z(n296) );
  XOR U280 ( .A(n298), .B(n276), .Z(n270) );
  XNOR U281 ( .A(p_input[15]), .B(p_input[79]), .Z(n276) );
  XOR U282 ( .A(n267), .B(n275), .Z(n298) );
  XOR U283 ( .A(n299), .B(n272), .Z(n275) );
  XNOR U284 ( .A(p_input[13]), .B(p_input[77]), .Z(n272) );
  XNOR U285 ( .A(p_input[14]), .B(p_input[78]), .Z(n299) );
  XNOR U286 ( .A(p_input[73]), .B(p_input[9]), .Z(n267) );
  XNOR U287 ( .A(n293), .B(n243), .Z(n295) );
  XOR U288 ( .A(n282), .B(n281), .Z(n243) );
  XOR U289 ( .A(n300), .B(n287), .Z(n281) );
  XNOR U290 ( .A(p_input[72]), .B(p_input[8]), .Z(n287) );
  XOR U291 ( .A(n278), .B(n286), .Z(n300) );
  XOR U292 ( .A(n301), .B(n283), .Z(n286) );
  XNOR U293 ( .A(p_input[6]), .B(p_input[70]), .Z(n283) );
  XNOR U294 ( .A(p_input[71]), .B(p_input[7]), .Z(n301) );
  XNOR U295 ( .A(p_input[2]), .B(p_input[66]), .Z(n278) );
  XOR U296 ( .A(n292), .B(n291), .Z(n282) );
  XNOR U297 ( .A(n302), .B(n288), .Z(n291) );
  XOR U298 ( .A(p_input[3]), .B(p_input[67]), .Z(n288) );
  XNOR U299 ( .A(p_input[4]), .B(p_input[68]), .Z(n302) );
  XNOR U300 ( .A(p_input[5]), .B(p_input[69]), .Z(n292) );
  XOR U301 ( .A(p_input[1]), .B(p_input[65]), .Z(n293) );
  AND U302 ( .A(n181), .B(n180), .Z(n138) );
  AND U303 ( .A(n214), .B(n213), .Z(n180) );
  AND U304 ( .A(n186), .B(n303), .Z(n213) );
  XOR U305 ( .A(n304), .B(n305), .Z(n186) );
  XOR U306 ( .A(n306), .B(n303), .Z(n305) );
  AND U307 ( .A(n194), .B(n307), .Z(n303) );
  XNOR U308 ( .A(n308), .B(n309), .Z(n194) );
  XNOR U309 ( .A(n310), .B(n307), .Z(n308) );
  AND U310 ( .A(n203), .B(n311), .Z(n307) );
  XNOR U311 ( .A(n312), .B(n313), .Z(n203) );
  XNOR U312 ( .A(n314), .B(n311), .Z(n312) );
  NOR U313 ( .A(n207), .B(n315), .Z(n311) );
  XNOR U314 ( .A(n316), .B(n317), .Z(n207) );
  XOR U315 ( .A(n318), .B(n315), .Z(n316) );
  XNOR U316 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[64]), .Z(n315) );
  AND U317 ( .A(n319), .B(n310), .Z(n306) );
  XOR U318 ( .A(n320), .B(n304), .Z(n310) );
  XOR U319 ( .A(n321), .B(n322), .Z(n320) );
  AND U320 ( .A(n323), .B(n324), .Z(n322) );
  XOR U321 ( .A(n321), .B(n325), .Z(n323) );
  XOR U322 ( .A(n304), .B(n309), .Z(n319) );
  XOR U323 ( .A(n326), .B(n327), .Z(n309) );
  AND U324 ( .A(n328), .B(n329), .Z(n327) );
  XOR U325 ( .A(n326), .B(n330), .Z(n328) );
  XOR U326 ( .A(n331), .B(n332), .Z(n304) );
  AND U327 ( .A(n333), .B(n314), .Z(n332) );
  XOR U328 ( .A(n334), .B(n325), .Z(n314) );
  XOR U329 ( .A(n335), .B(n336), .Z(n325) );
  AND U330 ( .A(n337), .B(n338), .Z(n336) );
  XOR U331 ( .A(n335), .B(n339), .Z(n337) );
  XOR U332 ( .A(n324), .B(n331), .Z(n334) );
  XOR U333 ( .A(n340), .B(n321), .Z(n324) );
  XOR U334 ( .A(n341), .B(n342), .Z(n321) );
  AND U335 ( .A(n343), .B(n344), .Z(n342) );
  XOR U336 ( .A(n341), .B(n345), .Z(n343) );
  XOR U337 ( .A(n346), .B(n347), .Z(n340) );
  AND U338 ( .A(n348), .B(n349), .Z(n347) );
  XOR U339 ( .A(n346), .B(n350), .Z(n348) );
  XOR U340 ( .A(n331), .B(n313), .Z(n333) );
  XOR U341 ( .A(n330), .B(n329), .Z(n313) );
  XOR U342 ( .A(n351), .B(n326), .Z(n329) );
  XOR U343 ( .A(n352), .B(n353), .Z(n326) );
  AND U344 ( .A(n354), .B(n355), .Z(n353) );
  XOR U345 ( .A(n352), .B(n356), .Z(n354) );
  XOR U346 ( .A(n357), .B(n358), .Z(n351) );
  AND U347 ( .A(n359), .B(n360), .Z(n358) );
  XOR U348 ( .A(n357), .B(n361), .Z(n359) );
  XOR U349 ( .A(n362), .B(n363), .Z(n330) );
  AND U350 ( .A(n364), .B(n365), .Z(n363) );
  XOR U351 ( .A(n362), .B(n366), .Z(n364) );
  XOR U352 ( .A(n367), .B(n368), .Z(n331) );
  AND U353 ( .A(n369), .B(n318), .Z(n368) );
  XOR U354 ( .A(n370), .B(n345), .Z(n318) );
  XOR U355 ( .A(n339), .B(n338), .Z(n345) );
  XOR U356 ( .A(n371), .B(n335), .Z(n338) );
  XOR U357 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n372), .Z(n335) );
  IV U358 ( .A(p_input[74]), .Z(n372) );
  XNOR U359 ( .A(\knn_comb_/min_val_out[0][11] ), .B(p_input[75]), .Z(n371) );
  XNOR U360 ( .A(\knn_comb_/min_val_out[0][12] ), .B(p_input[76]), .Z(n339) );
  XOR U361 ( .A(n344), .B(n367), .Z(n370) );
  XOR U362 ( .A(n373), .B(n350), .Z(n344) );
  XNOR U363 ( .A(\knn_comb_/min_val_out[0][15] ), .B(p_input[79]), .Z(n350) );
  XOR U364 ( .A(n341), .B(n349), .Z(n373) );
  XOR U365 ( .A(n374), .B(n346), .Z(n349) );
  XOR U366 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n375), .Z(n346) );
  IV U367 ( .A(p_input[77]), .Z(n375) );
  XNOR U368 ( .A(\knn_comb_/min_val_out[0][14] ), .B(p_input[78]), .Z(n374) );
  XNOR U369 ( .A(\knn_comb_/min_val_out[0][9] ), .B(p_input[73]), .Z(n341) );
  XNOR U370 ( .A(n367), .B(n317), .Z(n369) );
  XNOR U371 ( .A(n356), .B(n355), .Z(n317) );
  XOR U372 ( .A(n376), .B(n361), .Z(n355) );
  XNOR U373 ( .A(\knn_comb_/min_val_out[0][8] ), .B(p_input[72]), .Z(n361) );
  XOR U374 ( .A(n352), .B(n360), .Z(n376) );
  XOR U375 ( .A(n377), .B(n357), .Z(n360) );
  XOR U376 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n378), .Z(n357) );
  IV U377 ( .A(p_input[70]), .Z(n378) );
  XNOR U378 ( .A(\knn_comb_/min_val_out[0][7] ), .B(p_input[71]), .Z(n377) );
  XNOR U379 ( .A(\knn_comb_/min_val_out[0][2] ), .B(p_input[66]), .Z(n352) );
  XOR U380 ( .A(n366), .B(n365), .Z(n356) );
  XOR U381 ( .A(n379), .B(n362), .Z(n365) );
  XOR U382 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n380), .Z(n362) );
  IV U383 ( .A(p_input[67]), .Z(n380) );
  XNOR U384 ( .A(\knn_comb_/min_val_out[0][4] ), .B(p_input[68]), .Z(n379) );
  XNOR U385 ( .A(\knn_comb_/min_val_out[0][5] ), .B(p_input[69]), .Z(n366) );
  XOR U386 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n381), .Z(n367) );
  IV U387 ( .A(p_input[65]), .Z(n381) );
  AND U388 ( .A(n189), .B(n382), .Z(n214) );
  XOR U389 ( .A(n383), .B(n384), .Z(n189) );
  XOR U390 ( .A(n385), .B(n382), .Z(n384) );
  AND U391 ( .A(n197), .B(n386), .Z(n382) );
  XNOR U392 ( .A(n387), .B(n388), .Z(n197) );
  XOR U393 ( .A(n389), .B(n386), .Z(n387) );
  AND U394 ( .A(n206), .B(n390), .Z(n386) );
  XNOR U395 ( .A(n391), .B(n392), .Z(n206) );
  XOR U396 ( .A(n393), .B(n390), .Z(n391) );
  AND U397 ( .A(n210), .B(n394), .Z(n390) );
  XOR U398 ( .A(n395), .B(n394), .Z(n210) );
  XOR U399 ( .A(p_input[32]), .B(p_input[64]), .Z(n394) );
  XOR U400 ( .A(n396), .B(n397), .Z(n395) );
  NOR U401 ( .A(n398), .B(n388), .Z(n385) );
  XNOR U402 ( .A(n399), .B(n383), .Z(n388) );
  XOR U403 ( .A(n400), .B(n401), .Z(n399) );
  AND U404 ( .A(n402), .B(n403), .Z(n401) );
  XOR U405 ( .A(n400), .B(n404), .Z(n402) );
  XNOR U406 ( .A(n389), .B(n383), .Z(n398) );
  XOR U407 ( .A(n405), .B(n406), .Z(n389) );
  AND U408 ( .A(n407), .B(n408), .Z(n406) );
  XOR U409 ( .A(n405), .B(n409), .Z(n407) );
  XOR U410 ( .A(n410), .B(n411), .Z(n383) );
  NOR U411 ( .A(n412), .B(n392), .Z(n411) );
  XNOR U412 ( .A(n413), .B(n404), .Z(n392) );
  XOR U413 ( .A(n414), .B(n415), .Z(n404) );
  AND U414 ( .A(n416), .B(n417), .Z(n415) );
  XOR U415 ( .A(n414), .B(n418), .Z(n416) );
  XOR U416 ( .A(n403), .B(n410), .Z(n413) );
  XOR U417 ( .A(n419), .B(n400), .Z(n403) );
  XOR U418 ( .A(n420), .B(n421), .Z(n400) );
  AND U419 ( .A(n422), .B(n423), .Z(n421) );
  XOR U420 ( .A(n420), .B(n424), .Z(n422) );
  XOR U421 ( .A(n425), .B(n426), .Z(n419) );
  AND U422 ( .A(n427), .B(n428), .Z(n426) );
  XOR U423 ( .A(n425), .B(n429), .Z(n427) );
  XNOR U424 ( .A(n393), .B(n410), .Z(n412) );
  XOR U425 ( .A(n409), .B(n408), .Z(n393) );
  XOR U426 ( .A(n430), .B(n405), .Z(n408) );
  XOR U427 ( .A(n431), .B(n432), .Z(n405) );
  AND U428 ( .A(n433), .B(n434), .Z(n432) );
  XOR U429 ( .A(n431), .B(n435), .Z(n433) );
  XOR U430 ( .A(n436), .B(n437), .Z(n430) );
  AND U431 ( .A(n438), .B(n439), .Z(n437) );
  XOR U432 ( .A(n436), .B(n440), .Z(n438) );
  XNOR U433 ( .A(n441), .B(n442), .Z(n409) );
  AND U434 ( .A(n443), .B(n444), .Z(n442) );
  XNOR U435 ( .A(n441), .B(n445), .Z(n443) );
  XNOR U436 ( .A(n446), .B(n447), .Z(n410) );
  AND U437 ( .A(n448), .B(n397), .Z(n447) );
  XOR U438 ( .A(n449), .B(n424), .Z(n397) );
  XOR U439 ( .A(n418), .B(n417), .Z(n424) );
  XOR U440 ( .A(n450), .B(n414), .Z(n417) );
  XNOR U441 ( .A(p_input[42]), .B(p_input[74]), .Z(n414) );
  XNOR U442 ( .A(p_input[43]), .B(p_input[75]), .Z(n450) );
  XNOR U443 ( .A(p_input[44]), .B(p_input[76]), .Z(n418) );
  XNOR U444 ( .A(n423), .B(n446), .Z(n449) );
  XOR U445 ( .A(n451), .B(n429), .Z(n423) );
  XNOR U446 ( .A(p_input[47]), .B(p_input[79]), .Z(n429) );
  XOR U447 ( .A(n420), .B(n428), .Z(n451) );
  XOR U448 ( .A(n452), .B(n425), .Z(n428) );
  XNOR U449 ( .A(p_input[45]), .B(p_input[77]), .Z(n425) );
  XNOR U450 ( .A(p_input[46]), .B(p_input[78]), .Z(n452) );
  XNOR U451 ( .A(p_input[41]), .B(p_input[73]), .Z(n420) );
  XNOR U452 ( .A(n446), .B(n396), .Z(n448) );
  XOR U453 ( .A(n435), .B(n434), .Z(n396) );
  XOR U454 ( .A(n453), .B(n440), .Z(n434) );
  XNOR U455 ( .A(p_input[40]), .B(p_input[72]), .Z(n440) );
  XOR U456 ( .A(n431), .B(n439), .Z(n453) );
  XOR U457 ( .A(n454), .B(n436), .Z(n439) );
  XNOR U458 ( .A(p_input[38]), .B(p_input[70]), .Z(n436) );
  XNOR U459 ( .A(p_input[39]), .B(p_input[71]), .Z(n454) );
  XNOR U460 ( .A(p_input[34]), .B(p_input[66]), .Z(n431) );
  XOR U461 ( .A(n445), .B(n444), .Z(n435) );
  XNOR U462 ( .A(n455), .B(n441), .Z(n444) );
  XOR U463 ( .A(p_input[35]), .B(p_input[67]), .Z(n441) );
  XNOR U464 ( .A(p_input[36]), .B(p_input[68]), .Z(n455) );
  XNOR U465 ( .A(p_input[37]), .B(p_input[69]), .Z(n445) );
  XOR U466 ( .A(p_input[33]), .B(p_input[65]), .Z(n446) );
  AND U467 ( .A(n149), .B(n456), .Z(n181) );
  XOR U468 ( .A(n457), .B(n458), .Z(n149) );
  XOR U469 ( .A(n459), .B(n456), .Z(n458) );
  AND U470 ( .A(n159), .B(n460), .Z(n456) );
  XNOR U471 ( .A(n461), .B(n462), .Z(n159) );
  XOR U472 ( .A(n463), .B(n460), .Z(n461) );
  AND U473 ( .A(n170), .B(n464), .Z(n460) );
  XNOR U474 ( .A(n465), .B(n466), .Z(n170) );
  XOR U475 ( .A(n467), .B(n464), .Z(n465) );
  AND U476 ( .A(n176), .B(n468), .Z(n464) );
  XOR U477 ( .A(n469), .B(n468), .Z(n176) );
  XOR U478 ( .A(p_input[16]), .B(p_input[64]), .Z(n468) );
  XOR U479 ( .A(n470), .B(n471), .Z(n469) );
  NOR U480 ( .A(n472), .B(n462), .Z(n459) );
  XNOR U481 ( .A(n473), .B(n457), .Z(n462) );
  XOR U482 ( .A(n474), .B(n475), .Z(n473) );
  AND U483 ( .A(n476), .B(n477), .Z(n475) );
  XOR U484 ( .A(n474), .B(n478), .Z(n476) );
  XNOR U485 ( .A(n463), .B(n457), .Z(n472) );
  XOR U486 ( .A(n479), .B(n480), .Z(n463) );
  AND U487 ( .A(n481), .B(n482), .Z(n480) );
  XOR U488 ( .A(n479), .B(n483), .Z(n481) );
  XOR U489 ( .A(n484), .B(n485), .Z(n457) );
  NOR U490 ( .A(n486), .B(n466), .Z(n485) );
  XNOR U491 ( .A(n487), .B(n478), .Z(n466) );
  XOR U492 ( .A(n488), .B(n489), .Z(n478) );
  AND U493 ( .A(n490), .B(n491), .Z(n489) );
  XOR U494 ( .A(n488), .B(n492), .Z(n490) );
  XOR U495 ( .A(n477), .B(n484), .Z(n487) );
  XOR U496 ( .A(n493), .B(n474), .Z(n477) );
  XOR U497 ( .A(n494), .B(n495), .Z(n474) );
  AND U498 ( .A(n496), .B(n497), .Z(n495) );
  XOR U499 ( .A(n494), .B(n498), .Z(n496) );
  XOR U500 ( .A(n499), .B(n500), .Z(n493) );
  AND U501 ( .A(n501), .B(n502), .Z(n500) );
  XOR U502 ( .A(n499), .B(n503), .Z(n501) );
  XNOR U503 ( .A(n467), .B(n484), .Z(n486) );
  XOR U504 ( .A(n483), .B(n482), .Z(n467) );
  XOR U505 ( .A(n504), .B(n479), .Z(n482) );
  XOR U506 ( .A(n505), .B(n506), .Z(n479) );
  AND U507 ( .A(n507), .B(n508), .Z(n506) );
  XOR U508 ( .A(n505), .B(n509), .Z(n507) );
  XOR U509 ( .A(n510), .B(n511), .Z(n504) );
  AND U510 ( .A(n512), .B(n513), .Z(n511) );
  XOR U511 ( .A(n510), .B(n514), .Z(n512) );
  XNOR U512 ( .A(n515), .B(n516), .Z(n483) );
  AND U513 ( .A(n517), .B(n518), .Z(n516) );
  XNOR U514 ( .A(n515), .B(n519), .Z(n517) );
  XNOR U515 ( .A(n520), .B(n521), .Z(n484) );
  AND U516 ( .A(n522), .B(n471), .Z(n521) );
  XOR U517 ( .A(n523), .B(n498), .Z(n471) );
  XOR U518 ( .A(n492), .B(n491), .Z(n498) );
  XOR U519 ( .A(n524), .B(n488), .Z(n491) );
  XNOR U520 ( .A(p_input[26]), .B(p_input[74]), .Z(n488) );
  XNOR U521 ( .A(p_input[27]), .B(p_input[75]), .Z(n524) );
  XNOR U522 ( .A(p_input[28]), .B(p_input[76]), .Z(n492) );
  XNOR U523 ( .A(n497), .B(n520), .Z(n523) );
  XOR U524 ( .A(n525), .B(n503), .Z(n497) );
  XNOR U525 ( .A(p_input[31]), .B(p_input[79]), .Z(n503) );
  XOR U526 ( .A(n494), .B(n502), .Z(n525) );
  XOR U527 ( .A(n526), .B(n499), .Z(n502) );
  XNOR U528 ( .A(p_input[29]), .B(p_input[77]), .Z(n499) );
  XNOR U529 ( .A(p_input[30]), .B(p_input[78]), .Z(n526) );
  XNOR U530 ( .A(p_input[25]), .B(p_input[73]), .Z(n494) );
  XNOR U531 ( .A(n520), .B(n470), .Z(n522) );
  XOR U532 ( .A(n509), .B(n508), .Z(n470) );
  XOR U533 ( .A(n527), .B(n514), .Z(n508) );
  XNOR U534 ( .A(p_input[24]), .B(p_input[72]), .Z(n514) );
  XOR U535 ( .A(n505), .B(n513), .Z(n527) );
  XOR U536 ( .A(n528), .B(n510), .Z(n513) );
  XNOR U537 ( .A(p_input[22]), .B(p_input[70]), .Z(n510) );
  XNOR U538 ( .A(p_input[23]), .B(p_input[71]), .Z(n528) );
  XNOR U539 ( .A(p_input[18]), .B(p_input[66]), .Z(n505) );
  XOR U540 ( .A(n519), .B(n518), .Z(n509) );
  XNOR U541 ( .A(n529), .B(n515), .Z(n518) );
  XOR U542 ( .A(p_input[19]), .B(p_input[67]), .Z(n515) );
  XNOR U543 ( .A(p_input[20]), .B(p_input[68]), .Z(n529) );
  XNOR U544 ( .A(p_input[21]), .B(p_input[69]), .Z(n519) );
  XOR U545 ( .A(p_input[17]), .B(p_input[65]), .Z(n520) );
endmodule

