
module knn_comb_BMR_W32_K3_N8 ( p_input, o );
  input [287:0] p_input;
  output [95:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/min_val_out[0][16] , \knn_comb_/min_val_out[0][17] ,
         \knn_comb_/min_val_out[0][18] , \knn_comb_/min_val_out[0][19] ,
         \knn_comb_/min_val_out[0][20] , \knn_comb_/min_val_out[0][21] ,
         \knn_comb_/min_val_out[0][22] , \knn_comb_/min_val_out[0][23] ,
         \knn_comb_/min_val_out[0][24] , \knn_comb_/min_val_out[0][25] ,
         \knn_comb_/min_val_out[0][26] , \knn_comb_/min_val_out[0][27] ,
         \knn_comb_/min_val_out[0][28] , \knn_comb_/min_val_out[0][29] ,
         \knn_comb_/min_val_out[0][30] , \knn_comb_/min_val_out[0][31] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][16] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][17] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][18] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][19] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][20] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][21] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][22] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][23] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][24] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][25] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][26] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][27] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][28] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][29] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][30] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][31] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][31] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039;
  assign \knn_comb_/min_val_out[0][0]  = p_input[224];
  assign \knn_comb_/min_val_out[0][1]  = p_input[225];
  assign \knn_comb_/min_val_out[0][2]  = p_input[226];
  assign \knn_comb_/min_val_out[0][3]  = p_input[227];
  assign \knn_comb_/min_val_out[0][4]  = p_input[228];
  assign \knn_comb_/min_val_out[0][5]  = p_input[229];
  assign \knn_comb_/min_val_out[0][6]  = p_input[230];
  assign \knn_comb_/min_val_out[0][7]  = p_input[231];
  assign \knn_comb_/min_val_out[0][8]  = p_input[232];
  assign \knn_comb_/min_val_out[0][9]  = p_input[233];
  assign \knn_comb_/min_val_out[0][10]  = p_input[234];
  assign \knn_comb_/min_val_out[0][11]  = p_input[235];
  assign \knn_comb_/min_val_out[0][12]  = p_input[236];
  assign \knn_comb_/min_val_out[0][13]  = p_input[237];
  assign \knn_comb_/min_val_out[0][14]  = p_input[238];
  assign \knn_comb_/min_val_out[0][15]  = p_input[239];
  assign \knn_comb_/min_val_out[0][16]  = p_input[240];
  assign \knn_comb_/min_val_out[0][17]  = p_input[241];
  assign \knn_comb_/min_val_out[0][18]  = p_input[242];
  assign \knn_comb_/min_val_out[0][19]  = p_input[243];
  assign \knn_comb_/min_val_out[0][20]  = p_input[244];
  assign \knn_comb_/min_val_out[0][21]  = p_input[245];
  assign \knn_comb_/min_val_out[0][22]  = p_input[246];
  assign \knn_comb_/min_val_out[0][23]  = p_input[247];
  assign \knn_comb_/min_val_out[0][24]  = p_input[248];
  assign \knn_comb_/min_val_out[0][25]  = p_input[249];
  assign \knn_comb_/min_val_out[0][26]  = p_input[250];
  assign \knn_comb_/min_val_out[0][27]  = p_input[251];
  assign \knn_comb_/min_val_out[0][28]  = p_input[252];
  assign \knn_comb_/min_val_out[0][29]  = p_input[253];
  assign \knn_comb_/min_val_out[0][30]  = p_input[254];
  assign \knn_comb_/min_val_out[0][31]  = p_input[255];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][0]  = p_input[160];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][1]  = p_input[161];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][2]  = p_input[162];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][3]  = p_input[163];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][4]  = p_input[164];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][5]  = p_input[165];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][6]  = p_input[166];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][7]  = p_input[167];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][8]  = p_input[168];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][9]  = p_input[169];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][10]  = p_input[170];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][11]  = p_input[171];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][12]  = p_input[172];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][13]  = p_input[173];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][14]  = p_input[174];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][15]  = p_input[175];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][16]  = p_input[176];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][17]  = p_input[177];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][18]  = p_input[178];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][19]  = p_input[179];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][20]  = p_input[180];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][21]  = p_input[181];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][22]  = p_input[182];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][23]  = p_input[183];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][24]  = p_input[184];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][25]  = p_input[185];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][26]  = p_input[186];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][27]  = p_input[187];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][28]  = p_input[188];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][29]  = p_input[189];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][30]  = p_input[190];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][31]  = p_input[191];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][0]  = p_input[192];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][1]  = p_input[193];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][2]  = p_input[194];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][3]  = p_input[195];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][4]  = p_input[196];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][5]  = p_input[197];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][6]  = p_input[198];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][7]  = p_input[199];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][8]  = p_input[200];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][9]  = p_input[201];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][10]  = p_input[202];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][11]  = p_input[203];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][12]  = p_input[204];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][13]  = p_input[205];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][14]  = p_input[206];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][15]  = p_input[207];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][16]  = p_input[208];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][17]  = p_input[209];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][18]  = p_input[210];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][19]  = p_input[211];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][20]  = p_input[212];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][21]  = p_input[213];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][22]  = p_input[214];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][23]  = p_input[215];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][24]  = p_input[216];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][25]  = p_input[217];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][26]  = p_input[218];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][27]  = p_input[219];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][28]  = p_input[220];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][29]  = p_input[221];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][30]  = p_input[222];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][31]  = p_input[223];

  XOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  XOR U2 ( .A(n3), .B(n4), .Z(o[95]) );
  XOR U3 ( .A(n5), .B(n6), .Z(o[94]) );
  XOR U4 ( .A(n7), .B(n8), .Z(o[93]) );
  XOR U5 ( .A(n9), .B(n10), .Z(o[92]) );
  XOR U6 ( .A(n11), .B(n12), .Z(o[91]) );
  XOR U7 ( .A(n13), .B(n14), .Z(o[90]) );
  XOR U8 ( .A(n15), .B(n16), .Z(o[8]) );
  XOR U9 ( .A(n17), .B(n18), .Z(o[89]) );
  XOR U10 ( .A(n19), .B(n20), .Z(o[88]) );
  XOR U11 ( .A(n21), .B(n22), .Z(o[87]) );
  XOR U12 ( .A(n23), .B(n24), .Z(o[86]) );
  XOR U13 ( .A(n25), .B(n26), .Z(o[85]) );
  XOR U14 ( .A(n27), .B(n28), .Z(o[84]) );
  XOR U15 ( .A(n29), .B(n30), .Z(o[83]) );
  XOR U16 ( .A(n31), .B(n32), .Z(o[82]) );
  XOR U17 ( .A(n33), .B(n34), .Z(o[81]) );
  XOR U18 ( .A(n35), .B(n36), .Z(o[80]) );
  XOR U19 ( .A(n37), .B(n38), .Z(o[7]) );
  XOR U20 ( .A(n39), .B(n40), .Z(o[79]) );
  XOR U21 ( .A(n41), .B(n42), .Z(o[78]) );
  XOR U22 ( .A(n43), .B(n44), .Z(o[77]) );
  XOR U23 ( .A(n45), .B(n46), .Z(o[76]) );
  XOR U24 ( .A(n47), .B(n48), .Z(o[75]) );
  XOR U25 ( .A(n49), .B(n50), .Z(o[74]) );
  XOR U26 ( .A(n51), .B(n52), .Z(o[73]) );
  XOR U27 ( .A(n53), .B(n54), .Z(o[72]) );
  XOR U28 ( .A(n55), .B(n56), .Z(o[71]) );
  XOR U29 ( .A(n57), .B(n58), .Z(o[70]) );
  XOR U30 ( .A(n59), .B(n60), .Z(o[6]) );
  XOR U31 ( .A(n61), .B(n62), .Z(o[69]) );
  XOR U32 ( .A(n63), .B(n64), .Z(o[68]) );
  XOR U33 ( .A(n65), .B(n66), .Z(o[67]) );
  XOR U34 ( .A(n67), .B(n68), .Z(o[66]) );
  XOR U35 ( .A(n69), .B(n70), .Z(o[65]) );
  XOR U36 ( .A(n71), .B(n72), .Z(o[64]) );
  XOR U37 ( .A(n73), .B(n74), .Z(o[63]) );
  XOR U38 ( .A(n75), .B(n76), .Z(o[62]) );
  XOR U39 ( .A(n77), .B(n78), .Z(o[61]) );
  XOR U40 ( .A(n79), .B(n80), .Z(o[60]) );
  XOR U41 ( .A(n81), .B(n82), .Z(o[5]) );
  XOR U42 ( .A(n83), .B(n84), .Z(o[59]) );
  XOR U43 ( .A(n85), .B(n86), .Z(o[58]) );
  XOR U44 ( .A(n87), .B(n88), .Z(o[57]) );
  XOR U45 ( .A(n89), .B(n90), .Z(o[56]) );
  XOR U46 ( .A(n91), .B(n92), .Z(o[55]) );
  XOR U47 ( .A(n93), .B(n94), .Z(o[54]) );
  XOR U48 ( .A(n95), .B(n96), .Z(o[53]) );
  XOR U49 ( .A(n97), .B(n98), .Z(o[52]) );
  XOR U50 ( .A(n99), .B(n100), .Z(o[51]) );
  XOR U51 ( .A(n101), .B(n102), .Z(o[50]) );
  XOR U52 ( .A(n103), .B(n104), .Z(o[4]) );
  XOR U53 ( .A(n105), .B(n106), .Z(o[49]) );
  XOR U54 ( .A(n107), .B(n108), .Z(o[48]) );
  XOR U55 ( .A(n109), .B(n110), .Z(o[47]) );
  XOR U56 ( .A(n111), .B(n112), .Z(o[46]) );
  XOR U57 ( .A(n113), .B(n114), .Z(o[45]) );
  XOR U58 ( .A(n115), .B(n116), .Z(o[44]) );
  XOR U59 ( .A(n117), .B(n118), .Z(o[43]) );
  XOR U60 ( .A(n119), .B(n120), .Z(o[42]) );
  XOR U61 ( .A(n1), .B(n121), .Z(o[41]) );
  AND U62 ( .A(n122), .B(n123), .Z(n1) );
  XOR U63 ( .A(n2), .B(n121), .Z(n123) );
  XOR U64 ( .A(n124), .B(n51), .Z(n121) );
  AND U65 ( .A(n125), .B(n126), .Z(n51) );
  XNOR U66 ( .A(n127), .B(n52), .Z(n126) );
  XOR U67 ( .A(n128), .B(n129), .Z(n52) );
  AND U68 ( .A(n130), .B(n131), .Z(n129) );
  XOR U69 ( .A(p_input[9]), .B(n128), .Z(n131) );
  XOR U70 ( .A(n132), .B(n133), .Z(n128) );
  AND U71 ( .A(n134), .B(n135), .Z(n133) );
  IV U72 ( .A(n124), .Z(n127) );
  XOR U73 ( .A(n136), .B(n137), .Z(n124) );
  AND U74 ( .A(n138), .B(n139), .Z(n137) );
  XOR U75 ( .A(n140), .B(n141), .Z(n2) );
  AND U76 ( .A(n142), .B(n139), .Z(n141) );
  XNOR U77 ( .A(n143), .B(n136), .Z(n139) );
  XOR U78 ( .A(n144), .B(n145), .Z(n136) );
  AND U79 ( .A(n146), .B(n135), .Z(n145) );
  XNOR U80 ( .A(n147), .B(n132), .Z(n135) );
  XOR U81 ( .A(n148), .B(n149), .Z(n132) );
  AND U82 ( .A(n150), .B(n151), .Z(n149) );
  XOR U83 ( .A(p_input[41]), .B(n148), .Z(n151) );
  XOR U84 ( .A(n152), .B(n153), .Z(n148) );
  AND U85 ( .A(n154), .B(n155), .Z(n153) );
  IV U86 ( .A(n144), .Z(n147) );
  XOR U87 ( .A(n156), .B(n157), .Z(n144) );
  AND U88 ( .A(n158), .B(n159), .Z(n157) );
  IV U89 ( .A(n140), .Z(n143) );
  XNOR U90 ( .A(n160), .B(n161), .Z(n140) );
  AND U91 ( .A(n162), .B(n159), .Z(n161) );
  XNOR U92 ( .A(n160), .B(n156), .Z(n159) );
  XOR U93 ( .A(n163), .B(n164), .Z(n156) );
  AND U94 ( .A(n165), .B(n155), .Z(n164) );
  XNOR U95 ( .A(n166), .B(n152), .Z(n155) );
  XOR U96 ( .A(n167), .B(n168), .Z(n152) );
  AND U97 ( .A(n169), .B(n170), .Z(n168) );
  XOR U98 ( .A(p_input[73]), .B(n167), .Z(n170) );
  XOR U99 ( .A(n171), .B(n172), .Z(n167) );
  AND U100 ( .A(n173), .B(n174), .Z(n172) );
  IV U101 ( .A(n163), .Z(n166) );
  XOR U102 ( .A(n175), .B(n176), .Z(n163) );
  AND U103 ( .A(n177), .B(n178), .Z(n176) );
  XOR U104 ( .A(n179), .B(n180), .Z(n160) );
  AND U105 ( .A(n181), .B(n178), .Z(n180) );
  XNOR U106 ( .A(n179), .B(n175), .Z(n178) );
  XOR U107 ( .A(n182), .B(n183), .Z(n175) );
  AND U108 ( .A(n184), .B(n174), .Z(n183) );
  XNOR U109 ( .A(n185), .B(n171), .Z(n174) );
  XOR U110 ( .A(n186), .B(n187), .Z(n171) );
  AND U111 ( .A(n188), .B(n189), .Z(n187) );
  XOR U112 ( .A(p_input[105]), .B(n186), .Z(n189) );
  XOR U113 ( .A(n190), .B(n191), .Z(n186) );
  AND U114 ( .A(n192), .B(n193), .Z(n191) );
  IV U115 ( .A(n182), .Z(n185) );
  XOR U116 ( .A(n194), .B(n195), .Z(n182) );
  AND U117 ( .A(n196), .B(n197), .Z(n195) );
  XOR U118 ( .A(n198), .B(n199), .Z(n179) );
  AND U119 ( .A(n200), .B(n197), .Z(n199) );
  XNOR U120 ( .A(n198), .B(n194), .Z(n197) );
  XOR U121 ( .A(n201), .B(n202), .Z(n194) );
  AND U122 ( .A(n203), .B(n193), .Z(n202) );
  XNOR U123 ( .A(n204), .B(n190), .Z(n193) );
  XOR U124 ( .A(n205), .B(n206), .Z(n190) );
  AND U125 ( .A(n207), .B(n208), .Z(n206) );
  XOR U126 ( .A(p_input[137]), .B(n205), .Z(n208) );
  XOR U127 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(n209), .Z(
        n205) );
  AND U128 ( .A(n210), .B(n211), .Z(n209) );
  IV U129 ( .A(n201), .Z(n204) );
  XOR U130 ( .A(n212), .B(n213), .Z(n201) );
  AND U131 ( .A(n214), .B(n215), .Z(n213) );
  XOR U132 ( .A(n216), .B(n217), .Z(n198) );
  AND U133 ( .A(n218), .B(n215), .Z(n217) );
  XNOR U134 ( .A(n216), .B(n212), .Z(n215) );
  XNOR U135 ( .A(n219), .B(n220), .Z(n212) );
  AND U136 ( .A(n221), .B(n211), .Z(n220) );
  XNOR U137 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(n219), .Z(
        n211) );
  XNOR U138 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .B(n222), .Z(
        n219) );
  AND U139 ( .A(n223), .B(n224), .Z(n222) );
  XNOR U140 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n225), .Z(n216) );
  AND U141 ( .A(n226), .B(n224), .Z(n225) );
  XOR U142 ( .A(n227), .B(n228), .Z(n224) );
  XOR U143 ( .A(n15), .B(n229), .Z(o[40]) );
  AND U144 ( .A(n122), .B(n230), .Z(n15) );
  XOR U145 ( .A(n16), .B(n229), .Z(n230) );
  XOR U146 ( .A(n231), .B(n53), .Z(n229) );
  AND U147 ( .A(n125), .B(n232), .Z(n53) );
  XNOR U148 ( .A(n233), .B(n54), .Z(n232) );
  XOR U149 ( .A(n234), .B(n235), .Z(n54) );
  AND U150 ( .A(n130), .B(n236), .Z(n235) );
  XOR U151 ( .A(p_input[8]), .B(n234), .Z(n236) );
  XOR U152 ( .A(n237), .B(n238), .Z(n234) );
  AND U153 ( .A(n134), .B(n239), .Z(n238) );
  IV U154 ( .A(n231), .Z(n233) );
  XOR U155 ( .A(n240), .B(n241), .Z(n231) );
  AND U156 ( .A(n138), .B(n242), .Z(n241) );
  XOR U157 ( .A(n243), .B(n244), .Z(n16) );
  AND U158 ( .A(n142), .B(n242), .Z(n244) );
  XNOR U159 ( .A(n245), .B(n240), .Z(n242) );
  XOR U160 ( .A(n246), .B(n247), .Z(n240) );
  AND U161 ( .A(n146), .B(n239), .Z(n247) );
  XNOR U162 ( .A(n248), .B(n237), .Z(n239) );
  XOR U163 ( .A(n249), .B(n250), .Z(n237) );
  AND U164 ( .A(n150), .B(n251), .Z(n250) );
  XOR U165 ( .A(p_input[40]), .B(n249), .Z(n251) );
  XOR U166 ( .A(n252), .B(n253), .Z(n249) );
  AND U167 ( .A(n154), .B(n254), .Z(n253) );
  IV U168 ( .A(n246), .Z(n248) );
  XOR U169 ( .A(n255), .B(n256), .Z(n246) );
  AND U170 ( .A(n158), .B(n257), .Z(n256) );
  IV U171 ( .A(n243), .Z(n245) );
  XNOR U172 ( .A(n258), .B(n259), .Z(n243) );
  AND U173 ( .A(n162), .B(n257), .Z(n259) );
  XNOR U174 ( .A(n258), .B(n255), .Z(n257) );
  XOR U175 ( .A(n260), .B(n261), .Z(n255) );
  AND U176 ( .A(n165), .B(n254), .Z(n261) );
  XNOR U177 ( .A(n262), .B(n252), .Z(n254) );
  XOR U178 ( .A(n263), .B(n264), .Z(n252) );
  AND U179 ( .A(n169), .B(n265), .Z(n264) );
  XOR U180 ( .A(p_input[72]), .B(n263), .Z(n265) );
  XOR U181 ( .A(n266), .B(n267), .Z(n263) );
  AND U182 ( .A(n173), .B(n268), .Z(n267) );
  IV U183 ( .A(n260), .Z(n262) );
  XOR U184 ( .A(n269), .B(n270), .Z(n260) );
  AND U185 ( .A(n177), .B(n271), .Z(n270) );
  XOR U186 ( .A(n272), .B(n273), .Z(n258) );
  AND U187 ( .A(n181), .B(n271), .Z(n273) );
  XNOR U188 ( .A(n272), .B(n269), .Z(n271) );
  XOR U189 ( .A(n274), .B(n275), .Z(n269) );
  AND U190 ( .A(n184), .B(n268), .Z(n275) );
  XNOR U191 ( .A(n276), .B(n266), .Z(n268) );
  XOR U192 ( .A(n277), .B(n278), .Z(n266) );
  AND U193 ( .A(n188), .B(n279), .Z(n278) );
  XOR U194 ( .A(p_input[104]), .B(n277), .Z(n279) );
  XOR U195 ( .A(n280), .B(n281), .Z(n277) );
  AND U196 ( .A(n192), .B(n282), .Z(n281) );
  IV U197 ( .A(n274), .Z(n276) );
  XOR U198 ( .A(n283), .B(n284), .Z(n274) );
  AND U199 ( .A(n196), .B(n285), .Z(n284) );
  XOR U200 ( .A(n286), .B(n287), .Z(n272) );
  AND U201 ( .A(n200), .B(n285), .Z(n287) );
  XNOR U202 ( .A(n286), .B(n283), .Z(n285) );
  XOR U203 ( .A(n288), .B(n289), .Z(n283) );
  AND U204 ( .A(n203), .B(n282), .Z(n289) );
  XNOR U205 ( .A(n290), .B(n280), .Z(n282) );
  XOR U206 ( .A(n291), .B(n292), .Z(n280) );
  AND U207 ( .A(n207), .B(n293), .Z(n292) );
  XOR U208 ( .A(p_input[136]), .B(n291), .Z(n293) );
  XOR U209 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n294), .Z(
        n291) );
  AND U210 ( .A(n210), .B(n295), .Z(n294) );
  IV U211 ( .A(n288), .Z(n290) );
  XOR U212 ( .A(n296), .B(n297), .Z(n288) );
  AND U213 ( .A(n214), .B(n298), .Z(n297) );
  XOR U214 ( .A(n299), .B(n300), .Z(n286) );
  AND U215 ( .A(n218), .B(n298), .Z(n300) );
  XNOR U216 ( .A(n299), .B(n296), .Z(n298) );
  XNOR U217 ( .A(n301), .B(n302), .Z(n296) );
  AND U218 ( .A(n221), .B(n295), .Z(n302) );
  XNOR U219 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n301), .Z(
        n295) );
  XNOR U220 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .B(n303), .Z(
        n301) );
  AND U221 ( .A(n223), .B(n304), .Z(n303) );
  XNOR U222 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n305), .Z(n299) );
  AND U223 ( .A(n226), .B(n304), .Z(n305) );
  XOR U224 ( .A(n306), .B(n307), .Z(n304) );
  IV U225 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .Z(n307) );
  IV U226 ( .A(\knn_comb_/min_val_out[0][8] ), .Z(n306) );
  XOR U227 ( .A(n308), .B(n309), .Z(o[3]) );
  XOR U228 ( .A(n37), .B(n310), .Z(o[39]) );
  AND U229 ( .A(n122), .B(n311), .Z(n37) );
  XOR U230 ( .A(n38), .B(n310), .Z(n311) );
  XOR U231 ( .A(n312), .B(n55), .Z(n310) );
  AND U232 ( .A(n125), .B(n313), .Z(n55) );
  XNOR U233 ( .A(n314), .B(n56), .Z(n313) );
  XOR U234 ( .A(n315), .B(n316), .Z(n56) );
  AND U235 ( .A(n130), .B(n317), .Z(n316) );
  XOR U236 ( .A(p_input[7]), .B(n315), .Z(n317) );
  XOR U237 ( .A(n318), .B(n319), .Z(n315) );
  AND U238 ( .A(n134), .B(n320), .Z(n319) );
  IV U239 ( .A(n312), .Z(n314) );
  XOR U240 ( .A(n321), .B(n322), .Z(n312) );
  AND U241 ( .A(n138), .B(n323), .Z(n322) );
  XOR U242 ( .A(n324), .B(n325), .Z(n38) );
  AND U243 ( .A(n142), .B(n323), .Z(n325) );
  XNOR U244 ( .A(n326), .B(n321), .Z(n323) );
  XOR U245 ( .A(n327), .B(n328), .Z(n321) );
  AND U246 ( .A(n146), .B(n320), .Z(n328) );
  XNOR U247 ( .A(n329), .B(n318), .Z(n320) );
  XOR U248 ( .A(n330), .B(n331), .Z(n318) );
  AND U249 ( .A(n150), .B(n332), .Z(n331) );
  XOR U250 ( .A(p_input[39]), .B(n330), .Z(n332) );
  XOR U251 ( .A(n333), .B(n334), .Z(n330) );
  AND U252 ( .A(n154), .B(n335), .Z(n334) );
  IV U253 ( .A(n327), .Z(n329) );
  XOR U254 ( .A(n336), .B(n337), .Z(n327) );
  AND U255 ( .A(n158), .B(n338), .Z(n337) );
  IV U256 ( .A(n324), .Z(n326) );
  XNOR U257 ( .A(n339), .B(n340), .Z(n324) );
  AND U258 ( .A(n162), .B(n338), .Z(n340) );
  XNOR U259 ( .A(n339), .B(n336), .Z(n338) );
  XOR U260 ( .A(n341), .B(n342), .Z(n336) );
  AND U261 ( .A(n165), .B(n335), .Z(n342) );
  XNOR U262 ( .A(n343), .B(n333), .Z(n335) );
  XOR U263 ( .A(n344), .B(n345), .Z(n333) );
  AND U264 ( .A(n169), .B(n346), .Z(n345) );
  XOR U265 ( .A(p_input[71]), .B(n344), .Z(n346) );
  XOR U266 ( .A(n347), .B(n348), .Z(n344) );
  AND U267 ( .A(n173), .B(n349), .Z(n348) );
  IV U268 ( .A(n341), .Z(n343) );
  XOR U269 ( .A(n350), .B(n351), .Z(n341) );
  AND U270 ( .A(n177), .B(n352), .Z(n351) );
  XOR U271 ( .A(n353), .B(n354), .Z(n339) );
  AND U272 ( .A(n181), .B(n352), .Z(n354) );
  XNOR U273 ( .A(n353), .B(n350), .Z(n352) );
  XOR U274 ( .A(n355), .B(n356), .Z(n350) );
  AND U275 ( .A(n184), .B(n349), .Z(n356) );
  XNOR U276 ( .A(n357), .B(n347), .Z(n349) );
  XOR U277 ( .A(n358), .B(n359), .Z(n347) );
  AND U278 ( .A(n188), .B(n360), .Z(n359) );
  XOR U279 ( .A(p_input[103]), .B(n358), .Z(n360) );
  XOR U280 ( .A(n361), .B(n362), .Z(n358) );
  AND U281 ( .A(n192), .B(n363), .Z(n362) );
  IV U282 ( .A(n355), .Z(n357) );
  XOR U283 ( .A(n364), .B(n365), .Z(n355) );
  AND U284 ( .A(n196), .B(n366), .Z(n365) );
  XOR U285 ( .A(n367), .B(n368), .Z(n353) );
  AND U286 ( .A(n200), .B(n366), .Z(n368) );
  XNOR U287 ( .A(n367), .B(n364), .Z(n366) );
  XOR U288 ( .A(n369), .B(n370), .Z(n364) );
  AND U289 ( .A(n203), .B(n363), .Z(n370) );
  XNOR U290 ( .A(n371), .B(n361), .Z(n363) );
  XOR U291 ( .A(n372), .B(n373), .Z(n361) );
  AND U292 ( .A(n207), .B(n374), .Z(n373) );
  XOR U293 ( .A(p_input[135]), .B(n372), .Z(n374) );
  XOR U294 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(n375), .Z(
        n372) );
  AND U295 ( .A(n210), .B(n376), .Z(n375) );
  IV U296 ( .A(n369), .Z(n371) );
  XOR U297 ( .A(n377), .B(n378), .Z(n369) );
  AND U298 ( .A(n214), .B(n379), .Z(n378) );
  XOR U299 ( .A(n380), .B(n381), .Z(n367) );
  AND U300 ( .A(n218), .B(n379), .Z(n381) );
  XNOR U301 ( .A(n380), .B(n377), .Z(n379) );
  XNOR U302 ( .A(n382), .B(n383), .Z(n377) );
  AND U303 ( .A(n221), .B(n376), .Z(n383) );
  XNOR U304 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(n382), .Z(
        n376) );
  XNOR U305 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(n384), .Z(
        n382) );
  AND U306 ( .A(n223), .B(n385), .Z(n384) );
  XNOR U307 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n386), .Z(n380) );
  AND U308 ( .A(n226), .B(n385), .Z(n386) );
  XOR U309 ( .A(n387), .B(n388), .Z(n385) );
  XOR U310 ( .A(n59), .B(n389), .Z(o[38]) );
  AND U311 ( .A(n122), .B(n390), .Z(n59) );
  XOR U312 ( .A(n60), .B(n389), .Z(n390) );
  XOR U313 ( .A(n391), .B(n57), .Z(n389) );
  AND U314 ( .A(n125), .B(n392), .Z(n57) );
  XOR U315 ( .A(n58), .B(n391), .Z(n392) );
  XOR U316 ( .A(n393), .B(n394), .Z(n58) );
  AND U317 ( .A(n130), .B(n395), .Z(n394) );
  XOR U318 ( .A(p_input[6]), .B(n393), .Z(n395) );
  XNOR U319 ( .A(n396), .B(n397), .Z(n393) );
  AND U320 ( .A(n134), .B(n398), .Z(n397) );
  XOR U321 ( .A(n399), .B(n400), .Z(n391) );
  AND U322 ( .A(n138), .B(n401), .Z(n400) );
  XOR U323 ( .A(n402), .B(n403), .Z(n60) );
  AND U324 ( .A(n142), .B(n401), .Z(n403) );
  XNOR U325 ( .A(n404), .B(n402), .Z(n401) );
  IV U326 ( .A(n399), .Z(n404) );
  XOR U327 ( .A(n405), .B(n406), .Z(n399) );
  AND U328 ( .A(n146), .B(n398), .Z(n406) );
  XNOR U329 ( .A(n396), .B(n405), .Z(n398) );
  XNOR U330 ( .A(n407), .B(n408), .Z(n396) );
  AND U331 ( .A(n150), .B(n409), .Z(n408) );
  XOR U332 ( .A(p_input[38]), .B(n407), .Z(n409) );
  XNOR U333 ( .A(n410), .B(n411), .Z(n407) );
  AND U334 ( .A(n154), .B(n412), .Z(n411) );
  XOR U335 ( .A(n413), .B(n414), .Z(n405) );
  AND U336 ( .A(n158), .B(n415), .Z(n414) );
  XOR U337 ( .A(n416), .B(n417), .Z(n402) );
  AND U338 ( .A(n162), .B(n415), .Z(n417) );
  XNOR U339 ( .A(n418), .B(n416), .Z(n415) );
  IV U340 ( .A(n413), .Z(n418) );
  XOR U341 ( .A(n419), .B(n420), .Z(n413) );
  AND U342 ( .A(n165), .B(n412), .Z(n420) );
  XNOR U343 ( .A(n410), .B(n419), .Z(n412) );
  XNOR U344 ( .A(n421), .B(n422), .Z(n410) );
  AND U345 ( .A(n169), .B(n423), .Z(n422) );
  XOR U346 ( .A(p_input[70]), .B(n421), .Z(n423) );
  XNOR U347 ( .A(n424), .B(n425), .Z(n421) );
  AND U348 ( .A(n173), .B(n426), .Z(n425) );
  XOR U349 ( .A(n427), .B(n428), .Z(n419) );
  AND U350 ( .A(n177), .B(n429), .Z(n428) );
  XOR U351 ( .A(n430), .B(n431), .Z(n416) );
  AND U352 ( .A(n181), .B(n429), .Z(n431) );
  XNOR U353 ( .A(n432), .B(n430), .Z(n429) );
  IV U354 ( .A(n427), .Z(n432) );
  XOR U355 ( .A(n433), .B(n434), .Z(n427) );
  AND U356 ( .A(n184), .B(n426), .Z(n434) );
  XNOR U357 ( .A(n424), .B(n433), .Z(n426) );
  XNOR U358 ( .A(n435), .B(n436), .Z(n424) );
  AND U359 ( .A(n188), .B(n437), .Z(n436) );
  XOR U360 ( .A(p_input[102]), .B(n435), .Z(n437) );
  XNOR U361 ( .A(n438), .B(n439), .Z(n435) );
  AND U362 ( .A(n192), .B(n440), .Z(n439) );
  XOR U363 ( .A(n441), .B(n442), .Z(n433) );
  AND U364 ( .A(n196), .B(n443), .Z(n442) );
  XOR U365 ( .A(n444), .B(n445), .Z(n430) );
  AND U366 ( .A(n200), .B(n443), .Z(n445) );
  XNOR U367 ( .A(n446), .B(n444), .Z(n443) );
  IV U368 ( .A(n441), .Z(n446) );
  XOR U369 ( .A(n447), .B(n448), .Z(n441) );
  AND U370 ( .A(n203), .B(n440), .Z(n448) );
  XNOR U371 ( .A(n438), .B(n447), .Z(n440) );
  XNOR U372 ( .A(n449), .B(n450), .Z(n438) );
  AND U373 ( .A(n207), .B(n451), .Z(n450) );
  XOR U374 ( .A(p_input[134]), .B(n449), .Z(n451) );
  XOR U375 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(n452), .Z(
        n449) );
  AND U376 ( .A(n210), .B(n453), .Z(n452) );
  XOR U377 ( .A(n454), .B(n455), .Z(n447) );
  AND U378 ( .A(n214), .B(n456), .Z(n455) );
  XOR U379 ( .A(n457), .B(n458), .Z(n444) );
  AND U380 ( .A(n218), .B(n456), .Z(n458) );
  XNOR U381 ( .A(n459), .B(n457), .Z(n456) );
  IV U382 ( .A(n454), .Z(n459) );
  XOR U383 ( .A(n460), .B(n461), .Z(n454) );
  AND U384 ( .A(n221), .B(n453), .Z(n461) );
  XOR U385 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(n460), .Z(
        n453) );
  XOR U386 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .B(n462), .Z(
        n460) );
  AND U387 ( .A(n223), .B(n463), .Z(n462) );
  XOR U388 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n464), .Z(n457) );
  AND U389 ( .A(n226), .B(n463), .Z(n464) );
  XOR U390 ( .A(\knn_comb_/min_val_out[0][6] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .Z(n463) );
  XOR U391 ( .A(n81), .B(n465), .Z(o[37]) );
  AND U392 ( .A(n122), .B(n466), .Z(n81) );
  XOR U393 ( .A(n82), .B(n465), .Z(n466) );
  XOR U394 ( .A(n467), .B(n61), .Z(n465) );
  AND U395 ( .A(n125), .B(n468), .Z(n61) );
  XOR U396 ( .A(n62), .B(n467), .Z(n468) );
  XOR U397 ( .A(n469), .B(n470), .Z(n62) );
  AND U398 ( .A(n130), .B(n471), .Z(n470) );
  XOR U399 ( .A(p_input[5]), .B(n469), .Z(n471) );
  XNOR U400 ( .A(n472), .B(n473), .Z(n469) );
  AND U401 ( .A(n134), .B(n474), .Z(n473) );
  XOR U402 ( .A(n475), .B(n476), .Z(n467) );
  AND U403 ( .A(n138), .B(n477), .Z(n476) );
  XOR U404 ( .A(n478), .B(n479), .Z(n82) );
  AND U405 ( .A(n142), .B(n477), .Z(n479) );
  XNOR U406 ( .A(n480), .B(n478), .Z(n477) );
  IV U407 ( .A(n475), .Z(n480) );
  XOR U408 ( .A(n481), .B(n482), .Z(n475) );
  AND U409 ( .A(n146), .B(n474), .Z(n482) );
  XNOR U410 ( .A(n472), .B(n481), .Z(n474) );
  XNOR U411 ( .A(n483), .B(n484), .Z(n472) );
  AND U412 ( .A(n150), .B(n485), .Z(n484) );
  XOR U413 ( .A(p_input[37]), .B(n483), .Z(n485) );
  XNOR U414 ( .A(n486), .B(n487), .Z(n483) );
  AND U415 ( .A(n154), .B(n488), .Z(n487) );
  XOR U416 ( .A(n489), .B(n490), .Z(n481) );
  AND U417 ( .A(n158), .B(n491), .Z(n490) );
  XOR U418 ( .A(n492), .B(n493), .Z(n478) );
  AND U419 ( .A(n162), .B(n491), .Z(n493) );
  XNOR U420 ( .A(n494), .B(n492), .Z(n491) );
  IV U421 ( .A(n489), .Z(n494) );
  XOR U422 ( .A(n495), .B(n496), .Z(n489) );
  AND U423 ( .A(n165), .B(n488), .Z(n496) );
  XNOR U424 ( .A(n486), .B(n495), .Z(n488) );
  XNOR U425 ( .A(n497), .B(n498), .Z(n486) );
  AND U426 ( .A(n169), .B(n499), .Z(n498) );
  XOR U427 ( .A(p_input[69]), .B(n497), .Z(n499) );
  XNOR U428 ( .A(n500), .B(n501), .Z(n497) );
  AND U429 ( .A(n173), .B(n502), .Z(n501) );
  XOR U430 ( .A(n503), .B(n504), .Z(n495) );
  AND U431 ( .A(n177), .B(n505), .Z(n504) );
  XOR U432 ( .A(n506), .B(n507), .Z(n492) );
  AND U433 ( .A(n181), .B(n505), .Z(n507) );
  XNOR U434 ( .A(n508), .B(n506), .Z(n505) );
  IV U435 ( .A(n503), .Z(n508) );
  XOR U436 ( .A(n509), .B(n510), .Z(n503) );
  AND U437 ( .A(n184), .B(n502), .Z(n510) );
  XNOR U438 ( .A(n500), .B(n509), .Z(n502) );
  XNOR U439 ( .A(n511), .B(n512), .Z(n500) );
  AND U440 ( .A(n188), .B(n513), .Z(n512) );
  XOR U441 ( .A(p_input[101]), .B(n511), .Z(n513) );
  XNOR U442 ( .A(n514), .B(n515), .Z(n511) );
  AND U443 ( .A(n192), .B(n516), .Z(n515) );
  XOR U444 ( .A(n517), .B(n518), .Z(n509) );
  AND U445 ( .A(n196), .B(n519), .Z(n518) );
  XOR U446 ( .A(n520), .B(n521), .Z(n506) );
  AND U447 ( .A(n200), .B(n519), .Z(n521) );
  XNOR U448 ( .A(n522), .B(n520), .Z(n519) );
  IV U449 ( .A(n517), .Z(n522) );
  XOR U450 ( .A(n523), .B(n524), .Z(n517) );
  AND U451 ( .A(n203), .B(n516), .Z(n524) );
  XNOR U452 ( .A(n514), .B(n523), .Z(n516) );
  XNOR U453 ( .A(n525), .B(n526), .Z(n514) );
  AND U454 ( .A(n207), .B(n527), .Z(n526) );
  XOR U455 ( .A(p_input[133]), .B(n525), .Z(n527) );
  XOR U456 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n528), .Z(
        n525) );
  AND U457 ( .A(n210), .B(n529), .Z(n528) );
  XOR U458 ( .A(n530), .B(n531), .Z(n523) );
  AND U459 ( .A(n214), .B(n532), .Z(n531) );
  XOR U460 ( .A(n533), .B(n534), .Z(n520) );
  AND U461 ( .A(n218), .B(n532), .Z(n534) );
  XNOR U462 ( .A(n535), .B(n533), .Z(n532) );
  IV U463 ( .A(n530), .Z(n535) );
  XOR U464 ( .A(n536), .B(n537), .Z(n530) );
  AND U465 ( .A(n221), .B(n529), .Z(n537) );
  XOR U466 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n536), .Z(
        n529) );
  XOR U467 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(n538), .Z(
        n536) );
  AND U468 ( .A(n223), .B(n539), .Z(n538) );
  XOR U469 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n540), .Z(n533) );
  AND U470 ( .A(n226), .B(n539), .Z(n540) );
  XOR U471 ( .A(n541), .B(n542), .Z(n539) );
  IV U472 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .Z(n542) );
  IV U473 ( .A(\knn_comb_/min_val_out[0][5] ), .Z(n541) );
  XOR U474 ( .A(n103), .B(n543), .Z(o[36]) );
  AND U475 ( .A(n122), .B(n544), .Z(n103) );
  XOR U476 ( .A(n104), .B(n543), .Z(n544) );
  XOR U477 ( .A(n545), .B(n63), .Z(n543) );
  AND U478 ( .A(n125), .B(n546), .Z(n63) );
  XOR U479 ( .A(n64), .B(n545), .Z(n546) );
  XOR U480 ( .A(n547), .B(n548), .Z(n64) );
  AND U481 ( .A(n130), .B(n549), .Z(n548) );
  XOR U482 ( .A(p_input[4]), .B(n547), .Z(n549) );
  XNOR U483 ( .A(n550), .B(n551), .Z(n547) );
  AND U484 ( .A(n134), .B(n552), .Z(n551) );
  XOR U485 ( .A(n553), .B(n554), .Z(n545) );
  AND U486 ( .A(n138), .B(n555), .Z(n554) );
  XOR U487 ( .A(n556), .B(n557), .Z(n104) );
  AND U488 ( .A(n142), .B(n555), .Z(n557) );
  XNOR U489 ( .A(n558), .B(n556), .Z(n555) );
  IV U490 ( .A(n553), .Z(n558) );
  XOR U491 ( .A(n559), .B(n560), .Z(n553) );
  AND U492 ( .A(n146), .B(n552), .Z(n560) );
  XNOR U493 ( .A(n550), .B(n559), .Z(n552) );
  XNOR U494 ( .A(n561), .B(n562), .Z(n550) );
  AND U495 ( .A(n150), .B(n563), .Z(n562) );
  XOR U496 ( .A(p_input[36]), .B(n561), .Z(n563) );
  XNOR U497 ( .A(n564), .B(n565), .Z(n561) );
  AND U498 ( .A(n154), .B(n566), .Z(n565) );
  XOR U499 ( .A(n567), .B(n568), .Z(n559) );
  AND U500 ( .A(n158), .B(n569), .Z(n568) );
  XOR U501 ( .A(n570), .B(n571), .Z(n556) );
  AND U502 ( .A(n162), .B(n569), .Z(n571) );
  XNOR U503 ( .A(n572), .B(n570), .Z(n569) );
  IV U504 ( .A(n567), .Z(n572) );
  XOR U505 ( .A(n573), .B(n574), .Z(n567) );
  AND U506 ( .A(n165), .B(n566), .Z(n574) );
  XNOR U507 ( .A(n564), .B(n573), .Z(n566) );
  XNOR U508 ( .A(n575), .B(n576), .Z(n564) );
  AND U509 ( .A(n169), .B(n577), .Z(n576) );
  XOR U510 ( .A(p_input[68]), .B(n575), .Z(n577) );
  XNOR U511 ( .A(n578), .B(n579), .Z(n575) );
  AND U512 ( .A(n173), .B(n580), .Z(n579) );
  XOR U513 ( .A(n581), .B(n582), .Z(n573) );
  AND U514 ( .A(n177), .B(n583), .Z(n582) );
  XOR U515 ( .A(n584), .B(n585), .Z(n570) );
  AND U516 ( .A(n181), .B(n583), .Z(n585) );
  XNOR U517 ( .A(n586), .B(n584), .Z(n583) );
  IV U518 ( .A(n581), .Z(n586) );
  XOR U519 ( .A(n587), .B(n588), .Z(n581) );
  AND U520 ( .A(n184), .B(n580), .Z(n588) );
  XNOR U521 ( .A(n578), .B(n587), .Z(n580) );
  XNOR U522 ( .A(n589), .B(n590), .Z(n578) );
  AND U523 ( .A(n188), .B(n591), .Z(n590) );
  XOR U524 ( .A(p_input[100]), .B(n589), .Z(n591) );
  XNOR U525 ( .A(n592), .B(n593), .Z(n589) );
  AND U526 ( .A(n192), .B(n594), .Z(n593) );
  XOR U527 ( .A(n595), .B(n596), .Z(n587) );
  AND U528 ( .A(n196), .B(n597), .Z(n596) );
  XOR U529 ( .A(n598), .B(n599), .Z(n584) );
  AND U530 ( .A(n200), .B(n597), .Z(n599) );
  XNOR U531 ( .A(n600), .B(n598), .Z(n597) );
  IV U532 ( .A(n595), .Z(n600) );
  XOR U533 ( .A(n601), .B(n602), .Z(n595) );
  AND U534 ( .A(n203), .B(n594), .Z(n602) );
  XNOR U535 ( .A(n592), .B(n601), .Z(n594) );
  XNOR U536 ( .A(n603), .B(n604), .Z(n592) );
  AND U537 ( .A(n207), .B(n605), .Z(n604) );
  XOR U538 ( .A(p_input[132]), .B(n603), .Z(n605) );
  XOR U539 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(n606), .Z(
        n603) );
  AND U540 ( .A(n210), .B(n607), .Z(n606) );
  XOR U541 ( .A(n608), .B(n609), .Z(n601) );
  AND U542 ( .A(n214), .B(n610), .Z(n609) );
  XOR U543 ( .A(n611), .B(n612), .Z(n598) );
  AND U544 ( .A(n218), .B(n610), .Z(n612) );
  XNOR U545 ( .A(n613), .B(n611), .Z(n610) );
  IV U546 ( .A(n608), .Z(n613) );
  XOR U547 ( .A(n614), .B(n615), .Z(n608) );
  AND U548 ( .A(n221), .B(n607), .Z(n615) );
  XOR U549 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(n614), .Z(
        n607) );
  XOR U550 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(n616), .Z(
        n614) );
  AND U551 ( .A(n223), .B(n617), .Z(n616) );
  XOR U552 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n618), .Z(n611) );
  AND U553 ( .A(n226), .B(n617), .Z(n618) );
  XOR U554 ( .A(\knn_comb_/min_val_out[0][4] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .Z(n617) );
  XOR U555 ( .A(n308), .B(n619), .Z(o[35]) );
  AND U556 ( .A(n122), .B(n620), .Z(n308) );
  XOR U557 ( .A(n309), .B(n619), .Z(n620) );
  XOR U558 ( .A(n621), .B(n65), .Z(n619) );
  AND U559 ( .A(n125), .B(n622), .Z(n65) );
  XOR U560 ( .A(n66), .B(n621), .Z(n622) );
  XOR U561 ( .A(n623), .B(n624), .Z(n66) );
  AND U562 ( .A(n130), .B(n625), .Z(n624) );
  XOR U563 ( .A(p_input[3]), .B(n623), .Z(n625) );
  XNOR U564 ( .A(n626), .B(n627), .Z(n623) );
  AND U565 ( .A(n134), .B(n628), .Z(n627) );
  XOR U566 ( .A(n629), .B(n630), .Z(n621) );
  AND U567 ( .A(n138), .B(n631), .Z(n630) );
  XOR U568 ( .A(n632), .B(n633), .Z(n309) );
  AND U569 ( .A(n142), .B(n631), .Z(n633) );
  XNOR U570 ( .A(n634), .B(n632), .Z(n631) );
  IV U571 ( .A(n629), .Z(n634) );
  XOR U572 ( .A(n635), .B(n636), .Z(n629) );
  AND U573 ( .A(n146), .B(n628), .Z(n636) );
  XNOR U574 ( .A(n626), .B(n635), .Z(n628) );
  XNOR U575 ( .A(n637), .B(n638), .Z(n626) );
  AND U576 ( .A(n150), .B(n639), .Z(n638) );
  XOR U577 ( .A(p_input[35]), .B(n637), .Z(n639) );
  XNOR U578 ( .A(n640), .B(n641), .Z(n637) );
  AND U579 ( .A(n154), .B(n642), .Z(n641) );
  XOR U580 ( .A(n643), .B(n644), .Z(n635) );
  AND U581 ( .A(n158), .B(n645), .Z(n644) );
  XOR U582 ( .A(n646), .B(n647), .Z(n632) );
  AND U583 ( .A(n162), .B(n645), .Z(n647) );
  XNOR U584 ( .A(n648), .B(n646), .Z(n645) );
  IV U585 ( .A(n643), .Z(n648) );
  XOR U586 ( .A(n649), .B(n650), .Z(n643) );
  AND U587 ( .A(n165), .B(n642), .Z(n650) );
  XNOR U588 ( .A(n640), .B(n649), .Z(n642) );
  XNOR U589 ( .A(n651), .B(n652), .Z(n640) );
  AND U590 ( .A(n169), .B(n653), .Z(n652) );
  XOR U591 ( .A(p_input[67]), .B(n651), .Z(n653) );
  XNOR U592 ( .A(n654), .B(n655), .Z(n651) );
  AND U593 ( .A(n173), .B(n656), .Z(n655) );
  XOR U594 ( .A(n657), .B(n658), .Z(n649) );
  AND U595 ( .A(n177), .B(n659), .Z(n658) );
  XOR U596 ( .A(n660), .B(n661), .Z(n646) );
  AND U597 ( .A(n181), .B(n659), .Z(n661) );
  XNOR U598 ( .A(n662), .B(n660), .Z(n659) );
  IV U599 ( .A(n657), .Z(n662) );
  XOR U600 ( .A(n663), .B(n664), .Z(n657) );
  AND U601 ( .A(n184), .B(n656), .Z(n664) );
  XNOR U602 ( .A(n654), .B(n663), .Z(n656) );
  XNOR U603 ( .A(n665), .B(n666), .Z(n654) );
  AND U604 ( .A(n188), .B(n667), .Z(n666) );
  XOR U605 ( .A(p_input[99]), .B(n665), .Z(n667) );
  XNOR U606 ( .A(n668), .B(n669), .Z(n665) );
  AND U607 ( .A(n192), .B(n670), .Z(n669) );
  XOR U608 ( .A(n671), .B(n672), .Z(n663) );
  AND U609 ( .A(n196), .B(n673), .Z(n672) );
  XOR U610 ( .A(n674), .B(n675), .Z(n660) );
  AND U611 ( .A(n200), .B(n673), .Z(n675) );
  XNOR U612 ( .A(n676), .B(n674), .Z(n673) );
  IV U613 ( .A(n671), .Z(n676) );
  XOR U614 ( .A(n677), .B(n678), .Z(n671) );
  AND U615 ( .A(n203), .B(n670), .Z(n678) );
  XNOR U616 ( .A(n668), .B(n677), .Z(n670) );
  XNOR U617 ( .A(n679), .B(n680), .Z(n668) );
  AND U618 ( .A(n207), .B(n681), .Z(n680) );
  XOR U619 ( .A(p_input[131]), .B(n679), .Z(n681) );
  XOR U620 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(n682), .Z(
        n679) );
  AND U621 ( .A(n210), .B(n683), .Z(n682) );
  XOR U622 ( .A(n684), .B(n685), .Z(n677) );
  AND U623 ( .A(n214), .B(n686), .Z(n685) );
  XOR U624 ( .A(n687), .B(n688), .Z(n674) );
  AND U625 ( .A(n218), .B(n686), .Z(n688) );
  XNOR U626 ( .A(n689), .B(n687), .Z(n686) );
  IV U627 ( .A(n684), .Z(n689) );
  XOR U628 ( .A(n690), .B(n691), .Z(n684) );
  AND U629 ( .A(n221), .B(n683), .Z(n691) );
  XOR U630 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(n690), .Z(
        n683) );
  XOR U631 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .B(n692), .Z(
        n690) );
  AND U632 ( .A(n223), .B(n693), .Z(n692) );
  XOR U633 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n694), .Z(n687) );
  AND U634 ( .A(n226), .B(n693), .Z(n694) );
  XOR U635 ( .A(\knn_comb_/min_val_out[0][3] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .Z(n693) );
  XOR U636 ( .A(n695), .B(n696), .Z(o[34]) );
  XOR U637 ( .A(n697), .B(n698), .Z(o[33]) );
  XOR U638 ( .A(n699), .B(n700), .Z(o[32]) );
  XOR U639 ( .A(n73), .B(n701), .Z(o[31]) );
  AND U640 ( .A(n122), .B(n702), .Z(n73) );
  XOR U641 ( .A(n74), .B(n701), .Z(n702) );
  XOR U642 ( .A(n703), .B(n704), .Z(n701) );
  AND U643 ( .A(n142), .B(n705), .Z(n704) );
  XOR U644 ( .A(n706), .B(n3), .Z(n74) );
  AND U645 ( .A(n125), .B(n707), .Z(n3) );
  XOR U646 ( .A(n4), .B(n706), .Z(n707) );
  XOR U647 ( .A(n708), .B(n709), .Z(n4) );
  AND U648 ( .A(n130), .B(n710), .Z(n709) );
  XOR U649 ( .A(p_input[31]), .B(n708), .Z(n710) );
  XNOR U650 ( .A(n711), .B(n712), .Z(n708) );
  AND U651 ( .A(n134), .B(n713), .Z(n712) );
  XOR U652 ( .A(n714), .B(n715), .Z(n706) );
  AND U653 ( .A(n138), .B(n705), .Z(n715) );
  XNOR U654 ( .A(n716), .B(n703), .Z(n705) );
  XOR U655 ( .A(n717), .B(n718), .Z(n703) );
  AND U656 ( .A(n162), .B(n719), .Z(n718) );
  IV U657 ( .A(n714), .Z(n716) );
  XOR U658 ( .A(n720), .B(n721), .Z(n714) );
  AND U659 ( .A(n146), .B(n713), .Z(n721) );
  XNOR U660 ( .A(n711), .B(n720), .Z(n713) );
  XNOR U661 ( .A(n722), .B(n723), .Z(n711) );
  AND U662 ( .A(n150), .B(n724), .Z(n723) );
  XOR U663 ( .A(p_input[63]), .B(n722), .Z(n724) );
  XNOR U664 ( .A(n725), .B(n726), .Z(n722) );
  AND U665 ( .A(n154), .B(n727), .Z(n726) );
  XOR U666 ( .A(n728), .B(n729), .Z(n720) );
  AND U667 ( .A(n158), .B(n719), .Z(n729) );
  XNOR U668 ( .A(n730), .B(n717), .Z(n719) );
  XOR U669 ( .A(n731), .B(n732), .Z(n717) );
  AND U670 ( .A(n181), .B(n733), .Z(n732) );
  IV U671 ( .A(n728), .Z(n730) );
  XOR U672 ( .A(n734), .B(n735), .Z(n728) );
  AND U673 ( .A(n165), .B(n727), .Z(n735) );
  XNOR U674 ( .A(n725), .B(n734), .Z(n727) );
  XNOR U675 ( .A(n736), .B(n737), .Z(n725) );
  AND U676 ( .A(n169), .B(n738), .Z(n737) );
  XOR U677 ( .A(p_input[95]), .B(n736), .Z(n738) );
  XNOR U678 ( .A(n739), .B(n740), .Z(n736) );
  AND U679 ( .A(n173), .B(n741), .Z(n740) );
  XOR U680 ( .A(n742), .B(n743), .Z(n734) );
  AND U681 ( .A(n177), .B(n733), .Z(n743) );
  XNOR U682 ( .A(n744), .B(n731), .Z(n733) );
  XOR U683 ( .A(n745), .B(n746), .Z(n731) );
  AND U684 ( .A(n200), .B(n747), .Z(n746) );
  IV U685 ( .A(n742), .Z(n744) );
  XOR U686 ( .A(n748), .B(n749), .Z(n742) );
  AND U687 ( .A(n184), .B(n741), .Z(n749) );
  XNOR U688 ( .A(n739), .B(n748), .Z(n741) );
  XNOR U689 ( .A(n750), .B(n751), .Z(n739) );
  AND U690 ( .A(n188), .B(n752), .Z(n751) );
  XOR U691 ( .A(p_input[127]), .B(n750), .Z(n752) );
  XNOR U692 ( .A(n753), .B(n754), .Z(n750) );
  AND U693 ( .A(n192), .B(n755), .Z(n754) );
  XOR U694 ( .A(n756), .B(n757), .Z(n748) );
  AND U695 ( .A(n196), .B(n747), .Z(n757) );
  XNOR U696 ( .A(n758), .B(n745), .Z(n747) );
  XOR U697 ( .A(n759), .B(n760), .Z(n745) );
  AND U698 ( .A(n218), .B(n761), .Z(n760) );
  IV U699 ( .A(n756), .Z(n758) );
  XOR U700 ( .A(n762), .B(n763), .Z(n756) );
  AND U701 ( .A(n203), .B(n755), .Z(n763) );
  XNOR U702 ( .A(n753), .B(n762), .Z(n755) );
  XNOR U703 ( .A(n764), .B(n765), .Z(n753) );
  AND U704 ( .A(n207), .B(n766), .Z(n765) );
  XOR U705 ( .A(p_input[159]), .B(n764), .Z(n766) );
  XOR U706 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][31] ), .B(n767), .Z(
        n764) );
  AND U707 ( .A(n210), .B(n768), .Z(n767) );
  XOR U708 ( .A(n769), .B(n770), .Z(n762) );
  AND U709 ( .A(n214), .B(n761), .Z(n770) );
  XNOR U710 ( .A(n771), .B(n759), .Z(n761) );
  XOR U711 ( .A(\knn_comb_/min_val_out[0][31] ), .B(n772), .Z(n759) );
  AND U712 ( .A(n226), .B(n773), .Z(n772) );
  IV U713 ( .A(n769), .Z(n771) );
  XOR U714 ( .A(n774), .B(n775), .Z(n769) );
  AND U715 ( .A(n221), .B(n768), .Z(n775) );
  XOR U716 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][31] ), .B(n774), .Z(
        n768) );
  XOR U717 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .B(n776), .Z(
        n774) );
  AND U718 ( .A(n223), .B(n773), .Z(n776) );
  XOR U719 ( .A(n777), .B(n778), .Z(n773) );
  IV U720 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .Z(n778) );
  IV U721 ( .A(\knn_comb_/min_val_out[0][31] ), .Z(n777) );
  XOR U722 ( .A(n75), .B(n779), .Z(o[30]) );
  AND U723 ( .A(n122), .B(n780), .Z(n75) );
  XOR U724 ( .A(n76), .B(n779), .Z(n780) );
  XOR U725 ( .A(n781), .B(n782), .Z(n779) );
  AND U726 ( .A(n142), .B(n783), .Z(n782) );
  XOR U727 ( .A(n784), .B(n5), .Z(n76) );
  AND U728 ( .A(n125), .B(n785), .Z(n5) );
  XOR U729 ( .A(n6), .B(n784), .Z(n785) );
  XOR U730 ( .A(n786), .B(n787), .Z(n6) );
  AND U731 ( .A(n130), .B(n788), .Z(n787) );
  XOR U732 ( .A(p_input[30]), .B(n786), .Z(n788) );
  XNOR U733 ( .A(n789), .B(n790), .Z(n786) );
  AND U734 ( .A(n134), .B(n791), .Z(n790) );
  XOR U735 ( .A(n792), .B(n793), .Z(n784) );
  AND U736 ( .A(n138), .B(n783), .Z(n793) );
  XNOR U737 ( .A(n794), .B(n781), .Z(n783) );
  XOR U738 ( .A(n795), .B(n796), .Z(n781) );
  AND U739 ( .A(n162), .B(n797), .Z(n796) );
  IV U740 ( .A(n792), .Z(n794) );
  XOR U741 ( .A(n798), .B(n799), .Z(n792) );
  AND U742 ( .A(n146), .B(n791), .Z(n799) );
  XNOR U743 ( .A(n789), .B(n798), .Z(n791) );
  XNOR U744 ( .A(n800), .B(n801), .Z(n789) );
  AND U745 ( .A(n150), .B(n802), .Z(n801) );
  XOR U746 ( .A(p_input[62]), .B(n800), .Z(n802) );
  XNOR U747 ( .A(n803), .B(n804), .Z(n800) );
  AND U748 ( .A(n154), .B(n805), .Z(n804) );
  XOR U749 ( .A(n806), .B(n807), .Z(n798) );
  AND U750 ( .A(n158), .B(n797), .Z(n807) );
  XNOR U751 ( .A(n808), .B(n795), .Z(n797) );
  XOR U752 ( .A(n809), .B(n810), .Z(n795) );
  AND U753 ( .A(n181), .B(n811), .Z(n810) );
  IV U754 ( .A(n806), .Z(n808) );
  XOR U755 ( .A(n812), .B(n813), .Z(n806) );
  AND U756 ( .A(n165), .B(n805), .Z(n813) );
  XNOR U757 ( .A(n803), .B(n812), .Z(n805) );
  XNOR U758 ( .A(n814), .B(n815), .Z(n803) );
  AND U759 ( .A(n169), .B(n816), .Z(n815) );
  XOR U760 ( .A(p_input[94]), .B(n814), .Z(n816) );
  XNOR U761 ( .A(n817), .B(n818), .Z(n814) );
  AND U762 ( .A(n173), .B(n819), .Z(n818) );
  XOR U763 ( .A(n820), .B(n821), .Z(n812) );
  AND U764 ( .A(n177), .B(n811), .Z(n821) );
  XNOR U765 ( .A(n822), .B(n809), .Z(n811) );
  XOR U766 ( .A(n823), .B(n824), .Z(n809) );
  AND U767 ( .A(n200), .B(n825), .Z(n824) );
  IV U768 ( .A(n820), .Z(n822) );
  XOR U769 ( .A(n826), .B(n827), .Z(n820) );
  AND U770 ( .A(n184), .B(n819), .Z(n827) );
  XNOR U771 ( .A(n817), .B(n826), .Z(n819) );
  XNOR U772 ( .A(n828), .B(n829), .Z(n817) );
  AND U773 ( .A(n188), .B(n830), .Z(n829) );
  XOR U774 ( .A(p_input[126]), .B(n828), .Z(n830) );
  XNOR U775 ( .A(n831), .B(n832), .Z(n828) );
  AND U776 ( .A(n192), .B(n833), .Z(n832) );
  XOR U777 ( .A(n834), .B(n835), .Z(n826) );
  AND U778 ( .A(n196), .B(n825), .Z(n835) );
  XNOR U779 ( .A(n836), .B(n823), .Z(n825) );
  XOR U780 ( .A(n837), .B(n838), .Z(n823) );
  AND U781 ( .A(n218), .B(n839), .Z(n838) );
  IV U782 ( .A(n834), .Z(n836) );
  XOR U783 ( .A(n840), .B(n841), .Z(n834) );
  AND U784 ( .A(n203), .B(n833), .Z(n841) );
  XNOR U785 ( .A(n831), .B(n840), .Z(n833) );
  XNOR U786 ( .A(n842), .B(n843), .Z(n831) );
  AND U787 ( .A(n207), .B(n844), .Z(n843) );
  XOR U788 ( .A(p_input[158]), .B(n842), .Z(n844) );
  XOR U789 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][30] ), .B(n845), .Z(
        n842) );
  AND U790 ( .A(n210), .B(n846), .Z(n845) );
  XOR U791 ( .A(n847), .B(n848), .Z(n840) );
  AND U792 ( .A(n214), .B(n839), .Z(n848) );
  XNOR U793 ( .A(n849), .B(n837), .Z(n839) );
  XOR U794 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n850), .Z(n837) );
  AND U795 ( .A(n226), .B(n851), .Z(n850) );
  IV U796 ( .A(n847), .Z(n849) );
  XOR U797 ( .A(n852), .B(n853), .Z(n847) );
  AND U798 ( .A(n221), .B(n846), .Z(n853) );
  XOR U799 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][30] ), .B(n852), .Z(
        n846) );
  XOR U800 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .B(n854), .Z(
        n852) );
  AND U801 ( .A(n223), .B(n851), .Z(n854) );
  XOR U802 ( .A(n855), .B(n856), .Z(n851) );
  IV U803 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .Z(n856) );
  IV U804 ( .A(\knn_comb_/min_val_out[0][30] ), .Z(n855) );
  XOR U805 ( .A(n695), .B(n857), .Z(o[2]) );
  AND U806 ( .A(n122), .B(n858), .Z(n695) );
  XOR U807 ( .A(n696), .B(n857), .Z(n858) );
  XOR U808 ( .A(n859), .B(n860), .Z(n857) );
  AND U809 ( .A(n142), .B(n861), .Z(n860) );
  XOR U810 ( .A(n862), .B(n67), .Z(n696) );
  AND U811 ( .A(n125), .B(n863), .Z(n67) );
  XOR U812 ( .A(n68), .B(n862), .Z(n863) );
  XOR U813 ( .A(n864), .B(n865), .Z(n68) );
  AND U814 ( .A(n130), .B(n866), .Z(n865) );
  XOR U815 ( .A(p_input[2]), .B(n864), .Z(n866) );
  XNOR U816 ( .A(n867), .B(n868), .Z(n864) );
  AND U817 ( .A(n134), .B(n869), .Z(n868) );
  XOR U818 ( .A(n870), .B(n871), .Z(n862) );
  AND U819 ( .A(n138), .B(n861), .Z(n871) );
  XNOR U820 ( .A(n872), .B(n859), .Z(n861) );
  XOR U821 ( .A(n873), .B(n874), .Z(n859) );
  AND U822 ( .A(n162), .B(n875), .Z(n874) );
  IV U823 ( .A(n870), .Z(n872) );
  XOR U824 ( .A(n876), .B(n877), .Z(n870) );
  AND U825 ( .A(n146), .B(n869), .Z(n877) );
  XNOR U826 ( .A(n867), .B(n876), .Z(n869) );
  XNOR U827 ( .A(n878), .B(n879), .Z(n867) );
  AND U828 ( .A(n150), .B(n880), .Z(n879) );
  XOR U829 ( .A(p_input[34]), .B(n878), .Z(n880) );
  XNOR U830 ( .A(n881), .B(n882), .Z(n878) );
  AND U831 ( .A(n154), .B(n883), .Z(n882) );
  XOR U832 ( .A(n884), .B(n885), .Z(n876) );
  AND U833 ( .A(n158), .B(n875), .Z(n885) );
  XNOR U834 ( .A(n886), .B(n873), .Z(n875) );
  XOR U835 ( .A(n887), .B(n888), .Z(n873) );
  AND U836 ( .A(n181), .B(n889), .Z(n888) );
  IV U837 ( .A(n884), .Z(n886) );
  XOR U838 ( .A(n890), .B(n891), .Z(n884) );
  AND U839 ( .A(n165), .B(n883), .Z(n891) );
  XNOR U840 ( .A(n881), .B(n890), .Z(n883) );
  XNOR U841 ( .A(n892), .B(n893), .Z(n881) );
  AND U842 ( .A(n169), .B(n894), .Z(n893) );
  XOR U843 ( .A(p_input[66]), .B(n892), .Z(n894) );
  XNOR U844 ( .A(n895), .B(n896), .Z(n892) );
  AND U845 ( .A(n173), .B(n897), .Z(n896) );
  XOR U846 ( .A(n898), .B(n899), .Z(n890) );
  AND U847 ( .A(n177), .B(n889), .Z(n899) );
  XNOR U848 ( .A(n900), .B(n887), .Z(n889) );
  XOR U849 ( .A(n901), .B(n902), .Z(n887) );
  AND U850 ( .A(n200), .B(n903), .Z(n902) );
  IV U851 ( .A(n898), .Z(n900) );
  XOR U852 ( .A(n904), .B(n905), .Z(n898) );
  AND U853 ( .A(n184), .B(n897), .Z(n905) );
  XNOR U854 ( .A(n895), .B(n904), .Z(n897) );
  XNOR U855 ( .A(n906), .B(n907), .Z(n895) );
  AND U856 ( .A(n188), .B(n908), .Z(n907) );
  XOR U857 ( .A(p_input[98]), .B(n906), .Z(n908) );
  XNOR U858 ( .A(n909), .B(n910), .Z(n906) );
  AND U859 ( .A(n192), .B(n911), .Z(n910) );
  XOR U860 ( .A(n912), .B(n913), .Z(n904) );
  AND U861 ( .A(n196), .B(n903), .Z(n913) );
  XNOR U862 ( .A(n914), .B(n901), .Z(n903) );
  XOR U863 ( .A(n915), .B(n916), .Z(n901) );
  AND U864 ( .A(n218), .B(n917), .Z(n916) );
  IV U865 ( .A(n912), .Z(n914) );
  XOR U866 ( .A(n918), .B(n919), .Z(n912) );
  AND U867 ( .A(n203), .B(n911), .Z(n919) );
  XNOR U868 ( .A(n909), .B(n918), .Z(n911) );
  XNOR U869 ( .A(n920), .B(n921), .Z(n909) );
  AND U870 ( .A(n207), .B(n922), .Z(n921) );
  XOR U871 ( .A(p_input[130]), .B(n920), .Z(n922) );
  XOR U872 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n923), .Z(
        n920) );
  AND U873 ( .A(n210), .B(n924), .Z(n923) );
  XOR U874 ( .A(n925), .B(n926), .Z(n918) );
  AND U875 ( .A(n214), .B(n917), .Z(n926) );
  XNOR U876 ( .A(n927), .B(n915), .Z(n917) );
  XOR U877 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n928), .Z(n915) );
  AND U878 ( .A(n226), .B(n929), .Z(n928) );
  IV U879 ( .A(n925), .Z(n927) );
  XOR U880 ( .A(n930), .B(n931), .Z(n925) );
  AND U881 ( .A(n221), .B(n924), .Z(n931) );
  XOR U882 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n930), .Z(
        n924) );
  XOR U883 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .B(n932), .Z(
        n930) );
  AND U884 ( .A(n223), .B(n929), .Z(n932) );
  XOR U885 ( .A(\knn_comb_/min_val_out[0][2] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n929) );
  XOR U886 ( .A(n77), .B(n933), .Z(o[29]) );
  AND U887 ( .A(n122), .B(n934), .Z(n77) );
  XOR U888 ( .A(n78), .B(n933), .Z(n934) );
  XOR U889 ( .A(n935), .B(n936), .Z(n933) );
  AND U890 ( .A(n142), .B(n937), .Z(n936) );
  XOR U891 ( .A(n938), .B(n7), .Z(n78) );
  AND U892 ( .A(n125), .B(n939), .Z(n7) );
  XOR U893 ( .A(n8), .B(n938), .Z(n939) );
  XOR U894 ( .A(n940), .B(n941), .Z(n8) );
  AND U895 ( .A(n130), .B(n942), .Z(n941) );
  XOR U896 ( .A(p_input[29]), .B(n940), .Z(n942) );
  XNOR U897 ( .A(n943), .B(n944), .Z(n940) );
  AND U898 ( .A(n134), .B(n945), .Z(n944) );
  XOR U899 ( .A(n946), .B(n947), .Z(n938) );
  AND U900 ( .A(n138), .B(n937), .Z(n947) );
  XNOR U901 ( .A(n948), .B(n935), .Z(n937) );
  XOR U902 ( .A(n949), .B(n950), .Z(n935) );
  AND U903 ( .A(n162), .B(n951), .Z(n950) );
  IV U904 ( .A(n946), .Z(n948) );
  XOR U905 ( .A(n952), .B(n953), .Z(n946) );
  AND U906 ( .A(n146), .B(n945), .Z(n953) );
  XNOR U907 ( .A(n943), .B(n952), .Z(n945) );
  XNOR U908 ( .A(n954), .B(n955), .Z(n943) );
  AND U909 ( .A(n150), .B(n956), .Z(n955) );
  XOR U910 ( .A(p_input[61]), .B(n954), .Z(n956) );
  XNOR U911 ( .A(n957), .B(n958), .Z(n954) );
  AND U912 ( .A(n154), .B(n959), .Z(n958) );
  XOR U913 ( .A(n960), .B(n961), .Z(n952) );
  AND U914 ( .A(n158), .B(n951), .Z(n961) );
  XNOR U915 ( .A(n962), .B(n949), .Z(n951) );
  XOR U916 ( .A(n963), .B(n964), .Z(n949) );
  AND U917 ( .A(n181), .B(n965), .Z(n964) );
  IV U918 ( .A(n960), .Z(n962) );
  XOR U919 ( .A(n966), .B(n967), .Z(n960) );
  AND U920 ( .A(n165), .B(n959), .Z(n967) );
  XNOR U921 ( .A(n957), .B(n966), .Z(n959) );
  XNOR U922 ( .A(n968), .B(n969), .Z(n957) );
  AND U923 ( .A(n169), .B(n970), .Z(n969) );
  XOR U924 ( .A(p_input[93]), .B(n968), .Z(n970) );
  XNOR U925 ( .A(n971), .B(n972), .Z(n968) );
  AND U926 ( .A(n173), .B(n973), .Z(n972) );
  XOR U927 ( .A(n974), .B(n975), .Z(n966) );
  AND U928 ( .A(n177), .B(n965), .Z(n975) );
  XNOR U929 ( .A(n976), .B(n963), .Z(n965) );
  XOR U930 ( .A(n977), .B(n978), .Z(n963) );
  AND U931 ( .A(n200), .B(n979), .Z(n978) );
  IV U932 ( .A(n974), .Z(n976) );
  XOR U933 ( .A(n980), .B(n981), .Z(n974) );
  AND U934 ( .A(n184), .B(n973), .Z(n981) );
  XNOR U935 ( .A(n971), .B(n980), .Z(n973) );
  XNOR U936 ( .A(n982), .B(n983), .Z(n971) );
  AND U937 ( .A(n188), .B(n984), .Z(n983) );
  XOR U938 ( .A(p_input[125]), .B(n982), .Z(n984) );
  XNOR U939 ( .A(n985), .B(n986), .Z(n982) );
  AND U940 ( .A(n192), .B(n987), .Z(n986) );
  XOR U941 ( .A(n988), .B(n989), .Z(n980) );
  AND U942 ( .A(n196), .B(n979), .Z(n989) );
  XNOR U943 ( .A(n990), .B(n977), .Z(n979) );
  XOR U944 ( .A(n991), .B(n992), .Z(n977) );
  AND U945 ( .A(n218), .B(n993), .Z(n992) );
  IV U946 ( .A(n988), .Z(n990) );
  XOR U947 ( .A(n994), .B(n995), .Z(n988) );
  AND U948 ( .A(n203), .B(n987), .Z(n995) );
  XNOR U949 ( .A(n985), .B(n994), .Z(n987) );
  XNOR U950 ( .A(n996), .B(n997), .Z(n985) );
  AND U951 ( .A(n207), .B(n998), .Z(n997) );
  XOR U952 ( .A(p_input[157]), .B(n996), .Z(n998) );
  XOR U953 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][29] ), .B(n999), .Z(
        n996) );
  AND U954 ( .A(n210), .B(n1000), .Z(n999) );
  XOR U955 ( .A(n1001), .B(n1002), .Z(n994) );
  AND U956 ( .A(n214), .B(n993), .Z(n1002) );
  XNOR U957 ( .A(n1003), .B(n991), .Z(n993) );
  XOR U958 ( .A(\knn_comb_/min_val_out[0][29] ), .B(n1004), .Z(n991) );
  AND U959 ( .A(n226), .B(n1005), .Z(n1004) );
  IV U960 ( .A(n1001), .Z(n1003) );
  XOR U961 ( .A(n1006), .B(n1007), .Z(n1001) );
  AND U962 ( .A(n221), .B(n1000), .Z(n1007) );
  XOR U963 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][29] ), .B(n1006), 
        .Z(n1000) );
  XOR U964 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .B(n1008), 
        .Z(n1006) );
  AND U965 ( .A(n223), .B(n1005), .Z(n1008) );
  XOR U966 ( .A(\knn_comb_/min_val_out[0][29] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .Z(n1005) );
  XOR U967 ( .A(n79), .B(n1009), .Z(o[28]) );
  AND U968 ( .A(n122), .B(n1010), .Z(n79) );
  XOR U969 ( .A(n80), .B(n1009), .Z(n1010) );
  XOR U970 ( .A(n1011), .B(n1012), .Z(n1009) );
  AND U971 ( .A(n142), .B(n1013), .Z(n1012) );
  XOR U972 ( .A(n1014), .B(n9), .Z(n80) );
  AND U973 ( .A(n125), .B(n1015), .Z(n9) );
  XOR U974 ( .A(n10), .B(n1014), .Z(n1015) );
  XOR U975 ( .A(n1016), .B(n1017), .Z(n10) );
  AND U976 ( .A(n130), .B(n1018), .Z(n1017) );
  XOR U977 ( .A(p_input[28]), .B(n1016), .Z(n1018) );
  XNOR U978 ( .A(n1019), .B(n1020), .Z(n1016) );
  AND U979 ( .A(n134), .B(n1021), .Z(n1020) );
  XOR U980 ( .A(n1022), .B(n1023), .Z(n1014) );
  AND U981 ( .A(n138), .B(n1013), .Z(n1023) );
  XNOR U982 ( .A(n1024), .B(n1011), .Z(n1013) );
  XOR U983 ( .A(n1025), .B(n1026), .Z(n1011) );
  AND U984 ( .A(n162), .B(n1027), .Z(n1026) );
  IV U985 ( .A(n1022), .Z(n1024) );
  XOR U986 ( .A(n1028), .B(n1029), .Z(n1022) );
  AND U987 ( .A(n146), .B(n1021), .Z(n1029) );
  XNOR U988 ( .A(n1019), .B(n1028), .Z(n1021) );
  XNOR U989 ( .A(n1030), .B(n1031), .Z(n1019) );
  AND U990 ( .A(n150), .B(n1032), .Z(n1031) );
  XOR U991 ( .A(p_input[60]), .B(n1030), .Z(n1032) );
  XNOR U992 ( .A(n1033), .B(n1034), .Z(n1030) );
  AND U993 ( .A(n154), .B(n1035), .Z(n1034) );
  XOR U994 ( .A(n1036), .B(n1037), .Z(n1028) );
  AND U995 ( .A(n158), .B(n1027), .Z(n1037) );
  XNOR U996 ( .A(n1038), .B(n1025), .Z(n1027) );
  XOR U997 ( .A(n1039), .B(n1040), .Z(n1025) );
  AND U998 ( .A(n181), .B(n1041), .Z(n1040) );
  IV U999 ( .A(n1036), .Z(n1038) );
  XOR U1000 ( .A(n1042), .B(n1043), .Z(n1036) );
  AND U1001 ( .A(n165), .B(n1035), .Z(n1043) );
  XNOR U1002 ( .A(n1033), .B(n1042), .Z(n1035) );
  XNOR U1003 ( .A(n1044), .B(n1045), .Z(n1033) );
  AND U1004 ( .A(n169), .B(n1046), .Z(n1045) );
  XOR U1005 ( .A(p_input[92]), .B(n1044), .Z(n1046) );
  XNOR U1006 ( .A(n1047), .B(n1048), .Z(n1044) );
  AND U1007 ( .A(n173), .B(n1049), .Z(n1048) );
  XOR U1008 ( .A(n1050), .B(n1051), .Z(n1042) );
  AND U1009 ( .A(n177), .B(n1041), .Z(n1051) );
  XNOR U1010 ( .A(n1052), .B(n1039), .Z(n1041) );
  XOR U1011 ( .A(n1053), .B(n1054), .Z(n1039) );
  AND U1012 ( .A(n200), .B(n1055), .Z(n1054) );
  IV U1013 ( .A(n1050), .Z(n1052) );
  XOR U1014 ( .A(n1056), .B(n1057), .Z(n1050) );
  AND U1015 ( .A(n184), .B(n1049), .Z(n1057) );
  XNOR U1016 ( .A(n1047), .B(n1056), .Z(n1049) );
  XNOR U1017 ( .A(n1058), .B(n1059), .Z(n1047) );
  AND U1018 ( .A(n188), .B(n1060), .Z(n1059) );
  XOR U1019 ( .A(p_input[124]), .B(n1058), .Z(n1060) );
  XNOR U1020 ( .A(n1061), .B(n1062), .Z(n1058) );
  AND U1021 ( .A(n192), .B(n1063), .Z(n1062) );
  XOR U1022 ( .A(n1064), .B(n1065), .Z(n1056) );
  AND U1023 ( .A(n196), .B(n1055), .Z(n1065) );
  XNOR U1024 ( .A(n1066), .B(n1053), .Z(n1055) );
  XOR U1025 ( .A(n1067), .B(n1068), .Z(n1053) );
  AND U1026 ( .A(n218), .B(n1069), .Z(n1068) );
  IV U1027 ( .A(n1064), .Z(n1066) );
  XOR U1028 ( .A(n1070), .B(n1071), .Z(n1064) );
  AND U1029 ( .A(n203), .B(n1063), .Z(n1071) );
  XNOR U1030 ( .A(n1061), .B(n1070), .Z(n1063) );
  XNOR U1031 ( .A(n1072), .B(n1073), .Z(n1061) );
  AND U1032 ( .A(n207), .B(n1074), .Z(n1073) );
  XOR U1033 ( .A(p_input[156]), .B(n1072), .Z(n1074) );
  XOR U1034 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][28] ), .B(n1075), 
        .Z(n1072) );
  AND U1035 ( .A(n210), .B(n1076), .Z(n1075) );
  XOR U1036 ( .A(n1077), .B(n1078), .Z(n1070) );
  AND U1037 ( .A(n214), .B(n1069), .Z(n1078) );
  XNOR U1038 ( .A(n1079), .B(n1067), .Z(n1069) );
  XOR U1039 ( .A(\knn_comb_/min_val_out[0][28] ), .B(n1080), .Z(n1067) );
  AND U1040 ( .A(n226), .B(n1081), .Z(n1080) );
  IV U1041 ( .A(n1077), .Z(n1079) );
  XOR U1042 ( .A(n1082), .B(n1083), .Z(n1077) );
  AND U1043 ( .A(n221), .B(n1076), .Z(n1083) );
  XOR U1044 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][28] ), .B(n1082), 
        .Z(n1076) );
  XOR U1045 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .B(n1084), 
        .Z(n1082) );
  AND U1046 ( .A(n223), .B(n1081), .Z(n1084) );
  XOR U1047 ( .A(\knn_comb_/min_val_out[0][28] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .Z(n1081) );
  XOR U1048 ( .A(n83), .B(n1085), .Z(o[27]) );
  AND U1049 ( .A(n122), .B(n1086), .Z(n83) );
  XOR U1050 ( .A(n84), .B(n1085), .Z(n1086) );
  XOR U1051 ( .A(n1087), .B(n1088), .Z(n1085) );
  AND U1052 ( .A(n142), .B(n1089), .Z(n1088) );
  XOR U1053 ( .A(n1090), .B(n11), .Z(n84) );
  AND U1054 ( .A(n125), .B(n1091), .Z(n11) );
  XOR U1055 ( .A(n12), .B(n1090), .Z(n1091) );
  XOR U1056 ( .A(n1092), .B(n1093), .Z(n12) );
  AND U1057 ( .A(n130), .B(n1094), .Z(n1093) );
  XOR U1058 ( .A(p_input[27]), .B(n1092), .Z(n1094) );
  XNOR U1059 ( .A(n1095), .B(n1096), .Z(n1092) );
  AND U1060 ( .A(n134), .B(n1097), .Z(n1096) );
  XOR U1061 ( .A(n1098), .B(n1099), .Z(n1090) );
  AND U1062 ( .A(n138), .B(n1089), .Z(n1099) );
  XNOR U1063 ( .A(n1100), .B(n1087), .Z(n1089) );
  XOR U1064 ( .A(n1101), .B(n1102), .Z(n1087) );
  AND U1065 ( .A(n162), .B(n1103), .Z(n1102) );
  IV U1066 ( .A(n1098), .Z(n1100) );
  XOR U1067 ( .A(n1104), .B(n1105), .Z(n1098) );
  AND U1068 ( .A(n146), .B(n1097), .Z(n1105) );
  XNOR U1069 ( .A(n1095), .B(n1104), .Z(n1097) );
  XNOR U1070 ( .A(n1106), .B(n1107), .Z(n1095) );
  AND U1071 ( .A(n150), .B(n1108), .Z(n1107) );
  XOR U1072 ( .A(p_input[59]), .B(n1106), .Z(n1108) );
  XNOR U1073 ( .A(n1109), .B(n1110), .Z(n1106) );
  AND U1074 ( .A(n154), .B(n1111), .Z(n1110) );
  XOR U1075 ( .A(n1112), .B(n1113), .Z(n1104) );
  AND U1076 ( .A(n158), .B(n1103), .Z(n1113) );
  XNOR U1077 ( .A(n1114), .B(n1101), .Z(n1103) );
  XOR U1078 ( .A(n1115), .B(n1116), .Z(n1101) );
  AND U1079 ( .A(n181), .B(n1117), .Z(n1116) );
  IV U1080 ( .A(n1112), .Z(n1114) );
  XOR U1081 ( .A(n1118), .B(n1119), .Z(n1112) );
  AND U1082 ( .A(n165), .B(n1111), .Z(n1119) );
  XNOR U1083 ( .A(n1109), .B(n1118), .Z(n1111) );
  XNOR U1084 ( .A(n1120), .B(n1121), .Z(n1109) );
  AND U1085 ( .A(n169), .B(n1122), .Z(n1121) );
  XOR U1086 ( .A(p_input[91]), .B(n1120), .Z(n1122) );
  XNOR U1087 ( .A(n1123), .B(n1124), .Z(n1120) );
  AND U1088 ( .A(n173), .B(n1125), .Z(n1124) );
  XOR U1089 ( .A(n1126), .B(n1127), .Z(n1118) );
  AND U1090 ( .A(n177), .B(n1117), .Z(n1127) );
  XNOR U1091 ( .A(n1128), .B(n1115), .Z(n1117) );
  XOR U1092 ( .A(n1129), .B(n1130), .Z(n1115) );
  AND U1093 ( .A(n200), .B(n1131), .Z(n1130) );
  IV U1094 ( .A(n1126), .Z(n1128) );
  XOR U1095 ( .A(n1132), .B(n1133), .Z(n1126) );
  AND U1096 ( .A(n184), .B(n1125), .Z(n1133) );
  XNOR U1097 ( .A(n1123), .B(n1132), .Z(n1125) );
  XNOR U1098 ( .A(n1134), .B(n1135), .Z(n1123) );
  AND U1099 ( .A(n188), .B(n1136), .Z(n1135) );
  XOR U1100 ( .A(p_input[123]), .B(n1134), .Z(n1136) );
  XNOR U1101 ( .A(n1137), .B(n1138), .Z(n1134) );
  AND U1102 ( .A(n192), .B(n1139), .Z(n1138) );
  XOR U1103 ( .A(n1140), .B(n1141), .Z(n1132) );
  AND U1104 ( .A(n196), .B(n1131), .Z(n1141) );
  XNOR U1105 ( .A(n1142), .B(n1129), .Z(n1131) );
  XOR U1106 ( .A(n1143), .B(n1144), .Z(n1129) );
  AND U1107 ( .A(n218), .B(n1145), .Z(n1144) );
  IV U1108 ( .A(n1140), .Z(n1142) );
  XOR U1109 ( .A(n1146), .B(n1147), .Z(n1140) );
  AND U1110 ( .A(n203), .B(n1139), .Z(n1147) );
  XNOR U1111 ( .A(n1137), .B(n1146), .Z(n1139) );
  XNOR U1112 ( .A(n1148), .B(n1149), .Z(n1137) );
  AND U1113 ( .A(n207), .B(n1150), .Z(n1149) );
  XOR U1114 ( .A(p_input[155]), .B(n1148), .Z(n1150) );
  XOR U1115 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][27] ), .B(n1151), 
        .Z(n1148) );
  AND U1116 ( .A(n210), .B(n1152), .Z(n1151) );
  XOR U1117 ( .A(n1153), .B(n1154), .Z(n1146) );
  AND U1118 ( .A(n214), .B(n1145), .Z(n1154) );
  XNOR U1119 ( .A(n1155), .B(n1143), .Z(n1145) );
  XOR U1120 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n1156), .Z(n1143) );
  AND U1121 ( .A(n226), .B(n1157), .Z(n1156) );
  IV U1122 ( .A(n1153), .Z(n1155) );
  XOR U1123 ( .A(n1158), .B(n1159), .Z(n1153) );
  AND U1124 ( .A(n221), .B(n1152), .Z(n1159) );
  XOR U1125 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][27] ), .B(n1158), 
        .Z(n1152) );
  XOR U1126 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .B(n1160), 
        .Z(n1158) );
  AND U1127 ( .A(n223), .B(n1157), .Z(n1160) );
  XOR U1128 ( .A(n1161), .B(n1162), .Z(n1157) );
  IV U1129 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .Z(n1162) );
  IV U1130 ( .A(\knn_comb_/min_val_out[0][27] ), .Z(n1161) );
  XOR U1131 ( .A(n85), .B(n1163), .Z(o[26]) );
  AND U1132 ( .A(n122), .B(n1164), .Z(n85) );
  XOR U1133 ( .A(n86), .B(n1163), .Z(n1164) );
  XOR U1134 ( .A(n1165), .B(n1166), .Z(n1163) );
  AND U1135 ( .A(n142), .B(n1167), .Z(n1166) );
  XOR U1136 ( .A(n1168), .B(n13), .Z(n86) );
  AND U1137 ( .A(n125), .B(n1169), .Z(n13) );
  XOR U1138 ( .A(n14), .B(n1168), .Z(n1169) );
  XOR U1139 ( .A(n1170), .B(n1171), .Z(n14) );
  AND U1140 ( .A(n130), .B(n1172), .Z(n1171) );
  XOR U1141 ( .A(p_input[26]), .B(n1170), .Z(n1172) );
  XNOR U1142 ( .A(n1173), .B(n1174), .Z(n1170) );
  AND U1143 ( .A(n134), .B(n1175), .Z(n1174) );
  XOR U1144 ( .A(n1176), .B(n1177), .Z(n1168) );
  AND U1145 ( .A(n138), .B(n1167), .Z(n1177) );
  XNOR U1146 ( .A(n1178), .B(n1165), .Z(n1167) );
  XOR U1147 ( .A(n1179), .B(n1180), .Z(n1165) );
  AND U1148 ( .A(n162), .B(n1181), .Z(n1180) );
  IV U1149 ( .A(n1176), .Z(n1178) );
  XOR U1150 ( .A(n1182), .B(n1183), .Z(n1176) );
  AND U1151 ( .A(n146), .B(n1175), .Z(n1183) );
  XNOR U1152 ( .A(n1173), .B(n1182), .Z(n1175) );
  XNOR U1153 ( .A(n1184), .B(n1185), .Z(n1173) );
  AND U1154 ( .A(n150), .B(n1186), .Z(n1185) );
  XOR U1155 ( .A(p_input[58]), .B(n1184), .Z(n1186) );
  XNOR U1156 ( .A(n1187), .B(n1188), .Z(n1184) );
  AND U1157 ( .A(n154), .B(n1189), .Z(n1188) );
  XOR U1158 ( .A(n1190), .B(n1191), .Z(n1182) );
  AND U1159 ( .A(n158), .B(n1181), .Z(n1191) );
  XNOR U1160 ( .A(n1192), .B(n1179), .Z(n1181) );
  XOR U1161 ( .A(n1193), .B(n1194), .Z(n1179) );
  AND U1162 ( .A(n181), .B(n1195), .Z(n1194) );
  IV U1163 ( .A(n1190), .Z(n1192) );
  XOR U1164 ( .A(n1196), .B(n1197), .Z(n1190) );
  AND U1165 ( .A(n165), .B(n1189), .Z(n1197) );
  XNOR U1166 ( .A(n1187), .B(n1196), .Z(n1189) );
  XNOR U1167 ( .A(n1198), .B(n1199), .Z(n1187) );
  AND U1168 ( .A(n169), .B(n1200), .Z(n1199) );
  XOR U1169 ( .A(p_input[90]), .B(n1198), .Z(n1200) );
  XNOR U1170 ( .A(n1201), .B(n1202), .Z(n1198) );
  AND U1171 ( .A(n173), .B(n1203), .Z(n1202) );
  XOR U1172 ( .A(n1204), .B(n1205), .Z(n1196) );
  AND U1173 ( .A(n177), .B(n1195), .Z(n1205) );
  XNOR U1174 ( .A(n1206), .B(n1193), .Z(n1195) );
  XOR U1175 ( .A(n1207), .B(n1208), .Z(n1193) );
  AND U1176 ( .A(n200), .B(n1209), .Z(n1208) );
  IV U1177 ( .A(n1204), .Z(n1206) );
  XOR U1178 ( .A(n1210), .B(n1211), .Z(n1204) );
  AND U1179 ( .A(n184), .B(n1203), .Z(n1211) );
  XNOR U1180 ( .A(n1201), .B(n1210), .Z(n1203) );
  XNOR U1181 ( .A(n1212), .B(n1213), .Z(n1201) );
  AND U1182 ( .A(n188), .B(n1214), .Z(n1213) );
  XOR U1183 ( .A(p_input[122]), .B(n1212), .Z(n1214) );
  XNOR U1184 ( .A(n1215), .B(n1216), .Z(n1212) );
  AND U1185 ( .A(n192), .B(n1217), .Z(n1216) );
  XOR U1186 ( .A(n1218), .B(n1219), .Z(n1210) );
  AND U1187 ( .A(n196), .B(n1209), .Z(n1219) );
  XNOR U1188 ( .A(n1220), .B(n1207), .Z(n1209) );
  XOR U1189 ( .A(n1221), .B(n1222), .Z(n1207) );
  AND U1190 ( .A(n218), .B(n1223), .Z(n1222) );
  IV U1191 ( .A(n1218), .Z(n1220) );
  XOR U1192 ( .A(n1224), .B(n1225), .Z(n1218) );
  AND U1193 ( .A(n203), .B(n1217), .Z(n1225) );
  XNOR U1194 ( .A(n1215), .B(n1224), .Z(n1217) );
  XNOR U1195 ( .A(n1226), .B(n1227), .Z(n1215) );
  AND U1196 ( .A(n207), .B(n1228), .Z(n1227) );
  XOR U1197 ( .A(p_input[154]), .B(n1226), .Z(n1228) );
  XOR U1198 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][26] ), .B(n1229), 
        .Z(n1226) );
  AND U1199 ( .A(n210), .B(n1230), .Z(n1229) );
  XOR U1200 ( .A(n1231), .B(n1232), .Z(n1224) );
  AND U1201 ( .A(n214), .B(n1223), .Z(n1232) );
  XNOR U1202 ( .A(n1233), .B(n1221), .Z(n1223) );
  XOR U1203 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n1234), .Z(n1221) );
  AND U1204 ( .A(n226), .B(n1235), .Z(n1234) );
  IV U1205 ( .A(n1231), .Z(n1233) );
  XOR U1206 ( .A(n1236), .B(n1237), .Z(n1231) );
  AND U1207 ( .A(n221), .B(n1230), .Z(n1237) );
  XOR U1208 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][26] ), .B(n1236), 
        .Z(n1230) );
  XOR U1209 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .B(n1238), 
        .Z(n1236) );
  AND U1210 ( .A(n223), .B(n1235), .Z(n1238) );
  XOR U1211 ( .A(\knn_comb_/min_val_out[0][26] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .Z(n1235) );
  XOR U1212 ( .A(n87), .B(n1239), .Z(o[25]) );
  AND U1213 ( .A(n122), .B(n1240), .Z(n87) );
  XOR U1214 ( .A(n88), .B(n1239), .Z(n1240) );
  XOR U1215 ( .A(n1241), .B(n1242), .Z(n1239) );
  AND U1216 ( .A(n142), .B(n1243), .Z(n1242) );
  XOR U1217 ( .A(n1244), .B(n17), .Z(n88) );
  AND U1218 ( .A(n125), .B(n1245), .Z(n17) );
  XOR U1219 ( .A(n18), .B(n1244), .Z(n1245) );
  XOR U1220 ( .A(n1246), .B(n1247), .Z(n18) );
  AND U1221 ( .A(n130), .B(n1248), .Z(n1247) );
  XOR U1222 ( .A(p_input[25]), .B(n1246), .Z(n1248) );
  XNOR U1223 ( .A(n1249), .B(n1250), .Z(n1246) );
  AND U1224 ( .A(n134), .B(n1251), .Z(n1250) );
  XOR U1225 ( .A(n1252), .B(n1253), .Z(n1244) );
  AND U1226 ( .A(n138), .B(n1243), .Z(n1253) );
  XNOR U1227 ( .A(n1254), .B(n1241), .Z(n1243) );
  XOR U1228 ( .A(n1255), .B(n1256), .Z(n1241) );
  AND U1229 ( .A(n162), .B(n1257), .Z(n1256) );
  IV U1230 ( .A(n1252), .Z(n1254) );
  XOR U1231 ( .A(n1258), .B(n1259), .Z(n1252) );
  AND U1232 ( .A(n146), .B(n1251), .Z(n1259) );
  XNOR U1233 ( .A(n1249), .B(n1258), .Z(n1251) );
  XNOR U1234 ( .A(n1260), .B(n1261), .Z(n1249) );
  AND U1235 ( .A(n150), .B(n1262), .Z(n1261) );
  XOR U1236 ( .A(p_input[57]), .B(n1260), .Z(n1262) );
  XNOR U1237 ( .A(n1263), .B(n1264), .Z(n1260) );
  AND U1238 ( .A(n154), .B(n1265), .Z(n1264) );
  XOR U1239 ( .A(n1266), .B(n1267), .Z(n1258) );
  AND U1240 ( .A(n158), .B(n1257), .Z(n1267) );
  XNOR U1241 ( .A(n1268), .B(n1255), .Z(n1257) );
  XOR U1242 ( .A(n1269), .B(n1270), .Z(n1255) );
  AND U1243 ( .A(n181), .B(n1271), .Z(n1270) );
  IV U1244 ( .A(n1266), .Z(n1268) );
  XOR U1245 ( .A(n1272), .B(n1273), .Z(n1266) );
  AND U1246 ( .A(n165), .B(n1265), .Z(n1273) );
  XNOR U1247 ( .A(n1263), .B(n1272), .Z(n1265) );
  XNOR U1248 ( .A(n1274), .B(n1275), .Z(n1263) );
  AND U1249 ( .A(n169), .B(n1276), .Z(n1275) );
  XOR U1250 ( .A(p_input[89]), .B(n1274), .Z(n1276) );
  XNOR U1251 ( .A(n1277), .B(n1278), .Z(n1274) );
  AND U1252 ( .A(n173), .B(n1279), .Z(n1278) );
  XOR U1253 ( .A(n1280), .B(n1281), .Z(n1272) );
  AND U1254 ( .A(n177), .B(n1271), .Z(n1281) );
  XNOR U1255 ( .A(n1282), .B(n1269), .Z(n1271) );
  XOR U1256 ( .A(n1283), .B(n1284), .Z(n1269) );
  AND U1257 ( .A(n200), .B(n1285), .Z(n1284) );
  IV U1258 ( .A(n1280), .Z(n1282) );
  XOR U1259 ( .A(n1286), .B(n1287), .Z(n1280) );
  AND U1260 ( .A(n184), .B(n1279), .Z(n1287) );
  XNOR U1261 ( .A(n1277), .B(n1286), .Z(n1279) );
  XNOR U1262 ( .A(n1288), .B(n1289), .Z(n1277) );
  AND U1263 ( .A(n188), .B(n1290), .Z(n1289) );
  XOR U1264 ( .A(p_input[121]), .B(n1288), .Z(n1290) );
  XNOR U1265 ( .A(n1291), .B(n1292), .Z(n1288) );
  AND U1266 ( .A(n192), .B(n1293), .Z(n1292) );
  XOR U1267 ( .A(n1294), .B(n1295), .Z(n1286) );
  AND U1268 ( .A(n196), .B(n1285), .Z(n1295) );
  XNOR U1269 ( .A(n1296), .B(n1283), .Z(n1285) );
  XOR U1270 ( .A(n1297), .B(n1298), .Z(n1283) );
  AND U1271 ( .A(n218), .B(n1299), .Z(n1298) );
  IV U1272 ( .A(n1294), .Z(n1296) );
  XOR U1273 ( .A(n1300), .B(n1301), .Z(n1294) );
  AND U1274 ( .A(n203), .B(n1293), .Z(n1301) );
  XNOR U1275 ( .A(n1291), .B(n1300), .Z(n1293) );
  XNOR U1276 ( .A(n1302), .B(n1303), .Z(n1291) );
  AND U1277 ( .A(n207), .B(n1304), .Z(n1303) );
  XOR U1278 ( .A(p_input[153]), .B(n1302), .Z(n1304) );
  XOR U1279 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][25] ), .B(n1305), 
        .Z(n1302) );
  AND U1280 ( .A(n210), .B(n1306), .Z(n1305) );
  XOR U1281 ( .A(n1307), .B(n1308), .Z(n1300) );
  AND U1282 ( .A(n214), .B(n1299), .Z(n1308) );
  XNOR U1283 ( .A(n1309), .B(n1297), .Z(n1299) );
  XOR U1284 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n1310), .Z(n1297) );
  AND U1285 ( .A(n226), .B(n1311), .Z(n1310) );
  IV U1286 ( .A(n1307), .Z(n1309) );
  XOR U1287 ( .A(n1312), .B(n1313), .Z(n1307) );
  AND U1288 ( .A(n221), .B(n1306), .Z(n1313) );
  XOR U1289 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][25] ), .B(n1312), 
        .Z(n1306) );
  XOR U1290 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .B(n1314), 
        .Z(n1312) );
  AND U1291 ( .A(n223), .B(n1311), .Z(n1314) );
  XOR U1292 ( .A(\knn_comb_/min_val_out[0][25] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .Z(n1311) );
  XOR U1293 ( .A(n89), .B(n1315), .Z(o[24]) );
  AND U1294 ( .A(n122), .B(n1316), .Z(n89) );
  XOR U1295 ( .A(n90), .B(n1315), .Z(n1316) );
  XOR U1296 ( .A(n1317), .B(n1318), .Z(n1315) );
  AND U1297 ( .A(n142), .B(n1319), .Z(n1318) );
  XOR U1298 ( .A(n1320), .B(n19), .Z(n90) );
  AND U1299 ( .A(n125), .B(n1321), .Z(n19) );
  XOR U1300 ( .A(n20), .B(n1320), .Z(n1321) );
  XOR U1301 ( .A(n1322), .B(n1323), .Z(n20) );
  AND U1302 ( .A(n130), .B(n1324), .Z(n1323) );
  XOR U1303 ( .A(p_input[24]), .B(n1322), .Z(n1324) );
  XNOR U1304 ( .A(n1325), .B(n1326), .Z(n1322) );
  AND U1305 ( .A(n134), .B(n1327), .Z(n1326) );
  XOR U1306 ( .A(n1328), .B(n1329), .Z(n1320) );
  AND U1307 ( .A(n138), .B(n1319), .Z(n1329) );
  XNOR U1308 ( .A(n1330), .B(n1317), .Z(n1319) );
  XOR U1309 ( .A(n1331), .B(n1332), .Z(n1317) );
  AND U1310 ( .A(n162), .B(n1333), .Z(n1332) );
  IV U1311 ( .A(n1328), .Z(n1330) );
  XOR U1312 ( .A(n1334), .B(n1335), .Z(n1328) );
  AND U1313 ( .A(n146), .B(n1327), .Z(n1335) );
  XNOR U1314 ( .A(n1325), .B(n1334), .Z(n1327) );
  XNOR U1315 ( .A(n1336), .B(n1337), .Z(n1325) );
  AND U1316 ( .A(n150), .B(n1338), .Z(n1337) );
  XOR U1317 ( .A(p_input[56]), .B(n1336), .Z(n1338) );
  XNOR U1318 ( .A(n1339), .B(n1340), .Z(n1336) );
  AND U1319 ( .A(n154), .B(n1341), .Z(n1340) );
  XOR U1320 ( .A(n1342), .B(n1343), .Z(n1334) );
  AND U1321 ( .A(n158), .B(n1333), .Z(n1343) );
  XNOR U1322 ( .A(n1344), .B(n1331), .Z(n1333) );
  XOR U1323 ( .A(n1345), .B(n1346), .Z(n1331) );
  AND U1324 ( .A(n181), .B(n1347), .Z(n1346) );
  IV U1325 ( .A(n1342), .Z(n1344) );
  XOR U1326 ( .A(n1348), .B(n1349), .Z(n1342) );
  AND U1327 ( .A(n165), .B(n1341), .Z(n1349) );
  XNOR U1328 ( .A(n1339), .B(n1348), .Z(n1341) );
  XNOR U1329 ( .A(n1350), .B(n1351), .Z(n1339) );
  AND U1330 ( .A(n169), .B(n1352), .Z(n1351) );
  XOR U1331 ( .A(p_input[88]), .B(n1350), .Z(n1352) );
  XNOR U1332 ( .A(n1353), .B(n1354), .Z(n1350) );
  AND U1333 ( .A(n173), .B(n1355), .Z(n1354) );
  XOR U1334 ( .A(n1356), .B(n1357), .Z(n1348) );
  AND U1335 ( .A(n177), .B(n1347), .Z(n1357) );
  XNOR U1336 ( .A(n1358), .B(n1345), .Z(n1347) );
  XOR U1337 ( .A(n1359), .B(n1360), .Z(n1345) );
  AND U1338 ( .A(n200), .B(n1361), .Z(n1360) );
  IV U1339 ( .A(n1356), .Z(n1358) );
  XOR U1340 ( .A(n1362), .B(n1363), .Z(n1356) );
  AND U1341 ( .A(n184), .B(n1355), .Z(n1363) );
  XNOR U1342 ( .A(n1353), .B(n1362), .Z(n1355) );
  XNOR U1343 ( .A(n1364), .B(n1365), .Z(n1353) );
  AND U1344 ( .A(n188), .B(n1366), .Z(n1365) );
  XOR U1345 ( .A(p_input[120]), .B(n1364), .Z(n1366) );
  XNOR U1346 ( .A(n1367), .B(n1368), .Z(n1364) );
  AND U1347 ( .A(n192), .B(n1369), .Z(n1368) );
  XOR U1348 ( .A(n1370), .B(n1371), .Z(n1362) );
  AND U1349 ( .A(n196), .B(n1361), .Z(n1371) );
  XNOR U1350 ( .A(n1372), .B(n1359), .Z(n1361) );
  XOR U1351 ( .A(n1373), .B(n1374), .Z(n1359) );
  AND U1352 ( .A(n218), .B(n1375), .Z(n1374) );
  IV U1353 ( .A(n1370), .Z(n1372) );
  XOR U1354 ( .A(n1376), .B(n1377), .Z(n1370) );
  AND U1355 ( .A(n203), .B(n1369), .Z(n1377) );
  XNOR U1356 ( .A(n1367), .B(n1376), .Z(n1369) );
  XNOR U1357 ( .A(n1378), .B(n1379), .Z(n1367) );
  AND U1358 ( .A(n207), .B(n1380), .Z(n1379) );
  XOR U1359 ( .A(p_input[152]), .B(n1378), .Z(n1380) );
  XOR U1360 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][24] ), .B(n1381), 
        .Z(n1378) );
  AND U1361 ( .A(n210), .B(n1382), .Z(n1381) );
  XOR U1362 ( .A(n1383), .B(n1384), .Z(n1376) );
  AND U1363 ( .A(n214), .B(n1375), .Z(n1384) );
  XNOR U1364 ( .A(n1385), .B(n1373), .Z(n1375) );
  XOR U1365 ( .A(\knn_comb_/min_val_out[0][24] ), .B(n1386), .Z(n1373) );
  AND U1366 ( .A(n226), .B(n1387), .Z(n1386) );
  IV U1367 ( .A(n1383), .Z(n1385) );
  XOR U1368 ( .A(n1388), .B(n1389), .Z(n1383) );
  AND U1369 ( .A(n221), .B(n1382), .Z(n1389) );
  XOR U1370 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][24] ), .B(n1388), 
        .Z(n1382) );
  XOR U1371 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .B(n1390), 
        .Z(n1388) );
  AND U1372 ( .A(n223), .B(n1387), .Z(n1390) );
  XOR U1373 ( .A(\knn_comb_/min_val_out[0][24] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .Z(n1387) );
  XOR U1374 ( .A(n91), .B(n1391), .Z(o[23]) );
  AND U1375 ( .A(n122), .B(n1392), .Z(n91) );
  XOR U1376 ( .A(n92), .B(n1391), .Z(n1392) );
  XOR U1377 ( .A(n1393), .B(n1394), .Z(n1391) );
  AND U1378 ( .A(n142), .B(n1395), .Z(n1394) );
  XOR U1379 ( .A(n1396), .B(n21), .Z(n92) );
  AND U1380 ( .A(n125), .B(n1397), .Z(n21) );
  XOR U1381 ( .A(n22), .B(n1396), .Z(n1397) );
  XOR U1382 ( .A(n1398), .B(n1399), .Z(n22) );
  AND U1383 ( .A(n130), .B(n1400), .Z(n1399) );
  XOR U1384 ( .A(p_input[23]), .B(n1398), .Z(n1400) );
  XNOR U1385 ( .A(n1401), .B(n1402), .Z(n1398) );
  AND U1386 ( .A(n134), .B(n1403), .Z(n1402) );
  XOR U1387 ( .A(n1404), .B(n1405), .Z(n1396) );
  AND U1388 ( .A(n138), .B(n1395), .Z(n1405) );
  XNOR U1389 ( .A(n1406), .B(n1393), .Z(n1395) );
  XOR U1390 ( .A(n1407), .B(n1408), .Z(n1393) );
  AND U1391 ( .A(n162), .B(n1409), .Z(n1408) );
  IV U1392 ( .A(n1404), .Z(n1406) );
  XOR U1393 ( .A(n1410), .B(n1411), .Z(n1404) );
  AND U1394 ( .A(n146), .B(n1403), .Z(n1411) );
  XNOR U1395 ( .A(n1401), .B(n1410), .Z(n1403) );
  XNOR U1396 ( .A(n1412), .B(n1413), .Z(n1401) );
  AND U1397 ( .A(n150), .B(n1414), .Z(n1413) );
  XOR U1398 ( .A(p_input[55]), .B(n1412), .Z(n1414) );
  XNOR U1399 ( .A(n1415), .B(n1416), .Z(n1412) );
  AND U1400 ( .A(n154), .B(n1417), .Z(n1416) );
  XOR U1401 ( .A(n1418), .B(n1419), .Z(n1410) );
  AND U1402 ( .A(n158), .B(n1409), .Z(n1419) );
  XNOR U1403 ( .A(n1420), .B(n1407), .Z(n1409) );
  XOR U1404 ( .A(n1421), .B(n1422), .Z(n1407) );
  AND U1405 ( .A(n181), .B(n1423), .Z(n1422) );
  IV U1406 ( .A(n1418), .Z(n1420) );
  XOR U1407 ( .A(n1424), .B(n1425), .Z(n1418) );
  AND U1408 ( .A(n165), .B(n1417), .Z(n1425) );
  XNOR U1409 ( .A(n1415), .B(n1424), .Z(n1417) );
  XNOR U1410 ( .A(n1426), .B(n1427), .Z(n1415) );
  AND U1411 ( .A(n169), .B(n1428), .Z(n1427) );
  XOR U1412 ( .A(p_input[87]), .B(n1426), .Z(n1428) );
  XNOR U1413 ( .A(n1429), .B(n1430), .Z(n1426) );
  AND U1414 ( .A(n173), .B(n1431), .Z(n1430) );
  XOR U1415 ( .A(n1432), .B(n1433), .Z(n1424) );
  AND U1416 ( .A(n177), .B(n1423), .Z(n1433) );
  XNOR U1417 ( .A(n1434), .B(n1421), .Z(n1423) );
  XOR U1418 ( .A(n1435), .B(n1436), .Z(n1421) );
  AND U1419 ( .A(n200), .B(n1437), .Z(n1436) );
  IV U1420 ( .A(n1432), .Z(n1434) );
  XOR U1421 ( .A(n1438), .B(n1439), .Z(n1432) );
  AND U1422 ( .A(n184), .B(n1431), .Z(n1439) );
  XNOR U1423 ( .A(n1429), .B(n1438), .Z(n1431) );
  XNOR U1424 ( .A(n1440), .B(n1441), .Z(n1429) );
  AND U1425 ( .A(n188), .B(n1442), .Z(n1441) );
  XOR U1426 ( .A(p_input[119]), .B(n1440), .Z(n1442) );
  XNOR U1427 ( .A(n1443), .B(n1444), .Z(n1440) );
  AND U1428 ( .A(n192), .B(n1445), .Z(n1444) );
  XOR U1429 ( .A(n1446), .B(n1447), .Z(n1438) );
  AND U1430 ( .A(n196), .B(n1437), .Z(n1447) );
  XNOR U1431 ( .A(n1448), .B(n1435), .Z(n1437) );
  XOR U1432 ( .A(n1449), .B(n1450), .Z(n1435) );
  AND U1433 ( .A(n218), .B(n1451), .Z(n1450) );
  IV U1434 ( .A(n1446), .Z(n1448) );
  XOR U1435 ( .A(n1452), .B(n1453), .Z(n1446) );
  AND U1436 ( .A(n203), .B(n1445), .Z(n1453) );
  XNOR U1437 ( .A(n1443), .B(n1452), .Z(n1445) );
  XNOR U1438 ( .A(n1454), .B(n1455), .Z(n1443) );
  AND U1439 ( .A(n207), .B(n1456), .Z(n1455) );
  XOR U1440 ( .A(p_input[151]), .B(n1454), .Z(n1456) );
  XOR U1441 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][23] ), .B(n1457), 
        .Z(n1454) );
  AND U1442 ( .A(n210), .B(n1458), .Z(n1457) );
  XOR U1443 ( .A(n1459), .B(n1460), .Z(n1452) );
  AND U1444 ( .A(n214), .B(n1451), .Z(n1460) );
  XNOR U1445 ( .A(n1461), .B(n1449), .Z(n1451) );
  XOR U1446 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n1462), .Z(n1449) );
  AND U1447 ( .A(n226), .B(n1463), .Z(n1462) );
  IV U1448 ( .A(n1459), .Z(n1461) );
  XOR U1449 ( .A(n1464), .B(n1465), .Z(n1459) );
  AND U1450 ( .A(n221), .B(n1458), .Z(n1465) );
  XOR U1451 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][23] ), .B(n1464), 
        .Z(n1458) );
  XOR U1452 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .B(n1466), 
        .Z(n1464) );
  AND U1453 ( .A(n223), .B(n1463), .Z(n1466) );
  XOR U1454 ( .A(n1467), .B(n1468), .Z(n1463) );
  IV U1455 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .Z(n1468) );
  IV U1456 ( .A(\knn_comb_/min_val_out[0][23] ), .Z(n1467) );
  XOR U1457 ( .A(n93), .B(n1469), .Z(o[22]) );
  AND U1458 ( .A(n122), .B(n1470), .Z(n93) );
  XOR U1459 ( .A(n94), .B(n1469), .Z(n1470) );
  XOR U1460 ( .A(n1471), .B(n1472), .Z(n1469) );
  AND U1461 ( .A(n142), .B(n1473), .Z(n1472) );
  XOR U1462 ( .A(n1474), .B(n23), .Z(n94) );
  AND U1463 ( .A(n125), .B(n1475), .Z(n23) );
  XOR U1464 ( .A(n24), .B(n1474), .Z(n1475) );
  XOR U1465 ( .A(n1476), .B(n1477), .Z(n24) );
  AND U1466 ( .A(n130), .B(n1478), .Z(n1477) );
  XOR U1467 ( .A(p_input[22]), .B(n1476), .Z(n1478) );
  XNOR U1468 ( .A(n1479), .B(n1480), .Z(n1476) );
  AND U1469 ( .A(n134), .B(n1481), .Z(n1480) );
  XOR U1470 ( .A(n1482), .B(n1483), .Z(n1474) );
  AND U1471 ( .A(n138), .B(n1473), .Z(n1483) );
  XNOR U1472 ( .A(n1484), .B(n1471), .Z(n1473) );
  XOR U1473 ( .A(n1485), .B(n1486), .Z(n1471) );
  AND U1474 ( .A(n162), .B(n1487), .Z(n1486) );
  IV U1475 ( .A(n1482), .Z(n1484) );
  XOR U1476 ( .A(n1488), .B(n1489), .Z(n1482) );
  AND U1477 ( .A(n146), .B(n1481), .Z(n1489) );
  XNOR U1478 ( .A(n1479), .B(n1488), .Z(n1481) );
  XNOR U1479 ( .A(n1490), .B(n1491), .Z(n1479) );
  AND U1480 ( .A(n150), .B(n1492), .Z(n1491) );
  XOR U1481 ( .A(p_input[54]), .B(n1490), .Z(n1492) );
  XNOR U1482 ( .A(n1493), .B(n1494), .Z(n1490) );
  AND U1483 ( .A(n154), .B(n1495), .Z(n1494) );
  XOR U1484 ( .A(n1496), .B(n1497), .Z(n1488) );
  AND U1485 ( .A(n158), .B(n1487), .Z(n1497) );
  XNOR U1486 ( .A(n1498), .B(n1485), .Z(n1487) );
  XOR U1487 ( .A(n1499), .B(n1500), .Z(n1485) );
  AND U1488 ( .A(n181), .B(n1501), .Z(n1500) );
  IV U1489 ( .A(n1496), .Z(n1498) );
  XOR U1490 ( .A(n1502), .B(n1503), .Z(n1496) );
  AND U1491 ( .A(n165), .B(n1495), .Z(n1503) );
  XNOR U1492 ( .A(n1493), .B(n1502), .Z(n1495) );
  XNOR U1493 ( .A(n1504), .B(n1505), .Z(n1493) );
  AND U1494 ( .A(n169), .B(n1506), .Z(n1505) );
  XOR U1495 ( .A(p_input[86]), .B(n1504), .Z(n1506) );
  XNOR U1496 ( .A(n1507), .B(n1508), .Z(n1504) );
  AND U1497 ( .A(n173), .B(n1509), .Z(n1508) );
  XOR U1498 ( .A(n1510), .B(n1511), .Z(n1502) );
  AND U1499 ( .A(n177), .B(n1501), .Z(n1511) );
  XNOR U1500 ( .A(n1512), .B(n1499), .Z(n1501) );
  XOR U1501 ( .A(n1513), .B(n1514), .Z(n1499) );
  AND U1502 ( .A(n200), .B(n1515), .Z(n1514) );
  IV U1503 ( .A(n1510), .Z(n1512) );
  XOR U1504 ( .A(n1516), .B(n1517), .Z(n1510) );
  AND U1505 ( .A(n184), .B(n1509), .Z(n1517) );
  XNOR U1506 ( .A(n1507), .B(n1516), .Z(n1509) );
  XNOR U1507 ( .A(n1518), .B(n1519), .Z(n1507) );
  AND U1508 ( .A(n188), .B(n1520), .Z(n1519) );
  XOR U1509 ( .A(p_input[118]), .B(n1518), .Z(n1520) );
  XNOR U1510 ( .A(n1521), .B(n1522), .Z(n1518) );
  AND U1511 ( .A(n192), .B(n1523), .Z(n1522) );
  XOR U1512 ( .A(n1524), .B(n1525), .Z(n1516) );
  AND U1513 ( .A(n196), .B(n1515), .Z(n1525) );
  XNOR U1514 ( .A(n1526), .B(n1513), .Z(n1515) );
  XOR U1515 ( .A(n1527), .B(n1528), .Z(n1513) );
  AND U1516 ( .A(n218), .B(n1529), .Z(n1528) );
  IV U1517 ( .A(n1524), .Z(n1526) );
  XOR U1518 ( .A(n1530), .B(n1531), .Z(n1524) );
  AND U1519 ( .A(n203), .B(n1523), .Z(n1531) );
  XNOR U1520 ( .A(n1521), .B(n1530), .Z(n1523) );
  XNOR U1521 ( .A(n1532), .B(n1533), .Z(n1521) );
  AND U1522 ( .A(n207), .B(n1534), .Z(n1533) );
  XOR U1523 ( .A(p_input[150]), .B(n1532), .Z(n1534) );
  XOR U1524 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][22] ), .B(n1535), 
        .Z(n1532) );
  AND U1525 ( .A(n210), .B(n1536), .Z(n1535) );
  XOR U1526 ( .A(n1537), .B(n1538), .Z(n1530) );
  AND U1527 ( .A(n214), .B(n1529), .Z(n1538) );
  XNOR U1528 ( .A(n1539), .B(n1527), .Z(n1529) );
  XOR U1529 ( .A(\knn_comb_/min_val_out[0][22] ), .B(n1540), .Z(n1527) );
  AND U1530 ( .A(n226), .B(n1541), .Z(n1540) );
  IV U1531 ( .A(n1537), .Z(n1539) );
  XOR U1532 ( .A(n1542), .B(n1543), .Z(n1537) );
  AND U1533 ( .A(n221), .B(n1536), .Z(n1543) );
  XOR U1534 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][22] ), .B(n1542), 
        .Z(n1536) );
  XOR U1535 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .B(n1544), 
        .Z(n1542) );
  AND U1536 ( .A(n223), .B(n1541), .Z(n1544) );
  XOR U1537 ( .A(\knn_comb_/min_val_out[0][22] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .Z(n1541) );
  XOR U1538 ( .A(n95), .B(n1545), .Z(o[21]) );
  AND U1539 ( .A(n122), .B(n1546), .Z(n95) );
  XOR U1540 ( .A(n96), .B(n1545), .Z(n1546) );
  XOR U1541 ( .A(n1547), .B(n1548), .Z(n1545) );
  AND U1542 ( .A(n142), .B(n1549), .Z(n1548) );
  XOR U1543 ( .A(n1550), .B(n25), .Z(n96) );
  AND U1544 ( .A(n125), .B(n1551), .Z(n25) );
  XOR U1545 ( .A(n26), .B(n1550), .Z(n1551) );
  XOR U1546 ( .A(n1552), .B(n1553), .Z(n26) );
  AND U1547 ( .A(n130), .B(n1554), .Z(n1553) );
  XOR U1548 ( .A(p_input[21]), .B(n1552), .Z(n1554) );
  XNOR U1549 ( .A(n1555), .B(n1556), .Z(n1552) );
  AND U1550 ( .A(n134), .B(n1557), .Z(n1556) );
  XOR U1551 ( .A(n1558), .B(n1559), .Z(n1550) );
  AND U1552 ( .A(n138), .B(n1549), .Z(n1559) );
  XNOR U1553 ( .A(n1560), .B(n1547), .Z(n1549) );
  XOR U1554 ( .A(n1561), .B(n1562), .Z(n1547) );
  AND U1555 ( .A(n162), .B(n1563), .Z(n1562) );
  IV U1556 ( .A(n1558), .Z(n1560) );
  XOR U1557 ( .A(n1564), .B(n1565), .Z(n1558) );
  AND U1558 ( .A(n146), .B(n1557), .Z(n1565) );
  XNOR U1559 ( .A(n1555), .B(n1564), .Z(n1557) );
  XNOR U1560 ( .A(n1566), .B(n1567), .Z(n1555) );
  AND U1561 ( .A(n150), .B(n1568), .Z(n1567) );
  XOR U1562 ( .A(p_input[53]), .B(n1566), .Z(n1568) );
  XNOR U1563 ( .A(n1569), .B(n1570), .Z(n1566) );
  AND U1564 ( .A(n154), .B(n1571), .Z(n1570) );
  XOR U1565 ( .A(n1572), .B(n1573), .Z(n1564) );
  AND U1566 ( .A(n158), .B(n1563), .Z(n1573) );
  XNOR U1567 ( .A(n1574), .B(n1561), .Z(n1563) );
  XOR U1568 ( .A(n1575), .B(n1576), .Z(n1561) );
  AND U1569 ( .A(n181), .B(n1577), .Z(n1576) );
  IV U1570 ( .A(n1572), .Z(n1574) );
  XOR U1571 ( .A(n1578), .B(n1579), .Z(n1572) );
  AND U1572 ( .A(n165), .B(n1571), .Z(n1579) );
  XNOR U1573 ( .A(n1569), .B(n1578), .Z(n1571) );
  XNOR U1574 ( .A(n1580), .B(n1581), .Z(n1569) );
  AND U1575 ( .A(n169), .B(n1582), .Z(n1581) );
  XOR U1576 ( .A(p_input[85]), .B(n1580), .Z(n1582) );
  XNOR U1577 ( .A(n1583), .B(n1584), .Z(n1580) );
  AND U1578 ( .A(n173), .B(n1585), .Z(n1584) );
  XOR U1579 ( .A(n1586), .B(n1587), .Z(n1578) );
  AND U1580 ( .A(n177), .B(n1577), .Z(n1587) );
  XNOR U1581 ( .A(n1588), .B(n1575), .Z(n1577) );
  XOR U1582 ( .A(n1589), .B(n1590), .Z(n1575) );
  AND U1583 ( .A(n200), .B(n1591), .Z(n1590) );
  IV U1584 ( .A(n1586), .Z(n1588) );
  XOR U1585 ( .A(n1592), .B(n1593), .Z(n1586) );
  AND U1586 ( .A(n184), .B(n1585), .Z(n1593) );
  XNOR U1587 ( .A(n1583), .B(n1592), .Z(n1585) );
  XNOR U1588 ( .A(n1594), .B(n1595), .Z(n1583) );
  AND U1589 ( .A(n188), .B(n1596), .Z(n1595) );
  XOR U1590 ( .A(p_input[117]), .B(n1594), .Z(n1596) );
  XNOR U1591 ( .A(n1597), .B(n1598), .Z(n1594) );
  AND U1592 ( .A(n192), .B(n1599), .Z(n1598) );
  XOR U1593 ( .A(n1600), .B(n1601), .Z(n1592) );
  AND U1594 ( .A(n196), .B(n1591), .Z(n1601) );
  XNOR U1595 ( .A(n1602), .B(n1589), .Z(n1591) );
  XOR U1596 ( .A(n1603), .B(n1604), .Z(n1589) );
  AND U1597 ( .A(n218), .B(n1605), .Z(n1604) );
  IV U1598 ( .A(n1600), .Z(n1602) );
  XOR U1599 ( .A(n1606), .B(n1607), .Z(n1600) );
  AND U1600 ( .A(n203), .B(n1599), .Z(n1607) );
  XNOR U1601 ( .A(n1597), .B(n1606), .Z(n1599) );
  XNOR U1602 ( .A(n1608), .B(n1609), .Z(n1597) );
  AND U1603 ( .A(n207), .B(n1610), .Z(n1609) );
  XOR U1604 ( .A(p_input[149]), .B(n1608), .Z(n1610) );
  XOR U1605 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][21] ), .B(n1611), 
        .Z(n1608) );
  AND U1606 ( .A(n210), .B(n1612), .Z(n1611) );
  XOR U1607 ( .A(n1613), .B(n1614), .Z(n1606) );
  AND U1608 ( .A(n214), .B(n1605), .Z(n1614) );
  XNOR U1609 ( .A(n1615), .B(n1603), .Z(n1605) );
  XOR U1610 ( .A(\knn_comb_/min_val_out[0][21] ), .B(n1616), .Z(n1603) );
  AND U1611 ( .A(n226), .B(n1617), .Z(n1616) );
  IV U1612 ( .A(n1613), .Z(n1615) );
  XOR U1613 ( .A(n1618), .B(n1619), .Z(n1613) );
  AND U1614 ( .A(n221), .B(n1612), .Z(n1619) );
  XOR U1615 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][21] ), .B(n1618), 
        .Z(n1612) );
  XOR U1616 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .B(n1620), 
        .Z(n1618) );
  AND U1617 ( .A(n223), .B(n1617), .Z(n1620) );
  XOR U1618 ( .A(\knn_comb_/min_val_out[0][21] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .Z(n1617) );
  XOR U1619 ( .A(n97), .B(n1621), .Z(o[20]) );
  AND U1620 ( .A(n122), .B(n1622), .Z(n97) );
  XOR U1621 ( .A(n98), .B(n1621), .Z(n1622) );
  XOR U1622 ( .A(n1623), .B(n1624), .Z(n1621) );
  AND U1623 ( .A(n142), .B(n1625), .Z(n1624) );
  XOR U1624 ( .A(n1626), .B(n27), .Z(n98) );
  AND U1625 ( .A(n125), .B(n1627), .Z(n27) );
  XOR U1626 ( .A(n28), .B(n1626), .Z(n1627) );
  XOR U1627 ( .A(n1628), .B(n1629), .Z(n28) );
  AND U1628 ( .A(n130), .B(n1630), .Z(n1629) );
  XOR U1629 ( .A(p_input[20]), .B(n1628), .Z(n1630) );
  XNOR U1630 ( .A(n1631), .B(n1632), .Z(n1628) );
  AND U1631 ( .A(n134), .B(n1633), .Z(n1632) );
  XOR U1632 ( .A(n1634), .B(n1635), .Z(n1626) );
  AND U1633 ( .A(n138), .B(n1625), .Z(n1635) );
  XNOR U1634 ( .A(n1636), .B(n1623), .Z(n1625) );
  XOR U1635 ( .A(n1637), .B(n1638), .Z(n1623) );
  AND U1636 ( .A(n162), .B(n1639), .Z(n1638) );
  IV U1637 ( .A(n1634), .Z(n1636) );
  XOR U1638 ( .A(n1640), .B(n1641), .Z(n1634) );
  AND U1639 ( .A(n146), .B(n1633), .Z(n1641) );
  XNOR U1640 ( .A(n1631), .B(n1640), .Z(n1633) );
  XNOR U1641 ( .A(n1642), .B(n1643), .Z(n1631) );
  AND U1642 ( .A(n150), .B(n1644), .Z(n1643) );
  XOR U1643 ( .A(p_input[52]), .B(n1642), .Z(n1644) );
  XNOR U1644 ( .A(n1645), .B(n1646), .Z(n1642) );
  AND U1645 ( .A(n154), .B(n1647), .Z(n1646) );
  XOR U1646 ( .A(n1648), .B(n1649), .Z(n1640) );
  AND U1647 ( .A(n158), .B(n1639), .Z(n1649) );
  XNOR U1648 ( .A(n1650), .B(n1637), .Z(n1639) );
  XOR U1649 ( .A(n1651), .B(n1652), .Z(n1637) );
  AND U1650 ( .A(n181), .B(n1653), .Z(n1652) );
  IV U1651 ( .A(n1648), .Z(n1650) );
  XOR U1652 ( .A(n1654), .B(n1655), .Z(n1648) );
  AND U1653 ( .A(n165), .B(n1647), .Z(n1655) );
  XNOR U1654 ( .A(n1645), .B(n1654), .Z(n1647) );
  XNOR U1655 ( .A(n1656), .B(n1657), .Z(n1645) );
  AND U1656 ( .A(n169), .B(n1658), .Z(n1657) );
  XOR U1657 ( .A(p_input[84]), .B(n1656), .Z(n1658) );
  XNOR U1658 ( .A(n1659), .B(n1660), .Z(n1656) );
  AND U1659 ( .A(n173), .B(n1661), .Z(n1660) );
  XOR U1660 ( .A(n1662), .B(n1663), .Z(n1654) );
  AND U1661 ( .A(n177), .B(n1653), .Z(n1663) );
  XNOR U1662 ( .A(n1664), .B(n1651), .Z(n1653) );
  XOR U1663 ( .A(n1665), .B(n1666), .Z(n1651) );
  AND U1664 ( .A(n200), .B(n1667), .Z(n1666) );
  IV U1665 ( .A(n1662), .Z(n1664) );
  XOR U1666 ( .A(n1668), .B(n1669), .Z(n1662) );
  AND U1667 ( .A(n184), .B(n1661), .Z(n1669) );
  XNOR U1668 ( .A(n1659), .B(n1668), .Z(n1661) );
  XNOR U1669 ( .A(n1670), .B(n1671), .Z(n1659) );
  AND U1670 ( .A(n188), .B(n1672), .Z(n1671) );
  XOR U1671 ( .A(p_input[116]), .B(n1670), .Z(n1672) );
  XNOR U1672 ( .A(n1673), .B(n1674), .Z(n1670) );
  AND U1673 ( .A(n192), .B(n1675), .Z(n1674) );
  XOR U1674 ( .A(n1676), .B(n1677), .Z(n1668) );
  AND U1675 ( .A(n196), .B(n1667), .Z(n1677) );
  XNOR U1676 ( .A(n1678), .B(n1665), .Z(n1667) );
  XOR U1677 ( .A(n1679), .B(n1680), .Z(n1665) );
  AND U1678 ( .A(n218), .B(n1681), .Z(n1680) );
  IV U1679 ( .A(n1676), .Z(n1678) );
  XOR U1680 ( .A(n1682), .B(n1683), .Z(n1676) );
  AND U1681 ( .A(n203), .B(n1675), .Z(n1683) );
  XNOR U1682 ( .A(n1673), .B(n1682), .Z(n1675) );
  XNOR U1683 ( .A(n1684), .B(n1685), .Z(n1673) );
  AND U1684 ( .A(n207), .B(n1686), .Z(n1685) );
  XOR U1685 ( .A(p_input[148]), .B(n1684), .Z(n1686) );
  XOR U1686 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][20] ), .B(n1687), 
        .Z(n1684) );
  AND U1687 ( .A(n210), .B(n1688), .Z(n1687) );
  XOR U1688 ( .A(n1689), .B(n1690), .Z(n1682) );
  AND U1689 ( .A(n214), .B(n1681), .Z(n1690) );
  XNOR U1690 ( .A(n1691), .B(n1679), .Z(n1681) );
  XOR U1691 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n1692), .Z(n1679) );
  AND U1692 ( .A(n226), .B(n1693), .Z(n1692) );
  IV U1693 ( .A(n1689), .Z(n1691) );
  XOR U1694 ( .A(n1694), .B(n1695), .Z(n1689) );
  AND U1695 ( .A(n221), .B(n1688), .Z(n1695) );
  XOR U1696 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][20] ), .B(n1694), 
        .Z(n1688) );
  XOR U1697 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .B(n1696), 
        .Z(n1694) );
  AND U1698 ( .A(n223), .B(n1693), .Z(n1696) );
  XOR U1699 ( .A(n1697), .B(n1698), .Z(n1693) );
  IV U1700 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .Z(n1698) );
  IV U1701 ( .A(\knn_comb_/min_val_out[0][20] ), .Z(n1697) );
  XOR U1702 ( .A(n697), .B(n1699), .Z(o[1]) );
  AND U1703 ( .A(n122), .B(n1700), .Z(n697) );
  XOR U1704 ( .A(n698), .B(n1699), .Z(n1700) );
  XOR U1705 ( .A(n1701), .B(n1702), .Z(n1699) );
  AND U1706 ( .A(n142), .B(n1703), .Z(n1702) );
  XOR U1707 ( .A(n1704), .B(n69), .Z(n698) );
  AND U1708 ( .A(n125), .B(n1705), .Z(n69) );
  XOR U1709 ( .A(n70), .B(n1704), .Z(n1705) );
  XOR U1710 ( .A(n1706), .B(n1707), .Z(n70) );
  AND U1711 ( .A(n130), .B(n1708), .Z(n1707) );
  XOR U1712 ( .A(p_input[1]), .B(n1706), .Z(n1708) );
  XNOR U1713 ( .A(n1709), .B(n1710), .Z(n1706) );
  AND U1714 ( .A(n134), .B(n1711), .Z(n1710) );
  XOR U1715 ( .A(n1712), .B(n1713), .Z(n1704) );
  AND U1716 ( .A(n138), .B(n1703), .Z(n1713) );
  XNOR U1717 ( .A(n1714), .B(n1701), .Z(n1703) );
  XOR U1718 ( .A(n1715), .B(n1716), .Z(n1701) );
  AND U1719 ( .A(n162), .B(n1717), .Z(n1716) );
  IV U1720 ( .A(n1712), .Z(n1714) );
  XOR U1721 ( .A(n1718), .B(n1719), .Z(n1712) );
  AND U1722 ( .A(n146), .B(n1711), .Z(n1719) );
  XNOR U1723 ( .A(n1709), .B(n1718), .Z(n1711) );
  XNOR U1724 ( .A(n1720), .B(n1721), .Z(n1709) );
  AND U1725 ( .A(n150), .B(n1722), .Z(n1721) );
  XOR U1726 ( .A(p_input[33]), .B(n1720), .Z(n1722) );
  XNOR U1727 ( .A(n1723), .B(n1724), .Z(n1720) );
  AND U1728 ( .A(n154), .B(n1725), .Z(n1724) );
  XOR U1729 ( .A(n1726), .B(n1727), .Z(n1718) );
  AND U1730 ( .A(n158), .B(n1717), .Z(n1727) );
  XNOR U1731 ( .A(n1728), .B(n1715), .Z(n1717) );
  XOR U1732 ( .A(n1729), .B(n1730), .Z(n1715) );
  AND U1733 ( .A(n181), .B(n1731), .Z(n1730) );
  IV U1734 ( .A(n1726), .Z(n1728) );
  XOR U1735 ( .A(n1732), .B(n1733), .Z(n1726) );
  AND U1736 ( .A(n165), .B(n1725), .Z(n1733) );
  XNOR U1737 ( .A(n1723), .B(n1732), .Z(n1725) );
  XNOR U1738 ( .A(n1734), .B(n1735), .Z(n1723) );
  AND U1739 ( .A(n169), .B(n1736), .Z(n1735) );
  XOR U1740 ( .A(p_input[65]), .B(n1734), .Z(n1736) );
  XNOR U1741 ( .A(n1737), .B(n1738), .Z(n1734) );
  AND U1742 ( .A(n173), .B(n1739), .Z(n1738) );
  XOR U1743 ( .A(n1740), .B(n1741), .Z(n1732) );
  AND U1744 ( .A(n177), .B(n1731), .Z(n1741) );
  XNOR U1745 ( .A(n1742), .B(n1729), .Z(n1731) );
  XOR U1746 ( .A(n1743), .B(n1744), .Z(n1729) );
  AND U1747 ( .A(n200), .B(n1745), .Z(n1744) );
  IV U1748 ( .A(n1740), .Z(n1742) );
  XOR U1749 ( .A(n1746), .B(n1747), .Z(n1740) );
  AND U1750 ( .A(n184), .B(n1739), .Z(n1747) );
  XNOR U1751 ( .A(n1737), .B(n1746), .Z(n1739) );
  XNOR U1752 ( .A(n1748), .B(n1749), .Z(n1737) );
  AND U1753 ( .A(n188), .B(n1750), .Z(n1749) );
  XOR U1754 ( .A(p_input[97]), .B(n1748), .Z(n1750) );
  XNOR U1755 ( .A(n1751), .B(n1752), .Z(n1748) );
  AND U1756 ( .A(n192), .B(n1753), .Z(n1752) );
  XOR U1757 ( .A(n1754), .B(n1755), .Z(n1746) );
  AND U1758 ( .A(n196), .B(n1745), .Z(n1755) );
  XNOR U1759 ( .A(n1756), .B(n1743), .Z(n1745) );
  XOR U1760 ( .A(n1757), .B(n1758), .Z(n1743) );
  AND U1761 ( .A(n218), .B(n1759), .Z(n1758) );
  IV U1762 ( .A(n1754), .Z(n1756) );
  XOR U1763 ( .A(n1760), .B(n1761), .Z(n1754) );
  AND U1764 ( .A(n203), .B(n1753), .Z(n1761) );
  XNOR U1765 ( .A(n1751), .B(n1760), .Z(n1753) );
  XNOR U1766 ( .A(n1762), .B(n1763), .Z(n1751) );
  AND U1767 ( .A(n207), .B(n1764), .Z(n1763) );
  XOR U1768 ( .A(p_input[129]), .B(n1762), .Z(n1764) );
  XOR U1769 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n1765), 
        .Z(n1762) );
  AND U1770 ( .A(n210), .B(n1766), .Z(n1765) );
  XOR U1771 ( .A(n1767), .B(n1768), .Z(n1760) );
  AND U1772 ( .A(n214), .B(n1759), .Z(n1768) );
  XNOR U1773 ( .A(n1769), .B(n1757), .Z(n1759) );
  XOR U1774 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n1770), .Z(n1757) );
  AND U1775 ( .A(n226), .B(n1771), .Z(n1770) );
  IV U1776 ( .A(n1767), .Z(n1769) );
  XOR U1777 ( .A(n1772), .B(n1773), .Z(n1767) );
  AND U1778 ( .A(n221), .B(n1766), .Z(n1773) );
  XOR U1779 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n1772), 
        .Z(n1766) );
  XOR U1780 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(n1774), 
        .Z(n1772) );
  AND U1781 ( .A(n223), .B(n1771), .Z(n1774) );
  XOR U1782 ( .A(\knn_comb_/min_val_out[0][1] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n1771) );
  XOR U1783 ( .A(n99), .B(n1775), .Z(o[19]) );
  AND U1784 ( .A(n122), .B(n1776), .Z(n99) );
  XOR U1785 ( .A(n100), .B(n1775), .Z(n1776) );
  XOR U1786 ( .A(n1777), .B(n1778), .Z(n1775) );
  AND U1787 ( .A(n142), .B(n1779), .Z(n1778) );
  XOR U1788 ( .A(n1780), .B(n29), .Z(n100) );
  AND U1789 ( .A(n125), .B(n1781), .Z(n29) );
  XOR U1790 ( .A(n30), .B(n1780), .Z(n1781) );
  XOR U1791 ( .A(n1782), .B(n1783), .Z(n30) );
  AND U1792 ( .A(n130), .B(n1784), .Z(n1783) );
  XOR U1793 ( .A(p_input[19]), .B(n1782), .Z(n1784) );
  XNOR U1794 ( .A(n1785), .B(n1786), .Z(n1782) );
  AND U1795 ( .A(n134), .B(n1787), .Z(n1786) );
  XOR U1796 ( .A(n1788), .B(n1789), .Z(n1780) );
  AND U1797 ( .A(n138), .B(n1779), .Z(n1789) );
  XNOR U1798 ( .A(n1790), .B(n1777), .Z(n1779) );
  XOR U1799 ( .A(n1791), .B(n1792), .Z(n1777) );
  AND U1800 ( .A(n162), .B(n1793), .Z(n1792) );
  IV U1801 ( .A(n1788), .Z(n1790) );
  XOR U1802 ( .A(n1794), .B(n1795), .Z(n1788) );
  AND U1803 ( .A(n146), .B(n1787), .Z(n1795) );
  XNOR U1804 ( .A(n1785), .B(n1794), .Z(n1787) );
  XNOR U1805 ( .A(n1796), .B(n1797), .Z(n1785) );
  AND U1806 ( .A(n150), .B(n1798), .Z(n1797) );
  XOR U1807 ( .A(p_input[51]), .B(n1796), .Z(n1798) );
  XNOR U1808 ( .A(n1799), .B(n1800), .Z(n1796) );
  AND U1809 ( .A(n154), .B(n1801), .Z(n1800) );
  XOR U1810 ( .A(n1802), .B(n1803), .Z(n1794) );
  AND U1811 ( .A(n158), .B(n1793), .Z(n1803) );
  XNOR U1812 ( .A(n1804), .B(n1791), .Z(n1793) );
  XOR U1813 ( .A(n1805), .B(n1806), .Z(n1791) );
  AND U1814 ( .A(n181), .B(n1807), .Z(n1806) );
  IV U1815 ( .A(n1802), .Z(n1804) );
  XOR U1816 ( .A(n1808), .B(n1809), .Z(n1802) );
  AND U1817 ( .A(n165), .B(n1801), .Z(n1809) );
  XNOR U1818 ( .A(n1799), .B(n1808), .Z(n1801) );
  XNOR U1819 ( .A(n1810), .B(n1811), .Z(n1799) );
  AND U1820 ( .A(n169), .B(n1812), .Z(n1811) );
  XOR U1821 ( .A(p_input[83]), .B(n1810), .Z(n1812) );
  XNOR U1822 ( .A(n1813), .B(n1814), .Z(n1810) );
  AND U1823 ( .A(n173), .B(n1815), .Z(n1814) );
  XOR U1824 ( .A(n1816), .B(n1817), .Z(n1808) );
  AND U1825 ( .A(n177), .B(n1807), .Z(n1817) );
  XNOR U1826 ( .A(n1818), .B(n1805), .Z(n1807) );
  XOR U1827 ( .A(n1819), .B(n1820), .Z(n1805) );
  AND U1828 ( .A(n200), .B(n1821), .Z(n1820) );
  IV U1829 ( .A(n1816), .Z(n1818) );
  XOR U1830 ( .A(n1822), .B(n1823), .Z(n1816) );
  AND U1831 ( .A(n184), .B(n1815), .Z(n1823) );
  XNOR U1832 ( .A(n1813), .B(n1822), .Z(n1815) );
  XNOR U1833 ( .A(n1824), .B(n1825), .Z(n1813) );
  AND U1834 ( .A(n188), .B(n1826), .Z(n1825) );
  XOR U1835 ( .A(p_input[115]), .B(n1824), .Z(n1826) );
  XNOR U1836 ( .A(n1827), .B(n1828), .Z(n1824) );
  AND U1837 ( .A(n192), .B(n1829), .Z(n1828) );
  XOR U1838 ( .A(n1830), .B(n1831), .Z(n1822) );
  AND U1839 ( .A(n196), .B(n1821), .Z(n1831) );
  XNOR U1840 ( .A(n1832), .B(n1819), .Z(n1821) );
  XOR U1841 ( .A(n1833), .B(n1834), .Z(n1819) );
  AND U1842 ( .A(n218), .B(n1835), .Z(n1834) );
  IV U1843 ( .A(n1830), .Z(n1832) );
  XOR U1844 ( .A(n1836), .B(n1837), .Z(n1830) );
  AND U1845 ( .A(n203), .B(n1829), .Z(n1837) );
  XNOR U1846 ( .A(n1827), .B(n1836), .Z(n1829) );
  XNOR U1847 ( .A(n1838), .B(n1839), .Z(n1827) );
  AND U1848 ( .A(n207), .B(n1840), .Z(n1839) );
  XOR U1849 ( .A(p_input[147]), .B(n1838), .Z(n1840) );
  XOR U1850 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][19] ), .B(n1841), 
        .Z(n1838) );
  AND U1851 ( .A(n210), .B(n1842), .Z(n1841) );
  XOR U1852 ( .A(n1843), .B(n1844), .Z(n1836) );
  AND U1853 ( .A(n214), .B(n1835), .Z(n1844) );
  XNOR U1854 ( .A(n1845), .B(n1833), .Z(n1835) );
  XOR U1855 ( .A(\knn_comb_/min_val_out[0][19] ), .B(n1846), .Z(n1833) );
  AND U1856 ( .A(n226), .B(n1847), .Z(n1846) );
  IV U1857 ( .A(n1843), .Z(n1845) );
  XOR U1858 ( .A(n1848), .B(n1849), .Z(n1843) );
  AND U1859 ( .A(n221), .B(n1842), .Z(n1849) );
  XOR U1860 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][19] ), .B(n1848), 
        .Z(n1842) );
  XOR U1861 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .B(n1850), 
        .Z(n1848) );
  AND U1862 ( .A(n223), .B(n1847), .Z(n1850) );
  XOR U1863 ( .A(\knn_comb_/min_val_out[0][19] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .Z(n1847) );
  XOR U1864 ( .A(n101), .B(n1851), .Z(o[18]) );
  AND U1865 ( .A(n122), .B(n1852), .Z(n101) );
  XOR U1866 ( .A(n102), .B(n1851), .Z(n1852) );
  XOR U1867 ( .A(n1853), .B(n1854), .Z(n1851) );
  AND U1868 ( .A(n142), .B(n1855), .Z(n1854) );
  XOR U1869 ( .A(n1856), .B(n31), .Z(n102) );
  AND U1870 ( .A(n125), .B(n1857), .Z(n31) );
  XOR U1871 ( .A(n32), .B(n1856), .Z(n1857) );
  XOR U1872 ( .A(n1858), .B(n1859), .Z(n32) );
  AND U1873 ( .A(n130), .B(n1860), .Z(n1859) );
  XOR U1874 ( .A(p_input[18]), .B(n1858), .Z(n1860) );
  XNOR U1875 ( .A(n1861), .B(n1862), .Z(n1858) );
  AND U1876 ( .A(n134), .B(n1863), .Z(n1862) );
  XOR U1877 ( .A(n1864), .B(n1865), .Z(n1856) );
  AND U1878 ( .A(n138), .B(n1855), .Z(n1865) );
  XNOR U1879 ( .A(n1866), .B(n1853), .Z(n1855) );
  XOR U1880 ( .A(n1867), .B(n1868), .Z(n1853) );
  AND U1881 ( .A(n162), .B(n1869), .Z(n1868) );
  IV U1882 ( .A(n1864), .Z(n1866) );
  XOR U1883 ( .A(n1870), .B(n1871), .Z(n1864) );
  AND U1884 ( .A(n146), .B(n1863), .Z(n1871) );
  XNOR U1885 ( .A(n1861), .B(n1870), .Z(n1863) );
  XNOR U1886 ( .A(n1872), .B(n1873), .Z(n1861) );
  AND U1887 ( .A(n150), .B(n1874), .Z(n1873) );
  XOR U1888 ( .A(p_input[50]), .B(n1872), .Z(n1874) );
  XNOR U1889 ( .A(n1875), .B(n1876), .Z(n1872) );
  AND U1890 ( .A(n154), .B(n1877), .Z(n1876) );
  XOR U1891 ( .A(n1878), .B(n1879), .Z(n1870) );
  AND U1892 ( .A(n158), .B(n1869), .Z(n1879) );
  XNOR U1893 ( .A(n1880), .B(n1867), .Z(n1869) );
  XOR U1894 ( .A(n1881), .B(n1882), .Z(n1867) );
  AND U1895 ( .A(n181), .B(n1883), .Z(n1882) );
  IV U1896 ( .A(n1878), .Z(n1880) );
  XOR U1897 ( .A(n1884), .B(n1885), .Z(n1878) );
  AND U1898 ( .A(n165), .B(n1877), .Z(n1885) );
  XNOR U1899 ( .A(n1875), .B(n1884), .Z(n1877) );
  XNOR U1900 ( .A(n1886), .B(n1887), .Z(n1875) );
  AND U1901 ( .A(n169), .B(n1888), .Z(n1887) );
  XOR U1902 ( .A(p_input[82]), .B(n1886), .Z(n1888) );
  XNOR U1903 ( .A(n1889), .B(n1890), .Z(n1886) );
  AND U1904 ( .A(n173), .B(n1891), .Z(n1890) );
  XOR U1905 ( .A(n1892), .B(n1893), .Z(n1884) );
  AND U1906 ( .A(n177), .B(n1883), .Z(n1893) );
  XNOR U1907 ( .A(n1894), .B(n1881), .Z(n1883) );
  XOR U1908 ( .A(n1895), .B(n1896), .Z(n1881) );
  AND U1909 ( .A(n200), .B(n1897), .Z(n1896) );
  IV U1910 ( .A(n1892), .Z(n1894) );
  XOR U1911 ( .A(n1898), .B(n1899), .Z(n1892) );
  AND U1912 ( .A(n184), .B(n1891), .Z(n1899) );
  XNOR U1913 ( .A(n1889), .B(n1898), .Z(n1891) );
  XNOR U1914 ( .A(n1900), .B(n1901), .Z(n1889) );
  AND U1915 ( .A(n188), .B(n1902), .Z(n1901) );
  XOR U1916 ( .A(p_input[114]), .B(n1900), .Z(n1902) );
  XNOR U1917 ( .A(n1903), .B(n1904), .Z(n1900) );
  AND U1918 ( .A(n192), .B(n1905), .Z(n1904) );
  XOR U1919 ( .A(n1906), .B(n1907), .Z(n1898) );
  AND U1920 ( .A(n196), .B(n1897), .Z(n1907) );
  XNOR U1921 ( .A(n1908), .B(n1895), .Z(n1897) );
  XOR U1922 ( .A(n1909), .B(n1910), .Z(n1895) );
  AND U1923 ( .A(n218), .B(n1911), .Z(n1910) );
  IV U1924 ( .A(n1906), .Z(n1908) );
  XOR U1925 ( .A(n1912), .B(n1913), .Z(n1906) );
  AND U1926 ( .A(n203), .B(n1905), .Z(n1913) );
  XNOR U1927 ( .A(n1903), .B(n1912), .Z(n1905) );
  XNOR U1928 ( .A(n1914), .B(n1915), .Z(n1903) );
  AND U1929 ( .A(n207), .B(n1916), .Z(n1915) );
  XOR U1930 ( .A(p_input[146]), .B(n1914), .Z(n1916) );
  XOR U1931 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][18] ), .B(n1917), 
        .Z(n1914) );
  AND U1932 ( .A(n210), .B(n1918), .Z(n1917) );
  XOR U1933 ( .A(n1919), .B(n1920), .Z(n1912) );
  AND U1934 ( .A(n214), .B(n1911), .Z(n1920) );
  XNOR U1935 ( .A(n1921), .B(n1909), .Z(n1911) );
  XOR U1936 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n1922), .Z(n1909) );
  AND U1937 ( .A(n226), .B(n1923), .Z(n1922) );
  IV U1938 ( .A(n1919), .Z(n1921) );
  XOR U1939 ( .A(n1924), .B(n1925), .Z(n1919) );
  AND U1940 ( .A(n221), .B(n1918), .Z(n1925) );
  XOR U1941 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][18] ), .B(n1924), 
        .Z(n1918) );
  XOR U1942 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .B(n1926), 
        .Z(n1924) );
  AND U1943 ( .A(n223), .B(n1923), .Z(n1926) );
  XOR U1944 ( .A(\knn_comb_/min_val_out[0][18] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .Z(n1923) );
  XOR U1945 ( .A(n105), .B(n1927), .Z(o[17]) );
  AND U1946 ( .A(n122), .B(n1928), .Z(n105) );
  XOR U1947 ( .A(n106), .B(n1927), .Z(n1928) );
  XOR U1948 ( .A(n1929), .B(n1930), .Z(n1927) );
  AND U1949 ( .A(n142), .B(n1931), .Z(n1930) );
  XOR U1950 ( .A(n1932), .B(n33), .Z(n106) );
  AND U1951 ( .A(n125), .B(n1933), .Z(n33) );
  XOR U1952 ( .A(n34), .B(n1932), .Z(n1933) );
  XOR U1953 ( .A(n1934), .B(n1935), .Z(n34) );
  AND U1954 ( .A(n130), .B(n1936), .Z(n1935) );
  XOR U1955 ( .A(p_input[17]), .B(n1934), .Z(n1936) );
  XNOR U1956 ( .A(n1937), .B(n1938), .Z(n1934) );
  AND U1957 ( .A(n134), .B(n1939), .Z(n1938) );
  XOR U1958 ( .A(n1940), .B(n1941), .Z(n1932) );
  AND U1959 ( .A(n138), .B(n1931), .Z(n1941) );
  XNOR U1960 ( .A(n1942), .B(n1929), .Z(n1931) );
  XOR U1961 ( .A(n1943), .B(n1944), .Z(n1929) );
  AND U1962 ( .A(n162), .B(n1945), .Z(n1944) );
  IV U1963 ( .A(n1940), .Z(n1942) );
  XOR U1964 ( .A(n1946), .B(n1947), .Z(n1940) );
  AND U1965 ( .A(n146), .B(n1939), .Z(n1947) );
  XNOR U1966 ( .A(n1937), .B(n1946), .Z(n1939) );
  XNOR U1967 ( .A(n1948), .B(n1949), .Z(n1937) );
  AND U1968 ( .A(n150), .B(n1950), .Z(n1949) );
  XOR U1969 ( .A(p_input[49]), .B(n1948), .Z(n1950) );
  XNOR U1970 ( .A(n1951), .B(n1952), .Z(n1948) );
  AND U1971 ( .A(n154), .B(n1953), .Z(n1952) );
  XOR U1972 ( .A(n1954), .B(n1955), .Z(n1946) );
  AND U1973 ( .A(n158), .B(n1945), .Z(n1955) );
  XNOR U1974 ( .A(n1956), .B(n1943), .Z(n1945) );
  XOR U1975 ( .A(n1957), .B(n1958), .Z(n1943) );
  AND U1976 ( .A(n181), .B(n1959), .Z(n1958) );
  IV U1977 ( .A(n1954), .Z(n1956) );
  XOR U1978 ( .A(n1960), .B(n1961), .Z(n1954) );
  AND U1979 ( .A(n165), .B(n1953), .Z(n1961) );
  XNOR U1980 ( .A(n1951), .B(n1960), .Z(n1953) );
  XNOR U1981 ( .A(n1962), .B(n1963), .Z(n1951) );
  AND U1982 ( .A(n169), .B(n1964), .Z(n1963) );
  XOR U1983 ( .A(p_input[81]), .B(n1962), .Z(n1964) );
  XNOR U1984 ( .A(n1965), .B(n1966), .Z(n1962) );
  AND U1985 ( .A(n173), .B(n1967), .Z(n1966) );
  XOR U1986 ( .A(n1968), .B(n1969), .Z(n1960) );
  AND U1987 ( .A(n177), .B(n1959), .Z(n1969) );
  XNOR U1988 ( .A(n1970), .B(n1957), .Z(n1959) );
  XOR U1989 ( .A(n1971), .B(n1972), .Z(n1957) );
  AND U1990 ( .A(n200), .B(n1973), .Z(n1972) );
  IV U1991 ( .A(n1968), .Z(n1970) );
  XOR U1992 ( .A(n1974), .B(n1975), .Z(n1968) );
  AND U1993 ( .A(n184), .B(n1967), .Z(n1975) );
  XNOR U1994 ( .A(n1965), .B(n1974), .Z(n1967) );
  XNOR U1995 ( .A(n1976), .B(n1977), .Z(n1965) );
  AND U1996 ( .A(n188), .B(n1978), .Z(n1977) );
  XOR U1997 ( .A(p_input[113]), .B(n1976), .Z(n1978) );
  XNOR U1998 ( .A(n1979), .B(n1980), .Z(n1976) );
  AND U1999 ( .A(n192), .B(n1981), .Z(n1980) );
  XOR U2000 ( .A(n1982), .B(n1983), .Z(n1974) );
  AND U2001 ( .A(n196), .B(n1973), .Z(n1983) );
  XNOR U2002 ( .A(n1984), .B(n1971), .Z(n1973) );
  XOR U2003 ( .A(n1985), .B(n1986), .Z(n1971) );
  AND U2004 ( .A(n218), .B(n1987), .Z(n1986) );
  IV U2005 ( .A(n1982), .Z(n1984) );
  XOR U2006 ( .A(n1988), .B(n1989), .Z(n1982) );
  AND U2007 ( .A(n203), .B(n1981), .Z(n1989) );
  XNOR U2008 ( .A(n1979), .B(n1988), .Z(n1981) );
  XNOR U2009 ( .A(n1990), .B(n1991), .Z(n1979) );
  AND U2010 ( .A(n207), .B(n1992), .Z(n1991) );
  XOR U2011 ( .A(p_input[145]), .B(n1990), .Z(n1992) );
  XOR U2012 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][17] ), .B(n1993), 
        .Z(n1990) );
  AND U2013 ( .A(n210), .B(n1994), .Z(n1993) );
  XOR U2014 ( .A(n1995), .B(n1996), .Z(n1988) );
  AND U2015 ( .A(n214), .B(n1987), .Z(n1996) );
  XNOR U2016 ( .A(n1997), .B(n1985), .Z(n1987) );
  XOR U2017 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n1998), .Z(n1985) );
  AND U2018 ( .A(n226), .B(n1999), .Z(n1998) );
  IV U2019 ( .A(n1995), .Z(n1997) );
  XOR U2020 ( .A(n2000), .B(n2001), .Z(n1995) );
  AND U2021 ( .A(n221), .B(n1994), .Z(n2001) );
  XOR U2022 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][17] ), .B(n2000), 
        .Z(n1994) );
  XOR U2023 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .B(n2002), 
        .Z(n2000) );
  AND U2024 ( .A(n223), .B(n1999), .Z(n2002) );
  XOR U2025 ( .A(\knn_comb_/min_val_out[0][17] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .Z(n1999) );
  XOR U2026 ( .A(n107), .B(n2003), .Z(o[16]) );
  AND U2027 ( .A(n122), .B(n2004), .Z(n107) );
  XOR U2028 ( .A(n108), .B(n2003), .Z(n2004) );
  XOR U2029 ( .A(n2005), .B(n2006), .Z(n2003) );
  AND U2030 ( .A(n142), .B(n2007), .Z(n2006) );
  XOR U2031 ( .A(n2008), .B(n35), .Z(n108) );
  AND U2032 ( .A(n125), .B(n2009), .Z(n35) );
  XOR U2033 ( .A(n36), .B(n2008), .Z(n2009) );
  XOR U2034 ( .A(n2010), .B(n2011), .Z(n36) );
  AND U2035 ( .A(n130), .B(n2012), .Z(n2011) );
  XOR U2036 ( .A(p_input[16]), .B(n2010), .Z(n2012) );
  XNOR U2037 ( .A(n2013), .B(n2014), .Z(n2010) );
  AND U2038 ( .A(n134), .B(n2015), .Z(n2014) );
  XOR U2039 ( .A(n2016), .B(n2017), .Z(n2008) );
  AND U2040 ( .A(n138), .B(n2007), .Z(n2017) );
  XNOR U2041 ( .A(n2018), .B(n2005), .Z(n2007) );
  XOR U2042 ( .A(n2019), .B(n2020), .Z(n2005) );
  AND U2043 ( .A(n162), .B(n2021), .Z(n2020) );
  IV U2044 ( .A(n2016), .Z(n2018) );
  XOR U2045 ( .A(n2022), .B(n2023), .Z(n2016) );
  AND U2046 ( .A(n146), .B(n2015), .Z(n2023) );
  XNOR U2047 ( .A(n2013), .B(n2022), .Z(n2015) );
  XNOR U2048 ( .A(n2024), .B(n2025), .Z(n2013) );
  AND U2049 ( .A(n150), .B(n2026), .Z(n2025) );
  XOR U2050 ( .A(p_input[48]), .B(n2024), .Z(n2026) );
  XNOR U2051 ( .A(n2027), .B(n2028), .Z(n2024) );
  AND U2052 ( .A(n154), .B(n2029), .Z(n2028) );
  XOR U2053 ( .A(n2030), .B(n2031), .Z(n2022) );
  AND U2054 ( .A(n158), .B(n2021), .Z(n2031) );
  XNOR U2055 ( .A(n2032), .B(n2019), .Z(n2021) );
  XOR U2056 ( .A(n2033), .B(n2034), .Z(n2019) );
  AND U2057 ( .A(n181), .B(n2035), .Z(n2034) );
  IV U2058 ( .A(n2030), .Z(n2032) );
  XOR U2059 ( .A(n2036), .B(n2037), .Z(n2030) );
  AND U2060 ( .A(n165), .B(n2029), .Z(n2037) );
  XNOR U2061 ( .A(n2027), .B(n2036), .Z(n2029) );
  XNOR U2062 ( .A(n2038), .B(n2039), .Z(n2027) );
  AND U2063 ( .A(n169), .B(n2040), .Z(n2039) );
  XOR U2064 ( .A(p_input[80]), .B(n2038), .Z(n2040) );
  XNOR U2065 ( .A(n2041), .B(n2042), .Z(n2038) );
  AND U2066 ( .A(n173), .B(n2043), .Z(n2042) );
  XOR U2067 ( .A(n2044), .B(n2045), .Z(n2036) );
  AND U2068 ( .A(n177), .B(n2035), .Z(n2045) );
  XNOR U2069 ( .A(n2046), .B(n2033), .Z(n2035) );
  XOR U2070 ( .A(n2047), .B(n2048), .Z(n2033) );
  AND U2071 ( .A(n200), .B(n2049), .Z(n2048) );
  IV U2072 ( .A(n2044), .Z(n2046) );
  XOR U2073 ( .A(n2050), .B(n2051), .Z(n2044) );
  AND U2074 ( .A(n184), .B(n2043), .Z(n2051) );
  XNOR U2075 ( .A(n2041), .B(n2050), .Z(n2043) );
  XNOR U2076 ( .A(n2052), .B(n2053), .Z(n2041) );
  AND U2077 ( .A(n188), .B(n2054), .Z(n2053) );
  XOR U2078 ( .A(p_input[112]), .B(n2052), .Z(n2054) );
  XNOR U2079 ( .A(n2055), .B(n2056), .Z(n2052) );
  AND U2080 ( .A(n192), .B(n2057), .Z(n2056) );
  XOR U2081 ( .A(n2058), .B(n2059), .Z(n2050) );
  AND U2082 ( .A(n196), .B(n2049), .Z(n2059) );
  XNOR U2083 ( .A(n2060), .B(n2047), .Z(n2049) );
  XOR U2084 ( .A(n2061), .B(n2062), .Z(n2047) );
  AND U2085 ( .A(n218), .B(n2063), .Z(n2062) );
  IV U2086 ( .A(n2058), .Z(n2060) );
  XOR U2087 ( .A(n2064), .B(n2065), .Z(n2058) );
  AND U2088 ( .A(n203), .B(n2057), .Z(n2065) );
  XNOR U2089 ( .A(n2055), .B(n2064), .Z(n2057) );
  XNOR U2090 ( .A(n2066), .B(n2067), .Z(n2055) );
  AND U2091 ( .A(n207), .B(n2068), .Z(n2067) );
  XOR U2092 ( .A(p_input[144]), .B(n2066), .Z(n2068) );
  XOR U2093 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][16] ), .B(n2069), 
        .Z(n2066) );
  AND U2094 ( .A(n210), .B(n2070), .Z(n2069) );
  XOR U2095 ( .A(n2071), .B(n2072), .Z(n2064) );
  AND U2096 ( .A(n214), .B(n2063), .Z(n2072) );
  XNOR U2097 ( .A(n2073), .B(n2061), .Z(n2063) );
  XOR U2098 ( .A(\knn_comb_/min_val_out[0][16] ), .B(n2074), .Z(n2061) );
  AND U2099 ( .A(n226), .B(n2075), .Z(n2074) );
  IV U2100 ( .A(n2071), .Z(n2073) );
  XOR U2101 ( .A(n2076), .B(n2077), .Z(n2071) );
  AND U2102 ( .A(n221), .B(n2070), .Z(n2077) );
  XOR U2103 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][16] ), .B(n2076), 
        .Z(n2070) );
  XOR U2104 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .B(n2078), 
        .Z(n2076) );
  AND U2105 ( .A(n223), .B(n2075), .Z(n2078) );
  XOR U2106 ( .A(n2079), .B(n2080), .Z(n2075) );
  IV U2107 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .Z(n2080) );
  IV U2108 ( .A(\knn_comb_/min_val_out[0][16] ), .Z(n2079) );
  XOR U2109 ( .A(n109), .B(n2081), .Z(o[15]) );
  AND U2110 ( .A(n122), .B(n2082), .Z(n109) );
  XOR U2111 ( .A(n110), .B(n2081), .Z(n2082) );
  XOR U2112 ( .A(n2083), .B(n2084), .Z(n2081) );
  AND U2113 ( .A(n142), .B(n2085), .Z(n2084) );
  XOR U2114 ( .A(n2086), .B(n39), .Z(n110) );
  AND U2115 ( .A(n125), .B(n2087), .Z(n39) );
  XOR U2116 ( .A(n40), .B(n2086), .Z(n2087) );
  XOR U2117 ( .A(n2088), .B(n2089), .Z(n40) );
  AND U2118 ( .A(n130), .B(n2090), .Z(n2089) );
  XOR U2119 ( .A(p_input[15]), .B(n2088), .Z(n2090) );
  XNOR U2120 ( .A(n2091), .B(n2092), .Z(n2088) );
  AND U2121 ( .A(n134), .B(n2093), .Z(n2092) );
  XOR U2122 ( .A(n2094), .B(n2095), .Z(n2086) );
  AND U2123 ( .A(n138), .B(n2085), .Z(n2095) );
  XNOR U2124 ( .A(n2096), .B(n2083), .Z(n2085) );
  XOR U2125 ( .A(n2097), .B(n2098), .Z(n2083) );
  AND U2126 ( .A(n162), .B(n2099), .Z(n2098) );
  IV U2127 ( .A(n2094), .Z(n2096) );
  XOR U2128 ( .A(n2100), .B(n2101), .Z(n2094) );
  AND U2129 ( .A(n146), .B(n2093), .Z(n2101) );
  XNOR U2130 ( .A(n2091), .B(n2100), .Z(n2093) );
  XNOR U2131 ( .A(n2102), .B(n2103), .Z(n2091) );
  AND U2132 ( .A(n150), .B(n2104), .Z(n2103) );
  XOR U2133 ( .A(p_input[47]), .B(n2102), .Z(n2104) );
  XNOR U2134 ( .A(n2105), .B(n2106), .Z(n2102) );
  AND U2135 ( .A(n154), .B(n2107), .Z(n2106) );
  XOR U2136 ( .A(n2108), .B(n2109), .Z(n2100) );
  AND U2137 ( .A(n158), .B(n2099), .Z(n2109) );
  XNOR U2138 ( .A(n2110), .B(n2097), .Z(n2099) );
  XOR U2139 ( .A(n2111), .B(n2112), .Z(n2097) );
  AND U2140 ( .A(n181), .B(n2113), .Z(n2112) );
  IV U2141 ( .A(n2108), .Z(n2110) );
  XOR U2142 ( .A(n2114), .B(n2115), .Z(n2108) );
  AND U2143 ( .A(n165), .B(n2107), .Z(n2115) );
  XNOR U2144 ( .A(n2105), .B(n2114), .Z(n2107) );
  XNOR U2145 ( .A(n2116), .B(n2117), .Z(n2105) );
  AND U2146 ( .A(n169), .B(n2118), .Z(n2117) );
  XOR U2147 ( .A(p_input[79]), .B(n2116), .Z(n2118) );
  XNOR U2148 ( .A(n2119), .B(n2120), .Z(n2116) );
  AND U2149 ( .A(n173), .B(n2121), .Z(n2120) );
  XOR U2150 ( .A(n2122), .B(n2123), .Z(n2114) );
  AND U2151 ( .A(n177), .B(n2113), .Z(n2123) );
  XNOR U2152 ( .A(n2124), .B(n2111), .Z(n2113) );
  XOR U2153 ( .A(n2125), .B(n2126), .Z(n2111) );
  AND U2154 ( .A(n200), .B(n2127), .Z(n2126) );
  IV U2155 ( .A(n2122), .Z(n2124) );
  XOR U2156 ( .A(n2128), .B(n2129), .Z(n2122) );
  AND U2157 ( .A(n184), .B(n2121), .Z(n2129) );
  XNOR U2158 ( .A(n2119), .B(n2128), .Z(n2121) );
  XNOR U2159 ( .A(n2130), .B(n2131), .Z(n2119) );
  AND U2160 ( .A(n188), .B(n2132), .Z(n2131) );
  XOR U2161 ( .A(p_input[111]), .B(n2130), .Z(n2132) );
  XNOR U2162 ( .A(n2133), .B(n2134), .Z(n2130) );
  AND U2163 ( .A(n192), .B(n2135), .Z(n2134) );
  XOR U2164 ( .A(n2136), .B(n2137), .Z(n2128) );
  AND U2165 ( .A(n196), .B(n2127), .Z(n2137) );
  XNOR U2166 ( .A(n2138), .B(n2125), .Z(n2127) );
  XOR U2167 ( .A(n2139), .B(n2140), .Z(n2125) );
  AND U2168 ( .A(n218), .B(n2141), .Z(n2140) );
  IV U2169 ( .A(n2136), .Z(n2138) );
  XOR U2170 ( .A(n2142), .B(n2143), .Z(n2136) );
  AND U2171 ( .A(n203), .B(n2135), .Z(n2143) );
  XNOR U2172 ( .A(n2133), .B(n2142), .Z(n2135) );
  XNOR U2173 ( .A(n2144), .B(n2145), .Z(n2133) );
  AND U2174 ( .A(n207), .B(n2146), .Z(n2145) );
  XOR U2175 ( .A(p_input[143]), .B(n2144), .Z(n2146) );
  XOR U2176 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n2147), 
        .Z(n2144) );
  AND U2177 ( .A(n210), .B(n2148), .Z(n2147) );
  XOR U2178 ( .A(n2149), .B(n2150), .Z(n2142) );
  AND U2179 ( .A(n214), .B(n2141), .Z(n2150) );
  XNOR U2180 ( .A(n2151), .B(n2139), .Z(n2141) );
  XOR U2181 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n2152), .Z(n2139) );
  AND U2182 ( .A(n226), .B(n2153), .Z(n2152) );
  IV U2183 ( .A(n2149), .Z(n2151) );
  XOR U2184 ( .A(n2154), .B(n2155), .Z(n2149) );
  AND U2185 ( .A(n221), .B(n2148), .Z(n2155) );
  XOR U2186 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n2154), 
        .Z(n2148) );
  XOR U2187 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(n2156), 
        .Z(n2154) );
  AND U2188 ( .A(n223), .B(n2153), .Z(n2156) );
  XOR U2189 ( .A(n2157), .B(n2158), .Z(n2153) );
  IV U2190 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .Z(n2158) );
  IV U2191 ( .A(\knn_comb_/min_val_out[0][15] ), .Z(n2157) );
  XOR U2192 ( .A(n111), .B(n2159), .Z(o[14]) );
  AND U2193 ( .A(n122), .B(n2160), .Z(n111) );
  XOR U2194 ( .A(n112), .B(n2159), .Z(n2160) );
  XOR U2195 ( .A(n2161), .B(n2162), .Z(n2159) );
  AND U2196 ( .A(n142), .B(n2163), .Z(n2162) );
  XOR U2197 ( .A(n2164), .B(n41), .Z(n112) );
  AND U2198 ( .A(n125), .B(n2165), .Z(n41) );
  XOR U2199 ( .A(n42), .B(n2164), .Z(n2165) );
  XOR U2200 ( .A(n2166), .B(n2167), .Z(n42) );
  AND U2201 ( .A(n130), .B(n2168), .Z(n2167) );
  XOR U2202 ( .A(p_input[14]), .B(n2166), .Z(n2168) );
  XNOR U2203 ( .A(n2169), .B(n2170), .Z(n2166) );
  AND U2204 ( .A(n134), .B(n2171), .Z(n2170) );
  XOR U2205 ( .A(n2172), .B(n2173), .Z(n2164) );
  AND U2206 ( .A(n138), .B(n2163), .Z(n2173) );
  XNOR U2207 ( .A(n2174), .B(n2161), .Z(n2163) );
  XOR U2208 ( .A(n2175), .B(n2176), .Z(n2161) );
  AND U2209 ( .A(n162), .B(n2177), .Z(n2176) );
  IV U2210 ( .A(n2172), .Z(n2174) );
  XOR U2211 ( .A(n2178), .B(n2179), .Z(n2172) );
  AND U2212 ( .A(n146), .B(n2171), .Z(n2179) );
  XNOR U2213 ( .A(n2169), .B(n2178), .Z(n2171) );
  XNOR U2214 ( .A(n2180), .B(n2181), .Z(n2169) );
  AND U2215 ( .A(n150), .B(n2182), .Z(n2181) );
  XOR U2216 ( .A(p_input[46]), .B(n2180), .Z(n2182) );
  XNOR U2217 ( .A(n2183), .B(n2184), .Z(n2180) );
  AND U2218 ( .A(n154), .B(n2185), .Z(n2184) );
  XOR U2219 ( .A(n2186), .B(n2187), .Z(n2178) );
  AND U2220 ( .A(n158), .B(n2177), .Z(n2187) );
  XNOR U2221 ( .A(n2188), .B(n2175), .Z(n2177) );
  XOR U2222 ( .A(n2189), .B(n2190), .Z(n2175) );
  AND U2223 ( .A(n181), .B(n2191), .Z(n2190) );
  IV U2224 ( .A(n2186), .Z(n2188) );
  XOR U2225 ( .A(n2192), .B(n2193), .Z(n2186) );
  AND U2226 ( .A(n165), .B(n2185), .Z(n2193) );
  XNOR U2227 ( .A(n2183), .B(n2192), .Z(n2185) );
  XNOR U2228 ( .A(n2194), .B(n2195), .Z(n2183) );
  AND U2229 ( .A(n169), .B(n2196), .Z(n2195) );
  XOR U2230 ( .A(p_input[78]), .B(n2194), .Z(n2196) );
  XNOR U2231 ( .A(n2197), .B(n2198), .Z(n2194) );
  AND U2232 ( .A(n173), .B(n2199), .Z(n2198) );
  XOR U2233 ( .A(n2200), .B(n2201), .Z(n2192) );
  AND U2234 ( .A(n177), .B(n2191), .Z(n2201) );
  XNOR U2235 ( .A(n2202), .B(n2189), .Z(n2191) );
  XOR U2236 ( .A(n2203), .B(n2204), .Z(n2189) );
  AND U2237 ( .A(n200), .B(n2205), .Z(n2204) );
  IV U2238 ( .A(n2200), .Z(n2202) );
  XOR U2239 ( .A(n2206), .B(n2207), .Z(n2200) );
  AND U2240 ( .A(n184), .B(n2199), .Z(n2207) );
  XNOR U2241 ( .A(n2197), .B(n2206), .Z(n2199) );
  XNOR U2242 ( .A(n2208), .B(n2209), .Z(n2197) );
  AND U2243 ( .A(n188), .B(n2210), .Z(n2209) );
  XOR U2244 ( .A(p_input[110]), .B(n2208), .Z(n2210) );
  XNOR U2245 ( .A(n2211), .B(n2212), .Z(n2208) );
  AND U2246 ( .A(n192), .B(n2213), .Z(n2212) );
  XOR U2247 ( .A(n2214), .B(n2215), .Z(n2206) );
  AND U2248 ( .A(n196), .B(n2205), .Z(n2215) );
  XNOR U2249 ( .A(n2216), .B(n2203), .Z(n2205) );
  XOR U2250 ( .A(n2217), .B(n2218), .Z(n2203) );
  AND U2251 ( .A(n218), .B(n2219), .Z(n2218) );
  IV U2252 ( .A(n2214), .Z(n2216) );
  XOR U2253 ( .A(n2220), .B(n2221), .Z(n2214) );
  AND U2254 ( .A(n203), .B(n2213), .Z(n2221) );
  XNOR U2255 ( .A(n2211), .B(n2220), .Z(n2213) );
  XNOR U2256 ( .A(n2222), .B(n2223), .Z(n2211) );
  AND U2257 ( .A(n207), .B(n2224), .Z(n2223) );
  XOR U2258 ( .A(p_input[142]), .B(n2222), .Z(n2224) );
  XOR U2259 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n2225), 
        .Z(n2222) );
  AND U2260 ( .A(n210), .B(n2226), .Z(n2225) );
  XOR U2261 ( .A(n2227), .B(n2228), .Z(n2220) );
  AND U2262 ( .A(n214), .B(n2219), .Z(n2228) );
  XNOR U2263 ( .A(n2229), .B(n2217), .Z(n2219) );
  XOR U2264 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n2230), .Z(n2217) );
  AND U2265 ( .A(n226), .B(n2231), .Z(n2230) );
  IV U2266 ( .A(n2227), .Z(n2229) );
  XOR U2267 ( .A(n2232), .B(n2233), .Z(n2227) );
  AND U2268 ( .A(n221), .B(n2226), .Z(n2233) );
  XOR U2269 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n2232), 
        .Z(n2226) );
  XOR U2270 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(n2234), 
        .Z(n2232) );
  AND U2271 ( .A(n223), .B(n2231), .Z(n2234) );
  XOR U2272 ( .A(\knn_comb_/min_val_out[0][14] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n2231) );
  XOR U2273 ( .A(n113), .B(n2235), .Z(o[13]) );
  AND U2274 ( .A(n122), .B(n2236), .Z(n113) );
  XOR U2275 ( .A(n114), .B(n2235), .Z(n2236) );
  XOR U2276 ( .A(n2237), .B(n2238), .Z(n2235) );
  AND U2277 ( .A(n142), .B(n2239), .Z(n2238) );
  XOR U2278 ( .A(n2240), .B(n43), .Z(n114) );
  AND U2279 ( .A(n125), .B(n2241), .Z(n43) );
  XOR U2280 ( .A(n44), .B(n2240), .Z(n2241) );
  XOR U2281 ( .A(n2242), .B(n2243), .Z(n44) );
  AND U2282 ( .A(n130), .B(n2244), .Z(n2243) );
  XOR U2283 ( .A(p_input[13]), .B(n2242), .Z(n2244) );
  XNOR U2284 ( .A(n2245), .B(n2246), .Z(n2242) );
  AND U2285 ( .A(n134), .B(n2247), .Z(n2246) );
  XOR U2286 ( .A(n2248), .B(n2249), .Z(n2240) );
  AND U2287 ( .A(n138), .B(n2239), .Z(n2249) );
  XNOR U2288 ( .A(n2250), .B(n2237), .Z(n2239) );
  XOR U2289 ( .A(n2251), .B(n2252), .Z(n2237) );
  AND U2290 ( .A(n162), .B(n2253), .Z(n2252) );
  IV U2291 ( .A(n2248), .Z(n2250) );
  XOR U2292 ( .A(n2254), .B(n2255), .Z(n2248) );
  AND U2293 ( .A(n146), .B(n2247), .Z(n2255) );
  XNOR U2294 ( .A(n2245), .B(n2254), .Z(n2247) );
  XNOR U2295 ( .A(n2256), .B(n2257), .Z(n2245) );
  AND U2296 ( .A(n150), .B(n2258), .Z(n2257) );
  XOR U2297 ( .A(p_input[45]), .B(n2256), .Z(n2258) );
  XNOR U2298 ( .A(n2259), .B(n2260), .Z(n2256) );
  AND U2299 ( .A(n154), .B(n2261), .Z(n2260) );
  XOR U2300 ( .A(n2262), .B(n2263), .Z(n2254) );
  AND U2301 ( .A(n158), .B(n2253), .Z(n2263) );
  XNOR U2302 ( .A(n2264), .B(n2251), .Z(n2253) );
  XOR U2303 ( .A(n2265), .B(n2266), .Z(n2251) );
  AND U2304 ( .A(n181), .B(n2267), .Z(n2266) );
  IV U2305 ( .A(n2262), .Z(n2264) );
  XOR U2306 ( .A(n2268), .B(n2269), .Z(n2262) );
  AND U2307 ( .A(n165), .B(n2261), .Z(n2269) );
  XNOR U2308 ( .A(n2259), .B(n2268), .Z(n2261) );
  XNOR U2309 ( .A(n2270), .B(n2271), .Z(n2259) );
  AND U2310 ( .A(n169), .B(n2272), .Z(n2271) );
  XOR U2311 ( .A(p_input[77]), .B(n2270), .Z(n2272) );
  XNOR U2312 ( .A(n2273), .B(n2274), .Z(n2270) );
  AND U2313 ( .A(n173), .B(n2275), .Z(n2274) );
  XOR U2314 ( .A(n2276), .B(n2277), .Z(n2268) );
  AND U2315 ( .A(n177), .B(n2267), .Z(n2277) );
  XNOR U2316 ( .A(n2278), .B(n2265), .Z(n2267) );
  XOR U2317 ( .A(n2279), .B(n2280), .Z(n2265) );
  AND U2318 ( .A(n200), .B(n2281), .Z(n2280) );
  IV U2319 ( .A(n2276), .Z(n2278) );
  XOR U2320 ( .A(n2282), .B(n2283), .Z(n2276) );
  AND U2321 ( .A(n184), .B(n2275), .Z(n2283) );
  XNOR U2322 ( .A(n2273), .B(n2282), .Z(n2275) );
  XNOR U2323 ( .A(n2284), .B(n2285), .Z(n2273) );
  AND U2324 ( .A(n188), .B(n2286), .Z(n2285) );
  XOR U2325 ( .A(p_input[109]), .B(n2284), .Z(n2286) );
  XNOR U2326 ( .A(n2287), .B(n2288), .Z(n2284) );
  AND U2327 ( .A(n192), .B(n2289), .Z(n2288) );
  XOR U2328 ( .A(n2290), .B(n2291), .Z(n2282) );
  AND U2329 ( .A(n196), .B(n2281), .Z(n2291) );
  XNOR U2330 ( .A(n2292), .B(n2279), .Z(n2281) );
  XOR U2331 ( .A(n2293), .B(n2294), .Z(n2279) );
  AND U2332 ( .A(n218), .B(n2295), .Z(n2294) );
  IV U2333 ( .A(n2290), .Z(n2292) );
  XOR U2334 ( .A(n2296), .B(n2297), .Z(n2290) );
  AND U2335 ( .A(n203), .B(n2289), .Z(n2297) );
  XNOR U2336 ( .A(n2287), .B(n2296), .Z(n2289) );
  XNOR U2337 ( .A(n2298), .B(n2299), .Z(n2287) );
  AND U2338 ( .A(n207), .B(n2300), .Z(n2299) );
  XOR U2339 ( .A(p_input[141]), .B(n2298), .Z(n2300) );
  XOR U2340 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(n2301), 
        .Z(n2298) );
  AND U2341 ( .A(n210), .B(n2302), .Z(n2301) );
  XOR U2342 ( .A(n2303), .B(n2304), .Z(n2296) );
  AND U2343 ( .A(n214), .B(n2295), .Z(n2304) );
  XNOR U2344 ( .A(n2305), .B(n2293), .Z(n2295) );
  XOR U2345 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n2306), .Z(n2293) );
  AND U2346 ( .A(n226), .B(n2307), .Z(n2306) );
  IV U2347 ( .A(n2303), .Z(n2305) );
  XOR U2348 ( .A(n2308), .B(n2309), .Z(n2303) );
  AND U2349 ( .A(n221), .B(n2302), .Z(n2309) );
  XOR U2350 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(n2308), 
        .Z(n2302) );
  XOR U2351 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(n2310), 
        .Z(n2308) );
  AND U2352 ( .A(n223), .B(n2307), .Z(n2310) );
  XOR U2353 ( .A(\knn_comb_/min_val_out[0][13] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n2307) );
  XOR U2354 ( .A(n115), .B(n2311), .Z(o[12]) );
  AND U2355 ( .A(n122), .B(n2312), .Z(n115) );
  XOR U2356 ( .A(n116), .B(n2311), .Z(n2312) );
  XOR U2357 ( .A(n2313), .B(n2314), .Z(n2311) );
  AND U2358 ( .A(n142), .B(n2315), .Z(n2314) );
  XOR U2359 ( .A(n2316), .B(n45), .Z(n116) );
  AND U2360 ( .A(n125), .B(n2317), .Z(n45) );
  XOR U2361 ( .A(n46), .B(n2316), .Z(n2317) );
  XOR U2362 ( .A(n2318), .B(n2319), .Z(n46) );
  AND U2363 ( .A(n130), .B(n2320), .Z(n2319) );
  XOR U2364 ( .A(p_input[12]), .B(n2318), .Z(n2320) );
  XNOR U2365 ( .A(n2321), .B(n2322), .Z(n2318) );
  AND U2366 ( .A(n134), .B(n2323), .Z(n2322) );
  XOR U2367 ( .A(n2324), .B(n2325), .Z(n2316) );
  AND U2368 ( .A(n138), .B(n2315), .Z(n2325) );
  XNOR U2369 ( .A(n2326), .B(n2313), .Z(n2315) );
  XOR U2370 ( .A(n2327), .B(n2328), .Z(n2313) );
  AND U2371 ( .A(n162), .B(n2329), .Z(n2328) );
  IV U2372 ( .A(n2324), .Z(n2326) );
  XOR U2373 ( .A(n2330), .B(n2331), .Z(n2324) );
  AND U2374 ( .A(n146), .B(n2323), .Z(n2331) );
  XNOR U2375 ( .A(n2321), .B(n2330), .Z(n2323) );
  XNOR U2376 ( .A(n2332), .B(n2333), .Z(n2321) );
  AND U2377 ( .A(n150), .B(n2334), .Z(n2333) );
  XOR U2378 ( .A(p_input[44]), .B(n2332), .Z(n2334) );
  XNOR U2379 ( .A(n2335), .B(n2336), .Z(n2332) );
  AND U2380 ( .A(n154), .B(n2337), .Z(n2336) );
  XOR U2381 ( .A(n2338), .B(n2339), .Z(n2330) );
  AND U2382 ( .A(n158), .B(n2329), .Z(n2339) );
  XNOR U2383 ( .A(n2340), .B(n2327), .Z(n2329) );
  XOR U2384 ( .A(n2341), .B(n2342), .Z(n2327) );
  AND U2385 ( .A(n181), .B(n2343), .Z(n2342) );
  IV U2386 ( .A(n2338), .Z(n2340) );
  XOR U2387 ( .A(n2344), .B(n2345), .Z(n2338) );
  AND U2388 ( .A(n165), .B(n2337), .Z(n2345) );
  XNOR U2389 ( .A(n2335), .B(n2344), .Z(n2337) );
  XNOR U2390 ( .A(n2346), .B(n2347), .Z(n2335) );
  AND U2391 ( .A(n169), .B(n2348), .Z(n2347) );
  XOR U2392 ( .A(p_input[76]), .B(n2346), .Z(n2348) );
  XNOR U2393 ( .A(n2349), .B(n2350), .Z(n2346) );
  AND U2394 ( .A(n173), .B(n2351), .Z(n2350) );
  XOR U2395 ( .A(n2352), .B(n2353), .Z(n2344) );
  AND U2396 ( .A(n177), .B(n2343), .Z(n2353) );
  XNOR U2397 ( .A(n2354), .B(n2341), .Z(n2343) );
  XOR U2398 ( .A(n2355), .B(n2356), .Z(n2341) );
  AND U2399 ( .A(n200), .B(n2357), .Z(n2356) );
  IV U2400 ( .A(n2352), .Z(n2354) );
  XOR U2401 ( .A(n2358), .B(n2359), .Z(n2352) );
  AND U2402 ( .A(n184), .B(n2351), .Z(n2359) );
  XNOR U2403 ( .A(n2349), .B(n2358), .Z(n2351) );
  XNOR U2404 ( .A(n2360), .B(n2361), .Z(n2349) );
  AND U2405 ( .A(n188), .B(n2362), .Z(n2361) );
  XOR U2406 ( .A(p_input[108]), .B(n2360), .Z(n2362) );
  XNOR U2407 ( .A(n2363), .B(n2364), .Z(n2360) );
  AND U2408 ( .A(n192), .B(n2365), .Z(n2364) );
  XOR U2409 ( .A(n2366), .B(n2367), .Z(n2358) );
  AND U2410 ( .A(n196), .B(n2357), .Z(n2367) );
  XNOR U2411 ( .A(n2368), .B(n2355), .Z(n2357) );
  XOR U2412 ( .A(n2369), .B(n2370), .Z(n2355) );
  AND U2413 ( .A(n218), .B(n2371), .Z(n2370) );
  IV U2414 ( .A(n2366), .Z(n2368) );
  XOR U2415 ( .A(n2372), .B(n2373), .Z(n2366) );
  AND U2416 ( .A(n203), .B(n2365), .Z(n2373) );
  XNOR U2417 ( .A(n2363), .B(n2372), .Z(n2365) );
  XNOR U2418 ( .A(n2374), .B(n2375), .Z(n2363) );
  AND U2419 ( .A(n207), .B(n2376), .Z(n2375) );
  XOR U2420 ( .A(p_input[140]), .B(n2374), .Z(n2376) );
  XOR U2421 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n2377), 
        .Z(n2374) );
  AND U2422 ( .A(n210), .B(n2378), .Z(n2377) );
  XOR U2423 ( .A(n2379), .B(n2380), .Z(n2372) );
  AND U2424 ( .A(n214), .B(n2371), .Z(n2380) );
  XNOR U2425 ( .A(n2381), .B(n2369), .Z(n2371) );
  XOR U2426 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n2382), .Z(n2369) );
  AND U2427 ( .A(n226), .B(n2383), .Z(n2382) );
  IV U2428 ( .A(n2379), .Z(n2381) );
  XOR U2429 ( .A(n2384), .B(n2385), .Z(n2379) );
  AND U2430 ( .A(n221), .B(n2378), .Z(n2385) );
  XOR U2431 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n2384), 
        .Z(n2378) );
  XOR U2432 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(n2386), 
        .Z(n2384) );
  AND U2433 ( .A(n223), .B(n2383), .Z(n2386) );
  XOR U2434 ( .A(n2387), .B(n2388), .Z(n2383) );
  IV U2435 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n2388) );
  IV U2436 ( .A(\knn_comb_/min_val_out[0][12] ), .Z(n2387) );
  XOR U2437 ( .A(n117), .B(n2389), .Z(o[11]) );
  AND U2438 ( .A(n122), .B(n2390), .Z(n117) );
  XOR U2439 ( .A(n118), .B(n2389), .Z(n2390) );
  XOR U2440 ( .A(n2391), .B(n2392), .Z(n2389) );
  AND U2441 ( .A(n142), .B(n2393), .Z(n2392) );
  XOR U2442 ( .A(n2394), .B(n47), .Z(n118) );
  AND U2443 ( .A(n125), .B(n2395), .Z(n47) );
  XOR U2444 ( .A(n48), .B(n2394), .Z(n2395) );
  XOR U2445 ( .A(n2396), .B(n2397), .Z(n48) );
  AND U2446 ( .A(n130), .B(n2398), .Z(n2397) );
  XOR U2447 ( .A(p_input[11]), .B(n2396), .Z(n2398) );
  XNOR U2448 ( .A(n2399), .B(n2400), .Z(n2396) );
  AND U2449 ( .A(n134), .B(n2401), .Z(n2400) );
  XOR U2450 ( .A(n2402), .B(n2403), .Z(n2394) );
  AND U2451 ( .A(n138), .B(n2393), .Z(n2403) );
  XNOR U2452 ( .A(n2404), .B(n2391), .Z(n2393) );
  XOR U2453 ( .A(n2405), .B(n2406), .Z(n2391) );
  AND U2454 ( .A(n162), .B(n2407), .Z(n2406) );
  IV U2455 ( .A(n2402), .Z(n2404) );
  XOR U2456 ( .A(n2408), .B(n2409), .Z(n2402) );
  AND U2457 ( .A(n146), .B(n2401), .Z(n2409) );
  XNOR U2458 ( .A(n2399), .B(n2408), .Z(n2401) );
  XNOR U2459 ( .A(n2410), .B(n2411), .Z(n2399) );
  AND U2460 ( .A(n150), .B(n2412), .Z(n2411) );
  XOR U2461 ( .A(p_input[43]), .B(n2410), .Z(n2412) );
  XNOR U2462 ( .A(n2413), .B(n2414), .Z(n2410) );
  AND U2463 ( .A(n154), .B(n2415), .Z(n2414) );
  XOR U2464 ( .A(n2416), .B(n2417), .Z(n2408) );
  AND U2465 ( .A(n158), .B(n2407), .Z(n2417) );
  XNOR U2466 ( .A(n2418), .B(n2405), .Z(n2407) );
  XOR U2467 ( .A(n2419), .B(n2420), .Z(n2405) );
  AND U2468 ( .A(n181), .B(n2421), .Z(n2420) );
  IV U2469 ( .A(n2416), .Z(n2418) );
  XOR U2470 ( .A(n2422), .B(n2423), .Z(n2416) );
  AND U2471 ( .A(n165), .B(n2415), .Z(n2423) );
  XNOR U2472 ( .A(n2413), .B(n2422), .Z(n2415) );
  XNOR U2473 ( .A(n2424), .B(n2425), .Z(n2413) );
  AND U2474 ( .A(n169), .B(n2426), .Z(n2425) );
  XOR U2475 ( .A(p_input[75]), .B(n2424), .Z(n2426) );
  XNOR U2476 ( .A(n2427), .B(n2428), .Z(n2424) );
  AND U2477 ( .A(n173), .B(n2429), .Z(n2428) );
  XOR U2478 ( .A(n2430), .B(n2431), .Z(n2422) );
  AND U2479 ( .A(n177), .B(n2421), .Z(n2431) );
  XNOR U2480 ( .A(n2432), .B(n2419), .Z(n2421) );
  XOR U2481 ( .A(n2433), .B(n2434), .Z(n2419) );
  AND U2482 ( .A(n200), .B(n2435), .Z(n2434) );
  IV U2483 ( .A(n2430), .Z(n2432) );
  XOR U2484 ( .A(n2436), .B(n2437), .Z(n2430) );
  AND U2485 ( .A(n184), .B(n2429), .Z(n2437) );
  XNOR U2486 ( .A(n2427), .B(n2436), .Z(n2429) );
  XNOR U2487 ( .A(n2438), .B(n2439), .Z(n2427) );
  AND U2488 ( .A(n188), .B(n2440), .Z(n2439) );
  XOR U2489 ( .A(p_input[107]), .B(n2438), .Z(n2440) );
  XNOR U2490 ( .A(n2441), .B(n2442), .Z(n2438) );
  AND U2491 ( .A(n192), .B(n2443), .Z(n2442) );
  XOR U2492 ( .A(n2444), .B(n2445), .Z(n2436) );
  AND U2493 ( .A(n196), .B(n2435), .Z(n2445) );
  XNOR U2494 ( .A(n2446), .B(n2433), .Z(n2435) );
  XOR U2495 ( .A(n2447), .B(n2448), .Z(n2433) );
  AND U2496 ( .A(n218), .B(n2449), .Z(n2448) );
  IV U2497 ( .A(n2444), .Z(n2446) );
  XOR U2498 ( .A(n2450), .B(n2451), .Z(n2444) );
  AND U2499 ( .A(n203), .B(n2443), .Z(n2451) );
  XNOR U2500 ( .A(n2441), .B(n2450), .Z(n2443) );
  XNOR U2501 ( .A(n2452), .B(n2453), .Z(n2441) );
  AND U2502 ( .A(n207), .B(n2454), .Z(n2453) );
  XOR U2503 ( .A(p_input[139]), .B(n2452), .Z(n2454) );
  XOR U2504 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n2455), 
        .Z(n2452) );
  AND U2505 ( .A(n210), .B(n2456), .Z(n2455) );
  XOR U2506 ( .A(n2457), .B(n2458), .Z(n2450) );
  AND U2507 ( .A(n214), .B(n2449), .Z(n2458) );
  XNOR U2508 ( .A(n2459), .B(n2447), .Z(n2449) );
  XOR U2509 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n2460), .Z(n2447) );
  AND U2510 ( .A(n226), .B(n2461), .Z(n2460) );
  IV U2511 ( .A(n2457), .Z(n2459) );
  XOR U2512 ( .A(n2462), .B(n2463), .Z(n2457) );
  AND U2513 ( .A(n221), .B(n2456), .Z(n2463) );
  XOR U2514 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n2462), 
        .Z(n2456) );
  XOR U2515 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n2464), 
        .Z(n2462) );
  AND U2516 ( .A(n223), .B(n2461), .Z(n2464) );
  XOR U2517 ( .A(\knn_comb_/min_val_out[0][11] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n2461) );
  XOR U2518 ( .A(n119), .B(n2465), .Z(o[10]) );
  AND U2519 ( .A(n122), .B(n2466), .Z(n119) );
  XOR U2520 ( .A(n120), .B(n2465), .Z(n2466) );
  XOR U2521 ( .A(n2467), .B(n2468), .Z(n2465) );
  AND U2522 ( .A(n142), .B(n2469), .Z(n2468) );
  XOR U2523 ( .A(n2470), .B(n49), .Z(n120) );
  AND U2524 ( .A(n125), .B(n2471), .Z(n49) );
  XOR U2525 ( .A(n50), .B(n2470), .Z(n2471) );
  XOR U2526 ( .A(n2472), .B(n2473), .Z(n50) );
  AND U2527 ( .A(n130), .B(n2474), .Z(n2473) );
  XOR U2528 ( .A(p_input[10]), .B(n2472), .Z(n2474) );
  XNOR U2529 ( .A(n2475), .B(n2476), .Z(n2472) );
  AND U2530 ( .A(n134), .B(n2477), .Z(n2476) );
  XOR U2531 ( .A(n2478), .B(n2479), .Z(n2470) );
  AND U2532 ( .A(n138), .B(n2469), .Z(n2479) );
  XNOR U2533 ( .A(n2480), .B(n2467), .Z(n2469) );
  XOR U2534 ( .A(n2481), .B(n2482), .Z(n2467) );
  AND U2535 ( .A(n162), .B(n2483), .Z(n2482) );
  IV U2536 ( .A(n2478), .Z(n2480) );
  XOR U2537 ( .A(n2484), .B(n2485), .Z(n2478) );
  AND U2538 ( .A(n146), .B(n2477), .Z(n2485) );
  XNOR U2539 ( .A(n2475), .B(n2484), .Z(n2477) );
  XNOR U2540 ( .A(n2486), .B(n2487), .Z(n2475) );
  AND U2541 ( .A(n150), .B(n2488), .Z(n2487) );
  XOR U2542 ( .A(p_input[42]), .B(n2486), .Z(n2488) );
  XNOR U2543 ( .A(n2489), .B(n2490), .Z(n2486) );
  AND U2544 ( .A(n154), .B(n2491), .Z(n2490) );
  XOR U2545 ( .A(n2492), .B(n2493), .Z(n2484) );
  AND U2546 ( .A(n158), .B(n2483), .Z(n2493) );
  XNOR U2547 ( .A(n2494), .B(n2481), .Z(n2483) );
  XOR U2548 ( .A(n2495), .B(n2496), .Z(n2481) );
  AND U2549 ( .A(n181), .B(n2497), .Z(n2496) );
  IV U2550 ( .A(n2492), .Z(n2494) );
  XOR U2551 ( .A(n2498), .B(n2499), .Z(n2492) );
  AND U2552 ( .A(n165), .B(n2491), .Z(n2499) );
  XNOR U2553 ( .A(n2489), .B(n2498), .Z(n2491) );
  XNOR U2554 ( .A(n2500), .B(n2501), .Z(n2489) );
  AND U2555 ( .A(n169), .B(n2502), .Z(n2501) );
  XOR U2556 ( .A(p_input[74]), .B(n2500), .Z(n2502) );
  XNOR U2557 ( .A(n2503), .B(n2504), .Z(n2500) );
  AND U2558 ( .A(n173), .B(n2505), .Z(n2504) );
  XOR U2559 ( .A(n2506), .B(n2507), .Z(n2498) );
  AND U2560 ( .A(n177), .B(n2497), .Z(n2507) );
  XNOR U2561 ( .A(n2508), .B(n2495), .Z(n2497) );
  XOR U2562 ( .A(n2509), .B(n2510), .Z(n2495) );
  AND U2563 ( .A(n200), .B(n2511), .Z(n2510) );
  IV U2564 ( .A(n2506), .Z(n2508) );
  XOR U2565 ( .A(n2512), .B(n2513), .Z(n2506) );
  AND U2566 ( .A(n184), .B(n2505), .Z(n2513) );
  XNOR U2567 ( .A(n2503), .B(n2512), .Z(n2505) );
  XNOR U2568 ( .A(n2514), .B(n2515), .Z(n2503) );
  AND U2569 ( .A(n188), .B(n2516), .Z(n2515) );
  XOR U2570 ( .A(p_input[106]), .B(n2514), .Z(n2516) );
  XNOR U2571 ( .A(n2517), .B(n2518), .Z(n2514) );
  AND U2572 ( .A(n192), .B(n2519), .Z(n2518) );
  XOR U2573 ( .A(n2520), .B(n2521), .Z(n2512) );
  AND U2574 ( .A(n196), .B(n2511), .Z(n2521) );
  XNOR U2575 ( .A(n2522), .B(n2509), .Z(n2511) );
  XOR U2576 ( .A(n2523), .B(n2524), .Z(n2509) );
  AND U2577 ( .A(n218), .B(n2525), .Z(n2524) );
  IV U2578 ( .A(n2520), .Z(n2522) );
  XOR U2579 ( .A(n2526), .B(n2527), .Z(n2520) );
  AND U2580 ( .A(n203), .B(n2519), .Z(n2527) );
  XNOR U2581 ( .A(n2517), .B(n2526), .Z(n2519) );
  XNOR U2582 ( .A(n2528), .B(n2529), .Z(n2517) );
  AND U2583 ( .A(n207), .B(n2530), .Z(n2529) );
  XOR U2584 ( .A(p_input[138]), .B(n2528), .Z(n2530) );
  XOR U2585 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n2531), 
        .Z(n2528) );
  AND U2586 ( .A(n210), .B(n2532), .Z(n2531) );
  XOR U2587 ( .A(n2533), .B(n2534), .Z(n2526) );
  AND U2588 ( .A(n214), .B(n2525), .Z(n2534) );
  XNOR U2589 ( .A(n2535), .B(n2523), .Z(n2525) );
  XOR U2590 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n2536), .Z(n2523) );
  AND U2591 ( .A(n226), .B(n2537), .Z(n2536) );
  IV U2592 ( .A(n2533), .Z(n2535) );
  XOR U2593 ( .A(n2538), .B(n2539), .Z(n2533) );
  AND U2594 ( .A(n221), .B(n2532), .Z(n2539) );
  XOR U2595 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n2538), 
        .Z(n2532) );
  XOR U2596 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(n2540), 
        .Z(n2538) );
  AND U2597 ( .A(n223), .B(n2537), .Z(n2540) );
  XOR U2598 ( .A(\knn_comb_/min_val_out[0][10] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n2537) );
  XOR U2599 ( .A(n699), .B(n2541), .Z(o[0]) );
  AND U2600 ( .A(n122), .B(n2542), .Z(n699) );
  XOR U2601 ( .A(n700), .B(n2541), .Z(n2542) );
  XOR U2602 ( .A(n2543), .B(n2544), .Z(n2541) );
  AND U2603 ( .A(n142), .B(n2545), .Z(n2544) );
  XOR U2604 ( .A(n2546), .B(n71), .Z(n700) );
  AND U2605 ( .A(n125), .B(n2547), .Z(n71) );
  XOR U2606 ( .A(n72), .B(n2546), .Z(n2547) );
  XOR U2607 ( .A(n2548), .B(n2549), .Z(n72) );
  AND U2608 ( .A(n130), .B(n2550), .Z(n2549) );
  XOR U2609 ( .A(p_input[0]), .B(n2548), .Z(n2550) );
  XNOR U2610 ( .A(n2551), .B(n2552), .Z(n2548) );
  AND U2611 ( .A(n134), .B(n2553), .Z(n2552) );
  XOR U2612 ( .A(n2554), .B(n2555), .Z(n2546) );
  AND U2613 ( .A(n138), .B(n2545), .Z(n2555) );
  XNOR U2614 ( .A(n2556), .B(n2543), .Z(n2545) );
  XOR U2615 ( .A(n2557), .B(n2558), .Z(n2543) );
  AND U2616 ( .A(n162), .B(n2559), .Z(n2558) );
  IV U2617 ( .A(n2554), .Z(n2556) );
  XOR U2618 ( .A(n2560), .B(n2561), .Z(n2554) );
  AND U2619 ( .A(n146), .B(n2553), .Z(n2561) );
  XNOR U2620 ( .A(n2551), .B(n2560), .Z(n2553) );
  XNOR U2621 ( .A(n2562), .B(n2563), .Z(n2551) );
  AND U2622 ( .A(n150), .B(n2564), .Z(n2563) );
  XOR U2623 ( .A(p_input[32]), .B(n2562), .Z(n2564) );
  XNOR U2624 ( .A(n2565), .B(n2566), .Z(n2562) );
  AND U2625 ( .A(n154), .B(n2567), .Z(n2566) );
  XOR U2626 ( .A(n2568), .B(n2569), .Z(n2560) );
  AND U2627 ( .A(n158), .B(n2559), .Z(n2569) );
  XNOR U2628 ( .A(n2570), .B(n2557), .Z(n2559) );
  XOR U2629 ( .A(n2571), .B(n2572), .Z(n2557) );
  AND U2630 ( .A(n181), .B(n2573), .Z(n2572) );
  IV U2631 ( .A(n2568), .Z(n2570) );
  XOR U2632 ( .A(n2574), .B(n2575), .Z(n2568) );
  AND U2633 ( .A(n165), .B(n2567), .Z(n2575) );
  XNOR U2634 ( .A(n2565), .B(n2574), .Z(n2567) );
  XNOR U2635 ( .A(n2576), .B(n2577), .Z(n2565) );
  AND U2636 ( .A(n169), .B(n2578), .Z(n2577) );
  XOR U2637 ( .A(p_input[64]), .B(n2576), .Z(n2578) );
  XNOR U2638 ( .A(n2579), .B(n2580), .Z(n2576) );
  AND U2639 ( .A(n173), .B(n2581), .Z(n2580) );
  XOR U2640 ( .A(n2582), .B(n2583), .Z(n2574) );
  AND U2641 ( .A(n177), .B(n2573), .Z(n2583) );
  XNOR U2642 ( .A(n2584), .B(n2571), .Z(n2573) );
  XOR U2643 ( .A(n2585), .B(n2586), .Z(n2571) );
  AND U2644 ( .A(n200), .B(n2587), .Z(n2586) );
  IV U2645 ( .A(n2582), .Z(n2584) );
  XOR U2646 ( .A(n2588), .B(n2589), .Z(n2582) );
  AND U2647 ( .A(n184), .B(n2581), .Z(n2589) );
  XNOR U2648 ( .A(n2579), .B(n2588), .Z(n2581) );
  XNOR U2649 ( .A(n2590), .B(n2591), .Z(n2579) );
  AND U2650 ( .A(n188), .B(n2592), .Z(n2591) );
  XOR U2651 ( .A(p_input[96]), .B(n2590), .Z(n2592) );
  XNOR U2652 ( .A(n2593), .B(n2594), .Z(n2590) );
  AND U2653 ( .A(n192), .B(n2595), .Z(n2594) );
  XOR U2654 ( .A(n2596), .B(n2597), .Z(n2588) );
  AND U2655 ( .A(n196), .B(n2587), .Z(n2597) );
  XNOR U2656 ( .A(n2598), .B(n2585), .Z(n2587) );
  XOR U2657 ( .A(n2599), .B(n2600), .Z(n2585) );
  AND U2658 ( .A(n218), .B(n2601), .Z(n2600) );
  IV U2659 ( .A(n2596), .Z(n2598) );
  XOR U2660 ( .A(n2602), .B(n2603), .Z(n2596) );
  AND U2661 ( .A(n203), .B(n2595), .Z(n2603) );
  XNOR U2662 ( .A(n2593), .B(n2602), .Z(n2595) );
  XNOR U2663 ( .A(n2604), .B(n2605), .Z(n2593) );
  AND U2664 ( .A(n207), .B(n2606), .Z(n2605) );
  XOR U2665 ( .A(p_input[128]), .B(n2604), .Z(n2606) );
  XOR U2666 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(n2607), 
        .Z(n2604) );
  AND U2667 ( .A(n210), .B(n2608), .Z(n2607) );
  XOR U2668 ( .A(n2609), .B(n2610), .Z(n2602) );
  AND U2669 ( .A(n214), .B(n2601), .Z(n2610) );
  XNOR U2670 ( .A(n2611), .B(n2599), .Z(n2601) );
  XOR U2671 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n2612), .Z(n2599) );
  AND U2672 ( .A(n226), .B(n2613), .Z(n2612) );
  IV U2673 ( .A(n2609), .Z(n2611) );
  XOR U2674 ( .A(n2614), .B(n2615), .Z(n2609) );
  AND U2675 ( .A(n221), .B(n2608), .Z(n2615) );
  XOR U2676 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(n2614), 
        .Z(n2608) );
  XOR U2677 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(n2616), 
        .Z(n2614) );
  AND U2678 ( .A(n223), .B(n2613), .Z(n2616) );
  XOR U2679 ( .A(\knn_comb_/min_val_out[0][0] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n2613) );
  XNOR U2680 ( .A(n2617), .B(n2618), .Z(n122) );
  AND U2681 ( .A(n2619), .B(n2620), .Z(n2618) );
  XNOR U2682 ( .A(n2617), .B(n2621), .Z(n2620) );
  XOR U2683 ( .A(n2622), .B(n2623), .Z(n2621) );
  AND U2684 ( .A(n125), .B(n2624), .Z(n2623) );
  XNOR U2685 ( .A(n2622), .B(n2625), .Z(n2624) );
  IV U2686 ( .A(n2626), .Z(n2622) );
  XNOR U2687 ( .A(n2617), .B(n2627), .Z(n2619) );
  XOR U2688 ( .A(n2628), .B(n2629), .Z(n2627) );
  AND U2689 ( .A(n142), .B(n2630), .Z(n2629) );
  XOR U2690 ( .A(n2631), .B(n2632), .Z(n2617) );
  AND U2691 ( .A(n2633), .B(n2634), .Z(n2632) );
  XOR U2692 ( .A(n2635), .B(n2631), .Z(n2634) );
  XNOR U2693 ( .A(n2636), .B(n2637), .Z(n2635) );
  AND U2694 ( .A(n125), .B(n2638), .Z(n2637) );
  XNOR U2695 ( .A(n2639), .B(n2636), .Z(n2638) );
  XNOR U2696 ( .A(n2631), .B(n2640), .Z(n2633) );
  XOR U2697 ( .A(n2641), .B(n2642), .Z(n2640) );
  AND U2698 ( .A(n142), .B(n2643), .Z(n2642) );
  XOR U2699 ( .A(n2644), .B(n2645), .Z(n2631) );
  AND U2700 ( .A(n2646), .B(n2647), .Z(n2645) );
  XOR U2701 ( .A(n2648), .B(n2644), .Z(n2647) );
  XNOR U2702 ( .A(n2649), .B(n2650), .Z(n2648) );
  AND U2703 ( .A(n125), .B(n2651), .Z(n2650) );
  XNOR U2704 ( .A(n2652), .B(n2649), .Z(n2651) );
  XNOR U2705 ( .A(n2644), .B(n2653), .Z(n2646) );
  XOR U2706 ( .A(n2654), .B(n2655), .Z(n2653) );
  AND U2707 ( .A(n142), .B(n2656), .Z(n2655) );
  XOR U2708 ( .A(n2657), .B(n2658), .Z(n2644) );
  AND U2709 ( .A(n2659), .B(n2660), .Z(n2658) );
  XOR U2710 ( .A(n2661), .B(n2657), .Z(n2660) );
  XNOR U2711 ( .A(n2662), .B(n2663), .Z(n2661) );
  AND U2712 ( .A(n125), .B(n2664), .Z(n2663) );
  XNOR U2713 ( .A(n2665), .B(n2662), .Z(n2664) );
  XNOR U2714 ( .A(n2657), .B(n2666), .Z(n2659) );
  XOR U2715 ( .A(n2667), .B(n2668), .Z(n2666) );
  AND U2716 ( .A(n142), .B(n2669), .Z(n2668) );
  XOR U2717 ( .A(n2670), .B(n2671), .Z(n2657) );
  AND U2718 ( .A(n2672), .B(n2673), .Z(n2671) );
  XOR U2719 ( .A(n2670), .B(n2674), .Z(n2673) );
  XOR U2720 ( .A(n2675), .B(n2676), .Z(n2674) );
  AND U2721 ( .A(n125), .B(n2677), .Z(n2676) );
  XOR U2722 ( .A(n2678), .B(n2675), .Z(n2677) );
  XNOR U2723 ( .A(n2679), .B(n2670), .Z(n2672) );
  XNOR U2724 ( .A(n2680), .B(n2681), .Z(n2679) );
  AND U2725 ( .A(n142), .B(n2682), .Z(n2681) );
  AND U2726 ( .A(n2683), .B(n2684), .Z(n2670) );
  XNOR U2727 ( .A(n2685), .B(n2686), .Z(n2684) );
  AND U2728 ( .A(n125), .B(n2687), .Z(n2686) );
  XNOR U2729 ( .A(n2688), .B(n2685), .Z(n2687) );
  XNOR U2730 ( .A(n2689), .B(n2690), .Z(n125) );
  AND U2731 ( .A(n2691), .B(n2692), .Z(n2690) );
  XOR U2732 ( .A(n2625), .B(n2689), .Z(n2692) );
  XOR U2733 ( .A(n2693), .B(n2694), .Z(n2625) );
  AND U2734 ( .A(n130), .B(n2695), .Z(n2694) );
  XOR U2735 ( .A(n2696), .B(n2693), .Z(n2695) );
  XNOR U2736 ( .A(n2626), .B(n2689), .Z(n2691) );
  XOR U2737 ( .A(n2697), .B(n2698), .Z(n2626) );
  AND U2738 ( .A(n138), .B(n2630), .Z(n2698) );
  XOR U2739 ( .A(n2628), .B(n2697), .Z(n2630) );
  XOR U2740 ( .A(n2699), .B(n2700), .Z(n2689) );
  AND U2741 ( .A(n2701), .B(n2702), .Z(n2700) );
  XOR U2742 ( .A(n2639), .B(n2699), .Z(n2702) );
  XOR U2743 ( .A(n2703), .B(n2704), .Z(n2639) );
  AND U2744 ( .A(n130), .B(n2705), .Z(n2704) );
  XOR U2745 ( .A(n2706), .B(n2703), .Z(n2705) );
  XOR U2746 ( .A(n2699), .B(n2636), .Z(n2701) );
  XOR U2747 ( .A(n2707), .B(n2708), .Z(n2636) );
  AND U2748 ( .A(n138), .B(n2643), .Z(n2708) );
  XOR U2749 ( .A(n2707), .B(n2709), .Z(n2643) );
  XOR U2750 ( .A(n2710), .B(n2711), .Z(n2699) );
  AND U2751 ( .A(n2712), .B(n2713), .Z(n2711) );
  XOR U2752 ( .A(n2652), .B(n2710), .Z(n2713) );
  XOR U2753 ( .A(n2714), .B(n2715), .Z(n2652) );
  AND U2754 ( .A(n130), .B(n2716), .Z(n2715) );
  XNOR U2755 ( .A(n2717), .B(n2714), .Z(n2716) );
  XOR U2756 ( .A(n2710), .B(n2649), .Z(n2712) );
  XOR U2757 ( .A(n2718), .B(n2719), .Z(n2649) );
  AND U2758 ( .A(n138), .B(n2656), .Z(n2719) );
  XOR U2759 ( .A(n2718), .B(n2720), .Z(n2656) );
  XOR U2760 ( .A(n2721), .B(n2722), .Z(n2710) );
  AND U2761 ( .A(n2723), .B(n2724), .Z(n2722) );
  XOR U2762 ( .A(n2665), .B(n2721), .Z(n2724) );
  XOR U2763 ( .A(n2725), .B(n2726), .Z(n2665) );
  AND U2764 ( .A(n130), .B(n2727), .Z(n2726) );
  XOR U2765 ( .A(n2728), .B(n2725), .Z(n2727) );
  XOR U2766 ( .A(n2721), .B(n2662), .Z(n2723) );
  XOR U2767 ( .A(n2729), .B(n2730), .Z(n2662) );
  AND U2768 ( .A(n138), .B(n2669), .Z(n2730) );
  XOR U2769 ( .A(n2729), .B(n2731), .Z(n2669) );
  XOR U2770 ( .A(n2732), .B(n2733), .Z(n2721) );
  AND U2771 ( .A(n2734), .B(n2735), .Z(n2733) );
  XOR U2772 ( .A(n2732), .B(n2678), .Z(n2735) );
  XOR U2773 ( .A(n2736), .B(n2737), .Z(n2678) );
  AND U2774 ( .A(n130), .B(n2738), .Z(n2737) );
  XNOR U2775 ( .A(n2739), .B(n2736), .Z(n2738) );
  XNOR U2776 ( .A(n2675), .B(n2732), .Z(n2734) );
  XNOR U2777 ( .A(n2740), .B(n2741), .Z(n2675) );
  AND U2778 ( .A(n138), .B(n2682), .Z(n2741) );
  XOR U2779 ( .A(n2740), .B(n2680), .Z(n2682) );
  AND U2780 ( .A(n2685), .B(n2688), .Z(n2732) );
  XOR U2781 ( .A(n2742), .B(n2743), .Z(n2688) );
  AND U2782 ( .A(n130), .B(n2744), .Z(n2743) );
  XNOR U2783 ( .A(n2745), .B(n2746), .Z(n2744) );
  XNOR U2784 ( .A(n2747), .B(n2748), .Z(n130) );
  AND U2785 ( .A(n2749), .B(n2750), .Z(n2748) );
  XOR U2786 ( .A(n2696), .B(n2747), .Z(n2750) );
  AND U2787 ( .A(n2751), .B(n2752), .Z(n2696) );
  XNOR U2788 ( .A(n2693), .B(n2747), .Z(n2749) );
  XNOR U2789 ( .A(n2753), .B(n2754), .Z(n2693) );
  AND U2790 ( .A(n134), .B(n2755), .Z(n2754) );
  XNOR U2791 ( .A(n2756), .B(n2757), .Z(n2755) );
  XOR U2792 ( .A(n2758), .B(n2759), .Z(n2747) );
  AND U2793 ( .A(n2760), .B(n2761), .Z(n2759) );
  XNOR U2794 ( .A(n2758), .B(n2751), .Z(n2761) );
  IV U2795 ( .A(n2706), .Z(n2751) );
  XOR U2796 ( .A(n2762), .B(n2763), .Z(n2706) );
  XOR U2797 ( .A(n2764), .B(n2752), .Z(n2763) );
  AND U2798 ( .A(n2717), .B(n2765), .Z(n2752) );
  AND U2799 ( .A(n2766), .B(n2767), .Z(n2764) );
  XOR U2800 ( .A(n2768), .B(n2762), .Z(n2766) );
  XNOR U2801 ( .A(n2703), .B(n2758), .Z(n2760) );
  XNOR U2802 ( .A(n2769), .B(n2770), .Z(n2703) );
  AND U2803 ( .A(n134), .B(n2771), .Z(n2770) );
  XNOR U2804 ( .A(n2772), .B(n2773), .Z(n2771) );
  XOR U2805 ( .A(n2774), .B(n2775), .Z(n2758) );
  AND U2806 ( .A(n2776), .B(n2777), .Z(n2775) );
  XNOR U2807 ( .A(n2774), .B(n2717), .Z(n2777) );
  XOR U2808 ( .A(n2778), .B(n2767), .Z(n2717) );
  XNOR U2809 ( .A(n2779), .B(n2762), .Z(n2767) );
  XOR U2810 ( .A(n2780), .B(n2781), .Z(n2762) );
  AND U2811 ( .A(n2782), .B(n2783), .Z(n2781) );
  XOR U2812 ( .A(n2784), .B(n2780), .Z(n2782) );
  XNOR U2813 ( .A(n2785), .B(n2786), .Z(n2779) );
  AND U2814 ( .A(n2787), .B(n2788), .Z(n2786) );
  XOR U2815 ( .A(n2785), .B(n2789), .Z(n2787) );
  XNOR U2816 ( .A(n2768), .B(n2765), .Z(n2778) );
  AND U2817 ( .A(n2790), .B(n2791), .Z(n2765) );
  XOR U2818 ( .A(n2792), .B(n2793), .Z(n2768) );
  AND U2819 ( .A(n2794), .B(n2795), .Z(n2793) );
  XOR U2820 ( .A(n2792), .B(n2796), .Z(n2794) );
  XNOR U2821 ( .A(n2714), .B(n2774), .Z(n2776) );
  XNOR U2822 ( .A(n2797), .B(n2798), .Z(n2714) );
  AND U2823 ( .A(n134), .B(n2799), .Z(n2798) );
  XNOR U2824 ( .A(n2800), .B(n2801), .Z(n2799) );
  XOR U2825 ( .A(n2802), .B(n2803), .Z(n2774) );
  AND U2826 ( .A(n2804), .B(n2805), .Z(n2803) );
  XNOR U2827 ( .A(n2802), .B(n2790), .Z(n2805) );
  IV U2828 ( .A(n2728), .Z(n2790) );
  XNOR U2829 ( .A(n2806), .B(n2783), .Z(n2728) );
  XNOR U2830 ( .A(n2807), .B(n2789), .Z(n2783) );
  XOR U2831 ( .A(n2808), .B(n2809), .Z(n2789) );
  AND U2832 ( .A(n2810), .B(n2811), .Z(n2809) );
  XOR U2833 ( .A(n2808), .B(n2812), .Z(n2810) );
  XNOR U2834 ( .A(n2788), .B(n2780), .Z(n2807) );
  XOR U2835 ( .A(n2813), .B(n2814), .Z(n2780) );
  AND U2836 ( .A(n2815), .B(n2816), .Z(n2814) );
  XNOR U2837 ( .A(n2817), .B(n2813), .Z(n2815) );
  XNOR U2838 ( .A(n2818), .B(n2785), .Z(n2788) );
  XOR U2839 ( .A(n2819), .B(n2820), .Z(n2785) );
  AND U2840 ( .A(n2821), .B(n2822), .Z(n2820) );
  XOR U2841 ( .A(n2819), .B(n2823), .Z(n2821) );
  XNOR U2842 ( .A(n2824), .B(n2825), .Z(n2818) );
  AND U2843 ( .A(n2826), .B(n2827), .Z(n2825) );
  XNOR U2844 ( .A(n2824), .B(n2828), .Z(n2826) );
  XNOR U2845 ( .A(n2784), .B(n2791), .Z(n2806) );
  AND U2846 ( .A(n2739), .B(n2829), .Z(n2791) );
  XOR U2847 ( .A(n2796), .B(n2795), .Z(n2784) );
  XNOR U2848 ( .A(n2830), .B(n2792), .Z(n2795) );
  XOR U2849 ( .A(n2831), .B(n2832), .Z(n2792) );
  AND U2850 ( .A(n2833), .B(n2834), .Z(n2832) );
  XOR U2851 ( .A(n2831), .B(n2835), .Z(n2833) );
  XNOR U2852 ( .A(n2836), .B(n2837), .Z(n2830) );
  AND U2853 ( .A(n2838), .B(n2839), .Z(n2837) );
  XOR U2854 ( .A(n2836), .B(n2840), .Z(n2838) );
  XOR U2855 ( .A(n2841), .B(n2842), .Z(n2796) );
  AND U2856 ( .A(n2843), .B(n2844), .Z(n2842) );
  XOR U2857 ( .A(n2841), .B(n2845), .Z(n2843) );
  XNOR U2858 ( .A(n2725), .B(n2802), .Z(n2804) );
  XNOR U2859 ( .A(n2846), .B(n2847), .Z(n2725) );
  AND U2860 ( .A(n134), .B(n2848), .Z(n2847) );
  XNOR U2861 ( .A(n2849), .B(n2850), .Z(n2848) );
  XOR U2862 ( .A(n2851), .B(n2852), .Z(n2802) );
  AND U2863 ( .A(n2853), .B(n2854), .Z(n2852) );
  XNOR U2864 ( .A(n2851), .B(n2739), .Z(n2854) );
  XOR U2865 ( .A(n2855), .B(n2816), .Z(n2739) );
  XNOR U2866 ( .A(n2856), .B(n2823), .Z(n2816) );
  XOR U2867 ( .A(n2812), .B(n2811), .Z(n2823) );
  XNOR U2868 ( .A(n2857), .B(n2808), .Z(n2811) );
  XOR U2869 ( .A(n2858), .B(n2859), .Z(n2808) );
  AND U2870 ( .A(n2860), .B(n2861), .Z(n2859) );
  XNOR U2871 ( .A(n2862), .B(n2863), .Z(n2860) );
  IV U2872 ( .A(n2858), .Z(n2862) );
  XNOR U2873 ( .A(n2864), .B(n2865), .Z(n2857) );
  NOR U2874 ( .A(n2866), .B(n2867), .Z(n2865) );
  XNOR U2875 ( .A(n2864), .B(n2868), .Z(n2866) );
  XOR U2876 ( .A(n2869), .B(n2870), .Z(n2812) );
  NOR U2877 ( .A(n2871), .B(n2872), .Z(n2870) );
  XNOR U2878 ( .A(n2869), .B(n2873), .Z(n2871) );
  XNOR U2879 ( .A(n2822), .B(n2813), .Z(n2856) );
  XOR U2880 ( .A(n2874), .B(n2875), .Z(n2813) );
  AND U2881 ( .A(n2876), .B(n2877), .Z(n2875) );
  XOR U2882 ( .A(n2874), .B(n2878), .Z(n2876) );
  XOR U2883 ( .A(n2879), .B(n2828), .Z(n2822) );
  XOR U2884 ( .A(n2880), .B(n2881), .Z(n2828) );
  NOR U2885 ( .A(n2882), .B(n2883), .Z(n2881) );
  XOR U2886 ( .A(n2880), .B(n2884), .Z(n2882) );
  XNOR U2887 ( .A(n2827), .B(n2819), .Z(n2879) );
  XOR U2888 ( .A(n2885), .B(n2886), .Z(n2819) );
  AND U2889 ( .A(n2887), .B(n2888), .Z(n2886) );
  XOR U2890 ( .A(n2885), .B(n2889), .Z(n2887) );
  XNOR U2891 ( .A(n2890), .B(n2824), .Z(n2827) );
  XOR U2892 ( .A(n2891), .B(n2892), .Z(n2824) );
  AND U2893 ( .A(n2893), .B(n2894), .Z(n2892) );
  XNOR U2894 ( .A(n2895), .B(n2896), .Z(n2893) );
  IV U2895 ( .A(n2891), .Z(n2895) );
  XNOR U2896 ( .A(n2897), .B(n2898), .Z(n2890) );
  NOR U2897 ( .A(n2899), .B(n2900), .Z(n2898) );
  XOR U2898 ( .A(n2897), .B(n2901), .Z(n2899) );
  XOR U2899 ( .A(n2817), .B(n2829), .Z(n2855) );
  NOR U2900 ( .A(n2745), .B(n2902), .Z(n2829) );
  XNOR U2901 ( .A(n2835), .B(n2834), .Z(n2817) );
  XNOR U2902 ( .A(n2903), .B(n2840), .Z(n2834) );
  XNOR U2903 ( .A(n2904), .B(n2905), .Z(n2840) );
  NOR U2904 ( .A(n2906), .B(n2907), .Z(n2905) );
  XOR U2905 ( .A(n2904), .B(n2908), .Z(n2906) );
  XNOR U2906 ( .A(n2839), .B(n2831), .Z(n2903) );
  XOR U2907 ( .A(n2909), .B(n2910), .Z(n2831) );
  AND U2908 ( .A(n2911), .B(n2912), .Z(n2910) );
  XNOR U2909 ( .A(n2909), .B(n2913), .Z(n2911) );
  XNOR U2910 ( .A(n2914), .B(n2836), .Z(n2839) );
  XOR U2911 ( .A(n2915), .B(n2916), .Z(n2836) );
  AND U2912 ( .A(n2917), .B(n2918), .Z(n2916) );
  XNOR U2913 ( .A(n2919), .B(n2920), .Z(n2917) );
  IV U2914 ( .A(n2915), .Z(n2919) );
  XNOR U2915 ( .A(n2921), .B(n2922), .Z(n2914) );
  NOR U2916 ( .A(n2923), .B(n2924), .Z(n2922) );
  XNOR U2917 ( .A(n2921), .B(n2925), .Z(n2923) );
  XOR U2918 ( .A(n2845), .B(n2844), .Z(n2835) );
  XNOR U2919 ( .A(n2926), .B(n2841), .Z(n2844) );
  XOR U2920 ( .A(n2927), .B(n2928), .Z(n2841) );
  AND U2921 ( .A(n2929), .B(n2930), .Z(n2928) );
  XOR U2922 ( .A(n2927), .B(n2931), .Z(n2929) );
  XNOR U2923 ( .A(n2932), .B(n2933), .Z(n2926) );
  NOR U2924 ( .A(n2934), .B(n2935), .Z(n2933) );
  XNOR U2925 ( .A(n2932), .B(n2936), .Z(n2934) );
  XOR U2926 ( .A(n2937), .B(n2938), .Z(n2845) );
  NOR U2927 ( .A(n2939), .B(n2940), .Z(n2938) );
  XNOR U2928 ( .A(n2937), .B(n2941), .Z(n2939) );
  XNOR U2929 ( .A(n2736), .B(n2851), .Z(n2853) );
  XNOR U2930 ( .A(n2942), .B(n2943), .Z(n2736) );
  AND U2931 ( .A(n134), .B(n2944), .Z(n2943) );
  XNOR U2932 ( .A(n2945), .B(n2946), .Z(n2944) );
  AND U2933 ( .A(n2746), .B(n2745), .Z(n2851) );
  XOR U2934 ( .A(n2947), .B(n2902), .Z(n2745) );
  XNOR U2935 ( .A(p_input[0]), .B(p_input[256]), .Z(n2902) );
  XNOR U2936 ( .A(n2878), .B(n2877), .Z(n2947) );
  XNOR U2937 ( .A(n2948), .B(n2889), .Z(n2877) );
  XOR U2938 ( .A(n2863), .B(n2861), .Z(n2889) );
  XNOR U2939 ( .A(n2949), .B(n2868), .Z(n2861) );
  XOR U2940 ( .A(p_input[24]), .B(p_input[280]), .Z(n2868) );
  XOR U2941 ( .A(n2858), .B(n2867), .Z(n2949) );
  XOR U2942 ( .A(n2950), .B(n2864), .Z(n2867) );
  XOR U2943 ( .A(p_input[22]), .B(p_input[278]), .Z(n2864) );
  XOR U2944 ( .A(p_input[23]), .B(n2951), .Z(n2950) );
  XOR U2945 ( .A(p_input[18]), .B(p_input[274]), .Z(n2858) );
  XNOR U2946 ( .A(n2873), .B(n2872), .Z(n2863) );
  XOR U2947 ( .A(n2952), .B(n2869), .Z(n2872) );
  XOR U2948 ( .A(p_input[19]), .B(p_input[275]), .Z(n2869) );
  XOR U2949 ( .A(p_input[20]), .B(n2953), .Z(n2952) );
  XOR U2950 ( .A(p_input[21]), .B(p_input[277]), .Z(n2873) );
  XOR U2951 ( .A(n2888), .B(n2954), .Z(n2948) );
  IV U2952 ( .A(n2874), .Z(n2954) );
  XOR U2953 ( .A(p_input[1]), .B(p_input[257]), .Z(n2874) );
  XNOR U2954 ( .A(n2955), .B(n2896), .Z(n2888) );
  XNOR U2955 ( .A(n2884), .B(n2883), .Z(n2896) );
  XNOR U2956 ( .A(n2956), .B(n2880), .Z(n2883) );
  XNOR U2957 ( .A(p_input[26]), .B(p_input[282]), .Z(n2880) );
  XOR U2958 ( .A(p_input[27]), .B(n2957), .Z(n2956) );
  XOR U2959 ( .A(p_input[284]), .B(p_input[28]), .Z(n2884) );
  XOR U2960 ( .A(n2894), .B(n2958), .Z(n2955) );
  IV U2961 ( .A(n2885), .Z(n2958) );
  XOR U2962 ( .A(p_input[17]), .B(p_input[273]), .Z(n2885) );
  XOR U2963 ( .A(n2959), .B(n2901), .Z(n2894) );
  XNOR U2964 ( .A(p_input[287]), .B(p_input[31]), .Z(n2901) );
  XOR U2965 ( .A(n2891), .B(n2900), .Z(n2959) );
  XOR U2966 ( .A(n2960), .B(n2897), .Z(n2900) );
  XOR U2967 ( .A(p_input[285]), .B(p_input[29]), .Z(n2897) );
  XNOR U2968 ( .A(p_input[286]), .B(p_input[30]), .Z(n2960) );
  XOR U2969 ( .A(p_input[25]), .B(p_input[281]), .Z(n2891) );
  XNOR U2970 ( .A(n2913), .B(n2912), .Z(n2878) );
  XNOR U2971 ( .A(n2961), .B(n2920), .Z(n2912) );
  XNOR U2972 ( .A(n2908), .B(n2907), .Z(n2920) );
  XNOR U2973 ( .A(n2962), .B(n2904), .Z(n2907) );
  XNOR U2974 ( .A(p_input[11]), .B(p_input[267]), .Z(n2904) );
  XOR U2975 ( .A(p_input[12]), .B(n2963), .Z(n2962) );
  XOR U2976 ( .A(p_input[13]), .B(p_input[269]), .Z(n2908) );
  XNOR U2977 ( .A(n2918), .B(n2909), .Z(n2961) );
  XOR U2978 ( .A(p_input[258]), .B(p_input[2]), .Z(n2909) );
  XNOR U2979 ( .A(n2964), .B(n2925), .Z(n2918) );
  XNOR U2980 ( .A(p_input[16]), .B(n2965), .Z(n2925) );
  XOR U2981 ( .A(n2915), .B(n2924), .Z(n2964) );
  XOR U2982 ( .A(n2966), .B(n2921), .Z(n2924) );
  XOR U2983 ( .A(p_input[14]), .B(p_input[270]), .Z(n2921) );
  XOR U2984 ( .A(p_input[15]), .B(n2967), .Z(n2966) );
  XOR U2985 ( .A(p_input[10]), .B(p_input[266]), .Z(n2915) );
  XNOR U2986 ( .A(n2931), .B(n2930), .Z(n2913) );
  XNOR U2987 ( .A(n2968), .B(n2936), .Z(n2930) );
  XOR U2988 ( .A(p_input[265]), .B(p_input[9]), .Z(n2936) );
  XOR U2989 ( .A(n2927), .B(n2935), .Z(n2968) );
  XOR U2990 ( .A(n2969), .B(n2932), .Z(n2935) );
  XOR U2991 ( .A(p_input[263]), .B(p_input[7]), .Z(n2932) );
  XNOR U2992 ( .A(p_input[264]), .B(p_input[8]), .Z(n2969) );
  XOR U2993 ( .A(p_input[259]), .B(p_input[3]), .Z(n2927) );
  XNOR U2994 ( .A(n2941), .B(n2940), .Z(n2931) );
  XOR U2995 ( .A(n2970), .B(n2937), .Z(n2940) );
  XOR U2996 ( .A(p_input[260]), .B(p_input[4]), .Z(n2937) );
  XNOR U2997 ( .A(p_input[261]), .B(p_input[5]), .Z(n2970) );
  XOR U2998 ( .A(p_input[262]), .B(p_input[6]), .Z(n2941) );
  IV U2999 ( .A(n2742), .Z(n2746) );
  XOR U3000 ( .A(n2971), .B(n2972), .Z(n2742) );
  AND U3001 ( .A(n134), .B(n2973), .Z(n2972) );
  XNOR U3002 ( .A(n2974), .B(n2975), .Z(n134) );
  AND U3003 ( .A(n2976), .B(n2977), .Z(n2975) );
  XOR U3004 ( .A(n2757), .B(n2974), .Z(n2977) );
  XNOR U3005 ( .A(n2978), .B(n2974), .Z(n2976) );
  XOR U3006 ( .A(n2979), .B(n2980), .Z(n2974) );
  AND U3007 ( .A(n2981), .B(n2982), .Z(n2980) );
  XOR U3008 ( .A(n2772), .B(n2979), .Z(n2982) );
  XOR U3009 ( .A(n2979), .B(n2773), .Z(n2981) );
  XOR U3010 ( .A(n2983), .B(n2984), .Z(n2979) );
  AND U3011 ( .A(n2985), .B(n2986), .Z(n2984) );
  XOR U3012 ( .A(n2800), .B(n2983), .Z(n2986) );
  XOR U3013 ( .A(n2983), .B(n2801), .Z(n2985) );
  XOR U3014 ( .A(n2987), .B(n2988), .Z(n2983) );
  AND U3015 ( .A(n2989), .B(n2990), .Z(n2988) );
  XOR U3016 ( .A(n2849), .B(n2987), .Z(n2990) );
  XOR U3017 ( .A(n2987), .B(n2850), .Z(n2989) );
  XOR U3018 ( .A(n2991), .B(n2992), .Z(n2987) );
  AND U3019 ( .A(n2993), .B(n2994), .Z(n2992) );
  XOR U3020 ( .A(n2991), .B(n2945), .Z(n2994) );
  XNOR U3021 ( .A(n2995), .B(n2996), .Z(n2685) );
  AND U3022 ( .A(n138), .B(n2997), .Z(n2996) );
  XNOR U3023 ( .A(n2998), .B(n2999), .Z(n138) );
  AND U3024 ( .A(n3000), .B(n3001), .Z(n2999) );
  XOR U3025 ( .A(n2998), .B(n2697), .Z(n3001) );
  XNOR U3026 ( .A(n2998), .B(n2628), .Z(n3000) );
  XOR U3027 ( .A(n3002), .B(n3003), .Z(n2998) );
  AND U3028 ( .A(n3004), .B(n3005), .Z(n3003) );
  XNOR U3029 ( .A(n2707), .B(n3002), .Z(n3005) );
  XOR U3030 ( .A(n3002), .B(n2709), .Z(n3004) );
  XOR U3031 ( .A(n3006), .B(n3007), .Z(n3002) );
  AND U3032 ( .A(n3008), .B(n3009), .Z(n3007) );
  XNOR U3033 ( .A(n2718), .B(n3006), .Z(n3009) );
  XOR U3034 ( .A(n3006), .B(n2720), .Z(n3008) );
  IV U3035 ( .A(n2654), .Z(n2720) );
  XOR U3036 ( .A(n3010), .B(n3011), .Z(n3006) );
  AND U3037 ( .A(n3012), .B(n3013), .Z(n3011) );
  XOR U3038 ( .A(n3010), .B(n2731), .Z(n3012) );
  XOR U3039 ( .A(n3014), .B(n3015), .Z(n2683) );
  AND U3040 ( .A(n142), .B(n2997), .Z(n3015) );
  XNOR U3041 ( .A(n2995), .B(n3014), .Z(n2997) );
  XNOR U3042 ( .A(n3016), .B(n3017), .Z(n142) );
  AND U3043 ( .A(n3018), .B(n3019), .Z(n3017) );
  XNOR U3044 ( .A(n3020), .B(n3016), .Z(n3019) );
  IV U3045 ( .A(n2697), .Z(n3020) );
  XOR U3046 ( .A(n2978), .B(n3021), .Z(n2697) );
  AND U3047 ( .A(n146), .B(n3022), .Z(n3021) );
  XOR U3048 ( .A(n2756), .B(n2753), .Z(n3022) );
  XNOR U3049 ( .A(n2628), .B(n3016), .Z(n3018) );
  XNOR U3050 ( .A(n3023), .B(n3024), .Z(n2628) );
  AND U3051 ( .A(n162), .B(n3025), .Z(n3024) );
  XNOR U3052 ( .A(n3026), .B(n3027), .Z(n3025) );
  XOR U3053 ( .A(n3028), .B(n3029), .Z(n3016) );
  AND U3054 ( .A(n3030), .B(n3031), .Z(n3029) );
  XNOR U3055 ( .A(n3028), .B(n2707), .Z(n3031) );
  XOR U3056 ( .A(n2773), .B(n3032), .Z(n2707) );
  AND U3057 ( .A(n146), .B(n3033), .Z(n3032) );
  XOR U3058 ( .A(n2769), .B(n2773), .Z(n3033) );
  XNOR U3059 ( .A(n2641), .B(n3028), .Z(n3030) );
  IV U3060 ( .A(n2709), .Z(n2641) );
  XOR U3061 ( .A(n3034), .B(n3035), .Z(n2709) );
  AND U3062 ( .A(n162), .B(n3036), .Z(n3035) );
  XOR U3063 ( .A(n3037), .B(n3038), .Z(n3028) );
  AND U3064 ( .A(n3039), .B(n3040), .Z(n3038) );
  XNOR U3065 ( .A(n3037), .B(n2718), .Z(n3040) );
  XOR U3066 ( .A(n2801), .B(n3041), .Z(n2718) );
  AND U3067 ( .A(n146), .B(n3042), .Z(n3041) );
  XOR U3068 ( .A(n2797), .B(n2801), .Z(n3042) );
  XNOR U3069 ( .A(n2654), .B(n3037), .Z(n3039) );
  XNOR U3070 ( .A(n3043), .B(n3044), .Z(n2654) );
  AND U3071 ( .A(n162), .B(n3045), .Z(n3044) );
  XOR U3072 ( .A(n3010), .B(n3046), .Z(n3037) );
  AND U3073 ( .A(n3047), .B(n3013), .Z(n3046) );
  XNOR U3074 ( .A(n2729), .B(n3010), .Z(n3013) );
  XOR U3075 ( .A(n2850), .B(n3048), .Z(n2729) );
  AND U3076 ( .A(n146), .B(n3049), .Z(n3048) );
  XOR U3077 ( .A(n2846), .B(n2850), .Z(n3049) );
  XNOR U3078 ( .A(n2667), .B(n3010), .Z(n3047) );
  IV U3079 ( .A(n2731), .Z(n2667) );
  XOR U3080 ( .A(n3050), .B(n3051), .Z(n2731) );
  AND U3081 ( .A(n162), .B(n3052), .Z(n3051) );
  XOR U3082 ( .A(n3053), .B(n3054), .Z(n3010) );
  AND U3083 ( .A(n3055), .B(n3056), .Z(n3054) );
  XNOR U3084 ( .A(n3053), .B(n2740), .Z(n3056) );
  XOR U3085 ( .A(n2946), .B(n3057), .Z(n2740) );
  AND U3086 ( .A(n146), .B(n3058), .Z(n3057) );
  XOR U3087 ( .A(n2942), .B(n2946), .Z(n3058) );
  XNOR U3088 ( .A(n3059), .B(n3053), .Z(n3055) );
  IV U3089 ( .A(n2680), .Z(n3059) );
  XOR U3090 ( .A(n3060), .B(n3061), .Z(n2680) );
  AND U3091 ( .A(n162), .B(n3062), .Z(n3061) );
  AND U3092 ( .A(n3014), .B(n2995), .Z(n3053) );
  XNOR U3093 ( .A(n3063), .B(n3064), .Z(n2995) );
  AND U3094 ( .A(n146), .B(n2973), .Z(n3064) );
  XNOR U3095 ( .A(n2971), .B(n3063), .Z(n2973) );
  XNOR U3096 ( .A(n3065), .B(n3066), .Z(n146) );
  AND U3097 ( .A(n3067), .B(n3068), .Z(n3066) );
  XNOR U3098 ( .A(n3065), .B(n2753), .Z(n3068) );
  IV U3099 ( .A(n2757), .Z(n2753) );
  XOR U3100 ( .A(n3069), .B(n3070), .Z(n2757) );
  AND U3101 ( .A(n150), .B(n3071), .Z(n3070) );
  XOR U3102 ( .A(n3072), .B(n3069), .Z(n3071) );
  XNOR U3103 ( .A(n3065), .B(n2978), .Z(n3067) );
  IV U3104 ( .A(n2756), .Z(n2978) );
  XOR U3105 ( .A(n3026), .B(n3073), .Z(n2756) );
  AND U3106 ( .A(n158), .B(n3074), .Z(n3073) );
  XOR U3107 ( .A(n3026), .B(n3023), .Z(n3074) );
  XOR U3108 ( .A(n3075), .B(n3076), .Z(n3065) );
  AND U3109 ( .A(n3077), .B(n3078), .Z(n3076) );
  XNOR U3110 ( .A(n3075), .B(n2769), .Z(n3078) );
  IV U3111 ( .A(n2772), .Z(n2769) );
  XOR U3112 ( .A(n3079), .B(n3080), .Z(n2772) );
  AND U3113 ( .A(n150), .B(n3081), .Z(n3080) );
  XOR U3114 ( .A(n3082), .B(n3079), .Z(n3081) );
  XOR U3115 ( .A(n2773), .B(n3075), .Z(n3077) );
  XOR U3116 ( .A(n3083), .B(n3084), .Z(n2773) );
  AND U3117 ( .A(n158), .B(n3036), .Z(n3084) );
  XOR U3118 ( .A(n3083), .B(n3034), .Z(n3036) );
  XOR U3119 ( .A(n3085), .B(n3086), .Z(n3075) );
  AND U3120 ( .A(n3087), .B(n3088), .Z(n3086) );
  XNOR U3121 ( .A(n3085), .B(n2797), .Z(n3088) );
  IV U3122 ( .A(n2800), .Z(n2797) );
  XOR U3123 ( .A(n3089), .B(n3090), .Z(n2800) );
  AND U3124 ( .A(n150), .B(n3091), .Z(n3090) );
  XNOR U3125 ( .A(n3092), .B(n3089), .Z(n3091) );
  XOR U3126 ( .A(n2801), .B(n3085), .Z(n3087) );
  XOR U3127 ( .A(n3093), .B(n3094), .Z(n2801) );
  AND U3128 ( .A(n158), .B(n3045), .Z(n3094) );
  XOR U3129 ( .A(n3093), .B(n3043), .Z(n3045) );
  XOR U3130 ( .A(n3095), .B(n3096), .Z(n3085) );
  AND U3131 ( .A(n3097), .B(n3098), .Z(n3096) );
  XNOR U3132 ( .A(n3095), .B(n2846), .Z(n3098) );
  IV U3133 ( .A(n2849), .Z(n2846) );
  XOR U3134 ( .A(n3099), .B(n3100), .Z(n2849) );
  AND U3135 ( .A(n150), .B(n3101), .Z(n3100) );
  XOR U3136 ( .A(n3102), .B(n3099), .Z(n3101) );
  XOR U3137 ( .A(n2850), .B(n3095), .Z(n3097) );
  XOR U3138 ( .A(n3103), .B(n3104), .Z(n2850) );
  AND U3139 ( .A(n158), .B(n3052), .Z(n3104) );
  XOR U3140 ( .A(n3103), .B(n3050), .Z(n3052) );
  XOR U3141 ( .A(n2991), .B(n3105), .Z(n3095) );
  AND U3142 ( .A(n2993), .B(n3106), .Z(n3105) );
  XNOR U3143 ( .A(n2991), .B(n2942), .Z(n3106) );
  IV U3144 ( .A(n2945), .Z(n2942) );
  XOR U3145 ( .A(n3107), .B(n3108), .Z(n2945) );
  AND U3146 ( .A(n150), .B(n3109), .Z(n3108) );
  XNOR U3147 ( .A(n3110), .B(n3107), .Z(n3109) );
  XOR U3148 ( .A(n2946), .B(n2991), .Z(n2993) );
  XOR U3149 ( .A(n3111), .B(n3112), .Z(n2946) );
  AND U3150 ( .A(n158), .B(n3062), .Z(n3112) );
  XOR U3151 ( .A(n3111), .B(n3060), .Z(n3062) );
  AND U3152 ( .A(n3063), .B(n2971), .Z(n2991) );
  XNOR U3153 ( .A(n3113), .B(n3114), .Z(n2971) );
  AND U3154 ( .A(n150), .B(n3115), .Z(n3114) );
  XNOR U3155 ( .A(n3116), .B(n3113), .Z(n3115) );
  XNOR U3156 ( .A(n3117), .B(n3118), .Z(n150) );
  AND U3157 ( .A(n3119), .B(n3120), .Z(n3118) );
  XOR U3158 ( .A(n3072), .B(n3117), .Z(n3120) );
  AND U3159 ( .A(n3121), .B(n3122), .Z(n3072) );
  XNOR U3160 ( .A(n3069), .B(n3117), .Z(n3119) );
  XNOR U3161 ( .A(n3123), .B(n3124), .Z(n3069) );
  AND U3162 ( .A(n3125), .B(n154), .Z(n3124) );
  XOR U3163 ( .A(n3126), .B(n3127), .Z(n3117) );
  AND U3164 ( .A(n3128), .B(n3129), .Z(n3127) );
  XNOR U3165 ( .A(n3126), .B(n3121), .Z(n3129) );
  IV U3166 ( .A(n3082), .Z(n3121) );
  XOR U3167 ( .A(n3130), .B(n3131), .Z(n3082) );
  XOR U3168 ( .A(n3132), .B(n3122), .Z(n3131) );
  AND U3169 ( .A(n3092), .B(n3133), .Z(n3122) );
  AND U3170 ( .A(n3134), .B(n3135), .Z(n3132) );
  XOR U3171 ( .A(n3136), .B(n3130), .Z(n3134) );
  XNOR U3172 ( .A(n3079), .B(n3126), .Z(n3128) );
  XNOR U3173 ( .A(n3137), .B(n3138), .Z(n3079) );
  AND U3174 ( .A(n154), .B(n3139), .Z(n3138) );
  XNOR U3175 ( .A(n3140), .B(n3141), .Z(n3139) );
  XOR U3176 ( .A(n3142), .B(n3143), .Z(n3126) );
  AND U3177 ( .A(n3144), .B(n3145), .Z(n3143) );
  XNOR U3178 ( .A(n3142), .B(n3092), .Z(n3145) );
  XOR U3179 ( .A(n3146), .B(n3135), .Z(n3092) );
  XNOR U3180 ( .A(n3147), .B(n3130), .Z(n3135) );
  XOR U3181 ( .A(n3148), .B(n3149), .Z(n3130) );
  AND U3182 ( .A(n3150), .B(n3151), .Z(n3149) );
  XOR U3183 ( .A(n3152), .B(n3148), .Z(n3150) );
  XNOR U3184 ( .A(n3153), .B(n3154), .Z(n3147) );
  AND U3185 ( .A(n3155), .B(n3156), .Z(n3154) );
  XOR U3186 ( .A(n3153), .B(n3157), .Z(n3155) );
  XNOR U3187 ( .A(n3136), .B(n3133), .Z(n3146) );
  AND U3188 ( .A(n3158), .B(n3159), .Z(n3133) );
  XOR U3189 ( .A(n3160), .B(n3161), .Z(n3136) );
  AND U3190 ( .A(n3162), .B(n3163), .Z(n3161) );
  XOR U3191 ( .A(n3160), .B(n3164), .Z(n3162) );
  XNOR U3192 ( .A(n3089), .B(n3142), .Z(n3144) );
  XNOR U3193 ( .A(n3165), .B(n3166), .Z(n3089) );
  AND U3194 ( .A(n154), .B(n3167), .Z(n3166) );
  XNOR U3195 ( .A(n3168), .B(n3169), .Z(n3167) );
  XOR U3196 ( .A(n3170), .B(n3171), .Z(n3142) );
  AND U3197 ( .A(n3172), .B(n3173), .Z(n3171) );
  XNOR U3198 ( .A(n3170), .B(n3158), .Z(n3173) );
  IV U3199 ( .A(n3102), .Z(n3158) );
  XNOR U3200 ( .A(n3174), .B(n3151), .Z(n3102) );
  XNOR U3201 ( .A(n3175), .B(n3157), .Z(n3151) );
  XOR U3202 ( .A(n3176), .B(n3177), .Z(n3157) );
  AND U3203 ( .A(n3178), .B(n3179), .Z(n3177) );
  XOR U3204 ( .A(n3176), .B(n3180), .Z(n3178) );
  XNOR U3205 ( .A(n3156), .B(n3148), .Z(n3175) );
  XOR U3206 ( .A(n3181), .B(n3182), .Z(n3148) );
  AND U3207 ( .A(n3183), .B(n3184), .Z(n3182) );
  XNOR U3208 ( .A(n3185), .B(n3181), .Z(n3183) );
  XNOR U3209 ( .A(n3186), .B(n3153), .Z(n3156) );
  XOR U3210 ( .A(n3187), .B(n3188), .Z(n3153) );
  AND U3211 ( .A(n3189), .B(n3190), .Z(n3188) );
  XOR U3212 ( .A(n3187), .B(n3191), .Z(n3189) );
  XNOR U3213 ( .A(n3192), .B(n3193), .Z(n3186) );
  AND U3214 ( .A(n3194), .B(n3195), .Z(n3193) );
  XNOR U3215 ( .A(n3192), .B(n3196), .Z(n3194) );
  XNOR U3216 ( .A(n3152), .B(n3159), .Z(n3174) );
  AND U3217 ( .A(n3110), .B(n3197), .Z(n3159) );
  XOR U3218 ( .A(n3164), .B(n3163), .Z(n3152) );
  XNOR U3219 ( .A(n3198), .B(n3160), .Z(n3163) );
  XOR U3220 ( .A(n3199), .B(n3200), .Z(n3160) );
  AND U3221 ( .A(n3201), .B(n3202), .Z(n3200) );
  XOR U3222 ( .A(n3199), .B(n3203), .Z(n3201) );
  XNOR U3223 ( .A(n3204), .B(n3205), .Z(n3198) );
  AND U3224 ( .A(n3206), .B(n3207), .Z(n3205) );
  XOR U3225 ( .A(n3204), .B(n3208), .Z(n3206) );
  XOR U3226 ( .A(n3209), .B(n3210), .Z(n3164) );
  AND U3227 ( .A(n3211), .B(n3212), .Z(n3210) );
  XOR U3228 ( .A(n3209), .B(n3213), .Z(n3211) );
  XNOR U3229 ( .A(n3099), .B(n3170), .Z(n3172) );
  XNOR U3230 ( .A(n3214), .B(n3215), .Z(n3099) );
  AND U3231 ( .A(n154), .B(n3216), .Z(n3215) );
  XNOR U3232 ( .A(n3217), .B(n3218), .Z(n3216) );
  XOR U3233 ( .A(n3219), .B(n3220), .Z(n3170) );
  AND U3234 ( .A(n3221), .B(n3222), .Z(n3220) );
  XNOR U3235 ( .A(n3219), .B(n3110), .Z(n3222) );
  XOR U3236 ( .A(n3223), .B(n3184), .Z(n3110) );
  XNOR U3237 ( .A(n3224), .B(n3191), .Z(n3184) );
  XOR U3238 ( .A(n3180), .B(n3179), .Z(n3191) );
  XNOR U3239 ( .A(n3225), .B(n3176), .Z(n3179) );
  XOR U3240 ( .A(n3226), .B(n3227), .Z(n3176) );
  AND U3241 ( .A(n3228), .B(n3229), .Z(n3227) );
  XOR U3242 ( .A(n3226), .B(n3230), .Z(n3228) );
  XNOR U3243 ( .A(n3231), .B(n3232), .Z(n3225) );
  NOR U3244 ( .A(n3233), .B(n3234), .Z(n3232) );
  XNOR U3245 ( .A(n3231), .B(n3235), .Z(n3233) );
  XOR U3246 ( .A(n3236), .B(n3237), .Z(n3180) );
  NOR U3247 ( .A(n3238), .B(n3239), .Z(n3237) );
  XNOR U3248 ( .A(n3236), .B(n3240), .Z(n3238) );
  XNOR U3249 ( .A(n3190), .B(n3181), .Z(n3224) );
  XOR U3250 ( .A(n3241), .B(n3242), .Z(n3181) );
  NOR U3251 ( .A(n3243), .B(n3244), .Z(n3242) );
  XNOR U3252 ( .A(n3241), .B(n3245), .Z(n3243) );
  XOR U3253 ( .A(n3246), .B(n3196), .Z(n3190) );
  XNOR U3254 ( .A(n3247), .B(n3248), .Z(n3196) );
  NOR U3255 ( .A(n3249), .B(n3250), .Z(n3248) );
  XNOR U3256 ( .A(n3247), .B(n3251), .Z(n3249) );
  XNOR U3257 ( .A(n3195), .B(n3187), .Z(n3246) );
  XOR U3258 ( .A(n3252), .B(n3253), .Z(n3187) );
  AND U3259 ( .A(n3254), .B(n3255), .Z(n3253) );
  XOR U3260 ( .A(n3252), .B(n3256), .Z(n3254) );
  XNOR U3261 ( .A(n3257), .B(n3192), .Z(n3195) );
  XOR U3262 ( .A(n3258), .B(n3259), .Z(n3192) );
  AND U3263 ( .A(n3260), .B(n3261), .Z(n3259) );
  XOR U3264 ( .A(n3258), .B(n3262), .Z(n3260) );
  XNOR U3265 ( .A(n3263), .B(n3264), .Z(n3257) );
  NOR U3266 ( .A(n3265), .B(n3266), .Z(n3264) );
  XOR U3267 ( .A(n3263), .B(n3267), .Z(n3265) );
  XOR U3268 ( .A(n3185), .B(n3197), .Z(n3223) );
  NOR U3269 ( .A(n3116), .B(n3268), .Z(n3197) );
  XNOR U3270 ( .A(n3203), .B(n3202), .Z(n3185) );
  XNOR U3271 ( .A(n3269), .B(n3208), .Z(n3202) );
  XOR U3272 ( .A(n3270), .B(n3271), .Z(n3208) );
  NOR U3273 ( .A(n3272), .B(n3273), .Z(n3271) );
  XNOR U3274 ( .A(n3270), .B(n3274), .Z(n3272) );
  XNOR U3275 ( .A(n3207), .B(n3199), .Z(n3269) );
  XOR U3276 ( .A(n3275), .B(n3276), .Z(n3199) );
  AND U3277 ( .A(n3277), .B(n3278), .Z(n3276) );
  XNOR U3278 ( .A(n3275), .B(n3279), .Z(n3277) );
  XNOR U3279 ( .A(n3280), .B(n3204), .Z(n3207) );
  XOR U3280 ( .A(n3281), .B(n3282), .Z(n3204) );
  AND U3281 ( .A(n3283), .B(n3284), .Z(n3282) );
  XOR U3282 ( .A(n3281), .B(n3285), .Z(n3283) );
  XNOR U3283 ( .A(n3286), .B(n3287), .Z(n3280) );
  NOR U3284 ( .A(n3288), .B(n3289), .Z(n3287) );
  XOR U3285 ( .A(n3286), .B(n3290), .Z(n3288) );
  XOR U3286 ( .A(n3213), .B(n3212), .Z(n3203) );
  XNOR U3287 ( .A(n3291), .B(n3209), .Z(n3212) );
  XOR U3288 ( .A(n3292), .B(n3293), .Z(n3209) );
  AND U3289 ( .A(n3294), .B(n3295), .Z(n3293) );
  XOR U3290 ( .A(n3292), .B(n3296), .Z(n3294) );
  XNOR U3291 ( .A(n3297), .B(n3298), .Z(n3291) );
  NOR U3292 ( .A(n3299), .B(n3300), .Z(n3298) );
  XNOR U3293 ( .A(n3297), .B(n3301), .Z(n3299) );
  XOR U3294 ( .A(n3302), .B(n3303), .Z(n3213) );
  NOR U3295 ( .A(n3304), .B(n3305), .Z(n3303) );
  XNOR U3296 ( .A(n3302), .B(n3306), .Z(n3304) );
  XNOR U3297 ( .A(n3107), .B(n3219), .Z(n3221) );
  XNOR U3298 ( .A(n3307), .B(n3308), .Z(n3107) );
  AND U3299 ( .A(n154), .B(n3309), .Z(n3308) );
  XNOR U3300 ( .A(n3310), .B(n3311), .Z(n3309) );
  AND U3301 ( .A(n3113), .B(n3116), .Z(n3219) );
  XOR U3302 ( .A(n3312), .B(n3268), .Z(n3116) );
  XNOR U3303 ( .A(p_input[256]), .B(p_input[32]), .Z(n3268) );
  XOR U3304 ( .A(n3245), .B(n3244), .Z(n3312) );
  XOR U3305 ( .A(n3313), .B(n3256), .Z(n3244) );
  XOR U3306 ( .A(n3230), .B(n3229), .Z(n3256) );
  XNOR U3307 ( .A(n3314), .B(n3235), .Z(n3229) );
  XOR U3308 ( .A(p_input[280]), .B(p_input[56]), .Z(n3235) );
  XOR U3309 ( .A(n3226), .B(n3234), .Z(n3314) );
  XOR U3310 ( .A(n3315), .B(n3231), .Z(n3234) );
  XOR U3311 ( .A(p_input[278]), .B(p_input[54]), .Z(n3231) );
  XNOR U3312 ( .A(p_input[279]), .B(p_input[55]), .Z(n3315) );
  XNOR U3313 ( .A(n3316), .B(p_input[50]), .Z(n3226) );
  XNOR U3314 ( .A(n3240), .B(n3239), .Z(n3230) );
  XOR U3315 ( .A(n3317), .B(n3236), .Z(n3239) );
  XOR U3316 ( .A(p_input[275]), .B(p_input[51]), .Z(n3236) );
  XNOR U3317 ( .A(p_input[276]), .B(p_input[52]), .Z(n3317) );
  XOR U3318 ( .A(p_input[277]), .B(p_input[53]), .Z(n3240) );
  XNOR U3319 ( .A(n3255), .B(n3241), .Z(n3313) );
  XNOR U3320 ( .A(n3318), .B(p_input[33]), .Z(n3241) );
  XNOR U3321 ( .A(n3319), .B(n3262), .Z(n3255) );
  XNOR U3322 ( .A(n3251), .B(n3250), .Z(n3262) );
  XOR U3323 ( .A(n3320), .B(n3247), .Z(n3250) );
  XNOR U3324 ( .A(n3321), .B(p_input[58]), .Z(n3247) );
  XNOR U3325 ( .A(p_input[283]), .B(p_input[59]), .Z(n3320) );
  XOR U3326 ( .A(p_input[284]), .B(p_input[60]), .Z(n3251) );
  XNOR U3327 ( .A(n3261), .B(n3252), .Z(n3319) );
  XNOR U3328 ( .A(n3322), .B(p_input[49]), .Z(n3252) );
  XOR U3329 ( .A(n3323), .B(n3267), .Z(n3261) );
  XNOR U3330 ( .A(p_input[287]), .B(p_input[63]), .Z(n3267) );
  XOR U3331 ( .A(n3258), .B(n3266), .Z(n3323) );
  XOR U3332 ( .A(n3324), .B(n3263), .Z(n3266) );
  XOR U3333 ( .A(p_input[285]), .B(p_input[61]), .Z(n3263) );
  XNOR U3334 ( .A(p_input[286]), .B(p_input[62]), .Z(n3324) );
  XNOR U3335 ( .A(n3325), .B(p_input[57]), .Z(n3258) );
  XNOR U3336 ( .A(n3279), .B(n3278), .Z(n3245) );
  XNOR U3337 ( .A(n3326), .B(n3285), .Z(n3278) );
  XNOR U3338 ( .A(n3274), .B(n3273), .Z(n3285) );
  XOR U3339 ( .A(n3327), .B(n3270), .Z(n3273) );
  XNOR U3340 ( .A(n3328), .B(p_input[43]), .Z(n3270) );
  XNOR U3341 ( .A(p_input[268]), .B(p_input[44]), .Z(n3327) );
  XOR U3342 ( .A(p_input[269]), .B(p_input[45]), .Z(n3274) );
  XNOR U3343 ( .A(n3284), .B(n3275), .Z(n3326) );
  XOR U3344 ( .A(p_input[258]), .B(p_input[34]), .Z(n3275) );
  XOR U3345 ( .A(n3329), .B(n3290), .Z(n3284) );
  XNOR U3346 ( .A(p_input[272]), .B(p_input[48]), .Z(n3290) );
  XOR U3347 ( .A(n3281), .B(n3289), .Z(n3329) );
  XOR U3348 ( .A(n3330), .B(n3286), .Z(n3289) );
  XOR U3349 ( .A(p_input[270]), .B(p_input[46]), .Z(n3286) );
  XNOR U3350 ( .A(p_input[271]), .B(p_input[47]), .Z(n3330) );
  XNOR U3351 ( .A(n3331), .B(p_input[42]), .Z(n3281) );
  XNOR U3352 ( .A(n3296), .B(n3295), .Z(n3279) );
  XNOR U3353 ( .A(n3332), .B(n3301), .Z(n3295) );
  XOR U3354 ( .A(p_input[265]), .B(p_input[41]), .Z(n3301) );
  XOR U3355 ( .A(n3292), .B(n3300), .Z(n3332) );
  XOR U3356 ( .A(n3333), .B(n3297), .Z(n3300) );
  XOR U3357 ( .A(p_input[263]), .B(p_input[39]), .Z(n3297) );
  XNOR U3358 ( .A(p_input[264]), .B(p_input[40]), .Z(n3333) );
  XOR U3359 ( .A(p_input[259]), .B(p_input[35]), .Z(n3292) );
  XNOR U3360 ( .A(n3306), .B(n3305), .Z(n3296) );
  XOR U3361 ( .A(n3334), .B(n3302), .Z(n3305) );
  XOR U3362 ( .A(p_input[260]), .B(p_input[36]), .Z(n3302) );
  XNOR U3363 ( .A(p_input[261]), .B(p_input[37]), .Z(n3334) );
  XOR U3364 ( .A(p_input[262]), .B(p_input[38]), .Z(n3306) );
  XNOR U3365 ( .A(n3335), .B(n3336), .Z(n3113) );
  AND U3366 ( .A(n154), .B(n3337), .Z(n3336) );
  XNOR U3367 ( .A(n3338), .B(n3339), .Z(n154) );
  NOR U3368 ( .A(n3340), .B(n3341), .Z(n3339) );
  XNOR U3369 ( .A(n3342), .B(n3343), .Z(n3341) );
  AND U3370 ( .A(n3342), .B(n3123), .Z(n3340) );
  IV U3371 ( .A(n3338), .Z(n3342) );
  XOR U3372 ( .A(n3344), .B(n3345), .Z(n3338) );
  AND U3373 ( .A(n3346), .B(n3347), .Z(n3345) );
  XOR U3374 ( .A(n3140), .B(n3344), .Z(n3347) );
  XOR U3375 ( .A(n3344), .B(n3141), .Z(n3346) );
  XOR U3376 ( .A(n3348), .B(n3349), .Z(n3344) );
  AND U3377 ( .A(n3350), .B(n3351), .Z(n3349) );
  XOR U3378 ( .A(n3168), .B(n3348), .Z(n3351) );
  XOR U3379 ( .A(n3348), .B(n3169), .Z(n3350) );
  XOR U3380 ( .A(n3352), .B(n3353), .Z(n3348) );
  AND U3381 ( .A(n3354), .B(n3355), .Z(n3353) );
  XOR U3382 ( .A(n3217), .B(n3352), .Z(n3355) );
  XOR U3383 ( .A(n3352), .B(n3218), .Z(n3354) );
  XOR U3384 ( .A(n3356), .B(n3357), .Z(n3352) );
  AND U3385 ( .A(n3358), .B(n3359), .Z(n3357) );
  XOR U3386 ( .A(n3356), .B(n3310), .Z(n3359) );
  XNOR U3387 ( .A(n3360), .B(n3361), .Z(n3063) );
  AND U3388 ( .A(n158), .B(n3362), .Z(n3361) );
  XNOR U3389 ( .A(n3363), .B(n3364), .Z(n158) );
  AND U3390 ( .A(n3365), .B(n3366), .Z(n3364) );
  XNOR U3391 ( .A(n3363), .B(n3026), .Z(n3366) );
  XOR U3392 ( .A(n3363), .B(n3023), .Z(n3365) );
  XOR U3393 ( .A(n3367), .B(n3368), .Z(n3363) );
  AND U3394 ( .A(n3369), .B(n3370), .Z(n3368) );
  XNOR U3395 ( .A(n3083), .B(n3367), .Z(n3370) );
  XOR U3396 ( .A(n3367), .B(n3034), .Z(n3369) );
  XOR U3397 ( .A(n3371), .B(n3372), .Z(n3367) );
  AND U3398 ( .A(n3373), .B(n3374), .Z(n3372) );
  XNOR U3399 ( .A(n3093), .B(n3371), .Z(n3374) );
  XOR U3400 ( .A(n3371), .B(n3043), .Z(n3373) );
  XOR U3401 ( .A(n3375), .B(n3376), .Z(n3371) );
  AND U3402 ( .A(n3377), .B(n3378), .Z(n3376) );
  XOR U3403 ( .A(n3375), .B(n3050), .Z(n3377) );
  XOR U3404 ( .A(n3379), .B(n3380), .Z(n3014) );
  AND U3405 ( .A(n162), .B(n3362), .Z(n3380) );
  XNOR U3406 ( .A(n3360), .B(n3379), .Z(n3362) );
  XNOR U3407 ( .A(n3381), .B(n3382), .Z(n162) );
  AND U3408 ( .A(n3383), .B(n3384), .Z(n3382) );
  XNOR U3409 ( .A(n3026), .B(n3381), .Z(n3384) );
  XNOR U3410 ( .A(n3343), .B(n3385), .Z(n3026) );
  AND U3411 ( .A(n3125), .B(n165), .Z(n3385) );
  NOR U3412 ( .A(n3386), .B(n3387), .Z(n3125) );
  XOR U3413 ( .A(n3381), .B(n3023), .Z(n3383) );
  IV U3414 ( .A(n3027), .Z(n3023) );
  AND U3415 ( .A(n3388), .B(n3389), .Z(n3027) );
  XOR U3416 ( .A(n3390), .B(n3391), .Z(n3381) );
  AND U3417 ( .A(n3392), .B(n3393), .Z(n3391) );
  XNOR U3418 ( .A(n3390), .B(n3083), .Z(n3393) );
  XOR U3419 ( .A(n3141), .B(n3394), .Z(n3083) );
  AND U3420 ( .A(n165), .B(n3395), .Z(n3394) );
  XOR U3421 ( .A(n3137), .B(n3141), .Z(n3395) );
  XNOR U3422 ( .A(n3396), .B(n3390), .Z(n3392) );
  IV U3423 ( .A(n3034), .Z(n3396) );
  XOR U3424 ( .A(n3397), .B(n3398), .Z(n3034) );
  AND U3425 ( .A(n181), .B(n3399), .Z(n3398) );
  XOR U3426 ( .A(n3400), .B(n3401), .Z(n3390) );
  AND U3427 ( .A(n3402), .B(n3403), .Z(n3401) );
  XNOR U3428 ( .A(n3400), .B(n3093), .Z(n3403) );
  XOR U3429 ( .A(n3169), .B(n3404), .Z(n3093) );
  AND U3430 ( .A(n165), .B(n3405), .Z(n3404) );
  XOR U3431 ( .A(n3165), .B(n3169), .Z(n3405) );
  XOR U3432 ( .A(n3043), .B(n3400), .Z(n3402) );
  XOR U3433 ( .A(n3406), .B(n3407), .Z(n3043) );
  AND U3434 ( .A(n181), .B(n3408), .Z(n3407) );
  XOR U3435 ( .A(n3375), .B(n3409), .Z(n3400) );
  AND U3436 ( .A(n3410), .B(n3378), .Z(n3409) );
  XNOR U3437 ( .A(n3103), .B(n3375), .Z(n3378) );
  XOR U3438 ( .A(n3218), .B(n3411), .Z(n3103) );
  AND U3439 ( .A(n165), .B(n3412), .Z(n3411) );
  XOR U3440 ( .A(n3214), .B(n3218), .Z(n3412) );
  XNOR U3441 ( .A(n3413), .B(n3375), .Z(n3410) );
  IV U3442 ( .A(n3050), .Z(n3413) );
  XOR U3443 ( .A(n3414), .B(n3415), .Z(n3050) );
  AND U3444 ( .A(n181), .B(n3416), .Z(n3415) );
  XOR U3445 ( .A(n3417), .B(n3418), .Z(n3375) );
  AND U3446 ( .A(n3419), .B(n3420), .Z(n3418) );
  XNOR U3447 ( .A(n3417), .B(n3111), .Z(n3420) );
  XOR U3448 ( .A(n3311), .B(n3421), .Z(n3111) );
  AND U3449 ( .A(n165), .B(n3422), .Z(n3421) );
  XOR U3450 ( .A(n3307), .B(n3311), .Z(n3422) );
  XNOR U3451 ( .A(n3423), .B(n3417), .Z(n3419) );
  IV U3452 ( .A(n3060), .Z(n3423) );
  XOR U3453 ( .A(n3424), .B(n3425), .Z(n3060) );
  AND U3454 ( .A(n181), .B(n3426), .Z(n3425) );
  AND U3455 ( .A(n3379), .B(n3360), .Z(n3417) );
  XNOR U3456 ( .A(n3427), .B(n3428), .Z(n3360) );
  AND U3457 ( .A(n165), .B(n3337), .Z(n3428) );
  XNOR U3458 ( .A(n3335), .B(n3427), .Z(n3337) );
  XNOR U3459 ( .A(n3429), .B(n3430), .Z(n165) );
  NOR U3460 ( .A(n3431), .B(n3432), .Z(n3430) );
  XNOR U3461 ( .A(n3433), .B(n3343), .Z(n3432) );
  IV U3462 ( .A(n3387), .Z(n3343) );
  NOR U3463 ( .A(n3388), .B(n3389), .Z(n3387) );
  AND U3464 ( .A(n3433), .B(n3123), .Z(n3431) );
  IV U3465 ( .A(n3386), .Z(n3123) );
  AND U3466 ( .A(n3434), .B(n3435), .Z(n3386) );
  IV U3467 ( .A(n3436), .Z(n3434) );
  IV U3468 ( .A(n3429), .Z(n3433) );
  XOR U3469 ( .A(n3437), .B(n3438), .Z(n3429) );
  AND U3470 ( .A(n3439), .B(n3440), .Z(n3438) );
  XNOR U3471 ( .A(n3437), .B(n3137), .Z(n3440) );
  IV U3472 ( .A(n3140), .Z(n3137) );
  XOR U3473 ( .A(n3441), .B(n3442), .Z(n3140) );
  AND U3474 ( .A(n169), .B(n3443), .Z(n3442) );
  XOR U3475 ( .A(n3444), .B(n3441), .Z(n3443) );
  XOR U3476 ( .A(n3141), .B(n3437), .Z(n3439) );
  XOR U3477 ( .A(n3445), .B(n3446), .Z(n3141) );
  AND U3478 ( .A(n177), .B(n3399), .Z(n3446) );
  XOR U3479 ( .A(n3445), .B(n3397), .Z(n3399) );
  XOR U3480 ( .A(n3447), .B(n3448), .Z(n3437) );
  AND U3481 ( .A(n3449), .B(n3450), .Z(n3448) );
  XNOR U3482 ( .A(n3447), .B(n3165), .Z(n3450) );
  IV U3483 ( .A(n3168), .Z(n3165) );
  XOR U3484 ( .A(n3451), .B(n3452), .Z(n3168) );
  AND U3485 ( .A(n169), .B(n3453), .Z(n3452) );
  XNOR U3486 ( .A(n3454), .B(n3451), .Z(n3453) );
  XOR U3487 ( .A(n3169), .B(n3447), .Z(n3449) );
  XOR U3488 ( .A(n3455), .B(n3456), .Z(n3169) );
  AND U3489 ( .A(n177), .B(n3408), .Z(n3456) );
  XOR U3490 ( .A(n3455), .B(n3406), .Z(n3408) );
  XOR U3491 ( .A(n3457), .B(n3458), .Z(n3447) );
  AND U3492 ( .A(n3459), .B(n3460), .Z(n3458) );
  XNOR U3493 ( .A(n3457), .B(n3214), .Z(n3460) );
  IV U3494 ( .A(n3217), .Z(n3214) );
  XOR U3495 ( .A(n3461), .B(n3462), .Z(n3217) );
  AND U3496 ( .A(n169), .B(n3463), .Z(n3462) );
  XOR U3497 ( .A(n3464), .B(n3461), .Z(n3463) );
  XOR U3498 ( .A(n3218), .B(n3457), .Z(n3459) );
  XOR U3499 ( .A(n3465), .B(n3466), .Z(n3218) );
  AND U3500 ( .A(n177), .B(n3416), .Z(n3466) );
  XOR U3501 ( .A(n3465), .B(n3414), .Z(n3416) );
  XOR U3502 ( .A(n3356), .B(n3467), .Z(n3457) );
  AND U3503 ( .A(n3358), .B(n3468), .Z(n3467) );
  XNOR U3504 ( .A(n3356), .B(n3307), .Z(n3468) );
  IV U3505 ( .A(n3310), .Z(n3307) );
  XOR U3506 ( .A(n3469), .B(n3470), .Z(n3310) );
  AND U3507 ( .A(n169), .B(n3471), .Z(n3470) );
  XNOR U3508 ( .A(n3472), .B(n3469), .Z(n3471) );
  XOR U3509 ( .A(n3311), .B(n3356), .Z(n3358) );
  XOR U3510 ( .A(n3473), .B(n3474), .Z(n3311) );
  AND U3511 ( .A(n177), .B(n3426), .Z(n3474) );
  XOR U3512 ( .A(n3473), .B(n3424), .Z(n3426) );
  AND U3513 ( .A(n3427), .B(n3335), .Z(n3356) );
  XNOR U3514 ( .A(n3475), .B(n3476), .Z(n3335) );
  AND U3515 ( .A(n169), .B(n3477), .Z(n3476) );
  XNOR U3516 ( .A(n3478), .B(n3475), .Z(n3477) );
  XNOR U3517 ( .A(n3479), .B(n3480), .Z(n169) );
  NOR U3518 ( .A(n3481), .B(n3482), .Z(n3480) );
  XNOR U3519 ( .A(n3479), .B(n3436), .Z(n3482) );
  NOR U3520 ( .A(n3483), .B(n3484), .Z(n3436) );
  NOR U3521 ( .A(n3479), .B(n3435), .Z(n3481) );
  AND U3522 ( .A(n3485), .B(n3486), .Z(n3435) );
  XOR U3523 ( .A(n3487), .B(n3488), .Z(n3479) );
  AND U3524 ( .A(n3489), .B(n3490), .Z(n3488) );
  XNOR U3525 ( .A(n3487), .B(n3485), .Z(n3490) );
  IV U3526 ( .A(n3444), .Z(n3485) );
  XOR U3527 ( .A(n3491), .B(n3492), .Z(n3444) );
  XOR U3528 ( .A(n3493), .B(n3486), .Z(n3492) );
  AND U3529 ( .A(n3454), .B(n3494), .Z(n3486) );
  AND U3530 ( .A(n3495), .B(n3496), .Z(n3493) );
  XOR U3531 ( .A(n3497), .B(n3491), .Z(n3495) );
  XNOR U3532 ( .A(n3441), .B(n3487), .Z(n3489) );
  XNOR U3533 ( .A(n3498), .B(n3499), .Z(n3441) );
  AND U3534 ( .A(n173), .B(n3500), .Z(n3499) );
  XNOR U3535 ( .A(n3501), .B(n3502), .Z(n3500) );
  XOR U3536 ( .A(n3503), .B(n3504), .Z(n3487) );
  AND U3537 ( .A(n3505), .B(n3506), .Z(n3504) );
  XNOR U3538 ( .A(n3503), .B(n3454), .Z(n3506) );
  XOR U3539 ( .A(n3507), .B(n3496), .Z(n3454) );
  XNOR U3540 ( .A(n3508), .B(n3491), .Z(n3496) );
  XOR U3541 ( .A(n3509), .B(n3510), .Z(n3491) );
  AND U3542 ( .A(n3511), .B(n3512), .Z(n3510) );
  XOR U3543 ( .A(n3513), .B(n3509), .Z(n3511) );
  XNOR U3544 ( .A(n3514), .B(n3515), .Z(n3508) );
  AND U3545 ( .A(n3516), .B(n3517), .Z(n3515) );
  XOR U3546 ( .A(n3514), .B(n3518), .Z(n3516) );
  XNOR U3547 ( .A(n3497), .B(n3494), .Z(n3507) );
  AND U3548 ( .A(n3519), .B(n3520), .Z(n3494) );
  XOR U3549 ( .A(n3521), .B(n3522), .Z(n3497) );
  AND U3550 ( .A(n3523), .B(n3524), .Z(n3522) );
  XOR U3551 ( .A(n3521), .B(n3525), .Z(n3523) );
  XNOR U3552 ( .A(n3451), .B(n3503), .Z(n3505) );
  XNOR U3553 ( .A(n3526), .B(n3527), .Z(n3451) );
  AND U3554 ( .A(n173), .B(n3528), .Z(n3527) );
  XNOR U3555 ( .A(n3529), .B(n3530), .Z(n3528) );
  XOR U3556 ( .A(n3531), .B(n3532), .Z(n3503) );
  AND U3557 ( .A(n3533), .B(n3534), .Z(n3532) );
  XNOR U3558 ( .A(n3531), .B(n3519), .Z(n3534) );
  IV U3559 ( .A(n3464), .Z(n3519) );
  XNOR U3560 ( .A(n3535), .B(n3512), .Z(n3464) );
  XNOR U3561 ( .A(n3536), .B(n3518), .Z(n3512) );
  XOR U3562 ( .A(n3537), .B(n3538), .Z(n3518) );
  AND U3563 ( .A(n3539), .B(n3540), .Z(n3538) );
  XOR U3564 ( .A(n3537), .B(n3541), .Z(n3539) );
  XNOR U3565 ( .A(n3517), .B(n3509), .Z(n3536) );
  XOR U3566 ( .A(n3542), .B(n3543), .Z(n3509) );
  AND U3567 ( .A(n3544), .B(n3545), .Z(n3543) );
  XNOR U3568 ( .A(n3546), .B(n3542), .Z(n3544) );
  XNOR U3569 ( .A(n3547), .B(n3514), .Z(n3517) );
  XOR U3570 ( .A(n3548), .B(n3549), .Z(n3514) );
  AND U3571 ( .A(n3550), .B(n3551), .Z(n3549) );
  XOR U3572 ( .A(n3548), .B(n3552), .Z(n3550) );
  XNOR U3573 ( .A(n3553), .B(n3554), .Z(n3547) );
  AND U3574 ( .A(n3555), .B(n3556), .Z(n3554) );
  XNOR U3575 ( .A(n3553), .B(n3557), .Z(n3555) );
  XNOR U3576 ( .A(n3513), .B(n3520), .Z(n3535) );
  AND U3577 ( .A(n3472), .B(n3558), .Z(n3520) );
  XOR U3578 ( .A(n3525), .B(n3524), .Z(n3513) );
  XNOR U3579 ( .A(n3559), .B(n3521), .Z(n3524) );
  XOR U3580 ( .A(n3560), .B(n3561), .Z(n3521) );
  AND U3581 ( .A(n3562), .B(n3563), .Z(n3561) );
  XOR U3582 ( .A(n3560), .B(n3564), .Z(n3562) );
  XNOR U3583 ( .A(n3565), .B(n3566), .Z(n3559) );
  AND U3584 ( .A(n3567), .B(n3568), .Z(n3566) );
  XOR U3585 ( .A(n3565), .B(n3569), .Z(n3567) );
  XOR U3586 ( .A(n3570), .B(n3571), .Z(n3525) );
  AND U3587 ( .A(n3572), .B(n3573), .Z(n3571) );
  XOR U3588 ( .A(n3570), .B(n3574), .Z(n3572) );
  XNOR U3589 ( .A(n3461), .B(n3531), .Z(n3533) );
  XNOR U3590 ( .A(n3575), .B(n3576), .Z(n3461) );
  AND U3591 ( .A(n173), .B(n3577), .Z(n3576) );
  XNOR U3592 ( .A(n3578), .B(n3579), .Z(n3577) );
  XOR U3593 ( .A(n3580), .B(n3581), .Z(n3531) );
  AND U3594 ( .A(n3582), .B(n3583), .Z(n3581) );
  XNOR U3595 ( .A(n3580), .B(n3472), .Z(n3583) );
  XOR U3596 ( .A(n3584), .B(n3545), .Z(n3472) );
  XNOR U3597 ( .A(n3585), .B(n3552), .Z(n3545) );
  XOR U3598 ( .A(n3541), .B(n3540), .Z(n3552) );
  XNOR U3599 ( .A(n3586), .B(n3537), .Z(n3540) );
  XOR U3600 ( .A(n3587), .B(n3588), .Z(n3537) );
  AND U3601 ( .A(n3589), .B(n3590), .Z(n3588) );
  XOR U3602 ( .A(n3587), .B(n3591), .Z(n3589) );
  XNOR U3603 ( .A(n3592), .B(n3593), .Z(n3586) );
  NOR U3604 ( .A(n3594), .B(n3595), .Z(n3593) );
  XNOR U3605 ( .A(n3592), .B(n3596), .Z(n3594) );
  XOR U3606 ( .A(n3597), .B(n3598), .Z(n3541) );
  NOR U3607 ( .A(n3599), .B(n3600), .Z(n3598) );
  XNOR U3608 ( .A(n3597), .B(n3601), .Z(n3599) );
  XNOR U3609 ( .A(n3551), .B(n3542), .Z(n3585) );
  XOR U3610 ( .A(n3602), .B(n3603), .Z(n3542) );
  NOR U3611 ( .A(n3604), .B(n3605), .Z(n3603) );
  XNOR U3612 ( .A(n3602), .B(n3606), .Z(n3604) );
  XOR U3613 ( .A(n3607), .B(n3557), .Z(n3551) );
  XNOR U3614 ( .A(n3608), .B(n3609), .Z(n3557) );
  NOR U3615 ( .A(n3610), .B(n3611), .Z(n3609) );
  XNOR U3616 ( .A(n3608), .B(n3612), .Z(n3610) );
  XNOR U3617 ( .A(n3556), .B(n3548), .Z(n3607) );
  XOR U3618 ( .A(n3613), .B(n3614), .Z(n3548) );
  AND U3619 ( .A(n3615), .B(n3616), .Z(n3614) );
  XOR U3620 ( .A(n3613), .B(n3617), .Z(n3615) );
  XNOR U3621 ( .A(n3618), .B(n3553), .Z(n3556) );
  XOR U3622 ( .A(n3619), .B(n3620), .Z(n3553) );
  AND U3623 ( .A(n3621), .B(n3622), .Z(n3620) );
  XOR U3624 ( .A(n3619), .B(n3623), .Z(n3621) );
  XNOR U3625 ( .A(n3624), .B(n3625), .Z(n3618) );
  NOR U3626 ( .A(n3626), .B(n3627), .Z(n3625) );
  XOR U3627 ( .A(n3624), .B(n3628), .Z(n3626) );
  XOR U3628 ( .A(n3546), .B(n3558), .Z(n3584) );
  NOR U3629 ( .A(n3478), .B(n3629), .Z(n3558) );
  XNOR U3630 ( .A(n3564), .B(n3563), .Z(n3546) );
  XNOR U3631 ( .A(n3630), .B(n3569), .Z(n3563) );
  XOR U3632 ( .A(n3631), .B(n3632), .Z(n3569) );
  NOR U3633 ( .A(n3633), .B(n3634), .Z(n3632) );
  XNOR U3634 ( .A(n3631), .B(n3635), .Z(n3633) );
  XNOR U3635 ( .A(n3568), .B(n3560), .Z(n3630) );
  XOR U3636 ( .A(n3636), .B(n3637), .Z(n3560) );
  AND U3637 ( .A(n3638), .B(n3639), .Z(n3637) );
  XNOR U3638 ( .A(n3636), .B(n3640), .Z(n3638) );
  XNOR U3639 ( .A(n3641), .B(n3565), .Z(n3568) );
  XOR U3640 ( .A(n3642), .B(n3643), .Z(n3565) );
  AND U3641 ( .A(n3644), .B(n3645), .Z(n3643) );
  XOR U3642 ( .A(n3642), .B(n3646), .Z(n3644) );
  XNOR U3643 ( .A(n3647), .B(n3648), .Z(n3641) );
  NOR U3644 ( .A(n3649), .B(n3650), .Z(n3648) );
  XOR U3645 ( .A(n3647), .B(n3651), .Z(n3649) );
  XOR U3646 ( .A(n3574), .B(n3573), .Z(n3564) );
  XNOR U3647 ( .A(n3652), .B(n3570), .Z(n3573) );
  XOR U3648 ( .A(n3653), .B(n3654), .Z(n3570) );
  AND U3649 ( .A(n3655), .B(n3656), .Z(n3654) );
  XOR U3650 ( .A(n3653), .B(n3657), .Z(n3655) );
  XNOR U3651 ( .A(n3658), .B(n3659), .Z(n3652) );
  NOR U3652 ( .A(n3660), .B(n3661), .Z(n3659) );
  XNOR U3653 ( .A(n3658), .B(n3662), .Z(n3660) );
  XOR U3654 ( .A(n3663), .B(n3664), .Z(n3574) );
  NOR U3655 ( .A(n3665), .B(n3666), .Z(n3664) );
  XNOR U3656 ( .A(n3663), .B(n3667), .Z(n3665) );
  XNOR U3657 ( .A(n3469), .B(n3580), .Z(n3582) );
  XNOR U3658 ( .A(n3668), .B(n3669), .Z(n3469) );
  AND U3659 ( .A(n173), .B(n3670), .Z(n3669) );
  XNOR U3660 ( .A(n3671), .B(n3672), .Z(n3670) );
  AND U3661 ( .A(n3475), .B(n3478), .Z(n3580) );
  XOR U3662 ( .A(n3673), .B(n3629), .Z(n3478) );
  XNOR U3663 ( .A(p_input[256]), .B(p_input[64]), .Z(n3629) );
  XOR U3664 ( .A(n3606), .B(n3605), .Z(n3673) );
  XOR U3665 ( .A(n3674), .B(n3617), .Z(n3605) );
  XOR U3666 ( .A(n3591), .B(n3590), .Z(n3617) );
  XNOR U3667 ( .A(n3675), .B(n3596), .Z(n3590) );
  XOR U3668 ( .A(p_input[280]), .B(p_input[88]), .Z(n3596) );
  XOR U3669 ( .A(n3587), .B(n3595), .Z(n3675) );
  XOR U3670 ( .A(n3676), .B(n3592), .Z(n3595) );
  XOR U3671 ( .A(p_input[278]), .B(p_input[86]), .Z(n3592) );
  XNOR U3672 ( .A(p_input[279]), .B(p_input[87]), .Z(n3676) );
  XNOR U3673 ( .A(n3316), .B(p_input[82]), .Z(n3587) );
  XNOR U3674 ( .A(n3601), .B(n3600), .Z(n3591) );
  XOR U3675 ( .A(n3677), .B(n3597), .Z(n3600) );
  XOR U3676 ( .A(p_input[275]), .B(p_input[83]), .Z(n3597) );
  XNOR U3677 ( .A(p_input[276]), .B(p_input[84]), .Z(n3677) );
  XOR U3678 ( .A(p_input[277]), .B(p_input[85]), .Z(n3601) );
  XNOR U3679 ( .A(n3616), .B(n3602), .Z(n3674) );
  XNOR U3680 ( .A(n3318), .B(p_input[65]), .Z(n3602) );
  XNOR U3681 ( .A(n3678), .B(n3623), .Z(n3616) );
  XNOR U3682 ( .A(n3612), .B(n3611), .Z(n3623) );
  XOR U3683 ( .A(n3679), .B(n3608), .Z(n3611) );
  XNOR U3684 ( .A(n3321), .B(p_input[90]), .Z(n3608) );
  XNOR U3685 ( .A(p_input[283]), .B(p_input[91]), .Z(n3679) );
  XOR U3686 ( .A(p_input[284]), .B(p_input[92]), .Z(n3612) );
  XNOR U3687 ( .A(n3622), .B(n3613), .Z(n3678) );
  XNOR U3688 ( .A(n3322), .B(p_input[81]), .Z(n3613) );
  XOR U3689 ( .A(n3680), .B(n3628), .Z(n3622) );
  XNOR U3690 ( .A(p_input[287]), .B(p_input[95]), .Z(n3628) );
  XOR U3691 ( .A(n3619), .B(n3627), .Z(n3680) );
  XOR U3692 ( .A(n3681), .B(n3624), .Z(n3627) );
  XOR U3693 ( .A(p_input[285]), .B(p_input[93]), .Z(n3624) );
  XNOR U3694 ( .A(p_input[286]), .B(p_input[94]), .Z(n3681) );
  XNOR U3695 ( .A(n3325), .B(p_input[89]), .Z(n3619) );
  XNOR U3696 ( .A(n3640), .B(n3639), .Z(n3606) );
  XNOR U3697 ( .A(n3682), .B(n3646), .Z(n3639) );
  XNOR U3698 ( .A(n3635), .B(n3634), .Z(n3646) );
  XOR U3699 ( .A(n3683), .B(n3631), .Z(n3634) );
  XNOR U3700 ( .A(n3328), .B(p_input[75]), .Z(n3631) );
  XNOR U3701 ( .A(p_input[268]), .B(p_input[76]), .Z(n3683) );
  XOR U3702 ( .A(p_input[269]), .B(p_input[77]), .Z(n3635) );
  XNOR U3703 ( .A(n3645), .B(n3636), .Z(n3682) );
  XOR U3704 ( .A(p_input[258]), .B(p_input[66]), .Z(n3636) );
  XOR U3705 ( .A(n3684), .B(n3651), .Z(n3645) );
  XNOR U3706 ( .A(p_input[272]), .B(p_input[80]), .Z(n3651) );
  XOR U3707 ( .A(n3642), .B(n3650), .Z(n3684) );
  XOR U3708 ( .A(n3685), .B(n3647), .Z(n3650) );
  XOR U3709 ( .A(p_input[270]), .B(p_input[78]), .Z(n3647) );
  XNOR U3710 ( .A(p_input[271]), .B(p_input[79]), .Z(n3685) );
  XNOR U3711 ( .A(n3331), .B(p_input[74]), .Z(n3642) );
  XNOR U3712 ( .A(n3657), .B(n3656), .Z(n3640) );
  XNOR U3713 ( .A(n3686), .B(n3662), .Z(n3656) );
  XOR U3714 ( .A(p_input[265]), .B(p_input[73]), .Z(n3662) );
  XOR U3715 ( .A(n3653), .B(n3661), .Z(n3686) );
  XOR U3716 ( .A(n3687), .B(n3658), .Z(n3661) );
  XOR U3717 ( .A(p_input[263]), .B(p_input[71]), .Z(n3658) );
  XNOR U3718 ( .A(p_input[264]), .B(p_input[72]), .Z(n3687) );
  XOR U3719 ( .A(p_input[259]), .B(p_input[67]), .Z(n3653) );
  XNOR U3720 ( .A(n3667), .B(n3666), .Z(n3657) );
  XOR U3721 ( .A(n3688), .B(n3663), .Z(n3666) );
  XOR U3722 ( .A(p_input[260]), .B(p_input[68]), .Z(n3663) );
  XNOR U3723 ( .A(p_input[261]), .B(p_input[69]), .Z(n3688) );
  XOR U3724 ( .A(p_input[262]), .B(p_input[70]), .Z(n3667) );
  XNOR U3725 ( .A(n3689), .B(n3690), .Z(n3475) );
  AND U3726 ( .A(n173), .B(n3691), .Z(n3690) );
  XNOR U3727 ( .A(n3692), .B(n3693), .Z(n173) );
  NOR U3728 ( .A(n3694), .B(n3695), .Z(n3693) );
  XNOR U3729 ( .A(n3692), .B(n3696), .Z(n3695) );
  NOR U3730 ( .A(n3692), .B(n3484), .Z(n3694) );
  XOR U3731 ( .A(n3697), .B(n3698), .Z(n3692) );
  AND U3732 ( .A(n3699), .B(n3700), .Z(n3698) );
  XOR U3733 ( .A(n3501), .B(n3697), .Z(n3700) );
  XOR U3734 ( .A(n3697), .B(n3502), .Z(n3699) );
  XOR U3735 ( .A(n3701), .B(n3702), .Z(n3697) );
  AND U3736 ( .A(n3703), .B(n3704), .Z(n3702) );
  XOR U3737 ( .A(n3529), .B(n3701), .Z(n3704) );
  XOR U3738 ( .A(n3701), .B(n3530), .Z(n3703) );
  XOR U3739 ( .A(n3705), .B(n3706), .Z(n3701) );
  AND U3740 ( .A(n3707), .B(n3708), .Z(n3706) );
  XOR U3741 ( .A(n3578), .B(n3705), .Z(n3708) );
  XOR U3742 ( .A(n3705), .B(n3579), .Z(n3707) );
  XOR U3743 ( .A(n3709), .B(n3710), .Z(n3705) );
  AND U3744 ( .A(n3711), .B(n3712), .Z(n3710) );
  XOR U3745 ( .A(n3709), .B(n3671), .Z(n3712) );
  XNOR U3746 ( .A(n3713), .B(n3714), .Z(n3427) );
  AND U3747 ( .A(n177), .B(n3715), .Z(n3714) );
  XNOR U3748 ( .A(n3716), .B(n3717), .Z(n177) );
  NOR U3749 ( .A(n3718), .B(n3719), .Z(n3717) );
  XOR U3750 ( .A(n3389), .B(n3716), .Z(n3719) );
  NOR U3751 ( .A(n3716), .B(n3388), .Z(n3718) );
  XOR U3752 ( .A(n3720), .B(n3721), .Z(n3716) );
  AND U3753 ( .A(n3722), .B(n3723), .Z(n3721) );
  XNOR U3754 ( .A(n3445), .B(n3720), .Z(n3723) );
  XOR U3755 ( .A(n3720), .B(n3397), .Z(n3722) );
  XOR U3756 ( .A(n3724), .B(n3725), .Z(n3720) );
  AND U3757 ( .A(n3726), .B(n3727), .Z(n3725) );
  XNOR U3758 ( .A(n3455), .B(n3724), .Z(n3727) );
  XOR U3759 ( .A(n3724), .B(n3406), .Z(n3726) );
  XOR U3760 ( .A(n3728), .B(n3729), .Z(n3724) );
  AND U3761 ( .A(n3730), .B(n3731), .Z(n3729) );
  XOR U3762 ( .A(n3728), .B(n3414), .Z(n3730) );
  XOR U3763 ( .A(n3732), .B(n3733), .Z(n3379) );
  AND U3764 ( .A(n181), .B(n3715), .Z(n3733) );
  XNOR U3765 ( .A(n3713), .B(n3732), .Z(n3715) );
  XNOR U3766 ( .A(n3734), .B(n3735), .Z(n181) );
  NOR U3767 ( .A(n3736), .B(n3737), .Z(n3735) );
  XNOR U3768 ( .A(n3389), .B(n3738), .Z(n3737) );
  IV U3769 ( .A(n3734), .Z(n3738) );
  AND U3770 ( .A(n3739), .B(n3740), .Z(n3389) );
  NOR U3771 ( .A(n3734), .B(n3388), .Z(n3736) );
  AND U3772 ( .A(n3484), .B(n3483), .Z(n3388) );
  IV U3773 ( .A(n3696), .Z(n3483) );
  XOR U3774 ( .A(n3741), .B(n3742), .Z(n3734) );
  AND U3775 ( .A(n3743), .B(n3744), .Z(n3742) );
  XNOR U3776 ( .A(n3741), .B(n3445), .Z(n3744) );
  XOR U3777 ( .A(n3502), .B(n3745), .Z(n3445) );
  AND U3778 ( .A(n184), .B(n3746), .Z(n3745) );
  XOR U3779 ( .A(n3498), .B(n3502), .Z(n3746) );
  XNOR U3780 ( .A(n3747), .B(n3741), .Z(n3743) );
  IV U3781 ( .A(n3397), .Z(n3747) );
  XOR U3782 ( .A(n3748), .B(n3749), .Z(n3397) );
  AND U3783 ( .A(n200), .B(n3750), .Z(n3749) );
  XOR U3784 ( .A(n3751), .B(n3752), .Z(n3741) );
  AND U3785 ( .A(n3753), .B(n3754), .Z(n3752) );
  XNOR U3786 ( .A(n3751), .B(n3455), .Z(n3754) );
  XOR U3787 ( .A(n3530), .B(n3755), .Z(n3455) );
  AND U3788 ( .A(n184), .B(n3756), .Z(n3755) );
  XOR U3789 ( .A(n3526), .B(n3530), .Z(n3756) );
  XOR U3790 ( .A(n3406), .B(n3751), .Z(n3753) );
  XOR U3791 ( .A(n3757), .B(n3758), .Z(n3406) );
  AND U3792 ( .A(n200), .B(n3759), .Z(n3758) );
  XOR U3793 ( .A(n3728), .B(n3760), .Z(n3751) );
  AND U3794 ( .A(n3761), .B(n3731), .Z(n3760) );
  XNOR U3795 ( .A(n3465), .B(n3728), .Z(n3731) );
  XOR U3796 ( .A(n3579), .B(n3762), .Z(n3465) );
  AND U3797 ( .A(n184), .B(n3763), .Z(n3762) );
  XOR U3798 ( .A(n3575), .B(n3579), .Z(n3763) );
  XNOR U3799 ( .A(n3764), .B(n3728), .Z(n3761) );
  IV U3800 ( .A(n3414), .Z(n3764) );
  XOR U3801 ( .A(n3765), .B(n3766), .Z(n3414) );
  AND U3802 ( .A(n200), .B(n3767), .Z(n3766) );
  XOR U3803 ( .A(n3768), .B(n3769), .Z(n3728) );
  AND U3804 ( .A(n3770), .B(n3771), .Z(n3769) );
  XNOR U3805 ( .A(n3768), .B(n3473), .Z(n3771) );
  XOR U3806 ( .A(n3672), .B(n3772), .Z(n3473) );
  AND U3807 ( .A(n184), .B(n3773), .Z(n3772) );
  XOR U3808 ( .A(n3668), .B(n3672), .Z(n3773) );
  XNOR U3809 ( .A(n3774), .B(n3768), .Z(n3770) );
  IV U3810 ( .A(n3424), .Z(n3774) );
  XOR U3811 ( .A(n3775), .B(n3776), .Z(n3424) );
  AND U3812 ( .A(n200), .B(n3777), .Z(n3776) );
  AND U3813 ( .A(n3732), .B(n3713), .Z(n3768) );
  XNOR U3814 ( .A(n3778), .B(n3779), .Z(n3713) );
  AND U3815 ( .A(n184), .B(n3691), .Z(n3779) );
  XNOR U3816 ( .A(n3689), .B(n3778), .Z(n3691) );
  XNOR U3817 ( .A(n3780), .B(n3781), .Z(n184) );
  NOR U3818 ( .A(n3782), .B(n3783), .Z(n3781) );
  XNOR U3819 ( .A(n3780), .B(n3696), .Z(n3783) );
  NOR U3820 ( .A(n3739), .B(n3740), .Z(n3696) );
  NOR U3821 ( .A(n3780), .B(n3484), .Z(n3782) );
  AND U3822 ( .A(n3784), .B(n3785), .Z(n3484) );
  IV U3823 ( .A(n3786), .Z(n3784) );
  XOR U3824 ( .A(n3787), .B(n3788), .Z(n3780) );
  AND U3825 ( .A(n3789), .B(n3790), .Z(n3788) );
  XNOR U3826 ( .A(n3787), .B(n3498), .Z(n3790) );
  IV U3827 ( .A(n3501), .Z(n3498) );
  XOR U3828 ( .A(n3791), .B(n3792), .Z(n3501) );
  AND U3829 ( .A(n188), .B(n3793), .Z(n3792) );
  XOR U3830 ( .A(n3794), .B(n3791), .Z(n3793) );
  XOR U3831 ( .A(n3502), .B(n3787), .Z(n3789) );
  XOR U3832 ( .A(n3795), .B(n3796), .Z(n3502) );
  AND U3833 ( .A(n196), .B(n3750), .Z(n3796) );
  XOR U3834 ( .A(n3795), .B(n3748), .Z(n3750) );
  XOR U3835 ( .A(n3797), .B(n3798), .Z(n3787) );
  AND U3836 ( .A(n3799), .B(n3800), .Z(n3798) );
  XNOR U3837 ( .A(n3797), .B(n3526), .Z(n3800) );
  IV U3838 ( .A(n3529), .Z(n3526) );
  XOR U3839 ( .A(n3801), .B(n3802), .Z(n3529) );
  AND U3840 ( .A(n188), .B(n3803), .Z(n3802) );
  XNOR U3841 ( .A(n3804), .B(n3801), .Z(n3803) );
  XOR U3842 ( .A(n3530), .B(n3797), .Z(n3799) );
  XOR U3843 ( .A(n3805), .B(n3806), .Z(n3530) );
  AND U3844 ( .A(n196), .B(n3759), .Z(n3806) );
  XOR U3845 ( .A(n3805), .B(n3757), .Z(n3759) );
  XOR U3846 ( .A(n3807), .B(n3808), .Z(n3797) );
  AND U3847 ( .A(n3809), .B(n3810), .Z(n3808) );
  XNOR U3848 ( .A(n3807), .B(n3575), .Z(n3810) );
  IV U3849 ( .A(n3578), .Z(n3575) );
  XOR U3850 ( .A(n3811), .B(n3812), .Z(n3578) );
  AND U3851 ( .A(n188), .B(n3813), .Z(n3812) );
  XOR U3852 ( .A(n3814), .B(n3811), .Z(n3813) );
  XOR U3853 ( .A(n3579), .B(n3807), .Z(n3809) );
  XOR U3854 ( .A(n3815), .B(n3816), .Z(n3579) );
  AND U3855 ( .A(n196), .B(n3767), .Z(n3816) );
  XOR U3856 ( .A(n3815), .B(n3765), .Z(n3767) );
  XOR U3857 ( .A(n3709), .B(n3817), .Z(n3807) );
  AND U3858 ( .A(n3711), .B(n3818), .Z(n3817) );
  XNOR U3859 ( .A(n3709), .B(n3668), .Z(n3818) );
  IV U3860 ( .A(n3671), .Z(n3668) );
  XOR U3861 ( .A(n3819), .B(n3820), .Z(n3671) );
  AND U3862 ( .A(n188), .B(n3821), .Z(n3820) );
  XNOR U3863 ( .A(n3822), .B(n3819), .Z(n3821) );
  XOR U3864 ( .A(n3672), .B(n3709), .Z(n3711) );
  XOR U3865 ( .A(n3823), .B(n3824), .Z(n3672) );
  AND U3866 ( .A(n196), .B(n3777), .Z(n3824) );
  XOR U3867 ( .A(n3823), .B(n3775), .Z(n3777) );
  AND U3868 ( .A(n3778), .B(n3689), .Z(n3709) );
  XNOR U3869 ( .A(n3825), .B(n3826), .Z(n3689) );
  AND U3870 ( .A(n188), .B(n3827), .Z(n3826) );
  XNOR U3871 ( .A(n3828), .B(n3825), .Z(n3827) );
  XNOR U3872 ( .A(n3829), .B(n3830), .Z(n188) );
  NOR U3873 ( .A(n3831), .B(n3832), .Z(n3830) );
  XNOR U3874 ( .A(n3829), .B(n3786), .Z(n3832) );
  NOR U3875 ( .A(n3833), .B(n3834), .Z(n3786) );
  NOR U3876 ( .A(n3829), .B(n3785), .Z(n3831) );
  AND U3877 ( .A(n3835), .B(n3836), .Z(n3785) );
  XOR U3878 ( .A(n3837), .B(n3838), .Z(n3829) );
  AND U3879 ( .A(n3839), .B(n3840), .Z(n3838) );
  XNOR U3880 ( .A(n3837), .B(n3835), .Z(n3840) );
  IV U3881 ( .A(n3794), .Z(n3835) );
  XOR U3882 ( .A(n3841), .B(n3842), .Z(n3794) );
  XOR U3883 ( .A(n3843), .B(n3836), .Z(n3842) );
  AND U3884 ( .A(n3804), .B(n3844), .Z(n3836) );
  AND U3885 ( .A(n3845), .B(n3846), .Z(n3843) );
  XOR U3886 ( .A(n3847), .B(n3841), .Z(n3845) );
  XNOR U3887 ( .A(n3791), .B(n3837), .Z(n3839) );
  XNOR U3888 ( .A(n3848), .B(n3849), .Z(n3791) );
  AND U3889 ( .A(n192), .B(n3850), .Z(n3849) );
  XNOR U3890 ( .A(n3851), .B(n3852), .Z(n3850) );
  XOR U3891 ( .A(n3853), .B(n3854), .Z(n3837) );
  AND U3892 ( .A(n3855), .B(n3856), .Z(n3854) );
  XNOR U3893 ( .A(n3853), .B(n3804), .Z(n3856) );
  XOR U3894 ( .A(n3857), .B(n3846), .Z(n3804) );
  XNOR U3895 ( .A(n3858), .B(n3841), .Z(n3846) );
  XOR U3896 ( .A(n3859), .B(n3860), .Z(n3841) );
  AND U3897 ( .A(n3861), .B(n3862), .Z(n3860) );
  XOR U3898 ( .A(n3863), .B(n3859), .Z(n3861) );
  XNOR U3899 ( .A(n3864), .B(n3865), .Z(n3858) );
  AND U3900 ( .A(n3866), .B(n3867), .Z(n3865) );
  XOR U3901 ( .A(n3864), .B(n3868), .Z(n3866) );
  XNOR U3902 ( .A(n3847), .B(n3844), .Z(n3857) );
  AND U3903 ( .A(n3869), .B(n3870), .Z(n3844) );
  XOR U3904 ( .A(n3871), .B(n3872), .Z(n3847) );
  AND U3905 ( .A(n3873), .B(n3874), .Z(n3872) );
  XOR U3906 ( .A(n3871), .B(n3875), .Z(n3873) );
  XNOR U3907 ( .A(n3801), .B(n3853), .Z(n3855) );
  XNOR U3908 ( .A(n3876), .B(n3877), .Z(n3801) );
  AND U3909 ( .A(n192), .B(n3878), .Z(n3877) );
  XNOR U3910 ( .A(n3879), .B(n3880), .Z(n3878) );
  XOR U3911 ( .A(n3881), .B(n3882), .Z(n3853) );
  AND U3912 ( .A(n3883), .B(n3884), .Z(n3882) );
  XNOR U3913 ( .A(n3881), .B(n3869), .Z(n3884) );
  IV U3914 ( .A(n3814), .Z(n3869) );
  XNOR U3915 ( .A(n3885), .B(n3862), .Z(n3814) );
  XNOR U3916 ( .A(n3886), .B(n3868), .Z(n3862) );
  XOR U3917 ( .A(n3887), .B(n3888), .Z(n3868) );
  AND U3918 ( .A(n3889), .B(n3890), .Z(n3888) );
  XOR U3919 ( .A(n3887), .B(n3891), .Z(n3889) );
  XNOR U3920 ( .A(n3867), .B(n3859), .Z(n3886) );
  XOR U3921 ( .A(n3892), .B(n3893), .Z(n3859) );
  AND U3922 ( .A(n3894), .B(n3895), .Z(n3893) );
  XNOR U3923 ( .A(n3896), .B(n3892), .Z(n3894) );
  XNOR U3924 ( .A(n3897), .B(n3864), .Z(n3867) );
  XOR U3925 ( .A(n3898), .B(n3899), .Z(n3864) );
  AND U3926 ( .A(n3900), .B(n3901), .Z(n3899) );
  XOR U3927 ( .A(n3898), .B(n3902), .Z(n3900) );
  XNOR U3928 ( .A(n3903), .B(n3904), .Z(n3897) );
  AND U3929 ( .A(n3905), .B(n3906), .Z(n3904) );
  XNOR U3930 ( .A(n3903), .B(n3907), .Z(n3905) );
  XNOR U3931 ( .A(n3863), .B(n3870), .Z(n3885) );
  AND U3932 ( .A(n3822), .B(n3908), .Z(n3870) );
  XOR U3933 ( .A(n3875), .B(n3874), .Z(n3863) );
  XNOR U3934 ( .A(n3909), .B(n3871), .Z(n3874) );
  XOR U3935 ( .A(n3910), .B(n3911), .Z(n3871) );
  AND U3936 ( .A(n3912), .B(n3913), .Z(n3911) );
  XOR U3937 ( .A(n3910), .B(n3914), .Z(n3912) );
  XNOR U3938 ( .A(n3915), .B(n3916), .Z(n3909) );
  AND U3939 ( .A(n3917), .B(n3918), .Z(n3916) );
  XOR U3940 ( .A(n3915), .B(n3919), .Z(n3917) );
  XOR U3941 ( .A(n3920), .B(n3921), .Z(n3875) );
  AND U3942 ( .A(n3922), .B(n3923), .Z(n3921) );
  XOR U3943 ( .A(n3920), .B(n3924), .Z(n3922) );
  XNOR U3944 ( .A(n3811), .B(n3881), .Z(n3883) );
  XNOR U3945 ( .A(n3925), .B(n3926), .Z(n3811) );
  AND U3946 ( .A(n192), .B(n3927), .Z(n3926) );
  XNOR U3947 ( .A(n3928), .B(n3929), .Z(n3927) );
  XOR U3948 ( .A(n3930), .B(n3931), .Z(n3881) );
  AND U3949 ( .A(n3932), .B(n3933), .Z(n3931) );
  XNOR U3950 ( .A(n3930), .B(n3822), .Z(n3933) );
  XOR U3951 ( .A(n3934), .B(n3895), .Z(n3822) );
  XNOR U3952 ( .A(n3935), .B(n3902), .Z(n3895) );
  XOR U3953 ( .A(n3891), .B(n3890), .Z(n3902) );
  XNOR U3954 ( .A(n3936), .B(n3887), .Z(n3890) );
  XOR U3955 ( .A(n3937), .B(n3938), .Z(n3887) );
  AND U3956 ( .A(n3939), .B(n3940), .Z(n3938) );
  XNOR U3957 ( .A(n3941), .B(n3942), .Z(n3939) );
  IV U3958 ( .A(n3937), .Z(n3941) );
  XNOR U3959 ( .A(n3943), .B(n3944), .Z(n3936) );
  NOR U3960 ( .A(n3945), .B(n3946), .Z(n3944) );
  XNOR U3961 ( .A(n3943), .B(n3947), .Z(n3945) );
  XOR U3962 ( .A(n3948), .B(n3949), .Z(n3891) );
  NOR U3963 ( .A(n3950), .B(n3951), .Z(n3949) );
  XNOR U3964 ( .A(n3948), .B(n3952), .Z(n3950) );
  XNOR U3965 ( .A(n3901), .B(n3892), .Z(n3935) );
  XOR U3966 ( .A(n3953), .B(n3954), .Z(n3892) );
  AND U3967 ( .A(n3955), .B(n3956), .Z(n3954) );
  XOR U3968 ( .A(n3953), .B(n3957), .Z(n3955) );
  XOR U3969 ( .A(n3958), .B(n3907), .Z(n3901) );
  XOR U3970 ( .A(n3959), .B(n3960), .Z(n3907) );
  NOR U3971 ( .A(n3961), .B(n3962), .Z(n3960) );
  XOR U3972 ( .A(n3959), .B(n3963), .Z(n3961) );
  XNOR U3973 ( .A(n3906), .B(n3898), .Z(n3958) );
  XOR U3974 ( .A(n3964), .B(n3965), .Z(n3898) );
  AND U3975 ( .A(n3966), .B(n3967), .Z(n3965) );
  XOR U3976 ( .A(n3964), .B(n3968), .Z(n3966) );
  XNOR U3977 ( .A(n3969), .B(n3903), .Z(n3906) );
  XNOR U3978 ( .A(n3970), .B(n3971), .Z(n3903) );
  NOR U3979 ( .A(n3972), .B(n3973), .Z(n3971) );
  XOR U3980 ( .A(n3970), .B(n3974), .Z(n3972) );
  XNOR U3981 ( .A(n3975), .B(n3976), .Z(n3969) );
  NOR U3982 ( .A(n3977), .B(n3978), .Z(n3976) );
  XNOR U3983 ( .A(n3975), .B(n3979), .Z(n3977) );
  XOR U3984 ( .A(n3896), .B(n3908), .Z(n3934) );
  NOR U3985 ( .A(n3828), .B(n3980), .Z(n3908) );
  XNOR U3986 ( .A(n3914), .B(n3913), .Z(n3896) );
  XNOR U3987 ( .A(n3981), .B(n3919), .Z(n3913) );
  XNOR U3988 ( .A(n3982), .B(n3983), .Z(n3919) );
  NOR U3989 ( .A(n3984), .B(n3985), .Z(n3983) );
  XOR U3990 ( .A(n3982), .B(n3986), .Z(n3984) );
  XNOR U3991 ( .A(n3918), .B(n3910), .Z(n3981) );
  XOR U3992 ( .A(n3987), .B(n3988), .Z(n3910) );
  AND U3993 ( .A(n3989), .B(n3990), .Z(n3988) );
  XOR U3994 ( .A(n3987), .B(n3991), .Z(n3989) );
  XNOR U3995 ( .A(n3992), .B(n3915), .Z(n3918) );
  XOR U3996 ( .A(n3993), .B(n3994), .Z(n3915) );
  AND U3997 ( .A(n3995), .B(n3996), .Z(n3994) );
  XNOR U3998 ( .A(n3997), .B(n3998), .Z(n3995) );
  IV U3999 ( .A(n3993), .Z(n3997) );
  XNOR U4000 ( .A(n3999), .B(n4000), .Z(n3992) );
  NOR U4001 ( .A(n4001), .B(n4002), .Z(n4000) );
  XNOR U4002 ( .A(n3999), .B(n4003), .Z(n4001) );
  XOR U4003 ( .A(n3924), .B(n3923), .Z(n3914) );
  XNOR U4004 ( .A(n4004), .B(n3920), .Z(n3923) );
  XOR U4005 ( .A(n4005), .B(n4006), .Z(n3920) );
  NOR U4006 ( .A(n4007), .B(n4008), .Z(n4006) );
  XNOR U4007 ( .A(n4005), .B(n4009), .Z(n4007) );
  XNOR U4008 ( .A(n4010), .B(n4011), .Z(n4004) );
  NOR U4009 ( .A(n4012), .B(n4013), .Z(n4011) );
  XNOR U4010 ( .A(n4010), .B(n4014), .Z(n4012) );
  XOR U4011 ( .A(n4015), .B(n4016), .Z(n3924) );
  NOR U4012 ( .A(n4017), .B(n4018), .Z(n4016) );
  XNOR U4013 ( .A(n4015), .B(n4019), .Z(n4017) );
  XNOR U4014 ( .A(n3819), .B(n3930), .Z(n3932) );
  XNOR U4015 ( .A(n4020), .B(n4021), .Z(n3819) );
  AND U4016 ( .A(n192), .B(n4022), .Z(n4021) );
  XNOR U4017 ( .A(n4023), .B(n4024), .Z(n4022) );
  AND U4018 ( .A(n3825), .B(n3828), .Z(n3930) );
  XOR U4019 ( .A(n4025), .B(n3980), .Z(n3828) );
  XNOR U4020 ( .A(p_input[256]), .B(p_input[96]), .Z(n3980) );
  XNOR U4021 ( .A(n3957), .B(n3956), .Z(n4025) );
  XNOR U4022 ( .A(n4026), .B(n3968), .Z(n3956) );
  XOR U4023 ( .A(n3942), .B(n3940), .Z(n3968) );
  XNOR U4024 ( .A(n4027), .B(n3947), .Z(n3940) );
  XOR U4025 ( .A(p_input[120]), .B(p_input[280]), .Z(n3947) );
  XOR U4026 ( .A(n3937), .B(n3946), .Z(n4027) );
  XOR U4027 ( .A(n4028), .B(n3943), .Z(n3946) );
  XOR U4028 ( .A(p_input[118]), .B(p_input[278]), .Z(n3943) );
  XOR U4029 ( .A(p_input[119]), .B(n2951), .Z(n4028) );
  XOR U4030 ( .A(p_input[114]), .B(p_input[274]), .Z(n3937) );
  XNOR U4031 ( .A(n3952), .B(n3951), .Z(n3942) );
  XOR U4032 ( .A(n4029), .B(n3948), .Z(n3951) );
  XOR U4033 ( .A(p_input[115]), .B(p_input[275]), .Z(n3948) );
  XOR U4034 ( .A(p_input[116]), .B(n2953), .Z(n4029) );
  XOR U4035 ( .A(p_input[117]), .B(p_input[277]), .Z(n3952) );
  XNOR U4036 ( .A(n3967), .B(n3953), .Z(n4026) );
  XNOR U4037 ( .A(n3318), .B(p_input[97]), .Z(n3953) );
  XNOR U4038 ( .A(n4030), .B(n3974), .Z(n3967) );
  XNOR U4039 ( .A(n3963), .B(n3962), .Z(n3974) );
  XNOR U4040 ( .A(n4031), .B(n3959), .Z(n3962) );
  XNOR U4041 ( .A(p_input[122]), .B(p_input[282]), .Z(n3959) );
  XOR U4042 ( .A(p_input[123]), .B(n2957), .Z(n4031) );
  XOR U4043 ( .A(p_input[124]), .B(p_input[284]), .Z(n3963) );
  XNOR U4044 ( .A(n3973), .B(n4032), .Z(n4030) );
  IV U4045 ( .A(n3964), .Z(n4032) );
  XOR U4046 ( .A(p_input[113]), .B(p_input[273]), .Z(n3964) );
  XOR U4047 ( .A(n4033), .B(n3979), .Z(n3973) );
  XOR U4048 ( .A(p_input[127]), .B(p_input[287]), .Z(n3979) );
  XNOR U4049 ( .A(n3970), .B(n3978), .Z(n4033) );
  XOR U4050 ( .A(n4034), .B(n3975), .Z(n3978) );
  XOR U4051 ( .A(p_input[125]), .B(p_input[285]), .Z(n3975) );
  XNOR U4052 ( .A(p_input[126]), .B(p_input[286]), .Z(n4034) );
  XNOR U4053 ( .A(p_input[121]), .B(p_input[281]), .Z(n3970) );
  XOR U4054 ( .A(n3991), .B(n3990), .Z(n3957) );
  XNOR U4055 ( .A(n4035), .B(n3998), .Z(n3990) );
  XNOR U4056 ( .A(n3986), .B(n3985), .Z(n3998) );
  XNOR U4057 ( .A(n4036), .B(n3982), .Z(n3985) );
  XNOR U4058 ( .A(p_input[107]), .B(p_input[267]), .Z(n3982) );
  XOR U4059 ( .A(p_input[108]), .B(n2963), .Z(n4036) );
  XOR U4060 ( .A(p_input[109]), .B(p_input[269]), .Z(n3986) );
  XNOR U4061 ( .A(n3996), .B(n3987), .Z(n4035) );
  XOR U4062 ( .A(p_input[258]), .B(p_input[98]), .Z(n3987) );
  XNOR U4063 ( .A(n4037), .B(n4003), .Z(n3996) );
  XNOR U4064 ( .A(p_input[112]), .B(n2965), .Z(n4003) );
  XOR U4065 ( .A(n3993), .B(n4002), .Z(n4037) );
  XOR U4066 ( .A(n4038), .B(n3999), .Z(n4002) );
  XOR U4067 ( .A(p_input[110]), .B(p_input[270]), .Z(n3999) );
  XOR U4068 ( .A(p_input[111]), .B(n2967), .Z(n4038) );
  XOR U4069 ( .A(p_input[106]), .B(p_input[266]), .Z(n3993) );
  XNOR U4070 ( .A(n4009), .B(n4008), .Z(n3991) );
  XOR U4071 ( .A(n4039), .B(n4014), .Z(n4008) );
  XOR U4072 ( .A(p_input[105]), .B(p_input[265]), .Z(n4014) );
  XOR U4073 ( .A(n4005), .B(n4013), .Z(n4039) );
  XOR U4074 ( .A(n4040), .B(n4010), .Z(n4013) );
  XOR U4075 ( .A(p_input[103]), .B(p_input[263]), .Z(n4010) );
  XNOR U4076 ( .A(p_input[104]), .B(p_input[264]), .Z(n4040) );
  XOR U4077 ( .A(p_input[259]), .B(p_input[99]), .Z(n4005) );
  XNOR U4078 ( .A(n4019), .B(n4018), .Z(n4009) );
  XOR U4079 ( .A(n4041), .B(n4015), .Z(n4018) );
  XOR U4080 ( .A(p_input[100]), .B(p_input[260]), .Z(n4015) );
  XNOR U4081 ( .A(p_input[101]), .B(p_input[261]), .Z(n4041) );
  XOR U4082 ( .A(p_input[102]), .B(p_input[262]), .Z(n4019) );
  XNOR U4083 ( .A(n4042), .B(n4043), .Z(n3825) );
  AND U4084 ( .A(n192), .B(n4044), .Z(n4043) );
  XNOR U4085 ( .A(n4045), .B(n4046), .Z(n192) );
  NOR U4086 ( .A(n4047), .B(n4048), .Z(n4046) );
  XNOR U4087 ( .A(n4045), .B(n4049), .Z(n4048) );
  NOR U4088 ( .A(n4045), .B(n3834), .Z(n4047) );
  XOR U4089 ( .A(n4050), .B(n4051), .Z(n4045) );
  AND U4090 ( .A(n4052), .B(n4053), .Z(n4051) );
  XOR U4091 ( .A(n3851), .B(n4050), .Z(n4053) );
  XOR U4092 ( .A(n4050), .B(n3852), .Z(n4052) );
  XOR U4093 ( .A(n4054), .B(n4055), .Z(n4050) );
  AND U4094 ( .A(n4056), .B(n4057), .Z(n4055) );
  XOR U4095 ( .A(n3879), .B(n4054), .Z(n4057) );
  XOR U4096 ( .A(n4054), .B(n3880), .Z(n4056) );
  XOR U4097 ( .A(n4058), .B(n4059), .Z(n4054) );
  AND U4098 ( .A(n4060), .B(n4061), .Z(n4059) );
  XOR U4099 ( .A(n3928), .B(n4058), .Z(n4061) );
  XOR U4100 ( .A(n4058), .B(n3929), .Z(n4060) );
  XOR U4101 ( .A(n4062), .B(n4063), .Z(n4058) );
  AND U4102 ( .A(n4064), .B(n4065), .Z(n4063) );
  XOR U4103 ( .A(n4062), .B(n4023), .Z(n4065) );
  XNOR U4104 ( .A(n4066), .B(n4067), .Z(n3778) );
  AND U4105 ( .A(n196), .B(n4068), .Z(n4067) );
  XNOR U4106 ( .A(n4069), .B(n4070), .Z(n196) );
  NOR U4107 ( .A(n4071), .B(n4072), .Z(n4070) );
  XOR U4108 ( .A(n3740), .B(n4069), .Z(n4072) );
  NOR U4109 ( .A(n4069), .B(n3739), .Z(n4071) );
  XOR U4110 ( .A(n4073), .B(n4074), .Z(n4069) );
  AND U4111 ( .A(n4075), .B(n4076), .Z(n4074) );
  XNOR U4112 ( .A(n3795), .B(n4073), .Z(n4076) );
  XOR U4113 ( .A(n4073), .B(n3748), .Z(n4075) );
  XOR U4114 ( .A(n4077), .B(n4078), .Z(n4073) );
  AND U4115 ( .A(n4079), .B(n4080), .Z(n4078) );
  XNOR U4116 ( .A(n3805), .B(n4077), .Z(n4080) );
  XOR U4117 ( .A(n4077), .B(n3757), .Z(n4079) );
  XOR U4118 ( .A(n4081), .B(n4082), .Z(n4077) );
  AND U4119 ( .A(n4083), .B(n4084), .Z(n4082) );
  XOR U4120 ( .A(n4081), .B(n3765), .Z(n4083) );
  XOR U4121 ( .A(n4085), .B(n4086), .Z(n3732) );
  AND U4122 ( .A(n200), .B(n4068), .Z(n4086) );
  XNOR U4123 ( .A(n4066), .B(n4085), .Z(n4068) );
  XNOR U4124 ( .A(n4087), .B(n4088), .Z(n200) );
  NOR U4125 ( .A(n4089), .B(n4090), .Z(n4088) );
  XNOR U4126 ( .A(n3740), .B(n4091), .Z(n4090) );
  IV U4127 ( .A(n4087), .Z(n4091) );
  AND U4128 ( .A(n4092), .B(n4093), .Z(n3740) );
  NOR U4129 ( .A(n4087), .B(n3739), .Z(n4089) );
  AND U4130 ( .A(n3834), .B(n3833), .Z(n3739) );
  IV U4131 ( .A(n4049), .Z(n3833) );
  XOR U4132 ( .A(n4094), .B(n4095), .Z(n4087) );
  AND U4133 ( .A(n4096), .B(n4097), .Z(n4095) );
  XNOR U4134 ( .A(n4094), .B(n3795), .Z(n4097) );
  XOR U4135 ( .A(n3852), .B(n4098), .Z(n3795) );
  AND U4136 ( .A(n203), .B(n4099), .Z(n4098) );
  XOR U4137 ( .A(n3848), .B(n3852), .Z(n4099) );
  XNOR U4138 ( .A(n4100), .B(n4094), .Z(n4096) );
  IV U4139 ( .A(n3748), .Z(n4100) );
  XOR U4140 ( .A(n4101), .B(n4102), .Z(n3748) );
  AND U4141 ( .A(n218), .B(n4103), .Z(n4102) );
  XOR U4142 ( .A(n4104), .B(n4105), .Z(n4094) );
  AND U4143 ( .A(n4106), .B(n4107), .Z(n4105) );
  XNOR U4144 ( .A(n4104), .B(n3805), .Z(n4107) );
  XOR U4145 ( .A(n3880), .B(n4108), .Z(n3805) );
  AND U4146 ( .A(n203), .B(n4109), .Z(n4108) );
  XOR U4147 ( .A(n3876), .B(n3880), .Z(n4109) );
  XOR U4148 ( .A(n3757), .B(n4104), .Z(n4106) );
  XOR U4149 ( .A(n4110), .B(n4111), .Z(n3757) );
  AND U4150 ( .A(n218), .B(n4112), .Z(n4111) );
  XOR U4151 ( .A(n4081), .B(n4113), .Z(n4104) );
  AND U4152 ( .A(n4114), .B(n4084), .Z(n4113) );
  XNOR U4153 ( .A(n3815), .B(n4081), .Z(n4084) );
  XOR U4154 ( .A(n3929), .B(n4115), .Z(n3815) );
  AND U4155 ( .A(n203), .B(n4116), .Z(n4115) );
  XOR U4156 ( .A(n3925), .B(n3929), .Z(n4116) );
  XNOR U4157 ( .A(n4117), .B(n4081), .Z(n4114) );
  IV U4158 ( .A(n3765), .Z(n4117) );
  XOR U4159 ( .A(n4118), .B(n4119), .Z(n3765) );
  AND U4160 ( .A(n218), .B(n4120), .Z(n4119) );
  XOR U4161 ( .A(n4121), .B(n4122), .Z(n4081) );
  AND U4162 ( .A(n4123), .B(n4124), .Z(n4122) );
  XNOR U4163 ( .A(n4121), .B(n3823), .Z(n4124) );
  XOR U4164 ( .A(n4024), .B(n4125), .Z(n3823) );
  AND U4165 ( .A(n203), .B(n4126), .Z(n4125) );
  XOR U4166 ( .A(n4020), .B(n4024), .Z(n4126) );
  XNOR U4167 ( .A(n4127), .B(n4121), .Z(n4123) );
  IV U4168 ( .A(n3775), .Z(n4127) );
  XOR U4169 ( .A(n4128), .B(n4129), .Z(n3775) );
  AND U4170 ( .A(n218), .B(n4130), .Z(n4129) );
  AND U4171 ( .A(n4085), .B(n4066), .Z(n4121) );
  XNOR U4172 ( .A(n4131), .B(n4132), .Z(n4066) );
  AND U4173 ( .A(n203), .B(n4044), .Z(n4132) );
  XNOR U4174 ( .A(n4042), .B(n4131), .Z(n4044) );
  XNOR U4175 ( .A(n4133), .B(n4134), .Z(n203) );
  NOR U4176 ( .A(n4135), .B(n4136), .Z(n4134) );
  XNOR U4177 ( .A(n4133), .B(n4049), .Z(n4136) );
  NOR U4178 ( .A(n4092), .B(n4093), .Z(n4049) );
  NOR U4179 ( .A(n4133), .B(n3834), .Z(n4135) );
  AND U4180 ( .A(n4137), .B(n4138), .Z(n3834) );
  IV U4181 ( .A(n4139), .Z(n4137) );
  XOR U4182 ( .A(n4140), .B(n4141), .Z(n4133) );
  AND U4183 ( .A(n4142), .B(n4143), .Z(n4141) );
  XNOR U4184 ( .A(n4140), .B(n3848), .Z(n4143) );
  IV U4185 ( .A(n3851), .Z(n3848) );
  XOR U4186 ( .A(n4144), .B(n4145), .Z(n3851) );
  AND U4187 ( .A(n207), .B(n4146), .Z(n4145) );
  XOR U4188 ( .A(n4147), .B(n4144), .Z(n4146) );
  XOR U4189 ( .A(n3852), .B(n4140), .Z(n4142) );
  XOR U4190 ( .A(n4148), .B(n4149), .Z(n3852) );
  AND U4191 ( .A(n214), .B(n4103), .Z(n4149) );
  XOR U4192 ( .A(n4148), .B(n4101), .Z(n4103) );
  XOR U4193 ( .A(n4150), .B(n4151), .Z(n4140) );
  AND U4194 ( .A(n4152), .B(n4153), .Z(n4151) );
  XNOR U4195 ( .A(n4150), .B(n3876), .Z(n4153) );
  IV U4196 ( .A(n3879), .Z(n3876) );
  XOR U4197 ( .A(n4154), .B(n4155), .Z(n3879) );
  AND U4198 ( .A(n207), .B(n4156), .Z(n4155) );
  XNOR U4199 ( .A(n4157), .B(n4154), .Z(n4156) );
  XOR U4200 ( .A(n3880), .B(n4150), .Z(n4152) );
  XOR U4201 ( .A(n4158), .B(n4159), .Z(n3880) );
  AND U4202 ( .A(n214), .B(n4112), .Z(n4159) );
  XOR U4203 ( .A(n4158), .B(n4110), .Z(n4112) );
  XOR U4204 ( .A(n4160), .B(n4161), .Z(n4150) );
  AND U4205 ( .A(n4162), .B(n4163), .Z(n4161) );
  XNOR U4206 ( .A(n4160), .B(n3925), .Z(n4163) );
  IV U4207 ( .A(n3928), .Z(n3925) );
  XOR U4208 ( .A(n4164), .B(n4165), .Z(n3928) );
  AND U4209 ( .A(n207), .B(n4166), .Z(n4165) );
  XOR U4210 ( .A(n4167), .B(n4164), .Z(n4166) );
  XOR U4211 ( .A(n3929), .B(n4160), .Z(n4162) );
  XOR U4212 ( .A(n4168), .B(n4169), .Z(n3929) );
  AND U4213 ( .A(n214), .B(n4120), .Z(n4169) );
  XOR U4214 ( .A(n4168), .B(n4118), .Z(n4120) );
  XOR U4215 ( .A(n4062), .B(n4170), .Z(n4160) );
  AND U4216 ( .A(n4064), .B(n4171), .Z(n4170) );
  XNOR U4217 ( .A(n4062), .B(n4020), .Z(n4171) );
  IV U4218 ( .A(n4023), .Z(n4020) );
  XOR U4219 ( .A(n4172), .B(n4173), .Z(n4023) );
  AND U4220 ( .A(n207), .B(n4174), .Z(n4173) );
  XNOR U4221 ( .A(n4175), .B(n4172), .Z(n4174) );
  XOR U4222 ( .A(n4024), .B(n4062), .Z(n4064) );
  XOR U4223 ( .A(n4176), .B(n4177), .Z(n4024) );
  AND U4224 ( .A(n214), .B(n4130), .Z(n4177) );
  XOR U4225 ( .A(n4176), .B(n4128), .Z(n4130) );
  AND U4226 ( .A(n4131), .B(n4042), .Z(n4062) );
  XNOR U4227 ( .A(n4178), .B(n4179), .Z(n4042) );
  AND U4228 ( .A(n207), .B(n4180), .Z(n4179) );
  XNOR U4229 ( .A(n4181), .B(n4178), .Z(n4180) );
  XNOR U4230 ( .A(n4182), .B(n4183), .Z(n207) );
  NOR U4231 ( .A(n4184), .B(n4185), .Z(n4183) );
  XNOR U4232 ( .A(n4182), .B(n4139), .Z(n4185) );
  NOR U4233 ( .A(n4186), .B(n4187), .Z(n4139) );
  NOR U4234 ( .A(n4182), .B(n4138), .Z(n4184) );
  AND U4235 ( .A(n4188), .B(n4189), .Z(n4138) );
  XOR U4236 ( .A(n4190), .B(n4191), .Z(n4182) );
  AND U4237 ( .A(n4192), .B(n4193), .Z(n4191) );
  XNOR U4238 ( .A(n4190), .B(n4188), .Z(n4193) );
  IV U4239 ( .A(n4147), .Z(n4188) );
  XOR U4240 ( .A(n4194), .B(n4195), .Z(n4147) );
  XOR U4241 ( .A(n4196), .B(n4189), .Z(n4195) );
  AND U4242 ( .A(n4157), .B(n4197), .Z(n4189) );
  AND U4243 ( .A(n4198), .B(n4199), .Z(n4196) );
  XOR U4244 ( .A(n4200), .B(n4194), .Z(n4198) );
  XNOR U4245 ( .A(n4144), .B(n4190), .Z(n4192) );
  XNOR U4246 ( .A(n4201), .B(n4202), .Z(n4144) );
  AND U4247 ( .A(n210), .B(n4203), .Z(n4202) );
  XOR U4248 ( .A(n4204), .B(n4205), .Z(n4190) );
  AND U4249 ( .A(n4206), .B(n4207), .Z(n4205) );
  XNOR U4250 ( .A(n4204), .B(n4157), .Z(n4207) );
  XOR U4251 ( .A(n4208), .B(n4199), .Z(n4157) );
  XNOR U4252 ( .A(n4209), .B(n4194), .Z(n4199) );
  XOR U4253 ( .A(n4210), .B(n4211), .Z(n4194) );
  AND U4254 ( .A(n4212), .B(n4213), .Z(n4211) );
  XOR U4255 ( .A(n4214), .B(n4210), .Z(n4212) );
  XNOR U4256 ( .A(n4215), .B(n4216), .Z(n4209) );
  AND U4257 ( .A(n4217), .B(n4218), .Z(n4216) );
  XOR U4258 ( .A(n4215), .B(n4219), .Z(n4217) );
  XNOR U4259 ( .A(n4200), .B(n4197), .Z(n4208) );
  AND U4260 ( .A(n4220), .B(n4221), .Z(n4197) );
  XOR U4261 ( .A(n4222), .B(n4223), .Z(n4200) );
  AND U4262 ( .A(n4224), .B(n4225), .Z(n4223) );
  XOR U4263 ( .A(n4222), .B(n4226), .Z(n4224) );
  XNOR U4264 ( .A(n4154), .B(n4204), .Z(n4206) );
  XNOR U4265 ( .A(n4227), .B(n4228), .Z(n4154) );
  AND U4266 ( .A(n210), .B(n4229), .Z(n4228) );
  XOR U4267 ( .A(n4230), .B(n4231), .Z(n4204) );
  AND U4268 ( .A(n4232), .B(n4233), .Z(n4231) );
  XNOR U4269 ( .A(n4230), .B(n4220), .Z(n4233) );
  IV U4270 ( .A(n4167), .Z(n4220) );
  XNOR U4271 ( .A(n4234), .B(n4213), .Z(n4167) );
  XNOR U4272 ( .A(n4235), .B(n4219), .Z(n4213) );
  XOR U4273 ( .A(n4236), .B(n4237), .Z(n4219) );
  AND U4274 ( .A(n4238), .B(n4239), .Z(n4237) );
  XOR U4275 ( .A(n4236), .B(n4240), .Z(n4238) );
  XNOR U4276 ( .A(n4218), .B(n4210), .Z(n4235) );
  XOR U4277 ( .A(n4241), .B(n4242), .Z(n4210) );
  AND U4278 ( .A(n4243), .B(n4244), .Z(n4242) );
  XNOR U4279 ( .A(n4245), .B(n4241), .Z(n4243) );
  XNOR U4280 ( .A(n4246), .B(n4215), .Z(n4218) );
  XOR U4281 ( .A(n4247), .B(n4248), .Z(n4215) );
  AND U4282 ( .A(n4249), .B(n4250), .Z(n4248) );
  XOR U4283 ( .A(n4247), .B(n4251), .Z(n4249) );
  XNOR U4284 ( .A(n4252), .B(n4253), .Z(n4246) );
  AND U4285 ( .A(n4254), .B(n4255), .Z(n4253) );
  XNOR U4286 ( .A(n4252), .B(n4256), .Z(n4254) );
  XNOR U4287 ( .A(n4214), .B(n4221), .Z(n4234) );
  AND U4288 ( .A(n4175), .B(n4257), .Z(n4221) );
  XOR U4289 ( .A(n4226), .B(n4225), .Z(n4214) );
  XNOR U4290 ( .A(n4258), .B(n4222), .Z(n4225) );
  XOR U4291 ( .A(n4259), .B(n4260), .Z(n4222) );
  AND U4292 ( .A(n4261), .B(n4262), .Z(n4260) );
  XOR U4293 ( .A(n4259), .B(n4263), .Z(n4261) );
  XNOR U4294 ( .A(n4264), .B(n4265), .Z(n4258) );
  AND U4295 ( .A(n4266), .B(n4267), .Z(n4265) );
  XOR U4296 ( .A(n4264), .B(n4268), .Z(n4266) );
  XOR U4297 ( .A(n4269), .B(n4270), .Z(n4226) );
  AND U4298 ( .A(n4271), .B(n4272), .Z(n4270) );
  XOR U4299 ( .A(n4269), .B(n4273), .Z(n4271) );
  XNOR U4300 ( .A(n4164), .B(n4230), .Z(n4232) );
  XNOR U4301 ( .A(n4274), .B(n4275), .Z(n4164) );
  AND U4302 ( .A(n210), .B(n4276), .Z(n4275) );
  XNOR U4303 ( .A(n4277), .B(n4278), .Z(n4276) );
  XOR U4304 ( .A(n4279), .B(n4280), .Z(n4230) );
  AND U4305 ( .A(n4281), .B(n4282), .Z(n4280) );
  XNOR U4306 ( .A(n4279), .B(n4175), .Z(n4282) );
  XOR U4307 ( .A(n4283), .B(n4244), .Z(n4175) );
  XNOR U4308 ( .A(n4284), .B(n4251), .Z(n4244) );
  XOR U4309 ( .A(n4240), .B(n4239), .Z(n4251) );
  XNOR U4310 ( .A(n4285), .B(n4236), .Z(n4239) );
  XOR U4311 ( .A(n4286), .B(n4287), .Z(n4236) );
  AND U4312 ( .A(n4288), .B(n4289), .Z(n4287) );
  XNOR U4313 ( .A(n4290), .B(n4291), .Z(n4288) );
  IV U4314 ( .A(n4286), .Z(n4290) );
  XNOR U4315 ( .A(n4292), .B(n4293), .Z(n4285) );
  NOR U4316 ( .A(n4294), .B(n4295), .Z(n4293) );
  XNOR U4317 ( .A(n4292), .B(n4296), .Z(n4294) );
  XOR U4318 ( .A(n4297), .B(n4298), .Z(n4240) );
  NOR U4319 ( .A(n4299), .B(n4300), .Z(n4298) );
  XNOR U4320 ( .A(n4297), .B(n4301), .Z(n4299) );
  XNOR U4321 ( .A(n4250), .B(n4241), .Z(n4284) );
  XOR U4322 ( .A(n4302), .B(n4303), .Z(n4241) );
  AND U4323 ( .A(n4304), .B(n4305), .Z(n4303) );
  XOR U4324 ( .A(n4302), .B(n4306), .Z(n4304) );
  XOR U4325 ( .A(n4307), .B(n4256), .Z(n4250) );
  XOR U4326 ( .A(n4308), .B(n4309), .Z(n4256) );
  NOR U4327 ( .A(n4310), .B(n4311), .Z(n4309) );
  XOR U4328 ( .A(n4308), .B(n4312), .Z(n4310) );
  XNOR U4329 ( .A(n4255), .B(n4247), .Z(n4307) );
  XOR U4330 ( .A(n4313), .B(n4314), .Z(n4247) );
  AND U4331 ( .A(n4315), .B(n4316), .Z(n4314) );
  XOR U4332 ( .A(n4313), .B(n4317), .Z(n4315) );
  XNOR U4333 ( .A(n4318), .B(n4252), .Z(n4255) );
  XOR U4334 ( .A(n4319), .B(n4320), .Z(n4252) );
  AND U4335 ( .A(n4321), .B(n4322), .Z(n4320) );
  XNOR U4336 ( .A(n4323), .B(n4324), .Z(n4321) );
  IV U4337 ( .A(n4319), .Z(n4323) );
  XNOR U4338 ( .A(n4325), .B(n4326), .Z(n4318) );
  NOR U4339 ( .A(n4327), .B(n4328), .Z(n4326) );
  XNOR U4340 ( .A(n4325), .B(n4329), .Z(n4327) );
  XOR U4341 ( .A(n4245), .B(n4257), .Z(n4283) );
  NOR U4342 ( .A(n4181), .B(n4330), .Z(n4257) );
  XNOR U4343 ( .A(n4263), .B(n4262), .Z(n4245) );
  XNOR U4344 ( .A(n4331), .B(n4268), .Z(n4262) );
  XNOR U4345 ( .A(n4332), .B(n4333), .Z(n4268) );
  NOR U4346 ( .A(n4334), .B(n4335), .Z(n4333) );
  XOR U4347 ( .A(n4332), .B(n4336), .Z(n4334) );
  XNOR U4348 ( .A(n4267), .B(n4259), .Z(n4331) );
  XOR U4349 ( .A(n4337), .B(n4338), .Z(n4259) );
  AND U4350 ( .A(n4339), .B(n4340), .Z(n4338) );
  XNOR U4351 ( .A(n4341), .B(n4342), .Z(n4339) );
  XNOR U4352 ( .A(n4343), .B(n4264), .Z(n4267) );
  XOR U4353 ( .A(n4344), .B(n4345), .Z(n4264) );
  AND U4354 ( .A(n4346), .B(n4347), .Z(n4345) );
  XNOR U4355 ( .A(n4348), .B(n4349), .Z(n4346) );
  IV U4356 ( .A(n4344), .Z(n4348) );
  XNOR U4357 ( .A(n4350), .B(n4351), .Z(n4343) );
  NOR U4358 ( .A(n4352), .B(n4353), .Z(n4351) );
  XNOR U4359 ( .A(n4350), .B(n4354), .Z(n4352) );
  XOR U4360 ( .A(n4273), .B(n4272), .Z(n4263) );
  XNOR U4361 ( .A(n4355), .B(n4269), .Z(n4272) );
  XOR U4362 ( .A(n4356), .B(n4357), .Z(n4269) );
  AND U4363 ( .A(n4358), .B(n4359), .Z(n4357) );
  XOR U4364 ( .A(n4356), .B(n4360), .Z(n4358) );
  XNOR U4365 ( .A(n4361), .B(n4362), .Z(n4355) );
  NOR U4366 ( .A(n4363), .B(n4364), .Z(n4362) );
  XNOR U4367 ( .A(n4361), .B(n4365), .Z(n4363) );
  XOR U4368 ( .A(n4366), .B(n4367), .Z(n4273) );
  NOR U4369 ( .A(n4368), .B(n4369), .Z(n4367) );
  XNOR U4370 ( .A(n4366), .B(n4370), .Z(n4368) );
  XNOR U4371 ( .A(n4172), .B(n4279), .Z(n4281) );
  XNOR U4372 ( .A(n4371), .B(n4372), .Z(n4172) );
  AND U4373 ( .A(n210), .B(n4373), .Z(n4372) );
  AND U4374 ( .A(n4178), .B(n4181), .Z(n4279) );
  XOR U4375 ( .A(n4374), .B(n4330), .Z(n4181) );
  XNOR U4376 ( .A(p_input[128]), .B(p_input[256]), .Z(n4330) );
  XNOR U4377 ( .A(n4306), .B(n4305), .Z(n4374) );
  XNOR U4378 ( .A(n4375), .B(n4317), .Z(n4305) );
  XOR U4379 ( .A(n4291), .B(n4289), .Z(n4317) );
  XNOR U4380 ( .A(n4376), .B(n4296), .Z(n4289) );
  XOR U4381 ( .A(p_input[152]), .B(p_input[280]), .Z(n4296) );
  XOR U4382 ( .A(n4286), .B(n4295), .Z(n4376) );
  XOR U4383 ( .A(n4377), .B(n4292), .Z(n4295) );
  XOR U4384 ( .A(p_input[150]), .B(p_input[278]), .Z(n4292) );
  XOR U4385 ( .A(p_input[151]), .B(n2951), .Z(n4377) );
  XOR U4386 ( .A(p_input[146]), .B(p_input[274]), .Z(n4286) );
  XNOR U4387 ( .A(n4301), .B(n4300), .Z(n4291) );
  XOR U4388 ( .A(n4378), .B(n4297), .Z(n4300) );
  XOR U4389 ( .A(p_input[147]), .B(p_input[275]), .Z(n4297) );
  XOR U4390 ( .A(p_input[148]), .B(n2953), .Z(n4378) );
  XOR U4391 ( .A(p_input[149]), .B(p_input[277]), .Z(n4301) );
  XOR U4392 ( .A(n4316), .B(n4379), .Z(n4375) );
  IV U4393 ( .A(n4302), .Z(n4379) );
  XOR U4394 ( .A(p_input[129]), .B(p_input[257]), .Z(n4302) );
  XNOR U4395 ( .A(n4380), .B(n4324), .Z(n4316) );
  XNOR U4396 ( .A(n4312), .B(n4311), .Z(n4324) );
  XNOR U4397 ( .A(n4381), .B(n4308), .Z(n4311) );
  XNOR U4398 ( .A(p_input[154]), .B(p_input[282]), .Z(n4308) );
  XOR U4399 ( .A(p_input[155]), .B(n2957), .Z(n4381) );
  XOR U4400 ( .A(p_input[156]), .B(p_input[284]), .Z(n4312) );
  XOR U4401 ( .A(n4322), .B(n4382), .Z(n4380) );
  IV U4402 ( .A(n4313), .Z(n4382) );
  XOR U4403 ( .A(p_input[145]), .B(p_input[273]), .Z(n4313) );
  XNOR U4404 ( .A(n4383), .B(n4329), .Z(n4322) );
  XOR U4405 ( .A(p_input[159]), .B(p_input[287]), .Z(n4329) );
  XOR U4406 ( .A(n4319), .B(n4328), .Z(n4383) );
  XOR U4407 ( .A(n4384), .B(n4325), .Z(n4328) );
  XOR U4408 ( .A(p_input[157]), .B(p_input[285]), .Z(n4325) );
  XOR U4409 ( .A(p_input[158]), .B(n4385), .Z(n4384) );
  XOR U4410 ( .A(p_input[153]), .B(p_input[281]), .Z(n4319) );
  XOR U4411 ( .A(n4342), .B(n4340), .Z(n4306) );
  XNOR U4412 ( .A(n4386), .B(n4349), .Z(n4340) );
  XNOR U4413 ( .A(n4336), .B(n4335), .Z(n4349) );
  XNOR U4414 ( .A(n4387), .B(n4332), .Z(n4335) );
  XNOR U4415 ( .A(p_input[139]), .B(p_input[267]), .Z(n4332) );
  XOR U4416 ( .A(p_input[140]), .B(n2963), .Z(n4387) );
  XOR U4417 ( .A(p_input[141]), .B(p_input[269]), .Z(n4336) );
  XOR U4418 ( .A(n4347), .B(n4341), .Z(n4386) );
  IV U4419 ( .A(n4337), .Z(n4341) );
  XOR U4420 ( .A(p_input[130]), .B(p_input[258]), .Z(n4337) );
  XNOR U4421 ( .A(n4388), .B(n4354), .Z(n4347) );
  XNOR U4422 ( .A(p_input[144]), .B(n2965), .Z(n4354) );
  IV U4423 ( .A(p_input[272]), .Z(n2965) );
  XOR U4424 ( .A(n4344), .B(n4353), .Z(n4388) );
  XOR U4425 ( .A(n4389), .B(n4350), .Z(n4353) );
  XOR U4426 ( .A(p_input[142]), .B(p_input[270]), .Z(n4350) );
  XOR U4427 ( .A(p_input[143]), .B(n2967), .Z(n4389) );
  XOR U4428 ( .A(p_input[138]), .B(p_input[266]), .Z(n4344) );
  XOR U4429 ( .A(n4360), .B(n4359), .Z(n4342) );
  XNOR U4430 ( .A(n4390), .B(n4365), .Z(n4359) );
  XOR U4431 ( .A(p_input[137]), .B(p_input[265]), .Z(n4365) );
  XOR U4432 ( .A(n4356), .B(n4364), .Z(n4390) );
  XOR U4433 ( .A(n4391), .B(n4361), .Z(n4364) );
  XOR U4434 ( .A(p_input[135]), .B(p_input[263]), .Z(n4361) );
  XOR U4435 ( .A(p_input[136]), .B(n4392), .Z(n4391) );
  XOR U4436 ( .A(p_input[131]), .B(p_input[259]), .Z(n4356) );
  XNOR U4437 ( .A(n4370), .B(n4369), .Z(n4360) );
  XOR U4438 ( .A(n4393), .B(n4366), .Z(n4369) );
  XOR U4439 ( .A(p_input[132]), .B(p_input[260]), .Z(n4366) );
  XOR U4440 ( .A(p_input[133]), .B(n4394), .Z(n4393) );
  XOR U4441 ( .A(p_input[134]), .B(p_input[262]), .Z(n4370) );
  XNOR U4442 ( .A(n4395), .B(n4396), .Z(n4178) );
  AND U4443 ( .A(n210), .B(n4397), .Z(n4396) );
  XNOR U4444 ( .A(n4398), .B(n4399), .Z(n210) );
  NOR U4445 ( .A(n4400), .B(n4401), .Z(n4399) );
  XOR U4446 ( .A(n4398), .B(n4186), .Z(n4401) );
  XNOR U4447 ( .A(n4402), .B(n4403), .Z(n4131) );
  AND U4448 ( .A(n214), .B(n4404), .Z(n4403) );
  XNOR U4449 ( .A(n4405), .B(n4406), .Z(n214) );
  NOR U4450 ( .A(n4407), .B(n4408), .Z(n4406) );
  XOR U4451 ( .A(n4093), .B(n4405), .Z(n4408) );
  NOR U4452 ( .A(n4405), .B(n4092), .Z(n4407) );
  XOR U4453 ( .A(n4409), .B(n4410), .Z(n4405) );
  AND U4454 ( .A(n4411), .B(n4412), .Z(n4410) );
  XNOR U4455 ( .A(n4148), .B(n4409), .Z(n4412) );
  XOR U4456 ( .A(n4409), .B(n4101), .Z(n4411) );
  XOR U4457 ( .A(n4413), .B(n4414), .Z(n4409) );
  AND U4458 ( .A(n4415), .B(n4416), .Z(n4414) );
  XNOR U4459 ( .A(n4158), .B(n4413), .Z(n4416) );
  XOR U4460 ( .A(n4413), .B(n4110), .Z(n4415) );
  XOR U4461 ( .A(n4417), .B(n4418), .Z(n4413) );
  AND U4462 ( .A(n4419), .B(n4420), .Z(n4418) );
  XOR U4463 ( .A(n4417), .B(n4118), .Z(n4419) );
  XOR U4464 ( .A(n4421), .B(n4422), .Z(n4085) );
  AND U4465 ( .A(n218), .B(n4404), .Z(n4422) );
  XNOR U4466 ( .A(n4402), .B(n4421), .Z(n4404) );
  XNOR U4467 ( .A(n4423), .B(n4424), .Z(n218) );
  NOR U4468 ( .A(n4425), .B(n4426), .Z(n4424) );
  XNOR U4469 ( .A(n4093), .B(n4427), .Z(n4426) );
  IV U4470 ( .A(n4423), .Z(n4427) );
  AND U4471 ( .A(n4428), .B(n4429), .Z(n4093) );
  NOR U4472 ( .A(n4423), .B(n4092), .Z(n4425) );
  AND U4473 ( .A(n4186), .B(n4187), .Z(n4092) );
  IV U4474 ( .A(n4430), .Z(n4186) );
  XOR U4475 ( .A(n4431), .B(n4432), .Z(n4423) );
  AND U4476 ( .A(n4433), .B(n4434), .Z(n4432) );
  XNOR U4477 ( .A(n4431), .B(n4148), .Z(n4434) );
  XOR U4478 ( .A(n4435), .B(n4436), .Z(n4148) );
  AND U4479 ( .A(n221), .B(n4203), .Z(n4436) );
  XOR U4480 ( .A(n4201), .B(n4435), .Z(n4203) );
  XNOR U4481 ( .A(n4437), .B(n4431), .Z(n4433) );
  IV U4482 ( .A(n4101), .Z(n4437) );
  XOR U4483 ( .A(n4438), .B(n4439), .Z(n4101) );
  AND U4484 ( .A(n226), .B(n4440), .Z(n4439) );
  XOR U4485 ( .A(n4441), .B(n4442), .Z(n4431) );
  AND U4486 ( .A(n4443), .B(n4444), .Z(n4442) );
  XNOR U4487 ( .A(n4441), .B(n4158), .Z(n4444) );
  XOR U4488 ( .A(n4445), .B(n4446), .Z(n4158) );
  AND U4489 ( .A(n221), .B(n4229), .Z(n4446) );
  XOR U4490 ( .A(n4227), .B(n4445), .Z(n4229) );
  XOR U4491 ( .A(n4110), .B(n4441), .Z(n4443) );
  XOR U4492 ( .A(n4447), .B(n4448), .Z(n4110) );
  AND U4493 ( .A(n226), .B(n4449), .Z(n4448) );
  XOR U4494 ( .A(n4417), .B(n4450), .Z(n4441) );
  AND U4495 ( .A(n4451), .B(n4420), .Z(n4450) );
  XNOR U4496 ( .A(n4168), .B(n4417), .Z(n4420) );
  XOR U4497 ( .A(n4278), .B(n4452), .Z(n4168) );
  AND U4498 ( .A(n221), .B(n4453), .Z(n4452) );
  XOR U4499 ( .A(n4274), .B(n4278), .Z(n4453) );
  XNOR U4500 ( .A(n4454), .B(n4417), .Z(n4451) );
  IV U4501 ( .A(n4118), .Z(n4454) );
  XOR U4502 ( .A(n4455), .B(n4456), .Z(n4118) );
  AND U4503 ( .A(n226), .B(n4457), .Z(n4456) );
  XOR U4504 ( .A(n4458), .B(n4459), .Z(n4417) );
  AND U4505 ( .A(n4460), .B(n4461), .Z(n4459) );
  XNOR U4506 ( .A(n4458), .B(n4176), .Z(n4461) );
  XNOR U4507 ( .A(n4462), .B(n4463), .Z(n4176) );
  AND U4508 ( .A(n221), .B(n4373), .Z(n4463) );
  XOR U4509 ( .A(n4371), .B(n4464), .Z(n4373) );
  IV U4510 ( .A(n4462), .Z(n4464) );
  XNOR U4511 ( .A(n4465), .B(n4458), .Z(n4460) );
  IV U4512 ( .A(n4128), .Z(n4465) );
  XOR U4513 ( .A(n4466), .B(n4467), .Z(n4128) );
  AND U4514 ( .A(n226), .B(n4468), .Z(n4467) );
  AND U4515 ( .A(n4421), .B(n4402), .Z(n4458) );
  XNOR U4516 ( .A(n4469), .B(n4470), .Z(n4402) );
  AND U4517 ( .A(n221), .B(n4397), .Z(n4470) );
  XOR U4518 ( .A(n4471), .B(n4469), .Z(n4397) );
  XNOR U4519 ( .A(n4398), .B(n4472), .Z(n221) );
  NOR U4520 ( .A(n4400), .B(n4473), .Z(n4472) );
  XNOR U4521 ( .A(n4398), .B(n4430), .Z(n4473) );
  NOR U4522 ( .A(n4428), .B(n4429), .Z(n4430) );
  NOR U4523 ( .A(n4398), .B(n4187), .Z(n4400) );
  AND U4524 ( .A(n4201), .B(n4474), .Z(n4187) );
  XOR U4525 ( .A(n4475), .B(n4476), .Z(n4398) );
  AND U4526 ( .A(n4477), .B(n4478), .Z(n4476) );
  XNOR U4527 ( .A(n4201), .B(n4475), .Z(n4478) );
  XNOR U4528 ( .A(n4479), .B(n4480), .Z(n4201) );
  XOR U4529 ( .A(n4481), .B(n4474), .Z(n4480) );
  AND U4530 ( .A(n4227), .B(n4482), .Z(n4474) );
  AND U4531 ( .A(n4483), .B(n4484), .Z(n4481) );
  XOR U4532 ( .A(n4485), .B(n4479), .Z(n4483) );
  XOR U4533 ( .A(n4475), .B(n4435), .Z(n4477) );
  XOR U4534 ( .A(n4486), .B(n4487), .Z(n4435) );
  AND U4535 ( .A(n223), .B(n4440), .Z(n4487) );
  XOR U4536 ( .A(n4486), .B(n4438), .Z(n4440) );
  XOR U4537 ( .A(n4488), .B(n4489), .Z(n4475) );
  AND U4538 ( .A(n4490), .B(n4491), .Z(n4489) );
  XNOR U4539 ( .A(n4227), .B(n4488), .Z(n4491) );
  XOR U4540 ( .A(n4492), .B(n4484), .Z(n4227) );
  XNOR U4541 ( .A(n4493), .B(n4479), .Z(n4484) );
  XOR U4542 ( .A(n4494), .B(n4495), .Z(n4479) );
  AND U4543 ( .A(n4496), .B(n4497), .Z(n4495) );
  XOR U4544 ( .A(n4498), .B(n4494), .Z(n4496) );
  XNOR U4545 ( .A(n4499), .B(n4500), .Z(n4493) );
  AND U4546 ( .A(n4501), .B(n4502), .Z(n4500) );
  XOR U4547 ( .A(n4499), .B(n4503), .Z(n4501) );
  XNOR U4548 ( .A(n4485), .B(n4482), .Z(n4492) );
  AND U4549 ( .A(n4274), .B(n4504), .Z(n4482) );
  XOR U4550 ( .A(n4505), .B(n4506), .Z(n4485) );
  AND U4551 ( .A(n4507), .B(n4508), .Z(n4506) );
  XOR U4552 ( .A(n4505), .B(n4509), .Z(n4507) );
  XOR U4553 ( .A(n4488), .B(n4445), .Z(n4490) );
  XOR U4554 ( .A(n4510), .B(n4511), .Z(n4445) );
  AND U4555 ( .A(n223), .B(n4449), .Z(n4511) );
  XOR U4556 ( .A(n4510), .B(n4447), .Z(n4449) );
  XOR U4557 ( .A(n4512), .B(n4513), .Z(n4488) );
  AND U4558 ( .A(n4514), .B(n4515), .Z(n4513) );
  XNOR U4559 ( .A(n4274), .B(n4512), .Z(n4515) );
  IV U4560 ( .A(n4277), .Z(n4274) );
  XNOR U4561 ( .A(n4516), .B(n4497), .Z(n4277) );
  XNOR U4562 ( .A(n4517), .B(n4503), .Z(n4497) );
  XOR U4563 ( .A(n4518), .B(n4519), .Z(n4503) );
  AND U4564 ( .A(n4520), .B(n4521), .Z(n4519) );
  XOR U4565 ( .A(n4518), .B(n4522), .Z(n4520) );
  XNOR U4566 ( .A(n4502), .B(n4494), .Z(n4517) );
  XOR U4567 ( .A(n4523), .B(n4524), .Z(n4494) );
  AND U4568 ( .A(n4525), .B(n4526), .Z(n4524) );
  XNOR U4569 ( .A(n4527), .B(n4523), .Z(n4525) );
  XNOR U4570 ( .A(n4528), .B(n4499), .Z(n4502) );
  XOR U4571 ( .A(n4529), .B(n4530), .Z(n4499) );
  AND U4572 ( .A(n4531), .B(n4532), .Z(n4530) );
  XOR U4573 ( .A(n4529), .B(n4533), .Z(n4531) );
  XNOR U4574 ( .A(n4534), .B(n4535), .Z(n4528) );
  AND U4575 ( .A(n4536), .B(n4537), .Z(n4535) );
  XNOR U4576 ( .A(n4534), .B(n4538), .Z(n4536) );
  XNOR U4577 ( .A(n4498), .B(n4504), .Z(n4516) );
  AND U4578 ( .A(n4371), .B(n4539), .Z(n4504) );
  XOR U4579 ( .A(n4509), .B(n4508), .Z(n4498) );
  XNOR U4580 ( .A(n4540), .B(n4505), .Z(n4508) );
  XOR U4581 ( .A(n4541), .B(n4542), .Z(n4505) );
  AND U4582 ( .A(n4543), .B(n4544), .Z(n4542) );
  XOR U4583 ( .A(n4541), .B(n4545), .Z(n4543) );
  XNOR U4584 ( .A(n4546), .B(n4547), .Z(n4540) );
  AND U4585 ( .A(n4548), .B(n4549), .Z(n4547) );
  XOR U4586 ( .A(n4546), .B(n4550), .Z(n4548) );
  XOR U4587 ( .A(n4551), .B(n4552), .Z(n4509) );
  AND U4588 ( .A(n4553), .B(n4554), .Z(n4552) );
  XOR U4589 ( .A(n4551), .B(n4555), .Z(n4553) );
  XOR U4590 ( .A(n4512), .B(n4278), .Z(n4514) );
  XOR U4591 ( .A(n4556), .B(n4557), .Z(n4278) );
  AND U4592 ( .A(n223), .B(n4457), .Z(n4557) );
  XOR U4593 ( .A(n4556), .B(n4455), .Z(n4457) );
  XOR U4594 ( .A(n4558), .B(n4559), .Z(n4512) );
  AND U4595 ( .A(n4560), .B(n4561), .Z(n4559) );
  XNOR U4596 ( .A(n4558), .B(n4371), .Z(n4561) );
  XOR U4597 ( .A(n4562), .B(n4526), .Z(n4371) );
  XNOR U4598 ( .A(n4563), .B(n4533), .Z(n4526) );
  XOR U4599 ( .A(n4522), .B(n4521), .Z(n4533) );
  XNOR U4600 ( .A(n4564), .B(n4518), .Z(n4521) );
  XOR U4601 ( .A(n4565), .B(n4566), .Z(n4518) );
  AND U4602 ( .A(n4567), .B(n4568), .Z(n4566) );
  XOR U4603 ( .A(n4565), .B(n4569), .Z(n4567) );
  XNOR U4604 ( .A(n4570), .B(n4571), .Z(n4564) );
  NOR U4605 ( .A(n4572), .B(n4573), .Z(n4571) );
  XNOR U4606 ( .A(n4570), .B(n4574), .Z(n4572) );
  XOR U4607 ( .A(n4575), .B(n4576), .Z(n4522) );
  NOR U4608 ( .A(n4577), .B(n4578), .Z(n4576) );
  XNOR U4609 ( .A(n4575), .B(n4579), .Z(n4577) );
  XNOR U4610 ( .A(n4532), .B(n4523), .Z(n4563) );
  XOR U4611 ( .A(n4580), .B(n4581), .Z(n4523) );
  NOR U4612 ( .A(n4582), .B(n4583), .Z(n4581) );
  XNOR U4613 ( .A(n4580), .B(n4584), .Z(n4582) );
  XOR U4614 ( .A(n4585), .B(n4538), .Z(n4532) );
  XNOR U4615 ( .A(n4586), .B(n4587), .Z(n4538) );
  NOR U4616 ( .A(n4588), .B(n4589), .Z(n4587) );
  XNOR U4617 ( .A(n4586), .B(n4590), .Z(n4588) );
  XNOR U4618 ( .A(n4537), .B(n4529), .Z(n4585) );
  XOR U4619 ( .A(n4591), .B(n4592), .Z(n4529) );
  AND U4620 ( .A(n4593), .B(n4594), .Z(n4592) );
  XOR U4621 ( .A(n4591), .B(n4595), .Z(n4593) );
  XNOR U4622 ( .A(n4596), .B(n4534), .Z(n4537) );
  XOR U4623 ( .A(n4597), .B(n4598), .Z(n4534) );
  AND U4624 ( .A(n4599), .B(n4600), .Z(n4598) );
  XOR U4625 ( .A(n4597), .B(n4601), .Z(n4599) );
  XNOR U4626 ( .A(n4602), .B(n4603), .Z(n4596) );
  NOR U4627 ( .A(n4604), .B(n4605), .Z(n4603) );
  XOR U4628 ( .A(n4602), .B(n4606), .Z(n4604) );
  XOR U4629 ( .A(n4527), .B(n4539), .Z(n4562) );
  AND U4630 ( .A(n4471), .B(n4607), .Z(n4539) );
  IV U4631 ( .A(n4395), .Z(n4471) );
  XNOR U4632 ( .A(n4545), .B(n4544), .Z(n4527) );
  XNOR U4633 ( .A(n4608), .B(n4550), .Z(n4544) );
  XOR U4634 ( .A(n4609), .B(n4610), .Z(n4550) );
  NOR U4635 ( .A(n4611), .B(n4612), .Z(n4610) );
  XNOR U4636 ( .A(n4609), .B(n4613), .Z(n4611) );
  XNOR U4637 ( .A(n4549), .B(n4541), .Z(n4608) );
  XOR U4638 ( .A(n4614), .B(n4615), .Z(n4541) );
  AND U4639 ( .A(n4616), .B(n4617), .Z(n4615) );
  XNOR U4640 ( .A(n4614), .B(n4618), .Z(n4616) );
  XNOR U4641 ( .A(n4619), .B(n4546), .Z(n4549) );
  XOR U4642 ( .A(n4620), .B(n4621), .Z(n4546) );
  AND U4643 ( .A(n4622), .B(n4623), .Z(n4621) );
  XOR U4644 ( .A(n4620), .B(n4624), .Z(n4622) );
  XNOR U4645 ( .A(n4625), .B(n4626), .Z(n4619) );
  NOR U4646 ( .A(n4627), .B(n4628), .Z(n4626) );
  XOR U4647 ( .A(n4625), .B(n4629), .Z(n4627) );
  XOR U4648 ( .A(n4555), .B(n4554), .Z(n4545) );
  XNOR U4649 ( .A(n4630), .B(n4551), .Z(n4554) );
  XOR U4650 ( .A(n4631), .B(n4632), .Z(n4551) );
  AND U4651 ( .A(n4633), .B(n4634), .Z(n4632) );
  XOR U4652 ( .A(n4631), .B(n4635), .Z(n4633) );
  XNOR U4653 ( .A(n4636), .B(n4637), .Z(n4630) );
  NOR U4654 ( .A(n4638), .B(n4639), .Z(n4637) );
  XNOR U4655 ( .A(n4636), .B(n4640), .Z(n4638) );
  XOR U4656 ( .A(n4641), .B(n4642), .Z(n4555) );
  NOR U4657 ( .A(n4643), .B(n4644), .Z(n4642) );
  XNOR U4658 ( .A(n4641), .B(n4645), .Z(n4643) );
  XNOR U4659 ( .A(n4462), .B(n4558), .Z(n4560) );
  XNOR U4660 ( .A(n4646), .B(n4647), .Z(n4462) );
  AND U4661 ( .A(n223), .B(n4468), .Z(n4647) );
  XOR U4662 ( .A(n4646), .B(n4466), .Z(n4468) );
  AND U4663 ( .A(n4469), .B(n4395), .Z(n4558) );
  XNOR U4664 ( .A(n4648), .B(n4607), .Z(n4395) );
  XOR U4665 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(
        p_input[256]), .Z(n4607) );
  XOR U4666 ( .A(n4584), .B(n4583), .Z(n4648) );
  XOR U4667 ( .A(n4649), .B(n4595), .Z(n4583) );
  XOR U4668 ( .A(n4569), .B(n4568), .Z(n4595) );
  XNOR U4669 ( .A(n4650), .B(n4574), .Z(n4568) );
  XOR U4670 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][24] ), .B(
        p_input[280]), .Z(n4574) );
  XOR U4671 ( .A(n4565), .B(n4573), .Z(n4650) );
  XOR U4672 ( .A(n4651), .B(n4570), .Z(n4573) );
  XOR U4673 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][22] ), .B(
        p_input[278]), .Z(n4570) );
  XOR U4674 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][23] ), .B(n2951), 
        .Z(n4651) );
  XNOR U4675 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][18] ), .B(n3316), 
        .Z(n4565) );
  XNOR U4676 ( .A(n4579), .B(n4578), .Z(n4569) );
  XOR U4677 ( .A(n4652), .B(n4575), .Z(n4578) );
  XOR U4678 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][19] ), .B(
        p_input[275]), .Z(n4575) );
  XOR U4679 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][20] ), .B(n2953), 
        .Z(n4652) );
  XOR U4680 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][21] ), .B(
        p_input[277]), .Z(n4579) );
  XNOR U4681 ( .A(n4594), .B(n4580), .Z(n4649) );
  XNOR U4682 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n3318), 
        .Z(n4580) );
  XNOR U4683 ( .A(n4653), .B(n4601), .Z(n4594) );
  XNOR U4684 ( .A(n4590), .B(n4589), .Z(n4601) );
  XOR U4685 ( .A(n4654), .B(n4586), .Z(n4589) );
  XNOR U4686 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][26] ), .B(n3321), 
        .Z(n4586) );
  XOR U4687 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][27] ), .B(n2957), 
        .Z(n4654) );
  XOR U4688 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][28] ), .B(
        p_input[284]), .Z(n4590) );
  XNOR U4689 ( .A(n4600), .B(n4591), .Z(n4653) );
  XNOR U4690 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][17] ), .B(n3322), 
        .Z(n4591) );
  XOR U4691 ( .A(n4655), .B(n4606), .Z(n4600) );
  XNOR U4692 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][31] ), .B(
        p_input[287]), .Z(n4606) );
  XOR U4693 ( .A(n4597), .B(n4605), .Z(n4655) );
  XOR U4694 ( .A(n4656), .B(n4602), .Z(n4605) );
  XOR U4695 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][29] ), .B(
        p_input[285]), .Z(n4602) );
  XOR U4696 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][30] ), .B(n4385), 
        .Z(n4656) );
  XNOR U4697 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][25] ), .B(n3325), 
        .Z(n4597) );
  XNOR U4698 ( .A(n4618), .B(n4617), .Z(n4584) );
  XNOR U4699 ( .A(n4657), .B(n4624), .Z(n4617) );
  XNOR U4700 ( .A(n4613), .B(n4612), .Z(n4624) );
  XOR U4701 ( .A(n4658), .B(n4609), .Z(n4612) );
  XNOR U4702 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n3328), 
        .Z(n4609) );
  XOR U4703 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n2963), 
        .Z(n4658) );
  XOR U4704 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(
        p_input[269]), .Z(n4613) );
  XNOR U4705 ( .A(n4623), .B(n4614), .Z(n4657) );
  XOR U4706 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(
        p_input[258]), .Z(n4614) );
  XOR U4707 ( .A(n4659), .B(n4629), .Z(n4623) );
  XNOR U4708 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][16] ), .B(
        p_input[272]), .Z(n4629) );
  XOR U4709 ( .A(n4620), .B(n4628), .Z(n4659) );
  XOR U4710 ( .A(n4660), .B(n4625), .Z(n4628) );
  XOR U4711 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(
        p_input[270]), .Z(n4625) );
  XOR U4712 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n2967), 
        .Z(n4660) );
  XNOR U4713 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n3331), 
        .Z(n4620) );
  XNOR U4714 ( .A(n4635), .B(n4634), .Z(n4618) );
  XNOR U4715 ( .A(n4661), .B(n4640), .Z(n4634) );
  XOR U4716 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(
        p_input[265]), .Z(n4640) );
  XOR U4717 ( .A(n4631), .B(n4639), .Z(n4661) );
  XOR U4718 ( .A(n4662), .B(n4636), .Z(n4639) );
  XOR U4719 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(
        p_input[263]), .Z(n4636) );
  XOR U4720 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n4392), 
        .Z(n4662) );
  XOR U4721 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(
        p_input[259]), .Z(n4631) );
  XNOR U4722 ( .A(n4645), .B(n4644), .Z(n4635) );
  XOR U4723 ( .A(n4663), .B(n4641), .Z(n4644) );
  XOR U4724 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(
        p_input[260]), .Z(n4641) );
  XOR U4725 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n4394), 
        .Z(n4663) );
  XOR U4726 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(
        p_input[262]), .Z(n4645) );
  XNOR U4727 ( .A(n4664), .B(n4665), .Z(n4469) );
  AND U4728 ( .A(n223), .B(n4666), .Z(n4665) );
  XNOR U4729 ( .A(n4667), .B(n4668), .Z(n223) );
  NOR U4730 ( .A(n4669), .B(n4670), .Z(n4668) );
  XOR U4731 ( .A(n4429), .B(n4667), .Z(n4670) );
  NOR U4732 ( .A(n4667), .B(n4428), .Z(n4669) );
  XOR U4733 ( .A(n4671), .B(n4672), .Z(n4667) );
  AND U4734 ( .A(n4673), .B(n4674), .Z(n4672) );
  XNOR U4735 ( .A(n4486), .B(n4671), .Z(n4674) );
  XOR U4736 ( .A(n4671), .B(n4438), .Z(n4673) );
  XOR U4737 ( .A(n4675), .B(n4676), .Z(n4671) );
  AND U4738 ( .A(n4677), .B(n4678), .Z(n4676) );
  XNOR U4739 ( .A(n4510), .B(n4675), .Z(n4678) );
  XOR U4740 ( .A(n4675), .B(n4447), .Z(n4677) );
  XOR U4741 ( .A(n4679), .B(n4680), .Z(n4675) );
  AND U4742 ( .A(n4681), .B(n4682), .Z(n4680) );
  XOR U4743 ( .A(n4679), .B(n4455), .Z(n4681) );
  XOR U4744 ( .A(n4683), .B(n4684), .Z(n4421) );
  AND U4745 ( .A(n226), .B(n4666), .Z(n4684) );
  XOR U4746 ( .A(n4685), .B(n4683), .Z(n4666) );
  XNOR U4747 ( .A(n4686), .B(n4687), .Z(n226) );
  NOR U4748 ( .A(n4688), .B(n4689), .Z(n4687) );
  XNOR U4749 ( .A(n4429), .B(n4690), .Z(n4689) );
  IV U4750 ( .A(n4686), .Z(n4690) );
  AND U4751 ( .A(n4438), .B(n4691), .Z(n4429) );
  NOR U4752 ( .A(n4686), .B(n4428), .Z(n4688) );
  AND U4753 ( .A(n4486), .B(n4692), .Z(n4428) );
  XOR U4754 ( .A(n4693), .B(n4694), .Z(n4686) );
  AND U4755 ( .A(n4695), .B(n4696), .Z(n4694) );
  XNOR U4756 ( .A(n4693), .B(n4486), .Z(n4696) );
  XNOR U4757 ( .A(n4697), .B(n4698), .Z(n4486) );
  XOR U4758 ( .A(n4699), .B(n4692), .Z(n4698) );
  AND U4759 ( .A(n4510), .B(n4700), .Z(n4692) );
  AND U4760 ( .A(n4701), .B(n4702), .Z(n4699) );
  XOR U4761 ( .A(n4703), .B(n4697), .Z(n4701) );
  XNOR U4762 ( .A(n4704), .B(n4693), .Z(n4695) );
  IV U4763 ( .A(n4438), .Z(n4704) );
  XNOR U4764 ( .A(n4705), .B(n4706), .Z(n4438) );
  XOR U4765 ( .A(n4707), .B(n4691), .Z(n4706) );
  AND U4766 ( .A(n4447), .B(n4708), .Z(n4691) );
  AND U4767 ( .A(n4709), .B(n4710), .Z(n4707) );
  XNOR U4768 ( .A(n4705), .B(n4711), .Z(n4709) );
  XOR U4769 ( .A(n4712), .B(n4713), .Z(n4693) );
  AND U4770 ( .A(n4714), .B(n4715), .Z(n4713) );
  XNOR U4771 ( .A(n4712), .B(n4510), .Z(n4715) );
  XOR U4772 ( .A(n4716), .B(n4702), .Z(n4510) );
  XNOR U4773 ( .A(n4717), .B(n4697), .Z(n4702) );
  XOR U4774 ( .A(n4718), .B(n4719), .Z(n4697) );
  AND U4775 ( .A(n4720), .B(n4721), .Z(n4719) );
  XOR U4776 ( .A(n4722), .B(n4718), .Z(n4720) );
  XNOR U4777 ( .A(n4723), .B(n4724), .Z(n4717) );
  AND U4778 ( .A(n4725), .B(n4726), .Z(n4724) );
  XOR U4779 ( .A(n4723), .B(n4727), .Z(n4725) );
  XNOR U4780 ( .A(n4703), .B(n4700), .Z(n4716) );
  AND U4781 ( .A(n4556), .B(n4728), .Z(n4700) );
  XOR U4782 ( .A(n4729), .B(n4730), .Z(n4703) );
  AND U4783 ( .A(n4731), .B(n4732), .Z(n4730) );
  XOR U4784 ( .A(n4729), .B(n4733), .Z(n4731) );
  XOR U4785 ( .A(n4447), .B(n4712), .Z(n4714) );
  XNOR U4786 ( .A(n4734), .B(n4711), .Z(n4447) );
  XNOR U4787 ( .A(n4735), .B(n4736), .Z(n4711) );
  AND U4788 ( .A(n4737), .B(n4738), .Z(n4736) );
  XOR U4789 ( .A(n4735), .B(n4739), .Z(n4737) );
  XNOR U4790 ( .A(n4710), .B(n4708), .Z(n4734) );
  AND U4791 ( .A(n4455), .B(n4740), .Z(n4708) );
  XNOR U4792 ( .A(n4741), .B(n4705), .Z(n4710) );
  XOR U4793 ( .A(n4742), .B(n4743), .Z(n4705) );
  AND U4794 ( .A(n4744), .B(n4745), .Z(n4743) );
  XOR U4795 ( .A(n4742), .B(n4746), .Z(n4744) );
  XNOR U4796 ( .A(n4747), .B(n4748), .Z(n4741) );
  AND U4797 ( .A(n4749), .B(n4750), .Z(n4748) );
  XNOR U4798 ( .A(n4747), .B(n4751), .Z(n4749) );
  XOR U4799 ( .A(n4679), .B(n4752), .Z(n4712) );
  AND U4800 ( .A(n4753), .B(n4682), .Z(n4752) );
  XNOR U4801 ( .A(n4556), .B(n4679), .Z(n4682) );
  XOR U4802 ( .A(n4754), .B(n4721), .Z(n4556) );
  XNOR U4803 ( .A(n4755), .B(n4727), .Z(n4721) );
  XOR U4804 ( .A(n4756), .B(n4757), .Z(n4727) );
  AND U4805 ( .A(n4758), .B(n4759), .Z(n4757) );
  XOR U4806 ( .A(n4756), .B(n4760), .Z(n4758) );
  XNOR U4807 ( .A(n4726), .B(n4718), .Z(n4755) );
  XOR U4808 ( .A(n4761), .B(n4762), .Z(n4718) );
  AND U4809 ( .A(n4763), .B(n4764), .Z(n4762) );
  XNOR U4810 ( .A(n4765), .B(n4761), .Z(n4763) );
  XNOR U4811 ( .A(n4766), .B(n4723), .Z(n4726) );
  XOR U4812 ( .A(n4767), .B(n4768), .Z(n4723) );
  AND U4813 ( .A(n4769), .B(n4770), .Z(n4768) );
  XOR U4814 ( .A(n4767), .B(n4771), .Z(n4769) );
  XNOR U4815 ( .A(n4772), .B(n4773), .Z(n4766) );
  AND U4816 ( .A(n4774), .B(n4775), .Z(n4773) );
  XNOR U4817 ( .A(n4772), .B(n4776), .Z(n4774) );
  XNOR U4818 ( .A(n4722), .B(n4728), .Z(n4754) );
  AND U4819 ( .A(n4646), .B(n4777), .Z(n4728) );
  XOR U4820 ( .A(n4733), .B(n4732), .Z(n4722) );
  XNOR U4821 ( .A(n4778), .B(n4729), .Z(n4732) );
  XOR U4822 ( .A(n4779), .B(n4780), .Z(n4729) );
  AND U4823 ( .A(n4781), .B(n4782), .Z(n4780) );
  XOR U4824 ( .A(n4779), .B(n4783), .Z(n4781) );
  XNOR U4825 ( .A(n4784), .B(n4785), .Z(n4778) );
  AND U4826 ( .A(n4786), .B(n4787), .Z(n4785) );
  XOR U4827 ( .A(n4784), .B(n4788), .Z(n4786) );
  XOR U4828 ( .A(n4789), .B(n4790), .Z(n4733) );
  AND U4829 ( .A(n4791), .B(n4792), .Z(n4790) );
  XOR U4830 ( .A(n4789), .B(n4793), .Z(n4791) );
  XNOR U4831 ( .A(n4794), .B(n4679), .Z(n4753) );
  IV U4832 ( .A(n4455), .Z(n4794) );
  XOR U4833 ( .A(n4795), .B(n4746), .Z(n4455) );
  XOR U4834 ( .A(n4739), .B(n4738), .Z(n4746) );
  XNOR U4835 ( .A(n4796), .B(n4735), .Z(n4738) );
  XOR U4836 ( .A(n4797), .B(n4798), .Z(n4735) );
  AND U4837 ( .A(n4799), .B(n4800), .Z(n4798) );
  XOR U4838 ( .A(n4797), .B(n4801), .Z(n4799) );
  XNOR U4839 ( .A(n4802), .B(n4803), .Z(n4796) );
  AND U4840 ( .A(n4804), .B(n4805), .Z(n4803) );
  XOR U4841 ( .A(n4802), .B(n4806), .Z(n4804) );
  XOR U4842 ( .A(n4807), .B(n4808), .Z(n4739) );
  AND U4843 ( .A(n4809), .B(n4810), .Z(n4808) );
  XOR U4844 ( .A(n4807), .B(n4811), .Z(n4809) );
  XNOR U4845 ( .A(n4745), .B(n4740), .Z(n4795) );
  AND U4846 ( .A(n4466), .B(n4812), .Z(n4740) );
  XOR U4847 ( .A(n4813), .B(n4751), .Z(n4745) );
  XNOR U4848 ( .A(n4814), .B(n4815), .Z(n4751) );
  AND U4849 ( .A(n4816), .B(n4817), .Z(n4815) );
  XOR U4850 ( .A(n4814), .B(n4818), .Z(n4816) );
  XNOR U4851 ( .A(n4750), .B(n4742), .Z(n4813) );
  XOR U4852 ( .A(n4819), .B(n4820), .Z(n4742) );
  AND U4853 ( .A(n4821), .B(n4822), .Z(n4820) );
  XOR U4854 ( .A(n4819), .B(n4823), .Z(n4821) );
  XNOR U4855 ( .A(n4824), .B(n4747), .Z(n4750) );
  XOR U4856 ( .A(n4825), .B(n4826), .Z(n4747) );
  AND U4857 ( .A(n4827), .B(n4828), .Z(n4826) );
  XOR U4858 ( .A(n4825), .B(n4829), .Z(n4827) );
  XNOR U4859 ( .A(n4830), .B(n4831), .Z(n4824) );
  AND U4860 ( .A(n4832), .B(n4833), .Z(n4831) );
  XNOR U4861 ( .A(n4830), .B(n4834), .Z(n4832) );
  XOR U4862 ( .A(n4835), .B(n4836), .Z(n4679) );
  AND U4863 ( .A(n4837), .B(n4838), .Z(n4836) );
  XNOR U4864 ( .A(n4835), .B(n4646), .Z(n4838) );
  XOR U4865 ( .A(n4839), .B(n4764), .Z(n4646) );
  XNOR U4866 ( .A(n4840), .B(n4771), .Z(n4764) );
  XOR U4867 ( .A(n4760), .B(n4759), .Z(n4771) );
  XNOR U4868 ( .A(n4841), .B(n4756), .Z(n4759) );
  XOR U4869 ( .A(n4842), .B(n4843), .Z(n4756) );
  AND U4870 ( .A(n4844), .B(n4845), .Z(n4843) );
  XOR U4871 ( .A(n4842), .B(n4846), .Z(n4844) );
  XNOR U4872 ( .A(n4847), .B(n4848), .Z(n4841) );
  NOR U4873 ( .A(n4849), .B(n4850), .Z(n4848) );
  XNOR U4874 ( .A(n4847), .B(n4851), .Z(n4849) );
  XOR U4875 ( .A(n4852), .B(n4853), .Z(n4760) );
  NOR U4876 ( .A(n4854), .B(n4855), .Z(n4853) );
  XNOR U4877 ( .A(n4852), .B(n4856), .Z(n4854) );
  XNOR U4878 ( .A(n4770), .B(n4761), .Z(n4840) );
  XOR U4879 ( .A(n4857), .B(n4858), .Z(n4761) );
  NOR U4880 ( .A(n4859), .B(n4860), .Z(n4858) );
  XNOR U4881 ( .A(n4857), .B(n4861), .Z(n4859) );
  XOR U4882 ( .A(n4862), .B(n4776), .Z(n4770) );
  XNOR U4883 ( .A(n4863), .B(n4864), .Z(n4776) );
  NOR U4884 ( .A(n4865), .B(n4866), .Z(n4864) );
  XNOR U4885 ( .A(n4863), .B(n4867), .Z(n4865) );
  XNOR U4886 ( .A(n4775), .B(n4767), .Z(n4862) );
  XOR U4887 ( .A(n4868), .B(n4869), .Z(n4767) );
  AND U4888 ( .A(n4870), .B(n4871), .Z(n4869) );
  XOR U4889 ( .A(n4868), .B(n4872), .Z(n4870) );
  XNOR U4890 ( .A(n4873), .B(n4772), .Z(n4775) );
  XOR U4891 ( .A(n4874), .B(n4875), .Z(n4772) );
  AND U4892 ( .A(n4876), .B(n4877), .Z(n4875) );
  XOR U4893 ( .A(n4874), .B(n4878), .Z(n4876) );
  XNOR U4894 ( .A(n4879), .B(n4880), .Z(n4873) );
  NOR U4895 ( .A(n4881), .B(n4882), .Z(n4880) );
  XOR U4896 ( .A(n4879), .B(n4883), .Z(n4881) );
  XOR U4897 ( .A(n4765), .B(n4777), .Z(n4839) );
  AND U4898 ( .A(n4685), .B(n4884), .Z(n4777) );
  IV U4899 ( .A(n4664), .Z(n4685) );
  XNOR U4900 ( .A(n4783), .B(n4782), .Z(n4765) );
  XNOR U4901 ( .A(n4885), .B(n4788), .Z(n4782) );
  XOR U4902 ( .A(n4886), .B(n4887), .Z(n4788) );
  NOR U4903 ( .A(n4888), .B(n4889), .Z(n4887) );
  XNOR U4904 ( .A(n4886), .B(n4890), .Z(n4888) );
  XNOR U4905 ( .A(n4787), .B(n4779), .Z(n4885) );
  XOR U4906 ( .A(n4891), .B(n4892), .Z(n4779) );
  AND U4907 ( .A(n4893), .B(n4894), .Z(n4892) );
  XNOR U4908 ( .A(n4891), .B(n4895), .Z(n4893) );
  XNOR U4909 ( .A(n4896), .B(n4784), .Z(n4787) );
  XOR U4910 ( .A(n4897), .B(n4898), .Z(n4784) );
  AND U4911 ( .A(n4899), .B(n4900), .Z(n4898) );
  XOR U4912 ( .A(n4897), .B(n4901), .Z(n4899) );
  XNOR U4913 ( .A(n4902), .B(n4903), .Z(n4896) );
  NOR U4914 ( .A(n4904), .B(n4905), .Z(n4903) );
  XOR U4915 ( .A(n4902), .B(n4906), .Z(n4904) );
  XOR U4916 ( .A(n4793), .B(n4792), .Z(n4783) );
  XNOR U4917 ( .A(n4907), .B(n4789), .Z(n4792) );
  XOR U4918 ( .A(n4908), .B(n4909), .Z(n4789) );
  AND U4919 ( .A(n4910), .B(n4911), .Z(n4909) );
  XOR U4920 ( .A(n4908), .B(n4912), .Z(n4910) );
  XNOR U4921 ( .A(n4913), .B(n4914), .Z(n4907) );
  NOR U4922 ( .A(n4915), .B(n4916), .Z(n4914) );
  XNOR U4923 ( .A(n4913), .B(n4917), .Z(n4915) );
  XOR U4924 ( .A(n4918), .B(n4919), .Z(n4793) );
  NOR U4925 ( .A(n4920), .B(n4921), .Z(n4919) );
  XNOR U4926 ( .A(n4918), .B(n4922), .Z(n4920) );
  XNOR U4927 ( .A(n4923), .B(n4835), .Z(n4837) );
  IV U4928 ( .A(n4466), .Z(n4923) );
  XOR U4929 ( .A(n4924), .B(n4823), .Z(n4466) );
  XOR U4930 ( .A(n4801), .B(n4800), .Z(n4823) );
  XNOR U4931 ( .A(n4925), .B(n4806), .Z(n4800) );
  XOR U4932 ( .A(n4926), .B(n4927), .Z(n4806) );
  NOR U4933 ( .A(n4928), .B(n4929), .Z(n4927) );
  XNOR U4934 ( .A(n4926), .B(n4930), .Z(n4928) );
  XNOR U4935 ( .A(n4805), .B(n4797), .Z(n4925) );
  XOR U4936 ( .A(n4931), .B(n4932), .Z(n4797) );
  AND U4937 ( .A(n4933), .B(n4934), .Z(n4932) );
  XNOR U4938 ( .A(n4931), .B(n4935), .Z(n4933) );
  XNOR U4939 ( .A(n4936), .B(n4802), .Z(n4805) );
  XOR U4940 ( .A(n4937), .B(n4938), .Z(n4802) );
  AND U4941 ( .A(n4939), .B(n4940), .Z(n4938) );
  XOR U4942 ( .A(n4937), .B(n4941), .Z(n4939) );
  XNOR U4943 ( .A(n4942), .B(n4943), .Z(n4936) );
  NOR U4944 ( .A(n4944), .B(n4945), .Z(n4943) );
  XOR U4945 ( .A(n4942), .B(n4946), .Z(n4944) );
  XOR U4946 ( .A(n4811), .B(n4810), .Z(n4801) );
  XNOR U4947 ( .A(n4947), .B(n4807), .Z(n4810) );
  XOR U4948 ( .A(n4948), .B(n4949), .Z(n4807) );
  AND U4949 ( .A(n4950), .B(n4951), .Z(n4949) );
  XOR U4950 ( .A(n4948), .B(n4952), .Z(n4950) );
  XNOR U4951 ( .A(n4953), .B(n4954), .Z(n4947) );
  NOR U4952 ( .A(n4955), .B(n4956), .Z(n4954) );
  XNOR U4953 ( .A(n4953), .B(n4957), .Z(n4955) );
  XOR U4954 ( .A(n4958), .B(n4959), .Z(n4811) );
  NOR U4955 ( .A(n4960), .B(n4961), .Z(n4959) );
  XNOR U4956 ( .A(n4958), .B(n4962), .Z(n4960) );
  XNOR U4957 ( .A(n4822), .B(n4812), .Z(n4924) );
  AND U4958 ( .A(n4683), .B(n4963), .Z(n4812) );
  XNOR U4959 ( .A(n4964), .B(n4829), .Z(n4822) );
  XOR U4960 ( .A(n4818), .B(n4817), .Z(n4829) );
  XNOR U4961 ( .A(n4965), .B(n4814), .Z(n4817) );
  XOR U4962 ( .A(n4966), .B(n4967), .Z(n4814) );
  AND U4963 ( .A(n4968), .B(n4969), .Z(n4967) );
  XOR U4964 ( .A(n4966), .B(n4970), .Z(n4968) );
  XNOR U4965 ( .A(n4971), .B(n4972), .Z(n4965) );
  NOR U4966 ( .A(n4973), .B(n4974), .Z(n4972) );
  XNOR U4967 ( .A(n4971), .B(n4975), .Z(n4973) );
  XOR U4968 ( .A(n4976), .B(n4977), .Z(n4818) );
  NOR U4969 ( .A(n4978), .B(n4979), .Z(n4977) );
  XNOR U4970 ( .A(n4976), .B(n4980), .Z(n4978) );
  XNOR U4971 ( .A(n4828), .B(n4819), .Z(n4964) );
  XOR U4972 ( .A(n4981), .B(n4982), .Z(n4819) );
  NOR U4973 ( .A(n4983), .B(n4984), .Z(n4982) );
  XNOR U4974 ( .A(n4981), .B(n4985), .Z(n4983) );
  XOR U4975 ( .A(n4986), .B(n4834), .Z(n4828) );
  XNOR U4976 ( .A(n4987), .B(n4988), .Z(n4834) );
  NOR U4977 ( .A(n4989), .B(n4990), .Z(n4988) );
  XNOR U4978 ( .A(n4987), .B(n4991), .Z(n4989) );
  XNOR U4979 ( .A(n4833), .B(n4825), .Z(n4986) );
  XOR U4980 ( .A(n4992), .B(n4993), .Z(n4825) );
  AND U4981 ( .A(n4994), .B(n4995), .Z(n4993) );
  XOR U4982 ( .A(n4992), .B(n4996), .Z(n4994) );
  XNOR U4983 ( .A(n4997), .B(n4830), .Z(n4833) );
  XOR U4984 ( .A(n4998), .B(n4999), .Z(n4830) );
  AND U4985 ( .A(n5000), .B(n5001), .Z(n4999) );
  XOR U4986 ( .A(n4998), .B(n5002), .Z(n5000) );
  XNOR U4987 ( .A(n5003), .B(n5004), .Z(n4997) );
  NOR U4988 ( .A(n5005), .B(n5006), .Z(n5004) );
  XOR U4989 ( .A(n5003), .B(n5007), .Z(n5005) );
  AND U4990 ( .A(n4683), .B(n4664), .Z(n4835) );
  XNOR U4991 ( .A(n5008), .B(n4884), .Z(n4664) );
  XOR U4992 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(
        p_input[256]), .Z(n4884) );
  XOR U4993 ( .A(n4861), .B(n4860), .Z(n5008) );
  XOR U4994 ( .A(n5009), .B(n4872), .Z(n4860) );
  XOR U4995 ( .A(n4846), .B(n4845), .Z(n4872) );
  XNOR U4996 ( .A(n5010), .B(n4851), .Z(n4845) );
  XOR U4997 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .B(
        p_input[280]), .Z(n4851) );
  XOR U4998 ( .A(n4842), .B(n4850), .Z(n5010) );
  XOR U4999 ( .A(n5011), .B(n4847), .Z(n4850) );
  XOR U5000 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .B(
        p_input[278]), .Z(n4847) );
  XOR U5001 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .B(n2951), 
        .Z(n5011) );
  XNOR U5002 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .B(n3316), 
        .Z(n4842) );
  XNOR U5003 ( .A(n4856), .B(n4855), .Z(n4846) );
  XOR U5004 ( .A(n5012), .B(n4852), .Z(n4855) );
  XOR U5005 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .B(
        p_input[275]), .Z(n4852) );
  XOR U5006 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .B(n2953), 
        .Z(n5012) );
  XOR U5007 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .B(
        p_input[277]), .Z(n4856) );
  XNOR U5008 ( .A(n4871), .B(n4857), .Z(n5009) );
  XNOR U5009 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(n3318), 
        .Z(n4857) );
  XNOR U5010 ( .A(n5013), .B(n4878), .Z(n4871) );
  XNOR U5011 ( .A(n4867), .B(n4866), .Z(n4878) );
  XOR U5012 ( .A(n5014), .B(n4863), .Z(n4866) );
  XNOR U5013 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .B(n3321), 
        .Z(n4863) );
  XOR U5014 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .B(n2957), 
        .Z(n5014) );
  XOR U5015 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .B(
        p_input[284]), .Z(n4867) );
  XNOR U5016 ( .A(n4877), .B(n4868), .Z(n5013) );
  XNOR U5017 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .B(n3322), 
        .Z(n4868) );
  XOR U5018 ( .A(n5015), .B(n4883), .Z(n4877) );
  XNOR U5019 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .B(
        p_input[287]), .Z(n4883) );
  XOR U5020 ( .A(n4874), .B(n4882), .Z(n5015) );
  XOR U5021 ( .A(n5016), .B(n4879), .Z(n4882) );
  XOR U5022 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .B(
        p_input[285]), .Z(n4879) );
  XOR U5023 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .B(n4385), 
        .Z(n5016) );
  XNOR U5024 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .B(n3325), 
        .Z(n4874) );
  XNOR U5025 ( .A(n4895), .B(n4894), .Z(n4861) );
  XNOR U5026 ( .A(n5017), .B(n4901), .Z(n4894) );
  XNOR U5027 ( .A(n4890), .B(n4889), .Z(n4901) );
  XOR U5028 ( .A(n5018), .B(n4886), .Z(n4889) );
  XNOR U5029 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n3328), 
        .Z(n4886) );
  XOR U5030 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(n2963), 
        .Z(n5018) );
  XOR U5031 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(
        p_input[269]), .Z(n4890) );
  XNOR U5032 ( .A(n4900), .B(n4891), .Z(n5017) );
  XOR U5033 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .B(
        p_input[258]), .Z(n4891) );
  XOR U5034 ( .A(n5019), .B(n4906), .Z(n4900) );
  XNOR U5035 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .B(
        p_input[272]), .Z(n4906) );
  XOR U5036 ( .A(n4897), .B(n4905), .Z(n5019) );
  XOR U5037 ( .A(n5020), .B(n4902), .Z(n4905) );
  XOR U5038 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(
        p_input[270]), .Z(n4902) );
  XOR U5039 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(n2967), 
        .Z(n5020) );
  XNOR U5040 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(n3331), 
        .Z(n4897) );
  XNOR U5041 ( .A(n4912), .B(n4911), .Z(n4895) );
  XNOR U5042 ( .A(n5021), .B(n4917), .Z(n4911) );
  XNOR U5043 ( .A(n228), .B(p_input[265]), .Z(n4917) );
  IV U5044 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .Z(n228) );
  XOR U5045 ( .A(n4908), .B(n4916), .Z(n5021) );
  XOR U5046 ( .A(n5022), .B(n4913), .Z(n4916) );
  XNOR U5047 ( .A(n388), .B(p_input[263]), .Z(n4913) );
  IV U5048 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .Z(n388) );
  XOR U5049 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .B(n4392), 
        .Z(n5022) );
  XOR U5050 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .B(
        p_input[259]), .Z(n4908) );
  XNOR U5051 ( .A(n4922), .B(n4921), .Z(n4912) );
  XOR U5052 ( .A(n5023), .B(n4918), .Z(n4921) );
  XOR U5053 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(
        p_input[260]), .Z(n4918) );
  XOR U5054 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(n4394), 
        .Z(n5023) );
  XOR U5055 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .B(
        p_input[262]), .Z(n4922) );
  XOR U5056 ( .A(n5024), .B(n4985), .Z(n4683) );
  XNOR U5057 ( .A(n4935), .B(n4934), .Z(n4985) );
  XNOR U5058 ( .A(n5025), .B(n4941), .Z(n4934) );
  XNOR U5059 ( .A(n4930), .B(n4929), .Z(n4941) );
  XOR U5060 ( .A(n5026), .B(n4926), .Z(n4929) );
  XNOR U5061 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n3328), .Z(n4926) );
  IV U5062 ( .A(p_input[267]), .Z(n3328) );
  XOR U5063 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n2963), .Z(n5026) );
  IV U5064 ( .A(p_input[268]), .Z(n2963) );
  XOR U5065 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[269]), .Z(n4930)
         );
  XNOR U5066 ( .A(n4940), .B(n4931), .Z(n5025) );
  XOR U5067 ( .A(\knn_comb_/min_val_out[0][2] ), .B(p_input[258]), .Z(n4931)
         );
  XOR U5068 ( .A(n5027), .B(n4946), .Z(n4940) );
  XNOR U5069 ( .A(\knn_comb_/min_val_out[0][16] ), .B(p_input[272]), .Z(n4946)
         );
  XOR U5070 ( .A(n4937), .B(n4945), .Z(n5027) );
  XOR U5071 ( .A(n5028), .B(n4942), .Z(n4945) );
  XOR U5072 ( .A(\knn_comb_/min_val_out[0][14] ), .B(p_input[270]), .Z(n4942)
         );
  XOR U5073 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n2967), .Z(n5028) );
  IV U5074 ( .A(p_input[271]), .Z(n2967) );
  XNOR U5075 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n3331), .Z(n4937) );
  IV U5076 ( .A(p_input[266]), .Z(n3331) );
  XNOR U5077 ( .A(n4952), .B(n4951), .Z(n4935) );
  XNOR U5078 ( .A(n5029), .B(n4957), .Z(n4951) );
  XNOR U5079 ( .A(n227), .B(p_input[265]), .Z(n4957) );
  IV U5080 ( .A(\knn_comb_/min_val_out[0][9] ), .Z(n227) );
  XOR U5081 ( .A(n4948), .B(n4956), .Z(n5029) );
  XOR U5082 ( .A(n5030), .B(n4953), .Z(n4956) );
  XNOR U5083 ( .A(n387), .B(p_input[263]), .Z(n4953) );
  IV U5084 ( .A(\knn_comb_/min_val_out[0][7] ), .Z(n387) );
  XOR U5085 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n4392), .Z(n5030) );
  IV U5086 ( .A(p_input[264]), .Z(n4392) );
  XOR U5087 ( .A(\knn_comb_/min_val_out[0][3] ), .B(p_input[259]), .Z(n4948)
         );
  XNOR U5088 ( .A(n4962), .B(n4961), .Z(n4952) );
  XOR U5089 ( .A(n5031), .B(n4958), .Z(n4961) );
  XOR U5090 ( .A(\knn_comb_/min_val_out[0][4] ), .B(p_input[260]), .Z(n4958)
         );
  XOR U5091 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n4394), .Z(n5031) );
  IV U5092 ( .A(p_input[261]), .Z(n4394) );
  XOR U5093 ( .A(\knn_comb_/min_val_out[0][6] ), .B(p_input[262]), .Z(n4962)
         );
  XOR U5094 ( .A(n4984), .B(n4963), .Z(n5024) );
  XOR U5095 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[256]), .Z(n4963)
         );
  XOR U5096 ( .A(n5032), .B(n4996), .Z(n4984) );
  XOR U5097 ( .A(n4970), .B(n4969), .Z(n4996) );
  XNOR U5098 ( .A(n5033), .B(n4975), .Z(n4969) );
  XOR U5099 ( .A(\knn_comb_/min_val_out[0][24] ), .B(p_input[280]), .Z(n4975)
         );
  XOR U5100 ( .A(n4966), .B(n4974), .Z(n5033) );
  XOR U5101 ( .A(n5034), .B(n4971), .Z(n4974) );
  XOR U5102 ( .A(\knn_comb_/min_val_out[0][22] ), .B(p_input[278]), .Z(n4971)
         );
  XOR U5103 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n2951), .Z(n5034) );
  IV U5104 ( .A(p_input[279]), .Z(n2951) );
  XNOR U5105 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n3316), .Z(n4966) );
  IV U5106 ( .A(p_input[274]), .Z(n3316) );
  XNOR U5107 ( .A(n4980), .B(n4979), .Z(n4970) );
  XOR U5108 ( .A(n5035), .B(n4976), .Z(n4979) );
  XOR U5109 ( .A(\knn_comb_/min_val_out[0][19] ), .B(p_input[275]), .Z(n4976)
         );
  XOR U5110 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n2953), .Z(n5035) );
  IV U5111 ( .A(p_input[276]), .Z(n2953) );
  XOR U5112 ( .A(\knn_comb_/min_val_out[0][21] ), .B(p_input[277]), .Z(n4980)
         );
  XNOR U5113 ( .A(n4995), .B(n4981), .Z(n5032) );
  XNOR U5114 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n3318), .Z(n4981) );
  IV U5115 ( .A(p_input[257]), .Z(n3318) );
  XNOR U5116 ( .A(n5036), .B(n5002), .Z(n4995) );
  XNOR U5117 ( .A(n4991), .B(n4990), .Z(n5002) );
  XOR U5118 ( .A(n5037), .B(n4987), .Z(n4990) );
  XNOR U5119 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n3321), .Z(n4987) );
  IV U5120 ( .A(p_input[282]), .Z(n3321) );
  XOR U5121 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n2957), .Z(n5037) );
  IV U5122 ( .A(p_input[283]), .Z(n2957) );
  XOR U5123 ( .A(\knn_comb_/min_val_out[0][28] ), .B(p_input[284]), .Z(n4991)
         );
  XNOR U5124 ( .A(n5001), .B(n4992), .Z(n5036) );
  XNOR U5125 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n3322), .Z(n4992) );
  IV U5126 ( .A(p_input[273]), .Z(n3322) );
  XOR U5127 ( .A(n5038), .B(n5007), .Z(n5001) );
  XNOR U5128 ( .A(\knn_comb_/min_val_out[0][31] ), .B(p_input[287]), .Z(n5007)
         );
  XOR U5129 ( .A(n4998), .B(n5006), .Z(n5038) );
  XOR U5130 ( .A(n5039), .B(n5003), .Z(n5006) );
  XOR U5131 ( .A(\knn_comb_/min_val_out[0][29] ), .B(p_input[285]), .Z(n5003)
         );
  XOR U5132 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n4385), .Z(n5039) );
  IV U5133 ( .A(p_input[286]), .Z(n4385) );
  XNOR U5134 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n3325), .Z(n4998) );
  IV U5135 ( .A(p_input[281]), .Z(n3325) );
endmodule

