
module psi_BMR_b10000_n3 ( p_input, o );
  input [29999:0] p_input;
  output [9999:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582,
         n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592,
         n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602,
         n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612,
         n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622,
         n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632,
         n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642,
         n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652,
         n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662,
         n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672,
         n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682,
         n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692,
         n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702,
         n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712,
         n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722,
         n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732,
         n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742,
         n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752,
         n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762,
         n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772,
         n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782,
         n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792,
         n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802,
         n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812,
         n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822,
         n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832,
         n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842,
         n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852,
         n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862,
         n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872,
         n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882,
         n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892,
         n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902,
         n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912,
         n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922,
         n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932,
         n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942,
         n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952,
         n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962,
         n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972,
         n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982,
         n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992,
         n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002,
         n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012,
         n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022,
         n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032,
         n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042,
         n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052,
         n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062,
         n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072,
         n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082,
         n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092,
         n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102,
         n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112,
         n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122,
         n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132,
         n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142,
         n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152,
         n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162,
         n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172,
         n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182,
         n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192,
         n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202,
         n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212,
         n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222,
         n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232,
         n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242,
         n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252,
         n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262,
         n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272,
         n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282,
         n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292,
         n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302,
         n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312,
         n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322,
         n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332,
         n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342,
         n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352,
         n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362,
         n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372,
         n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382,
         n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392,
         n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402,
         n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412,
         n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422,
         n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432,
         n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442,
         n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452,
         n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462,
         n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472,
         n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482,
         n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492,
         n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502,
         n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512,
         n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522,
         n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532,
         n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542,
         n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552,
         n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562,
         n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572,
         n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582,
         n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592,
         n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602,
         n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612,
         n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622,
         n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632,
         n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642,
         n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652,
         n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662,
         n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672,
         n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682,
         n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692,
         n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702,
         n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712,
         n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722,
         n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732,
         n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742,
         n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752,
         n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762,
         n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772,
         n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782,
         n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792,
         n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802,
         n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812,
         n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822,
         n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832,
         n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842,
         n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852,
         n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862,
         n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872,
         n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882,
         n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892,
         n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902,
         n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912,
         n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922,
         n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932,
         n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942,
         n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952,
         n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962,
         n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972,
         n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982,
         n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992,
         n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000;

  AND U1 ( .A(n1), .B(p_input[9]), .Z(o[9]) );
  AND U2 ( .A(p_input[20009]), .B(p_input[10009]), .Z(n1) );
  AND U3 ( .A(n2), .B(p_input[99]), .Z(o[99]) );
  AND U4 ( .A(p_input[20099]), .B(p_input[10099]), .Z(n2) );
  AND U5 ( .A(n3), .B(p_input[999]), .Z(o[999]) );
  AND U6 ( .A(p_input[20999]), .B(p_input[10999]), .Z(n3) );
  AND U7 ( .A(n4), .B(p_input[9999]), .Z(o[9999]) );
  AND U8 ( .A(p_input[29999]), .B(p_input[19999]), .Z(n4) );
  AND U9 ( .A(n5), .B(p_input[9998]), .Z(o[9998]) );
  AND U10 ( .A(p_input[29998]), .B(p_input[19998]), .Z(n5) );
  AND U11 ( .A(n6), .B(p_input[9997]), .Z(o[9997]) );
  AND U12 ( .A(p_input[29997]), .B(p_input[19997]), .Z(n6) );
  AND U13 ( .A(n7), .B(p_input[9996]), .Z(o[9996]) );
  AND U14 ( .A(p_input[29996]), .B(p_input[19996]), .Z(n7) );
  AND U15 ( .A(n8), .B(p_input[9995]), .Z(o[9995]) );
  AND U16 ( .A(p_input[29995]), .B(p_input[19995]), .Z(n8) );
  AND U17 ( .A(n9), .B(p_input[9994]), .Z(o[9994]) );
  AND U18 ( .A(p_input[29994]), .B(p_input[19994]), .Z(n9) );
  AND U19 ( .A(n10), .B(p_input[9993]), .Z(o[9993]) );
  AND U20 ( .A(p_input[29993]), .B(p_input[19993]), .Z(n10) );
  AND U21 ( .A(n11), .B(p_input[9992]), .Z(o[9992]) );
  AND U22 ( .A(p_input[29992]), .B(p_input[19992]), .Z(n11) );
  AND U23 ( .A(n12), .B(p_input[9991]), .Z(o[9991]) );
  AND U24 ( .A(p_input[29991]), .B(p_input[19991]), .Z(n12) );
  AND U25 ( .A(n13), .B(p_input[9990]), .Z(o[9990]) );
  AND U26 ( .A(p_input[29990]), .B(p_input[19990]), .Z(n13) );
  AND U27 ( .A(n14), .B(p_input[998]), .Z(o[998]) );
  AND U28 ( .A(p_input[20998]), .B(p_input[10998]), .Z(n14) );
  AND U29 ( .A(n15), .B(p_input[9989]), .Z(o[9989]) );
  AND U30 ( .A(p_input[29989]), .B(p_input[19989]), .Z(n15) );
  AND U31 ( .A(n16), .B(p_input[9988]), .Z(o[9988]) );
  AND U32 ( .A(p_input[29988]), .B(p_input[19988]), .Z(n16) );
  AND U33 ( .A(n17), .B(p_input[9987]), .Z(o[9987]) );
  AND U34 ( .A(p_input[29987]), .B(p_input[19987]), .Z(n17) );
  AND U35 ( .A(n18), .B(p_input[9986]), .Z(o[9986]) );
  AND U36 ( .A(p_input[29986]), .B(p_input[19986]), .Z(n18) );
  AND U37 ( .A(n19), .B(p_input[9985]), .Z(o[9985]) );
  AND U38 ( .A(p_input[29985]), .B(p_input[19985]), .Z(n19) );
  AND U39 ( .A(n20), .B(p_input[9984]), .Z(o[9984]) );
  AND U40 ( .A(p_input[29984]), .B(p_input[19984]), .Z(n20) );
  AND U41 ( .A(n21), .B(p_input[9983]), .Z(o[9983]) );
  AND U42 ( .A(p_input[29983]), .B(p_input[19983]), .Z(n21) );
  AND U43 ( .A(n22), .B(p_input[9982]), .Z(o[9982]) );
  AND U44 ( .A(p_input[29982]), .B(p_input[19982]), .Z(n22) );
  AND U45 ( .A(n23), .B(p_input[9981]), .Z(o[9981]) );
  AND U46 ( .A(p_input[29981]), .B(p_input[19981]), .Z(n23) );
  AND U47 ( .A(n24), .B(p_input[9980]), .Z(o[9980]) );
  AND U48 ( .A(p_input[29980]), .B(p_input[19980]), .Z(n24) );
  AND U49 ( .A(n25), .B(p_input[997]), .Z(o[997]) );
  AND U50 ( .A(p_input[20997]), .B(p_input[10997]), .Z(n25) );
  AND U51 ( .A(n26), .B(p_input[9979]), .Z(o[9979]) );
  AND U52 ( .A(p_input[29979]), .B(p_input[19979]), .Z(n26) );
  AND U53 ( .A(n27), .B(p_input[9978]), .Z(o[9978]) );
  AND U54 ( .A(p_input[29978]), .B(p_input[19978]), .Z(n27) );
  AND U55 ( .A(n28), .B(p_input[9977]), .Z(o[9977]) );
  AND U56 ( .A(p_input[29977]), .B(p_input[19977]), .Z(n28) );
  AND U57 ( .A(n29), .B(p_input[9976]), .Z(o[9976]) );
  AND U58 ( .A(p_input[29976]), .B(p_input[19976]), .Z(n29) );
  AND U59 ( .A(n30), .B(p_input[9975]), .Z(o[9975]) );
  AND U60 ( .A(p_input[29975]), .B(p_input[19975]), .Z(n30) );
  AND U61 ( .A(n31), .B(p_input[9974]), .Z(o[9974]) );
  AND U62 ( .A(p_input[29974]), .B(p_input[19974]), .Z(n31) );
  AND U63 ( .A(n32), .B(p_input[9973]), .Z(o[9973]) );
  AND U64 ( .A(p_input[29973]), .B(p_input[19973]), .Z(n32) );
  AND U65 ( .A(n33), .B(p_input[9972]), .Z(o[9972]) );
  AND U66 ( .A(p_input[29972]), .B(p_input[19972]), .Z(n33) );
  AND U67 ( .A(n34), .B(p_input[9971]), .Z(o[9971]) );
  AND U68 ( .A(p_input[29971]), .B(p_input[19971]), .Z(n34) );
  AND U69 ( .A(n35), .B(p_input[9970]), .Z(o[9970]) );
  AND U70 ( .A(p_input[29970]), .B(p_input[19970]), .Z(n35) );
  AND U71 ( .A(n36), .B(p_input[996]), .Z(o[996]) );
  AND U72 ( .A(p_input[20996]), .B(p_input[10996]), .Z(n36) );
  AND U73 ( .A(n37), .B(p_input[9969]), .Z(o[9969]) );
  AND U74 ( .A(p_input[29969]), .B(p_input[19969]), .Z(n37) );
  AND U75 ( .A(n38), .B(p_input[9968]), .Z(o[9968]) );
  AND U76 ( .A(p_input[29968]), .B(p_input[19968]), .Z(n38) );
  AND U77 ( .A(n39), .B(p_input[9967]), .Z(o[9967]) );
  AND U78 ( .A(p_input[29967]), .B(p_input[19967]), .Z(n39) );
  AND U79 ( .A(n40), .B(p_input[9966]), .Z(o[9966]) );
  AND U80 ( .A(p_input[29966]), .B(p_input[19966]), .Z(n40) );
  AND U81 ( .A(n41), .B(p_input[9965]), .Z(o[9965]) );
  AND U82 ( .A(p_input[29965]), .B(p_input[19965]), .Z(n41) );
  AND U83 ( .A(n42), .B(p_input[9964]), .Z(o[9964]) );
  AND U84 ( .A(p_input[29964]), .B(p_input[19964]), .Z(n42) );
  AND U85 ( .A(n43), .B(p_input[9963]), .Z(o[9963]) );
  AND U86 ( .A(p_input[29963]), .B(p_input[19963]), .Z(n43) );
  AND U87 ( .A(n44), .B(p_input[9962]), .Z(o[9962]) );
  AND U88 ( .A(p_input[29962]), .B(p_input[19962]), .Z(n44) );
  AND U89 ( .A(n45), .B(p_input[9961]), .Z(o[9961]) );
  AND U90 ( .A(p_input[29961]), .B(p_input[19961]), .Z(n45) );
  AND U91 ( .A(n46), .B(p_input[9960]), .Z(o[9960]) );
  AND U92 ( .A(p_input[29960]), .B(p_input[19960]), .Z(n46) );
  AND U93 ( .A(n47), .B(p_input[995]), .Z(o[995]) );
  AND U94 ( .A(p_input[20995]), .B(p_input[10995]), .Z(n47) );
  AND U95 ( .A(n48), .B(p_input[9959]), .Z(o[9959]) );
  AND U96 ( .A(p_input[29959]), .B(p_input[19959]), .Z(n48) );
  AND U97 ( .A(n49), .B(p_input[9958]), .Z(o[9958]) );
  AND U98 ( .A(p_input[29958]), .B(p_input[19958]), .Z(n49) );
  AND U99 ( .A(n50), .B(p_input[9957]), .Z(o[9957]) );
  AND U100 ( .A(p_input[29957]), .B(p_input[19957]), .Z(n50) );
  AND U101 ( .A(n51), .B(p_input[9956]), .Z(o[9956]) );
  AND U102 ( .A(p_input[29956]), .B(p_input[19956]), .Z(n51) );
  AND U103 ( .A(n52), .B(p_input[9955]), .Z(o[9955]) );
  AND U104 ( .A(p_input[29955]), .B(p_input[19955]), .Z(n52) );
  AND U105 ( .A(n53), .B(p_input[9954]), .Z(o[9954]) );
  AND U106 ( .A(p_input[29954]), .B(p_input[19954]), .Z(n53) );
  AND U107 ( .A(n54), .B(p_input[9953]), .Z(o[9953]) );
  AND U108 ( .A(p_input[29953]), .B(p_input[19953]), .Z(n54) );
  AND U109 ( .A(n55), .B(p_input[9952]), .Z(o[9952]) );
  AND U110 ( .A(p_input[29952]), .B(p_input[19952]), .Z(n55) );
  AND U111 ( .A(n56), .B(p_input[9951]), .Z(o[9951]) );
  AND U112 ( .A(p_input[29951]), .B(p_input[19951]), .Z(n56) );
  AND U113 ( .A(n57), .B(p_input[9950]), .Z(o[9950]) );
  AND U114 ( .A(p_input[29950]), .B(p_input[19950]), .Z(n57) );
  AND U115 ( .A(n58), .B(p_input[994]), .Z(o[994]) );
  AND U116 ( .A(p_input[20994]), .B(p_input[10994]), .Z(n58) );
  AND U117 ( .A(n59), .B(p_input[9949]), .Z(o[9949]) );
  AND U118 ( .A(p_input[29949]), .B(p_input[19949]), .Z(n59) );
  AND U119 ( .A(n60), .B(p_input[9948]), .Z(o[9948]) );
  AND U120 ( .A(p_input[29948]), .B(p_input[19948]), .Z(n60) );
  AND U121 ( .A(n61), .B(p_input[9947]), .Z(o[9947]) );
  AND U122 ( .A(p_input[29947]), .B(p_input[19947]), .Z(n61) );
  AND U123 ( .A(n62), .B(p_input[9946]), .Z(o[9946]) );
  AND U124 ( .A(p_input[29946]), .B(p_input[19946]), .Z(n62) );
  AND U125 ( .A(n63), .B(p_input[9945]), .Z(o[9945]) );
  AND U126 ( .A(p_input[29945]), .B(p_input[19945]), .Z(n63) );
  AND U127 ( .A(n64), .B(p_input[9944]), .Z(o[9944]) );
  AND U128 ( .A(p_input[29944]), .B(p_input[19944]), .Z(n64) );
  AND U129 ( .A(n65), .B(p_input[9943]), .Z(o[9943]) );
  AND U130 ( .A(p_input[29943]), .B(p_input[19943]), .Z(n65) );
  AND U131 ( .A(n66), .B(p_input[9942]), .Z(o[9942]) );
  AND U132 ( .A(p_input[29942]), .B(p_input[19942]), .Z(n66) );
  AND U133 ( .A(n67), .B(p_input[9941]), .Z(o[9941]) );
  AND U134 ( .A(p_input[29941]), .B(p_input[19941]), .Z(n67) );
  AND U135 ( .A(n68), .B(p_input[9940]), .Z(o[9940]) );
  AND U136 ( .A(p_input[29940]), .B(p_input[19940]), .Z(n68) );
  AND U137 ( .A(n69), .B(p_input[993]), .Z(o[993]) );
  AND U138 ( .A(p_input[20993]), .B(p_input[10993]), .Z(n69) );
  AND U139 ( .A(n70), .B(p_input[9939]), .Z(o[9939]) );
  AND U140 ( .A(p_input[29939]), .B(p_input[19939]), .Z(n70) );
  AND U141 ( .A(n71), .B(p_input[9938]), .Z(o[9938]) );
  AND U142 ( .A(p_input[29938]), .B(p_input[19938]), .Z(n71) );
  AND U143 ( .A(n72), .B(p_input[9937]), .Z(o[9937]) );
  AND U144 ( .A(p_input[29937]), .B(p_input[19937]), .Z(n72) );
  AND U145 ( .A(n73), .B(p_input[9936]), .Z(o[9936]) );
  AND U146 ( .A(p_input[29936]), .B(p_input[19936]), .Z(n73) );
  AND U147 ( .A(n74), .B(p_input[9935]), .Z(o[9935]) );
  AND U148 ( .A(p_input[29935]), .B(p_input[19935]), .Z(n74) );
  AND U149 ( .A(n75), .B(p_input[9934]), .Z(o[9934]) );
  AND U150 ( .A(p_input[29934]), .B(p_input[19934]), .Z(n75) );
  AND U151 ( .A(n76), .B(p_input[9933]), .Z(o[9933]) );
  AND U152 ( .A(p_input[29933]), .B(p_input[19933]), .Z(n76) );
  AND U153 ( .A(n77), .B(p_input[9932]), .Z(o[9932]) );
  AND U154 ( .A(p_input[29932]), .B(p_input[19932]), .Z(n77) );
  AND U155 ( .A(n78), .B(p_input[9931]), .Z(o[9931]) );
  AND U156 ( .A(p_input[29931]), .B(p_input[19931]), .Z(n78) );
  AND U157 ( .A(n79), .B(p_input[9930]), .Z(o[9930]) );
  AND U158 ( .A(p_input[29930]), .B(p_input[19930]), .Z(n79) );
  AND U159 ( .A(n80), .B(p_input[992]), .Z(o[992]) );
  AND U160 ( .A(p_input[20992]), .B(p_input[10992]), .Z(n80) );
  AND U161 ( .A(n81), .B(p_input[9929]), .Z(o[9929]) );
  AND U162 ( .A(p_input[29929]), .B(p_input[19929]), .Z(n81) );
  AND U163 ( .A(n82), .B(p_input[9928]), .Z(o[9928]) );
  AND U164 ( .A(p_input[29928]), .B(p_input[19928]), .Z(n82) );
  AND U165 ( .A(n83), .B(p_input[9927]), .Z(o[9927]) );
  AND U166 ( .A(p_input[29927]), .B(p_input[19927]), .Z(n83) );
  AND U167 ( .A(n84), .B(p_input[9926]), .Z(o[9926]) );
  AND U168 ( .A(p_input[29926]), .B(p_input[19926]), .Z(n84) );
  AND U169 ( .A(n85), .B(p_input[9925]), .Z(o[9925]) );
  AND U170 ( .A(p_input[29925]), .B(p_input[19925]), .Z(n85) );
  AND U171 ( .A(n86), .B(p_input[9924]), .Z(o[9924]) );
  AND U172 ( .A(p_input[29924]), .B(p_input[19924]), .Z(n86) );
  AND U173 ( .A(n87), .B(p_input[9923]), .Z(o[9923]) );
  AND U174 ( .A(p_input[29923]), .B(p_input[19923]), .Z(n87) );
  AND U175 ( .A(n88), .B(p_input[9922]), .Z(o[9922]) );
  AND U176 ( .A(p_input[29922]), .B(p_input[19922]), .Z(n88) );
  AND U177 ( .A(n89), .B(p_input[9921]), .Z(o[9921]) );
  AND U178 ( .A(p_input[29921]), .B(p_input[19921]), .Z(n89) );
  AND U179 ( .A(n90), .B(p_input[9920]), .Z(o[9920]) );
  AND U180 ( .A(p_input[29920]), .B(p_input[19920]), .Z(n90) );
  AND U181 ( .A(n91), .B(p_input[991]), .Z(o[991]) );
  AND U182 ( .A(p_input[20991]), .B(p_input[10991]), .Z(n91) );
  AND U183 ( .A(n92), .B(p_input[9919]), .Z(o[9919]) );
  AND U184 ( .A(p_input[29919]), .B(p_input[19919]), .Z(n92) );
  AND U185 ( .A(n93), .B(p_input[9918]), .Z(o[9918]) );
  AND U186 ( .A(p_input[29918]), .B(p_input[19918]), .Z(n93) );
  AND U187 ( .A(n94), .B(p_input[9917]), .Z(o[9917]) );
  AND U188 ( .A(p_input[29917]), .B(p_input[19917]), .Z(n94) );
  AND U189 ( .A(n95), .B(p_input[9916]), .Z(o[9916]) );
  AND U190 ( .A(p_input[29916]), .B(p_input[19916]), .Z(n95) );
  AND U191 ( .A(n96), .B(p_input[9915]), .Z(o[9915]) );
  AND U192 ( .A(p_input[29915]), .B(p_input[19915]), .Z(n96) );
  AND U193 ( .A(n97), .B(p_input[9914]), .Z(o[9914]) );
  AND U194 ( .A(p_input[29914]), .B(p_input[19914]), .Z(n97) );
  AND U195 ( .A(n98), .B(p_input[9913]), .Z(o[9913]) );
  AND U196 ( .A(p_input[29913]), .B(p_input[19913]), .Z(n98) );
  AND U197 ( .A(n99), .B(p_input[9912]), .Z(o[9912]) );
  AND U198 ( .A(p_input[29912]), .B(p_input[19912]), .Z(n99) );
  AND U199 ( .A(n100), .B(p_input[9911]), .Z(o[9911]) );
  AND U200 ( .A(p_input[29911]), .B(p_input[19911]), .Z(n100) );
  AND U201 ( .A(n101), .B(p_input[9910]), .Z(o[9910]) );
  AND U202 ( .A(p_input[29910]), .B(p_input[19910]), .Z(n101) );
  AND U203 ( .A(n102), .B(p_input[990]), .Z(o[990]) );
  AND U204 ( .A(p_input[20990]), .B(p_input[10990]), .Z(n102) );
  AND U205 ( .A(n103), .B(p_input[9909]), .Z(o[9909]) );
  AND U206 ( .A(p_input[29909]), .B(p_input[19909]), .Z(n103) );
  AND U207 ( .A(n104), .B(p_input[9908]), .Z(o[9908]) );
  AND U208 ( .A(p_input[29908]), .B(p_input[19908]), .Z(n104) );
  AND U209 ( .A(n105), .B(p_input[9907]), .Z(o[9907]) );
  AND U210 ( .A(p_input[29907]), .B(p_input[19907]), .Z(n105) );
  AND U211 ( .A(n106), .B(p_input[9906]), .Z(o[9906]) );
  AND U212 ( .A(p_input[29906]), .B(p_input[19906]), .Z(n106) );
  AND U213 ( .A(n107), .B(p_input[9905]), .Z(o[9905]) );
  AND U214 ( .A(p_input[29905]), .B(p_input[19905]), .Z(n107) );
  AND U215 ( .A(n108), .B(p_input[9904]), .Z(o[9904]) );
  AND U216 ( .A(p_input[29904]), .B(p_input[19904]), .Z(n108) );
  AND U217 ( .A(n109), .B(p_input[9903]), .Z(o[9903]) );
  AND U218 ( .A(p_input[29903]), .B(p_input[19903]), .Z(n109) );
  AND U219 ( .A(n110), .B(p_input[9902]), .Z(o[9902]) );
  AND U220 ( .A(p_input[29902]), .B(p_input[19902]), .Z(n110) );
  AND U221 ( .A(n111), .B(p_input[9901]), .Z(o[9901]) );
  AND U222 ( .A(p_input[29901]), .B(p_input[19901]), .Z(n111) );
  AND U223 ( .A(n112), .B(p_input[9900]), .Z(o[9900]) );
  AND U224 ( .A(p_input[29900]), .B(p_input[19900]), .Z(n112) );
  AND U225 ( .A(n113), .B(p_input[98]), .Z(o[98]) );
  AND U226 ( .A(p_input[20098]), .B(p_input[10098]), .Z(n113) );
  AND U227 ( .A(n114), .B(p_input[989]), .Z(o[989]) );
  AND U228 ( .A(p_input[20989]), .B(p_input[10989]), .Z(n114) );
  AND U229 ( .A(n115), .B(p_input[9899]), .Z(o[9899]) );
  AND U230 ( .A(p_input[29899]), .B(p_input[19899]), .Z(n115) );
  AND U231 ( .A(n116), .B(p_input[9898]), .Z(o[9898]) );
  AND U232 ( .A(p_input[29898]), .B(p_input[19898]), .Z(n116) );
  AND U233 ( .A(n117), .B(p_input[9897]), .Z(o[9897]) );
  AND U234 ( .A(p_input[29897]), .B(p_input[19897]), .Z(n117) );
  AND U235 ( .A(n118), .B(p_input[9896]), .Z(o[9896]) );
  AND U236 ( .A(p_input[29896]), .B(p_input[19896]), .Z(n118) );
  AND U237 ( .A(n119), .B(p_input[9895]), .Z(o[9895]) );
  AND U238 ( .A(p_input[29895]), .B(p_input[19895]), .Z(n119) );
  AND U239 ( .A(n120), .B(p_input[9894]), .Z(o[9894]) );
  AND U240 ( .A(p_input[29894]), .B(p_input[19894]), .Z(n120) );
  AND U241 ( .A(n121), .B(p_input[9893]), .Z(o[9893]) );
  AND U242 ( .A(p_input[29893]), .B(p_input[19893]), .Z(n121) );
  AND U243 ( .A(n122), .B(p_input[9892]), .Z(o[9892]) );
  AND U244 ( .A(p_input[29892]), .B(p_input[19892]), .Z(n122) );
  AND U245 ( .A(n123), .B(p_input[9891]), .Z(o[9891]) );
  AND U246 ( .A(p_input[29891]), .B(p_input[19891]), .Z(n123) );
  AND U247 ( .A(n124), .B(p_input[9890]), .Z(o[9890]) );
  AND U248 ( .A(p_input[29890]), .B(p_input[19890]), .Z(n124) );
  AND U249 ( .A(n125), .B(p_input[988]), .Z(o[988]) );
  AND U250 ( .A(p_input[20988]), .B(p_input[10988]), .Z(n125) );
  AND U251 ( .A(n126), .B(p_input[9889]), .Z(o[9889]) );
  AND U252 ( .A(p_input[29889]), .B(p_input[19889]), .Z(n126) );
  AND U253 ( .A(n127), .B(p_input[9888]), .Z(o[9888]) );
  AND U254 ( .A(p_input[29888]), .B(p_input[19888]), .Z(n127) );
  AND U255 ( .A(n128), .B(p_input[9887]), .Z(o[9887]) );
  AND U256 ( .A(p_input[29887]), .B(p_input[19887]), .Z(n128) );
  AND U257 ( .A(n129), .B(p_input[9886]), .Z(o[9886]) );
  AND U258 ( .A(p_input[29886]), .B(p_input[19886]), .Z(n129) );
  AND U259 ( .A(n130), .B(p_input[9885]), .Z(o[9885]) );
  AND U260 ( .A(p_input[29885]), .B(p_input[19885]), .Z(n130) );
  AND U261 ( .A(n131), .B(p_input[9884]), .Z(o[9884]) );
  AND U262 ( .A(p_input[29884]), .B(p_input[19884]), .Z(n131) );
  AND U263 ( .A(n132), .B(p_input[9883]), .Z(o[9883]) );
  AND U264 ( .A(p_input[29883]), .B(p_input[19883]), .Z(n132) );
  AND U265 ( .A(n133), .B(p_input[9882]), .Z(o[9882]) );
  AND U266 ( .A(p_input[29882]), .B(p_input[19882]), .Z(n133) );
  AND U267 ( .A(n134), .B(p_input[9881]), .Z(o[9881]) );
  AND U268 ( .A(p_input[29881]), .B(p_input[19881]), .Z(n134) );
  AND U269 ( .A(n135), .B(p_input[9880]), .Z(o[9880]) );
  AND U270 ( .A(p_input[29880]), .B(p_input[19880]), .Z(n135) );
  AND U271 ( .A(n136), .B(p_input[987]), .Z(o[987]) );
  AND U272 ( .A(p_input[20987]), .B(p_input[10987]), .Z(n136) );
  AND U273 ( .A(n137), .B(p_input[9879]), .Z(o[9879]) );
  AND U274 ( .A(p_input[29879]), .B(p_input[19879]), .Z(n137) );
  AND U275 ( .A(n138), .B(p_input[9878]), .Z(o[9878]) );
  AND U276 ( .A(p_input[29878]), .B(p_input[19878]), .Z(n138) );
  AND U277 ( .A(n139), .B(p_input[9877]), .Z(o[9877]) );
  AND U278 ( .A(p_input[29877]), .B(p_input[19877]), .Z(n139) );
  AND U279 ( .A(n140), .B(p_input[9876]), .Z(o[9876]) );
  AND U280 ( .A(p_input[29876]), .B(p_input[19876]), .Z(n140) );
  AND U281 ( .A(n141), .B(p_input[9875]), .Z(o[9875]) );
  AND U282 ( .A(p_input[29875]), .B(p_input[19875]), .Z(n141) );
  AND U283 ( .A(n142), .B(p_input[9874]), .Z(o[9874]) );
  AND U284 ( .A(p_input[29874]), .B(p_input[19874]), .Z(n142) );
  AND U285 ( .A(n143), .B(p_input[9873]), .Z(o[9873]) );
  AND U286 ( .A(p_input[29873]), .B(p_input[19873]), .Z(n143) );
  AND U287 ( .A(n144), .B(p_input[9872]), .Z(o[9872]) );
  AND U288 ( .A(p_input[29872]), .B(p_input[19872]), .Z(n144) );
  AND U289 ( .A(n145), .B(p_input[9871]), .Z(o[9871]) );
  AND U290 ( .A(p_input[29871]), .B(p_input[19871]), .Z(n145) );
  AND U291 ( .A(n146), .B(p_input[9870]), .Z(o[9870]) );
  AND U292 ( .A(p_input[29870]), .B(p_input[19870]), .Z(n146) );
  AND U293 ( .A(n147), .B(p_input[986]), .Z(o[986]) );
  AND U294 ( .A(p_input[20986]), .B(p_input[10986]), .Z(n147) );
  AND U295 ( .A(n148), .B(p_input[9869]), .Z(o[9869]) );
  AND U296 ( .A(p_input[29869]), .B(p_input[19869]), .Z(n148) );
  AND U297 ( .A(n149), .B(p_input[9868]), .Z(o[9868]) );
  AND U298 ( .A(p_input[29868]), .B(p_input[19868]), .Z(n149) );
  AND U299 ( .A(n150), .B(p_input[9867]), .Z(o[9867]) );
  AND U300 ( .A(p_input[29867]), .B(p_input[19867]), .Z(n150) );
  AND U301 ( .A(n151), .B(p_input[9866]), .Z(o[9866]) );
  AND U302 ( .A(p_input[29866]), .B(p_input[19866]), .Z(n151) );
  AND U303 ( .A(n152), .B(p_input[9865]), .Z(o[9865]) );
  AND U304 ( .A(p_input[29865]), .B(p_input[19865]), .Z(n152) );
  AND U305 ( .A(n153), .B(p_input[9864]), .Z(o[9864]) );
  AND U306 ( .A(p_input[29864]), .B(p_input[19864]), .Z(n153) );
  AND U307 ( .A(n154), .B(p_input[9863]), .Z(o[9863]) );
  AND U308 ( .A(p_input[29863]), .B(p_input[19863]), .Z(n154) );
  AND U309 ( .A(n155), .B(p_input[9862]), .Z(o[9862]) );
  AND U310 ( .A(p_input[29862]), .B(p_input[19862]), .Z(n155) );
  AND U311 ( .A(n156), .B(p_input[9861]), .Z(o[9861]) );
  AND U312 ( .A(p_input[29861]), .B(p_input[19861]), .Z(n156) );
  AND U313 ( .A(n157), .B(p_input[9860]), .Z(o[9860]) );
  AND U314 ( .A(p_input[29860]), .B(p_input[19860]), .Z(n157) );
  AND U315 ( .A(n158), .B(p_input[985]), .Z(o[985]) );
  AND U316 ( .A(p_input[20985]), .B(p_input[10985]), .Z(n158) );
  AND U317 ( .A(n159), .B(p_input[9859]), .Z(o[9859]) );
  AND U318 ( .A(p_input[29859]), .B(p_input[19859]), .Z(n159) );
  AND U319 ( .A(n160), .B(p_input[9858]), .Z(o[9858]) );
  AND U320 ( .A(p_input[29858]), .B(p_input[19858]), .Z(n160) );
  AND U321 ( .A(n161), .B(p_input[9857]), .Z(o[9857]) );
  AND U322 ( .A(p_input[29857]), .B(p_input[19857]), .Z(n161) );
  AND U323 ( .A(n162), .B(p_input[9856]), .Z(o[9856]) );
  AND U324 ( .A(p_input[29856]), .B(p_input[19856]), .Z(n162) );
  AND U325 ( .A(n163), .B(p_input[9855]), .Z(o[9855]) );
  AND U326 ( .A(p_input[29855]), .B(p_input[19855]), .Z(n163) );
  AND U327 ( .A(n164), .B(p_input[9854]), .Z(o[9854]) );
  AND U328 ( .A(p_input[29854]), .B(p_input[19854]), .Z(n164) );
  AND U329 ( .A(n165), .B(p_input[9853]), .Z(o[9853]) );
  AND U330 ( .A(p_input[29853]), .B(p_input[19853]), .Z(n165) );
  AND U331 ( .A(n166), .B(p_input[9852]), .Z(o[9852]) );
  AND U332 ( .A(p_input[29852]), .B(p_input[19852]), .Z(n166) );
  AND U333 ( .A(n167), .B(p_input[9851]), .Z(o[9851]) );
  AND U334 ( .A(p_input[29851]), .B(p_input[19851]), .Z(n167) );
  AND U335 ( .A(n168), .B(p_input[9850]), .Z(o[9850]) );
  AND U336 ( .A(p_input[29850]), .B(p_input[19850]), .Z(n168) );
  AND U337 ( .A(n169), .B(p_input[984]), .Z(o[984]) );
  AND U338 ( .A(p_input[20984]), .B(p_input[10984]), .Z(n169) );
  AND U339 ( .A(n170), .B(p_input[9849]), .Z(o[9849]) );
  AND U340 ( .A(p_input[29849]), .B(p_input[19849]), .Z(n170) );
  AND U341 ( .A(n171), .B(p_input[9848]), .Z(o[9848]) );
  AND U342 ( .A(p_input[29848]), .B(p_input[19848]), .Z(n171) );
  AND U343 ( .A(n172), .B(p_input[9847]), .Z(o[9847]) );
  AND U344 ( .A(p_input[29847]), .B(p_input[19847]), .Z(n172) );
  AND U345 ( .A(n173), .B(p_input[9846]), .Z(o[9846]) );
  AND U346 ( .A(p_input[29846]), .B(p_input[19846]), .Z(n173) );
  AND U347 ( .A(n174), .B(p_input[9845]), .Z(o[9845]) );
  AND U348 ( .A(p_input[29845]), .B(p_input[19845]), .Z(n174) );
  AND U349 ( .A(n175), .B(p_input[9844]), .Z(o[9844]) );
  AND U350 ( .A(p_input[29844]), .B(p_input[19844]), .Z(n175) );
  AND U351 ( .A(n176), .B(p_input[9843]), .Z(o[9843]) );
  AND U352 ( .A(p_input[29843]), .B(p_input[19843]), .Z(n176) );
  AND U353 ( .A(n177), .B(p_input[9842]), .Z(o[9842]) );
  AND U354 ( .A(p_input[29842]), .B(p_input[19842]), .Z(n177) );
  AND U355 ( .A(n178), .B(p_input[9841]), .Z(o[9841]) );
  AND U356 ( .A(p_input[29841]), .B(p_input[19841]), .Z(n178) );
  AND U357 ( .A(n179), .B(p_input[9840]), .Z(o[9840]) );
  AND U358 ( .A(p_input[29840]), .B(p_input[19840]), .Z(n179) );
  AND U359 ( .A(n180), .B(p_input[983]), .Z(o[983]) );
  AND U360 ( .A(p_input[20983]), .B(p_input[10983]), .Z(n180) );
  AND U361 ( .A(n181), .B(p_input[9839]), .Z(o[9839]) );
  AND U362 ( .A(p_input[29839]), .B(p_input[19839]), .Z(n181) );
  AND U363 ( .A(n182), .B(p_input[9838]), .Z(o[9838]) );
  AND U364 ( .A(p_input[29838]), .B(p_input[19838]), .Z(n182) );
  AND U365 ( .A(n183), .B(p_input[9837]), .Z(o[9837]) );
  AND U366 ( .A(p_input[29837]), .B(p_input[19837]), .Z(n183) );
  AND U367 ( .A(n184), .B(p_input[9836]), .Z(o[9836]) );
  AND U368 ( .A(p_input[29836]), .B(p_input[19836]), .Z(n184) );
  AND U369 ( .A(n185), .B(p_input[9835]), .Z(o[9835]) );
  AND U370 ( .A(p_input[29835]), .B(p_input[19835]), .Z(n185) );
  AND U371 ( .A(n186), .B(p_input[9834]), .Z(o[9834]) );
  AND U372 ( .A(p_input[29834]), .B(p_input[19834]), .Z(n186) );
  AND U373 ( .A(n187), .B(p_input[9833]), .Z(o[9833]) );
  AND U374 ( .A(p_input[29833]), .B(p_input[19833]), .Z(n187) );
  AND U375 ( .A(n188), .B(p_input[9832]), .Z(o[9832]) );
  AND U376 ( .A(p_input[29832]), .B(p_input[19832]), .Z(n188) );
  AND U377 ( .A(n189), .B(p_input[9831]), .Z(o[9831]) );
  AND U378 ( .A(p_input[29831]), .B(p_input[19831]), .Z(n189) );
  AND U379 ( .A(n190), .B(p_input[9830]), .Z(o[9830]) );
  AND U380 ( .A(p_input[29830]), .B(p_input[19830]), .Z(n190) );
  AND U381 ( .A(n191), .B(p_input[982]), .Z(o[982]) );
  AND U382 ( .A(p_input[20982]), .B(p_input[10982]), .Z(n191) );
  AND U383 ( .A(n192), .B(p_input[9829]), .Z(o[9829]) );
  AND U384 ( .A(p_input[29829]), .B(p_input[19829]), .Z(n192) );
  AND U385 ( .A(n193), .B(p_input[9828]), .Z(o[9828]) );
  AND U386 ( .A(p_input[29828]), .B(p_input[19828]), .Z(n193) );
  AND U387 ( .A(n194), .B(p_input[9827]), .Z(o[9827]) );
  AND U388 ( .A(p_input[29827]), .B(p_input[19827]), .Z(n194) );
  AND U389 ( .A(n195), .B(p_input[9826]), .Z(o[9826]) );
  AND U390 ( .A(p_input[29826]), .B(p_input[19826]), .Z(n195) );
  AND U391 ( .A(n196), .B(p_input[9825]), .Z(o[9825]) );
  AND U392 ( .A(p_input[29825]), .B(p_input[19825]), .Z(n196) );
  AND U393 ( .A(n197), .B(p_input[9824]), .Z(o[9824]) );
  AND U394 ( .A(p_input[29824]), .B(p_input[19824]), .Z(n197) );
  AND U395 ( .A(n198), .B(p_input[9823]), .Z(o[9823]) );
  AND U396 ( .A(p_input[29823]), .B(p_input[19823]), .Z(n198) );
  AND U397 ( .A(n199), .B(p_input[9822]), .Z(o[9822]) );
  AND U398 ( .A(p_input[29822]), .B(p_input[19822]), .Z(n199) );
  AND U399 ( .A(n200), .B(p_input[9821]), .Z(o[9821]) );
  AND U400 ( .A(p_input[29821]), .B(p_input[19821]), .Z(n200) );
  AND U401 ( .A(n201), .B(p_input[9820]), .Z(o[9820]) );
  AND U402 ( .A(p_input[29820]), .B(p_input[19820]), .Z(n201) );
  AND U403 ( .A(n202), .B(p_input[981]), .Z(o[981]) );
  AND U404 ( .A(p_input[20981]), .B(p_input[10981]), .Z(n202) );
  AND U405 ( .A(n203), .B(p_input[9819]), .Z(o[9819]) );
  AND U406 ( .A(p_input[29819]), .B(p_input[19819]), .Z(n203) );
  AND U407 ( .A(n204), .B(p_input[9818]), .Z(o[9818]) );
  AND U408 ( .A(p_input[29818]), .B(p_input[19818]), .Z(n204) );
  AND U409 ( .A(n205), .B(p_input[9817]), .Z(o[9817]) );
  AND U410 ( .A(p_input[29817]), .B(p_input[19817]), .Z(n205) );
  AND U411 ( .A(n206), .B(p_input[9816]), .Z(o[9816]) );
  AND U412 ( .A(p_input[29816]), .B(p_input[19816]), .Z(n206) );
  AND U413 ( .A(n207), .B(p_input[9815]), .Z(o[9815]) );
  AND U414 ( .A(p_input[29815]), .B(p_input[19815]), .Z(n207) );
  AND U415 ( .A(n208), .B(p_input[9814]), .Z(o[9814]) );
  AND U416 ( .A(p_input[29814]), .B(p_input[19814]), .Z(n208) );
  AND U417 ( .A(n209), .B(p_input[9813]), .Z(o[9813]) );
  AND U418 ( .A(p_input[29813]), .B(p_input[19813]), .Z(n209) );
  AND U419 ( .A(n210), .B(p_input[9812]), .Z(o[9812]) );
  AND U420 ( .A(p_input[29812]), .B(p_input[19812]), .Z(n210) );
  AND U421 ( .A(n211), .B(p_input[9811]), .Z(o[9811]) );
  AND U422 ( .A(p_input[29811]), .B(p_input[19811]), .Z(n211) );
  AND U423 ( .A(n212), .B(p_input[9810]), .Z(o[9810]) );
  AND U424 ( .A(p_input[29810]), .B(p_input[19810]), .Z(n212) );
  AND U425 ( .A(n213), .B(p_input[980]), .Z(o[980]) );
  AND U426 ( .A(p_input[20980]), .B(p_input[10980]), .Z(n213) );
  AND U427 ( .A(n214), .B(p_input[9809]), .Z(o[9809]) );
  AND U428 ( .A(p_input[29809]), .B(p_input[19809]), .Z(n214) );
  AND U429 ( .A(n215), .B(p_input[9808]), .Z(o[9808]) );
  AND U430 ( .A(p_input[29808]), .B(p_input[19808]), .Z(n215) );
  AND U431 ( .A(n216), .B(p_input[9807]), .Z(o[9807]) );
  AND U432 ( .A(p_input[29807]), .B(p_input[19807]), .Z(n216) );
  AND U433 ( .A(n217), .B(p_input[9806]), .Z(o[9806]) );
  AND U434 ( .A(p_input[29806]), .B(p_input[19806]), .Z(n217) );
  AND U435 ( .A(n218), .B(p_input[9805]), .Z(o[9805]) );
  AND U436 ( .A(p_input[29805]), .B(p_input[19805]), .Z(n218) );
  AND U437 ( .A(n219), .B(p_input[9804]), .Z(o[9804]) );
  AND U438 ( .A(p_input[29804]), .B(p_input[19804]), .Z(n219) );
  AND U439 ( .A(n220), .B(p_input[9803]), .Z(o[9803]) );
  AND U440 ( .A(p_input[29803]), .B(p_input[19803]), .Z(n220) );
  AND U441 ( .A(n221), .B(p_input[9802]), .Z(o[9802]) );
  AND U442 ( .A(p_input[29802]), .B(p_input[19802]), .Z(n221) );
  AND U443 ( .A(n222), .B(p_input[9801]), .Z(o[9801]) );
  AND U444 ( .A(p_input[29801]), .B(p_input[19801]), .Z(n222) );
  AND U445 ( .A(n223), .B(p_input[9800]), .Z(o[9800]) );
  AND U446 ( .A(p_input[29800]), .B(p_input[19800]), .Z(n223) );
  AND U447 ( .A(n224), .B(p_input[97]), .Z(o[97]) );
  AND U448 ( .A(p_input[20097]), .B(p_input[10097]), .Z(n224) );
  AND U449 ( .A(n225), .B(p_input[979]), .Z(o[979]) );
  AND U450 ( .A(p_input[20979]), .B(p_input[10979]), .Z(n225) );
  AND U451 ( .A(n226), .B(p_input[9799]), .Z(o[9799]) );
  AND U452 ( .A(p_input[29799]), .B(p_input[19799]), .Z(n226) );
  AND U453 ( .A(n227), .B(p_input[9798]), .Z(o[9798]) );
  AND U454 ( .A(p_input[29798]), .B(p_input[19798]), .Z(n227) );
  AND U455 ( .A(n228), .B(p_input[9797]), .Z(o[9797]) );
  AND U456 ( .A(p_input[29797]), .B(p_input[19797]), .Z(n228) );
  AND U457 ( .A(n229), .B(p_input[9796]), .Z(o[9796]) );
  AND U458 ( .A(p_input[29796]), .B(p_input[19796]), .Z(n229) );
  AND U459 ( .A(n230), .B(p_input[9795]), .Z(o[9795]) );
  AND U460 ( .A(p_input[29795]), .B(p_input[19795]), .Z(n230) );
  AND U461 ( .A(n231), .B(p_input[9794]), .Z(o[9794]) );
  AND U462 ( .A(p_input[29794]), .B(p_input[19794]), .Z(n231) );
  AND U463 ( .A(n232), .B(p_input[9793]), .Z(o[9793]) );
  AND U464 ( .A(p_input[29793]), .B(p_input[19793]), .Z(n232) );
  AND U465 ( .A(n233), .B(p_input[9792]), .Z(o[9792]) );
  AND U466 ( .A(p_input[29792]), .B(p_input[19792]), .Z(n233) );
  AND U467 ( .A(n234), .B(p_input[9791]), .Z(o[9791]) );
  AND U468 ( .A(p_input[29791]), .B(p_input[19791]), .Z(n234) );
  AND U469 ( .A(n235), .B(p_input[9790]), .Z(o[9790]) );
  AND U470 ( .A(p_input[29790]), .B(p_input[19790]), .Z(n235) );
  AND U471 ( .A(n236), .B(p_input[978]), .Z(o[978]) );
  AND U472 ( .A(p_input[20978]), .B(p_input[10978]), .Z(n236) );
  AND U473 ( .A(n237), .B(p_input[9789]), .Z(o[9789]) );
  AND U474 ( .A(p_input[29789]), .B(p_input[19789]), .Z(n237) );
  AND U475 ( .A(n238), .B(p_input[9788]), .Z(o[9788]) );
  AND U476 ( .A(p_input[29788]), .B(p_input[19788]), .Z(n238) );
  AND U477 ( .A(n239), .B(p_input[9787]), .Z(o[9787]) );
  AND U478 ( .A(p_input[29787]), .B(p_input[19787]), .Z(n239) );
  AND U479 ( .A(n240), .B(p_input[9786]), .Z(o[9786]) );
  AND U480 ( .A(p_input[29786]), .B(p_input[19786]), .Z(n240) );
  AND U481 ( .A(n241), .B(p_input[9785]), .Z(o[9785]) );
  AND U482 ( .A(p_input[29785]), .B(p_input[19785]), .Z(n241) );
  AND U483 ( .A(n242), .B(p_input[9784]), .Z(o[9784]) );
  AND U484 ( .A(p_input[29784]), .B(p_input[19784]), .Z(n242) );
  AND U485 ( .A(n243), .B(p_input[9783]), .Z(o[9783]) );
  AND U486 ( .A(p_input[29783]), .B(p_input[19783]), .Z(n243) );
  AND U487 ( .A(n244), .B(p_input[9782]), .Z(o[9782]) );
  AND U488 ( .A(p_input[29782]), .B(p_input[19782]), .Z(n244) );
  AND U489 ( .A(n245), .B(p_input[9781]), .Z(o[9781]) );
  AND U490 ( .A(p_input[29781]), .B(p_input[19781]), .Z(n245) );
  AND U491 ( .A(n246), .B(p_input[9780]), .Z(o[9780]) );
  AND U492 ( .A(p_input[29780]), .B(p_input[19780]), .Z(n246) );
  AND U493 ( .A(n247), .B(p_input[977]), .Z(o[977]) );
  AND U494 ( .A(p_input[20977]), .B(p_input[10977]), .Z(n247) );
  AND U495 ( .A(n248), .B(p_input[9779]), .Z(o[9779]) );
  AND U496 ( .A(p_input[29779]), .B(p_input[19779]), .Z(n248) );
  AND U497 ( .A(n249), .B(p_input[9778]), .Z(o[9778]) );
  AND U498 ( .A(p_input[29778]), .B(p_input[19778]), .Z(n249) );
  AND U499 ( .A(n250), .B(p_input[9777]), .Z(o[9777]) );
  AND U500 ( .A(p_input[29777]), .B(p_input[19777]), .Z(n250) );
  AND U501 ( .A(n251), .B(p_input[9776]), .Z(o[9776]) );
  AND U502 ( .A(p_input[29776]), .B(p_input[19776]), .Z(n251) );
  AND U503 ( .A(n252), .B(p_input[9775]), .Z(o[9775]) );
  AND U504 ( .A(p_input[29775]), .B(p_input[19775]), .Z(n252) );
  AND U505 ( .A(n253), .B(p_input[9774]), .Z(o[9774]) );
  AND U506 ( .A(p_input[29774]), .B(p_input[19774]), .Z(n253) );
  AND U507 ( .A(n254), .B(p_input[9773]), .Z(o[9773]) );
  AND U508 ( .A(p_input[29773]), .B(p_input[19773]), .Z(n254) );
  AND U509 ( .A(n255), .B(p_input[9772]), .Z(o[9772]) );
  AND U510 ( .A(p_input[29772]), .B(p_input[19772]), .Z(n255) );
  AND U511 ( .A(n256), .B(p_input[9771]), .Z(o[9771]) );
  AND U512 ( .A(p_input[29771]), .B(p_input[19771]), .Z(n256) );
  AND U513 ( .A(n257), .B(p_input[9770]), .Z(o[9770]) );
  AND U514 ( .A(p_input[29770]), .B(p_input[19770]), .Z(n257) );
  AND U515 ( .A(n258), .B(p_input[976]), .Z(o[976]) );
  AND U516 ( .A(p_input[20976]), .B(p_input[10976]), .Z(n258) );
  AND U517 ( .A(n259), .B(p_input[9769]), .Z(o[9769]) );
  AND U518 ( .A(p_input[29769]), .B(p_input[19769]), .Z(n259) );
  AND U519 ( .A(n260), .B(p_input[9768]), .Z(o[9768]) );
  AND U520 ( .A(p_input[29768]), .B(p_input[19768]), .Z(n260) );
  AND U521 ( .A(n261), .B(p_input[9767]), .Z(o[9767]) );
  AND U522 ( .A(p_input[29767]), .B(p_input[19767]), .Z(n261) );
  AND U523 ( .A(n262), .B(p_input[9766]), .Z(o[9766]) );
  AND U524 ( .A(p_input[29766]), .B(p_input[19766]), .Z(n262) );
  AND U525 ( .A(n263), .B(p_input[9765]), .Z(o[9765]) );
  AND U526 ( .A(p_input[29765]), .B(p_input[19765]), .Z(n263) );
  AND U527 ( .A(n264), .B(p_input[9764]), .Z(o[9764]) );
  AND U528 ( .A(p_input[29764]), .B(p_input[19764]), .Z(n264) );
  AND U529 ( .A(n265), .B(p_input[9763]), .Z(o[9763]) );
  AND U530 ( .A(p_input[29763]), .B(p_input[19763]), .Z(n265) );
  AND U531 ( .A(n266), .B(p_input[9762]), .Z(o[9762]) );
  AND U532 ( .A(p_input[29762]), .B(p_input[19762]), .Z(n266) );
  AND U533 ( .A(n267), .B(p_input[9761]), .Z(o[9761]) );
  AND U534 ( .A(p_input[29761]), .B(p_input[19761]), .Z(n267) );
  AND U535 ( .A(n268), .B(p_input[9760]), .Z(o[9760]) );
  AND U536 ( .A(p_input[29760]), .B(p_input[19760]), .Z(n268) );
  AND U537 ( .A(n269), .B(p_input[975]), .Z(o[975]) );
  AND U538 ( .A(p_input[20975]), .B(p_input[10975]), .Z(n269) );
  AND U539 ( .A(n270), .B(p_input[9759]), .Z(o[9759]) );
  AND U540 ( .A(p_input[29759]), .B(p_input[19759]), .Z(n270) );
  AND U541 ( .A(n271), .B(p_input[9758]), .Z(o[9758]) );
  AND U542 ( .A(p_input[29758]), .B(p_input[19758]), .Z(n271) );
  AND U543 ( .A(n272), .B(p_input[9757]), .Z(o[9757]) );
  AND U544 ( .A(p_input[29757]), .B(p_input[19757]), .Z(n272) );
  AND U545 ( .A(n273), .B(p_input[9756]), .Z(o[9756]) );
  AND U546 ( .A(p_input[29756]), .B(p_input[19756]), .Z(n273) );
  AND U547 ( .A(n274), .B(p_input[9755]), .Z(o[9755]) );
  AND U548 ( .A(p_input[29755]), .B(p_input[19755]), .Z(n274) );
  AND U549 ( .A(n275), .B(p_input[9754]), .Z(o[9754]) );
  AND U550 ( .A(p_input[29754]), .B(p_input[19754]), .Z(n275) );
  AND U551 ( .A(n276), .B(p_input[9753]), .Z(o[9753]) );
  AND U552 ( .A(p_input[29753]), .B(p_input[19753]), .Z(n276) );
  AND U553 ( .A(n277), .B(p_input[9752]), .Z(o[9752]) );
  AND U554 ( .A(p_input[29752]), .B(p_input[19752]), .Z(n277) );
  AND U555 ( .A(n278), .B(p_input[9751]), .Z(o[9751]) );
  AND U556 ( .A(p_input[29751]), .B(p_input[19751]), .Z(n278) );
  AND U557 ( .A(n279), .B(p_input[9750]), .Z(o[9750]) );
  AND U558 ( .A(p_input[29750]), .B(p_input[19750]), .Z(n279) );
  AND U559 ( .A(n280), .B(p_input[974]), .Z(o[974]) );
  AND U560 ( .A(p_input[20974]), .B(p_input[10974]), .Z(n280) );
  AND U561 ( .A(n281), .B(p_input[9749]), .Z(o[9749]) );
  AND U562 ( .A(p_input[29749]), .B(p_input[19749]), .Z(n281) );
  AND U563 ( .A(n282), .B(p_input[9748]), .Z(o[9748]) );
  AND U564 ( .A(p_input[29748]), .B(p_input[19748]), .Z(n282) );
  AND U565 ( .A(n283), .B(p_input[9747]), .Z(o[9747]) );
  AND U566 ( .A(p_input[29747]), .B(p_input[19747]), .Z(n283) );
  AND U567 ( .A(n284), .B(p_input[9746]), .Z(o[9746]) );
  AND U568 ( .A(p_input[29746]), .B(p_input[19746]), .Z(n284) );
  AND U569 ( .A(n285), .B(p_input[9745]), .Z(o[9745]) );
  AND U570 ( .A(p_input[29745]), .B(p_input[19745]), .Z(n285) );
  AND U571 ( .A(n286), .B(p_input[9744]), .Z(o[9744]) );
  AND U572 ( .A(p_input[29744]), .B(p_input[19744]), .Z(n286) );
  AND U573 ( .A(n287), .B(p_input[9743]), .Z(o[9743]) );
  AND U574 ( .A(p_input[29743]), .B(p_input[19743]), .Z(n287) );
  AND U575 ( .A(n288), .B(p_input[9742]), .Z(o[9742]) );
  AND U576 ( .A(p_input[29742]), .B(p_input[19742]), .Z(n288) );
  AND U577 ( .A(n289), .B(p_input[9741]), .Z(o[9741]) );
  AND U578 ( .A(p_input[29741]), .B(p_input[19741]), .Z(n289) );
  AND U579 ( .A(n290), .B(p_input[9740]), .Z(o[9740]) );
  AND U580 ( .A(p_input[29740]), .B(p_input[19740]), .Z(n290) );
  AND U581 ( .A(n291), .B(p_input[973]), .Z(o[973]) );
  AND U582 ( .A(p_input[20973]), .B(p_input[10973]), .Z(n291) );
  AND U583 ( .A(n292), .B(p_input[9739]), .Z(o[9739]) );
  AND U584 ( .A(p_input[29739]), .B(p_input[19739]), .Z(n292) );
  AND U585 ( .A(n293), .B(p_input[9738]), .Z(o[9738]) );
  AND U586 ( .A(p_input[29738]), .B(p_input[19738]), .Z(n293) );
  AND U587 ( .A(n294), .B(p_input[9737]), .Z(o[9737]) );
  AND U588 ( .A(p_input[29737]), .B(p_input[19737]), .Z(n294) );
  AND U589 ( .A(n295), .B(p_input[9736]), .Z(o[9736]) );
  AND U590 ( .A(p_input[29736]), .B(p_input[19736]), .Z(n295) );
  AND U591 ( .A(n296), .B(p_input[9735]), .Z(o[9735]) );
  AND U592 ( .A(p_input[29735]), .B(p_input[19735]), .Z(n296) );
  AND U593 ( .A(n297), .B(p_input[9734]), .Z(o[9734]) );
  AND U594 ( .A(p_input[29734]), .B(p_input[19734]), .Z(n297) );
  AND U595 ( .A(n298), .B(p_input[9733]), .Z(o[9733]) );
  AND U596 ( .A(p_input[29733]), .B(p_input[19733]), .Z(n298) );
  AND U597 ( .A(n299), .B(p_input[9732]), .Z(o[9732]) );
  AND U598 ( .A(p_input[29732]), .B(p_input[19732]), .Z(n299) );
  AND U599 ( .A(n300), .B(p_input[9731]), .Z(o[9731]) );
  AND U600 ( .A(p_input[29731]), .B(p_input[19731]), .Z(n300) );
  AND U601 ( .A(n301), .B(p_input[9730]), .Z(o[9730]) );
  AND U602 ( .A(p_input[29730]), .B(p_input[19730]), .Z(n301) );
  AND U603 ( .A(n302), .B(p_input[972]), .Z(o[972]) );
  AND U604 ( .A(p_input[20972]), .B(p_input[10972]), .Z(n302) );
  AND U605 ( .A(n303), .B(p_input[9729]), .Z(o[9729]) );
  AND U606 ( .A(p_input[29729]), .B(p_input[19729]), .Z(n303) );
  AND U607 ( .A(n304), .B(p_input[9728]), .Z(o[9728]) );
  AND U608 ( .A(p_input[29728]), .B(p_input[19728]), .Z(n304) );
  AND U609 ( .A(n305), .B(p_input[9727]), .Z(o[9727]) );
  AND U610 ( .A(p_input[29727]), .B(p_input[19727]), .Z(n305) );
  AND U611 ( .A(n306), .B(p_input[9726]), .Z(o[9726]) );
  AND U612 ( .A(p_input[29726]), .B(p_input[19726]), .Z(n306) );
  AND U613 ( .A(n307), .B(p_input[9725]), .Z(o[9725]) );
  AND U614 ( .A(p_input[29725]), .B(p_input[19725]), .Z(n307) );
  AND U615 ( .A(n308), .B(p_input[9724]), .Z(o[9724]) );
  AND U616 ( .A(p_input[29724]), .B(p_input[19724]), .Z(n308) );
  AND U617 ( .A(n309), .B(p_input[9723]), .Z(o[9723]) );
  AND U618 ( .A(p_input[29723]), .B(p_input[19723]), .Z(n309) );
  AND U619 ( .A(n310), .B(p_input[9722]), .Z(o[9722]) );
  AND U620 ( .A(p_input[29722]), .B(p_input[19722]), .Z(n310) );
  AND U621 ( .A(n311), .B(p_input[9721]), .Z(o[9721]) );
  AND U622 ( .A(p_input[29721]), .B(p_input[19721]), .Z(n311) );
  AND U623 ( .A(n312), .B(p_input[9720]), .Z(o[9720]) );
  AND U624 ( .A(p_input[29720]), .B(p_input[19720]), .Z(n312) );
  AND U625 ( .A(n313), .B(p_input[971]), .Z(o[971]) );
  AND U626 ( .A(p_input[20971]), .B(p_input[10971]), .Z(n313) );
  AND U627 ( .A(n314), .B(p_input[9719]), .Z(o[9719]) );
  AND U628 ( .A(p_input[29719]), .B(p_input[19719]), .Z(n314) );
  AND U629 ( .A(n315), .B(p_input[9718]), .Z(o[9718]) );
  AND U630 ( .A(p_input[29718]), .B(p_input[19718]), .Z(n315) );
  AND U631 ( .A(n316), .B(p_input[9717]), .Z(o[9717]) );
  AND U632 ( .A(p_input[29717]), .B(p_input[19717]), .Z(n316) );
  AND U633 ( .A(n317), .B(p_input[9716]), .Z(o[9716]) );
  AND U634 ( .A(p_input[29716]), .B(p_input[19716]), .Z(n317) );
  AND U635 ( .A(n318), .B(p_input[9715]), .Z(o[9715]) );
  AND U636 ( .A(p_input[29715]), .B(p_input[19715]), .Z(n318) );
  AND U637 ( .A(n319), .B(p_input[9714]), .Z(o[9714]) );
  AND U638 ( .A(p_input[29714]), .B(p_input[19714]), .Z(n319) );
  AND U639 ( .A(n320), .B(p_input[9713]), .Z(o[9713]) );
  AND U640 ( .A(p_input[29713]), .B(p_input[19713]), .Z(n320) );
  AND U641 ( .A(n321), .B(p_input[9712]), .Z(o[9712]) );
  AND U642 ( .A(p_input[29712]), .B(p_input[19712]), .Z(n321) );
  AND U643 ( .A(n322), .B(p_input[9711]), .Z(o[9711]) );
  AND U644 ( .A(p_input[29711]), .B(p_input[19711]), .Z(n322) );
  AND U645 ( .A(n323), .B(p_input[9710]), .Z(o[9710]) );
  AND U646 ( .A(p_input[29710]), .B(p_input[19710]), .Z(n323) );
  AND U647 ( .A(n324), .B(p_input[970]), .Z(o[970]) );
  AND U648 ( .A(p_input[20970]), .B(p_input[10970]), .Z(n324) );
  AND U649 ( .A(n325), .B(p_input[9709]), .Z(o[9709]) );
  AND U650 ( .A(p_input[29709]), .B(p_input[19709]), .Z(n325) );
  AND U651 ( .A(n326), .B(p_input[9708]), .Z(o[9708]) );
  AND U652 ( .A(p_input[29708]), .B(p_input[19708]), .Z(n326) );
  AND U653 ( .A(n327), .B(p_input[9707]), .Z(o[9707]) );
  AND U654 ( .A(p_input[29707]), .B(p_input[19707]), .Z(n327) );
  AND U655 ( .A(n328), .B(p_input[9706]), .Z(o[9706]) );
  AND U656 ( .A(p_input[29706]), .B(p_input[19706]), .Z(n328) );
  AND U657 ( .A(n329), .B(p_input[9705]), .Z(o[9705]) );
  AND U658 ( .A(p_input[29705]), .B(p_input[19705]), .Z(n329) );
  AND U659 ( .A(n330), .B(p_input[9704]), .Z(o[9704]) );
  AND U660 ( .A(p_input[29704]), .B(p_input[19704]), .Z(n330) );
  AND U661 ( .A(n331), .B(p_input[9703]), .Z(o[9703]) );
  AND U662 ( .A(p_input[29703]), .B(p_input[19703]), .Z(n331) );
  AND U663 ( .A(n332), .B(p_input[9702]), .Z(o[9702]) );
  AND U664 ( .A(p_input[29702]), .B(p_input[19702]), .Z(n332) );
  AND U665 ( .A(n333), .B(p_input[9701]), .Z(o[9701]) );
  AND U666 ( .A(p_input[29701]), .B(p_input[19701]), .Z(n333) );
  AND U667 ( .A(n334), .B(p_input[9700]), .Z(o[9700]) );
  AND U668 ( .A(p_input[29700]), .B(p_input[19700]), .Z(n334) );
  AND U669 ( .A(n335), .B(p_input[96]), .Z(o[96]) );
  AND U670 ( .A(p_input[20096]), .B(p_input[10096]), .Z(n335) );
  AND U671 ( .A(n336), .B(p_input[969]), .Z(o[969]) );
  AND U672 ( .A(p_input[20969]), .B(p_input[10969]), .Z(n336) );
  AND U673 ( .A(n337), .B(p_input[9699]), .Z(o[9699]) );
  AND U674 ( .A(p_input[29699]), .B(p_input[19699]), .Z(n337) );
  AND U675 ( .A(n338), .B(p_input[9698]), .Z(o[9698]) );
  AND U676 ( .A(p_input[29698]), .B(p_input[19698]), .Z(n338) );
  AND U677 ( .A(n339), .B(p_input[9697]), .Z(o[9697]) );
  AND U678 ( .A(p_input[29697]), .B(p_input[19697]), .Z(n339) );
  AND U679 ( .A(n340), .B(p_input[9696]), .Z(o[9696]) );
  AND U680 ( .A(p_input[29696]), .B(p_input[19696]), .Z(n340) );
  AND U681 ( .A(n341), .B(p_input[9695]), .Z(o[9695]) );
  AND U682 ( .A(p_input[29695]), .B(p_input[19695]), .Z(n341) );
  AND U683 ( .A(n342), .B(p_input[9694]), .Z(o[9694]) );
  AND U684 ( .A(p_input[29694]), .B(p_input[19694]), .Z(n342) );
  AND U685 ( .A(n343), .B(p_input[9693]), .Z(o[9693]) );
  AND U686 ( .A(p_input[29693]), .B(p_input[19693]), .Z(n343) );
  AND U687 ( .A(n344), .B(p_input[9692]), .Z(o[9692]) );
  AND U688 ( .A(p_input[29692]), .B(p_input[19692]), .Z(n344) );
  AND U689 ( .A(n345), .B(p_input[9691]), .Z(o[9691]) );
  AND U690 ( .A(p_input[29691]), .B(p_input[19691]), .Z(n345) );
  AND U691 ( .A(n346), .B(p_input[9690]), .Z(o[9690]) );
  AND U692 ( .A(p_input[29690]), .B(p_input[19690]), .Z(n346) );
  AND U693 ( .A(n347), .B(p_input[968]), .Z(o[968]) );
  AND U694 ( .A(p_input[20968]), .B(p_input[10968]), .Z(n347) );
  AND U695 ( .A(n348), .B(p_input[9689]), .Z(o[9689]) );
  AND U696 ( .A(p_input[29689]), .B(p_input[19689]), .Z(n348) );
  AND U697 ( .A(n349), .B(p_input[9688]), .Z(o[9688]) );
  AND U698 ( .A(p_input[29688]), .B(p_input[19688]), .Z(n349) );
  AND U699 ( .A(n350), .B(p_input[9687]), .Z(o[9687]) );
  AND U700 ( .A(p_input[29687]), .B(p_input[19687]), .Z(n350) );
  AND U701 ( .A(n351), .B(p_input[9686]), .Z(o[9686]) );
  AND U702 ( .A(p_input[29686]), .B(p_input[19686]), .Z(n351) );
  AND U703 ( .A(n352), .B(p_input[9685]), .Z(o[9685]) );
  AND U704 ( .A(p_input[29685]), .B(p_input[19685]), .Z(n352) );
  AND U705 ( .A(n353), .B(p_input[9684]), .Z(o[9684]) );
  AND U706 ( .A(p_input[29684]), .B(p_input[19684]), .Z(n353) );
  AND U707 ( .A(n354), .B(p_input[9683]), .Z(o[9683]) );
  AND U708 ( .A(p_input[29683]), .B(p_input[19683]), .Z(n354) );
  AND U709 ( .A(n355), .B(p_input[9682]), .Z(o[9682]) );
  AND U710 ( .A(p_input[29682]), .B(p_input[19682]), .Z(n355) );
  AND U711 ( .A(n356), .B(p_input[9681]), .Z(o[9681]) );
  AND U712 ( .A(p_input[29681]), .B(p_input[19681]), .Z(n356) );
  AND U713 ( .A(n357), .B(p_input[9680]), .Z(o[9680]) );
  AND U714 ( .A(p_input[29680]), .B(p_input[19680]), .Z(n357) );
  AND U715 ( .A(n358), .B(p_input[967]), .Z(o[967]) );
  AND U716 ( .A(p_input[20967]), .B(p_input[10967]), .Z(n358) );
  AND U717 ( .A(n359), .B(p_input[9679]), .Z(o[9679]) );
  AND U718 ( .A(p_input[29679]), .B(p_input[19679]), .Z(n359) );
  AND U719 ( .A(n360), .B(p_input[9678]), .Z(o[9678]) );
  AND U720 ( .A(p_input[29678]), .B(p_input[19678]), .Z(n360) );
  AND U721 ( .A(n361), .B(p_input[9677]), .Z(o[9677]) );
  AND U722 ( .A(p_input[29677]), .B(p_input[19677]), .Z(n361) );
  AND U723 ( .A(n362), .B(p_input[9676]), .Z(o[9676]) );
  AND U724 ( .A(p_input[29676]), .B(p_input[19676]), .Z(n362) );
  AND U725 ( .A(n363), .B(p_input[9675]), .Z(o[9675]) );
  AND U726 ( .A(p_input[29675]), .B(p_input[19675]), .Z(n363) );
  AND U727 ( .A(n364), .B(p_input[9674]), .Z(o[9674]) );
  AND U728 ( .A(p_input[29674]), .B(p_input[19674]), .Z(n364) );
  AND U729 ( .A(n365), .B(p_input[9673]), .Z(o[9673]) );
  AND U730 ( .A(p_input[29673]), .B(p_input[19673]), .Z(n365) );
  AND U731 ( .A(n366), .B(p_input[9672]), .Z(o[9672]) );
  AND U732 ( .A(p_input[29672]), .B(p_input[19672]), .Z(n366) );
  AND U733 ( .A(n367), .B(p_input[9671]), .Z(o[9671]) );
  AND U734 ( .A(p_input[29671]), .B(p_input[19671]), .Z(n367) );
  AND U735 ( .A(n368), .B(p_input[9670]), .Z(o[9670]) );
  AND U736 ( .A(p_input[29670]), .B(p_input[19670]), .Z(n368) );
  AND U737 ( .A(n369), .B(p_input[966]), .Z(o[966]) );
  AND U738 ( .A(p_input[20966]), .B(p_input[10966]), .Z(n369) );
  AND U739 ( .A(n370), .B(p_input[9669]), .Z(o[9669]) );
  AND U740 ( .A(p_input[29669]), .B(p_input[19669]), .Z(n370) );
  AND U741 ( .A(n371), .B(p_input[9668]), .Z(o[9668]) );
  AND U742 ( .A(p_input[29668]), .B(p_input[19668]), .Z(n371) );
  AND U743 ( .A(n372), .B(p_input[9667]), .Z(o[9667]) );
  AND U744 ( .A(p_input[29667]), .B(p_input[19667]), .Z(n372) );
  AND U745 ( .A(n373), .B(p_input[9666]), .Z(o[9666]) );
  AND U746 ( .A(p_input[29666]), .B(p_input[19666]), .Z(n373) );
  AND U747 ( .A(n374), .B(p_input[9665]), .Z(o[9665]) );
  AND U748 ( .A(p_input[29665]), .B(p_input[19665]), .Z(n374) );
  AND U749 ( .A(n375), .B(p_input[9664]), .Z(o[9664]) );
  AND U750 ( .A(p_input[29664]), .B(p_input[19664]), .Z(n375) );
  AND U751 ( .A(n376), .B(p_input[9663]), .Z(o[9663]) );
  AND U752 ( .A(p_input[29663]), .B(p_input[19663]), .Z(n376) );
  AND U753 ( .A(n377), .B(p_input[9662]), .Z(o[9662]) );
  AND U754 ( .A(p_input[29662]), .B(p_input[19662]), .Z(n377) );
  AND U755 ( .A(n378), .B(p_input[9661]), .Z(o[9661]) );
  AND U756 ( .A(p_input[29661]), .B(p_input[19661]), .Z(n378) );
  AND U757 ( .A(n379), .B(p_input[9660]), .Z(o[9660]) );
  AND U758 ( .A(p_input[29660]), .B(p_input[19660]), .Z(n379) );
  AND U759 ( .A(n380), .B(p_input[965]), .Z(o[965]) );
  AND U760 ( .A(p_input[20965]), .B(p_input[10965]), .Z(n380) );
  AND U761 ( .A(n381), .B(p_input[9659]), .Z(o[9659]) );
  AND U762 ( .A(p_input[29659]), .B(p_input[19659]), .Z(n381) );
  AND U763 ( .A(n382), .B(p_input[9658]), .Z(o[9658]) );
  AND U764 ( .A(p_input[29658]), .B(p_input[19658]), .Z(n382) );
  AND U765 ( .A(n383), .B(p_input[9657]), .Z(o[9657]) );
  AND U766 ( .A(p_input[29657]), .B(p_input[19657]), .Z(n383) );
  AND U767 ( .A(n384), .B(p_input[9656]), .Z(o[9656]) );
  AND U768 ( .A(p_input[29656]), .B(p_input[19656]), .Z(n384) );
  AND U769 ( .A(n385), .B(p_input[9655]), .Z(o[9655]) );
  AND U770 ( .A(p_input[29655]), .B(p_input[19655]), .Z(n385) );
  AND U771 ( .A(n386), .B(p_input[9654]), .Z(o[9654]) );
  AND U772 ( .A(p_input[29654]), .B(p_input[19654]), .Z(n386) );
  AND U773 ( .A(n387), .B(p_input[9653]), .Z(o[9653]) );
  AND U774 ( .A(p_input[29653]), .B(p_input[19653]), .Z(n387) );
  AND U775 ( .A(n388), .B(p_input[9652]), .Z(o[9652]) );
  AND U776 ( .A(p_input[29652]), .B(p_input[19652]), .Z(n388) );
  AND U777 ( .A(n389), .B(p_input[9651]), .Z(o[9651]) );
  AND U778 ( .A(p_input[29651]), .B(p_input[19651]), .Z(n389) );
  AND U779 ( .A(n390), .B(p_input[9650]), .Z(o[9650]) );
  AND U780 ( .A(p_input[29650]), .B(p_input[19650]), .Z(n390) );
  AND U781 ( .A(n391), .B(p_input[964]), .Z(o[964]) );
  AND U782 ( .A(p_input[20964]), .B(p_input[10964]), .Z(n391) );
  AND U783 ( .A(n392), .B(p_input[9649]), .Z(o[9649]) );
  AND U784 ( .A(p_input[29649]), .B(p_input[19649]), .Z(n392) );
  AND U785 ( .A(n393), .B(p_input[9648]), .Z(o[9648]) );
  AND U786 ( .A(p_input[29648]), .B(p_input[19648]), .Z(n393) );
  AND U787 ( .A(n394), .B(p_input[9647]), .Z(o[9647]) );
  AND U788 ( .A(p_input[29647]), .B(p_input[19647]), .Z(n394) );
  AND U789 ( .A(n395), .B(p_input[9646]), .Z(o[9646]) );
  AND U790 ( .A(p_input[29646]), .B(p_input[19646]), .Z(n395) );
  AND U791 ( .A(n396), .B(p_input[9645]), .Z(o[9645]) );
  AND U792 ( .A(p_input[29645]), .B(p_input[19645]), .Z(n396) );
  AND U793 ( .A(n397), .B(p_input[9644]), .Z(o[9644]) );
  AND U794 ( .A(p_input[29644]), .B(p_input[19644]), .Z(n397) );
  AND U795 ( .A(n398), .B(p_input[9643]), .Z(o[9643]) );
  AND U796 ( .A(p_input[29643]), .B(p_input[19643]), .Z(n398) );
  AND U797 ( .A(n399), .B(p_input[9642]), .Z(o[9642]) );
  AND U798 ( .A(p_input[29642]), .B(p_input[19642]), .Z(n399) );
  AND U799 ( .A(n400), .B(p_input[9641]), .Z(o[9641]) );
  AND U800 ( .A(p_input[29641]), .B(p_input[19641]), .Z(n400) );
  AND U801 ( .A(n401), .B(p_input[9640]), .Z(o[9640]) );
  AND U802 ( .A(p_input[29640]), .B(p_input[19640]), .Z(n401) );
  AND U803 ( .A(n402), .B(p_input[963]), .Z(o[963]) );
  AND U804 ( .A(p_input[20963]), .B(p_input[10963]), .Z(n402) );
  AND U805 ( .A(n403), .B(p_input[9639]), .Z(o[9639]) );
  AND U806 ( .A(p_input[29639]), .B(p_input[19639]), .Z(n403) );
  AND U807 ( .A(n404), .B(p_input[9638]), .Z(o[9638]) );
  AND U808 ( .A(p_input[29638]), .B(p_input[19638]), .Z(n404) );
  AND U809 ( .A(n405), .B(p_input[9637]), .Z(o[9637]) );
  AND U810 ( .A(p_input[29637]), .B(p_input[19637]), .Z(n405) );
  AND U811 ( .A(n406), .B(p_input[9636]), .Z(o[9636]) );
  AND U812 ( .A(p_input[29636]), .B(p_input[19636]), .Z(n406) );
  AND U813 ( .A(n407), .B(p_input[9635]), .Z(o[9635]) );
  AND U814 ( .A(p_input[29635]), .B(p_input[19635]), .Z(n407) );
  AND U815 ( .A(n408), .B(p_input[9634]), .Z(o[9634]) );
  AND U816 ( .A(p_input[29634]), .B(p_input[19634]), .Z(n408) );
  AND U817 ( .A(n409), .B(p_input[9633]), .Z(o[9633]) );
  AND U818 ( .A(p_input[29633]), .B(p_input[19633]), .Z(n409) );
  AND U819 ( .A(n410), .B(p_input[9632]), .Z(o[9632]) );
  AND U820 ( .A(p_input[29632]), .B(p_input[19632]), .Z(n410) );
  AND U821 ( .A(n411), .B(p_input[9631]), .Z(o[9631]) );
  AND U822 ( .A(p_input[29631]), .B(p_input[19631]), .Z(n411) );
  AND U823 ( .A(n412), .B(p_input[9630]), .Z(o[9630]) );
  AND U824 ( .A(p_input[29630]), .B(p_input[19630]), .Z(n412) );
  AND U825 ( .A(n413), .B(p_input[962]), .Z(o[962]) );
  AND U826 ( .A(p_input[20962]), .B(p_input[10962]), .Z(n413) );
  AND U827 ( .A(n414), .B(p_input[9629]), .Z(o[9629]) );
  AND U828 ( .A(p_input[29629]), .B(p_input[19629]), .Z(n414) );
  AND U829 ( .A(n415), .B(p_input[9628]), .Z(o[9628]) );
  AND U830 ( .A(p_input[29628]), .B(p_input[19628]), .Z(n415) );
  AND U831 ( .A(n416), .B(p_input[9627]), .Z(o[9627]) );
  AND U832 ( .A(p_input[29627]), .B(p_input[19627]), .Z(n416) );
  AND U833 ( .A(n417), .B(p_input[9626]), .Z(o[9626]) );
  AND U834 ( .A(p_input[29626]), .B(p_input[19626]), .Z(n417) );
  AND U835 ( .A(n418), .B(p_input[9625]), .Z(o[9625]) );
  AND U836 ( .A(p_input[29625]), .B(p_input[19625]), .Z(n418) );
  AND U837 ( .A(n419), .B(p_input[9624]), .Z(o[9624]) );
  AND U838 ( .A(p_input[29624]), .B(p_input[19624]), .Z(n419) );
  AND U839 ( .A(n420), .B(p_input[9623]), .Z(o[9623]) );
  AND U840 ( .A(p_input[29623]), .B(p_input[19623]), .Z(n420) );
  AND U841 ( .A(n421), .B(p_input[9622]), .Z(o[9622]) );
  AND U842 ( .A(p_input[29622]), .B(p_input[19622]), .Z(n421) );
  AND U843 ( .A(n422), .B(p_input[9621]), .Z(o[9621]) );
  AND U844 ( .A(p_input[29621]), .B(p_input[19621]), .Z(n422) );
  AND U845 ( .A(n423), .B(p_input[9620]), .Z(o[9620]) );
  AND U846 ( .A(p_input[29620]), .B(p_input[19620]), .Z(n423) );
  AND U847 ( .A(n424), .B(p_input[961]), .Z(o[961]) );
  AND U848 ( .A(p_input[20961]), .B(p_input[10961]), .Z(n424) );
  AND U849 ( .A(n425), .B(p_input[9619]), .Z(o[9619]) );
  AND U850 ( .A(p_input[29619]), .B(p_input[19619]), .Z(n425) );
  AND U851 ( .A(n426), .B(p_input[9618]), .Z(o[9618]) );
  AND U852 ( .A(p_input[29618]), .B(p_input[19618]), .Z(n426) );
  AND U853 ( .A(n427), .B(p_input[9617]), .Z(o[9617]) );
  AND U854 ( .A(p_input[29617]), .B(p_input[19617]), .Z(n427) );
  AND U855 ( .A(n428), .B(p_input[9616]), .Z(o[9616]) );
  AND U856 ( .A(p_input[29616]), .B(p_input[19616]), .Z(n428) );
  AND U857 ( .A(n429), .B(p_input[9615]), .Z(o[9615]) );
  AND U858 ( .A(p_input[29615]), .B(p_input[19615]), .Z(n429) );
  AND U859 ( .A(n430), .B(p_input[9614]), .Z(o[9614]) );
  AND U860 ( .A(p_input[29614]), .B(p_input[19614]), .Z(n430) );
  AND U861 ( .A(n431), .B(p_input[9613]), .Z(o[9613]) );
  AND U862 ( .A(p_input[29613]), .B(p_input[19613]), .Z(n431) );
  AND U863 ( .A(n432), .B(p_input[9612]), .Z(o[9612]) );
  AND U864 ( .A(p_input[29612]), .B(p_input[19612]), .Z(n432) );
  AND U865 ( .A(n433), .B(p_input[9611]), .Z(o[9611]) );
  AND U866 ( .A(p_input[29611]), .B(p_input[19611]), .Z(n433) );
  AND U867 ( .A(n434), .B(p_input[9610]), .Z(o[9610]) );
  AND U868 ( .A(p_input[29610]), .B(p_input[19610]), .Z(n434) );
  AND U869 ( .A(n435), .B(p_input[960]), .Z(o[960]) );
  AND U870 ( .A(p_input[20960]), .B(p_input[10960]), .Z(n435) );
  AND U871 ( .A(n436), .B(p_input[9609]), .Z(o[9609]) );
  AND U872 ( .A(p_input[29609]), .B(p_input[19609]), .Z(n436) );
  AND U873 ( .A(n437), .B(p_input[9608]), .Z(o[9608]) );
  AND U874 ( .A(p_input[29608]), .B(p_input[19608]), .Z(n437) );
  AND U875 ( .A(n438), .B(p_input[9607]), .Z(o[9607]) );
  AND U876 ( .A(p_input[29607]), .B(p_input[19607]), .Z(n438) );
  AND U877 ( .A(n439), .B(p_input[9606]), .Z(o[9606]) );
  AND U878 ( .A(p_input[29606]), .B(p_input[19606]), .Z(n439) );
  AND U879 ( .A(n440), .B(p_input[9605]), .Z(o[9605]) );
  AND U880 ( .A(p_input[29605]), .B(p_input[19605]), .Z(n440) );
  AND U881 ( .A(n441), .B(p_input[9604]), .Z(o[9604]) );
  AND U882 ( .A(p_input[29604]), .B(p_input[19604]), .Z(n441) );
  AND U883 ( .A(n442), .B(p_input[9603]), .Z(o[9603]) );
  AND U884 ( .A(p_input[29603]), .B(p_input[19603]), .Z(n442) );
  AND U885 ( .A(n443), .B(p_input[9602]), .Z(o[9602]) );
  AND U886 ( .A(p_input[29602]), .B(p_input[19602]), .Z(n443) );
  AND U887 ( .A(n444), .B(p_input[9601]), .Z(o[9601]) );
  AND U888 ( .A(p_input[29601]), .B(p_input[19601]), .Z(n444) );
  AND U889 ( .A(n445), .B(p_input[9600]), .Z(o[9600]) );
  AND U890 ( .A(p_input[29600]), .B(p_input[19600]), .Z(n445) );
  AND U891 ( .A(n446), .B(p_input[95]), .Z(o[95]) );
  AND U892 ( .A(p_input[20095]), .B(p_input[10095]), .Z(n446) );
  AND U893 ( .A(n447), .B(p_input[959]), .Z(o[959]) );
  AND U894 ( .A(p_input[20959]), .B(p_input[10959]), .Z(n447) );
  AND U895 ( .A(n448), .B(p_input[9599]), .Z(o[9599]) );
  AND U896 ( .A(p_input[29599]), .B(p_input[19599]), .Z(n448) );
  AND U897 ( .A(n449), .B(p_input[9598]), .Z(o[9598]) );
  AND U898 ( .A(p_input[29598]), .B(p_input[19598]), .Z(n449) );
  AND U899 ( .A(n450), .B(p_input[9597]), .Z(o[9597]) );
  AND U900 ( .A(p_input[29597]), .B(p_input[19597]), .Z(n450) );
  AND U901 ( .A(n451), .B(p_input[9596]), .Z(o[9596]) );
  AND U902 ( .A(p_input[29596]), .B(p_input[19596]), .Z(n451) );
  AND U903 ( .A(n452), .B(p_input[9595]), .Z(o[9595]) );
  AND U904 ( .A(p_input[29595]), .B(p_input[19595]), .Z(n452) );
  AND U905 ( .A(n453), .B(p_input[9594]), .Z(o[9594]) );
  AND U906 ( .A(p_input[29594]), .B(p_input[19594]), .Z(n453) );
  AND U907 ( .A(n454), .B(p_input[9593]), .Z(o[9593]) );
  AND U908 ( .A(p_input[29593]), .B(p_input[19593]), .Z(n454) );
  AND U909 ( .A(n455), .B(p_input[9592]), .Z(o[9592]) );
  AND U910 ( .A(p_input[29592]), .B(p_input[19592]), .Z(n455) );
  AND U911 ( .A(n456), .B(p_input[9591]), .Z(o[9591]) );
  AND U912 ( .A(p_input[29591]), .B(p_input[19591]), .Z(n456) );
  AND U913 ( .A(n457), .B(p_input[9590]), .Z(o[9590]) );
  AND U914 ( .A(p_input[29590]), .B(p_input[19590]), .Z(n457) );
  AND U915 ( .A(n458), .B(p_input[958]), .Z(o[958]) );
  AND U916 ( .A(p_input[20958]), .B(p_input[10958]), .Z(n458) );
  AND U917 ( .A(n459), .B(p_input[9589]), .Z(o[9589]) );
  AND U918 ( .A(p_input[29589]), .B(p_input[19589]), .Z(n459) );
  AND U919 ( .A(n460), .B(p_input[9588]), .Z(o[9588]) );
  AND U920 ( .A(p_input[29588]), .B(p_input[19588]), .Z(n460) );
  AND U921 ( .A(n461), .B(p_input[9587]), .Z(o[9587]) );
  AND U922 ( .A(p_input[29587]), .B(p_input[19587]), .Z(n461) );
  AND U923 ( .A(n462), .B(p_input[9586]), .Z(o[9586]) );
  AND U924 ( .A(p_input[29586]), .B(p_input[19586]), .Z(n462) );
  AND U925 ( .A(n463), .B(p_input[9585]), .Z(o[9585]) );
  AND U926 ( .A(p_input[29585]), .B(p_input[19585]), .Z(n463) );
  AND U927 ( .A(n464), .B(p_input[9584]), .Z(o[9584]) );
  AND U928 ( .A(p_input[29584]), .B(p_input[19584]), .Z(n464) );
  AND U929 ( .A(n465), .B(p_input[9583]), .Z(o[9583]) );
  AND U930 ( .A(p_input[29583]), .B(p_input[19583]), .Z(n465) );
  AND U931 ( .A(n466), .B(p_input[9582]), .Z(o[9582]) );
  AND U932 ( .A(p_input[29582]), .B(p_input[19582]), .Z(n466) );
  AND U933 ( .A(n467), .B(p_input[9581]), .Z(o[9581]) );
  AND U934 ( .A(p_input[29581]), .B(p_input[19581]), .Z(n467) );
  AND U935 ( .A(n468), .B(p_input[9580]), .Z(o[9580]) );
  AND U936 ( .A(p_input[29580]), .B(p_input[19580]), .Z(n468) );
  AND U937 ( .A(n469), .B(p_input[957]), .Z(o[957]) );
  AND U938 ( .A(p_input[20957]), .B(p_input[10957]), .Z(n469) );
  AND U939 ( .A(n470), .B(p_input[9579]), .Z(o[9579]) );
  AND U940 ( .A(p_input[29579]), .B(p_input[19579]), .Z(n470) );
  AND U941 ( .A(n471), .B(p_input[9578]), .Z(o[9578]) );
  AND U942 ( .A(p_input[29578]), .B(p_input[19578]), .Z(n471) );
  AND U943 ( .A(n472), .B(p_input[9577]), .Z(o[9577]) );
  AND U944 ( .A(p_input[29577]), .B(p_input[19577]), .Z(n472) );
  AND U945 ( .A(n473), .B(p_input[9576]), .Z(o[9576]) );
  AND U946 ( .A(p_input[29576]), .B(p_input[19576]), .Z(n473) );
  AND U947 ( .A(n474), .B(p_input[9575]), .Z(o[9575]) );
  AND U948 ( .A(p_input[29575]), .B(p_input[19575]), .Z(n474) );
  AND U949 ( .A(n475), .B(p_input[9574]), .Z(o[9574]) );
  AND U950 ( .A(p_input[29574]), .B(p_input[19574]), .Z(n475) );
  AND U951 ( .A(n476), .B(p_input[9573]), .Z(o[9573]) );
  AND U952 ( .A(p_input[29573]), .B(p_input[19573]), .Z(n476) );
  AND U953 ( .A(n477), .B(p_input[9572]), .Z(o[9572]) );
  AND U954 ( .A(p_input[29572]), .B(p_input[19572]), .Z(n477) );
  AND U955 ( .A(n478), .B(p_input[9571]), .Z(o[9571]) );
  AND U956 ( .A(p_input[29571]), .B(p_input[19571]), .Z(n478) );
  AND U957 ( .A(n479), .B(p_input[9570]), .Z(o[9570]) );
  AND U958 ( .A(p_input[29570]), .B(p_input[19570]), .Z(n479) );
  AND U959 ( .A(n480), .B(p_input[956]), .Z(o[956]) );
  AND U960 ( .A(p_input[20956]), .B(p_input[10956]), .Z(n480) );
  AND U961 ( .A(n481), .B(p_input[9569]), .Z(o[9569]) );
  AND U962 ( .A(p_input[29569]), .B(p_input[19569]), .Z(n481) );
  AND U963 ( .A(n482), .B(p_input[9568]), .Z(o[9568]) );
  AND U964 ( .A(p_input[29568]), .B(p_input[19568]), .Z(n482) );
  AND U965 ( .A(n483), .B(p_input[9567]), .Z(o[9567]) );
  AND U966 ( .A(p_input[29567]), .B(p_input[19567]), .Z(n483) );
  AND U967 ( .A(n484), .B(p_input[9566]), .Z(o[9566]) );
  AND U968 ( .A(p_input[29566]), .B(p_input[19566]), .Z(n484) );
  AND U969 ( .A(n485), .B(p_input[9565]), .Z(o[9565]) );
  AND U970 ( .A(p_input[29565]), .B(p_input[19565]), .Z(n485) );
  AND U971 ( .A(n486), .B(p_input[9564]), .Z(o[9564]) );
  AND U972 ( .A(p_input[29564]), .B(p_input[19564]), .Z(n486) );
  AND U973 ( .A(n487), .B(p_input[9563]), .Z(o[9563]) );
  AND U974 ( .A(p_input[29563]), .B(p_input[19563]), .Z(n487) );
  AND U975 ( .A(n488), .B(p_input[9562]), .Z(o[9562]) );
  AND U976 ( .A(p_input[29562]), .B(p_input[19562]), .Z(n488) );
  AND U977 ( .A(n489), .B(p_input[9561]), .Z(o[9561]) );
  AND U978 ( .A(p_input[29561]), .B(p_input[19561]), .Z(n489) );
  AND U979 ( .A(n490), .B(p_input[9560]), .Z(o[9560]) );
  AND U980 ( .A(p_input[29560]), .B(p_input[19560]), .Z(n490) );
  AND U981 ( .A(n491), .B(p_input[955]), .Z(o[955]) );
  AND U982 ( .A(p_input[20955]), .B(p_input[10955]), .Z(n491) );
  AND U983 ( .A(n492), .B(p_input[9559]), .Z(o[9559]) );
  AND U984 ( .A(p_input[29559]), .B(p_input[19559]), .Z(n492) );
  AND U985 ( .A(n493), .B(p_input[9558]), .Z(o[9558]) );
  AND U986 ( .A(p_input[29558]), .B(p_input[19558]), .Z(n493) );
  AND U987 ( .A(n494), .B(p_input[9557]), .Z(o[9557]) );
  AND U988 ( .A(p_input[29557]), .B(p_input[19557]), .Z(n494) );
  AND U989 ( .A(n495), .B(p_input[9556]), .Z(o[9556]) );
  AND U990 ( .A(p_input[29556]), .B(p_input[19556]), .Z(n495) );
  AND U991 ( .A(n496), .B(p_input[9555]), .Z(o[9555]) );
  AND U992 ( .A(p_input[29555]), .B(p_input[19555]), .Z(n496) );
  AND U993 ( .A(n497), .B(p_input[9554]), .Z(o[9554]) );
  AND U994 ( .A(p_input[29554]), .B(p_input[19554]), .Z(n497) );
  AND U995 ( .A(n498), .B(p_input[9553]), .Z(o[9553]) );
  AND U996 ( .A(p_input[29553]), .B(p_input[19553]), .Z(n498) );
  AND U997 ( .A(n499), .B(p_input[9552]), .Z(o[9552]) );
  AND U998 ( .A(p_input[29552]), .B(p_input[19552]), .Z(n499) );
  AND U999 ( .A(n500), .B(p_input[9551]), .Z(o[9551]) );
  AND U1000 ( .A(p_input[29551]), .B(p_input[19551]), .Z(n500) );
  AND U1001 ( .A(n501), .B(p_input[9550]), .Z(o[9550]) );
  AND U1002 ( .A(p_input[29550]), .B(p_input[19550]), .Z(n501) );
  AND U1003 ( .A(n502), .B(p_input[954]), .Z(o[954]) );
  AND U1004 ( .A(p_input[20954]), .B(p_input[10954]), .Z(n502) );
  AND U1005 ( .A(n503), .B(p_input[9549]), .Z(o[9549]) );
  AND U1006 ( .A(p_input[29549]), .B(p_input[19549]), .Z(n503) );
  AND U1007 ( .A(n504), .B(p_input[9548]), .Z(o[9548]) );
  AND U1008 ( .A(p_input[29548]), .B(p_input[19548]), .Z(n504) );
  AND U1009 ( .A(n505), .B(p_input[9547]), .Z(o[9547]) );
  AND U1010 ( .A(p_input[29547]), .B(p_input[19547]), .Z(n505) );
  AND U1011 ( .A(n506), .B(p_input[9546]), .Z(o[9546]) );
  AND U1012 ( .A(p_input[29546]), .B(p_input[19546]), .Z(n506) );
  AND U1013 ( .A(n507), .B(p_input[9545]), .Z(o[9545]) );
  AND U1014 ( .A(p_input[29545]), .B(p_input[19545]), .Z(n507) );
  AND U1015 ( .A(n508), .B(p_input[9544]), .Z(o[9544]) );
  AND U1016 ( .A(p_input[29544]), .B(p_input[19544]), .Z(n508) );
  AND U1017 ( .A(n509), .B(p_input[9543]), .Z(o[9543]) );
  AND U1018 ( .A(p_input[29543]), .B(p_input[19543]), .Z(n509) );
  AND U1019 ( .A(n510), .B(p_input[9542]), .Z(o[9542]) );
  AND U1020 ( .A(p_input[29542]), .B(p_input[19542]), .Z(n510) );
  AND U1021 ( .A(n511), .B(p_input[9541]), .Z(o[9541]) );
  AND U1022 ( .A(p_input[29541]), .B(p_input[19541]), .Z(n511) );
  AND U1023 ( .A(n512), .B(p_input[9540]), .Z(o[9540]) );
  AND U1024 ( .A(p_input[29540]), .B(p_input[19540]), .Z(n512) );
  AND U1025 ( .A(n513), .B(p_input[953]), .Z(o[953]) );
  AND U1026 ( .A(p_input[20953]), .B(p_input[10953]), .Z(n513) );
  AND U1027 ( .A(n514), .B(p_input[9539]), .Z(o[9539]) );
  AND U1028 ( .A(p_input[29539]), .B(p_input[19539]), .Z(n514) );
  AND U1029 ( .A(n515), .B(p_input[9538]), .Z(o[9538]) );
  AND U1030 ( .A(p_input[29538]), .B(p_input[19538]), .Z(n515) );
  AND U1031 ( .A(n516), .B(p_input[9537]), .Z(o[9537]) );
  AND U1032 ( .A(p_input[29537]), .B(p_input[19537]), .Z(n516) );
  AND U1033 ( .A(n517), .B(p_input[9536]), .Z(o[9536]) );
  AND U1034 ( .A(p_input[29536]), .B(p_input[19536]), .Z(n517) );
  AND U1035 ( .A(n518), .B(p_input[9535]), .Z(o[9535]) );
  AND U1036 ( .A(p_input[29535]), .B(p_input[19535]), .Z(n518) );
  AND U1037 ( .A(n519), .B(p_input[9534]), .Z(o[9534]) );
  AND U1038 ( .A(p_input[29534]), .B(p_input[19534]), .Z(n519) );
  AND U1039 ( .A(n520), .B(p_input[9533]), .Z(o[9533]) );
  AND U1040 ( .A(p_input[29533]), .B(p_input[19533]), .Z(n520) );
  AND U1041 ( .A(n521), .B(p_input[9532]), .Z(o[9532]) );
  AND U1042 ( .A(p_input[29532]), .B(p_input[19532]), .Z(n521) );
  AND U1043 ( .A(n522), .B(p_input[9531]), .Z(o[9531]) );
  AND U1044 ( .A(p_input[29531]), .B(p_input[19531]), .Z(n522) );
  AND U1045 ( .A(n523), .B(p_input[9530]), .Z(o[9530]) );
  AND U1046 ( .A(p_input[29530]), .B(p_input[19530]), .Z(n523) );
  AND U1047 ( .A(n524), .B(p_input[952]), .Z(o[952]) );
  AND U1048 ( .A(p_input[20952]), .B(p_input[10952]), .Z(n524) );
  AND U1049 ( .A(n525), .B(p_input[9529]), .Z(o[9529]) );
  AND U1050 ( .A(p_input[29529]), .B(p_input[19529]), .Z(n525) );
  AND U1051 ( .A(n526), .B(p_input[9528]), .Z(o[9528]) );
  AND U1052 ( .A(p_input[29528]), .B(p_input[19528]), .Z(n526) );
  AND U1053 ( .A(n527), .B(p_input[9527]), .Z(o[9527]) );
  AND U1054 ( .A(p_input[29527]), .B(p_input[19527]), .Z(n527) );
  AND U1055 ( .A(n528), .B(p_input[9526]), .Z(o[9526]) );
  AND U1056 ( .A(p_input[29526]), .B(p_input[19526]), .Z(n528) );
  AND U1057 ( .A(n529), .B(p_input[9525]), .Z(o[9525]) );
  AND U1058 ( .A(p_input[29525]), .B(p_input[19525]), .Z(n529) );
  AND U1059 ( .A(n530), .B(p_input[9524]), .Z(o[9524]) );
  AND U1060 ( .A(p_input[29524]), .B(p_input[19524]), .Z(n530) );
  AND U1061 ( .A(n531), .B(p_input[9523]), .Z(o[9523]) );
  AND U1062 ( .A(p_input[29523]), .B(p_input[19523]), .Z(n531) );
  AND U1063 ( .A(n532), .B(p_input[9522]), .Z(o[9522]) );
  AND U1064 ( .A(p_input[29522]), .B(p_input[19522]), .Z(n532) );
  AND U1065 ( .A(n533), .B(p_input[9521]), .Z(o[9521]) );
  AND U1066 ( .A(p_input[29521]), .B(p_input[19521]), .Z(n533) );
  AND U1067 ( .A(n534), .B(p_input[9520]), .Z(o[9520]) );
  AND U1068 ( .A(p_input[29520]), .B(p_input[19520]), .Z(n534) );
  AND U1069 ( .A(n535), .B(p_input[951]), .Z(o[951]) );
  AND U1070 ( .A(p_input[20951]), .B(p_input[10951]), .Z(n535) );
  AND U1071 ( .A(n536), .B(p_input[9519]), .Z(o[9519]) );
  AND U1072 ( .A(p_input[29519]), .B(p_input[19519]), .Z(n536) );
  AND U1073 ( .A(n537), .B(p_input[9518]), .Z(o[9518]) );
  AND U1074 ( .A(p_input[29518]), .B(p_input[19518]), .Z(n537) );
  AND U1075 ( .A(n538), .B(p_input[9517]), .Z(o[9517]) );
  AND U1076 ( .A(p_input[29517]), .B(p_input[19517]), .Z(n538) );
  AND U1077 ( .A(n539), .B(p_input[9516]), .Z(o[9516]) );
  AND U1078 ( .A(p_input[29516]), .B(p_input[19516]), .Z(n539) );
  AND U1079 ( .A(n540), .B(p_input[9515]), .Z(o[9515]) );
  AND U1080 ( .A(p_input[29515]), .B(p_input[19515]), .Z(n540) );
  AND U1081 ( .A(n541), .B(p_input[9514]), .Z(o[9514]) );
  AND U1082 ( .A(p_input[29514]), .B(p_input[19514]), .Z(n541) );
  AND U1083 ( .A(n542), .B(p_input[9513]), .Z(o[9513]) );
  AND U1084 ( .A(p_input[29513]), .B(p_input[19513]), .Z(n542) );
  AND U1085 ( .A(n543), .B(p_input[9512]), .Z(o[9512]) );
  AND U1086 ( .A(p_input[29512]), .B(p_input[19512]), .Z(n543) );
  AND U1087 ( .A(n544), .B(p_input[9511]), .Z(o[9511]) );
  AND U1088 ( .A(p_input[29511]), .B(p_input[19511]), .Z(n544) );
  AND U1089 ( .A(n545), .B(p_input[9510]), .Z(o[9510]) );
  AND U1090 ( .A(p_input[29510]), .B(p_input[19510]), .Z(n545) );
  AND U1091 ( .A(n546), .B(p_input[950]), .Z(o[950]) );
  AND U1092 ( .A(p_input[20950]), .B(p_input[10950]), .Z(n546) );
  AND U1093 ( .A(n547), .B(p_input[9509]), .Z(o[9509]) );
  AND U1094 ( .A(p_input[29509]), .B(p_input[19509]), .Z(n547) );
  AND U1095 ( .A(n548), .B(p_input[9508]), .Z(o[9508]) );
  AND U1096 ( .A(p_input[29508]), .B(p_input[19508]), .Z(n548) );
  AND U1097 ( .A(n549), .B(p_input[9507]), .Z(o[9507]) );
  AND U1098 ( .A(p_input[29507]), .B(p_input[19507]), .Z(n549) );
  AND U1099 ( .A(n550), .B(p_input[9506]), .Z(o[9506]) );
  AND U1100 ( .A(p_input[29506]), .B(p_input[19506]), .Z(n550) );
  AND U1101 ( .A(n551), .B(p_input[9505]), .Z(o[9505]) );
  AND U1102 ( .A(p_input[29505]), .B(p_input[19505]), .Z(n551) );
  AND U1103 ( .A(n552), .B(p_input[9504]), .Z(o[9504]) );
  AND U1104 ( .A(p_input[29504]), .B(p_input[19504]), .Z(n552) );
  AND U1105 ( .A(n553), .B(p_input[9503]), .Z(o[9503]) );
  AND U1106 ( .A(p_input[29503]), .B(p_input[19503]), .Z(n553) );
  AND U1107 ( .A(n554), .B(p_input[9502]), .Z(o[9502]) );
  AND U1108 ( .A(p_input[29502]), .B(p_input[19502]), .Z(n554) );
  AND U1109 ( .A(n555), .B(p_input[9501]), .Z(o[9501]) );
  AND U1110 ( .A(p_input[29501]), .B(p_input[19501]), .Z(n555) );
  AND U1111 ( .A(n556), .B(p_input[9500]), .Z(o[9500]) );
  AND U1112 ( .A(p_input[29500]), .B(p_input[19500]), .Z(n556) );
  AND U1113 ( .A(n557), .B(p_input[94]), .Z(o[94]) );
  AND U1114 ( .A(p_input[20094]), .B(p_input[10094]), .Z(n557) );
  AND U1115 ( .A(n558), .B(p_input[949]), .Z(o[949]) );
  AND U1116 ( .A(p_input[20949]), .B(p_input[10949]), .Z(n558) );
  AND U1117 ( .A(n559), .B(p_input[9499]), .Z(o[9499]) );
  AND U1118 ( .A(p_input[29499]), .B(p_input[19499]), .Z(n559) );
  AND U1119 ( .A(n560), .B(p_input[9498]), .Z(o[9498]) );
  AND U1120 ( .A(p_input[29498]), .B(p_input[19498]), .Z(n560) );
  AND U1121 ( .A(n561), .B(p_input[9497]), .Z(o[9497]) );
  AND U1122 ( .A(p_input[29497]), .B(p_input[19497]), .Z(n561) );
  AND U1123 ( .A(n562), .B(p_input[9496]), .Z(o[9496]) );
  AND U1124 ( .A(p_input[29496]), .B(p_input[19496]), .Z(n562) );
  AND U1125 ( .A(n563), .B(p_input[9495]), .Z(o[9495]) );
  AND U1126 ( .A(p_input[29495]), .B(p_input[19495]), .Z(n563) );
  AND U1127 ( .A(n564), .B(p_input[9494]), .Z(o[9494]) );
  AND U1128 ( .A(p_input[29494]), .B(p_input[19494]), .Z(n564) );
  AND U1129 ( .A(n565), .B(p_input[9493]), .Z(o[9493]) );
  AND U1130 ( .A(p_input[29493]), .B(p_input[19493]), .Z(n565) );
  AND U1131 ( .A(n566), .B(p_input[9492]), .Z(o[9492]) );
  AND U1132 ( .A(p_input[29492]), .B(p_input[19492]), .Z(n566) );
  AND U1133 ( .A(n567), .B(p_input[9491]), .Z(o[9491]) );
  AND U1134 ( .A(p_input[29491]), .B(p_input[19491]), .Z(n567) );
  AND U1135 ( .A(n568), .B(p_input[9490]), .Z(o[9490]) );
  AND U1136 ( .A(p_input[29490]), .B(p_input[19490]), .Z(n568) );
  AND U1137 ( .A(n569), .B(p_input[948]), .Z(o[948]) );
  AND U1138 ( .A(p_input[20948]), .B(p_input[10948]), .Z(n569) );
  AND U1139 ( .A(n570), .B(p_input[9489]), .Z(o[9489]) );
  AND U1140 ( .A(p_input[29489]), .B(p_input[19489]), .Z(n570) );
  AND U1141 ( .A(n571), .B(p_input[9488]), .Z(o[9488]) );
  AND U1142 ( .A(p_input[29488]), .B(p_input[19488]), .Z(n571) );
  AND U1143 ( .A(n572), .B(p_input[9487]), .Z(o[9487]) );
  AND U1144 ( .A(p_input[29487]), .B(p_input[19487]), .Z(n572) );
  AND U1145 ( .A(n573), .B(p_input[9486]), .Z(o[9486]) );
  AND U1146 ( .A(p_input[29486]), .B(p_input[19486]), .Z(n573) );
  AND U1147 ( .A(n574), .B(p_input[9485]), .Z(o[9485]) );
  AND U1148 ( .A(p_input[29485]), .B(p_input[19485]), .Z(n574) );
  AND U1149 ( .A(n575), .B(p_input[9484]), .Z(o[9484]) );
  AND U1150 ( .A(p_input[29484]), .B(p_input[19484]), .Z(n575) );
  AND U1151 ( .A(n576), .B(p_input[9483]), .Z(o[9483]) );
  AND U1152 ( .A(p_input[29483]), .B(p_input[19483]), .Z(n576) );
  AND U1153 ( .A(n577), .B(p_input[9482]), .Z(o[9482]) );
  AND U1154 ( .A(p_input[29482]), .B(p_input[19482]), .Z(n577) );
  AND U1155 ( .A(n578), .B(p_input[9481]), .Z(o[9481]) );
  AND U1156 ( .A(p_input[29481]), .B(p_input[19481]), .Z(n578) );
  AND U1157 ( .A(n579), .B(p_input[9480]), .Z(o[9480]) );
  AND U1158 ( .A(p_input[29480]), .B(p_input[19480]), .Z(n579) );
  AND U1159 ( .A(n580), .B(p_input[947]), .Z(o[947]) );
  AND U1160 ( .A(p_input[20947]), .B(p_input[10947]), .Z(n580) );
  AND U1161 ( .A(n581), .B(p_input[9479]), .Z(o[9479]) );
  AND U1162 ( .A(p_input[29479]), .B(p_input[19479]), .Z(n581) );
  AND U1163 ( .A(n582), .B(p_input[9478]), .Z(o[9478]) );
  AND U1164 ( .A(p_input[29478]), .B(p_input[19478]), .Z(n582) );
  AND U1165 ( .A(n583), .B(p_input[9477]), .Z(o[9477]) );
  AND U1166 ( .A(p_input[29477]), .B(p_input[19477]), .Z(n583) );
  AND U1167 ( .A(n584), .B(p_input[9476]), .Z(o[9476]) );
  AND U1168 ( .A(p_input[29476]), .B(p_input[19476]), .Z(n584) );
  AND U1169 ( .A(n585), .B(p_input[9475]), .Z(o[9475]) );
  AND U1170 ( .A(p_input[29475]), .B(p_input[19475]), .Z(n585) );
  AND U1171 ( .A(n586), .B(p_input[9474]), .Z(o[9474]) );
  AND U1172 ( .A(p_input[29474]), .B(p_input[19474]), .Z(n586) );
  AND U1173 ( .A(n587), .B(p_input[9473]), .Z(o[9473]) );
  AND U1174 ( .A(p_input[29473]), .B(p_input[19473]), .Z(n587) );
  AND U1175 ( .A(n588), .B(p_input[9472]), .Z(o[9472]) );
  AND U1176 ( .A(p_input[29472]), .B(p_input[19472]), .Z(n588) );
  AND U1177 ( .A(n589), .B(p_input[9471]), .Z(o[9471]) );
  AND U1178 ( .A(p_input[29471]), .B(p_input[19471]), .Z(n589) );
  AND U1179 ( .A(n590), .B(p_input[9470]), .Z(o[9470]) );
  AND U1180 ( .A(p_input[29470]), .B(p_input[19470]), .Z(n590) );
  AND U1181 ( .A(n591), .B(p_input[946]), .Z(o[946]) );
  AND U1182 ( .A(p_input[20946]), .B(p_input[10946]), .Z(n591) );
  AND U1183 ( .A(n592), .B(p_input[9469]), .Z(o[9469]) );
  AND U1184 ( .A(p_input[29469]), .B(p_input[19469]), .Z(n592) );
  AND U1185 ( .A(n593), .B(p_input[9468]), .Z(o[9468]) );
  AND U1186 ( .A(p_input[29468]), .B(p_input[19468]), .Z(n593) );
  AND U1187 ( .A(n594), .B(p_input[9467]), .Z(o[9467]) );
  AND U1188 ( .A(p_input[29467]), .B(p_input[19467]), .Z(n594) );
  AND U1189 ( .A(n595), .B(p_input[9466]), .Z(o[9466]) );
  AND U1190 ( .A(p_input[29466]), .B(p_input[19466]), .Z(n595) );
  AND U1191 ( .A(n596), .B(p_input[9465]), .Z(o[9465]) );
  AND U1192 ( .A(p_input[29465]), .B(p_input[19465]), .Z(n596) );
  AND U1193 ( .A(n597), .B(p_input[9464]), .Z(o[9464]) );
  AND U1194 ( .A(p_input[29464]), .B(p_input[19464]), .Z(n597) );
  AND U1195 ( .A(n598), .B(p_input[9463]), .Z(o[9463]) );
  AND U1196 ( .A(p_input[29463]), .B(p_input[19463]), .Z(n598) );
  AND U1197 ( .A(n599), .B(p_input[9462]), .Z(o[9462]) );
  AND U1198 ( .A(p_input[29462]), .B(p_input[19462]), .Z(n599) );
  AND U1199 ( .A(n600), .B(p_input[9461]), .Z(o[9461]) );
  AND U1200 ( .A(p_input[29461]), .B(p_input[19461]), .Z(n600) );
  AND U1201 ( .A(n601), .B(p_input[9460]), .Z(o[9460]) );
  AND U1202 ( .A(p_input[29460]), .B(p_input[19460]), .Z(n601) );
  AND U1203 ( .A(n602), .B(p_input[945]), .Z(o[945]) );
  AND U1204 ( .A(p_input[20945]), .B(p_input[10945]), .Z(n602) );
  AND U1205 ( .A(n603), .B(p_input[9459]), .Z(o[9459]) );
  AND U1206 ( .A(p_input[29459]), .B(p_input[19459]), .Z(n603) );
  AND U1207 ( .A(n604), .B(p_input[9458]), .Z(o[9458]) );
  AND U1208 ( .A(p_input[29458]), .B(p_input[19458]), .Z(n604) );
  AND U1209 ( .A(n605), .B(p_input[9457]), .Z(o[9457]) );
  AND U1210 ( .A(p_input[29457]), .B(p_input[19457]), .Z(n605) );
  AND U1211 ( .A(n606), .B(p_input[9456]), .Z(o[9456]) );
  AND U1212 ( .A(p_input[29456]), .B(p_input[19456]), .Z(n606) );
  AND U1213 ( .A(n607), .B(p_input[9455]), .Z(o[9455]) );
  AND U1214 ( .A(p_input[29455]), .B(p_input[19455]), .Z(n607) );
  AND U1215 ( .A(n608), .B(p_input[9454]), .Z(o[9454]) );
  AND U1216 ( .A(p_input[29454]), .B(p_input[19454]), .Z(n608) );
  AND U1217 ( .A(n609), .B(p_input[9453]), .Z(o[9453]) );
  AND U1218 ( .A(p_input[29453]), .B(p_input[19453]), .Z(n609) );
  AND U1219 ( .A(n610), .B(p_input[9452]), .Z(o[9452]) );
  AND U1220 ( .A(p_input[29452]), .B(p_input[19452]), .Z(n610) );
  AND U1221 ( .A(n611), .B(p_input[9451]), .Z(o[9451]) );
  AND U1222 ( .A(p_input[29451]), .B(p_input[19451]), .Z(n611) );
  AND U1223 ( .A(n612), .B(p_input[9450]), .Z(o[9450]) );
  AND U1224 ( .A(p_input[29450]), .B(p_input[19450]), .Z(n612) );
  AND U1225 ( .A(n613), .B(p_input[944]), .Z(o[944]) );
  AND U1226 ( .A(p_input[20944]), .B(p_input[10944]), .Z(n613) );
  AND U1227 ( .A(n614), .B(p_input[9449]), .Z(o[9449]) );
  AND U1228 ( .A(p_input[29449]), .B(p_input[19449]), .Z(n614) );
  AND U1229 ( .A(n615), .B(p_input[9448]), .Z(o[9448]) );
  AND U1230 ( .A(p_input[29448]), .B(p_input[19448]), .Z(n615) );
  AND U1231 ( .A(n616), .B(p_input[9447]), .Z(o[9447]) );
  AND U1232 ( .A(p_input[29447]), .B(p_input[19447]), .Z(n616) );
  AND U1233 ( .A(n617), .B(p_input[9446]), .Z(o[9446]) );
  AND U1234 ( .A(p_input[29446]), .B(p_input[19446]), .Z(n617) );
  AND U1235 ( .A(n618), .B(p_input[9445]), .Z(o[9445]) );
  AND U1236 ( .A(p_input[29445]), .B(p_input[19445]), .Z(n618) );
  AND U1237 ( .A(n619), .B(p_input[9444]), .Z(o[9444]) );
  AND U1238 ( .A(p_input[29444]), .B(p_input[19444]), .Z(n619) );
  AND U1239 ( .A(n620), .B(p_input[9443]), .Z(o[9443]) );
  AND U1240 ( .A(p_input[29443]), .B(p_input[19443]), .Z(n620) );
  AND U1241 ( .A(n621), .B(p_input[9442]), .Z(o[9442]) );
  AND U1242 ( .A(p_input[29442]), .B(p_input[19442]), .Z(n621) );
  AND U1243 ( .A(n622), .B(p_input[9441]), .Z(o[9441]) );
  AND U1244 ( .A(p_input[29441]), .B(p_input[19441]), .Z(n622) );
  AND U1245 ( .A(n623), .B(p_input[9440]), .Z(o[9440]) );
  AND U1246 ( .A(p_input[29440]), .B(p_input[19440]), .Z(n623) );
  AND U1247 ( .A(n624), .B(p_input[943]), .Z(o[943]) );
  AND U1248 ( .A(p_input[20943]), .B(p_input[10943]), .Z(n624) );
  AND U1249 ( .A(n625), .B(p_input[9439]), .Z(o[9439]) );
  AND U1250 ( .A(p_input[29439]), .B(p_input[19439]), .Z(n625) );
  AND U1251 ( .A(n626), .B(p_input[9438]), .Z(o[9438]) );
  AND U1252 ( .A(p_input[29438]), .B(p_input[19438]), .Z(n626) );
  AND U1253 ( .A(n627), .B(p_input[9437]), .Z(o[9437]) );
  AND U1254 ( .A(p_input[29437]), .B(p_input[19437]), .Z(n627) );
  AND U1255 ( .A(n628), .B(p_input[9436]), .Z(o[9436]) );
  AND U1256 ( .A(p_input[29436]), .B(p_input[19436]), .Z(n628) );
  AND U1257 ( .A(n629), .B(p_input[9435]), .Z(o[9435]) );
  AND U1258 ( .A(p_input[29435]), .B(p_input[19435]), .Z(n629) );
  AND U1259 ( .A(n630), .B(p_input[9434]), .Z(o[9434]) );
  AND U1260 ( .A(p_input[29434]), .B(p_input[19434]), .Z(n630) );
  AND U1261 ( .A(n631), .B(p_input[9433]), .Z(o[9433]) );
  AND U1262 ( .A(p_input[29433]), .B(p_input[19433]), .Z(n631) );
  AND U1263 ( .A(n632), .B(p_input[9432]), .Z(o[9432]) );
  AND U1264 ( .A(p_input[29432]), .B(p_input[19432]), .Z(n632) );
  AND U1265 ( .A(n633), .B(p_input[9431]), .Z(o[9431]) );
  AND U1266 ( .A(p_input[29431]), .B(p_input[19431]), .Z(n633) );
  AND U1267 ( .A(n634), .B(p_input[9430]), .Z(o[9430]) );
  AND U1268 ( .A(p_input[29430]), .B(p_input[19430]), .Z(n634) );
  AND U1269 ( .A(n635), .B(p_input[942]), .Z(o[942]) );
  AND U1270 ( .A(p_input[20942]), .B(p_input[10942]), .Z(n635) );
  AND U1271 ( .A(n636), .B(p_input[9429]), .Z(o[9429]) );
  AND U1272 ( .A(p_input[29429]), .B(p_input[19429]), .Z(n636) );
  AND U1273 ( .A(n637), .B(p_input[9428]), .Z(o[9428]) );
  AND U1274 ( .A(p_input[29428]), .B(p_input[19428]), .Z(n637) );
  AND U1275 ( .A(n638), .B(p_input[9427]), .Z(o[9427]) );
  AND U1276 ( .A(p_input[29427]), .B(p_input[19427]), .Z(n638) );
  AND U1277 ( .A(n639), .B(p_input[9426]), .Z(o[9426]) );
  AND U1278 ( .A(p_input[29426]), .B(p_input[19426]), .Z(n639) );
  AND U1279 ( .A(n640), .B(p_input[9425]), .Z(o[9425]) );
  AND U1280 ( .A(p_input[29425]), .B(p_input[19425]), .Z(n640) );
  AND U1281 ( .A(n641), .B(p_input[9424]), .Z(o[9424]) );
  AND U1282 ( .A(p_input[29424]), .B(p_input[19424]), .Z(n641) );
  AND U1283 ( .A(n642), .B(p_input[9423]), .Z(o[9423]) );
  AND U1284 ( .A(p_input[29423]), .B(p_input[19423]), .Z(n642) );
  AND U1285 ( .A(n643), .B(p_input[9422]), .Z(o[9422]) );
  AND U1286 ( .A(p_input[29422]), .B(p_input[19422]), .Z(n643) );
  AND U1287 ( .A(n644), .B(p_input[9421]), .Z(o[9421]) );
  AND U1288 ( .A(p_input[29421]), .B(p_input[19421]), .Z(n644) );
  AND U1289 ( .A(n645), .B(p_input[9420]), .Z(o[9420]) );
  AND U1290 ( .A(p_input[29420]), .B(p_input[19420]), .Z(n645) );
  AND U1291 ( .A(n646), .B(p_input[941]), .Z(o[941]) );
  AND U1292 ( .A(p_input[20941]), .B(p_input[10941]), .Z(n646) );
  AND U1293 ( .A(n647), .B(p_input[9419]), .Z(o[9419]) );
  AND U1294 ( .A(p_input[29419]), .B(p_input[19419]), .Z(n647) );
  AND U1295 ( .A(n648), .B(p_input[9418]), .Z(o[9418]) );
  AND U1296 ( .A(p_input[29418]), .B(p_input[19418]), .Z(n648) );
  AND U1297 ( .A(n649), .B(p_input[9417]), .Z(o[9417]) );
  AND U1298 ( .A(p_input[29417]), .B(p_input[19417]), .Z(n649) );
  AND U1299 ( .A(n650), .B(p_input[9416]), .Z(o[9416]) );
  AND U1300 ( .A(p_input[29416]), .B(p_input[19416]), .Z(n650) );
  AND U1301 ( .A(n651), .B(p_input[9415]), .Z(o[9415]) );
  AND U1302 ( .A(p_input[29415]), .B(p_input[19415]), .Z(n651) );
  AND U1303 ( .A(n652), .B(p_input[9414]), .Z(o[9414]) );
  AND U1304 ( .A(p_input[29414]), .B(p_input[19414]), .Z(n652) );
  AND U1305 ( .A(n653), .B(p_input[9413]), .Z(o[9413]) );
  AND U1306 ( .A(p_input[29413]), .B(p_input[19413]), .Z(n653) );
  AND U1307 ( .A(n654), .B(p_input[9412]), .Z(o[9412]) );
  AND U1308 ( .A(p_input[29412]), .B(p_input[19412]), .Z(n654) );
  AND U1309 ( .A(n655), .B(p_input[9411]), .Z(o[9411]) );
  AND U1310 ( .A(p_input[29411]), .B(p_input[19411]), .Z(n655) );
  AND U1311 ( .A(n656), .B(p_input[9410]), .Z(o[9410]) );
  AND U1312 ( .A(p_input[29410]), .B(p_input[19410]), .Z(n656) );
  AND U1313 ( .A(n657), .B(p_input[940]), .Z(o[940]) );
  AND U1314 ( .A(p_input[20940]), .B(p_input[10940]), .Z(n657) );
  AND U1315 ( .A(n658), .B(p_input[9409]), .Z(o[9409]) );
  AND U1316 ( .A(p_input[29409]), .B(p_input[19409]), .Z(n658) );
  AND U1317 ( .A(n659), .B(p_input[9408]), .Z(o[9408]) );
  AND U1318 ( .A(p_input[29408]), .B(p_input[19408]), .Z(n659) );
  AND U1319 ( .A(n660), .B(p_input[9407]), .Z(o[9407]) );
  AND U1320 ( .A(p_input[29407]), .B(p_input[19407]), .Z(n660) );
  AND U1321 ( .A(n661), .B(p_input[9406]), .Z(o[9406]) );
  AND U1322 ( .A(p_input[29406]), .B(p_input[19406]), .Z(n661) );
  AND U1323 ( .A(n662), .B(p_input[9405]), .Z(o[9405]) );
  AND U1324 ( .A(p_input[29405]), .B(p_input[19405]), .Z(n662) );
  AND U1325 ( .A(n663), .B(p_input[9404]), .Z(o[9404]) );
  AND U1326 ( .A(p_input[29404]), .B(p_input[19404]), .Z(n663) );
  AND U1327 ( .A(n664), .B(p_input[9403]), .Z(o[9403]) );
  AND U1328 ( .A(p_input[29403]), .B(p_input[19403]), .Z(n664) );
  AND U1329 ( .A(n665), .B(p_input[9402]), .Z(o[9402]) );
  AND U1330 ( .A(p_input[29402]), .B(p_input[19402]), .Z(n665) );
  AND U1331 ( .A(n666), .B(p_input[9401]), .Z(o[9401]) );
  AND U1332 ( .A(p_input[29401]), .B(p_input[19401]), .Z(n666) );
  AND U1333 ( .A(n667), .B(p_input[9400]), .Z(o[9400]) );
  AND U1334 ( .A(p_input[29400]), .B(p_input[19400]), .Z(n667) );
  AND U1335 ( .A(n668), .B(p_input[93]), .Z(o[93]) );
  AND U1336 ( .A(p_input[20093]), .B(p_input[10093]), .Z(n668) );
  AND U1337 ( .A(n669), .B(p_input[939]), .Z(o[939]) );
  AND U1338 ( .A(p_input[20939]), .B(p_input[10939]), .Z(n669) );
  AND U1339 ( .A(n670), .B(p_input[9399]), .Z(o[9399]) );
  AND U1340 ( .A(p_input[29399]), .B(p_input[19399]), .Z(n670) );
  AND U1341 ( .A(n671), .B(p_input[9398]), .Z(o[9398]) );
  AND U1342 ( .A(p_input[29398]), .B(p_input[19398]), .Z(n671) );
  AND U1343 ( .A(n672), .B(p_input[9397]), .Z(o[9397]) );
  AND U1344 ( .A(p_input[29397]), .B(p_input[19397]), .Z(n672) );
  AND U1345 ( .A(n673), .B(p_input[9396]), .Z(o[9396]) );
  AND U1346 ( .A(p_input[29396]), .B(p_input[19396]), .Z(n673) );
  AND U1347 ( .A(n674), .B(p_input[9395]), .Z(o[9395]) );
  AND U1348 ( .A(p_input[29395]), .B(p_input[19395]), .Z(n674) );
  AND U1349 ( .A(n675), .B(p_input[9394]), .Z(o[9394]) );
  AND U1350 ( .A(p_input[29394]), .B(p_input[19394]), .Z(n675) );
  AND U1351 ( .A(n676), .B(p_input[9393]), .Z(o[9393]) );
  AND U1352 ( .A(p_input[29393]), .B(p_input[19393]), .Z(n676) );
  AND U1353 ( .A(n677), .B(p_input[9392]), .Z(o[9392]) );
  AND U1354 ( .A(p_input[29392]), .B(p_input[19392]), .Z(n677) );
  AND U1355 ( .A(n678), .B(p_input[9391]), .Z(o[9391]) );
  AND U1356 ( .A(p_input[29391]), .B(p_input[19391]), .Z(n678) );
  AND U1357 ( .A(n679), .B(p_input[9390]), .Z(o[9390]) );
  AND U1358 ( .A(p_input[29390]), .B(p_input[19390]), .Z(n679) );
  AND U1359 ( .A(n680), .B(p_input[938]), .Z(o[938]) );
  AND U1360 ( .A(p_input[20938]), .B(p_input[10938]), .Z(n680) );
  AND U1361 ( .A(n681), .B(p_input[9389]), .Z(o[9389]) );
  AND U1362 ( .A(p_input[29389]), .B(p_input[19389]), .Z(n681) );
  AND U1363 ( .A(n682), .B(p_input[9388]), .Z(o[9388]) );
  AND U1364 ( .A(p_input[29388]), .B(p_input[19388]), .Z(n682) );
  AND U1365 ( .A(n683), .B(p_input[9387]), .Z(o[9387]) );
  AND U1366 ( .A(p_input[29387]), .B(p_input[19387]), .Z(n683) );
  AND U1367 ( .A(n684), .B(p_input[9386]), .Z(o[9386]) );
  AND U1368 ( .A(p_input[29386]), .B(p_input[19386]), .Z(n684) );
  AND U1369 ( .A(n685), .B(p_input[9385]), .Z(o[9385]) );
  AND U1370 ( .A(p_input[29385]), .B(p_input[19385]), .Z(n685) );
  AND U1371 ( .A(n686), .B(p_input[9384]), .Z(o[9384]) );
  AND U1372 ( .A(p_input[29384]), .B(p_input[19384]), .Z(n686) );
  AND U1373 ( .A(n687), .B(p_input[9383]), .Z(o[9383]) );
  AND U1374 ( .A(p_input[29383]), .B(p_input[19383]), .Z(n687) );
  AND U1375 ( .A(n688), .B(p_input[9382]), .Z(o[9382]) );
  AND U1376 ( .A(p_input[29382]), .B(p_input[19382]), .Z(n688) );
  AND U1377 ( .A(n689), .B(p_input[9381]), .Z(o[9381]) );
  AND U1378 ( .A(p_input[29381]), .B(p_input[19381]), .Z(n689) );
  AND U1379 ( .A(n690), .B(p_input[9380]), .Z(o[9380]) );
  AND U1380 ( .A(p_input[29380]), .B(p_input[19380]), .Z(n690) );
  AND U1381 ( .A(n691), .B(p_input[937]), .Z(o[937]) );
  AND U1382 ( .A(p_input[20937]), .B(p_input[10937]), .Z(n691) );
  AND U1383 ( .A(n692), .B(p_input[9379]), .Z(o[9379]) );
  AND U1384 ( .A(p_input[29379]), .B(p_input[19379]), .Z(n692) );
  AND U1385 ( .A(n693), .B(p_input[9378]), .Z(o[9378]) );
  AND U1386 ( .A(p_input[29378]), .B(p_input[19378]), .Z(n693) );
  AND U1387 ( .A(n694), .B(p_input[9377]), .Z(o[9377]) );
  AND U1388 ( .A(p_input[29377]), .B(p_input[19377]), .Z(n694) );
  AND U1389 ( .A(n695), .B(p_input[9376]), .Z(o[9376]) );
  AND U1390 ( .A(p_input[29376]), .B(p_input[19376]), .Z(n695) );
  AND U1391 ( .A(n696), .B(p_input[9375]), .Z(o[9375]) );
  AND U1392 ( .A(p_input[29375]), .B(p_input[19375]), .Z(n696) );
  AND U1393 ( .A(n697), .B(p_input[9374]), .Z(o[9374]) );
  AND U1394 ( .A(p_input[29374]), .B(p_input[19374]), .Z(n697) );
  AND U1395 ( .A(n698), .B(p_input[9373]), .Z(o[9373]) );
  AND U1396 ( .A(p_input[29373]), .B(p_input[19373]), .Z(n698) );
  AND U1397 ( .A(n699), .B(p_input[9372]), .Z(o[9372]) );
  AND U1398 ( .A(p_input[29372]), .B(p_input[19372]), .Z(n699) );
  AND U1399 ( .A(n700), .B(p_input[9371]), .Z(o[9371]) );
  AND U1400 ( .A(p_input[29371]), .B(p_input[19371]), .Z(n700) );
  AND U1401 ( .A(n701), .B(p_input[9370]), .Z(o[9370]) );
  AND U1402 ( .A(p_input[29370]), .B(p_input[19370]), .Z(n701) );
  AND U1403 ( .A(n702), .B(p_input[936]), .Z(o[936]) );
  AND U1404 ( .A(p_input[20936]), .B(p_input[10936]), .Z(n702) );
  AND U1405 ( .A(n703), .B(p_input[9369]), .Z(o[9369]) );
  AND U1406 ( .A(p_input[29369]), .B(p_input[19369]), .Z(n703) );
  AND U1407 ( .A(n704), .B(p_input[9368]), .Z(o[9368]) );
  AND U1408 ( .A(p_input[29368]), .B(p_input[19368]), .Z(n704) );
  AND U1409 ( .A(n705), .B(p_input[9367]), .Z(o[9367]) );
  AND U1410 ( .A(p_input[29367]), .B(p_input[19367]), .Z(n705) );
  AND U1411 ( .A(n706), .B(p_input[9366]), .Z(o[9366]) );
  AND U1412 ( .A(p_input[29366]), .B(p_input[19366]), .Z(n706) );
  AND U1413 ( .A(n707), .B(p_input[9365]), .Z(o[9365]) );
  AND U1414 ( .A(p_input[29365]), .B(p_input[19365]), .Z(n707) );
  AND U1415 ( .A(n708), .B(p_input[9364]), .Z(o[9364]) );
  AND U1416 ( .A(p_input[29364]), .B(p_input[19364]), .Z(n708) );
  AND U1417 ( .A(n709), .B(p_input[9363]), .Z(o[9363]) );
  AND U1418 ( .A(p_input[29363]), .B(p_input[19363]), .Z(n709) );
  AND U1419 ( .A(n710), .B(p_input[9362]), .Z(o[9362]) );
  AND U1420 ( .A(p_input[29362]), .B(p_input[19362]), .Z(n710) );
  AND U1421 ( .A(n711), .B(p_input[9361]), .Z(o[9361]) );
  AND U1422 ( .A(p_input[29361]), .B(p_input[19361]), .Z(n711) );
  AND U1423 ( .A(n712), .B(p_input[9360]), .Z(o[9360]) );
  AND U1424 ( .A(p_input[29360]), .B(p_input[19360]), .Z(n712) );
  AND U1425 ( .A(n713), .B(p_input[935]), .Z(o[935]) );
  AND U1426 ( .A(p_input[20935]), .B(p_input[10935]), .Z(n713) );
  AND U1427 ( .A(n714), .B(p_input[9359]), .Z(o[9359]) );
  AND U1428 ( .A(p_input[29359]), .B(p_input[19359]), .Z(n714) );
  AND U1429 ( .A(n715), .B(p_input[9358]), .Z(o[9358]) );
  AND U1430 ( .A(p_input[29358]), .B(p_input[19358]), .Z(n715) );
  AND U1431 ( .A(n716), .B(p_input[9357]), .Z(o[9357]) );
  AND U1432 ( .A(p_input[29357]), .B(p_input[19357]), .Z(n716) );
  AND U1433 ( .A(n717), .B(p_input[9356]), .Z(o[9356]) );
  AND U1434 ( .A(p_input[29356]), .B(p_input[19356]), .Z(n717) );
  AND U1435 ( .A(n718), .B(p_input[9355]), .Z(o[9355]) );
  AND U1436 ( .A(p_input[29355]), .B(p_input[19355]), .Z(n718) );
  AND U1437 ( .A(n719), .B(p_input[9354]), .Z(o[9354]) );
  AND U1438 ( .A(p_input[29354]), .B(p_input[19354]), .Z(n719) );
  AND U1439 ( .A(n720), .B(p_input[9353]), .Z(o[9353]) );
  AND U1440 ( .A(p_input[29353]), .B(p_input[19353]), .Z(n720) );
  AND U1441 ( .A(n721), .B(p_input[9352]), .Z(o[9352]) );
  AND U1442 ( .A(p_input[29352]), .B(p_input[19352]), .Z(n721) );
  AND U1443 ( .A(n722), .B(p_input[9351]), .Z(o[9351]) );
  AND U1444 ( .A(p_input[29351]), .B(p_input[19351]), .Z(n722) );
  AND U1445 ( .A(n723), .B(p_input[9350]), .Z(o[9350]) );
  AND U1446 ( .A(p_input[29350]), .B(p_input[19350]), .Z(n723) );
  AND U1447 ( .A(n724), .B(p_input[934]), .Z(o[934]) );
  AND U1448 ( .A(p_input[20934]), .B(p_input[10934]), .Z(n724) );
  AND U1449 ( .A(n725), .B(p_input[9349]), .Z(o[9349]) );
  AND U1450 ( .A(p_input[29349]), .B(p_input[19349]), .Z(n725) );
  AND U1451 ( .A(n726), .B(p_input[9348]), .Z(o[9348]) );
  AND U1452 ( .A(p_input[29348]), .B(p_input[19348]), .Z(n726) );
  AND U1453 ( .A(n727), .B(p_input[9347]), .Z(o[9347]) );
  AND U1454 ( .A(p_input[29347]), .B(p_input[19347]), .Z(n727) );
  AND U1455 ( .A(n728), .B(p_input[9346]), .Z(o[9346]) );
  AND U1456 ( .A(p_input[29346]), .B(p_input[19346]), .Z(n728) );
  AND U1457 ( .A(n729), .B(p_input[9345]), .Z(o[9345]) );
  AND U1458 ( .A(p_input[29345]), .B(p_input[19345]), .Z(n729) );
  AND U1459 ( .A(n730), .B(p_input[9344]), .Z(o[9344]) );
  AND U1460 ( .A(p_input[29344]), .B(p_input[19344]), .Z(n730) );
  AND U1461 ( .A(n731), .B(p_input[9343]), .Z(o[9343]) );
  AND U1462 ( .A(p_input[29343]), .B(p_input[19343]), .Z(n731) );
  AND U1463 ( .A(n732), .B(p_input[9342]), .Z(o[9342]) );
  AND U1464 ( .A(p_input[29342]), .B(p_input[19342]), .Z(n732) );
  AND U1465 ( .A(n733), .B(p_input[9341]), .Z(o[9341]) );
  AND U1466 ( .A(p_input[29341]), .B(p_input[19341]), .Z(n733) );
  AND U1467 ( .A(n734), .B(p_input[9340]), .Z(o[9340]) );
  AND U1468 ( .A(p_input[29340]), .B(p_input[19340]), .Z(n734) );
  AND U1469 ( .A(n735), .B(p_input[933]), .Z(o[933]) );
  AND U1470 ( .A(p_input[20933]), .B(p_input[10933]), .Z(n735) );
  AND U1471 ( .A(n736), .B(p_input[9339]), .Z(o[9339]) );
  AND U1472 ( .A(p_input[29339]), .B(p_input[19339]), .Z(n736) );
  AND U1473 ( .A(n737), .B(p_input[9338]), .Z(o[9338]) );
  AND U1474 ( .A(p_input[29338]), .B(p_input[19338]), .Z(n737) );
  AND U1475 ( .A(n738), .B(p_input[9337]), .Z(o[9337]) );
  AND U1476 ( .A(p_input[29337]), .B(p_input[19337]), .Z(n738) );
  AND U1477 ( .A(n739), .B(p_input[9336]), .Z(o[9336]) );
  AND U1478 ( .A(p_input[29336]), .B(p_input[19336]), .Z(n739) );
  AND U1479 ( .A(n740), .B(p_input[9335]), .Z(o[9335]) );
  AND U1480 ( .A(p_input[29335]), .B(p_input[19335]), .Z(n740) );
  AND U1481 ( .A(n741), .B(p_input[9334]), .Z(o[9334]) );
  AND U1482 ( .A(p_input[29334]), .B(p_input[19334]), .Z(n741) );
  AND U1483 ( .A(n742), .B(p_input[9333]), .Z(o[9333]) );
  AND U1484 ( .A(p_input[29333]), .B(p_input[19333]), .Z(n742) );
  AND U1485 ( .A(n743), .B(p_input[9332]), .Z(o[9332]) );
  AND U1486 ( .A(p_input[29332]), .B(p_input[19332]), .Z(n743) );
  AND U1487 ( .A(n744), .B(p_input[9331]), .Z(o[9331]) );
  AND U1488 ( .A(p_input[29331]), .B(p_input[19331]), .Z(n744) );
  AND U1489 ( .A(n745), .B(p_input[9330]), .Z(o[9330]) );
  AND U1490 ( .A(p_input[29330]), .B(p_input[19330]), .Z(n745) );
  AND U1491 ( .A(n746), .B(p_input[932]), .Z(o[932]) );
  AND U1492 ( .A(p_input[20932]), .B(p_input[10932]), .Z(n746) );
  AND U1493 ( .A(n747), .B(p_input[9329]), .Z(o[9329]) );
  AND U1494 ( .A(p_input[29329]), .B(p_input[19329]), .Z(n747) );
  AND U1495 ( .A(n748), .B(p_input[9328]), .Z(o[9328]) );
  AND U1496 ( .A(p_input[29328]), .B(p_input[19328]), .Z(n748) );
  AND U1497 ( .A(n749), .B(p_input[9327]), .Z(o[9327]) );
  AND U1498 ( .A(p_input[29327]), .B(p_input[19327]), .Z(n749) );
  AND U1499 ( .A(n750), .B(p_input[9326]), .Z(o[9326]) );
  AND U1500 ( .A(p_input[29326]), .B(p_input[19326]), .Z(n750) );
  AND U1501 ( .A(n751), .B(p_input[9325]), .Z(o[9325]) );
  AND U1502 ( .A(p_input[29325]), .B(p_input[19325]), .Z(n751) );
  AND U1503 ( .A(n752), .B(p_input[9324]), .Z(o[9324]) );
  AND U1504 ( .A(p_input[29324]), .B(p_input[19324]), .Z(n752) );
  AND U1505 ( .A(n753), .B(p_input[9323]), .Z(o[9323]) );
  AND U1506 ( .A(p_input[29323]), .B(p_input[19323]), .Z(n753) );
  AND U1507 ( .A(n754), .B(p_input[9322]), .Z(o[9322]) );
  AND U1508 ( .A(p_input[29322]), .B(p_input[19322]), .Z(n754) );
  AND U1509 ( .A(n755), .B(p_input[9321]), .Z(o[9321]) );
  AND U1510 ( .A(p_input[29321]), .B(p_input[19321]), .Z(n755) );
  AND U1511 ( .A(n756), .B(p_input[9320]), .Z(o[9320]) );
  AND U1512 ( .A(p_input[29320]), .B(p_input[19320]), .Z(n756) );
  AND U1513 ( .A(n757), .B(p_input[931]), .Z(o[931]) );
  AND U1514 ( .A(p_input[20931]), .B(p_input[10931]), .Z(n757) );
  AND U1515 ( .A(n758), .B(p_input[9319]), .Z(o[9319]) );
  AND U1516 ( .A(p_input[29319]), .B(p_input[19319]), .Z(n758) );
  AND U1517 ( .A(n759), .B(p_input[9318]), .Z(o[9318]) );
  AND U1518 ( .A(p_input[29318]), .B(p_input[19318]), .Z(n759) );
  AND U1519 ( .A(n760), .B(p_input[9317]), .Z(o[9317]) );
  AND U1520 ( .A(p_input[29317]), .B(p_input[19317]), .Z(n760) );
  AND U1521 ( .A(n761), .B(p_input[9316]), .Z(o[9316]) );
  AND U1522 ( .A(p_input[29316]), .B(p_input[19316]), .Z(n761) );
  AND U1523 ( .A(n762), .B(p_input[9315]), .Z(o[9315]) );
  AND U1524 ( .A(p_input[29315]), .B(p_input[19315]), .Z(n762) );
  AND U1525 ( .A(n763), .B(p_input[9314]), .Z(o[9314]) );
  AND U1526 ( .A(p_input[29314]), .B(p_input[19314]), .Z(n763) );
  AND U1527 ( .A(n764), .B(p_input[9313]), .Z(o[9313]) );
  AND U1528 ( .A(p_input[29313]), .B(p_input[19313]), .Z(n764) );
  AND U1529 ( .A(n765), .B(p_input[9312]), .Z(o[9312]) );
  AND U1530 ( .A(p_input[29312]), .B(p_input[19312]), .Z(n765) );
  AND U1531 ( .A(n766), .B(p_input[9311]), .Z(o[9311]) );
  AND U1532 ( .A(p_input[29311]), .B(p_input[19311]), .Z(n766) );
  AND U1533 ( .A(n767), .B(p_input[9310]), .Z(o[9310]) );
  AND U1534 ( .A(p_input[29310]), .B(p_input[19310]), .Z(n767) );
  AND U1535 ( .A(n768), .B(p_input[930]), .Z(o[930]) );
  AND U1536 ( .A(p_input[20930]), .B(p_input[10930]), .Z(n768) );
  AND U1537 ( .A(n769), .B(p_input[9309]), .Z(o[9309]) );
  AND U1538 ( .A(p_input[29309]), .B(p_input[19309]), .Z(n769) );
  AND U1539 ( .A(n770), .B(p_input[9308]), .Z(o[9308]) );
  AND U1540 ( .A(p_input[29308]), .B(p_input[19308]), .Z(n770) );
  AND U1541 ( .A(n771), .B(p_input[9307]), .Z(o[9307]) );
  AND U1542 ( .A(p_input[29307]), .B(p_input[19307]), .Z(n771) );
  AND U1543 ( .A(n772), .B(p_input[9306]), .Z(o[9306]) );
  AND U1544 ( .A(p_input[29306]), .B(p_input[19306]), .Z(n772) );
  AND U1545 ( .A(n773), .B(p_input[9305]), .Z(o[9305]) );
  AND U1546 ( .A(p_input[29305]), .B(p_input[19305]), .Z(n773) );
  AND U1547 ( .A(n774), .B(p_input[9304]), .Z(o[9304]) );
  AND U1548 ( .A(p_input[29304]), .B(p_input[19304]), .Z(n774) );
  AND U1549 ( .A(n775), .B(p_input[9303]), .Z(o[9303]) );
  AND U1550 ( .A(p_input[29303]), .B(p_input[19303]), .Z(n775) );
  AND U1551 ( .A(n776), .B(p_input[9302]), .Z(o[9302]) );
  AND U1552 ( .A(p_input[29302]), .B(p_input[19302]), .Z(n776) );
  AND U1553 ( .A(n777), .B(p_input[9301]), .Z(o[9301]) );
  AND U1554 ( .A(p_input[29301]), .B(p_input[19301]), .Z(n777) );
  AND U1555 ( .A(n778), .B(p_input[9300]), .Z(o[9300]) );
  AND U1556 ( .A(p_input[29300]), .B(p_input[19300]), .Z(n778) );
  AND U1557 ( .A(n779), .B(p_input[92]), .Z(o[92]) );
  AND U1558 ( .A(p_input[20092]), .B(p_input[10092]), .Z(n779) );
  AND U1559 ( .A(n780), .B(p_input[929]), .Z(o[929]) );
  AND U1560 ( .A(p_input[20929]), .B(p_input[10929]), .Z(n780) );
  AND U1561 ( .A(n781), .B(p_input[9299]), .Z(o[9299]) );
  AND U1562 ( .A(p_input[29299]), .B(p_input[19299]), .Z(n781) );
  AND U1563 ( .A(n782), .B(p_input[9298]), .Z(o[9298]) );
  AND U1564 ( .A(p_input[29298]), .B(p_input[19298]), .Z(n782) );
  AND U1565 ( .A(n783), .B(p_input[9297]), .Z(o[9297]) );
  AND U1566 ( .A(p_input[29297]), .B(p_input[19297]), .Z(n783) );
  AND U1567 ( .A(n784), .B(p_input[9296]), .Z(o[9296]) );
  AND U1568 ( .A(p_input[29296]), .B(p_input[19296]), .Z(n784) );
  AND U1569 ( .A(n785), .B(p_input[9295]), .Z(o[9295]) );
  AND U1570 ( .A(p_input[29295]), .B(p_input[19295]), .Z(n785) );
  AND U1571 ( .A(n786), .B(p_input[9294]), .Z(o[9294]) );
  AND U1572 ( .A(p_input[29294]), .B(p_input[19294]), .Z(n786) );
  AND U1573 ( .A(n787), .B(p_input[9293]), .Z(o[9293]) );
  AND U1574 ( .A(p_input[29293]), .B(p_input[19293]), .Z(n787) );
  AND U1575 ( .A(n788), .B(p_input[9292]), .Z(o[9292]) );
  AND U1576 ( .A(p_input[29292]), .B(p_input[19292]), .Z(n788) );
  AND U1577 ( .A(n789), .B(p_input[9291]), .Z(o[9291]) );
  AND U1578 ( .A(p_input[29291]), .B(p_input[19291]), .Z(n789) );
  AND U1579 ( .A(n790), .B(p_input[9290]), .Z(o[9290]) );
  AND U1580 ( .A(p_input[29290]), .B(p_input[19290]), .Z(n790) );
  AND U1581 ( .A(n791), .B(p_input[928]), .Z(o[928]) );
  AND U1582 ( .A(p_input[20928]), .B(p_input[10928]), .Z(n791) );
  AND U1583 ( .A(n792), .B(p_input[9289]), .Z(o[9289]) );
  AND U1584 ( .A(p_input[29289]), .B(p_input[19289]), .Z(n792) );
  AND U1585 ( .A(n793), .B(p_input[9288]), .Z(o[9288]) );
  AND U1586 ( .A(p_input[29288]), .B(p_input[19288]), .Z(n793) );
  AND U1587 ( .A(n794), .B(p_input[9287]), .Z(o[9287]) );
  AND U1588 ( .A(p_input[29287]), .B(p_input[19287]), .Z(n794) );
  AND U1589 ( .A(n795), .B(p_input[9286]), .Z(o[9286]) );
  AND U1590 ( .A(p_input[29286]), .B(p_input[19286]), .Z(n795) );
  AND U1591 ( .A(n796), .B(p_input[9285]), .Z(o[9285]) );
  AND U1592 ( .A(p_input[29285]), .B(p_input[19285]), .Z(n796) );
  AND U1593 ( .A(n797), .B(p_input[9284]), .Z(o[9284]) );
  AND U1594 ( .A(p_input[29284]), .B(p_input[19284]), .Z(n797) );
  AND U1595 ( .A(n798), .B(p_input[9283]), .Z(o[9283]) );
  AND U1596 ( .A(p_input[29283]), .B(p_input[19283]), .Z(n798) );
  AND U1597 ( .A(n799), .B(p_input[9282]), .Z(o[9282]) );
  AND U1598 ( .A(p_input[29282]), .B(p_input[19282]), .Z(n799) );
  AND U1599 ( .A(n800), .B(p_input[9281]), .Z(o[9281]) );
  AND U1600 ( .A(p_input[29281]), .B(p_input[19281]), .Z(n800) );
  AND U1601 ( .A(n801), .B(p_input[9280]), .Z(o[9280]) );
  AND U1602 ( .A(p_input[29280]), .B(p_input[19280]), .Z(n801) );
  AND U1603 ( .A(n802), .B(p_input[927]), .Z(o[927]) );
  AND U1604 ( .A(p_input[20927]), .B(p_input[10927]), .Z(n802) );
  AND U1605 ( .A(n803), .B(p_input[9279]), .Z(o[9279]) );
  AND U1606 ( .A(p_input[29279]), .B(p_input[19279]), .Z(n803) );
  AND U1607 ( .A(n804), .B(p_input[9278]), .Z(o[9278]) );
  AND U1608 ( .A(p_input[29278]), .B(p_input[19278]), .Z(n804) );
  AND U1609 ( .A(n805), .B(p_input[9277]), .Z(o[9277]) );
  AND U1610 ( .A(p_input[29277]), .B(p_input[19277]), .Z(n805) );
  AND U1611 ( .A(n806), .B(p_input[9276]), .Z(o[9276]) );
  AND U1612 ( .A(p_input[29276]), .B(p_input[19276]), .Z(n806) );
  AND U1613 ( .A(n807), .B(p_input[9275]), .Z(o[9275]) );
  AND U1614 ( .A(p_input[29275]), .B(p_input[19275]), .Z(n807) );
  AND U1615 ( .A(n808), .B(p_input[9274]), .Z(o[9274]) );
  AND U1616 ( .A(p_input[29274]), .B(p_input[19274]), .Z(n808) );
  AND U1617 ( .A(n809), .B(p_input[9273]), .Z(o[9273]) );
  AND U1618 ( .A(p_input[29273]), .B(p_input[19273]), .Z(n809) );
  AND U1619 ( .A(n810), .B(p_input[9272]), .Z(o[9272]) );
  AND U1620 ( .A(p_input[29272]), .B(p_input[19272]), .Z(n810) );
  AND U1621 ( .A(n811), .B(p_input[9271]), .Z(o[9271]) );
  AND U1622 ( .A(p_input[29271]), .B(p_input[19271]), .Z(n811) );
  AND U1623 ( .A(n812), .B(p_input[9270]), .Z(o[9270]) );
  AND U1624 ( .A(p_input[29270]), .B(p_input[19270]), .Z(n812) );
  AND U1625 ( .A(n813), .B(p_input[926]), .Z(o[926]) );
  AND U1626 ( .A(p_input[20926]), .B(p_input[10926]), .Z(n813) );
  AND U1627 ( .A(n814), .B(p_input[9269]), .Z(o[9269]) );
  AND U1628 ( .A(p_input[29269]), .B(p_input[19269]), .Z(n814) );
  AND U1629 ( .A(n815), .B(p_input[9268]), .Z(o[9268]) );
  AND U1630 ( .A(p_input[29268]), .B(p_input[19268]), .Z(n815) );
  AND U1631 ( .A(n816), .B(p_input[9267]), .Z(o[9267]) );
  AND U1632 ( .A(p_input[29267]), .B(p_input[19267]), .Z(n816) );
  AND U1633 ( .A(n817), .B(p_input[9266]), .Z(o[9266]) );
  AND U1634 ( .A(p_input[29266]), .B(p_input[19266]), .Z(n817) );
  AND U1635 ( .A(n818), .B(p_input[9265]), .Z(o[9265]) );
  AND U1636 ( .A(p_input[29265]), .B(p_input[19265]), .Z(n818) );
  AND U1637 ( .A(n819), .B(p_input[9264]), .Z(o[9264]) );
  AND U1638 ( .A(p_input[29264]), .B(p_input[19264]), .Z(n819) );
  AND U1639 ( .A(n820), .B(p_input[9263]), .Z(o[9263]) );
  AND U1640 ( .A(p_input[29263]), .B(p_input[19263]), .Z(n820) );
  AND U1641 ( .A(n821), .B(p_input[9262]), .Z(o[9262]) );
  AND U1642 ( .A(p_input[29262]), .B(p_input[19262]), .Z(n821) );
  AND U1643 ( .A(n822), .B(p_input[9261]), .Z(o[9261]) );
  AND U1644 ( .A(p_input[29261]), .B(p_input[19261]), .Z(n822) );
  AND U1645 ( .A(n823), .B(p_input[9260]), .Z(o[9260]) );
  AND U1646 ( .A(p_input[29260]), .B(p_input[19260]), .Z(n823) );
  AND U1647 ( .A(n824), .B(p_input[925]), .Z(o[925]) );
  AND U1648 ( .A(p_input[20925]), .B(p_input[10925]), .Z(n824) );
  AND U1649 ( .A(n825), .B(p_input[9259]), .Z(o[9259]) );
  AND U1650 ( .A(p_input[29259]), .B(p_input[19259]), .Z(n825) );
  AND U1651 ( .A(n826), .B(p_input[9258]), .Z(o[9258]) );
  AND U1652 ( .A(p_input[29258]), .B(p_input[19258]), .Z(n826) );
  AND U1653 ( .A(n827), .B(p_input[9257]), .Z(o[9257]) );
  AND U1654 ( .A(p_input[29257]), .B(p_input[19257]), .Z(n827) );
  AND U1655 ( .A(n828), .B(p_input[9256]), .Z(o[9256]) );
  AND U1656 ( .A(p_input[29256]), .B(p_input[19256]), .Z(n828) );
  AND U1657 ( .A(n829), .B(p_input[9255]), .Z(o[9255]) );
  AND U1658 ( .A(p_input[29255]), .B(p_input[19255]), .Z(n829) );
  AND U1659 ( .A(n830), .B(p_input[9254]), .Z(o[9254]) );
  AND U1660 ( .A(p_input[29254]), .B(p_input[19254]), .Z(n830) );
  AND U1661 ( .A(n831), .B(p_input[9253]), .Z(o[9253]) );
  AND U1662 ( .A(p_input[29253]), .B(p_input[19253]), .Z(n831) );
  AND U1663 ( .A(n832), .B(p_input[9252]), .Z(o[9252]) );
  AND U1664 ( .A(p_input[29252]), .B(p_input[19252]), .Z(n832) );
  AND U1665 ( .A(n833), .B(p_input[9251]), .Z(o[9251]) );
  AND U1666 ( .A(p_input[29251]), .B(p_input[19251]), .Z(n833) );
  AND U1667 ( .A(n834), .B(p_input[9250]), .Z(o[9250]) );
  AND U1668 ( .A(p_input[29250]), .B(p_input[19250]), .Z(n834) );
  AND U1669 ( .A(n835), .B(p_input[924]), .Z(o[924]) );
  AND U1670 ( .A(p_input[20924]), .B(p_input[10924]), .Z(n835) );
  AND U1671 ( .A(n836), .B(p_input[9249]), .Z(o[9249]) );
  AND U1672 ( .A(p_input[29249]), .B(p_input[19249]), .Z(n836) );
  AND U1673 ( .A(n837), .B(p_input[9248]), .Z(o[9248]) );
  AND U1674 ( .A(p_input[29248]), .B(p_input[19248]), .Z(n837) );
  AND U1675 ( .A(n838), .B(p_input[9247]), .Z(o[9247]) );
  AND U1676 ( .A(p_input[29247]), .B(p_input[19247]), .Z(n838) );
  AND U1677 ( .A(n839), .B(p_input[9246]), .Z(o[9246]) );
  AND U1678 ( .A(p_input[29246]), .B(p_input[19246]), .Z(n839) );
  AND U1679 ( .A(n840), .B(p_input[9245]), .Z(o[9245]) );
  AND U1680 ( .A(p_input[29245]), .B(p_input[19245]), .Z(n840) );
  AND U1681 ( .A(n841), .B(p_input[9244]), .Z(o[9244]) );
  AND U1682 ( .A(p_input[29244]), .B(p_input[19244]), .Z(n841) );
  AND U1683 ( .A(n842), .B(p_input[9243]), .Z(o[9243]) );
  AND U1684 ( .A(p_input[29243]), .B(p_input[19243]), .Z(n842) );
  AND U1685 ( .A(n843), .B(p_input[9242]), .Z(o[9242]) );
  AND U1686 ( .A(p_input[29242]), .B(p_input[19242]), .Z(n843) );
  AND U1687 ( .A(n844), .B(p_input[9241]), .Z(o[9241]) );
  AND U1688 ( .A(p_input[29241]), .B(p_input[19241]), .Z(n844) );
  AND U1689 ( .A(n845), .B(p_input[9240]), .Z(o[9240]) );
  AND U1690 ( .A(p_input[29240]), .B(p_input[19240]), .Z(n845) );
  AND U1691 ( .A(n846), .B(p_input[923]), .Z(o[923]) );
  AND U1692 ( .A(p_input[20923]), .B(p_input[10923]), .Z(n846) );
  AND U1693 ( .A(n847), .B(p_input[9239]), .Z(o[9239]) );
  AND U1694 ( .A(p_input[29239]), .B(p_input[19239]), .Z(n847) );
  AND U1695 ( .A(n848), .B(p_input[9238]), .Z(o[9238]) );
  AND U1696 ( .A(p_input[29238]), .B(p_input[19238]), .Z(n848) );
  AND U1697 ( .A(n849), .B(p_input[9237]), .Z(o[9237]) );
  AND U1698 ( .A(p_input[29237]), .B(p_input[19237]), .Z(n849) );
  AND U1699 ( .A(n850), .B(p_input[9236]), .Z(o[9236]) );
  AND U1700 ( .A(p_input[29236]), .B(p_input[19236]), .Z(n850) );
  AND U1701 ( .A(n851), .B(p_input[9235]), .Z(o[9235]) );
  AND U1702 ( .A(p_input[29235]), .B(p_input[19235]), .Z(n851) );
  AND U1703 ( .A(n852), .B(p_input[9234]), .Z(o[9234]) );
  AND U1704 ( .A(p_input[29234]), .B(p_input[19234]), .Z(n852) );
  AND U1705 ( .A(n853), .B(p_input[9233]), .Z(o[9233]) );
  AND U1706 ( .A(p_input[29233]), .B(p_input[19233]), .Z(n853) );
  AND U1707 ( .A(n854), .B(p_input[9232]), .Z(o[9232]) );
  AND U1708 ( .A(p_input[29232]), .B(p_input[19232]), .Z(n854) );
  AND U1709 ( .A(n855), .B(p_input[9231]), .Z(o[9231]) );
  AND U1710 ( .A(p_input[29231]), .B(p_input[19231]), .Z(n855) );
  AND U1711 ( .A(n856), .B(p_input[9230]), .Z(o[9230]) );
  AND U1712 ( .A(p_input[29230]), .B(p_input[19230]), .Z(n856) );
  AND U1713 ( .A(n857), .B(p_input[922]), .Z(o[922]) );
  AND U1714 ( .A(p_input[20922]), .B(p_input[10922]), .Z(n857) );
  AND U1715 ( .A(n858), .B(p_input[9229]), .Z(o[9229]) );
  AND U1716 ( .A(p_input[29229]), .B(p_input[19229]), .Z(n858) );
  AND U1717 ( .A(n859), .B(p_input[9228]), .Z(o[9228]) );
  AND U1718 ( .A(p_input[29228]), .B(p_input[19228]), .Z(n859) );
  AND U1719 ( .A(n860), .B(p_input[9227]), .Z(o[9227]) );
  AND U1720 ( .A(p_input[29227]), .B(p_input[19227]), .Z(n860) );
  AND U1721 ( .A(n861), .B(p_input[9226]), .Z(o[9226]) );
  AND U1722 ( .A(p_input[29226]), .B(p_input[19226]), .Z(n861) );
  AND U1723 ( .A(n862), .B(p_input[9225]), .Z(o[9225]) );
  AND U1724 ( .A(p_input[29225]), .B(p_input[19225]), .Z(n862) );
  AND U1725 ( .A(n863), .B(p_input[9224]), .Z(o[9224]) );
  AND U1726 ( .A(p_input[29224]), .B(p_input[19224]), .Z(n863) );
  AND U1727 ( .A(n864), .B(p_input[9223]), .Z(o[9223]) );
  AND U1728 ( .A(p_input[29223]), .B(p_input[19223]), .Z(n864) );
  AND U1729 ( .A(n865), .B(p_input[9222]), .Z(o[9222]) );
  AND U1730 ( .A(p_input[29222]), .B(p_input[19222]), .Z(n865) );
  AND U1731 ( .A(n866), .B(p_input[9221]), .Z(o[9221]) );
  AND U1732 ( .A(p_input[29221]), .B(p_input[19221]), .Z(n866) );
  AND U1733 ( .A(n867), .B(p_input[9220]), .Z(o[9220]) );
  AND U1734 ( .A(p_input[29220]), .B(p_input[19220]), .Z(n867) );
  AND U1735 ( .A(n868), .B(p_input[921]), .Z(o[921]) );
  AND U1736 ( .A(p_input[20921]), .B(p_input[10921]), .Z(n868) );
  AND U1737 ( .A(n869), .B(p_input[9219]), .Z(o[9219]) );
  AND U1738 ( .A(p_input[29219]), .B(p_input[19219]), .Z(n869) );
  AND U1739 ( .A(n870), .B(p_input[9218]), .Z(o[9218]) );
  AND U1740 ( .A(p_input[29218]), .B(p_input[19218]), .Z(n870) );
  AND U1741 ( .A(n871), .B(p_input[9217]), .Z(o[9217]) );
  AND U1742 ( .A(p_input[29217]), .B(p_input[19217]), .Z(n871) );
  AND U1743 ( .A(n872), .B(p_input[9216]), .Z(o[9216]) );
  AND U1744 ( .A(p_input[29216]), .B(p_input[19216]), .Z(n872) );
  AND U1745 ( .A(n873), .B(p_input[9215]), .Z(o[9215]) );
  AND U1746 ( .A(p_input[29215]), .B(p_input[19215]), .Z(n873) );
  AND U1747 ( .A(n874), .B(p_input[9214]), .Z(o[9214]) );
  AND U1748 ( .A(p_input[29214]), .B(p_input[19214]), .Z(n874) );
  AND U1749 ( .A(n875), .B(p_input[9213]), .Z(o[9213]) );
  AND U1750 ( .A(p_input[29213]), .B(p_input[19213]), .Z(n875) );
  AND U1751 ( .A(n876), .B(p_input[9212]), .Z(o[9212]) );
  AND U1752 ( .A(p_input[29212]), .B(p_input[19212]), .Z(n876) );
  AND U1753 ( .A(n877), .B(p_input[9211]), .Z(o[9211]) );
  AND U1754 ( .A(p_input[29211]), .B(p_input[19211]), .Z(n877) );
  AND U1755 ( .A(n878), .B(p_input[9210]), .Z(o[9210]) );
  AND U1756 ( .A(p_input[29210]), .B(p_input[19210]), .Z(n878) );
  AND U1757 ( .A(n879), .B(p_input[920]), .Z(o[920]) );
  AND U1758 ( .A(p_input[20920]), .B(p_input[10920]), .Z(n879) );
  AND U1759 ( .A(n880), .B(p_input[9209]), .Z(o[9209]) );
  AND U1760 ( .A(p_input[29209]), .B(p_input[19209]), .Z(n880) );
  AND U1761 ( .A(n881), .B(p_input[9208]), .Z(o[9208]) );
  AND U1762 ( .A(p_input[29208]), .B(p_input[19208]), .Z(n881) );
  AND U1763 ( .A(n882), .B(p_input[9207]), .Z(o[9207]) );
  AND U1764 ( .A(p_input[29207]), .B(p_input[19207]), .Z(n882) );
  AND U1765 ( .A(n883), .B(p_input[9206]), .Z(o[9206]) );
  AND U1766 ( .A(p_input[29206]), .B(p_input[19206]), .Z(n883) );
  AND U1767 ( .A(n884), .B(p_input[9205]), .Z(o[9205]) );
  AND U1768 ( .A(p_input[29205]), .B(p_input[19205]), .Z(n884) );
  AND U1769 ( .A(n885), .B(p_input[9204]), .Z(o[9204]) );
  AND U1770 ( .A(p_input[29204]), .B(p_input[19204]), .Z(n885) );
  AND U1771 ( .A(n886), .B(p_input[9203]), .Z(o[9203]) );
  AND U1772 ( .A(p_input[29203]), .B(p_input[19203]), .Z(n886) );
  AND U1773 ( .A(n887), .B(p_input[9202]), .Z(o[9202]) );
  AND U1774 ( .A(p_input[29202]), .B(p_input[19202]), .Z(n887) );
  AND U1775 ( .A(n888), .B(p_input[9201]), .Z(o[9201]) );
  AND U1776 ( .A(p_input[29201]), .B(p_input[19201]), .Z(n888) );
  AND U1777 ( .A(n889), .B(p_input[9200]), .Z(o[9200]) );
  AND U1778 ( .A(p_input[29200]), .B(p_input[19200]), .Z(n889) );
  AND U1779 ( .A(n890), .B(p_input[91]), .Z(o[91]) );
  AND U1780 ( .A(p_input[20091]), .B(p_input[10091]), .Z(n890) );
  AND U1781 ( .A(n891), .B(p_input[919]), .Z(o[919]) );
  AND U1782 ( .A(p_input[20919]), .B(p_input[10919]), .Z(n891) );
  AND U1783 ( .A(n892), .B(p_input[9199]), .Z(o[9199]) );
  AND U1784 ( .A(p_input[29199]), .B(p_input[19199]), .Z(n892) );
  AND U1785 ( .A(n893), .B(p_input[9198]), .Z(o[9198]) );
  AND U1786 ( .A(p_input[29198]), .B(p_input[19198]), .Z(n893) );
  AND U1787 ( .A(n894), .B(p_input[9197]), .Z(o[9197]) );
  AND U1788 ( .A(p_input[29197]), .B(p_input[19197]), .Z(n894) );
  AND U1789 ( .A(n895), .B(p_input[9196]), .Z(o[9196]) );
  AND U1790 ( .A(p_input[29196]), .B(p_input[19196]), .Z(n895) );
  AND U1791 ( .A(n896), .B(p_input[9195]), .Z(o[9195]) );
  AND U1792 ( .A(p_input[29195]), .B(p_input[19195]), .Z(n896) );
  AND U1793 ( .A(n897), .B(p_input[9194]), .Z(o[9194]) );
  AND U1794 ( .A(p_input[29194]), .B(p_input[19194]), .Z(n897) );
  AND U1795 ( .A(n898), .B(p_input[9193]), .Z(o[9193]) );
  AND U1796 ( .A(p_input[29193]), .B(p_input[19193]), .Z(n898) );
  AND U1797 ( .A(n899), .B(p_input[9192]), .Z(o[9192]) );
  AND U1798 ( .A(p_input[29192]), .B(p_input[19192]), .Z(n899) );
  AND U1799 ( .A(n900), .B(p_input[9191]), .Z(o[9191]) );
  AND U1800 ( .A(p_input[29191]), .B(p_input[19191]), .Z(n900) );
  AND U1801 ( .A(n901), .B(p_input[9190]), .Z(o[9190]) );
  AND U1802 ( .A(p_input[29190]), .B(p_input[19190]), .Z(n901) );
  AND U1803 ( .A(n902), .B(p_input[918]), .Z(o[918]) );
  AND U1804 ( .A(p_input[20918]), .B(p_input[10918]), .Z(n902) );
  AND U1805 ( .A(n903), .B(p_input[9189]), .Z(o[9189]) );
  AND U1806 ( .A(p_input[29189]), .B(p_input[19189]), .Z(n903) );
  AND U1807 ( .A(n904), .B(p_input[9188]), .Z(o[9188]) );
  AND U1808 ( .A(p_input[29188]), .B(p_input[19188]), .Z(n904) );
  AND U1809 ( .A(n905), .B(p_input[9187]), .Z(o[9187]) );
  AND U1810 ( .A(p_input[29187]), .B(p_input[19187]), .Z(n905) );
  AND U1811 ( .A(n906), .B(p_input[9186]), .Z(o[9186]) );
  AND U1812 ( .A(p_input[29186]), .B(p_input[19186]), .Z(n906) );
  AND U1813 ( .A(n907), .B(p_input[9185]), .Z(o[9185]) );
  AND U1814 ( .A(p_input[29185]), .B(p_input[19185]), .Z(n907) );
  AND U1815 ( .A(n908), .B(p_input[9184]), .Z(o[9184]) );
  AND U1816 ( .A(p_input[29184]), .B(p_input[19184]), .Z(n908) );
  AND U1817 ( .A(n909), .B(p_input[9183]), .Z(o[9183]) );
  AND U1818 ( .A(p_input[29183]), .B(p_input[19183]), .Z(n909) );
  AND U1819 ( .A(n910), .B(p_input[9182]), .Z(o[9182]) );
  AND U1820 ( .A(p_input[29182]), .B(p_input[19182]), .Z(n910) );
  AND U1821 ( .A(n911), .B(p_input[9181]), .Z(o[9181]) );
  AND U1822 ( .A(p_input[29181]), .B(p_input[19181]), .Z(n911) );
  AND U1823 ( .A(n912), .B(p_input[9180]), .Z(o[9180]) );
  AND U1824 ( .A(p_input[29180]), .B(p_input[19180]), .Z(n912) );
  AND U1825 ( .A(n913), .B(p_input[917]), .Z(o[917]) );
  AND U1826 ( .A(p_input[20917]), .B(p_input[10917]), .Z(n913) );
  AND U1827 ( .A(n914), .B(p_input[9179]), .Z(o[9179]) );
  AND U1828 ( .A(p_input[29179]), .B(p_input[19179]), .Z(n914) );
  AND U1829 ( .A(n915), .B(p_input[9178]), .Z(o[9178]) );
  AND U1830 ( .A(p_input[29178]), .B(p_input[19178]), .Z(n915) );
  AND U1831 ( .A(n916), .B(p_input[9177]), .Z(o[9177]) );
  AND U1832 ( .A(p_input[29177]), .B(p_input[19177]), .Z(n916) );
  AND U1833 ( .A(n917), .B(p_input[9176]), .Z(o[9176]) );
  AND U1834 ( .A(p_input[29176]), .B(p_input[19176]), .Z(n917) );
  AND U1835 ( .A(n918), .B(p_input[9175]), .Z(o[9175]) );
  AND U1836 ( .A(p_input[29175]), .B(p_input[19175]), .Z(n918) );
  AND U1837 ( .A(n919), .B(p_input[9174]), .Z(o[9174]) );
  AND U1838 ( .A(p_input[29174]), .B(p_input[19174]), .Z(n919) );
  AND U1839 ( .A(n920), .B(p_input[9173]), .Z(o[9173]) );
  AND U1840 ( .A(p_input[29173]), .B(p_input[19173]), .Z(n920) );
  AND U1841 ( .A(n921), .B(p_input[9172]), .Z(o[9172]) );
  AND U1842 ( .A(p_input[29172]), .B(p_input[19172]), .Z(n921) );
  AND U1843 ( .A(n922), .B(p_input[9171]), .Z(o[9171]) );
  AND U1844 ( .A(p_input[29171]), .B(p_input[19171]), .Z(n922) );
  AND U1845 ( .A(n923), .B(p_input[9170]), .Z(o[9170]) );
  AND U1846 ( .A(p_input[29170]), .B(p_input[19170]), .Z(n923) );
  AND U1847 ( .A(n924), .B(p_input[916]), .Z(o[916]) );
  AND U1848 ( .A(p_input[20916]), .B(p_input[10916]), .Z(n924) );
  AND U1849 ( .A(n925), .B(p_input[9169]), .Z(o[9169]) );
  AND U1850 ( .A(p_input[29169]), .B(p_input[19169]), .Z(n925) );
  AND U1851 ( .A(n926), .B(p_input[9168]), .Z(o[9168]) );
  AND U1852 ( .A(p_input[29168]), .B(p_input[19168]), .Z(n926) );
  AND U1853 ( .A(n927), .B(p_input[9167]), .Z(o[9167]) );
  AND U1854 ( .A(p_input[29167]), .B(p_input[19167]), .Z(n927) );
  AND U1855 ( .A(n928), .B(p_input[9166]), .Z(o[9166]) );
  AND U1856 ( .A(p_input[29166]), .B(p_input[19166]), .Z(n928) );
  AND U1857 ( .A(n929), .B(p_input[9165]), .Z(o[9165]) );
  AND U1858 ( .A(p_input[29165]), .B(p_input[19165]), .Z(n929) );
  AND U1859 ( .A(n930), .B(p_input[9164]), .Z(o[9164]) );
  AND U1860 ( .A(p_input[29164]), .B(p_input[19164]), .Z(n930) );
  AND U1861 ( .A(n931), .B(p_input[9163]), .Z(o[9163]) );
  AND U1862 ( .A(p_input[29163]), .B(p_input[19163]), .Z(n931) );
  AND U1863 ( .A(n932), .B(p_input[9162]), .Z(o[9162]) );
  AND U1864 ( .A(p_input[29162]), .B(p_input[19162]), .Z(n932) );
  AND U1865 ( .A(n933), .B(p_input[9161]), .Z(o[9161]) );
  AND U1866 ( .A(p_input[29161]), .B(p_input[19161]), .Z(n933) );
  AND U1867 ( .A(n934), .B(p_input[9160]), .Z(o[9160]) );
  AND U1868 ( .A(p_input[29160]), .B(p_input[19160]), .Z(n934) );
  AND U1869 ( .A(n935), .B(p_input[915]), .Z(o[915]) );
  AND U1870 ( .A(p_input[20915]), .B(p_input[10915]), .Z(n935) );
  AND U1871 ( .A(n936), .B(p_input[9159]), .Z(o[9159]) );
  AND U1872 ( .A(p_input[29159]), .B(p_input[19159]), .Z(n936) );
  AND U1873 ( .A(n937), .B(p_input[9158]), .Z(o[9158]) );
  AND U1874 ( .A(p_input[29158]), .B(p_input[19158]), .Z(n937) );
  AND U1875 ( .A(n938), .B(p_input[9157]), .Z(o[9157]) );
  AND U1876 ( .A(p_input[29157]), .B(p_input[19157]), .Z(n938) );
  AND U1877 ( .A(n939), .B(p_input[9156]), .Z(o[9156]) );
  AND U1878 ( .A(p_input[29156]), .B(p_input[19156]), .Z(n939) );
  AND U1879 ( .A(n940), .B(p_input[9155]), .Z(o[9155]) );
  AND U1880 ( .A(p_input[29155]), .B(p_input[19155]), .Z(n940) );
  AND U1881 ( .A(n941), .B(p_input[9154]), .Z(o[9154]) );
  AND U1882 ( .A(p_input[29154]), .B(p_input[19154]), .Z(n941) );
  AND U1883 ( .A(n942), .B(p_input[9153]), .Z(o[9153]) );
  AND U1884 ( .A(p_input[29153]), .B(p_input[19153]), .Z(n942) );
  AND U1885 ( .A(n943), .B(p_input[9152]), .Z(o[9152]) );
  AND U1886 ( .A(p_input[29152]), .B(p_input[19152]), .Z(n943) );
  AND U1887 ( .A(n944), .B(p_input[9151]), .Z(o[9151]) );
  AND U1888 ( .A(p_input[29151]), .B(p_input[19151]), .Z(n944) );
  AND U1889 ( .A(n945), .B(p_input[9150]), .Z(o[9150]) );
  AND U1890 ( .A(p_input[29150]), .B(p_input[19150]), .Z(n945) );
  AND U1891 ( .A(n946), .B(p_input[914]), .Z(o[914]) );
  AND U1892 ( .A(p_input[20914]), .B(p_input[10914]), .Z(n946) );
  AND U1893 ( .A(n947), .B(p_input[9149]), .Z(o[9149]) );
  AND U1894 ( .A(p_input[29149]), .B(p_input[19149]), .Z(n947) );
  AND U1895 ( .A(n948), .B(p_input[9148]), .Z(o[9148]) );
  AND U1896 ( .A(p_input[29148]), .B(p_input[19148]), .Z(n948) );
  AND U1897 ( .A(n949), .B(p_input[9147]), .Z(o[9147]) );
  AND U1898 ( .A(p_input[29147]), .B(p_input[19147]), .Z(n949) );
  AND U1899 ( .A(n950), .B(p_input[9146]), .Z(o[9146]) );
  AND U1900 ( .A(p_input[29146]), .B(p_input[19146]), .Z(n950) );
  AND U1901 ( .A(n951), .B(p_input[9145]), .Z(o[9145]) );
  AND U1902 ( .A(p_input[29145]), .B(p_input[19145]), .Z(n951) );
  AND U1903 ( .A(n952), .B(p_input[9144]), .Z(o[9144]) );
  AND U1904 ( .A(p_input[29144]), .B(p_input[19144]), .Z(n952) );
  AND U1905 ( .A(n953), .B(p_input[9143]), .Z(o[9143]) );
  AND U1906 ( .A(p_input[29143]), .B(p_input[19143]), .Z(n953) );
  AND U1907 ( .A(n954), .B(p_input[9142]), .Z(o[9142]) );
  AND U1908 ( .A(p_input[29142]), .B(p_input[19142]), .Z(n954) );
  AND U1909 ( .A(n955), .B(p_input[9141]), .Z(o[9141]) );
  AND U1910 ( .A(p_input[29141]), .B(p_input[19141]), .Z(n955) );
  AND U1911 ( .A(n956), .B(p_input[9140]), .Z(o[9140]) );
  AND U1912 ( .A(p_input[29140]), .B(p_input[19140]), .Z(n956) );
  AND U1913 ( .A(n957), .B(p_input[913]), .Z(o[913]) );
  AND U1914 ( .A(p_input[20913]), .B(p_input[10913]), .Z(n957) );
  AND U1915 ( .A(n958), .B(p_input[9139]), .Z(o[9139]) );
  AND U1916 ( .A(p_input[29139]), .B(p_input[19139]), .Z(n958) );
  AND U1917 ( .A(n959), .B(p_input[9138]), .Z(o[9138]) );
  AND U1918 ( .A(p_input[29138]), .B(p_input[19138]), .Z(n959) );
  AND U1919 ( .A(n960), .B(p_input[9137]), .Z(o[9137]) );
  AND U1920 ( .A(p_input[29137]), .B(p_input[19137]), .Z(n960) );
  AND U1921 ( .A(n961), .B(p_input[9136]), .Z(o[9136]) );
  AND U1922 ( .A(p_input[29136]), .B(p_input[19136]), .Z(n961) );
  AND U1923 ( .A(n962), .B(p_input[9135]), .Z(o[9135]) );
  AND U1924 ( .A(p_input[29135]), .B(p_input[19135]), .Z(n962) );
  AND U1925 ( .A(n963), .B(p_input[9134]), .Z(o[9134]) );
  AND U1926 ( .A(p_input[29134]), .B(p_input[19134]), .Z(n963) );
  AND U1927 ( .A(n964), .B(p_input[9133]), .Z(o[9133]) );
  AND U1928 ( .A(p_input[29133]), .B(p_input[19133]), .Z(n964) );
  AND U1929 ( .A(n965), .B(p_input[9132]), .Z(o[9132]) );
  AND U1930 ( .A(p_input[29132]), .B(p_input[19132]), .Z(n965) );
  AND U1931 ( .A(n966), .B(p_input[9131]), .Z(o[9131]) );
  AND U1932 ( .A(p_input[29131]), .B(p_input[19131]), .Z(n966) );
  AND U1933 ( .A(n967), .B(p_input[9130]), .Z(o[9130]) );
  AND U1934 ( .A(p_input[29130]), .B(p_input[19130]), .Z(n967) );
  AND U1935 ( .A(n968), .B(p_input[912]), .Z(o[912]) );
  AND U1936 ( .A(p_input[20912]), .B(p_input[10912]), .Z(n968) );
  AND U1937 ( .A(n969), .B(p_input[9129]), .Z(o[9129]) );
  AND U1938 ( .A(p_input[29129]), .B(p_input[19129]), .Z(n969) );
  AND U1939 ( .A(n970), .B(p_input[9128]), .Z(o[9128]) );
  AND U1940 ( .A(p_input[29128]), .B(p_input[19128]), .Z(n970) );
  AND U1941 ( .A(n971), .B(p_input[9127]), .Z(o[9127]) );
  AND U1942 ( .A(p_input[29127]), .B(p_input[19127]), .Z(n971) );
  AND U1943 ( .A(n972), .B(p_input[9126]), .Z(o[9126]) );
  AND U1944 ( .A(p_input[29126]), .B(p_input[19126]), .Z(n972) );
  AND U1945 ( .A(n973), .B(p_input[9125]), .Z(o[9125]) );
  AND U1946 ( .A(p_input[29125]), .B(p_input[19125]), .Z(n973) );
  AND U1947 ( .A(n974), .B(p_input[9124]), .Z(o[9124]) );
  AND U1948 ( .A(p_input[29124]), .B(p_input[19124]), .Z(n974) );
  AND U1949 ( .A(n975), .B(p_input[9123]), .Z(o[9123]) );
  AND U1950 ( .A(p_input[29123]), .B(p_input[19123]), .Z(n975) );
  AND U1951 ( .A(n976), .B(p_input[9122]), .Z(o[9122]) );
  AND U1952 ( .A(p_input[29122]), .B(p_input[19122]), .Z(n976) );
  AND U1953 ( .A(n977), .B(p_input[9121]), .Z(o[9121]) );
  AND U1954 ( .A(p_input[29121]), .B(p_input[19121]), .Z(n977) );
  AND U1955 ( .A(n978), .B(p_input[9120]), .Z(o[9120]) );
  AND U1956 ( .A(p_input[29120]), .B(p_input[19120]), .Z(n978) );
  AND U1957 ( .A(n979), .B(p_input[911]), .Z(o[911]) );
  AND U1958 ( .A(p_input[20911]), .B(p_input[10911]), .Z(n979) );
  AND U1959 ( .A(n980), .B(p_input[9119]), .Z(o[9119]) );
  AND U1960 ( .A(p_input[29119]), .B(p_input[19119]), .Z(n980) );
  AND U1961 ( .A(n981), .B(p_input[9118]), .Z(o[9118]) );
  AND U1962 ( .A(p_input[29118]), .B(p_input[19118]), .Z(n981) );
  AND U1963 ( .A(n982), .B(p_input[9117]), .Z(o[9117]) );
  AND U1964 ( .A(p_input[29117]), .B(p_input[19117]), .Z(n982) );
  AND U1965 ( .A(n983), .B(p_input[9116]), .Z(o[9116]) );
  AND U1966 ( .A(p_input[29116]), .B(p_input[19116]), .Z(n983) );
  AND U1967 ( .A(n984), .B(p_input[9115]), .Z(o[9115]) );
  AND U1968 ( .A(p_input[29115]), .B(p_input[19115]), .Z(n984) );
  AND U1969 ( .A(n985), .B(p_input[9114]), .Z(o[9114]) );
  AND U1970 ( .A(p_input[29114]), .B(p_input[19114]), .Z(n985) );
  AND U1971 ( .A(n986), .B(p_input[9113]), .Z(o[9113]) );
  AND U1972 ( .A(p_input[29113]), .B(p_input[19113]), .Z(n986) );
  AND U1973 ( .A(n987), .B(p_input[9112]), .Z(o[9112]) );
  AND U1974 ( .A(p_input[29112]), .B(p_input[19112]), .Z(n987) );
  AND U1975 ( .A(n988), .B(p_input[9111]), .Z(o[9111]) );
  AND U1976 ( .A(p_input[29111]), .B(p_input[19111]), .Z(n988) );
  AND U1977 ( .A(n989), .B(p_input[9110]), .Z(o[9110]) );
  AND U1978 ( .A(p_input[29110]), .B(p_input[19110]), .Z(n989) );
  AND U1979 ( .A(n990), .B(p_input[910]), .Z(o[910]) );
  AND U1980 ( .A(p_input[20910]), .B(p_input[10910]), .Z(n990) );
  AND U1981 ( .A(n991), .B(p_input[9109]), .Z(o[9109]) );
  AND U1982 ( .A(p_input[29109]), .B(p_input[19109]), .Z(n991) );
  AND U1983 ( .A(n992), .B(p_input[9108]), .Z(o[9108]) );
  AND U1984 ( .A(p_input[29108]), .B(p_input[19108]), .Z(n992) );
  AND U1985 ( .A(n993), .B(p_input[9107]), .Z(o[9107]) );
  AND U1986 ( .A(p_input[29107]), .B(p_input[19107]), .Z(n993) );
  AND U1987 ( .A(n994), .B(p_input[9106]), .Z(o[9106]) );
  AND U1988 ( .A(p_input[29106]), .B(p_input[19106]), .Z(n994) );
  AND U1989 ( .A(n995), .B(p_input[9105]), .Z(o[9105]) );
  AND U1990 ( .A(p_input[29105]), .B(p_input[19105]), .Z(n995) );
  AND U1991 ( .A(n996), .B(p_input[9104]), .Z(o[9104]) );
  AND U1992 ( .A(p_input[29104]), .B(p_input[19104]), .Z(n996) );
  AND U1993 ( .A(n997), .B(p_input[9103]), .Z(o[9103]) );
  AND U1994 ( .A(p_input[29103]), .B(p_input[19103]), .Z(n997) );
  AND U1995 ( .A(n998), .B(p_input[9102]), .Z(o[9102]) );
  AND U1996 ( .A(p_input[29102]), .B(p_input[19102]), .Z(n998) );
  AND U1997 ( .A(n999), .B(p_input[9101]), .Z(o[9101]) );
  AND U1998 ( .A(p_input[29101]), .B(p_input[19101]), .Z(n999) );
  AND U1999 ( .A(n1000), .B(p_input[9100]), .Z(o[9100]) );
  AND U2000 ( .A(p_input[29100]), .B(p_input[19100]), .Z(n1000) );
  AND U2001 ( .A(n1001), .B(p_input[90]), .Z(o[90]) );
  AND U2002 ( .A(p_input[20090]), .B(p_input[10090]), .Z(n1001) );
  AND U2003 ( .A(n1002), .B(p_input[909]), .Z(o[909]) );
  AND U2004 ( .A(p_input[20909]), .B(p_input[10909]), .Z(n1002) );
  AND U2005 ( .A(n1003), .B(p_input[9099]), .Z(o[9099]) );
  AND U2006 ( .A(p_input[29099]), .B(p_input[19099]), .Z(n1003) );
  AND U2007 ( .A(n1004), .B(p_input[9098]), .Z(o[9098]) );
  AND U2008 ( .A(p_input[29098]), .B(p_input[19098]), .Z(n1004) );
  AND U2009 ( .A(n1005), .B(p_input[9097]), .Z(o[9097]) );
  AND U2010 ( .A(p_input[29097]), .B(p_input[19097]), .Z(n1005) );
  AND U2011 ( .A(n1006), .B(p_input[9096]), .Z(o[9096]) );
  AND U2012 ( .A(p_input[29096]), .B(p_input[19096]), .Z(n1006) );
  AND U2013 ( .A(n1007), .B(p_input[9095]), .Z(o[9095]) );
  AND U2014 ( .A(p_input[29095]), .B(p_input[19095]), .Z(n1007) );
  AND U2015 ( .A(n1008), .B(p_input[9094]), .Z(o[9094]) );
  AND U2016 ( .A(p_input[29094]), .B(p_input[19094]), .Z(n1008) );
  AND U2017 ( .A(n1009), .B(p_input[9093]), .Z(o[9093]) );
  AND U2018 ( .A(p_input[29093]), .B(p_input[19093]), .Z(n1009) );
  AND U2019 ( .A(n1010), .B(p_input[9092]), .Z(o[9092]) );
  AND U2020 ( .A(p_input[29092]), .B(p_input[19092]), .Z(n1010) );
  AND U2021 ( .A(n1011), .B(p_input[9091]), .Z(o[9091]) );
  AND U2022 ( .A(p_input[29091]), .B(p_input[19091]), .Z(n1011) );
  AND U2023 ( .A(n1012), .B(p_input[9090]), .Z(o[9090]) );
  AND U2024 ( .A(p_input[29090]), .B(p_input[19090]), .Z(n1012) );
  AND U2025 ( .A(n1013), .B(p_input[908]), .Z(o[908]) );
  AND U2026 ( .A(p_input[20908]), .B(p_input[10908]), .Z(n1013) );
  AND U2027 ( .A(n1014), .B(p_input[9089]), .Z(o[9089]) );
  AND U2028 ( .A(p_input[29089]), .B(p_input[19089]), .Z(n1014) );
  AND U2029 ( .A(n1015), .B(p_input[9088]), .Z(o[9088]) );
  AND U2030 ( .A(p_input[29088]), .B(p_input[19088]), .Z(n1015) );
  AND U2031 ( .A(n1016), .B(p_input[9087]), .Z(o[9087]) );
  AND U2032 ( .A(p_input[29087]), .B(p_input[19087]), .Z(n1016) );
  AND U2033 ( .A(n1017), .B(p_input[9086]), .Z(o[9086]) );
  AND U2034 ( .A(p_input[29086]), .B(p_input[19086]), .Z(n1017) );
  AND U2035 ( .A(n1018), .B(p_input[9085]), .Z(o[9085]) );
  AND U2036 ( .A(p_input[29085]), .B(p_input[19085]), .Z(n1018) );
  AND U2037 ( .A(n1019), .B(p_input[9084]), .Z(o[9084]) );
  AND U2038 ( .A(p_input[29084]), .B(p_input[19084]), .Z(n1019) );
  AND U2039 ( .A(n1020), .B(p_input[9083]), .Z(o[9083]) );
  AND U2040 ( .A(p_input[29083]), .B(p_input[19083]), .Z(n1020) );
  AND U2041 ( .A(n1021), .B(p_input[9082]), .Z(o[9082]) );
  AND U2042 ( .A(p_input[29082]), .B(p_input[19082]), .Z(n1021) );
  AND U2043 ( .A(n1022), .B(p_input[9081]), .Z(o[9081]) );
  AND U2044 ( .A(p_input[29081]), .B(p_input[19081]), .Z(n1022) );
  AND U2045 ( .A(n1023), .B(p_input[9080]), .Z(o[9080]) );
  AND U2046 ( .A(p_input[29080]), .B(p_input[19080]), .Z(n1023) );
  AND U2047 ( .A(n1024), .B(p_input[907]), .Z(o[907]) );
  AND U2048 ( .A(p_input[20907]), .B(p_input[10907]), .Z(n1024) );
  AND U2049 ( .A(n1025), .B(p_input[9079]), .Z(o[9079]) );
  AND U2050 ( .A(p_input[29079]), .B(p_input[19079]), .Z(n1025) );
  AND U2051 ( .A(n1026), .B(p_input[9078]), .Z(o[9078]) );
  AND U2052 ( .A(p_input[29078]), .B(p_input[19078]), .Z(n1026) );
  AND U2053 ( .A(n1027), .B(p_input[9077]), .Z(o[9077]) );
  AND U2054 ( .A(p_input[29077]), .B(p_input[19077]), .Z(n1027) );
  AND U2055 ( .A(n1028), .B(p_input[9076]), .Z(o[9076]) );
  AND U2056 ( .A(p_input[29076]), .B(p_input[19076]), .Z(n1028) );
  AND U2057 ( .A(n1029), .B(p_input[9075]), .Z(o[9075]) );
  AND U2058 ( .A(p_input[29075]), .B(p_input[19075]), .Z(n1029) );
  AND U2059 ( .A(n1030), .B(p_input[9074]), .Z(o[9074]) );
  AND U2060 ( .A(p_input[29074]), .B(p_input[19074]), .Z(n1030) );
  AND U2061 ( .A(n1031), .B(p_input[9073]), .Z(o[9073]) );
  AND U2062 ( .A(p_input[29073]), .B(p_input[19073]), .Z(n1031) );
  AND U2063 ( .A(n1032), .B(p_input[9072]), .Z(o[9072]) );
  AND U2064 ( .A(p_input[29072]), .B(p_input[19072]), .Z(n1032) );
  AND U2065 ( .A(n1033), .B(p_input[9071]), .Z(o[9071]) );
  AND U2066 ( .A(p_input[29071]), .B(p_input[19071]), .Z(n1033) );
  AND U2067 ( .A(n1034), .B(p_input[9070]), .Z(o[9070]) );
  AND U2068 ( .A(p_input[29070]), .B(p_input[19070]), .Z(n1034) );
  AND U2069 ( .A(n1035), .B(p_input[906]), .Z(o[906]) );
  AND U2070 ( .A(p_input[20906]), .B(p_input[10906]), .Z(n1035) );
  AND U2071 ( .A(n1036), .B(p_input[9069]), .Z(o[9069]) );
  AND U2072 ( .A(p_input[29069]), .B(p_input[19069]), .Z(n1036) );
  AND U2073 ( .A(n1037), .B(p_input[9068]), .Z(o[9068]) );
  AND U2074 ( .A(p_input[29068]), .B(p_input[19068]), .Z(n1037) );
  AND U2075 ( .A(n1038), .B(p_input[9067]), .Z(o[9067]) );
  AND U2076 ( .A(p_input[29067]), .B(p_input[19067]), .Z(n1038) );
  AND U2077 ( .A(n1039), .B(p_input[9066]), .Z(o[9066]) );
  AND U2078 ( .A(p_input[29066]), .B(p_input[19066]), .Z(n1039) );
  AND U2079 ( .A(n1040), .B(p_input[9065]), .Z(o[9065]) );
  AND U2080 ( .A(p_input[29065]), .B(p_input[19065]), .Z(n1040) );
  AND U2081 ( .A(n1041), .B(p_input[9064]), .Z(o[9064]) );
  AND U2082 ( .A(p_input[29064]), .B(p_input[19064]), .Z(n1041) );
  AND U2083 ( .A(n1042), .B(p_input[9063]), .Z(o[9063]) );
  AND U2084 ( .A(p_input[29063]), .B(p_input[19063]), .Z(n1042) );
  AND U2085 ( .A(n1043), .B(p_input[9062]), .Z(o[9062]) );
  AND U2086 ( .A(p_input[29062]), .B(p_input[19062]), .Z(n1043) );
  AND U2087 ( .A(n1044), .B(p_input[9061]), .Z(o[9061]) );
  AND U2088 ( .A(p_input[29061]), .B(p_input[19061]), .Z(n1044) );
  AND U2089 ( .A(n1045), .B(p_input[9060]), .Z(o[9060]) );
  AND U2090 ( .A(p_input[29060]), .B(p_input[19060]), .Z(n1045) );
  AND U2091 ( .A(n1046), .B(p_input[905]), .Z(o[905]) );
  AND U2092 ( .A(p_input[20905]), .B(p_input[10905]), .Z(n1046) );
  AND U2093 ( .A(n1047), .B(p_input[9059]), .Z(o[9059]) );
  AND U2094 ( .A(p_input[29059]), .B(p_input[19059]), .Z(n1047) );
  AND U2095 ( .A(n1048), .B(p_input[9058]), .Z(o[9058]) );
  AND U2096 ( .A(p_input[29058]), .B(p_input[19058]), .Z(n1048) );
  AND U2097 ( .A(n1049), .B(p_input[9057]), .Z(o[9057]) );
  AND U2098 ( .A(p_input[29057]), .B(p_input[19057]), .Z(n1049) );
  AND U2099 ( .A(n1050), .B(p_input[9056]), .Z(o[9056]) );
  AND U2100 ( .A(p_input[29056]), .B(p_input[19056]), .Z(n1050) );
  AND U2101 ( .A(n1051), .B(p_input[9055]), .Z(o[9055]) );
  AND U2102 ( .A(p_input[29055]), .B(p_input[19055]), .Z(n1051) );
  AND U2103 ( .A(n1052), .B(p_input[9054]), .Z(o[9054]) );
  AND U2104 ( .A(p_input[29054]), .B(p_input[19054]), .Z(n1052) );
  AND U2105 ( .A(n1053), .B(p_input[9053]), .Z(o[9053]) );
  AND U2106 ( .A(p_input[29053]), .B(p_input[19053]), .Z(n1053) );
  AND U2107 ( .A(n1054), .B(p_input[9052]), .Z(o[9052]) );
  AND U2108 ( .A(p_input[29052]), .B(p_input[19052]), .Z(n1054) );
  AND U2109 ( .A(n1055), .B(p_input[9051]), .Z(o[9051]) );
  AND U2110 ( .A(p_input[29051]), .B(p_input[19051]), .Z(n1055) );
  AND U2111 ( .A(n1056), .B(p_input[9050]), .Z(o[9050]) );
  AND U2112 ( .A(p_input[29050]), .B(p_input[19050]), .Z(n1056) );
  AND U2113 ( .A(n1057), .B(p_input[904]), .Z(o[904]) );
  AND U2114 ( .A(p_input[20904]), .B(p_input[10904]), .Z(n1057) );
  AND U2115 ( .A(n1058), .B(p_input[9049]), .Z(o[9049]) );
  AND U2116 ( .A(p_input[29049]), .B(p_input[19049]), .Z(n1058) );
  AND U2117 ( .A(n1059), .B(p_input[9048]), .Z(o[9048]) );
  AND U2118 ( .A(p_input[29048]), .B(p_input[19048]), .Z(n1059) );
  AND U2119 ( .A(n1060), .B(p_input[9047]), .Z(o[9047]) );
  AND U2120 ( .A(p_input[29047]), .B(p_input[19047]), .Z(n1060) );
  AND U2121 ( .A(n1061), .B(p_input[9046]), .Z(o[9046]) );
  AND U2122 ( .A(p_input[29046]), .B(p_input[19046]), .Z(n1061) );
  AND U2123 ( .A(n1062), .B(p_input[9045]), .Z(o[9045]) );
  AND U2124 ( .A(p_input[29045]), .B(p_input[19045]), .Z(n1062) );
  AND U2125 ( .A(n1063), .B(p_input[9044]), .Z(o[9044]) );
  AND U2126 ( .A(p_input[29044]), .B(p_input[19044]), .Z(n1063) );
  AND U2127 ( .A(n1064), .B(p_input[9043]), .Z(o[9043]) );
  AND U2128 ( .A(p_input[29043]), .B(p_input[19043]), .Z(n1064) );
  AND U2129 ( .A(n1065), .B(p_input[9042]), .Z(o[9042]) );
  AND U2130 ( .A(p_input[29042]), .B(p_input[19042]), .Z(n1065) );
  AND U2131 ( .A(n1066), .B(p_input[9041]), .Z(o[9041]) );
  AND U2132 ( .A(p_input[29041]), .B(p_input[19041]), .Z(n1066) );
  AND U2133 ( .A(n1067), .B(p_input[9040]), .Z(o[9040]) );
  AND U2134 ( .A(p_input[29040]), .B(p_input[19040]), .Z(n1067) );
  AND U2135 ( .A(n1068), .B(p_input[903]), .Z(o[903]) );
  AND U2136 ( .A(p_input[20903]), .B(p_input[10903]), .Z(n1068) );
  AND U2137 ( .A(n1069), .B(p_input[9039]), .Z(o[9039]) );
  AND U2138 ( .A(p_input[29039]), .B(p_input[19039]), .Z(n1069) );
  AND U2139 ( .A(n1070), .B(p_input[9038]), .Z(o[9038]) );
  AND U2140 ( .A(p_input[29038]), .B(p_input[19038]), .Z(n1070) );
  AND U2141 ( .A(n1071), .B(p_input[9037]), .Z(o[9037]) );
  AND U2142 ( .A(p_input[29037]), .B(p_input[19037]), .Z(n1071) );
  AND U2143 ( .A(n1072), .B(p_input[9036]), .Z(o[9036]) );
  AND U2144 ( .A(p_input[29036]), .B(p_input[19036]), .Z(n1072) );
  AND U2145 ( .A(n1073), .B(p_input[9035]), .Z(o[9035]) );
  AND U2146 ( .A(p_input[29035]), .B(p_input[19035]), .Z(n1073) );
  AND U2147 ( .A(n1074), .B(p_input[9034]), .Z(o[9034]) );
  AND U2148 ( .A(p_input[29034]), .B(p_input[19034]), .Z(n1074) );
  AND U2149 ( .A(n1075), .B(p_input[9033]), .Z(o[9033]) );
  AND U2150 ( .A(p_input[29033]), .B(p_input[19033]), .Z(n1075) );
  AND U2151 ( .A(n1076), .B(p_input[9032]), .Z(o[9032]) );
  AND U2152 ( .A(p_input[29032]), .B(p_input[19032]), .Z(n1076) );
  AND U2153 ( .A(n1077), .B(p_input[9031]), .Z(o[9031]) );
  AND U2154 ( .A(p_input[29031]), .B(p_input[19031]), .Z(n1077) );
  AND U2155 ( .A(n1078), .B(p_input[9030]), .Z(o[9030]) );
  AND U2156 ( .A(p_input[29030]), .B(p_input[19030]), .Z(n1078) );
  AND U2157 ( .A(n1079), .B(p_input[902]), .Z(o[902]) );
  AND U2158 ( .A(p_input[20902]), .B(p_input[10902]), .Z(n1079) );
  AND U2159 ( .A(n1080), .B(p_input[9029]), .Z(o[9029]) );
  AND U2160 ( .A(p_input[29029]), .B(p_input[19029]), .Z(n1080) );
  AND U2161 ( .A(n1081), .B(p_input[9028]), .Z(o[9028]) );
  AND U2162 ( .A(p_input[29028]), .B(p_input[19028]), .Z(n1081) );
  AND U2163 ( .A(n1082), .B(p_input[9027]), .Z(o[9027]) );
  AND U2164 ( .A(p_input[29027]), .B(p_input[19027]), .Z(n1082) );
  AND U2165 ( .A(n1083), .B(p_input[9026]), .Z(o[9026]) );
  AND U2166 ( .A(p_input[29026]), .B(p_input[19026]), .Z(n1083) );
  AND U2167 ( .A(n1084), .B(p_input[9025]), .Z(o[9025]) );
  AND U2168 ( .A(p_input[29025]), .B(p_input[19025]), .Z(n1084) );
  AND U2169 ( .A(n1085), .B(p_input[9024]), .Z(o[9024]) );
  AND U2170 ( .A(p_input[29024]), .B(p_input[19024]), .Z(n1085) );
  AND U2171 ( .A(n1086), .B(p_input[9023]), .Z(o[9023]) );
  AND U2172 ( .A(p_input[29023]), .B(p_input[19023]), .Z(n1086) );
  AND U2173 ( .A(n1087), .B(p_input[9022]), .Z(o[9022]) );
  AND U2174 ( .A(p_input[29022]), .B(p_input[19022]), .Z(n1087) );
  AND U2175 ( .A(n1088), .B(p_input[9021]), .Z(o[9021]) );
  AND U2176 ( .A(p_input[29021]), .B(p_input[19021]), .Z(n1088) );
  AND U2177 ( .A(n1089), .B(p_input[9020]), .Z(o[9020]) );
  AND U2178 ( .A(p_input[29020]), .B(p_input[19020]), .Z(n1089) );
  AND U2179 ( .A(n1090), .B(p_input[901]), .Z(o[901]) );
  AND U2180 ( .A(p_input[20901]), .B(p_input[10901]), .Z(n1090) );
  AND U2181 ( .A(n1091), .B(p_input[9019]), .Z(o[9019]) );
  AND U2182 ( .A(p_input[29019]), .B(p_input[19019]), .Z(n1091) );
  AND U2183 ( .A(n1092), .B(p_input[9018]), .Z(o[9018]) );
  AND U2184 ( .A(p_input[29018]), .B(p_input[19018]), .Z(n1092) );
  AND U2185 ( .A(n1093), .B(p_input[9017]), .Z(o[9017]) );
  AND U2186 ( .A(p_input[29017]), .B(p_input[19017]), .Z(n1093) );
  AND U2187 ( .A(n1094), .B(p_input[9016]), .Z(o[9016]) );
  AND U2188 ( .A(p_input[29016]), .B(p_input[19016]), .Z(n1094) );
  AND U2189 ( .A(n1095), .B(p_input[9015]), .Z(o[9015]) );
  AND U2190 ( .A(p_input[29015]), .B(p_input[19015]), .Z(n1095) );
  AND U2191 ( .A(n1096), .B(p_input[9014]), .Z(o[9014]) );
  AND U2192 ( .A(p_input[29014]), .B(p_input[19014]), .Z(n1096) );
  AND U2193 ( .A(n1097), .B(p_input[9013]), .Z(o[9013]) );
  AND U2194 ( .A(p_input[29013]), .B(p_input[19013]), .Z(n1097) );
  AND U2195 ( .A(n1098), .B(p_input[9012]), .Z(o[9012]) );
  AND U2196 ( .A(p_input[29012]), .B(p_input[19012]), .Z(n1098) );
  AND U2197 ( .A(n1099), .B(p_input[9011]), .Z(o[9011]) );
  AND U2198 ( .A(p_input[29011]), .B(p_input[19011]), .Z(n1099) );
  AND U2199 ( .A(n1100), .B(p_input[9010]), .Z(o[9010]) );
  AND U2200 ( .A(p_input[29010]), .B(p_input[19010]), .Z(n1100) );
  AND U2201 ( .A(n1101), .B(p_input[900]), .Z(o[900]) );
  AND U2202 ( .A(p_input[20900]), .B(p_input[10900]), .Z(n1101) );
  AND U2203 ( .A(n1102), .B(p_input[9009]), .Z(o[9009]) );
  AND U2204 ( .A(p_input[29009]), .B(p_input[19009]), .Z(n1102) );
  AND U2205 ( .A(n1103), .B(p_input[9008]), .Z(o[9008]) );
  AND U2206 ( .A(p_input[29008]), .B(p_input[19008]), .Z(n1103) );
  AND U2207 ( .A(n1104), .B(p_input[9007]), .Z(o[9007]) );
  AND U2208 ( .A(p_input[29007]), .B(p_input[19007]), .Z(n1104) );
  AND U2209 ( .A(n1105), .B(p_input[9006]), .Z(o[9006]) );
  AND U2210 ( .A(p_input[29006]), .B(p_input[19006]), .Z(n1105) );
  AND U2211 ( .A(n1106), .B(p_input[9005]), .Z(o[9005]) );
  AND U2212 ( .A(p_input[29005]), .B(p_input[19005]), .Z(n1106) );
  AND U2213 ( .A(n1107), .B(p_input[9004]), .Z(o[9004]) );
  AND U2214 ( .A(p_input[29004]), .B(p_input[19004]), .Z(n1107) );
  AND U2215 ( .A(n1108), .B(p_input[9003]), .Z(o[9003]) );
  AND U2216 ( .A(p_input[29003]), .B(p_input[19003]), .Z(n1108) );
  AND U2217 ( .A(n1109), .B(p_input[9002]), .Z(o[9002]) );
  AND U2218 ( .A(p_input[29002]), .B(p_input[19002]), .Z(n1109) );
  AND U2219 ( .A(n1110), .B(p_input[9001]), .Z(o[9001]) );
  AND U2220 ( .A(p_input[29001]), .B(p_input[19001]), .Z(n1110) );
  AND U2221 ( .A(n1111), .B(p_input[9000]), .Z(o[9000]) );
  AND U2222 ( .A(p_input[29000]), .B(p_input[19000]), .Z(n1111) );
  AND U2223 ( .A(n1112), .B(p_input[8]), .Z(o[8]) );
  AND U2224 ( .A(p_input[20008]), .B(p_input[10008]), .Z(n1112) );
  AND U2225 ( .A(n1113), .B(p_input[89]), .Z(o[89]) );
  AND U2226 ( .A(p_input[20089]), .B(p_input[10089]), .Z(n1113) );
  AND U2227 ( .A(n1114), .B(p_input[899]), .Z(o[899]) );
  AND U2228 ( .A(p_input[20899]), .B(p_input[10899]), .Z(n1114) );
  AND U2229 ( .A(n1115), .B(p_input[8999]), .Z(o[8999]) );
  AND U2230 ( .A(p_input[28999]), .B(p_input[18999]), .Z(n1115) );
  AND U2231 ( .A(n1116), .B(p_input[8998]), .Z(o[8998]) );
  AND U2232 ( .A(p_input[28998]), .B(p_input[18998]), .Z(n1116) );
  AND U2233 ( .A(n1117), .B(p_input[8997]), .Z(o[8997]) );
  AND U2234 ( .A(p_input[28997]), .B(p_input[18997]), .Z(n1117) );
  AND U2235 ( .A(n1118), .B(p_input[8996]), .Z(o[8996]) );
  AND U2236 ( .A(p_input[28996]), .B(p_input[18996]), .Z(n1118) );
  AND U2237 ( .A(n1119), .B(p_input[8995]), .Z(o[8995]) );
  AND U2238 ( .A(p_input[28995]), .B(p_input[18995]), .Z(n1119) );
  AND U2239 ( .A(n1120), .B(p_input[8994]), .Z(o[8994]) );
  AND U2240 ( .A(p_input[28994]), .B(p_input[18994]), .Z(n1120) );
  AND U2241 ( .A(n1121), .B(p_input[8993]), .Z(o[8993]) );
  AND U2242 ( .A(p_input[28993]), .B(p_input[18993]), .Z(n1121) );
  AND U2243 ( .A(n1122), .B(p_input[8992]), .Z(o[8992]) );
  AND U2244 ( .A(p_input[28992]), .B(p_input[18992]), .Z(n1122) );
  AND U2245 ( .A(n1123), .B(p_input[8991]), .Z(o[8991]) );
  AND U2246 ( .A(p_input[28991]), .B(p_input[18991]), .Z(n1123) );
  AND U2247 ( .A(n1124), .B(p_input[8990]), .Z(o[8990]) );
  AND U2248 ( .A(p_input[28990]), .B(p_input[18990]), .Z(n1124) );
  AND U2249 ( .A(n1125), .B(p_input[898]), .Z(o[898]) );
  AND U2250 ( .A(p_input[20898]), .B(p_input[10898]), .Z(n1125) );
  AND U2251 ( .A(n1126), .B(p_input[8989]), .Z(o[8989]) );
  AND U2252 ( .A(p_input[28989]), .B(p_input[18989]), .Z(n1126) );
  AND U2253 ( .A(n1127), .B(p_input[8988]), .Z(o[8988]) );
  AND U2254 ( .A(p_input[28988]), .B(p_input[18988]), .Z(n1127) );
  AND U2255 ( .A(n1128), .B(p_input[8987]), .Z(o[8987]) );
  AND U2256 ( .A(p_input[28987]), .B(p_input[18987]), .Z(n1128) );
  AND U2257 ( .A(n1129), .B(p_input[8986]), .Z(o[8986]) );
  AND U2258 ( .A(p_input[28986]), .B(p_input[18986]), .Z(n1129) );
  AND U2259 ( .A(n1130), .B(p_input[8985]), .Z(o[8985]) );
  AND U2260 ( .A(p_input[28985]), .B(p_input[18985]), .Z(n1130) );
  AND U2261 ( .A(n1131), .B(p_input[8984]), .Z(o[8984]) );
  AND U2262 ( .A(p_input[28984]), .B(p_input[18984]), .Z(n1131) );
  AND U2263 ( .A(n1132), .B(p_input[8983]), .Z(o[8983]) );
  AND U2264 ( .A(p_input[28983]), .B(p_input[18983]), .Z(n1132) );
  AND U2265 ( .A(n1133), .B(p_input[8982]), .Z(o[8982]) );
  AND U2266 ( .A(p_input[28982]), .B(p_input[18982]), .Z(n1133) );
  AND U2267 ( .A(n1134), .B(p_input[8981]), .Z(o[8981]) );
  AND U2268 ( .A(p_input[28981]), .B(p_input[18981]), .Z(n1134) );
  AND U2269 ( .A(n1135), .B(p_input[8980]), .Z(o[8980]) );
  AND U2270 ( .A(p_input[28980]), .B(p_input[18980]), .Z(n1135) );
  AND U2271 ( .A(n1136), .B(p_input[897]), .Z(o[897]) );
  AND U2272 ( .A(p_input[20897]), .B(p_input[10897]), .Z(n1136) );
  AND U2273 ( .A(n1137), .B(p_input[8979]), .Z(o[8979]) );
  AND U2274 ( .A(p_input[28979]), .B(p_input[18979]), .Z(n1137) );
  AND U2275 ( .A(n1138), .B(p_input[8978]), .Z(o[8978]) );
  AND U2276 ( .A(p_input[28978]), .B(p_input[18978]), .Z(n1138) );
  AND U2277 ( .A(n1139), .B(p_input[8977]), .Z(o[8977]) );
  AND U2278 ( .A(p_input[28977]), .B(p_input[18977]), .Z(n1139) );
  AND U2279 ( .A(n1140), .B(p_input[8976]), .Z(o[8976]) );
  AND U2280 ( .A(p_input[28976]), .B(p_input[18976]), .Z(n1140) );
  AND U2281 ( .A(n1141), .B(p_input[8975]), .Z(o[8975]) );
  AND U2282 ( .A(p_input[28975]), .B(p_input[18975]), .Z(n1141) );
  AND U2283 ( .A(n1142), .B(p_input[8974]), .Z(o[8974]) );
  AND U2284 ( .A(p_input[28974]), .B(p_input[18974]), .Z(n1142) );
  AND U2285 ( .A(n1143), .B(p_input[8973]), .Z(o[8973]) );
  AND U2286 ( .A(p_input[28973]), .B(p_input[18973]), .Z(n1143) );
  AND U2287 ( .A(n1144), .B(p_input[8972]), .Z(o[8972]) );
  AND U2288 ( .A(p_input[28972]), .B(p_input[18972]), .Z(n1144) );
  AND U2289 ( .A(n1145), .B(p_input[8971]), .Z(o[8971]) );
  AND U2290 ( .A(p_input[28971]), .B(p_input[18971]), .Z(n1145) );
  AND U2291 ( .A(n1146), .B(p_input[8970]), .Z(o[8970]) );
  AND U2292 ( .A(p_input[28970]), .B(p_input[18970]), .Z(n1146) );
  AND U2293 ( .A(n1147), .B(p_input[896]), .Z(o[896]) );
  AND U2294 ( .A(p_input[20896]), .B(p_input[10896]), .Z(n1147) );
  AND U2295 ( .A(n1148), .B(p_input[8969]), .Z(o[8969]) );
  AND U2296 ( .A(p_input[28969]), .B(p_input[18969]), .Z(n1148) );
  AND U2297 ( .A(n1149), .B(p_input[8968]), .Z(o[8968]) );
  AND U2298 ( .A(p_input[28968]), .B(p_input[18968]), .Z(n1149) );
  AND U2299 ( .A(n1150), .B(p_input[8967]), .Z(o[8967]) );
  AND U2300 ( .A(p_input[28967]), .B(p_input[18967]), .Z(n1150) );
  AND U2301 ( .A(n1151), .B(p_input[8966]), .Z(o[8966]) );
  AND U2302 ( .A(p_input[28966]), .B(p_input[18966]), .Z(n1151) );
  AND U2303 ( .A(n1152), .B(p_input[8965]), .Z(o[8965]) );
  AND U2304 ( .A(p_input[28965]), .B(p_input[18965]), .Z(n1152) );
  AND U2305 ( .A(n1153), .B(p_input[8964]), .Z(o[8964]) );
  AND U2306 ( .A(p_input[28964]), .B(p_input[18964]), .Z(n1153) );
  AND U2307 ( .A(n1154), .B(p_input[8963]), .Z(o[8963]) );
  AND U2308 ( .A(p_input[28963]), .B(p_input[18963]), .Z(n1154) );
  AND U2309 ( .A(n1155), .B(p_input[8962]), .Z(o[8962]) );
  AND U2310 ( .A(p_input[28962]), .B(p_input[18962]), .Z(n1155) );
  AND U2311 ( .A(n1156), .B(p_input[8961]), .Z(o[8961]) );
  AND U2312 ( .A(p_input[28961]), .B(p_input[18961]), .Z(n1156) );
  AND U2313 ( .A(n1157), .B(p_input[8960]), .Z(o[8960]) );
  AND U2314 ( .A(p_input[28960]), .B(p_input[18960]), .Z(n1157) );
  AND U2315 ( .A(n1158), .B(p_input[895]), .Z(o[895]) );
  AND U2316 ( .A(p_input[20895]), .B(p_input[10895]), .Z(n1158) );
  AND U2317 ( .A(n1159), .B(p_input[8959]), .Z(o[8959]) );
  AND U2318 ( .A(p_input[28959]), .B(p_input[18959]), .Z(n1159) );
  AND U2319 ( .A(n1160), .B(p_input[8958]), .Z(o[8958]) );
  AND U2320 ( .A(p_input[28958]), .B(p_input[18958]), .Z(n1160) );
  AND U2321 ( .A(n1161), .B(p_input[8957]), .Z(o[8957]) );
  AND U2322 ( .A(p_input[28957]), .B(p_input[18957]), .Z(n1161) );
  AND U2323 ( .A(n1162), .B(p_input[8956]), .Z(o[8956]) );
  AND U2324 ( .A(p_input[28956]), .B(p_input[18956]), .Z(n1162) );
  AND U2325 ( .A(n1163), .B(p_input[8955]), .Z(o[8955]) );
  AND U2326 ( .A(p_input[28955]), .B(p_input[18955]), .Z(n1163) );
  AND U2327 ( .A(n1164), .B(p_input[8954]), .Z(o[8954]) );
  AND U2328 ( .A(p_input[28954]), .B(p_input[18954]), .Z(n1164) );
  AND U2329 ( .A(n1165), .B(p_input[8953]), .Z(o[8953]) );
  AND U2330 ( .A(p_input[28953]), .B(p_input[18953]), .Z(n1165) );
  AND U2331 ( .A(n1166), .B(p_input[8952]), .Z(o[8952]) );
  AND U2332 ( .A(p_input[28952]), .B(p_input[18952]), .Z(n1166) );
  AND U2333 ( .A(n1167), .B(p_input[8951]), .Z(o[8951]) );
  AND U2334 ( .A(p_input[28951]), .B(p_input[18951]), .Z(n1167) );
  AND U2335 ( .A(n1168), .B(p_input[8950]), .Z(o[8950]) );
  AND U2336 ( .A(p_input[28950]), .B(p_input[18950]), .Z(n1168) );
  AND U2337 ( .A(n1169), .B(p_input[894]), .Z(o[894]) );
  AND U2338 ( .A(p_input[20894]), .B(p_input[10894]), .Z(n1169) );
  AND U2339 ( .A(n1170), .B(p_input[8949]), .Z(o[8949]) );
  AND U2340 ( .A(p_input[28949]), .B(p_input[18949]), .Z(n1170) );
  AND U2341 ( .A(n1171), .B(p_input[8948]), .Z(o[8948]) );
  AND U2342 ( .A(p_input[28948]), .B(p_input[18948]), .Z(n1171) );
  AND U2343 ( .A(n1172), .B(p_input[8947]), .Z(o[8947]) );
  AND U2344 ( .A(p_input[28947]), .B(p_input[18947]), .Z(n1172) );
  AND U2345 ( .A(n1173), .B(p_input[8946]), .Z(o[8946]) );
  AND U2346 ( .A(p_input[28946]), .B(p_input[18946]), .Z(n1173) );
  AND U2347 ( .A(n1174), .B(p_input[8945]), .Z(o[8945]) );
  AND U2348 ( .A(p_input[28945]), .B(p_input[18945]), .Z(n1174) );
  AND U2349 ( .A(n1175), .B(p_input[8944]), .Z(o[8944]) );
  AND U2350 ( .A(p_input[28944]), .B(p_input[18944]), .Z(n1175) );
  AND U2351 ( .A(n1176), .B(p_input[8943]), .Z(o[8943]) );
  AND U2352 ( .A(p_input[28943]), .B(p_input[18943]), .Z(n1176) );
  AND U2353 ( .A(n1177), .B(p_input[8942]), .Z(o[8942]) );
  AND U2354 ( .A(p_input[28942]), .B(p_input[18942]), .Z(n1177) );
  AND U2355 ( .A(n1178), .B(p_input[8941]), .Z(o[8941]) );
  AND U2356 ( .A(p_input[28941]), .B(p_input[18941]), .Z(n1178) );
  AND U2357 ( .A(n1179), .B(p_input[8940]), .Z(o[8940]) );
  AND U2358 ( .A(p_input[28940]), .B(p_input[18940]), .Z(n1179) );
  AND U2359 ( .A(n1180), .B(p_input[893]), .Z(o[893]) );
  AND U2360 ( .A(p_input[20893]), .B(p_input[10893]), .Z(n1180) );
  AND U2361 ( .A(n1181), .B(p_input[8939]), .Z(o[8939]) );
  AND U2362 ( .A(p_input[28939]), .B(p_input[18939]), .Z(n1181) );
  AND U2363 ( .A(n1182), .B(p_input[8938]), .Z(o[8938]) );
  AND U2364 ( .A(p_input[28938]), .B(p_input[18938]), .Z(n1182) );
  AND U2365 ( .A(n1183), .B(p_input[8937]), .Z(o[8937]) );
  AND U2366 ( .A(p_input[28937]), .B(p_input[18937]), .Z(n1183) );
  AND U2367 ( .A(n1184), .B(p_input[8936]), .Z(o[8936]) );
  AND U2368 ( .A(p_input[28936]), .B(p_input[18936]), .Z(n1184) );
  AND U2369 ( .A(n1185), .B(p_input[8935]), .Z(o[8935]) );
  AND U2370 ( .A(p_input[28935]), .B(p_input[18935]), .Z(n1185) );
  AND U2371 ( .A(n1186), .B(p_input[8934]), .Z(o[8934]) );
  AND U2372 ( .A(p_input[28934]), .B(p_input[18934]), .Z(n1186) );
  AND U2373 ( .A(n1187), .B(p_input[8933]), .Z(o[8933]) );
  AND U2374 ( .A(p_input[28933]), .B(p_input[18933]), .Z(n1187) );
  AND U2375 ( .A(n1188), .B(p_input[8932]), .Z(o[8932]) );
  AND U2376 ( .A(p_input[28932]), .B(p_input[18932]), .Z(n1188) );
  AND U2377 ( .A(n1189), .B(p_input[8931]), .Z(o[8931]) );
  AND U2378 ( .A(p_input[28931]), .B(p_input[18931]), .Z(n1189) );
  AND U2379 ( .A(n1190), .B(p_input[8930]), .Z(o[8930]) );
  AND U2380 ( .A(p_input[28930]), .B(p_input[18930]), .Z(n1190) );
  AND U2381 ( .A(n1191), .B(p_input[892]), .Z(o[892]) );
  AND U2382 ( .A(p_input[20892]), .B(p_input[10892]), .Z(n1191) );
  AND U2383 ( .A(n1192), .B(p_input[8929]), .Z(o[8929]) );
  AND U2384 ( .A(p_input[28929]), .B(p_input[18929]), .Z(n1192) );
  AND U2385 ( .A(n1193), .B(p_input[8928]), .Z(o[8928]) );
  AND U2386 ( .A(p_input[28928]), .B(p_input[18928]), .Z(n1193) );
  AND U2387 ( .A(n1194), .B(p_input[8927]), .Z(o[8927]) );
  AND U2388 ( .A(p_input[28927]), .B(p_input[18927]), .Z(n1194) );
  AND U2389 ( .A(n1195), .B(p_input[8926]), .Z(o[8926]) );
  AND U2390 ( .A(p_input[28926]), .B(p_input[18926]), .Z(n1195) );
  AND U2391 ( .A(n1196), .B(p_input[8925]), .Z(o[8925]) );
  AND U2392 ( .A(p_input[28925]), .B(p_input[18925]), .Z(n1196) );
  AND U2393 ( .A(n1197), .B(p_input[8924]), .Z(o[8924]) );
  AND U2394 ( .A(p_input[28924]), .B(p_input[18924]), .Z(n1197) );
  AND U2395 ( .A(n1198), .B(p_input[8923]), .Z(o[8923]) );
  AND U2396 ( .A(p_input[28923]), .B(p_input[18923]), .Z(n1198) );
  AND U2397 ( .A(n1199), .B(p_input[8922]), .Z(o[8922]) );
  AND U2398 ( .A(p_input[28922]), .B(p_input[18922]), .Z(n1199) );
  AND U2399 ( .A(n1200), .B(p_input[8921]), .Z(o[8921]) );
  AND U2400 ( .A(p_input[28921]), .B(p_input[18921]), .Z(n1200) );
  AND U2401 ( .A(n1201), .B(p_input[8920]), .Z(o[8920]) );
  AND U2402 ( .A(p_input[28920]), .B(p_input[18920]), .Z(n1201) );
  AND U2403 ( .A(n1202), .B(p_input[891]), .Z(o[891]) );
  AND U2404 ( .A(p_input[20891]), .B(p_input[10891]), .Z(n1202) );
  AND U2405 ( .A(n1203), .B(p_input[8919]), .Z(o[8919]) );
  AND U2406 ( .A(p_input[28919]), .B(p_input[18919]), .Z(n1203) );
  AND U2407 ( .A(n1204), .B(p_input[8918]), .Z(o[8918]) );
  AND U2408 ( .A(p_input[28918]), .B(p_input[18918]), .Z(n1204) );
  AND U2409 ( .A(n1205), .B(p_input[8917]), .Z(o[8917]) );
  AND U2410 ( .A(p_input[28917]), .B(p_input[18917]), .Z(n1205) );
  AND U2411 ( .A(n1206), .B(p_input[8916]), .Z(o[8916]) );
  AND U2412 ( .A(p_input[28916]), .B(p_input[18916]), .Z(n1206) );
  AND U2413 ( .A(n1207), .B(p_input[8915]), .Z(o[8915]) );
  AND U2414 ( .A(p_input[28915]), .B(p_input[18915]), .Z(n1207) );
  AND U2415 ( .A(n1208), .B(p_input[8914]), .Z(o[8914]) );
  AND U2416 ( .A(p_input[28914]), .B(p_input[18914]), .Z(n1208) );
  AND U2417 ( .A(n1209), .B(p_input[8913]), .Z(o[8913]) );
  AND U2418 ( .A(p_input[28913]), .B(p_input[18913]), .Z(n1209) );
  AND U2419 ( .A(n1210), .B(p_input[8912]), .Z(o[8912]) );
  AND U2420 ( .A(p_input[28912]), .B(p_input[18912]), .Z(n1210) );
  AND U2421 ( .A(n1211), .B(p_input[8911]), .Z(o[8911]) );
  AND U2422 ( .A(p_input[28911]), .B(p_input[18911]), .Z(n1211) );
  AND U2423 ( .A(n1212), .B(p_input[8910]), .Z(o[8910]) );
  AND U2424 ( .A(p_input[28910]), .B(p_input[18910]), .Z(n1212) );
  AND U2425 ( .A(n1213), .B(p_input[890]), .Z(o[890]) );
  AND U2426 ( .A(p_input[20890]), .B(p_input[10890]), .Z(n1213) );
  AND U2427 ( .A(n1214), .B(p_input[8909]), .Z(o[8909]) );
  AND U2428 ( .A(p_input[28909]), .B(p_input[18909]), .Z(n1214) );
  AND U2429 ( .A(n1215), .B(p_input[8908]), .Z(o[8908]) );
  AND U2430 ( .A(p_input[28908]), .B(p_input[18908]), .Z(n1215) );
  AND U2431 ( .A(n1216), .B(p_input[8907]), .Z(o[8907]) );
  AND U2432 ( .A(p_input[28907]), .B(p_input[18907]), .Z(n1216) );
  AND U2433 ( .A(n1217), .B(p_input[8906]), .Z(o[8906]) );
  AND U2434 ( .A(p_input[28906]), .B(p_input[18906]), .Z(n1217) );
  AND U2435 ( .A(n1218), .B(p_input[8905]), .Z(o[8905]) );
  AND U2436 ( .A(p_input[28905]), .B(p_input[18905]), .Z(n1218) );
  AND U2437 ( .A(n1219), .B(p_input[8904]), .Z(o[8904]) );
  AND U2438 ( .A(p_input[28904]), .B(p_input[18904]), .Z(n1219) );
  AND U2439 ( .A(n1220), .B(p_input[8903]), .Z(o[8903]) );
  AND U2440 ( .A(p_input[28903]), .B(p_input[18903]), .Z(n1220) );
  AND U2441 ( .A(n1221), .B(p_input[8902]), .Z(o[8902]) );
  AND U2442 ( .A(p_input[28902]), .B(p_input[18902]), .Z(n1221) );
  AND U2443 ( .A(n1222), .B(p_input[8901]), .Z(o[8901]) );
  AND U2444 ( .A(p_input[28901]), .B(p_input[18901]), .Z(n1222) );
  AND U2445 ( .A(n1223), .B(p_input[8900]), .Z(o[8900]) );
  AND U2446 ( .A(p_input[28900]), .B(p_input[18900]), .Z(n1223) );
  AND U2447 ( .A(n1224), .B(p_input[88]), .Z(o[88]) );
  AND U2448 ( .A(p_input[20088]), .B(p_input[10088]), .Z(n1224) );
  AND U2449 ( .A(n1225), .B(p_input[889]), .Z(o[889]) );
  AND U2450 ( .A(p_input[20889]), .B(p_input[10889]), .Z(n1225) );
  AND U2451 ( .A(n1226), .B(p_input[8899]), .Z(o[8899]) );
  AND U2452 ( .A(p_input[28899]), .B(p_input[18899]), .Z(n1226) );
  AND U2453 ( .A(n1227), .B(p_input[8898]), .Z(o[8898]) );
  AND U2454 ( .A(p_input[28898]), .B(p_input[18898]), .Z(n1227) );
  AND U2455 ( .A(n1228), .B(p_input[8897]), .Z(o[8897]) );
  AND U2456 ( .A(p_input[28897]), .B(p_input[18897]), .Z(n1228) );
  AND U2457 ( .A(n1229), .B(p_input[8896]), .Z(o[8896]) );
  AND U2458 ( .A(p_input[28896]), .B(p_input[18896]), .Z(n1229) );
  AND U2459 ( .A(n1230), .B(p_input[8895]), .Z(o[8895]) );
  AND U2460 ( .A(p_input[28895]), .B(p_input[18895]), .Z(n1230) );
  AND U2461 ( .A(n1231), .B(p_input[8894]), .Z(o[8894]) );
  AND U2462 ( .A(p_input[28894]), .B(p_input[18894]), .Z(n1231) );
  AND U2463 ( .A(n1232), .B(p_input[8893]), .Z(o[8893]) );
  AND U2464 ( .A(p_input[28893]), .B(p_input[18893]), .Z(n1232) );
  AND U2465 ( .A(n1233), .B(p_input[8892]), .Z(o[8892]) );
  AND U2466 ( .A(p_input[28892]), .B(p_input[18892]), .Z(n1233) );
  AND U2467 ( .A(n1234), .B(p_input[8891]), .Z(o[8891]) );
  AND U2468 ( .A(p_input[28891]), .B(p_input[18891]), .Z(n1234) );
  AND U2469 ( .A(n1235), .B(p_input[8890]), .Z(o[8890]) );
  AND U2470 ( .A(p_input[28890]), .B(p_input[18890]), .Z(n1235) );
  AND U2471 ( .A(n1236), .B(p_input[888]), .Z(o[888]) );
  AND U2472 ( .A(p_input[20888]), .B(p_input[10888]), .Z(n1236) );
  AND U2473 ( .A(n1237), .B(p_input[8889]), .Z(o[8889]) );
  AND U2474 ( .A(p_input[28889]), .B(p_input[18889]), .Z(n1237) );
  AND U2475 ( .A(n1238), .B(p_input[8888]), .Z(o[8888]) );
  AND U2476 ( .A(p_input[28888]), .B(p_input[18888]), .Z(n1238) );
  AND U2477 ( .A(n1239), .B(p_input[8887]), .Z(o[8887]) );
  AND U2478 ( .A(p_input[28887]), .B(p_input[18887]), .Z(n1239) );
  AND U2479 ( .A(n1240), .B(p_input[8886]), .Z(o[8886]) );
  AND U2480 ( .A(p_input[28886]), .B(p_input[18886]), .Z(n1240) );
  AND U2481 ( .A(n1241), .B(p_input[8885]), .Z(o[8885]) );
  AND U2482 ( .A(p_input[28885]), .B(p_input[18885]), .Z(n1241) );
  AND U2483 ( .A(n1242), .B(p_input[8884]), .Z(o[8884]) );
  AND U2484 ( .A(p_input[28884]), .B(p_input[18884]), .Z(n1242) );
  AND U2485 ( .A(n1243), .B(p_input[8883]), .Z(o[8883]) );
  AND U2486 ( .A(p_input[28883]), .B(p_input[18883]), .Z(n1243) );
  AND U2487 ( .A(n1244), .B(p_input[8882]), .Z(o[8882]) );
  AND U2488 ( .A(p_input[28882]), .B(p_input[18882]), .Z(n1244) );
  AND U2489 ( .A(n1245), .B(p_input[8881]), .Z(o[8881]) );
  AND U2490 ( .A(p_input[28881]), .B(p_input[18881]), .Z(n1245) );
  AND U2491 ( .A(n1246), .B(p_input[8880]), .Z(o[8880]) );
  AND U2492 ( .A(p_input[28880]), .B(p_input[18880]), .Z(n1246) );
  AND U2493 ( .A(n1247), .B(p_input[887]), .Z(o[887]) );
  AND U2494 ( .A(p_input[20887]), .B(p_input[10887]), .Z(n1247) );
  AND U2495 ( .A(n1248), .B(p_input[8879]), .Z(o[8879]) );
  AND U2496 ( .A(p_input[28879]), .B(p_input[18879]), .Z(n1248) );
  AND U2497 ( .A(n1249), .B(p_input[8878]), .Z(o[8878]) );
  AND U2498 ( .A(p_input[28878]), .B(p_input[18878]), .Z(n1249) );
  AND U2499 ( .A(n1250), .B(p_input[8877]), .Z(o[8877]) );
  AND U2500 ( .A(p_input[28877]), .B(p_input[18877]), .Z(n1250) );
  AND U2501 ( .A(n1251), .B(p_input[8876]), .Z(o[8876]) );
  AND U2502 ( .A(p_input[28876]), .B(p_input[18876]), .Z(n1251) );
  AND U2503 ( .A(n1252), .B(p_input[8875]), .Z(o[8875]) );
  AND U2504 ( .A(p_input[28875]), .B(p_input[18875]), .Z(n1252) );
  AND U2505 ( .A(n1253), .B(p_input[8874]), .Z(o[8874]) );
  AND U2506 ( .A(p_input[28874]), .B(p_input[18874]), .Z(n1253) );
  AND U2507 ( .A(n1254), .B(p_input[8873]), .Z(o[8873]) );
  AND U2508 ( .A(p_input[28873]), .B(p_input[18873]), .Z(n1254) );
  AND U2509 ( .A(n1255), .B(p_input[8872]), .Z(o[8872]) );
  AND U2510 ( .A(p_input[28872]), .B(p_input[18872]), .Z(n1255) );
  AND U2511 ( .A(n1256), .B(p_input[8871]), .Z(o[8871]) );
  AND U2512 ( .A(p_input[28871]), .B(p_input[18871]), .Z(n1256) );
  AND U2513 ( .A(n1257), .B(p_input[8870]), .Z(o[8870]) );
  AND U2514 ( .A(p_input[28870]), .B(p_input[18870]), .Z(n1257) );
  AND U2515 ( .A(n1258), .B(p_input[886]), .Z(o[886]) );
  AND U2516 ( .A(p_input[20886]), .B(p_input[10886]), .Z(n1258) );
  AND U2517 ( .A(n1259), .B(p_input[8869]), .Z(o[8869]) );
  AND U2518 ( .A(p_input[28869]), .B(p_input[18869]), .Z(n1259) );
  AND U2519 ( .A(n1260), .B(p_input[8868]), .Z(o[8868]) );
  AND U2520 ( .A(p_input[28868]), .B(p_input[18868]), .Z(n1260) );
  AND U2521 ( .A(n1261), .B(p_input[8867]), .Z(o[8867]) );
  AND U2522 ( .A(p_input[28867]), .B(p_input[18867]), .Z(n1261) );
  AND U2523 ( .A(n1262), .B(p_input[8866]), .Z(o[8866]) );
  AND U2524 ( .A(p_input[28866]), .B(p_input[18866]), .Z(n1262) );
  AND U2525 ( .A(n1263), .B(p_input[8865]), .Z(o[8865]) );
  AND U2526 ( .A(p_input[28865]), .B(p_input[18865]), .Z(n1263) );
  AND U2527 ( .A(n1264), .B(p_input[8864]), .Z(o[8864]) );
  AND U2528 ( .A(p_input[28864]), .B(p_input[18864]), .Z(n1264) );
  AND U2529 ( .A(n1265), .B(p_input[8863]), .Z(o[8863]) );
  AND U2530 ( .A(p_input[28863]), .B(p_input[18863]), .Z(n1265) );
  AND U2531 ( .A(n1266), .B(p_input[8862]), .Z(o[8862]) );
  AND U2532 ( .A(p_input[28862]), .B(p_input[18862]), .Z(n1266) );
  AND U2533 ( .A(n1267), .B(p_input[8861]), .Z(o[8861]) );
  AND U2534 ( .A(p_input[28861]), .B(p_input[18861]), .Z(n1267) );
  AND U2535 ( .A(n1268), .B(p_input[8860]), .Z(o[8860]) );
  AND U2536 ( .A(p_input[28860]), .B(p_input[18860]), .Z(n1268) );
  AND U2537 ( .A(n1269), .B(p_input[885]), .Z(o[885]) );
  AND U2538 ( .A(p_input[20885]), .B(p_input[10885]), .Z(n1269) );
  AND U2539 ( .A(n1270), .B(p_input[8859]), .Z(o[8859]) );
  AND U2540 ( .A(p_input[28859]), .B(p_input[18859]), .Z(n1270) );
  AND U2541 ( .A(n1271), .B(p_input[8858]), .Z(o[8858]) );
  AND U2542 ( .A(p_input[28858]), .B(p_input[18858]), .Z(n1271) );
  AND U2543 ( .A(n1272), .B(p_input[8857]), .Z(o[8857]) );
  AND U2544 ( .A(p_input[28857]), .B(p_input[18857]), .Z(n1272) );
  AND U2545 ( .A(n1273), .B(p_input[8856]), .Z(o[8856]) );
  AND U2546 ( .A(p_input[28856]), .B(p_input[18856]), .Z(n1273) );
  AND U2547 ( .A(n1274), .B(p_input[8855]), .Z(o[8855]) );
  AND U2548 ( .A(p_input[28855]), .B(p_input[18855]), .Z(n1274) );
  AND U2549 ( .A(n1275), .B(p_input[8854]), .Z(o[8854]) );
  AND U2550 ( .A(p_input[28854]), .B(p_input[18854]), .Z(n1275) );
  AND U2551 ( .A(n1276), .B(p_input[8853]), .Z(o[8853]) );
  AND U2552 ( .A(p_input[28853]), .B(p_input[18853]), .Z(n1276) );
  AND U2553 ( .A(n1277), .B(p_input[8852]), .Z(o[8852]) );
  AND U2554 ( .A(p_input[28852]), .B(p_input[18852]), .Z(n1277) );
  AND U2555 ( .A(n1278), .B(p_input[8851]), .Z(o[8851]) );
  AND U2556 ( .A(p_input[28851]), .B(p_input[18851]), .Z(n1278) );
  AND U2557 ( .A(n1279), .B(p_input[8850]), .Z(o[8850]) );
  AND U2558 ( .A(p_input[28850]), .B(p_input[18850]), .Z(n1279) );
  AND U2559 ( .A(n1280), .B(p_input[884]), .Z(o[884]) );
  AND U2560 ( .A(p_input[20884]), .B(p_input[10884]), .Z(n1280) );
  AND U2561 ( .A(n1281), .B(p_input[8849]), .Z(o[8849]) );
  AND U2562 ( .A(p_input[28849]), .B(p_input[18849]), .Z(n1281) );
  AND U2563 ( .A(n1282), .B(p_input[8848]), .Z(o[8848]) );
  AND U2564 ( .A(p_input[28848]), .B(p_input[18848]), .Z(n1282) );
  AND U2565 ( .A(n1283), .B(p_input[8847]), .Z(o[8847]) );
  AND U2566 ( .A(p_input[28847]), .B(p_input[18847]), .Z(n1283) );
  AND U2567 ( .A(n1284), .B(p_input[8846]), .Z(o[8846]) );
  AND U2568 ( .A(p_input[28846]), .B(p_input[18846]), .Z(n1284) );
  AND U2569 ( .A(n1285), .B(p_input[8845]), .Z(o[8845]) );
  AND U2570 ( .A(p_input[28845]), .B(p_input[18845]), .Z(n1285) );
  AND U2571 ( .A(n1286), .B(p_input[8844]), .Z(o[8844]) );
  AND U2572 ( .A(p_input[28844]), .B(p_input[18844]), .Z(n1286) );
  AND U2573 ( .A(n1287), .B(p_input[8843]), .Z(o[8843]) );
  AND U2574 ( .A(p_input[28843]), .B(p_input[18843]), .Z(n1287) );
  AND U2575 ( .A(n1288), .B(p_input[8842]), .Z(o[8842]) );
  AND U2576 ( .A(p_input[28842]), .B(p_input[18842]), .Z(n1288) );
  AND U2577 ( .A(n1289), .B(p_input[8841]), .Z(o[8841]) );
  AND U2578 ( .A(p_input[28841]), .B(p_input[18841]), .Z(n1289) );
  AND U2579 ( .A(n1290), .B(p_input[8840]), .Z(o[8840]) );
  AND U2580 ( .A(p_input[28840]), .B(p_input[18840]), .Z(n1290) );
  AND U2581 ( .A(n1291), .B(p_input[883]), .Z(o[883]) );
  AND U2582 ( .A(p_input[20883]), .B(p_input[10883]), .Z(n1291) );
  AND U2583 ( .A(n1292), .B(p_input[8839]), .Z(o[8839]) );
  AND U2584 ( .A(p_input[28839]), .B(p_input[18839]), .Z(n1292) );
  AND U2585 ( .A(n1293), .B(p_input[8838]), .Z(o[8838]) );
  AND U2586 ( .A(p_input[28838]), .B(p_input[18838]), .Z(n1293) );
  AND U2587 ( .A(n1294), .B(p_input[8837]), .Z(o[8837]) );
  AND U2588 ( .A(p_input[28837]), .B(p_input[18837]), .Z(n1294) );
  AND U2589 ( .A(n1295), .B(p_input[8836]), .Z(o[8836]) );
  AND U2590 ( .A(p_input[28836]), .B(p_input[18836]), .Z(n1295) );
  AND U2591 ( .A(n1296), .B(p_input[8835]), .Z(o[8835]) );
  AND U2592 ( .A(p_input[28835]), .B(p_input[18835]), .Z(n1296) );
  AND U2593 ( .A(n1297), .B(p_input[8834]), .Z(o[8834]) );
  AND U2594 ( .A(p_input[28834]), .B(p_input[18834]), .Z(n1297) );
  AND U2595 ( .A(n1298), .B(p_input[8833]), .Z(o[8833]) );
  AND U2596 ( .A(p_input[28833]), .B(p_input[18833]), .Z(n1298) );
  AND U2597 ( .A(n1299), .B(p_input[8832]), .Z(o[8832]) );
  AND U2598 ( .A(p_input[28832]), .B(p_input[18832]), .Z(n1299) );
  AND U2599 ( .A(n1300), .B(p_input[8831]), .Z(o[8831]) );
  AND U2600 ( .A(p_input[28831]), .B(p_input[18831]), .Z(n1300) );
  AND U2601 ( .A(n1301), .B(p_input[8830]), .Z(o[8830]) );
  AND U2602 ( .A(p_input[28830]), .B(p_input[18830]), .Z(n1301) );
  AND U2603 ( .A(n1302), .B(p_input[882]), .Z(o[882]) );
  AND U2604 ( .A(p_input[20882]), .B(p_input[10882]), .Z(n1302) );
  AND U2605 ( .A(n1303), .B(p_input[8829]), .Z(o[8829]) );
  AND U2606 ( .A(p_input[28829]), .B(p_input[18829]), .Z(n1303) );
  AND U2607 ( .A(n1304), .B(p_input[8828]), .Z(o[8828]) );
  AND U2608 ( .A(p_input[28828]), .B(p_input[18828]), .Z(n1304) );
  AND U2609 ( .A(n1305), .B(p_input[8827]), .Z(o[8827]) );
  AND U2610 ( .A(p_input[28827]), .B(p_input[18827]), .Z(n1305) );
  AND U2611 ( .A(n1306), .B(p_input[8826]), .Z(o[8826]) );
  AND U2612 ( .A(p_input[28826]), .B(p_input[18826]), .Z(n1306) );
  AND U2613 ( .A(n1307), .B(p_input[8825]), .Z(o[8825]) );
  AND U2614 ( .A(p_input[28825]), .B(p_input[18825]), .Z(n1307) );
  AND U2615 ( .A(n1308), .B(p_input[8824]), .Z(o[8824]) );
  AND U2616 ( .A(p_input[28824]), .B(p_input[18824]), .Z(n1308) );
  AND U2617 ( .A(n1309), .B(p_input[8823]), .Z(o[8823]) );
  AND U2618 ( .A(p_input[28823]), .B(p_input[18823]), .Z(n1309) );
  AND U2619 ( .A(n1310), .B(p_input[8822]), .Z(o[8822]) );
  AND U2620 ( .A(p_input[28822]), .B(p_input[18822]), .Z(n1310) );
  AND U2621 ( .A(n1311), .B(p_input[8821]), .Z(o[8821]) );
  AND U2622 ( .A(p_input[28821]), .B(p_input[18821]), .Z(n1311) );
  AND U2623 ( .A(n1312), .B(p_input[8820]), .Z(o[8820]) );
  AND U2624 ( .A(p_input[28820]), .B(p_input[18820]), .Z(n1312) );
  AND U2625 ( .A(n1313), .B(p_input[881]), .Z(o[881]) );
  AND U2626 ( .A(p_input[20881]), .B(p_input[10881]), .Z(n1313) );
  AND U2627 ( .A(n1314), .B(p_input[8819]), .Z(o[8819]) );
  AND U2628 ( .A(p_input[28819]), .B(p_input[18819]), .Z(n1314) );
  AND U2629 ( .A(n1315), .B(p_input[8818]), .Z(o[8818]) );
  AND U2630 ( .A(p_input[28818]), .B(p_input[18818]), .Z(n1315) );
  AND U2631 ( .A(n1316), .B(p_input[8817]), .Z(o[8817]) );
  AND U2632 ( .A(p_input[28817]), .B(p_input[18817]), .Z(n1316) );
  AND U2633 ( .A(n1317), .B(p_input[8816]), .Z(o[8816]) );
  AND U2634 ( .A(p_input[28816]), .B(p_input[18816]), .Z(n1317) );
  AND U2635 ( .A(n1318), .B(p_input[8815]), .Z(o[8815]) );
  AND U2636 ( .A(p_input[28815]), .B(p_input[18815]), .Z(n1318) );
  AND U2637 ( .A(n1319), .B(p_input[8814]), .Z(o[8814]) );
  AND U2638 ( .A(p_input[28814]), .B(p_input[18814]), .Z(n1319) );
  AND U2639 ( .A(n1320), .B(p_input[8813]), .Z(o[8813]) );
  AND U2640 ( .A(p_input[28813]), .B(p_input[18813]), .Z(n1320) );
  AND U2641 ( .A(n1321), .B(p_input[8812]), .Z(o[8812]) );
  AND U2642 ( .A(p_input[28812]), .B(p_input[18812]), .Z(n1321) );
  AND U2643 ( .A(n1322), .B(p_input[8811]), .Z(o[8811]) );
  AND U2644 ( .A(p_input[28811]), .B(p_input[18811]), .Z(n1322) );
  AND U2645 ( .A(n1323), .B(p_input[8810]), .Z(o[8810]) );
  AND U2646 ( .A(p_input[28810]), .B(p_input[18810]), .Z(n1323) );
  AND U2647 ( .A(n1324), .B(p_input[880]), .Z(o[880]) );
  AND U2648 ( .A(p_input[20880]), .B(p_input[10880]), .Z(n1324) );
  AND U2649 ( .A(n1325), .B(p_input[8809]), .Z(o[8809]) );
  AND U2650 ( .A(p_input[28809]), .B(p_input[18809]), .Z(n1325) );
  AND U2651 ( .A(n1326), .B(p_input[8808]), .Z(o[8808]) );
  AND U2652 ( .A(p_input[28808]), .B(p_input[18808]), .Z(n1326) );
  AND U2653 ( .A(n1327), .B(p_input[8807]), .Z(o[8807]) );
  AND U2654 ( .A(p_input[28807]), .B(p_input[18807]), .Z(n1327) );
  AND U2655 ( .A(n1328), .B(p_input[8806]), .Z(o[8806]) );
  AND U2656 ( .A(p_input[28806]), .B(p_input[18806]), .Z(n1328) );
  AND U2657 ( .A(n1329), .B(p_input[8805]), .Z(o[8805]) );
  AND U2658 ( .A(p_input[28805]), .B(p_input[18805]), .Z(n1329) );
  AND U2659 ( .A(n1330), .B(p_input[8804]), .Z(o[8804]) );
  AND U2660 ( .A(p_input[28804]), .B(p_input[18804]), .Z(n1330) );
  AND U2661 ( .A(n1331), .B(p_input[8803]), .Z(o[8803]) );
  AND U2662 ( .A(p_input[28803]), .B(p_input[18803]), .Z(n1331) );
  AND U2663 ( .A(n1332), .B(p_input[8802]), .Z(o[8802]) );
  AND U2664 ( .A(p_input[28802]), .B(p_input[18802]), .Z(n1332) );
  AND U2665 ( .A(n1333), .B(p_input[8801]), .Z(o[8801]) );
  AND U2666 ( .A(p_input[28801]), .B(p_input[18801]), .Z(n1333) );
  AND U2667 ( .A(n1334), .B(p_input[8800]), .Z(o[8800]) );
  AND U2668 ( .A(p_input[28800]), .B(p_input[18800]), .Z(n1334) );
  AND U2669 ( .A(n1335), .B(p_input[87]), .Z(o[87]) );
  AND U2670 ( .A(p_input[20087]), .B(p_input[10087]), .Z(n1335) );
  AND U2671 ( .A(n1336), .B(p_input[879]), .Z(o[879]) );
  AND U2672 ( .A(p_input[20879]), .B(p_input[10879]), .Z(n1336) );
  AND U2673 ( .A(n1337), .B(p_input[8799]), .Z(o[8799]) );
  AND U2674 ( .A(p_input[28799]), .B(p_input[18799]), .Z(n1337) );
  AND U2675 ( .A(n1338), .B(p_input[8798]), .Z(o[8798]) );
  AND U2676 ( .A(p_input[28798]), .B(p_input[18798]), .Z(n1338) );
  AND U2677 ( .A(n1339), .B(p_input[8797]), .Z(o[8797]) );
  AND U2678 ( .A(p_input[28797]), .B(p_input[18797]), .Z(n1339) );
  AND U2679 ( .A(n1340), .B(p_input[8796]), .Z(o[8796]) );
  AND U2680 ( .A(p_input[28796]), .B(p_input[18796]), .Z(n1340) );
  AND U2681 ( .A(n1341), .B(p_input[8795]), .Z(o[8795]) );
  AND U2682 ( .A(p_input[28795]), .B(p_input[18795]), .Z(n1341) );
  AND U2683 ( .A(n1342), .B(p_input[8794]), .Z(o[8794]) );
  AND U2684 ( .A(p_input[28794]), .B(p_input[18794]), .Z(n1342) );
  AND U2685 ( .A(n1343), .B(p_input[8793]), .Z(o[8793]) );
  AND U2686 ( .A(p_input[28793]), .B(p_input[18793]), .Z(n1343) );
  AND U2687 ( .A(n1344), .B(p_input[8792]), .Z(o[8792]) );
  AND U2688 ( .A(p_input[28792]), .B(p_input[18792]), .Z(n1344) );
  AND U2689 ( .A(n1345), .B(p_input[8791]), .Z(o[8791]) );
  AND U2690 ( .A(p_input[28791]), .B(p_input[18791]), .Z(n1345) );
  AND U2691 ( .A(n1346), .B(p_input[8790]), .Z(o[8790]) );
  AND U2692 ( .A(p_input[28790]), .B(p_input[18790]), .Z(n1346) );
  AND U2693 ( .A(n1347), .B(p_input[878]), .Z(o[878]) );
  AND U2694 ( .A(p_input[20878]), .B(p_input[10878]), .Z(n1347) );
  AND U2695 ( .A(n1348), .B(p_input[8789]), .Z(o[8789]) );
  AND U2696 ( .A(p_input[28789]), .B(p_input[18789]), .Z(n1348) );
  AND U2697 ( .A(n1349), .B(p_input[8788]), .Z(o[8788]) );
  AND U2698 ( .A(p_input[28788]), .B(p_input[18788]), .Z(n1349) );
  AND U2699 ( .A(n1350), .B(p_input[8787]), .Z(o[8787]) );
  AND U2700 ( .A(p_input[28787]), .B(p_input[18787]), .Z(n1350) );
  AND U2701 ( .A(n1351), .B(p_input[8786]), .Z(o[8786]) );
  AND U2702 ( .A(p_input[28786]), .B(p_input[18786]), .Z(n1351) );
  AND U2703 ( .A(n1352), .B(p_input[8785]), .Z(o[8785]) );
  AND U2704 ( .A(p_input[28785]), .B(p_input[18785]), .Z(n1352) );
  AND U2705 ( .A(n1353), .B(p_input[8784]), .Z(o[8784]) );
  AND U2706 ( .A(p_input[28784]), .B(p_input[18784]), .Z(n1353) );
  AND U2707 ( .A(n1354), .B(p_input[8783]), .Z(o[8783]) );
  AND U2708 ( .A(p_input[28783]), .B(p_input[18783]), .Z(n1354) );
  AND U2709 ( .A(n1355), .B(p_input[8782]), .Z(o[8782]) );
  AND U2710 ( .A(p_input[28782]), .B(p_input[18782]), .Z(n1355) );
  AND U2711 ( .A(n1356), .B(p_input[8781]), .Z(o[8781]) );
  AND U2712 ( .A(p_input[28781]), .B(p_input[18781]), .Z(n1356) );
  AND U2713 ( .A(n1357), .B(p_input[8780]), .Z(o[8780]) );
  AND U2714 ( .A(p_input[28780]), .B(p_input[18780]), .Z(n1357) );
  AND U2715 ( .A(n1358), .B(p_input[877]), .Z(o[877]) );
  AND U2716 ( .A(p_input[20877]), .B(p_input[10877]), .Z(n1358) );
  AND U2717 ( .A(n1359), .B(p_input[8779]), .Z(o[8779]) );
  AND U2718 ( .A(p_input[28779]), .B(p_input[18779]), .Z(n1359) );
  AND U2719 ( .A(n1360), .B(p_input[8778]), .Z(o[8778]) );
  AND U2720 ( .A(p_input[28778]), .B(p_input[18778]), .Z(n1360) );
  AND U2721 ( .A(n1361), .B(p_input[8777]), .Z(o[8777]) );
  AND U2722 ( .A(p_input[28777]), .B(p_input[18777]), .Z(n1361) );
  AND U2723 ( .A(n1362), .B(p_input[8776]), .Z(o[8776]) );
  AND U2724 ( .A(p_input[28776]), .B(p_input[18776]), .Z(n1362) );
  AND U2725 ( .A(n1363), .B(p_input[8775]), .Z(o[8775]) );
  AND U2726 ( .A(p_input[28775]), .B(p_input[18775]), .Z(n1363) );
  AND U2727 ( .A(n1364), .B(p_input[8774]), .Z(o[8774]) );
  AND U2728 ( .A(p_input[28774]), .B(p_input[18774]), .Z(n1364) );
  AND U2729 ( .A(n1365), .B(p_input[8773]), .Z(o[8773]) );
  AND U2730 ( .A(p_input[28773]), .B(p_input[18773]), .Z(n1365) );
  AND U2731 ( .A(n1366), .B(p_input[8772]), .Z(o[8772]) );
  AND U2732 ( .A(p_input[28772]), .B(p_input[18772]), .Z(n1366) );
  AND U2733 ( .A(n1367), .B(p_input[8771]), .Z(o[8771]) );
  AND U2734 ( .A(p_input[28771]), .B(p_input[18771]), .Z(n1367) );
  AND U2735 ( .A(n1368), .B(p_input[8770]), .Z(o[8770]) );
  AND U2736 ( .A(p_input[28770]), .B(p_input[18770]), .Z(n1368) );
  AND U2737 ( .A(n1369), .B(p_input[876]), .Z(o[876]) );
  AND U2738 ( .A(p_input[20876]), .B(p_input[10876]), .Z(n1369) );
  AND U2739 ( .A(n1370), .B(p_input[8769]), .Z(o[8769]) );
  AND U2740 ( .A(p_input[28769]), .B(p_input[18769]), .Z(n1370) );
  AND U2741 ( .A(n1371), .B(p_input[8768]), .Z(o[8768]) );
  AND U2742 ( .A(p_input[28768]), .B(p_input[18768]), .Z(n1371) );
  AND U2743 ( .A(n1372), .B(p_input[8767]), .Z(o[8767]) );
  AND U2744 ( .A(p_input[28767]), .B(p_input[18767]), .Z(n1372) );
  AND U2745 ( .A(n1373), .B(p_input[8766]), .Z(o[8766]) );
  AND U2746 ( .A(p_input[28766]), .B(p_input[18766]), .Z(n1373) );
  AND U2747 ( .A(n1374), .B(p_input[8765]), .Z(o[8765]) );
  AND U2748 ( .A(p_input[28765]), .B(p_input[18765]), .Z(n1374) );
  AND U2749 ( .A(n1375), .B(p_input[8764]), .Z(o[8764]) );
  AND U2750 ( .A(p_input[28764]), .B(p_input[18764]), .Z(n1375) );
  AND U2751 ( .A(n1376), .B(p_input[8763]), .Z(o[8763]) );
  AND U2752 ( .A(p_input[28763]), .B(p_input[18763]), .Z(n1376) );
  AND U2753 ( .A(n1377), .B(p_input[8762]), .Z(o[8762]) );
  AND U2754 ( .A(p_input[28762]), .B(p_input[18762]), .Z(n1377) );
  AND U2755 ( .A(n1378), .B(p_input[8761]), .Z(o[8761]) );
  AND U2756 ( .A(p_input[28761]), .B(p_input[18761]), .Z(n1378) );
  AND U2757 ( .A(n1379), .B(p_input[8760]), .Z(o[8760]) );
  AND U2758 ( .A(p_input[28760]), .B(p_input[18760]), .Z(n1379) );
  AND U2759 ( .A(n1380), .B(p_input[875]), .Z(o[875]) );
  AND U2760 ( .A(p_input[20875]), .B(p_input[10875]), .Z(n1380) );
  AND U2761 ( .A(n1381), .B(p_input[8759]), .Z(o[8759]) );
  AND U2762 ( .A(p_input[28759]), .B(p_input[18759]), .Z(n1381) );
  AND U2763 ( .A(n1382), .B(p_input[8758]), .Z(o[8758]) );
  AND U2764 ( .A(p_input[28758]), .B(p_input[18758]), .Z(n1382) );
  AND U2765 ( .A(n1383), .B(p_input[8757]), .Z(o[8757]) );
  AND U2766 ( .A(p_input[28757]), .B(p_input[18757]), .Z(n1383) );
  AND U2767 ( .A(n1384), .B(p_input[8756]), .Z(o[8756]) );
  AND U2768 ( .A(p_input[28756]), .B(p_input[18756]), .Z(n1384) );
  AND U2769 ( .A(n1385), .B(p_input[8755]), .Z(o[8755]) );
  AND U2770 ( .A(p_input[28755]), .B(p_input[18755]), .Z(n1385) );
  AND U2771 ( .A(n1386), .B(p_input[8754]), .Z(o[8754]) );
  AND U2772 ( .A(p_input[28754]), .B(p_input[18754]), .Z(n1386) );
  AND U2773 ( .A(n1387), .B(p_input[8753]), .Z(o[8753]) );
  AND U2774 ( .A(p_input[28753]), .B(p_input[18753]), .Z(n1387) );
  AND U2775 ( .A(n1388), .B(p_input[8752]), .Z(o[8752]) );
  AND U2776 ( .A(p_input[28752]), .B(p_input[18752]), .Z(n1388) );
  AND U2777 ( .A(n1389), .B(p_input[8751]), .Z(o[8751]) );
  AND U2778 ( .A(p_input[28751]), .B(p_input[18751]), .Z(n1389) );
  AND U2779 ( .A(n1390), .B(p_input[8750]), .Z(o[8750]) );
  AND U2780 ( .A(p_input[28750]), .B(p_input[18750]), .Z(n1390) );
  AND U2781 ( .A(n1391), .B(p_input[874]), .Z(o[874]) );
  AND U2782 ( .A(p_input[20874]), .B(p_input[10874]), .Z(n1391) );
  AND U2783 ( .A(n1392), .B(p_input[8749]), .Z(o[8749]) );
  AND U2784 ( .A(p_input[28749]), .B(p_input[18749]), .Z(n1392) );
  AND U2785 ( .A(n1393), .B(p_input[8748]), .Z(o[8748]) );
  AND U2786 ( .A(p_input[28748]), .B(p_input[18748]), .Z(n1393) );
  AND U2787 ( .A(n1394), .B(p_input[8747]), .Z(o[8747]) );
  AND U2788 ( .A(p_input[28747]), .B(p_input[18747]), .Z(n1394) );
  AND U2789 ( .A(n1395), .B(p_input[8746]), .Z(o[8746]) );
  AND U2790 ( .A(p_input[28746]), .B(p_input[18746]), .Z(n1395) );
  AND U2791 ( .A(n1396), .B(p_input[8745]), .Z(o[8745]) );
  AND U2792 ( .A(p_input[28745]), .B(p_input[18745]), .Z(n1396) );
  AND U2793 ( .A(n1397), .B(p_input[8744]), .Z(o[8744]) );
  AND U2794 ( .A(p_input[28744]), .B(p_input[18744]), .Z(n1397) );
  AND U2795 ( .A(n1398), .B(p_input[8743]), .Z(o[8743]) );
  AND U2796 ( .A(p_input[28743]), .B(p_input[18743]), .Z(n1398) );
  AND U2797 ( .A(n1399), .B(p_input[8742]), .Z(o[8742]) );
  AND U2798 ( .A(p_input[28742]), .B(p_input[18742]), .Z(n1399) );
  AND U2799 ( .A(n1400), .B(p_input[8741]), .Z(o[8741]) );
  AND U2800 ( .A(p_input[28741]), .B(p_input[18741]), .Z(n1400) );
  AND U2801 ( .A(n1401), .B(p_input[8740]), .Z(o[8740]) );
  AND U2802 ( .A(p_input[28740]), .B(p_input[18740]), .Z(n1401) );
  AND U2803 ( .A(n1402), .B(p_input[873]), .Z(o[873]) );
  AND U2804 ( .A(p_input[20873]), .B(p_input[10873]), .Z(n1402) );
  AND U2805 ( .A(n1403), .B(p_input[8739]), .Z(o[8739]) );
  AND U2806 ( .A(p_input[28739]), .B(p_input[18739]), .Z(n1403) );
  AND U2807 ( .A(n1404), .B(p_input[8738]), .Z(o[8738]) );
  AND U2808 ( .A(p_input[28738]), .B(p_input[18738]), .Z(n1404) );
  AND U2809 ( .A(n1405), .B(p_input[8737]), .Z(o[8737]) );
  AND U2810 ( .A(p_input[28737]), .B(p_input[18737]), .Z(n1405) );
  AND U2811 ( .A(n1406), .B(p_input[8736]), .Z(o[8736]) );
  AND U2812 ( .A(p_input[28736]), .B(p_input[18736]), .Z(n1406) );
  AND U2813 ( .A(n1407), .B(p_input[8735]), .Z(o[8735]) );
  AND U2814 ( .A(p_input[28735]), .B(p_input[18735]), .Z(n1407) );
  AND U2815 ( .A(n1408), .B(p_input[8734]), .Z(o[8734]) );
  AND U2816 ( .A(p_input[28734]), .B(p_input[18734]), .Z(n1408) );
  AND U2817 ( .A(n1409), .B(p_input[8733]), .Z(o[8733]) );
  AND U2818 ( .A(p_input[28733]), .B(p_input[18733]), .Z(n1409) );
  AND U2819 ( .A(n1410), .B(p_input[8732]), .Z(o[8732]) );
  AND U2820 ( .A(p_input[28732]), .B(p_input[18732]), .Z(n1410) );
  AND U2821 ( .A(n1411), .B(p_input[8731]), .Z(o[8731]) );
  AND U2822 ( .A(p_input[28731]), .B(p_input[18731]), .Z(n1411) );
  AND U2823 ( .A(n1412), .B(p_input[8730]), .Z(o[8730]) );
  AND U2824 ( .A(p_input[28730]), .B(p_input[18730]), .Z(n1412) );
  AND U2825 ( .A(n1413), .B(p_input[872]), .Z(o[872]) );
  AND U2826 ( .A(p_input[20872]), .B(p_input[10872]), .Z(n1413) );
  AND U2827 ( .A(n1414), .B(p_input[8729]), .Z(o[8729]) );
  AND U2828 ( .A(p_input[28729]), .B(p_input[18729]), .Z(n1414) );
  AND U2829 ( .A(n1415), .B(p_input[8728]), .Z(o[8728]) );
  AND U2830 ( .A(p_input[28728]), .B(p_input[18728]), .Z(n1415) );
  AND U2831 ( .A(n1416), .B(p_input[8727]), .Z(o[8727]) );
  AND U2832 ( .A(p_input[28727]), .B(p_input[18727]), .Z(n1416) );
  AND U2833 ( .A(n1417), .B(p_input[8726]), .Z(o[8726]) );
  AND U2834 ( .A(p_input[28726]), .B(p_input[18726]), .Z(n1417) );
  AND U2835 ( .A(n1418), .B(p_input[8725]), .Z(o[8725]) );
  AND U2836 ( .A(p_input[28725]), .B(p_input[18725]), .Z(n1418) );
  AND U2837 ( .A(n1419), .B(p_input[8724]), .Z(o[8724]) );
  AND U2838 ( .A(p_input[28724]), .B(p_input[18724]), .Z(n1419) );
  AND U2839 ( .A(n1420), .B(p_input[8723]), .Z(o[8723]) );
  AND U2840 ( .A(p_input[28723]), .B(p_input[18723]), .Z(n1420) );
  AND U2841 ( .A(n1421), .B(p_input[8722]), .Z(o[8722]) );
  AND U2842 ( .A(p_input[28722]), .B(p_input[18722]), .Z(n1421) );
  AND U2843 ( .A(n1422), .B(p_input[8721]), .Z(o[8721]) );
  AND U2844 ( .A(p_input[28721]), .B(p_input[18721]), .Z(n1422) );
  AND U2845 ( .A(n1423), .B(p_input[8720]), .Z(o[8720]) );
  AND U2846 ( .A(p_input[28720]), .B(p_input[18720]), .Z(n1423) );
  AND U2847 ( .A(n1424), .B(p_input[871]), .Z(o[871]) );
  AND U2848 ( .A(p_input[20871]), .B(p_input[10871]), .Z(n1424) );
  AND U2849 ( .A(n1425), .B(p_input[8719]), .Z(o[8719]) );
  AND U2850 ( .A(p_input[28719]), .B(p_input[18719]), .Z(n1425) );
  AND U2851 ( .A(n1426), .B(p_input[8718]), .Z(o[8718]) );
  AND U2852 ( .A(p_input[28718]), .B(p_input[18718]), .Z(n1426) );
  AND U2853 ( .A(n1427), .B(p_input[8717]), .Z(o[8717]) );
  AND U2854 ( .A(p_input[28717]), .B(p_input[18717]), .Z(n1427) );
  AND U2855 ( .A(n1428), .B(p_input[8716]), .Z(o[8716]) );
  AND U2856 ( .A(p_input[28716]), .B(p_input[18716]), .Z(n1428) );
  AND U2857 ( .A(n1429), .B(p_input[8715]), .Z(o[8715]) );
  AND U2858 ( .A(p_input[28715]), .B(p_input[18715]), .Z(n1429) );
  AND U2859 ( .A(n1430), .B(p_input[8714]), .Z(o[8714]) );
  AND U2860 ( .A(p_input[28714]), .B(p_input[18714]), .Z(n1430) );
  AND U2861 ( .A(n1431), .B(p_input[8713]), .Z(o[8713]) );
  AND U2862 ( .A(p_input[28713]), .B(p_input[18713]), .Z(n1431) );
  AND U2863 ( .A(n1432), .B(p_input[8712]), .Z(o[8712]) );
  AND U2864 ( .A(p_input[28712]), .B(p_input[18712]), .Z(n1432) );
  AND U2865 ( .A(n1433), .B(p_input[8711]), .Z(o[8711]) );
  AND U2866 ( .A(p_input[28711]), .B(p_input[18711]), .Z(n1433) );
  AND U2867 ( .A(n1434), .B(p_input[8710]), .Z(o[8710]) );
  AND U2868 ( .A(p_input[28710]), .B(p_input[18710]), .Z(n1434) );
  AND U2869 ( .A(n1435), .B(p_input[870]), .Z(o[870]) );
  AND U2870 ( .A(p_input[20870]), .B(p_input[10870]), .Z(n1435) );
  AND U2871 ( .A(n1436), .B(p_input[8709]), .Z(o[8709]) );
  AND U2872 ( .A(p_input[28709]), .B(p_input[18709]), .Z(n1436) );
  AND U2873 ( .A(n1437), .B(p_input[8708]), .Z(o[8708]) );
  AND U2874 ( .A(p_input[28708]), .B(p_input[18708]), .Z(n1437) );
  AND U2875 ( .A(n1438), .B(p_input[8707]), .Z(o[8707]) );
  AND U2876 ( .A(p_input[28707]), .B(p_input[18707]), .Z(n1438) );
  AND U2877 ( .A(n1439), .B(p_input[8706]), .Z(o[8706]) );
  AND U2878 ( .A(p_input[28706]), .B(p_input[18706]), .Z(n1439) );
  AND U2879 ( .A(n1440), .B(p_input[8705]), .Z(o[8705]) );
  AND U2880 ( .A(p_input[28705]), .B(p_input[18705]), .Z(n1440) );
  AND U2881 ( .A(n1441), .B(p_input[8704]), .Z(o[8704]) );
  AND U2882 ( .A(p_input[28704]), .B(p_input[18704]), .Z(n1441) );
  AND U2883 ( .A(n1442), .B(p_input[8703]), .Z(o[8703]) );
  AND U2884 ( .A(p_input[28703]), .B(p_input[18703]), .Z(n1442) );
  AND U2885 ( .A(n1443), .B(p_input[8702]), .Z(o[8702]) );
  AND U2886 ( .A(p_input[28702]), .B(p_input[18702]), .Z(n1443) );
  AND U2887 ( .A(n1444), .B(p_input[8701]), .Z(o[8701]) );
  AND U2888 ( .A(p_input[28701]), .B(p_input[18701]), .Z(n1444) );
  AND U2889 ( .A(n1445), .B(p_input[8700]), .Z(o[8700]) );
  AND U2890 ( .A(p_input[28700]), .B(p_input[18700]), .Z(n1445) );
  AND U2891 ( .A(n1446), .B(p_input[86]), .Z(o[86]) );
  AND U2892 ( .A(p_input[20086]), .B(p_input[10086]), .Z(n1446) );
  AND U2893 ( .A(n1447), .B(p_input[869]), .Z(o[869]) );
  AND U2894 ( .A(p_input[20869]), .B(p_input[10869]), .Z(n1447) );
  AND U2895 ( .A(n1448), .B(p_input[8699]), .Z(o[8699]) );
  AND U2896 ( .A(p_input[28699]), .B(p_input[18699]), .Z(n1448) );
  AND U2897 ( .A(n1449), .B(p_input[8698]), .Z(o[8698]) );
  AND U2898 ( .A(p_input[28698]), .B(p_input[18698]), .Z(n1449) );
  AND U2899 ( .A(n1450), .B(p_input[8697]), .Z(o[8697]) );
  AND U2900 ( .A(p_input[28697]), .B(p_input[18697]), .Z(n1450) );
  AND U2901 ( .A(n1451), .B(p_input[8696]), .Z(o[8696]) );
  AND U2902 ( .A(p_input[28696]), .B(p_input[18696]), .Z(n1451) );
  AND U2903 ( .A(n1452), .B(p_input[8695]), .Z(o[8695]) );
  AND U2904 ( .A(p_input[28695]), .B(p_input[18695]), .Z(n1452) );
  AND U2905 ( .A(n1453), .B(p_input[8694]), .Z(o[8694]) );
  AND U2906 ( .A(p_input[28694]), .B(p_input[18694]), .Z(n1453) );
  AND U2907 ( .A(n1454), .B(p_input[8693]), .Z(o[8693]) );
  AND U2908 ( .A(p_input[28693]), .B(p_input[18693]), .Z(n1454) );
  AND U2909 ( .A(n1455), .B(p_input[8692]), .Z(o[8692]) );
  AND U2910 ( .A(p_input[28692]), .B(p_input[18692]), .Z(n1455) );
  AND U2911 ( .A(n1456), .B(p_input[8691]), .Z(o[8691]) );
  AND U2912 ( .A(p_input[28691]), .B(p_input[18691]), .Z(n1456) );
  AND U2913 ( .A(n1457), .B(p_input[8690]), .Z(o[8690]) );
  AND U2914 ( .A(p_input[28690]), .B(p_input[18690]), .Z(n1457) );
  AND U2915 ( .A(n1458), .B(p_input[868]), .Z(o[868]) );
  AND U2916 ( .A(p_input[20868]), .B(p_input[10868]), .Z(n1458) );
  AND U2917 ( .A(n1459), .B(p_input[8689]), .Z(o[8689]) );
  AND U2918 ( .A(p_input[28689]), .B(p_input[18689]), .Z(n1459) );
  AND U2919 ( .A(n1460), .B(p_input[8688]), .Z(o[8688]) );
  AND U2920 ( .A(p_input[28688]), .B(p_input[18688]), .Z(n1460) );
  AND U2921 ( .A(n1461), .B(p_input[8687]), .Z(o[8687]) );
  AND U2922 ( .A(p_input[28687]), .B(p_input[18687]), .Z(n1461) );
  AND U2923 ( .A(n1462), .B(p_input[8686]), .Z(o[8686]) );
  AND U2924 ( .A(p_input[28686]), .B(p_input[18686]), .Z(n1462) );
  AND U2925 ( .A(n1463), .B(p_input[8685]), .Z(o[8685]) );
  AND U2926 ( .A(p_input[28685]), .B(p_input[18685]), .Z(n1463) );
  AND U2927 ( .A(n1464), .B(p_input[8684]), .Z(o[8684]) );
  AND U2928 ( .A(p_input[28684]), .B(p_input[18684]), .Z(n1464) );
  AND U2929 ( .A(n1465), .B(p_input[8683]), .Z(o[8683]) );
  AND U2930 ( .A(p_input[28683]), .B(p_input[18683]), .Z(n1465) );
  AND U2931 ( .A(n1466), .B(p_input[8682]), .Z(o[8682]) );
  AND U2932 ( .A(p_input[28682]), .B(p_input[18682]), .Z(n1466) );
  AND U2933 ( .A(n1467), .B(p_input[8681]), .Z(o[8681]) );
  AND U2934 ( .A(p_input[28681]), .B(p_input[18681]), .Z(n1467) );
  AND U2935 ( .A(n1468), .B(p_input[8680]), .Z(o[8680]) );
  AND U2936 ( .A(p_input[28680]), .B(p_input[18680]), .Z(n1468) );
  AND U2937 ( .A(n1469), .B(p_input[867]), .Z(o[867]) );
  AND U2938 ( .A(p_input[20867]), .B(p_input[10867]), .Z(n1469) );
  AND U2939 ( .A(n1470), .B(p_input[8679]), .Z(o[8679]) );
  AND U2940 ( .A(p_input[28679]), .B(p_input[18679]), .Z(n1470) );
  AND U2941 ( .A(n1471), .B(p_input[8678]), .Z(o[8678]) );
  AND U2942 ( .A(p_input[28678]), .B(p_input[18678]), .Z(n1471) );
  AND U2943 ( .A(n1472), .B(p_input[8677]), .Z(o[8677]) );
  AND U2944 ( .A(p_input[28677]), .B(p_input[18677]), .Z(n1472) );
  AND U2945 ( .A(n1473), .B(p_input[8676]), .Z(o[8676]) );
  AND U2946 ( .A(p_input[28676]), .B(p_input[18676]), .Z(n1473) );
  AND U2947 ( .A(n1474), .B(p_input[8675]), .Z(o[8675]) );
  AND U2948 ( .A(p_input[28675]), .B(p_input[18675]), .Z(n1474) );
  AND U2949 ( .A(n1475), .B(p_input[8674]), .Z(o[8674]) );
  AND U2950 ( .A(p_input[28674]), .B(p_input[18674]), .Z(n1475) );
  AND U2951 ( .A(n1476), .B(p_input[8673]), .Z(o[8673]) );
  AND U2952 ( .A(p_input[28673]), .B(p_input[18673]), .Z(n1476) );
  AND U2953 ( .A(n1477), .B(p_input[8672]), .Z(o[8672]) );
  AND U2954 ( .A(p_input[28672]), .B(p_input[18672]), .Z(n1477) );
  AND U2955 ( .A(n1478), .B(p_input[8671]), .Z(o[8671]) );
  AND U2956 ( .A(p_input[28671]), .B(p_input[18671]), .Z(n1478) );
  AND U2957 ( .A(n1479), .B(p_input[8670]), .Z(o[8670]) );
  AND U2958 ( .A(p_input[28670]), .B(p_input[18670]), .Z(n1479) );
  AND U2959 ( .A(n1480), .B(p_input[866]), .Z(o[866]) );
  AND U2960 ( .A(p_input[20866]), .B(p_input[10866]), .Z(n1480) );
  AND U2961 ( .A(n1481), .B(p_input[8669]), .Z(o[8669]) );
  AND U2962 ( .A(p_input[28669]), .B(p_input[18669]), .Z(n1481) );
  AND U2963 ( .A(n1482), .B(p_input[8668]), .Z(o[8668]) );
  AND U2964 ( .A(p_input[28668]), .B(p_input[18668]), .Z(n1482) );
  AND U2965 ( .A(n1483), .B(p_input[8667]), .Z(o[8667]) );
  AND U2966 ( .A(p_input[28667]), .B(p_input[18667]), .Z(n1483) );
  AND U2967 ( .A(n1484), .B(p_input[8666]), .Z(o[8666]) );
  AND U2968 ( .A(p_input[28666]), .B(p_input[18666]), .Z(n1484) );
  AND U2969 ( .A(n1485), .B(p_input[8665]), .Z(o[8665]) );
  AND U2970 ( .A(p_input[28665]), .B(p_input[18665]), .Z(n1485) );
  AND U2971 ( .A(n1486), .B(p_input[8664]), .Z(o[8664]) );
  AND U2972 ( .A(p_input[28664]), .B(p_input[18664]), .Z(n1486) );
  AND U2973 ( .A(n1487), .B(p_input[8663]), .Z(o[8663]) );
  AND U2974 ( .A(p_input[28663]), .B(p_input[18663]), .Z(n1487) );
  AND U2975 ( .A(n1488), .B(p_input[8662]), .Z(o[8662]) );
  AND U2976 ( .A(p_input[28662]), .B(p_input[18662]), .Z(n1488) );
  AND U2977 ( .A(n1489), .B(p_input[8661]), .Z(o[8661]) );
  AND U2978 ( .A(p_input[28661]), .B(p_input[18661]), .Z(n1489) );
  AND U2979 ( .A(n1490), .B(p_input[8660]), .Z(o[8660]) );
  AND U2980 ( .A(p_input[28660]), .B(p_input[18660]), .Z(n1490) );
  AND U2981 ( .A(n1491), .B(p_input[865]), .Z(o[865]) );
  AND U2982 ( .A(p_input[20865]), .B(p_input[10865]), .Z(n1491) );
  AND U2983 ( .A(n1492), .B(p_input[8659]), .Z(o[8659]) );
  AND U2984 ( .A(p_input[28659]), .B(p_input[18659]), .Z(n1492) );
  AND U2985 ( .A(n1493), .B(p_input[8658]), .Z(o[8658]) );
  AND U2986 ( .A(p_input[28658]), .B(p_input[18658]), .Z(n1493) );
  AND U2987 ( .A(n1494), .B(p_input[8657]), .Z(o[8657]) );
  AND U2988 ( .A(p_input[28657]), .B(p_input[18657]), .Z(n1494) );
  AND U2989 ( .A(n1495), .B(p_input[8656]), .Z(o[8656]) );
  AND U2990 ( .A(p_input[28656]), .B(p_input[18656]), .Z(n1495) );
  AND U2991 ( .A(n1496), .B(p_input[8655]), .Z(o[8655]) );
  AND U2992 ( .A(p_input[28655]), .B(p_input[18655]), .Z(n1496) );
  AND U2993 ( .A(n1497), .B(p_input[8654]), .Z(o[8654]) );
  AND U2994 ( .A(p_input[28654]), .B(p_input[18654]), .Z(n1497) );
  AND U2995 ( .A(n1498), .B(p_input[8653]), .Z(o[8653]) );
  AND U2996 ( .A(p_input[28653]), .B(p_input[18653]), .Z(n1498) );
  AND U2997 ( .A(n1499), .B(p_input[8652]), .Z(o[8652]) );
  AND U2998 ( .A(p_input[28652]), .B(p_input[18652]), .Z(n1499) );
  AND U2999 ( .A(n1500), .B(p_input[8651]), .Z(o[8651]) );
  AND U3000 ( .A(p_input[28651]), .B(p_input[18651]), .Z(n1500) );
  AND U3001 ( .A(n1501), .B(p_input[8650]), .Z(o[8650]) );
  AND U3002 ( .A(p_input[28650]), .B(p_input[18650]), .Z(n1501) );
  AND U3003 ( .A(n1502), .B(p_input[864]), .Z(o[864]) );
  AND U3004 ( .A(p_input[20864]), .B(p_input[10864]), .Z(n1502) );
  AND U3005 ( .A(n1503), .B(p_input[8649]), .Z(o[8649]) );
  AND U3006 ( .A(p_input[28649]), .B(p_input[18649]), .Z(n1503) );
  AND U3007 ( .A(n1504), .B(p_input[8648]), .Z(o[8648]) );
  AND U3008 ( .A(p_input[28648]), .B(p_input[18648]), .Z(n1504) );
  AND U3009 ( .A(n1505), .B(p_input[8647]), .Z(o[8647]) );
  AND U3010 ( .A(p_input[28647]), .B(p_input[18647]), .Z(n1505) );
  AND U3011 ( .A(n1506), .B(p_input[8646]), .Z(o[8646]) );
  AND U3012 ( .A(p_input[28646]), .B(p_input[18646]), .Z(n1506) );
  AND U3013 ( .A(n1507), .B(p_input[8645]), .Z(o[8645]) );
  AND U3014 ( .A(p_input[28645]), .B(p_input[18645]), .Z(n1507) );
  AND U3015 ( .A(n1508), .B(p_input[8644]), .Z(o[8644]) );
  AND U3016 ( .A(p_input[28644]), .B(p_input[18644]), .Z(n1508) );
  AND U3017 ( .A(n1509), .B(p_input[8643]), .Z(o[8643]) );
  AND U3018 ( .A(p_input[28643]), .B(p_input[18643]), .Z(n1509) );
  AND U3019 ( .A(n1510), .B(p_input[8642]), .Z(o[8642]) );
  AND U3020 ( .A(p_input[28642]), .B(p_input[18642]), .Z(n1510) );
  AND U3021 ( .A(n1511), .B(p_input[8641]), .Z(o[8641]) );
  AND U3022 ( .A(p_input[28641]), .B(p_input[18641]), .Z(n1511) );
  AND U3023 ( .A(n1512), .B(p_input[8640]), .Z(o[8640]) );
  AND U3024 ( .A(p_input[28640]), .B(p_input[18640]), .Z(n1512) );
  AND U3025 ( .A(n1513), .B(p_input[863]), .Z(o[863]) );
  AND U3026 ( .A(p_input[20863]), .B(p_input[10863]), .Z(n1513) );
  AND U3027 ( .A(n1514), .B(p_input[8639]), .Z(o[8639]) );
  AND U3028 ( .A(p_input[28639]), .B(p_input[18639]), .Z(n1514) );
  AND U3029 ( .A(n1515), .B(p_input[8638]), .Z(o[8638]) );
  AND U3030 ( .A(p_input[28638]), .B(p_input[18638]), .Z(n1515) );
  AND U3031 ( .A(n1516), .B(p_input[8637]), .Z(o[8637]) );
  AND U3032 ( .A(p_input[28637]), .B(p_input[18637]), .Z(n1516) );
  AND U3033 ( .A(n1517), .B(p_input[8636]), .Z(o[8636]) );
  AND U3034 ( .A(p_input[28636]), .B(p_input[18636]), .Z(n1517) );
  AND U3035 ( .A(n1518), .B(p_input[8635]), .Z(o[8635]) );
  AND U3036 ( .A(p_input[28635]), .B(p_input[18635]), .Z(n1518) );
  AND U3037 ( .A(n1519), .B(p_input[8634]), .Z(o[8634]) );
  AND U3038 ( .A(p_input[28634]), .B(p_input[18634]), .Z(n1519) );
  AND U3039 ( .A(n1520), .B(p_input[8633]), .Z(o[8633]) );
  AND U3040 ( .A(p_input[28633]), .B(p_input[18633]), .Z(n1520) );
  AND U3041 ( .A(n1521), .B(p_input[8632]), .Z(o[8632]) );
  AND U3042 ( .A(p_input[28632]), .B(p_input[18632]), .Z(n1521) );
  AND U3043 ( .A(n1522), .B(p_input[8631]), .Z(o[8631]) );
  AND U3044 ( .A(p_input[28631]), .B(p_input[18631]), .Z(n1522) );
  AND U3045 ( .A(n1523), .B(p_input[8630]), .Z(o[8630]) );
  AND U3046 ( .A(p_input[28630]), .B(p_input[18630]), .Z(n1523) );
  AND U3047 ( .A(n1524), .B(p_input[862]), .Z(o[862]) );
  AND U3048 ( .A(p_input[20862]), .B(p_input[10862]), .Z(n1524) );
  AND U3049 ( .A(n1525), .B(p_input[8629]), .Z(o[8629]) );
  AND U3050 ( .A(p_input[28629]), .B(p_input[18629]), .Z(n1525) );
  AND U3051 ( .A(n1526), .B(p_input[8628]), .Z(o[8628]) );
  AND U3052 ( .A(p_input[28628]), .B(p_input[18628]), .Z(n1526) );
  AND U3053 ( .A(n1527), .B(p_input[8627]), .Z(o[8627]) );
  AND U3054 ( .A(p_input[28627]), .B(p_input[18627]), .Z(n1527) );
  AND U3055 ( .A(n1528), .B(p_input[8626]), .Z(o[8626]) );
  AND U3056 ( .A(p_input[28626]), .B(p_input[18626]), .Z(n1528) );
  AND U3057 ( .A(n1529), .B(p_input[8625]), .Z(o[8625]) );
  AND U3058 ( .A(p_input[28625]), .B(p_input[18625]), .Z(n1529) );
  AND U3059 ( .A(n1530), .B(p_input[8624]), .Z(o[8624]) );
  AND U3060 ( .A(p_input[28624]), .B(p_input[18624]), .Z(n1530) );
  AND U3061 ( .A(n1531), .B(p_input[8623]), .Z(o[8623]) );
  AND U3062 ( .A(p_input[28623]), .B(p_input[18623]), .Z(n1531) );
  AND U3063 ( .A(n1532), .B(p_input[8622]), .Z(o[8622]) );
  AND U3064 ( .A(p_input[28622]), .B(p_input[18622]), .Z(n1532) );
  AND U3065 ( .A(n1533), .B(p_input[8621]), .Z(o[8621]) );
  AND U3066 ( .A(p_input[28621]), .B(p_input[18621]), .Z(n1533) );
  AND U3067 ( .A(n1534), .B(p_input[8620]), .Z(o[8620]) );
  AND U3068 ( .A(p_input[28620]), .B(p_input[18620]), .Z(n1534) );
  AND U3069 ( .A(n1535), .B(p_input[861]), .Z(o[861]) );
  AND U3070 ( .A(p_input[20861]), .B(p_input[10861]), .Z(n1535) );
  AND U3071 ( .A(n1536), .B(p_input[8619]), .Z(o[8619]) );
  AND U3072 ( .A(p_input[28619]), .B(p_input[18619]), .Z(n1536) );
  AND U3073 ( .A(n1537), .B(p_input[8618]), .Z(o[8618]) );
  AND U3074 ( .A(p_input[28618]), .B(p_input[18618]), .Z(n1537) );
  AND U3075 ( .A(n1538), .B(p_input[8617]), .Z(o[8617]) );
  AND U3076 ( .A(p_input[28617]), .B(p_input[18617]), .Z(n1538) );
  AND U3077 ( .A(n1539), .B(p_input[8616]), .Z(o[8616]) );
  AND U3078 ( .A(p_input[28616]), .B(p_input[18616]), .Z(n1539) );
  AND U3079 ( .A(n1540), .B(p_input[8615]), .Z(o[8615]) );
  AND U3080 ( .A(p_input[28615]), .B(p_input[18615]), .Z(n1540) );
  AND U3081 ( .A(n1541), .B(p_input[8614]), .Z(o[8614]) );
  AND U3082 ( .A(p_input[28614]), .B(p_input[18614]), .Z(n1541) );
  AND U3083 ( .A(n1542), .B(p_input[8613]), .Z(o[8613]) );
  AND U3084 ( .A(p_input[28613]), .B(p_input[18613]), .Z(n1542) );
  AND U3085 ( .A(n1543), .B(p_input[8612]), .Z(o[8612]) );
  AND U3086 ( .A(p_input[28612]), .B(p_input[18612]), .Z(n1543) );
  AND U3087 ( .A(n1544), .B(p_input[8611]), .Z(o[8611]) );
  AND U3088 ( .A(p_input[28611]), .B(p_input[18611]), .Z(n1544) );
  AND U3089 ( .A(n1545), .B(p_input[8610]), .Z(o[8610]) );
  AND U3090 ( .A(p_input[28610]), .B(p_input[18610]), .Z(n1545) );
  AND U3091 ( .A(n1546), .B(p_input[860]), .Z(o[860]) );
  AND U3092 ( .A(p_input[20860]), .B(p_input[10860]), .Z(n1546) );
  AND U3093 ( .A(n1547), .B(p_input[8609]), .Z(o[8609]) );
  AND U3094 ( .A(p_input[28609]), .B(p_input[18609]), .Z(n1547) );
  AND U3095 ( .A(n1548), .B(p_input[8608]), .Z(o[8608]) );
  AND U3096 ( .A(p_input[28608]), .B(p_input[18608]), .Z(n1548) );
  AND U3097 ( .A(n1549), .B(p_input[8607]), .Z(o[8607]) );
  AND U3098 ( .A(p_input[28607]), .B(p_input[18607]), .Z(n1549) );
  AND U3099 ( .A(n1550), .B(p_input[8606]), .Z(o[8606]) );
  AND U3100 ( .A(p_input[28606]), .B(p_input[18606]), .Z(n1550) );
  AND U3101 ( .A(n1551), .B(p_input[8605]), .Z(o[8605]) );
  AND U3102 ( .A(p_input[28605]), .B(p_input[18605]), .Z(n1551) );
  AND U3103 ( .A(n1552), .B(p_input[8604]), .Z(o[8604]) );
  AND U3104 ( .A(p_input[28604]), .B(p_input[18604]), .Z(n1552) );
  AND U3105 ( .A(n1553), .B(p_input[8603]), .Z(o[8603]) );
  AND U3106 ( .A(p_input[28603]), .B(p_input[18603]), .Z(n1553) );
  AND U3107 ( .A(n1554), .B(p_input[8602]), .Z(o[8602]) );
  AND U3108 ( .A(p_input[28602]), .B(p_input[18602]), .Z(n1554) );
  AND U3109 ( .A(n1555), .B(p_input[8601]), .Z(o[8601]) );
  AND U3110 ( .A(p_input[28601]), .B(p_input[18601]), .Z(n1555) );
  AND U3111 ( .A(n1556), .B(p_input[8600]), .Z(o[8600]) );
  AND U3112 ( .A(p_input[28600]), .B(p_input[18600]), .Z(n1556) );
  AND U3113 ( .A(n1557), .B(p_input[85]), .Z(o[85]) );
  AND U3114 ( .A(p_input[20085]), .B(p_input[10085]), .Z(n1557) );
  AND U3115 ( .A(n1558), .B(p_input[859]), .Z(o[859]) );
  AND U3116 ( .A(p_input[20859]), .B(p_input[10859]), .Z(n1558) );
  AND U3117 ( .A(n1559), .B(p_input[8599]), .Z(o[8599]) );
  AND U3118 ( .A(p_input[28599]), .B(p_input[18599]), .Z(n1559) );
  AND U3119 ( .A(n1560), .B(p_input[8598]), .Z(o[8598]) );
  AND U3120 ( .A(p_input[28598]), .B(p_input[18598]), .Z(n1560) );
  AND U3121 ( .A(n1561), .B(p_input[8597]), .Z(o[8597]) );
  AND U3122 ( .A(p_input[28597]), .B(p_input[18597]), .Z(n1561) );
  AND U3123 ( .A(n1562), .B(p_input[8596]), .Z(o[8596]) );
  AND U3124 ( .A(p_input[28596]), .B(p_input[18596]), .Z(n1562) );
  AND U3125 ( .A(n1563), .B(p_input[8595]), .Z(o[8595]) );
  AND U3126 ( .A(p_input[28595]), .B(p_input[18595]), .Z(n1563) );
  AND U3127 ( .A(n1564), .B(p_input[8594]), .Z(o[8594]) );
  AND U3128 ( .A(p_input[28594]), .B(p_input[18594]), .Z(n1564) );
  AND U3129 ( .A(n1565), .B(p_input[8593]), .Z(o[8593]) );
  AND U3130 ( .A(p_input[28593]), .B(p_input[18593]), .Z(n1565) );
  AND U3131 ( .A(n1566), .B(p_input[8592]), .Z(o[8592]) );
  AND U3132 ( .A(p_input[28592]), .B(p_input[18592]), .Z(n1566) );
  AND U3133 ( .A(n1567), .B(p_input[8591]), .Z(o[8591]) );
  AND U3134 ( .A(p_input[28591]), .B(p_input[18591]), .Z(n1567) );
  AND U3135 ( .A(n1568), .B(p_input[8590]), .Z(o[8590]) );
  AND U3136 ( .A(p_input[28590]), .B(p_input[18590]), .Z(n1568) );
  AND U3137 ( .A(n1569), .B(p_input[858]), .Z(o[858]) );
  AND U3138 ( .A(p_input[20858]), .B(p_input[10858]), .Z(n1569) );
  AND U3139 ( .A(n1570), .B(p_input[8589]), .Z(o[8589]) );
  AND U3140 ( .A(p_input[28589]), .B(p_input[18589]), .Z(n1570) );
  AND U3141 ( .A(n1571), .B(p_input[8588]), .Z(o[8588]) );
  AND U3142 ( .A(p_input[28588]), .B(p_input[18588]), .Z(n1571) );
  AND U3143 ( .A(n1572), .B(p_input[8587]), .Z(o[8587]) );
  AND U3144 ( .A(p_input[28587]), .B(p_input[18587]), .Z(n1572) );
  AND U3145 ( .A(n1573), .B(p_input[8586]), .Z(o[8586]) );
  AND U3146 ( .A(p_input[28586]), .B(p_input[18586]), .Z(n1573) );
  AND U3147 ( .A(n1574), .B(p_input[8585]), .Z(o[8585]) );
  AND U3148 ( .A(p_input[28585]), .B(p_input[18585]), .Z(n1574) );
  AND U3149 ( .A(n1575), .B(p_input[8584]), .Z(o[8584]) );
  AND U3150 ( .A(p_input[28584]), .B(p_input[18584]), .Z(n1575) );
  AND U3151 ( .A(n1576), .B(p_input[8583]), .Z(o[8583]) );
  AND U3152 ( .A(p_input[28583]), .B(p_input[18583]), .Z(n1576) );
  AND U3153 ( .A(n1577), .B(p_input[8582]), .Z(o[8582]) );
  AND U3154 ( .A(p_input[28582]), .B(p_input[18582]), .Z(n1577) );
  AND U3155 ( .A(n1578), .B(p_input[8581]), .Z(o[8581]) );
  AND U3156 ( .A(p_input[28581]), .B(p_input[18581]), .Z(n1578) );
  AND U3157 ( .A(n1579), .B(p_input[8580]), .Z(o[8580]) );
  AND U3158 ( .A(p_input[28580]), .B(p_input[18580]), .Z(n1579) );
  AND U3159 ( .A(n1580), .B(p_input[857]), .Z(o[857]) );
  AND U3160 ( .A(p_input[20857]), .B(p_input[10857]), .Z(n1580) );
  AND U3161 ( .A(n1581), .B(p_input[8579]), .Z(o[8579]) );
  AND U3162 ( .A(p_input[28579]), .B(p_input[18579]), .Z(n1581) );
  AND U3163 ( .A(n1582), .B(p_input[8578]), .Z(o[8578]) );
  AND U3164 ( .A(p_input[28578]), .B(p_input[18578]), .Z(n1582) );
  AND U3165 ( .A(n1583), .B(p_input[8577]), .Z(o[8577]) );
  AND U3166 ( .A(p_input[28577]), .B(p_input[18577]), .Z(n1583) );
  AND U3167 ( .A(n1584), .B(p_input[8576]), .Z(o[8576]) );
  AND U3168 ( .A(p_input[28576]), .B(p_input[18576]), .Z(n1584) );
  AND U3169 ( .A(n1585), .B(p_input[8575]), .Z(o[8575]) );
  AND U3170 ( .A(p_input[28575]), .B(p_input[18575]), .Z(n1585) );
  AND U3171 ( .A(n1586), .B(p_input[8574]), .Z(o[8574]) );
  AND U3172 ( .A(p_input[28574]), .B(p_input[18574]), .Z(n1586) );
  AND U3173 ( .A(n1587), .B(p_input[8573]), .Z(o[8573]) );
  AND U3174 ( .A(p_input[28573]), .B(p_input[18573]), .Z(n1587) );
  AND U3175 ( .A(n1588), .B(p_input[8572]), .Z(o[8572]) );
  AND U3176 ( .A(p_input[28572]), .B(p_input[18572]), .Z(n1588) );
  AND U3177 ( .A(n1589), .B(p_input[8571]), .Z(o[8571]) );
  AND U3178 ( .A(p_input[28571]), .B(p_input[18571]), .Z(n1589) );
  AND U3179 ( .A(n1590), .B(p_input[8570]), .Z(o[8570]) );
  AND U3180 ( .A(p_input[28570]), .B(p_input[18570]), .Z(n1590) );
  AND U3181 ( .A(n1591), .B(p_input[856]), .Z(o[856]) );
  AND U3182 ( .A(p_input[20856]), .B(p_input[10856]), .Z(n1591) );
  AND U3183 ( .A(n1592), .B(p_input[8569]), .Z(o[8569]) );
  AND U3184 ( .A(p_input[28569]), .B(p_input[18569]), .Z(n1592) );
  AND U3185 ( .A(n1593), .B(p_input[8568]), .Z(o[8568]) );
  AND U3186 ( .A(p_input[28568]), .B(p_input[18568]), .Z(n1593) );
  AND U3187 ( .A(n1594), .B(p_input[8567]), .Z(o[8567]) );
  AND U3188 ( .A(p_input[28567]), .B(p_input[18567]), .Z(n1594) );
  AND U3189 ( .A(n1595), .B(p_input[8566]), .Z(o[8566]) );
  AND U3190 ( .A(p_input[28566]), .B(p_input[18566]), .Z(n1595) );
  AND U3191 ( .A(n1596), .B(p_input[8565]), .Z(o[8565]) );
  AND U3192 ( .A(p_input[28565]), .B(p_input[18565]), .Z(n1596) );
  AND U3193 ( .A(n1597), .B(p_input[8564]), .Z(o[8564]) );
  AND U3194 ( .A(p_input[28564]), .B(p_input[18564]), .Z(n1597) );
  AND U3195 ( .A(n1598), .B(p_input[8563]), .Z(o[8563]) );
  AND U3196 ( .A(p_input[28563]), .B(p_input[18563]), .Z(n1598) );
  AND U3197 ( .A(n1599), .B(p_input[8562]), .Z(o[8562]) );
  AND U3198 ( .A(p_input[28562]), .B(p_input[18562]), .Z(n1599) );
  AND U3199 ( .A(n1600), .B(p_input[8561]), .Z(o[8561]) );
  AND U3200 ( .A(p_input[28561]), .B(p_input[18561]), .Z(n1600) );
  AND U3201 ( .A(n1601), .B(p_input[8560]), .Z(o[8560]) );
  AND U3202 ( .A(p_input[28560]), .B(p_input[18560]), .Z(n1601) );
  AND U3203 ( .A(n1602), .B(p_input[855]), .Z(o[855]) );
  AND U3204 ( .A(p_input[20855]), .B(p_input[10855]), .Z(n1602) );
  AND U3205 ( .A(n1603), .B(p_input[8559]), .Z(o[8559]) );
  AND U3206 ( .A(p_input[28559]), .B(p_input[18559]), .Z(n1603) );
  AND U3207 ( .A(n1604), .B(p_input[8558]), .Z(o[8558]) );
  AND U3208 ( .A(p_input[28558]), .B(p_input[18558]), .Z(n1604) );
  AND U3209 ( .A(n1605), .B(p_input[8557]), .Z(o[8557]) );
  AND U3210 ( .A(p_input[28557]), .B(p_input[18557]), .Z(n1605) );
  AND U3211 ( .A(n1606), .B(p_input[8556]), .Z(o[8556]) );
  AND U3212 ( .A(p_input[28556]), .B(p_input[18556]), .Z(n1606) );
  AND U3213 ( .A(n1607), .B(p_input[8555]), .Z(o[8555]) );
  AND U3214 ( .A(p_input[28555]), .B(p_input[18555]), .Z(n1607) );
  AND U3215 ( .A(n1608), .B(p_input[8554]), .Z(o[8554]) );
  AND U3216 ( .A(p_input[28554]), .B(p_input[18554]), .Z(n1608) );
  AND U3217 ( .A(n1609), .B(p_input[8553]), .Z(o[8553]) );
  AND U3218 ( .A(p_input[28553]), .B(p_input[18553]), .Z(n1609) );
  AND U3219 ( .A(n1610), .B(p_input[8552]), .Z(o[8552]) );
  AND U3220 ( .A(p_input[28552]), .B(p_input[18552]), .Z(n1610) );
  AND U3221 ( .A(n1611), .B(p_input[8551]), .Z(o[8551]) );
  AND U3222 ( .A(p_input[28551]), .B(p_input[18551]), .Z(n1611) );
  AND U3223 ( .A(n1612), .B(p_input[8550]), .Z(o[8550]) );
  AND U3224 ( .A(p_input[28550]), .B(p_input[18550]), .Z(n1612) );
  AND U3225 ( .A(n1613), .B(p_input[854]), .Z(o[854]) );
  AND U3226 ( .A(p_input[20854]), .B(p_input[10854]), .Z(n1613) );
  AND U3227 ( .A(n1614), .B(p_input[8549]), .Z(o[8549]) );
  AND U3228 ( .A(p_input[28549]), .B(p_input[18549]), .Z(n1614) );
  AND U3229 ( .A(n1615), .B(p_input[8548]), .Z(o[8548]) );
  AND U3230 ( .A(p_input[28548]), .B(p_input[18548]), .Z(n1615) );
  AND U3231 ( .A(n1616), .B(p_input[8547]), .Z(o[8547]) );
  AND U3232 ( .A(p_input[28547]), .B(p_input[18547]), .Z(n1616) );
  AND U3233 ( .A(n1617), .B(p_input[8546]), .Z(o[8546]) );
  AND U3234 ( .A(p_input[28546]), .B(p_input[18546]), .Z(n1617) );
  AND U3235 ( .A(n1618), .B(p_input[8545]), .Z(o[8545]) );
  AND U3236 ( .A(p_input[28545]), .B(p_input[18545]), .Z(n1618) );
  AND U3237 ( .A(n1619), .B(p_input[8544]), .Z(o[8544]) );
  AND U3238 ( .A(p_input[28544]), .B(p_input[18544]), .Z(n1619) );
  AND U3239 ( .A(n1620), .B(p_input[8543]), .Z(o[8543]) );
  AND U3240 ( .A(p_input[28543]), .B(p_input[18543]), .Z(n1620) );
  AND U3241 ( .A(n1621), .B(p_input[8542]), .Z(o[8542]) );
  AND U3242 ( .A(p_input[28542]), .B(p_input[18542]), .Z(n1621) );
  AND U3243 ( .A(n1622), .B(p_input[8541]), .Z(o[8541]) );
  AND U3244 ( .A(p_input[28541]), .B(p_input[18541]), .Z(n1622) );
  AND U3245 ( .A(n1623), .B(p_input[8540]), .Z(o[8540]) );
  AND U3246 ( .A(p_input[28540]), .B(p_input[18540]), .Z(n1623) );
  AND U3247 ( .A(n1624), .B(p_input[853]), .Z(o[853]) );
  AND U3248 ( .A(p_input[20853]), .B(p_input[10853]), .Z(n1624) );
  AND U3249 ( .A(n1625), .B(p_input[8539]), .Z(o[8539]) );
  AND U3250 ( .A(p_input[28539]), .B(p_input[18539]), .Z(n1625) );
  AND U3251 ( .A(n1626), .B(p_input[8538]), .Z(o[8538]) );
  AND U3252 ( .A(p_input[28538]), .B(p_input[18538]), .Z(n1626) );
  AND U3253 ( .A(n1627), .B(p_input[8537]), .Z(o[8537]) );
  AND U3254 ( .A(p_input[28537]), .B(p_input[18537]), .Z(n1627) );
  AND U3255 ( .A(n1628), .B(p_input[8536]), .Z(o[8536]) );
  AND U3256 ( .A(p_input[28536]), .B(p_input[18536]), .Z(n1628) );
  AND U3257 ( .A(n1629), .B(p_input[8535]), .Z(o[8535]) );
  AND U3258 ( .A(p_input[28535]), .B(p_input[18535]), .Z(n1629) );
  AND U3259 ( .A(n1630), .B(p_input[8534]), .Z(o[8534]) );
  AND U3260 ( .A(p_input[28534]), .B(p_input[18534]), .Z(n1630) );
  AND U3261 ( .A(n1631), .B(p_input[8533]), .Z(o[8533]) );
  AND U3262 ( .A(p_input[28533]), .B(p_input[18533]), .Z(n1631) );
  AND U3263 ( .A(n1632), .B(p_input[8532]), .Z(o[8532]) );
  AND U3264 ( .A(p_input[28532]), .B(p_input[18532]), .Z(n1632) );
  AND U3265 ( .A(n1633), .B(p_input[8531]), .Z(o[8531]) );
  AND U3266 ( .A(p_input[28531]), .B(p_input[18531]), .Z(n1633) );
  AND U3267 ( .A(n1634), .B(p_input[8530]), .Z(o[8530]) );
  AND U3268 ( .A(p_input[28530]), .B(p_input[18530]), .Z(n1634) );
  AND U3269 ( .A(n1635), .B(p_input[852]), .Z(o[852]) );
  AND U3270 ( .A(p_input[20852]), .B(p_input[10852]), .Z(n1635) );
  AND U3271 ( .A(n1636), .B(p_input[8529]), .Z(o[8529]) );
  AND U3272 ( .A(p_input[28529]), .B(p_input[18529]), .Z(n1636) );
  AND U3273 ( .A(n1637), .B(p_input[8528]), .Z(o[8528]) );
  AND U3274 ( .A(p_input[28528]), .B(p_input[18528]), .Z(n1637) );
  AND U3275 ( .A(n1638), .B(p_input[8527]), .Z(o[8527]) );
  AND U3276 ( .A(p_input[28527]), .B(p_input[18527]), .Z(n1638) );
  AND U3277 ( .A(n1639), .B(p_input[8526]), .Z(o[8526]) );
  AND U3278 ( .A(p_input[28526]), .B(p_input[18526]), .Z(n1639) );
  AND U3279 ( .A(n1640), .B(p_input[8525]), .Z(o[8525]) );
  AND U3280 ( .A(p_input[28525]), .B(p_input[18525]), .Z(n1640) );
  AND U3281 ( .A(n1641), .B(p_input[8524]), .Z(o[8524]) );
  AND U3282 ( .A(p_input[28524]), .B(p_input[18524]), .Z(n1641) );
  AND U3283 ( .A(n1642), .B(p_input[8523]), .Z(o[8523]) );
  AND U3284 ( .A(p_input[28523]), .B(p_input[18523]), .Z(n1642) );
  AND U3285 ( .A(n1643), .B(p_input[8522]), .Z(o[8522]) );
  AND U3286 ( .A(p_input[28522]), .B(p_input[18522]), .Z(n1643) );
  AND U3287 ( .A(n1644), .B(p_input[8521]), .Z(o[8521]) );
  AND U3288 ( .A(p_input[28521]), .B(p_input[18521]), .Z(n1644) );
  AND U3289 ( .A(n1645), .B(p_input[8520]), .Z(o[8520]) );
  AND U3290 ( .A(p_input[28520]), .B(p_input[18520]), .Z(n1645) );
  AND U3291 ( .A(n1646), .B(p_input[851]), .Z(o[851]) );
  AND U3292 ( .A(p_input[20851]), .B(p_input[10851]), .Z(n1646) );
  AND U3293 ( .A(n1647), .B(p_input[8519]), .Z(o[8519]) );
  AND U3294 ( .A(p_input[28519]), .B(p_input[18519]), .Z(n1647) );
  AND U3295 ( .A(n1648), .B(p_input[8518]), .Z(o[8518]) );
  AND U3296 ( .A(p_input[28518]), .B(p_input[18518]), .Z(n1648) );
  AND U3297 ( .A(n1649), .B(p_input[8517]), .Z(o[8517]) );
  AND U3298 ( .A(p_input[28517]), .B(p_input[18517]), .Z(n1649) );
  AND U3299 ( .A(n1650), .B(p_input[8516]), .Z(o[8516]) );
  AND U3300 ( .A(p_input[28516]), .B(p_input[18516]), .Z(n1650) );
  AND U3301 ( .A(n1651), .B(p_input[8515]), .Z(o[8515]) );
  AND U3302 ( .A(p_input[28515]), .B(p_input[18515]), .Z(n1651) );
  AND U3303 ( .A(n1652), .B(p_input[8514]), .Z(o[8514]) );
  AND U3304 ( .A(p_input[28514]), .B(p_input[18514]), .Z(n1652) );
  AND U3305 ( .A(n1653), .B(p_input[8513]), .Z(o[8513]) );
  AND U3306 ( .A(p_input[28513]), .B(p_input[18513]), .Z(n1653) );
  AND U3307 ( .A(n1654), .B(p_input[8512]), .Z(o[8512]) );
  AND U3308 ( .A(p_input[28512]), .B(p_input[18512]), .Z(n1654) );
  AND U3309 ( .A(n1655), .B(p_input[8511]), .Z(o[8511]) );
  AND U3310 ( .A(p_input[28511]), .B(p_input[18511]), .Z(n1655) );
  AND U3311 ( .A(n1656), .B(p_input[8510]), .Z(o[8510]) );
  AND U3312 ( .A(p_input[28510]), .B(p_input[18510]), .Z(n1656) );
  AND U3313 ( .A(n1657), .B(p_input[850]), .Z(o[850]) );
  AND U3314 ( .A(p_input[20850]), .B(p_input[10850]), .Z(n1657) );
  AND U3315 ( .A(n1658), .B(p_input[8509]), .Z(o[8509]) );
  AND U3316 ( .A(p_input[28509]), .B(p_input[18509]), .Z(n1658) );
  AND U3317 ( .A(n1659), .B(p_input[8508]), .Z(o[8508]) );
  AND U3318 ( .A(p_input[28508]), .B(p_input[18508]), .Z(n1659) );
  AND U3319 ( .A(n1660), .B(p_input[8507]), .Z(o[8507]) );
  AND U3320 ( .A(p_input[28507]), .B(p_input[18507]), .Z(n1660) );
  AND U3321 ( .A(n1661), .B(p_input[8506]), .Z(o[8506]) );
  AND U3322 ( .A(p_input[28506]), .B(p_input[18506]), .Z(n1661) );
  AND U3323 ( .A(n1662), .B(p_input[8505]), .Z(o[8505]) );
  AND U3324 ( .A(p_input[28505]), .B(p_input[18505]), .Z(n1662) );
  AND U3325 ( .A(n1663), .B(p_input[8504]), .Z(o[8504]) );
  AND U3326 ( .A(p_input[28504]), .B(p_input[18504]), .Z(n1663) );
  AND U3327 ( .A(n1664), .B(p_input[8503]), .Z(o[8503]) );
  AND U3328 ( .A(p_input[28503]), .B(p_input[18503]), .Z(n1664) );
  AND U3329 ( .A(n1665), .B(p_input[8502]), .Z(o[8502]) );
  AND U3330 ( .A(p_input[28502]), .B(p_input[18502]), .Z(n1665) );
  AND U3331 ( .A(n1666), .B(p_input[8501]), .Z(o[8501]) );
  AND U3332 ( .A(p_input[28501]), .B(p_input[18501]), .Z(n1666) );
  AND U3333 ( .A(n1667), .B(p_input[8500]), .Z(o[8500]) );
  AND U3334 ( .A(p_input[28500]), .B(p_input[18500]), .Z(n1667) );
  AND U3335 ( .A(n1668), .B(p_input[84]), .Z(o[84]) );
  AND U3336 ( .A(p_input[20084]), .B(p_input[10084]), .Z(n1668) );
  AND U3337 ( .A(n1669), .B(p_input[849]), .Z(o[849]) );
  AND U3338 ( .A(p_input[20849]), .B(p_input[10849]), .Z(n1669) );
  AND U3339 ( .A(n1670), .B(p_input[8499]), .Z(o[8499]) );
  AND U3340 ( .A(p_input[28499]), .B(p_input[18499]), .Z(n1670) );
  AND U3341 ( .A(n1671), .B(p_input[8498]), .Z(o[8498]) );
  AND U3342 ( .A(p_input[28498]), .B(p_input[18498]), .Z(n1671) );
  AND U3343 ( .A(n1672), .B(p_input[8497]), .Z(o[8497]) );
  AND U3344 ( .A(p_input[28497]), .B(p_input[18497]), .Z(n1672) );
  AND U3345 ( .A(n1673), .B(p_input[8496]), .Z(o[8496]) );
  AND U3346 ( .A(p_input[28496]), .B(p_input[18496]), .Z(n1673) );
  AND U3347 ( .A(n1674), .B(p_input[8495]), .Z(o[8495]) );
  AND U3348 ( .A(p_input[28495]), .B(p_input[18495]), .Z(n1674) );
  AND U3349 ( .A(n1675), .B(p_input[8494]), .Z(o[8494]) );
  AND U3350 ( .A(p_input[28494]), .B(p_input[18494]), .Z(n1675) );
  AND U3351 ( .A(n1676), .B(p_input[8493]), .Z(o[8493]) );
  AND U3352 ( .A(p_input[28493]), .B(p_input[18493]), .Z(n1676) );
  AND U3353 ( .A(n1677), .B(p_input[8492]), .Z(o[8492]) );
  AND U3354 ( .A(p_input[28492]), .B(p_input[18492]), .Z(n1677) );
  AND U3355 ( .A(n1678), .B(p_input[8491]), .Z(o[8491]) );
  AND U3356 ( .A(p_input[28491]), .B(p_input[18491]), .Z(n1678) );
  AND U3357 ( .A(n1679), .B(p_input[8490]), .Z(o[8490]) );
  AND U3358 ( .A(p_input[28490]), .B(p_input[18490]), .Z(n1679) );
  AND U3359 ( .A(n1680), .B(p_input[848]), .Z(o[848]) );
  AND U3360 ( .A(p_input[20848]), .B(p_input[10848]), .Z(n1680) );
  AND U3361 ( .A(n1681), .B(p_input[8489]), .Z(o[8489]) );
  AND U3362 ( .A(p_input[28489]), .B(p_input[18489]), .Z(n1681) );
  AND U3363 ( .A(n1682), .B(p_input[8488]), .Z(o[8488]) );
  AND U3364 ( .A(p_input[28488]), .B(p_input[18488]), .Z(n1682) );
  AND U3365 ( .A(n1683), .B(p_input[8487]), .Z(o[8487]) );
  AND U3366 ( .A(p_input[28487]), .B(p_input[18487]), .Z(n1683) );
  AND U3367 ( .A(n1684), .B(p_input[8486]), .Z(o[8486]) );
  AND U3368 ( .A(p_input[28486]), .B(p_input[18486]), .Z(n1684) );
  AND U3369 ( .A(n1685), .B(p_input[8485]), .Z(o[8485]) );
  AND U3370 ( .A(p_input[28485]), .B(p_input[18485]), .Z(n1685) );
  AND U3371 ( .A(n1686), .B(p_input[8484]), .Z(o[8484]) );
  AND U3372 ( .A(p_input[28484]), .B(p_input[18484]), .Z(n1686) );
  AND U3373 ( .A(n1687), .B(p_input[8483]), .Z(o[8483]) );
  AND U3374 ( .A(p_input[28483]), .B(p_input[18483]), .Z(n1687) );
  AND U3375 ( .A(n1688), .B(p_input[8482]), .Z(o[8482]) );
  AND U3376 ( .A(p_input[28482]), .B(p_input[18482]), .Z(n1688) );
  AND U3377 ( .A(n1689), .B(p_input[8481]), .Z(o[8481]) );
  AND U3378 ( .A(p_input[28481]), .B(p_input[18481]), .Z(n1689) );
  AND U3379 ( .A(n1690), .B(p_input[8480]), .Z(o[8480]) );
  AND U3380 ( .A(p_input[28480]), .B(p_input[18480]), .Z(n1690) );
  AND U3381 ( .A(n1691), .B(p_input[847]), .Z(o[847]) );
  AND U3382 ( .A(p_input[20847]), .B(p_input[10847]), .Z(n1691) );
  AND U3383 ( .A(n1692), .B(p_input[8479]), .Z(o[8479]) );
  AND U3384 ( .A(p_input[28479]), .B(p_input[18479]), .Z(n1692) );
  AND U3385 ( .A(n1693), .B(p_input[8478]), .Z(o[8478]) );
  AND U3386 ( .A(p_input[28478]), .B(p_input[18478]), .Z(n1693) );
  AND U3387 ( .A(n1694), .B(p_input[8477]), .Z(o[8477]) );
  AND U3388 ( .A(p_input[28477]), .B(p_input[18477]), .Z(n1694) );
  AND U3389 ( .A(n1695), .B(p_input[8476]), .Z(o[8476]) );
  AND U3390 ( .A(p_input[28476]), .B(p_input[18476]), .Z(n1695) );
  AND U3391 ( .A(n1696), .B(p_input[8475]), .Z(o[8475]) );
  AND U3392 ( .A(p_input[28475]), .B(p_input[18475]), .Z(n1696) );
  AND U3393 ( .A(n1697), .B(p_input[8474]), .Z(o[8474]) );
  AND U3394 ( .A(p_input[28474]), .B(p_input[18474]), .Z(n1697) );
  AND U3395 ( .A(n1698), .B(p_input[8473]), .Z(o[8473]) );
  AND U3396 ( .A(p_input[28473]), .B(p_input[18473]), .Z(n1698) );
  AND U3397 ( .A(n1699), .B(p_input[8472]), .Z(o[8472]) );
  AND U3398 ( .A(p_input[28472]), .B(p_input[18472]), .Z(n1699) );
  AND U3399 ( .A(n1700), .B(p_input[8471]), .Z(o[8471]) );
  AND U3400 ( .A(p_input[28471]), .B(p_input[18471]), .Z(n1700) );
  AND U3401 ( .A(n1701), .B(p_input[8470]), .Z(o[8470]) );
  AND U3402 ( .A(p_input[28470]), .B(p_input[18470]), .Z(n1701) );
  AND U3403 ( .A(n1702), .B(p_input[846]), .Z(o[846]) );
  AND U3404 ( .A(p_input[20846]), .B(p_input[10846]), .Z(n1702) );
  AND U3405 ( .A(n1703), .B(p_input[8469]), .Z(o[8469]) );
  AND U3406 ( .A(p_input[28469]), .B(p_input[18469]), .Z(n1703) );
  AND U3407 ( .A(n1704), .B(p_input[8468]), .Z(o[8468]) );
  AND U3408 ( .A(p_input[28468]), .B(p_input[18468]), .Z(n1704) );
  AND U3409 ( .A(n1705), .B(p_input[8467]), .Z(o[8467]) );
  AND U3410 ( .A(p_input[28467]), .B(p_input[18467]), .Z(n1705) );
  AND U3411 ( .A(n1706), .B(p_input[8466]), .Z(o[8466]) );
  AND U3412 ( .A(p_input[28466]), .B(p_input[18466]), .Z(n1706) );
  AND U3413 ( .A(n1707), .B(p_input[8465]), .Z(o[8465]) );
  AND U3414 ( .A(p_input[28465]), .B(p_input[18465]), .Z(n1707) );
  AND U3415 ( .A(n1708), .B(p_input[8464]), .Z(o[8464]) );
  AND U3416 ( .A(p_input[28464]), .B(p_input[18464]), .Z(n1708) );
  AND U3417 ( .A(n1709), .B(p_input[8463]), .Z(o[8463]) );
  AND U3418 ( .A(p_input[28463]), .B(p_input[18463]), .Z(n1709) );
  AND U3419 ( .A(n1710), .B(p_input[8462]), .Z(o[8462]) );
  AND U3420 ( .A(p_input[28462]), .B(p_input[18462]), .Z(n1710) );
  AND U3421 ( .A(n1711), .B(p_input[8461]), .Z(o[8461]) );
  AND U3422 ( .A(p_input[28461]), .B(p_input[18461]), .Z(n1711) );
  AND U3423 ( .A(n1712), .B(p_input[8460]), .Z(o[8460]) );
  AND U3424 ( .A(p_input[28460]), .B(p_input[18460]), .Z(n1712) );
  AND U3425 ( .A(n1713), .B(p_input[845]), .Z(o[845]) );
  AND U3426 ( .A(p_input[20845]), .B(p_input[10845]), .Z(n1713) );
  AND U3427 ( .A(n1714), .B(p_input[8459]), .Z(o[8459]) );
  AND U3428 ( .A(p_input[28459]), .B(p_input[18459]), .Z(n1714) );
  AND U3429 ( .A(n1715), .B(p_input[8458]), .Z(o[8458]) );
  AND U3430 ( .A(p_input[28458]), .B(p_input[18458]), .Z(n1715) );
  AND U3431 ( .A(n1716), .B(p_input[8457]), .Z(o[8457]) );
  AND U3432 ( .A(p_input[28457]), .B(p_input[18457]), .Z(n1716) );
  AND U3433 ( .A(n1717), .B(p_input[8456]), .Z(o[8456]) );
  AND U3434 ( .A(p_input[28456]), .B(p_input[18456]), .Z(n1717) );
  AND U3435 ( .A(n1718), .B(p_input[8455]), .Z(o[8455]) );
  AND U3436 ( .A(p_input[28455]), .B(p_input[18455]), .Z(n1718) );
  AND U3437 ( .A(n1719), .B(p_input[8454]), .Z(o[8454]) );
  AND U3438 ( .A(p_input[28454]), .B(p_input[18454]), .Z(n1719) );
  AND U3439 ( .A(n1720), .B(p_input[8453]), .Z(o[8453]) );
  AND U3440 ( .A(p_input[28453]), .B(p_input[18453]), .Z(n1720) );
  AND U3441 ( .A(n1721), .B(p_input[8452]), .Z(o[8452]) );
  AND U3442 ( .A(p_input[28452]), .B(p_input[18452]), .Z(n1721) );
  AND U3443 ( .A(n1722), .B(p_input[8451]), .Z(o[8451]) );
  AND U3444 ( .A(p_input[28451]), .B(p_input[18451]), .Z(n1722) );
  AND U3445 ( .A(n1723), .B(p_input[8450]), .Z(o[8450]) );
  AND U3446 ( .A(p_input[28450]), .B(p_input[18450]), .Z(n1723) );
  AND U3447 ( .A(n1724), .B(p_input[844]), .Z(o[844]) );
  AND U3448 ( .A(p_input[20844]), .B(p_input[10844]), .Z(n1724) );
  AND U3449 ( .A(n1725), .B(p_input[8449]), .Z(o[8449]) );
  AND U3450 ( .A(p_input[28449]), .B(p_input[18449]), .Z(n1725) );
  AND U3451 ( .A(n1726), .B(p_input[8448]), .Z(o[8448]) );
  AND U3452 ( .A(p_input[28448]), .B(p_input[18448]), .Z(n1726) );
  AND U3453 ( .A(n1727), .B(p_input[8447]), .Z(o[8447]) );
  AND U3454 ( .A(p_input[28447]), .B(p_input[18447]), .Z(n1727) );
  AND U3455 ( .A(n1728), .B(p_input[8446]), .Z(o[8446]) );
  AND U3456 ( .A(p_input[28446]), .B(p_input[18446]), .Z(n1728) );
  AND U3457 ( .A(n1729), .B(p_input[8445]), .Z(o[8445]) );
  AND U3458 ( .A(p_input[28445]), .B(p_input[18445]), .Z(n1729) );
  AND U3459 ( .A(n1730), .B(p_input[8444]), .Z(o[8444]) );
  AND U3460 ( .A(p_input[28444]), .B(p_input[18444]), .Z(n1730) );
  AND U3461 ( .A(n1731), .B(p_input[8443]), .Z(o[8443]) );
  AND U3462 ( .A(p_input[28443]), .B(p_input[18443]), .Z(n1731) );
  AND U3463 ( .A(n1732), .B(p_input[8442]), .Z(o[8442]) );
  AND U3464 ( .A(p_input[28442]), .B(p_input[18442]), .Z(n1732) );
  AND U3465 ( .A(n1733), .B(p_input[8441]), .Z(o[8441]) );
  AND U3466 ( .A(p_input[28441]), .B(p_input[18441]), .Z(n1733) );
  AND U3467 ( .A(n1734), .B(p_input[8440]), .Z(o[8440]) );
  AND U3468 ( .A(p_input[28440]), .B(p_input[18440]), .Z(n1734) );
  AND U3469 ( .A(n1735), .B(p_input[843]), .Z(o[843]) );
  AND U3470 ( .A(p_input[20843]), .B(p_input[10843]), .Z(n1735) );
  AND U3471 ( .A(n1736), .B(p_input[8439]), .Z(o[8439]) );
  AND U3472 ( .A(p_input[28439]), .B(p_input[18439]), .Z(n1736) );
  AND U3473 ( .A(n1737), .B(p_input[8438]), .Z(o[8438]) );
  AND U3474 ( .A(p_input[28438]), .B(p_input[18438]), .Z(n1737) );
  AND U3475 ( .A(n1738), .B(p_input[8437]), .Z(o[8437]) );
  AND U3476 ( .A(p_input[28437]), .B(p_input[18437]), .Z(n1738) );
  AND U3477 ( .A(n1739), .B(p_input[8436]), .Z(o[8436]) );
  AND U3478 ( .A(p_input[28436]), .B(p_input[18436]), .Z(n1739) );
  AND U3479 ( .A(n1740), .B(p_input[8435]), .Z(o[8435]) );
  AND U3480 ( .A(p_input[28435]), .B(p_input[18435]), .Z(n1740) );
  AND U3481 ( .A(n1741), .B(p_input[8434]), .Z(o[8434]) );
  AND U3482 ( .A(p_input[28434]), .B(p_input[18434]), .Z(n1741) );
  AND U3483 ( .A(n1742), .B(p_input[8433]), .Z(o[8433]) );
  AND U3484 ( .A(p_input[28433]), .B(p_input[18433]), .Z(n1742) );
  AND U3485 ( .A(n1743), .B(p_input[8432]), .Z(o[8432]) );
  AND U3486 ( .A(p_input[28432]), .B(p_input[18432]), .Z(n1743) );
  AND U3487 ( .A(n1744), .B(p_input[8431]), .Z(o[8431]) );
  AND U3488 ( .A(p_input[28431]), .B(p_input[18431]), .Z(n1744) );
  AND U3489 ( .A(n1745), .B(p_input[8430]), .Z(o[8430]) );
  AND U3490 ( .A(p_input[28430]), .B(p_input[18430]), .Z(n1745) );
  AND U3491 ( .A(n1746), .B(p_input[842]), .Z(o[842]) );
  AND U3492 ( .A(p_input[20842]), .B(p_input[10842]), .Z(n1746) );
  AND U3493 ( .A(n1747), .B(p_input[8429]), .Z(o[8429]) );
  AND U3494 ( .A(p_input[28429]), .B(p_input[18429]), .Z(n1747) );
  AND U3495 ( .A(n1748), .B(p_input[8428]), .Z(o[8428]) );
  AND U3496 ( .A(p_input[28428]), .B(p_input[18428]), .Z(n1748) );
  AND U3497 ( .A(n1749), .B(p_input[8427]), .Z(o[8427]) );
  AND U3498 ( .A(p_input[28427]), .B(p_input[18427]), .Z(n1749) );
  AND U3499 ( .A(n1750), .B(p_input[8426]), .Z(o[8426]) );
  AND U3500 ( .A(p_input[28426]), .B(p_input[18426]), .Z(n1750) );
  AND U3501 ( .A(n1751), .B(p_input[8425]), .Z(o[8425]) );
  AND U3502 ( .A(p_input[28425]), .B(p_input[18425]), .Z(n1751) );
  AND U3503 ( .A(n1752), .B(p_input[8424]), .Z(o[8424]) );
  AND U3504 ( .A(p_input[28424]), .B(p_input[18424]), .Z(n1752) );
  AND U3505 ( .A(n1753), .B(p_input[8423]), .Z(o[8423]) );
  AND U3506 ( .A(p_input[28423]), .B(p_input[18423]), .Z(n1753) );
  AND U3507 ( .A(n1754), .B(p_input[8422]), .Z(o[8422]) );
  AND U3508 ( .A(p_input[28422]), .B(p_input[18422]), .Z(n1754) );
  AND U3509 ( .A(n1755), .B(p_input[8421]), .Z(o[8421]) );
  AND U3510 ( .A(p_input[28421]), .B(p_input[18421]), .Z(n1755) );
  AND U3511 ( .A(n1756), .B(p_input[8420]), .Z(o[8420]) );
  AND U3512 ( .A(p_input[28420]), .B(p_input[18420]), .Z(n1756) );
  AND U3513 ( .A(n1757), .B(p_input[841]), .Z(o[841]) );
  AND U3514 ( .A(p_input[20841]), .B(p_input[10841]), .Z(n1757) );
  AND U3515 ( .A(n1758), .B(p_input[8419]), .Z(o[8419]) );
  AND U3516 ( .A(p_input[28419]), .B(p_input[18419]), .Z(n1758) );
  AND U3517 ( .A(n1759), .B(p_input[8418]), .Z(o[8418]) );
  AND U3518 ( .A(p_input[28418]), .B(p_input[18418]), .Z(n1759) );
  AND U3519 ( .A(n1760), .B(p_input[8417]), .Z(o[8417]) );
  AND U3520 ( .A(p_input[28417]), .B(p_input[18417]), .Z(n1760) );
  AND U3521 ( .A(n1761), .B(p_input[8416]), .Z(o[8416]) );
  AND U3522 ( .A(p_input[28416]), .B(p_input[18416]), .Z(n1761) );
  AND U3523 ( .A(n1762), .B(p_input[8415]), .Z(o[8415]) );
  AND U3524 ( .A(p_input[28415]), .B(p_input[18415]), .Z(n1762) );
  AND U3525 ( .A(n1763), .B(p_input[8414]), .Z(o[8414]) );
  AND U3526 ( .A(p_input[28414]), .B(p_input[18414]), .Z(n1763) );
  AND U3527 ( .A(n1764), .B(p_input[8413]), .Z(o[8413]) );
  AND U3528 ( .A(p_input[28413]), .B(p_input[18413]), .Z(n1764) );
  AND U3529 ( .A(n1765), .B(p_input[8412]), .Z(o[8412]) );
  AND U3530 ( .A(p_input[28412]), .B(p_input[18412]), .Z(n1765) );
  AND U3531 ( .A(n1766), .B(p_input[8411]), .Z(o[8411]) );
  AND U3532 ( .A(p_input[28411]), .B(p_input[18411]), .Z(n1766) );
  AND U3533 ( .A(n1767), .B(p_input[8410]), .Z(o[8410]) );
  AND U3534 ( .A(p_input[28410]), .B(p_input[18410]), .Z(n1767) );
  AND U3535 ( .A(n1768), .B(p_input[840]), .Z(o[840]) );
  AND U3536 ( .A(p_input[20840]), .B(p_input[10840]), .Z(n1768) );
  AND U3537 ( .A(n1769), .B(p_input[8409]), .Z(o[8409]) );
  AND U3538 ( .A(p_input[28409]), .B(p_input[18409]), .Z(n1769) );
  AND U3539 ( .A(n1770), .B(p_input[8408]), .Z(o[8408]) );
  AND U3540 ( .A(p_input[28408]), .B(p_input[18408]), .Z(n1770) );
  AND U3541 ( .A(n1771), .B(p_input[8407]), .Z(o[8407]) );
  AND U3542 ( .A(p_input[28407]), .B(p_input[18407]), .Z(n1771) );
  AND U3543 ( .A(n1772), .B(p_input[8406]), .Z(o[8406]) );
  AND U3544 ( .A(p_input[28406]), .B(p_input[18406]), .Z(n1772) );
  AND U3545 ( .A(n1773), .B(p_input[8405]), .Z(o[8405]) );
  AND U3546 ( .A(p_input[28405]), .B(p_input[18405]), .Z(n1773) );
  AND U3547 ( .A(n1774), .B(p_input[8404]), .Z(o[8404]) );
  AND U3548 ( .A(p_input[28404]), .B(p_input[18404]), .Z(n1774) );
  AND U3549 ( .A(n1775), .B(p_input[8403]), .Z(o[8403]) );
  AND U3550 ( .A(p_input[28403]), .B(p_input[18403]), .Z(n1775) );
  AND U3551 ( .A(n1776), .B(p_input[8402]), .Z(o[8402]) );
  AND U3552 ( .A(p_input[28402]), .B(p_input[18402]), .Z(n1776) );
  AND U3553 ( .A(n1777), .B(p_input[8401]), .Z(o[8401]) );
  AND U3554 ( .A(p_input[28401]), .B(p_input[18401]), .Z(n1777) );
  AND U3555 ( .A(n1778), .B(p_input[8400]), .Z(o[8400]) );
  AND U3556 ( .A(p_input[28400]), .B(p_input[18400]), .Z(n1778) );
  AND U3557 ( .A(n1779), .B(p_input[83]), .Z(o[83]) );
  AND U3558 ( .A(p_input[20083]), .B(p_input[10083]), .Z(n1779) );
  AND U3559 ( .A(n1780), .B(p_input[839]), .Z(o[839]) );
  AND U3560 ( .A(p_input[20839]), .B(p_input[10839]), .Z(n1780) );
  AND U3561 ( .A(n1781), .B(p_input[8399]), .Z(o[8399]) );
  AND U3562 ( .A(p_input[28399]), .B(p_input[18399]), .Z(n1781) );
  AND U3563 ( .A(n1782), .B(p_input[8398]), .Z(o[8398]) );
  AND U3564 ( .A(p_input[28398]), .B(p_input[18398]), .Z(n1782) );
  AND U3565 ( .A(n1783), .B(p_input[8397]), .Z(o[8397]) );
  AND U3566 ( .A(p_input[28397]), .B(p_input[18397]), .Z(n1783) );
  AND U3567 ( .A(n1784), .B(p_input[8396]), .Z(o[8396]) );
  AND U3568 ( .A(p_input[28396]), .B(p_input[18396]), .Z(n1784) );
  AND U3569 ( .A(n1785), .B(p_input[8395]), .Z(o[8395]) );
  AND U3570 ( .A(p_input[28395]), .B(p_input[18395]), .Z(n1785) );
  AND U3571 ( .A(n1786), .B(p_input[8394]), .Z(o[8394]) );
  AND U3572 ( .A(p_input[28394]), .B(p_input[18394]), .Z(n1786) );
  AND U3573 ( .A(n1787), .B(p_input[8393]), .Z(o[8393]) );
  AND U3574 ( .A(p_input[28393]), .B(p_input[18393]), .Z(n1787) );
  AND U3575 ( .A(n1788), .B(p_input[8392]), .Z(o[8392]) );
  AND U3576 ( .A(p_input[28392]), .B(p_input[18392]), .Z(n1788) );
  AND U3577 ( .A(n1789), .B(p_input[8391]), .Z(o[8391]) );
  AND U3578 ( .A(p_input[28391]), .B(p_input[18391]), .Z(n1789) );
  AND U3579 ( .A(n1790), .B(p_input[8390]), .Z(o[8390]) );
  AND U3580 ( .A(p_input[28390]), .B(p_input[18390]), .Z(n1790) );
  AND U3581 ( .A(n1791), .B(p_input[838]), .Z(o[838]) );
  AND U3582 ( .A(p_input[20838]), .B(p_input[10838]), .Z(n1791) );
  AND U3583 ( .A(n1792), .B(p_input[8389]), .Z(o[8389]) );
  AND U3584 ( .A(p_input[28389]), .B(p_input[18389]), .Z(n1792) );
  AND U3585 ( .A(n1793), .B(p_input[8388]), .Z(o[8388]) );
  AND U3586 ( .A(p_input[28388]), .B(p_input[18388]), .Z(n1793) );
  AND U3587 ( .A(n1794), .B(p_input[8387]), .Z(o[8387]) );
  AND U3588 ( .A(p_input[28387]), .B(p_input[18387]), .Z(n1794) );
  AND U3589 ( .A(n1795), .B(p_input[8386]), .Z(o[8386]) );
  AND U3590 ( .A(p_input[28386]), .B(p_input[18386]), .Z(n1795) );
  AND U3591 ( .A(n1796), .B(p_input[8385]), .Z(o[8385]) );
  AND U3592 ( .A(p_input[28385]), .B(p_input[18385]), .Z(n1796) );
  AND U3593 ( .A(n1797), .B(p_input[8384]), .Z(o[8384]) );
  AND U3594 ( .A(p_input[28384]), .B(p_input[18384]), .Z(n1797) );
  AND U3595 ( .A(n1798), .B(p_input[8383]), .Z(o[8383]) );
  AND U3596 ( .A(p_input[28383]), .B(p_input[18383]), .Z(n1798) );
  AND U3597 ( .A(n1799), .B(p_input[8382]), .Z(o[8382]) );
  AND U3598 ( .A(p_input[28382]), .B(p_input[18382]), .Z(n1799) );
  AND U3599 ( .A(n1800), .B(p_input[8381]), .Z(o[8381]) );
  AND U3600 ( .A(p_input[28381]), .B(p_input[18381]), .Z(n1800) );
  AND U3601 ( .A(n1801), .B(p_input[8380]), .Z(o[8380]) );
  AND U3602 ( .A(p_input[28380]), .B(p_input[18380]), .Z(n1801) );
  AND U3603 ( .A(n1802), .B(p_input[837]), .Z(o[837]) );
  AND U3604 ( .A(p_input[20837]), .B(p_input[10837]), .Z(n1802) );
  AND U3605 ( .A(n1803), .B(p_input[8379]), .Z(o[8379]) );
  AND U3606 ( .A(p_input[28379]), .B(p_input[18379]), .Z(n1803) );
  AND U3607 ( .A(n1804), .B(p_input[8378]), .Z(o[8378]) );
  AND U3608 ( .A(p_input[28378]), .B(p_input[18378]), .Z(n1804) );
  AND U3609 ( .A(n1805), .B(p_input[8377]), .Z(o[8377]) );
  AND U3610 ( .A(p_input[28377]), .B(p_input[18377]), .Z(n1805) );
  AND U3611 ( .A(n1806), .B(p_input[8376]), .Z(o[8376]) );
  AND U3612 ( .A(p_input[28376]), .B(p_input[18376]), .Z(n1806) );
  AND U3613 ( .A(n1807), .B(p_input[8375]), .Z(o[8375]) );
  AND U3614 ( .A(p_input[28375]), .B(p_input[18375]), .Z(n1807) );
  AND U3615 ( .A(n1808), .B(p_input[8374]), .Z(o[8374]) );
  AND U3616 ( .A(p_input[28374]), .B(p_input[18374]), .Z(n1808) );
  AND U3617 ( .A(n1809), .B(p_input[8373]), .Z(o[8373]) );
  AND U3618 ( .A(p_input[28373]), .B(p_input[18373]), .Z(n1809) );
  AND U3619 ( .A(n1810), .B(p_input[8372]), .Z(o[8372]) );
  AND U3620 ( .A(p_input[28372]), .B(p_input[18372]), .Z(n1810) );
  AND U3621 ( .A(n1811), .B(p_input[8371]), .Z(o[8371]) );
  AND U3622 ( .A(p_input[28371]), .B(p_input[18371]), .Z(n1811) );
  AND U3623 ( .A(n1812), .B(p_input[8370]), .Z(o[8370]) );
  AND U3624 ( .A(p_input[28370]), .B(p_input[18370]), .Z(n1812) );
  AND U3625 ( .A(n1813), .B(p_input[836]), .Z(o[836]) );
  AND U3626 ( .A(p_input[20836]), .B(p_input[10836]), .Z(n1813) );
  AND U3627 ( .A(n1814), .B(p_input[8369]), .Z(o[8369]) );
  AND U3628 ( .A(p_input[28369]), .B(p_input[18369]), .Z(n1814) );
  AND U3629 ( .A(n1815), .B(p_input[8368]), .Z(o[8368]) );
  AND U3630 ( .A(p_input[28368]), .B(p_input[18368]), .Z(n1815) );
  AND U3631 ( .A(n1816), .B(p_input[8367]), .Z(o[8367]) );
  AND U3632 ( .A(p_input[28367]), .B(p_input[18367]), .Z(n1816) );
  AND U3633 ( .A(n1817), .B(p_input[8366]), .Z(o[8366]) );
  AND U3634 ( .A(p_input[28366]), .B(p_input[18366]), .Z(n1817) );
  AND U3635 ( .A(n1818), .B(p_input[8365]), .Z(o[8365]) );
  AND U3636 ( .A(p_input[28365]), .B(p_input[18365]), .Z(n1818) );
  AND U3637 ( .A(n1819), .B(p_input[8364]), .Z(o[8364]) );
  AND U3638 ( .A(p_input[28364]), .B(p_input[18364]), .Z(n1819) );
  AND U3639 ( .A(n1820), .B(p_input[8363]), .Z(o[8363]) );
  AND U3640 ( .A(p_input[28363]), .B(p_input[18363]), .Z(n1820) );
  AND U3641 ( .A(n1821), .B(p_input[8362]), .Z(o[8362]) );
  AND U3642 ( .A(p_input[28362]), .B(p_input[18362]), .Z(n1821) );
  AND U3643 ( .A(n1822), .B(p_input[8361]), .Z(o[8361]) );
  AND U3644 ( .A(p_input[28361]), .B(p_input[18361]), .Z(n1822) );
  AND U3645 ( .A(n1823), .B(p_input[8360]), .Z(o[8360]) );
  AND U3646 ( .A(p_input[28360]), .B(p_input[18360]), .Z(n1823) );
  AND U3647 ( .A(n1824), .B(p_input[835]), .Z(o[835]) );
  AND U3648 ( .A(p_input[20835]), .B(p_input[10835]), .Z(n1824) );
  AND U3649 ( .A(n1825), .B(p_input[8359]), .Z(o[8359]) );
  AND U3650 ( .A(p_input[28359]), .B(p_input[18359]), .Z(n1825) );
  AND U3651 ( .A(n1826), .B(p_input[8358]), .Z(o[8358]) );
  AND U3652 ( .A(p_input[28358]), .B(p_input[18358]), .Z(n1826) );
  AND U3653 ( .A(n1827), .B(p_input[8357]), .Z(o[8357]) );
  AND U3654 ( .A(p_input[28357]), .B(p_input[18357]), .Z(n1827) );
  AND U3655 ( .A(n1828), .B(p_input[8356]), .Z(o[8356]) );
  AND U3656 ( .A(p_input[28356]), .B(p_input[18356]), .Z(n1828) );
  AND U3657 ( .A(n1829), .B(p_input[8355]), .Z(o[8355]) );
  AND U3658 ( .A(p_input[28355]), .B(p_input[18355]), .Z(n1829) );
  AND U3659 ( .A(n1830), .B(p_input[8354]), .Z(o[8354]) );
  AND U3660 ( .A(p_input[28354]), .B(p_input[18354]), .Z(n1830) );
  AND U3661 ( .A(n1831), .B(p_input[8353]), .Z(o[8353]) );
  AND U3662 ( .A(p_input[28353]), .B(p_input[18353]), .Z(n1831) );
  AND U3663 ( .A(n1832), .B(p_input[8352]), .Z(o[8352]) );
  AND U3664 ( .A(p_input[28352]), .B(p_input[18352]), .Z(n1832) );
  AND U3665 ( .A(n1833), .B(p_input[8351]), .Z(o[8351]) );
  AND U3666 ( .A(p_input[28351]), .B(p_input[18351]), .Z(n1833) );
  AND U3667 ( .A(n1834), .B(p_input[8350]), .Z(o[8350]) );
  AND U3668 ( .A(p_input[28350]), .B(p_input[18350]), .Z(n1834) );
  AND U3669 ( .A(n1835), .B(p_input[834]), .Z(o[834]) );
  AND U3670 ( .A(p_input[20834]), .B(p_input[10834]), .Z(n1835) );
  AND U3671 ( .A(n1836), .B(p_input[8349]), .Z(o[8349]) );
  AND U3672 ( .A(p_input[28349]), .B(p_input[18349]), .Z(n1836) );
  AND U3673 ( .A(n1837), .B(p_input[8348]), .Z(o[8348]) );
  AND U3674 ( .A(p_input[28348]), .B(p_input[18348]), .Z(n1837) );
  AND U3675 ( .A(n1838), .B(p_input[8347]), .Z(o[8347]) );
  AND U3676 ( .A(p_input[28347]), .B(p_input[18347]), .Z(n1838) );
  AND U3677 ( .A(n1839), .B(p_input[8346]), .Z(o[8346]) );
  AND U3678 ( .A(p_input[28346]), .B(p_input[18346]), .Z(n1839) );
  AND U3679 ( .A(n1840), .B(p_input[8345]), .Z(o[8345]) );
  AND U3680 ( .A(p_input[28345]), .B(p_input[18345]), .Z(n1840) );
  AND U3681 ( .A(n1841), .B(p_input[8344]), .Z(o[8344]) );
  AND U3682 ( .A(p_input[28344]), .B(p_input[18344]), .Z(n1841) );
  AND U3683 ( .A(n1842), .B(p_input[8343]), .Z(o[8343]) );
  AND U3684 ( .A(p_input[28343]), .B(p_input[18343]), .Z(n1842) );
  AND U3685 ( .A(n1843), .B(p_input[8342]), .Z(o[8342]) );
  AND U3686 ( .A(p_input[28342]), .B(p_input[18342]), .Z(n1843) );
  AND U3687 ( .A(n1844), .B(p_input[8341]), .Z(o[8341]) );
  AND U3688 ( .A(p_input[28341]), .B(p_input[18341]), .Z(n1844) );
  AND U3689 ( .A(n1845), .B(p_input[8340]), .Z(o[8340]) );
  AND U3690 ( .A(p_input[28340]), .B(p_input[18340]), .Z(n1845) );
  AND U3691 ( .A(n1846), .B(p_input[833]), .Z(o[833]) );
  AND U3692 ( .A(p_input[20833]), .B(p_input[10833]), .Z(n1846) );
  AND U3693 ( .A(n1847), .B(p_input[8339]), .Z(o[8339]) );
  AND U3694 ( .A(p_input[28339]), .B(p_input[18339]), .Z(n1847) );
  AND U3695 ( .A(n1848), .B(p_input[8338]), .Z(o[8338]) );
  AND U3696 ( .A(p_input[28338]), .B(p_input[18338]), .Z(n1848) );
  AND U3697 ( .A(n1849), .B(p_input[8337]), .Z(o[8337]) );
  AND U3698 ( .A(p_input[28337]), .B(p_input[18337]), .Z(n1849) );
  AND U3699 ( .A(n1850), .B(p_input[8336]), .Z(o[8336]) );
  AND U3700 ( .A(p_input[28336]), .B(p_input[18336]), .Z(n1850) );
  AND U3701 ( .A(n1851), .B(p_input[8335]), .Z(o[8335]) );
  AND U3702 ( .A(p_input[28335]), .B(p_input[18335]), .Z(n1851) );
  AND U3703 ( .A(n1852), .B(p_input[8334]), .Z(o[8334]) );
  AND U3704 ( .A(p_input[28334]), .B(p_input[18334]), .Z(n1852) );
  AND U3705 ( .A(n1853), .B(p_input[8333]), .Z(o[8333]) );
  AND U3706 ( .A(p_input[28333]), .B(p_input[18333]), .Z(n1853) );
  AND U3707 ( .A(n1854), .B(p_input[8332]), .Z(o[8332]) );
  AND U3708 ( .A(p_input[28332]), .B(p_input[18332]), .Z(n1854) );
  AND U3709 ( .A(n1855), .B(p_input[8331]), .Z(o[8331]) );
  AND U3710 ( .A(p_input[28331]), .B(p_input[18331]), .Z(n1855) );
  AND U3711 ( .A(n1856), .B(p_input[8330]), .Z(o[8330]) );
  AND U3712 ( .A(p_input[28330]), .B(p_input[18330]), .Z(n1856) );
  AND U3713 ( .A(n1857), .B(p_input[832]), .Z(o[832]) );
  AND U3714 ( .A(p_input[20832]), .B(p_input[10832]), .Z(n1857) );
  AND U3715 ( .A(n1858), .B(p_input[8329]), .Z(o[8329]) );
  AND U3716 ( .A(p_input[28329]), .B(p_input[18329]), .Z(n1858) );
  AND U3717 ( .A(n1859), .B(p_input[8328]), .Z(o[8328]) );
  AND U3718 ( .A(p_input[28328]), .B(p_input[18328]), .Z(n1859) );
  AND U3719 ( .A(n1860), .B(p_input[8327]), .Z(o[8327]) );
  AND U3720 ( .A(p_input[28327]), .B(p_input[18327]), .Z(n1860) );
  AND U3721 ( .A(n1861), .B(p_input[8326]), .Z(o[8326]) );
  AND U3722 ( .A(p_input[28326]), .B(p_input[18326]), .Z(n1861) );
  AND U3723 ( .A(n1862), .B(p_input[8325]), .Z(o[8325]) );
  AND U3724 ( .A(p_input[28325]), .B(p_input[18325]), .Z(n1862) );
  AND U3725 ( .A(n1863), .B(p_input[8324]), .Z(o[8324]) );
  AND U3726 ( .A(p_input[28324]), .B(p_input[18324]), .Z(n1863) );
  AND U3727 ( .A(n1864), .B(p_input[8323]), .Z(o[8323]) );
  AND U3728 ( .A(p_input[28323]), .B(p_input[18323]), .Z(n1864) );
  AND U3729 ( .A(n1865), .B(p_input[8322]), .Z(o[8322]) );
  AND U3730 ( .A(p_input[28322]), .B(p_input[18322]), .Z(n1865) );
  AND U3731 ( .A(n1866), .B(p_input[8321]), .Z(o[8321]) );
  AND U3732 ( .A(p_input[28321]), .B(p_input[18321]), .Z(n1866) );
  AND U3733 ( .A(n1867), .B(p_input[8320]), .Z(o[8320]) );
  AND U3734 ( .A(p_input[28320]), .B(p_input[18320]), .Z(n1867) );
  AND U3735 ( .A(n1868), .B(p_input[831]), .Z(o[831]) );
  AND U3736 ( .A(p_input[20831]), .B(p_input[10831]), .Z(n1868) );
  AND U3737 ( .A(n1869), .B(p_input[8319]), .Z(o[8319]) );
  AND U3738 ( .A(p_input[28319]), .B(p_input[18319]), .Z(n1869) );
  AND U3739 ( .A(n1870), .B(p_input[8318]), .Z(o[8318]) );
  AND U3740 ( .A(p_input[28318]), .B(p_input[18318]), .Z(n1870) );
  AND U3741 ( .A(n1871), .B(p_input[8317]), .Z(o[8317]) );
  AND U3742 ( .A(p_input[28317]), .B(p_input[18317]), .Z(n1871) );
  AND U3743 ( .A(n1872), .B(p_input[8316]), .Z(o[8316]) );
  AND U3744 ( .A(p_input[28316]), .B(p_input[18316]), .Z(n1872) );
  AND U3745 ( .A(n1873), .B(p_input[8315]), .Z(o[8315]) );
  AND U3746 ( .A(p_input[28315]), .B(p_input[18315]), .Z(n1873) );
  AND U3747 ( .A(n1874), .B(p_input[8314]), .Z(o[8314]) );
  AND U3748 ( .A(p_input[28314]), .B(p_input[18314]), .Z(n1874) );
  AND U3749 ( .A(n1875), .B(p_input[8313]), .Z(o[8313]) );
  AND U3750 ( .A(p_input[28313]), .B(p_input[18313]), .Z(n1875) );
  AND U3751 ( .A(n1876), .B(p_input[8312]), .Z(o[8312]) );
  AND U3752 ( .A(p_input[28312]), .B(p_input[18312]), .Z(n1876) );
  AND U3753 ( .A(n1877), .B(p_input[8311]), .Z(o[8311]) );
  AND U3754 ( .A(p_input[28311]), .B(p_input[18311]), .Z(n1877) );
  AND U3755 ( .A(n1878), .B(p_input[8310]), .Z(o[8310]) );
  AND U3756 ( .A(p_input[28310]), .B(p_input[18310]), .Z(n1878) );
  AND U3757 ( .A(n1879), .B(p_input[830]), .Z(o[830]) );
  AND U3758 ( .A(p_input[20830]), .B(p_input[10830]), .Z(n1879) );
  AND U3759 ( .A(n1880), .B(p_input[8309]), .Z(o[8309]) );
  AND U3760 ( .A(p_input[28309]), .B(p_input[18309]), .Z(n1880) );
  AND U3761 ( .A(n1881), .B(p_input[8308]), .Z(o[8308]) );
  AND U3762 ( .A(p_input[28308]), .B(p_input[18308]), .Z(n1881) );
  AND U3763 ( .A(n1882), .B(p_input[8307]), .Z(o[8307]) );
  AND U3764 ( .A(p_input[28307]), .B(p_input[18307]), .Z(n1882) );
  AND U3765 ( .A(n1883), .B(p_input[8306]), .Z(o[8306]) );
  AND U3766 ( .A(p_input[28306]), .B(p_input[18306]), .Z(n1883) );
  AND U3767 ( .A(n1884), .B(p_input[8305]), .Z(o[8305]) );
  AND U3768 ( .A(p_input[28305]), .B(p_input[18305]), .Z(n1884) );
  AND U3769 ( .A(n1885), .B(p_input[8304]), .Z(o[8304]) );
  AND U3770 ( .A(p_input[28304]), .B(p_input[18304]), .Z(n1885) );
  AND U3771 ( .A(n1886), .B(p_input[8303]), .Z(o[8303]) );
  AND U3772 ( .A(p_input[28303]), .B(p_input[18303]), .Z(n1886) );
  AND U3773 ( .A(n1887), .B(p_input[8302]), .Z(o[8302]) );
  AND U3774 ( .A(p_input[28302]), .B(p_input[18302]), .Z(n1887) );
  AND U3775 ( .A(n1888), .B(p_input[8301]), .Z(o[8301]) );
  AND U3776 ( .A(p_input[28301]), .B(p_input[18301]), .Z(n1888) );
  AND U3777 ( .A(n1889), .B(p_input[8300]), .Z(o[8300]) );
  AND U3778 ( .A(p_input[28300]), .B(p_input[18300]), .Z(n1889) );
  AND U3779 ( .A(n1890), .B(p_input[82]), .Z(o[82]) );
  AND U3780 ( .A(p_input[20082]), .B(p_input[10082]), .Z(n1890) );
  AND U3781 ( .A(n1891), .B(p_input[829]), .Z(o[829]) );
  AND U3782 ( .A(p_input[20829]), .B(p_input[10829]), .Z(n1891) );
  AND U3783 ( .A(n1892), .B(p_input[8299]), .Z(o[8299]) );
  AND U3784 ( .A(p_input[28299]), .B(p_input[18299]), .Z(n1892) );
  AND U3785 ( .A(n1893), .B(p_input[8298]), .Z(o[8298]) );
  AND U3786 ( .A(p_input[28298]), .B(p_input[18298]), .Z(n1893) );
  AND U3787 ( .A(n1894), .B(p_input[8297]), .Z(o[8297]) );
  AND U3788 ( .A(p_input[28297]), .B(p_input[18297]), .Z(n1894) );
  AND U3789 ( .A(n1895), .B(p_input[8296]), .Z(o[8296]) );
  AND U3790 ( .A(p_input[28296]), .B(p_input[18296]), .Z(n1895) );
  AND U3791 ( .A(n1896), .B(p_input[8295]), .Z(o[8295]) );
  AND U3792 ( .A(p_input[28295]), .B(p_input[18295]), .Z(n1896) );
  AND U3793 ( .A(n1897), .B(p_input[8294]), .Z(o[8294]) );
  AND U3794 ( .A(p_input[28294]), .B(p_input[18294]), .Z(n1897) );
  AND U3795 ( .A(n1898), .B(p_input[8293]), .Z(o[8293]) );
  AND U3796 ( .A(p_input[28293]), .B(p_input[18293]), .Z(n1898) );
  AND U3797 ( .A(n1899), .B(p_input[8292]), .Z(o[8292]) );
  AND U3798 ( .A(p_input[28292]), .B(p_input[18292]), .Z(n1899) );
  AND U3799 ( .A(n1900), .B(p_input[8291]), .Z(o[8291]) );
  AND U3800 ( .A(p_input[28291]), .B(p_input[18291]), .Z(n1900) );
  AND U3801 ( .A(n1901), .B(p_input[8290]), .Z(o[8290]) );
  AND U3802 ( .A(p_input[28290]), .B(p_input[18290]), .Z(n1901) );
  AND U3803 ( .A(n1902), .B(p_input[828]), .Z(o[828]) );
  AND U3804 ( .A(p_input[20828]), .B(p_input[10828]), .Z(n1902) );
  AND U3805 ( .A(n1903), .B(p_input[8289]), .Z(o[8289]) );
  AND U3806 ( .A(p_input[28289]), .B(p_input[18289]), .Z(n1903) );
  AND U3807 ( .A(n1904), .B(p_input[8288]), .Z(o[8288]) );
  AND U3808 ( .A(p_input[28288]), .B(p_input[18288]), .Z(n1904) );
  AND U3809 ( .A(n1905), .B(p_input[8287]), .Z(o[8287]) );
  AND U3810 ( .A(p_input[28287]), .B(p_input[18287]), .Z(n1905) );
  AND U3811 ( .A(n1906), .B(p_input[8286]), .Z(o[8286]) );
  AND U3812 ( .A(p_input[28286]), .B(p_input[18286]), .Z(n1906) );
  AND U3813 ( .A(n1907), .B(p_input[8285]), .Z(o[8285]) );
  AND U3814 ( .A(p_input[28285]), .B(p_input[18285]), .Z(n1907) );
  AND U3815 ( .A(n1908), .B(p_input[8284]), .Z(o[8284]) );
  AND U3816 ( .A(p_input[28284]), .B(p_input[18284]), .Z(n1908) );
  AND U3817 ( .A(n1909), .B(p_input[8283]), .Z(o[8283]) );
  AND U3818 ( .A(p_input[28283]), .B(p_input[18283]), .Z(n1909) );
  AND U3819 ( .A(n1910), .B(p_input[8282]), .Z(o[8282]) );
  AND U3820 ( .A(p_input[28282]), .B(p_input[18282]), .Z(n1910) );
  AND U3821 ( .A(n1911), .B(p_input[8281]), .Z(o[8281]) );
  AND U3822 ( .A(p_input[28281]), .B(p_input[18281]), .Z(n1911) );
  AND U3823 ( .A(n1912), .B(p_input[8280]), .Z(o[8280]) );
  AND U3824 ( .A(p_input[28280]), .B(p_input[18280]), .Z(n1912) );
  AND U3825 ( .A(n1913), .B(p_input[827]), .Z(o[827]) );
  AND U3826 ( .A(p_input[20827]), .B(p_input[10827]), .Z(n1913) );
  AND U3827 ( .A(n1914), .B(p_input[8279]), .Z(o[8279]) );
  AND U3828 ( .A(p_input[28279]), .B(p_input[18279]), .Z(n1914) );
  AND U3829 ( .A(n1915), .B(p_input[8278]), .Z(o[8278]) );
  AND U3830 ( .A(p_input[28278]), .B(p_input[18278]), .Z(n1915) );
  AND U3831 ( .A(n1916), .B(p_input[8277]), .Z(o[8277]) );
  AND U3832 ( .A(p_input[28277]), .B(p_input[18277]), .Z(n1916) );
  AND U3833 ( .A(n1917), .B(p_input[8276]), .Z(o[8276]) );
  AND U3834 ( .A(p_input[28276]), .B(p_input[18276]), .Z(n1917) );
  AND U3835 ( .A(n1918), .B(p_input[8275]), .Z(o[8275]) );
  AND U3836 ( .A(p_input[28275]), .B(p_input[18275]), .Z(n1918) );
  AND U3837 ( .A(n1919), .B(p_input[8274]), .Z(o[8274]) );
  AND U3838 ( .A(p_input[28274]), .B(p_input[18274]), .Z(n1919) );
  AND U3839 ( .A(n1920), .B(p_input[8273]), .Z(o[8273]) );
  AND U3840 ( .A(p_input[28273]), .B(p_input[18273]), .Z(n1920) );
  AND U3841 ( .A(n1921), .B(p_input[8272]), .Z(o[8272]) );
  AND U3842 ( .A(p_input[28272]), .B(p_input[18272]), .Z(n1921) );
  AND U3843 ( .A(n1922), .B(p_input[8271]), .Z(o[8271]) );
  AND U3844 ( .A(p_input[28271]), .B(p_input[18271]), .Z(n1922) );
  AND U3845 ( .A(n1923), .B(p_input[8270]), .Z(o[8270]) );
  AND U3846 ( .A(p_input[28270]), .B(p_input[18270]), .Z(n1923) );
  AND U3847 ( .A(n1924), .B(p_input[826]), .Z(o[826]) );
  AND U3848 ( .A(p_input[20826]), .B(p_input[10826]), .Z(n1924) );
  AND U3849 ( .A(n1925), .B(p_input[8269]), .Z(o[8269]) );
  AND U3850 ( .A(p_input[28269]), .B(p_input[18269]), .Z(n1925) );
  AND U3851 ( .A(n1926), .B(p_input[8268]), .Z(o[8268]) );
  AND U3852 ( .A(p_input[28268]), .B(p_input[18268]), .Z(n1926) );
  AND U3853 ( .A(n1927), .B(p_input[8267]), .Z(o[8267]) );
  AND U3854 ( .A(p_input[28267]), .B(p_input[18267]), .Z(n1927) );
  AND U3855 ( .A(n1928), .B(p_input[8266]), .Z(o[8266]) );
  AND U3856 ( .A(p_input[28266]), .B(p_input[18266]), .Z(n1928) );
  AND U3857 ( .A(n1929), .B(p_input[8265]), .Z(o[8265]) );
  AND U3858 ( .A(p_input[28265]), .B(p_input[18265]), .Z(n1929) );
  AND U3859 ( .A(n1930), .B(p_input[8264]), .Z(o[8264]) );
  AND U3860 ( .A(p_input[28264]), .B(p_input[18264]), .Z(n1930) );
  AND U3861 ( .A(n1931), .B(p_input[8263]), .Z(o[8263]) );
  AND U3862 ( .A(p_input[28263]), .B(p_input[18263]), .Z(n1931) );
  AND U3863 ( .A(n1932), .B(p_input[8262]), .Z(o[8262]) );
  AND U3864 ( .A(p_input[28262]), .B(p_input[18262]), .Z(n1932) );
  AND U3865 ( .A(n1933), .B(p_input[8261]), .Z(o[8261]) );
  AND U3866 ( .A(p_input[28261]), .B(p_input[18261]), .Z(n1933) );
  AND U3867 ( .A(n1934), .B(p_input[8260]), .Z(o[8260]) );
  AND U3868 ( .A(p_input[28260]), .B(p_input[18260]), .Z(n1934) );
  AND U3869 ( .A(n1935), .B(p_input[825]), .Z(o[825]) );
  AND U3870 ( .A(p_input[20825]), .B(p_input[10825]), .Z(n1935) );
  AND U3871 ( .A(n1936), .B(p_input[8259]), .Z(o[8259]) );
  AND U3872 ( .A(p_input[28259]), .B(p_input[18259]), .Z(n1936) );
  AND U3873 ( .A(n1937), .B(p_input[8258]), .Z(o[8258]) );
  AND U3874 ( .A(p_input[28258]), .B(p_input[18258]), .Z(n1937) );
  AND U3875 ( .A(n1938), .B(p_input[8257]), .Z(o[8257]) );
  AND U3876 ( .A(p_input[28257]), .B(p_input[18257]), .Z(n1938) );
  AND U3877 ( .A(n1939), .B(p_input[8256]), .Z(o[8256]) );
  AND U3878 ( .A(p_input[28256]), .B(p_input[18256]), .Z(n1939) );
  AND U3879 ( .A(n1940), .B(p_input[8255]), .Z(o[8255]) );
  AND U3880 ( .A(p_input[28255]), .B(p_input[18255]), .Z(n1940) );
  AND U3881 ( .A(n1941), .B(p_input[8254]), .Z(o[8254]) );
  AND U3882 ( .A(p_input[28254]), .B(p_input[18254]), .Z(n1941) );
  AND U3883 ( .A(n1942), .B(p_input[8253]), .Z(o[8253]) );
  AND U3884 ( .A(p_input[28253]), .B(p_input[18253]), .Z(n1942) );
  AND U3885 ( .A(n1943), .B(p_input[8252]), .Z(o[8252]) );
  AND U3886 ( .A(p_input[28252]), .B(p_input[18252]), .Z(n1943) );
  AND U3887 ( .A(n1944), .B(p_input[8251]), .Z(o[8251]) );
  AND U3888 ( .A(p_input[28251]), .B(p_input[18251]), .Z(n1944) );
  AND U3889 ( .A(n1945), .B(p_input[8250]), .Z(o[8250]) );
  AND U3890 ( .A(p_input[28250]), .B(p_input[18250]), .Z(n1945) );
  AND U3891 ( .A(n1946), .B(p_input[824]), .Z(o[824]) );
  AND U3892 ( .A(p_input[20824]), .B(p_input[10824]), .Z(n1946) );
  AND U3893 ( .A(n1947), .B(p_input[8249]), .Z(o[8249]) );
  AND U3894 ( .A(p_input[28249]), .B(p_input[18249]), .Z(n1947) );
  AND U3895 ( .A(n1948), .B(p_input[8248]), .Z(o[8248]) );
  AND U3896 ( .A(p_input[28248]), .B(p_input[18248]), .Z(n1948) );
  AND U3897 ( .A(n1949), .B(p_input[8247]), .Z(o[8247]) );
  AND U3898 ( .A(p_input[28247]), .B(p_input[18247]), .Z(n1949) );
  AND U3899 ( .A(n1950), .B(p_input[8246]), .Z(o[8246]) );
  AND U3900 ( .A(p_input[28246]), .B(p_input[18246]), .Z(n1950) );
  AND U3901 ( .A(n1951), .B(p_input[8245]), .Z(o[8245]) );
  AND U3902 ( .A(p_input[28245]), .B(p_input[18245]), .Z(n1951) );
  AND U3903 ( .A(n1952), .B(p_input[8244]), .Z(o[8244]) );
  AND U3904 ( .A(p_input[28244]), .B(p_input[18244]), .Z(n1952) );
  AND U3905 ( .A(n1953), .B(p_input[8243]), .Z(o[8243]) );
  AND U3906 ( .A(p_input[28243]), .B(p_input[18243]), .Z(n1953) );
  AND U3907 ( .A(n1954), .B(p_input[8242]), .Z(o[8242]) );
  AND U3908 ( .A(p_input[28242]), .B(p_input[18242]), .Z(n1954) );
  AND U3909 ( .A(n1955), .B(p_input[8241]), .Z(o[8241]) );
  AND U3910 ( .A(p_input[28241]), .B(p_input[18241]), .Z(n1955) );
  AND U3911 ( .A(n1956), .B(p_input[8240]), .Z(o[8240]) );
  AND U3912 ( .A(p_input[28240]), .B(p_input[18240]), .Z(n1956) );
  AND U3913 ( .A(n1957), .B(p_input[823]), .Z(o[823]) );
  AND U3914 ( .A(p_input[20823]), .B(p_input[10823]), .Z(n1957) );
  AND U3915 ( .A(n1958), .B(p_input[8239]), .Z(o[8239]) );
  AND U3916 ( .A(p_input[28239]), .B(p_input[18239]), .Z(n1958) );
  AND U3917 ( .A(n1959), .B(p_input[8238]), .Z(o[8238]) );
  AND U3918 ( .A(p_input[28238]), .B(p_input[18238]), .Z(n1959) );
  AND U3919 ( .A(n1960), .B(p_input[8237]), .Z(o[8237]) );
  AND U3920 ( .A(p_input[28237]), .B(p_input[18237]), .Z(n1960) );
  AND U3921 ( .A(n1961), .B(p_input[8236]), .Z(o[8236]) );
  AND U3922 ( .A(p_input[28236]), .B(p_input[18236]), .Z(n1961) );
  AND U3923 ( .A(n1962), .B(p_input[8235]), .Z(o[8235]) );
  AND U3924 ( .A(p_input[28235]), .B(p_input[18235]), .Z(n1962) );
  AND U3925 ( .A(n1963), .B(p_input[8234]), .Z(o[8234]) );
  AND U3926 ( .A(p_input[28234]), .B(p_input[18234]), .Z(n1963) );
  AND U3927 ( .A(n1964), .B(p_input[8233]), .Z(o[8233]) );
  AND U3928 ( .A(p_input[28233]), .B(p_input[18233]), .Z(n1964) );
  AND U3929 ( .A(n1965), .B(p_input[8232]), .Z(o[8232]) );
  AND U3930 ( .A(p_input[28232]), .B(p_input[18232]), .Z(n1965) );
  AND U3931 ( .A(n1966), .B(p_input[8231]), .Z(o[8231]) );
  AND U3932 ( .A(p_input[28231]), .B(p_input[18231]), .Z(n1966) );
  AND U3933 ( .A(n1967), .B(p_input[8230]), .Z(o[8230]) );
  AND U3934 ( .A(p_input[28230]), .B(p_input[18230]), .Z(n1967) );
  AND U3935 ( .A(n1968), .B(p_input[822]), .Z(o[822]) );
  AND U3936 ( .A(p_input[20822]), .B(p_input[10822]), .Z(n1968) );
  AND U3937 ( .A(n1969), .B(p_input[8229]), .Z(o[8229]) );
  AND U3938 ( .A(p_input[28229]), .B(p_input[18229]), .Z(n1969) );
  AND U3939 ( .A(n1970), .B(p_input[8228]), .Z(o[8228]) );
  AND U3940 ( .A(p_input[28228]), .B(p_input[18228]), .Z(n1970) );
  AND U3941 ( .A(n1971), .B(p_input[8227]), .Z(o[8227]) );
  AND U3942 ( .A(p_input[28227]), .B(p_input[18227]), .Z(n1971) );
  AND U3943 ( .A(n1972), .B(p_input[8226]), .Z(o[8226]) );
  AND U3944 ( .A(p_input[28226]), .B(p_input[18226]), .Z(n1972) );
  AND U3945 ( .A(n1973), .B(p_input[8225]), .Z(o[8225]) );
  AND U3946 ( .A(p_input[28225]), .B(p_input[18225]), .Z(n1973) );
  AND U3947 ( .A(n1974), .B(p_input[8224]), .Z(o[8224]) );
  AND U3948 ( .A(p_input[28224]), .B(p_input[18224]), .Z(n1974) );
  AND U3949 ( .A(n1975), .B(p_input[8223]), .Z(o[8223]) );
  AND U3950 ( .A(p_input[28223]), .B(p_input[18223]), .Z(n1975) );
  AND U3951 ( .A(n1976), .B(p_input[8222]), .Z(o[8222]) );
  AND U3952 ( .A(p_input[28222]), .B(p_input[18222]), .Z(n1976) );
  AND U3953 ( .A(n1977), .B(p_input[8221]), .Z(o[8221]) );
  AND U3954 ( .A(p_input[28221]), .B(p_input[18221]), .Z(n1977) );
  AND U3955 ( .A(n1978), .B(p_input[8220]), .Z(o[8220]) );
  AND U3956 ( .A(p_input[28220]), .B(p_input[18220]), .Z(n1978) );
  AND U3957 ( .A(n1979), .B(p_input[821]), .Z(o[821]) );
  AND U3958 ( .A(p_input[20821]), .B(p_input[10821]), .Z(n1979) );
  AND U3959 ( .A(n1980), .B(p_input[8219]), .Z(o[8219]) );
  AND U3960 ( .A(p_input[28219]), .B(p_input[18219]), .Z(n1980) );
  AND U3961 ( .A(n1981), .B(p_input[8218]), .Z(o[8218]) );
  AND U3962 ( .A(p_input[28218]), .B(p_input[18218]), .Z(n1981) );
  AND U3963 ( .A(n1982), .B(p_input[8217]), .Z(o[8217]) );
  AND U3964 ( .A(p_input[28217]), .B(p_input[18217]), .Z(n1982) );
  AND U3965 ( .A(n1983), .B(p_input[8216]), .Z(o[8216]) );
  AND U3966 ( .A(p_input[28216]), .B(p_input[18216]), .Z(n1983) );
  AND U3967 ( .A(n1984), .B(p_input[8215]), .Z(o[8215]) );
  AND U3968 ( .A(p_input[28215]), .B(p_input[18215]), .Z(n1984) );
  AND U3969 ( .A(n1985), .B(p_input[8214]), .Z(o[8214]) );
  AND U3970 ( .A(p_input[28214]), .B(p_input[18214]), .Z(n1985) );
  AND U3971 ( .A(n1986), .B(p_input[8213]), .Z(o[8213]) );
  AND U3972 ( .A(p_input[28213]), .B(p_input[18213]), .Z(n1986) );
  AND U3973 ( .A(n1987), .B(p_input[8212]), .Z(o[8212]) );
  AND U3974 ( .A(p_input[28212]), .B(p_input[18212]), .Z(n1987) );
  AND U3975 ( .A(n1988), .B(p_input[8211]), .Z(o[8211]) );
  AND U3976 ( .A(p_input[28211]), .B(p_input[18211]), .Z(n1988) );
  AND U3977 ( .A(n1989), .B(p_input[8210]), .Z(o[8210]) );
  AND U3978 ( .A(p_input[28210]), .B(p_input[18210]), .Z(n1989) );
  AND U3979 ( .A(n1990), .B(p_input[820]), .Z(o[820]) );
  AND U3980 ( .A(p_input[20820]), .B(p_input[10820]), .Z(n1990) );
  AND U3981 ( .A(n1991), .B(p_input[8209]), .Z(o[8209]) );
  AND U3982 ( .A(p_input[28209]), .B(p_input[18209]), .Z(n1991) );
  AND U3983 ( .A(n1992), .B(p_input[8208]), .Z(o[8208]) );
  AND U3984 ( .A(p_input[28208]), .B(p_input[18208]), .Z(n1992) );
  AND U3985 ( .A(n1993), .B(p_input[8207]), .Z(o[8207]) );
  AND U3986 ( .A(p_input[28207]), .B(p_input[18207]), .Z(n1993) );
  AND U3987 ( .A(n1994), .B(p_input[8206]), .Z(o[8206]) );
  AND U3988 ( .A(p_input[28206]), .B(p_input[18206]), .Z(n1994) );
  AND U3989 ( .A(n1995), .B(p_input[8205]), .Z(o[8205]) );
  AND U3990 ( .A(p_input[28205]), .B(p_input[18205]), .Z(n1995) );
  AND U3991 ( .A(n1996), .B(p_input[8204]), .Z(o[8204]) );
  AND U3992 ( .A(p_input[28204]), .B(p_input[18204]), .Z(n1996) );
  AND U3993 ( .A(n1997), .B(p_input[8203]), .Z(o[8203]) );
  AND U3994 ( .A(p_input[28203]), .B(p_input[18203]), .Z(n1997) );
  AND U3995 ( .A(n1998), .B(p_input[8202]), .Z(o[8202]) );
  AND U3996 ( .A(p_input[28202]), .B(p_input[18202]), .Z(n1998) );
  AND U3997 ( .A(n1999), .B(p_input[8201]), .Z(o[8201]) );
  AND U3998 ( .A(p_input[28201]), .B(p_input[18201]), .Z(n1999) );
  AND U3999 ( .A(n2000), .B(p_input[8200]), .Z(o[8200]) );
  AND U4000 ( .A(p_input[28200]), .B(p_input[18200]), .Z(n2000) );
  AND U4001 ( .A(n2001), .B(p_input[81]), .Z(o[81]) );
  AND U4002 ( .A(p_input[20081]), .B(p_input[10081]), .Z(n2001) );
  AND U4003 ( .A(n2002), .B(p_input[819]), .Z(o[819]) );
  AND U4004 ( .A(p_input[20819]), .B(p_input[10819]), .Z(n2002) );
  AND U4005 ( .A(n2003), .B(p_input[8199]), .Z(o[8199]) );
  AND U4006 ( .A(p_input[28199]), .B(p_input[18199]), .Z(n2003) );
  AND U4007 ( .A(n2004), .B(p_input[8198]), .Z(o[8198]) );
  AND U4008 ( .A(p_input[28198]), .B(p_input[18198]), .Z(n2004) );
  AND U4009 ( .A(n2005), .B(p_input[8197]), .Z(o[8197]) );
  AND U4010 ( .A(p_input[28197]), .B(p_input[18197]), .Z(n2005) );
  AND U4011 ( .A(n2006), .B(p_input[8196]), .Z(o[8196]) );
  AND U4012 ( .A(p_input[28196]), .B(p_input[18196]), .Z(n2006) );
  AND U4013 ( .A(n2007), .B(p_input[8195]), .Z(o[8195]) );
  AND U4014 ( .A(p_input[28195]), .B(p_input[18195]), .Z(n2007) );
  AND U4015 ( .A(n2008), .B(p_input[8194]), .Z(o[8194]) );
  AND U4016 ( .A(p_input[28194]), .B(p_input[18194]), .Z(n2008) );
  AND U4017 ( .A(n2009), .B(p_input[8193]), .Z(o[8193]) );
  AND U4018 ( .A(p_input[28193]), .B(p_input[18193]), .Z(n2009) );
  AND U4019 ( .A(n2010), .B(p_input[8192]), .Z(o[8192]) );
  AND U4020 ( .A(p_input[28192]), .B(p_input[18192]), .Z(n2010) );
  AND U4021 ( .A(n2011), .B(p_input[8191]), .Z(o[8191]) );
  AND U4022 ( .A(p_input[28191]), .B(p_input[18191]), .Z(n2011) );
  AND U4023 ( .A(n2012), .B(p_input[8190]), .Z(o[8190]) );
  AND U4024 ( .A(p_input[28190]), .B(p_input[18190]), .Z(n2012) );
  AND U4025 ( .A(n2013), .B(p_input[818]), .Z(o[818]) );
  AND U4026 ( .A(p_input[20818]), .B(p_input[10818]), .Z(n2013) );
  AND U4027 ( .A(n2014), .B(p_input[8189]), .Z(o[8189]) );
  AND U4028 ( .A(p_input[28189]), .B(p_input[18189]), .Z(n2014) );
  AND U4029 ( .A(n2015), .B(p_input[8188]), .Z(o[8188]) );
  AND U4030 ( .A(p_input[28188]), .B(p_input[18188]), .Z(n2015) );
  AND U4031 ( .A(n2016), .B(p_input[8187]), .Z(o[8187]) );
  AND U4032 ( .A(p_input[28187]), .B(p_input[18187]), .Z(n2016) );
  AND U4033 ( .A(n2017), .B(p_input[8186]), .Z(o[8186]) );
  AND U4034 ( .A(p_input[28186]), .B(p_input[18186]), .Z(n2017) );
  AND U4035 ( .A(n2018), .B(p_input[8185]), .Z(o[8185]) );
  AND U4036 ( .A(p_input[28185]), .B(p_input[18185]), .Z(n2018) );
  AND U4037 ( .A(n2019), .B(p_input[8184]), .Z(o[8184]) );
  AND U4038 ( .A(p_input[28184]), .B(p_input[18184]), .Z(n2019) );
  AND U4039 ( .A(n2020), .B(p_input[8183]), .Z(o[8183]) );
  AND U4040 ( .A(p_input[28183]), .B(p_input[18183]), .Z(n2020) );
  AND U4041 ( .A(n2021), .B(p_input[8182]), .Z(o[8182]) );
  AND U4042 ( .A(p_input[28182]), .B(p_input[18182]), .Z(n2021) );
  AND U4043 ( .A(n2022), .B(p_input[8181]), .Z(o[8181]) );
  AND U4044 ( .A(p_input[28181]), .B(p_input[18181]), .Z(n2022) );
  AND U4045 ( .A(n2023), .B(p_input[8180]), .Z(o[8180]) );
  AND U4046 ( .A(p_input[28180]), .B(p_input[18180]), .Z(n2023) );
  AND U4047 ( .A(n2024), .B(p_input[817]), .Z(o[817]) );
  AND U4048 ( .A(p_input[20817]), .B(p_input[10817]), .Z(n2024) );
  AND U4049 ( .A(n2025), .B(p_input[8179]), .Z(o[8179]) );
  AND U4050 ( .A(p_input[28179]), .B(p_input[18179]), .Z(n2025) );
  AND U4051 ( .A(n2026), .B(p_input[8178]), .Z(o[8178]) );
  AND U4052 ( .A(p_input[28178]), .B(p_input[18178]), .Z(n2026) );
  AND U4053 ( .A(n2027), .B(p_input[8177]), .Z(o[8177]) );
  AND U4054 ( .A(p_input[28177]), .B(p_input[18177]), .Z(n2027) );
  AND U4055 ( .A(n2028), .B(p_input[8176]), .Z(o[8176]) );
  AND U4056 ( .A(p_input[28176]), .B(p_input[18176]), .Z(n2028) );
  AND U4057 ( .A(n2029), .B(p_input[8175]), .Z(o[8175]) );
  AND U4058 ( .A(p_input[28175]), .B(p_input[18175]), .Z(n2029) );
  AND U4059 ( .A(n2030), .B(p_input[8174]), .Z(o[8174]) );
  AND U4060 ( .A(p_input[28174]), .B(p_input[18174]), .Z(n2030) );
  AND U4061 ( .A(n2031), .B(p_input[8173]), .Z(o[8173]) );
  AND U4062 ( .A(p_input[28173]), .B(p_input[18173]), .Z(n2031) );
  AND U4063 ( .A(n2032), .B(p_input[8172]), .Z(o[8172]) );
  AND U4064 ( .A(p_input[28172]), .B(p_input[18172]), .Z(n2032) );
  AND U4065 ( .A(n2033), .B(p_input[8171]), .Z(o[8171]) );
  AND U4066 ( .A(p_input[28171]), .B(p_input[18171]), .Z(n2033) );
  AND U4067 ( .A(n2034), .B(p_input[8170]), .Z(o[8170]) );
  AND U4068 ( .A(p_input[28170]), .B(p_input[18170]), .Z(n2034) );
  AND U4069 ( .A(n2035), .B(p_input[816]), .Z(o[816]) );
  AND U4070 ( .A(p_input[20816]), .B(p_input[10816]), .Z(n2035) );
  AND U4071 ( .A(n2036), .B(p_input[8169]), .Z(o[8169]) );
  AND U4072 ( .A(p_input[28169]), .B(p_input[18169]), .Z(n2036) );
  AND U4073 ( .A(n2037), .B(p_input[8168]), .Z(o[8168]) );
  AND U4074 ( .A(p_input[28168]), .B(p_input[18168]), .Z(n2037) );
  AND U4075 ( .A(n2038), .B(p_input[8167]), .Z(o[8167]) );
  AND U4076 ( .A(p_input[28167]), .B(p_input[18167]), .Z(n2038) );
  AND U4077 ( .A(n2039), .B(p_input[8166]), .Z(o[8166]) );
  AND U4078 ( .A(p_input[28166]), .B(p_input[18166]), .Z(n2039) );
  AND U4079 ( .A(n2040), .B(p_input[8165]), .Z(o[8165]) );
  AND U4080 ( .A(p_input[28165]), .B(p_input[18165]), .Z(n2040) );
  AND U4081 ( .A(n2041), .B(p_input[8164]), .Z(o[8164]) );
  AND U4082 ( .A(p_input[28164]), .B(p_input[18164]), .Z(n2041) );
  AND U4083 ( .A(n2042), .B(p_input[8163]), .Z(o[8163]) );
  AND U4084 ( .A(p_input[28163]), .B(p_input[18163]), .Z(n2042) );
  AND U4085 ( .A(n2043), .B(p_input[8162]), .Z(o[8162]) );
  AND U4086 ( .A(p_input[28162]), .B(p_input[18162]), .Z(n2043) );
  AND U4087 ( .A(n2044), .B(p_input[8161]), .Z(o[8161]) );
  AND U4088 ( .A(p_input[28161]), .B(p_input[18161]), .Z(n2044) );
  AND U4089 ( .A(n2045), .B(p_input[8160]), .Z(o[8160]) );
  AND U4090 ( .A(p_input[28160]), .B(p_input[18160]), .Z(n2045) );
  AND U4091 ( .A(n2046), .B(p_input[815]), .Z(o[815]) );
  AND U4092 ( .A(p_input[20815]), .B(p_input[10815]), .Z(n2046) );
  AND U4093 ( .A(n2047), .B(p_input[8159]), .Z(o[8159]) );
  AND U4094 ( .A(p_input[28159]), .B(p_input[18159]), .Z(n2047) );
  AND U4095 ( .A(n2048), .B(p_input[8158]), .Z(o[8158]) );
  AND U4096 ( .A(p_input[28158]), .B(p_input[18158]), .Z(n2048) );
  AND U4097 ( .A(n2049), .B(p_input[8157]), .Z(o[8157]) );
  AND U4098 ( .A(p_input[28157]), .B(p_input[18157]), .Z(n2049) );
  AND U4099 ( .A(n2050), .B(p_input[8156]), .Z(o[8156]) );
  AND U4100 ( .A(p_input[28156]), .B(p_input[18156]), .Z(n2050) );
  AND U4101 ( .A(n2051), .B(p_input[8155]), .Z(o[8155]) );
  AND U4102 ( .A(p_input[28155]), .B(p_input[18155]), .Z(n2051) );
  AND U4103 ( .A(n2052), .B(p_input[8154]), .Z(o[8154]) );
  AND U4104 ( .A(p_input[28154]), .B(p_input[18154]), .Z(n2052) );
  AND U4105 ( .A(n2053), .B(p_input[8153]), .Z(o[8153]) );
  AND U4106 ( .A(p_input[28153]), .B(p_input[18153]), .Z(n2053) );
  AND U4107 ( .A(n2054), .B(p_input[8152]), .Z(o[8152]) );
  AND U4108 ( .A(p_input[28152]), .B(p_input[18152]), .Z(n2054) );
  AND U4109 ( .A(n2055), .B(p_input[8151]), .Z(o[8151]) );
  AND U4110 ( .A(p_input[28151]), .B(p_input[18151]), .Z(n2055) );
  AND U4111 ( .A(n2056), .B(p_input[8150]), .Z(o[8150]) );
  AND U4112 ( .A(p_input[28150]), .B(p_input[18150]), .Z(n2056) );
  AND U4113 ( .A(n2057), .B(p_input[814]), .Z(o[814]) );
  AND U4114 ( .A(p_input[20814]), .B(p_input[10814]), .Z(n2057) );
  AND U4115 ( .A(n2058), .B(p_input[8149]), .Z(o[8149]) );
  AND U4116 ( .A(p_input[28149]), .B(p_input[18149]), .Z(n2058) );
  AND U4117 ( .A(n2059), .B(p_input[8148]), .Z(o[8148]) );
  AND U4118 ( .A(p_input[28148]), .B(p_input[18148]), .Z(n2059) );
  AND U4119 ( .A(n2060), .B(p_input[8147]), .Z(o[8147]) );
  AND U4120 ( .A(p_input[28147]), .B(p_input[18147]), .Z(n2060) );
  AND U4121 ( .A(n2061), .B(p_input[8146]), .Z(o[8146]) );
  AND U4122 ( .A(p_input[28146]), .B(p_input[18146]), .Z(n2061) );
  AND U4123 ( .A(n2062), .B(p_input[8145]), .Z(o[8145]) );
  AND U4124 ( .A(p_input[28145]), .B(p_input[18145]), .Z(n2062) );
  AND U4125 ( .A(n2063), .B(p_input[8144]), .Z(o[8144]) );
  AND U4126 ( .A(p_input[28144]), .B(p_input[18144]), .Z(n2063) );
  AND U4127 ( .A(n2064), .B(p_input[8143]), .Z(o[8143]) );
  AND U4128 ( .A(p_input[28143]), .B(p_input[18143]), .Z(n2064) );
  AND U4129 ( .A(n2065), .B(p_input[8142]), .Z(o[8142]) );
  AND U4130 ( .A(p_input[28142]), .B(p_input[18142]), .Z(n2065) );
  AND U4131 ( .A(n2066), .B(p_input[8141]), .Z(o[8141]) );
  AND U4132 ( .A(p_input[28141]), .B(p_input[18141]), .Z(n2066) );
  AND U4133 ( .A(n2067), .B(p_input[8140]), .Z(o[8140]) );
  AND U4134 ( .A(p_input[28140]), .B(p_input[18140]), .Z(n2067) );
  AND U4135 ( .A(n2068), .B(p_input[813]), .Z(o[813]) );
  AND U4136 ( .A(p_input[20813]), .B(p_input[10813]), .Z(n2068) );
  AND U4137 ( .A(n2069), .B(p_input[8139]), .Z(o[8139]) );
  AND U4138 ( .A(p_input[28139]), .B(p_input[18139]), .Z(n2069) );
  AND U4139 ( .A(n2070), .B(p_input[8138]), .Z(o[8138]) );
  AND U4140 ( .A(p_input[28138]), .B(p_input[18138]), .Z(n2070) );
  AND U4141 ( .A(n2071), .B(p_input[8137]), .Z(o[8137]) );
  AND U4142 ( .A(p_input[28137]), .B(p_input[18137]), .Z(n2071) );
  AND U4143 ( .A(n2072), .B(p_input[8136]), .Z(o[8136]) );
  AND U4144 ( .A(p_input[28136]), .B(p_input[18136]), .Z(n2072) );
  AND U4145 ( .A(n2073), .B(p_input[8135]), .Z(o[8135]) );
  AND U4146 ( .A(p_input[28135]), .B(p_input[18135]), .Z(n2073) );
  AND U4147 ( .A(n2074), .B(p_input[8134]), .Z(o[8134]) );
  AND U4148 ( .A(p_input[28134]), .B(p_input[18134]), .Z(n2074) );
  AND U4149 ( .A(n2075), .B(p_input[8133]), .Z(o[8133]) );
  AND U4150 ( .A(p_input[28133]), .B(p_input[18133]), .Z(n2075) );
  AND U4151 ( .A(n2076), .B(p_input[8132]), .Z(o[8132]) );
  AND U4152 ( .A(p_input[28132]), .B(p_input[18132]), .Z(n2076) );
  AND U4153 ( .A(n2077), .B(p_input[8131]), .Z(o[8131]) );
  AND U4154 ( .A(p_input[28131]), .B(p_input[18131]), .Z(n2077) );
  AND U4155 ( .A(n2078), .B(p_input[8130]), .Z(o[8130]) );
  AND U4156 ( .A(p_input[28130]), .B(p_input[18130]), .Z(n2078) );
  AND U4157 ( .A(n2079), .B(p_input[812]), .Z(o[812]) );
  AND U4158 ( .A(p_input[20812]), .B(p_input[10812]), .Z(n2079) );
  AND U4159 ( .A(n2080), .B(p_input[8129]), .Z(o[8129]) );
  AND U4160 ( .A(p_input[28129]), .B(p_input[18129]), .Z(n2080) );
  AND U4161 ( .A(n2081), .B(p_input[8128]), .Z(o[8128]) );
  AND U4162 ( .A(p_input[28128]), .B(p_input[18128]), .Z(n2081) );
  AND U4163 ( .A(n2082), .B(p_input[8127]), .Z(o[8127]) );
  AND U4164 ( .A(p_input[28127]), .B(p_input[18127]), .Z(n2082) );
  AND U4165 ( .A(n2083), .B(p_input[8126]), .Z(o[8126]) );
  AND U4166 ( .A(p_input[28126]), .B(p_input[18126]), .Z(n2083) );
  AND U4167 ( .A(n2084), .B(p_input[8125]), .Z(o[8125]) );
  AND U4168 ( .A(p_input[28125]), .B(p_input[18125]), .Z(n2084) );
  AND U4169 ( .A(n2085), .B(p_input[8124]), .Z(o[8124]) );
  AND U4170 ( .A(p_input[28124]), .B(p_input[18124]), .Z(n2085) );
  AND U4171 ( .A(n2086), .B(p_input[8123]), .Z(o[8123]) );
  AND U4172 ( .A(p_input[28123]), .B(p_input[18123]), .Z(n2086) );
  AND U4173 ( .A(n2087), .B(p_input[8122]), .Z(o[8122]) );
  AND U4174 ( .A(p_input[28122]), .B(p_input[18122]), .Z(n2087) );
  AND U4175 ( .A(n2088), .B(p_input[8121]), .Z(o[8121]) );
  AND U4176 ( .A(p_input[28121]), .B(p_input[18121]), .Z(n2088) );
  AND U4177 ( .A(n2089), .B(p_input[8120]), .Z(o[8120]) );
  AND U4178 ( .A(p_input[28120]), .B(p_input[18120]), .Z(n2089) );
  AND U4179 ( .A(n2090), .B(p_input[811]), .Z(o[811]) );
  AND U4180 ( .A(p_input[20811]), .B(p_input[10811]), .Z(n2090) );
  AND U4181 ( .A(n2091), .B(p_input[8119]), .Z(o[8119]) );
  AND U4182 ( .A(p_input[28119]), .B(p_input[18119]), .Z(n2091) );
  AND U4183 ( .A(n2092), .B(p_input[8118]), .Z(o[8118]) );
  AND U4184 ( .A(p_input[28118]), .B(p_input[18118]), .Z(n2092) );
  AND U4185 ( .A(n2093), .B(p_input[8117]), .Z(o[8117]) );
  AND U4186 ( .A(p_input[28117]), .B(p_input[18117]), .Z(n2093) );
  AND U4187 ( .A(n2094), .B(p_input[8116]), .Z(o[8116]) );
  AND U4188 ( .A(p_input[28116]), .B(p_input[18116]), .Z(n2094) );
  AND U4189 ( .A(n2095), .B(p_input[8115]), .Z(o[8115]) );
  AND U4190 ( .A(p_input[28115]), .B(p_input[18115]), .Z(n2095) );
  AND U4191 ( .A(n2096), .B(p_input[8114]), .Z(o[8114]) );
  AND U4192 ( .A(p_input[28114]), .B(p_input[18114]), .Z(n2096) );
  AND U4193 ( .A(n2097), .B(p_input[8113]), .Z(o[8113]) );
  AND U4194 ( .A(p_input[28113]), .B(p_input[18113]), .Z(n2097) );
  AND U4195 ( .A(n2098), .B(p_input[8112]), .Z(o[8112]) );
  AND U4196 ( .A(p_input[28112]), .B(p_input[18112]), .Z(n2098) );
  AND U4197 ( .A(n2099), .B(p_input[8111]), .Z(o[8111]) );
  AND U4198 ( .A(p_input[28111]), .B(p_input[18111]), .Z(n2099) );
  AND U4199 ( .A(n2100), .B(p_input[8110]), .Z(o[8110]) );
  AND U4200 ( .A(p_input[28110]), .B(p_input[18110]), .Z(n2100) );
  AND U4201 ( .A(n2101), .B(p_input[810]), .Z(o[810]) );
  AND U4202 ( .A(p_input[20810]), .B(p_input[10810]), .Z(n2101) );
  AND U4203 ( .A(n2102), .B(p_input[8109]), .Z(o[8109]) );
  AND U4204 ( .A(p_input[28109]), .B(p_input[18109]), .Z(n2102) );
  AND U4205 ( .A(n2103), .B(p_input[8108]), .Z(o[8108]) );
  AND U4206 ( .A(p_input[28108]), .B(p_input[18108]), .Z(n2103) );
  AND U4207 ( .A(n2104), .B(p_input[8107]), .Z(o[8107]) );
  AND U4208 ( .A(p_input[28107]), .B(p_input[18107]), .Z(n2104) );
  AND U4209 ( .A(n2105), .B(p_input[8106]), .Z(o[8106]) );
  AND U4210 ( .A(p_input[28106]), .B(p_input[18106]), .Z(n2105) );
  AND U4211 ( .A(n2106), .B(p_input[8105]), .Z(o[8105]) );
  AND U4212 ( .A(p_input[28105]), .B(p_input[18105]), .Z(n2106) );
  AND U4213 ( .A(n2107), .B(p_input[8104]), .Z(o[8104]) );
  AND U4214 ( .A(p_input[28104]), .B(p_input[18104]), .Z(n2107) );
  AND U4215 ( .A(n2108), .B(p_input[8103]), .Z(o[8103]) );
  AND U4216 ( .A(p_input[28103]), .B(p_input[18103]), .Z(n2108) );
  AND U4217 ( .A(n2109), .B(p_input[8102]), .Z(o[8102]) );
  AND U4218 ( .A(p_input[28102]), .B(p_input[18102]), .Z(n2109) );
  AND U4219 ( .A(n2110), .B(p_input[8101]), .Z(o[8101]) );
  AND U4220 ( .A(p_input[28101]), .B(p_input[18101]), .Z(n2110) );
  AND U4221 ( .A(n2111), .B(p_input[8100]), .Z(o[8100]) );
  AND U4222 ( .A(p_input[28100]), .B(p_input[18100]), .Z(n2111) );
  AND U4223 ( .A(n2112), .B(p_input[80]), .Z(o[80]) );
  AND U4224 ( .A(p_input[20080]), .B(p_input[10080]), .Z(n2112) );
  AND U4225 ( .A(n2113), .B(p_input[809]), .Z(o[809]) );
  AND U4226 ( .A(p_input[20809]), .B(p_input[10809]), .Z(n2113) );
  AND U4227 ( .A(n2114), .B(p_input[8099]), .Z(o[8099]) );
  AND U4228 ( .A(p_input[28099]), .B(p_input[18099]), .Z(n2114) );
  AND U4229 ( .A(n2115), .B(p_input[8098]), .Z(o[8098]) );
  AND U4230 ( .A(p_input[28098]), .B(p_input[18098]), .Z(n2115) );
  AND U4231 ( .A(n2116), .B(p_input[8097]), .Z(o[8097]) );
  AND U4232 ( .A(p_input[28097]), .B(p_input[18097]), .Z(n2116) );
  AND U4233 ( .A(n2117), .B(p_input[8096]), .Z(o[8096]) );
  AND U4234 ( .A(p_input[28096]), .B(p_input[18096]), .Z(n2117) );
  AND U4235 ( .A(n2118), .B(p_input[8095]), .Z(o[8095]) );
  AND U4236 ( .A(p_input[28095]), .B(p_input[18095]), .Z(n2118) );
  AND U4237 ( .A(n2119), .B(p_input[8094]), .Z(o[8094]) );
  AND U4238 ( .A(p_input[28094]), .B(p_input[18094]), .Z(n2119) );
  AND U4239 ( .A(n2120), .B(p_input[8093]), .Z(o[8093]) );
  AND U4240 ( .A(p_input[28093]), .B(p_input[18093]), .Z(n2120) );
  AND U4241 ( .A(n2121), .B(p_input[8092]), .Z(o[8092]) );
  AND U4242 ( .A(p_input[28092]), .B(p_input[18092]), .Z(n2121) );
  AND U4243 ( .A(n2122), .B(p_input[8091]), .Z(o[8091]) );
  AND U4244 ( .A(p_input[28091]), .B(p_input[18091]), .Z(n2122) );
  AND U4245 ( .A(n2123), .B(p_input[8090]), .Z(o[8090]) );
  AND U4246 ( .A(p_input[28090]), .B(p_input[18090]), .Z(n2123) );
  AND U4247 ( .A(n2124), .B(p_input[808]), .Z(o[808]) );
  AND U4248 ( .A(p_input[20808]), .B(p_input[10808]), .Z(n2124) );
  AND U4249 ( .A(n2125), .B(p_input[8089]), .Z(o[8089]) );
  AND U4250 ( .A(p_input[28089]), .B(p_input[18089]), .Z(n2125) );
  AND U4251 ( .A(n2126), .B(p_input[8088]), .Z(o[8088]) );
  AND U4252 ( .A(p_input[28088]), .B(p_input[18088]), .Z(n2126) );
  AND U4253 ( .A(n2127), .B(p_input[8087]), .Z(o[8087]) );
  AND U4254 ( .A(p_input[28087]), .B(p_input[18087]), .Z(n2127) );
  AND U4255 ( .A(n2128), .B(p_input[8086]), .Z(o[8086]) );
  AND U4256 ( .A(p_input[28086]), .B(p_input[18086]), .Z(n2128) );
  AND U4257 ( .A(n2129), .B(p_input[8085]), .Z(o[8085]) );
  AND U4258 ( .A(p_input[28085]), .B(p_input[18085]), .Z(n2129) );
  AND U4259 ( .A(n2130), .B(p_input[8084]), .Z(o[8084]) );
  AND U4260 ( .A(p_input[28084]), .B(p_input[18084]), .Z(n2130) );
  AND U4261 ( .A(n2131), .B(p_input[8083]), .Z(o[8083]) );
  AND U4262 ( .A(p_input[28083]), .B(p_input[18083]), .Z(n2131) );
  AND U4263 ( .A(n2132), .B(p_input[8082]), .Z(o[8082]) );
  AND U4264 ( .A(p_input[28082]), .B(p_input[18082]), .Z(n2132) );
  AND U4265 ( .A(n2133), .B(p_input[8081]), .Z(o[8081]) );
  AND U4266 ( .A(p_input[28081]), .B(p_input[18081]), .Z(n2133) );
  AND U4267 ( .A(n2134), .B(p_input[8080]), .Z(o[8080]) );
  AND U4268 ( .A(p_input[28080]), .B(p_input[18080]), .Z(n2134) );
  AND U4269 ( .A(n2135), .B(p_input[807]), .Z(o[807]) );
  AND U4270 ( .A(p_input[20807]), .B(p_input[10807]), .Z(n2135) );
  AND U4271 ( .A(n2136), .B(p_input[8079]), .Z(o[8079]) );
  AND U4272 ( .A(p_input[28079]), .B(p_input[18079]), .Z(n2136) );
  AND U4273 ( .A(n2137), .B(p_input[8078]), .Z(o[8078]) );
  AND U4274 ( .A(p_input[28078]), .B(p_input[18078]), .Z(n2137) );
  AND U4275 ( .A(n2138), .B(p_input[8077]), .Z(o[8077]) );
  AND U4276 ( .A(p_input[28077]), .B(p_input[18077]), .Z(n2138) );
  AND U4277 ( .A(n2139), .B(p_input[8076]), .Z(o[8076]) );
  AND U4278 ( .A(p_input[28076]), .B(p_input[18076]), .Z(n2139) );
  AND U4279 ( .A(n2140), .B(p_input[8075]), .Z(o[8075]) );
  AND U4280 ( .A(p_input[28075]), .B(p_input[18075]), .Z(n2140) );
  AND U4281 ( .A(n2141), .B(p_input[8074]), .Z(o[8074]) );
  AND U4282 ( .A(p_input[28074]), .B(p_input[18074]), .Z(n2141) );
  AND U4283 ( .A(n2142), .B(p_input[8073]), .Z(o[8073]) );
  AND U4284 ( .A(p_input[28073]), .B(p_input[18073]), .Z(n2142) );
  AND U4285 ( .A(n2143), .B(p_input[8072]), .Z(o[8072]) );
  AND U4286 ( .A(p_input[28072]), .B(p_input[18072]), .Z(n2143) );
  AND U4287 ( .A(n2144), .B(p_input[8071]), .Z(o[8071]) );
  AND U4288 ( .A(p_input[28071]), .B(p_input[18071]), .Z(n2144) );
  AND U4289 ( .A(n2145), .B(p_input[8070]), .Z(o[8070]) );
  AND U4290 ( .A(p_input[28070]), .B(p_input[18070]), .Z(n2145) );
  AND U4291 ( .A(n2146), .B(p_input[806]), .Z(o[806]) );
  AND U4292 ( .A(p_input[20806]), .B(p_input[10806]), .Z(n2146) );
  AND U4293 ( .A(n2147), .B(p_input[8069]), .Z(o[8069]) );
  AND U4294 ( .A(p_input[28069]), .B(p_input[18069]), .Z(n2147) );
  AND U4295 ( .A(n2148), .B(p_input[8068]), .Z(o[8068]) );
  AND U4296 ( .A(p_input[28068]), .B(p_input[18068]), .Z(n2148) );
  AND U4297 ( .A(n2149), .B(p_input[8067]), .Z(o[8067]) );
  AND U4298 ( .A(p_input[28067]), .B(p_input[18067]), .Z(n2149) );
  AND U4299 ( .A(n2150), .B(p_input[8066]), .Z(o[8066]) );
  AND U4300 ( .A(p_input[28066]), .B(p_input[18066]), .Z(n2150) );
  AND U4301 ( .A(n2151), .B(p_input[8065]), .Z(o[8065]) );
  AND U4302 ( .A(p_input[28065]), .B(p_input[18065]), .Z(n2151) );
  AND U4303 ( .A(n2152), .B(p_input[8064]), .Z(o[8064]) );
  AND U4304 ( .A(p_input[28064]), .B(p_input[18064]), .Z(n2152) );
  AND U4305 ( .A(n2153), .B(p_input[8063]), .Z(o[8063]) );
  AND U4306 ( .A(p_input[28063]), .B(p_input[18063]), .Z(n2153) );
  AND U4307 ( .A(n2154), .B(p_input[8062]), .Z(o[8062]) );
  AND U4308 ( .A(p_input[28062]), .B(p_input[18062]), .Z(n2154) );
  AND U4309 ( .A(n2155), .B(p_input[8061]), .Z(o[8061]) );
  AND U4310 ( .A(p_input[28061]), .B(p_input[18061]), .Z(n2155) );
  AND U4311 ( .A(n2156), .B(p_input[8060]), .Z(o[8060]) );
  AND U4312 ( .A(p_input[28060]), .B(p_input[18060]), .Z(n2156) );
  AND U4313 ( .A(n2157), .B(p_input[805]), .Z(o[805]) );
  AND U4314 ( .A(p_input[20805]), .B(p_input[10805]), .Z(n2157) );
  AND U4315 ( .A(n2158), .B(p_input[8059]), .Z(o[8059]) );
  AND U4316 ( .A(p_input[28059]), .B(p_input[18059]), .Z(n2158) );
  AND U4317 ( .A(n2159), .B(p_input[8058]), .Z(o[8058]) );
  AND U4318 ( .A(p_input[28058]), .B(p_input[18058]), .Z(n2159) );
  AND U4319 ( .A(n2160), .B(p_input[8057]), .Z(o[8057]) );
  AND U4320 ( .A(p_input[28057]), .B(p_input[18057]), .Z(n2160) );
  AND U4321 ( .A(n2161), .B(p_input[8056]), .Z(o[8056]) );
  AND U4322 ( .A(p_input[28056]), .B(p_input[18056]), .Z(n2161) );
  AND U4323 ( .A(n2162), .B(p_input[8055]), .Z(o[8055]) );
  AND U4324 ( .A(p_input[28055]), .B(p_input[18055]), .Z(n2162) );
  AND U4325 ( .A(n2163), .B(p_input[8054]), .Z(o[8054]) );
  AND U4326 ( .A(p_input[28054]), .B(p_input[18054]), .Z(n2163) );
  AND U4327 ( .A(n2164), .B(p_input[8053]), .Z(o[8053]) );
  AND U4328 ( .A(p_input[28053]), .B(p_input[18053]), .Z(n2164) );
  AND U4329 ( .A(n2165), .B(p_input[8052]), .Z(o[8052]) );
  AND U4330 ( .A(p_input[28052]), .B(p_input[18052]), .Z(n2165) );
  AND U4331 ( .A(n2166), .B(p_input[8051]), .Z(o[8051]) );
  AND U4332 ( .A(p_input[28051]), .B(p_input[18051]), .Z(n2166) );
  AND U4333 ( .A(n2167), .B(p_input[8050]), .Z(o[8050]) );
  AND U4334 ( .A(p_input[28050]), .B(p_input[18050]), .Z(n2167) );
  AND U4335 ( .A(n2168), .B(p_input[804]), .Z(o[804]) );
  AND U4336 ( .A(p_input[20804]), .B(p_input[10804]), .Z(n2168) );
  AND U4337 ( .A(n2169), .B(p_input[8049]), .Z(o[8049]) );
  AND U4338 ( .A(p_input[28049]), .B(p_input[18049]), .Z(n2169) );
  AND U4339 ( .A(n2170), .B(p_input[8048]), .Z(o[8048]) );
  AND U4340 ( .A(p_input[28048]), .B(p_input[18048]), .Z(n2170) );
  AND U4341 ( .A(n2171), .B(p_input[8047]), .Z(o[8047]) );
  AND U4342 ( .A(p_input[28047]), .B(p_input[18047]), .Z(n2171) );
  AND U4343 ( .A(n2172), .B(p_input[8046]), .Z(o[8046]) );
  AND U4344 ( .A(p_input[28046]), .B(p_input[18046]), .Z(n2172) );
  AND U4345 ( .A(n2173), .B(p_input[8045]), .Z(o[8045]) );
  AND U4346 ( .A(p_input[28045]), .B(p_input[18045]), .Z(n2173) );
  AND U4347 ( .A(n2174), .B(p_input[8044]), .Z(o[8044]) );
  AND U4348 ( .A(p_input[28044]), .B(p_input[18044]), .Z(n2174) );
  AND U4349 ( .A(n2175), .B(p_input[8043]), .Z(o[8043]) );
  AND U4350 ( .A(p_input[28043]), .B(p_input[18043]), .Z(n2175) );
  AND U4351 ( .A(n2176), .B(p_input[8042]), .Z(o[8042]) );
  AND U4352 ( .A(p_input[28042]), .B(p_input[18042]), .Z(n2176) );
  AND U4353 ( .A(n2177), .B(p_input[8041]), .Z(o[8041]) );
  AND U4354 ( .A(p_input[28041]), .B(p_input[18041]), .Z(n2177) );
  AND U4355 ( .A(n2178), .B(p_input[8040]), .Z(o[8040]) );
  AND U4356 ( .A(p_input[28040]), .B(p_input[18040]), .Z(n2178) );
  AND U4357 ( .A(n2179), .B(p_input[803]), .Z(o[803]) );
  AND U4358 ( .A(p_input[20803]), .B(p_input[10803]), .Z(n2179) );
  AND U4359 ( .A(n2180), .B(p_input[8039]), .Z(o[8039]) );
  AND U4360 ( .A(p_input[28039]), .B(p_input[18039]), .Z(n2180) );
  AND U4361 ( .A(n2181), .B(p_input[8038]), .Z(o[8038]) );
  AND U4362 ( .A(p_input[28038]), .B(p_input[18038]), .Z(n2181) );
  AND U4363 ( .A(n2182), .B(p_input[8037]), .Z(o[8037]) );
  AND U4364 ( .A(p_input[28037]), .B(p_input[18037]), .Z(n2182) );
  AND U4365 ( .A(n2183), .B(p_input[8036]), .Z(o[8036]) );
  AND U4366 ( .A(p_input[28036]), .B(p_input[18036]), .Z(n2183) );
  AND U4367 ( .A(n2184), .B(p_input[8035]), .Z(o[8035]) );
  AND U4368 ( .A(p_input[28035]), .B(p_input[18035]), .Z(n2184) );
  AND U4369 ( .A(n2185), .B(p_input[8034]), .Z(o[8034]) );
  AND U4370 ( .A(p_input[28034]), .B(p_input[18034]), .Z(n2185) );
  AND U4371 ( .A(n2186), .B(p_input[8033]), .Z(o[8033]) );
  AND U4372 ( .A(p_input[28033]), .B(p_input[18033]), .Z(n2186) );
  AND U4373 ( .A(n2187), .B(p_input[8032]), .Z(o[8032]) );
  AND U4374 ( .A(p_input[28032]), .B(p_input[18032]), .Z(n2187) );
  AND U4375 ( .A(n2188), .B(p_input[8031]), .Z(o[8031]) );
  AND U4376 ( .A(p_input[28031]), .B(p_input[18031]), .Z(n2188) );
  AND U4377 ( .A(n2189), .B(p_input[8030]), .Z(o[8030]) );
  AND U4378 ( .A(p_input[28030]), .B(p_input[18030]), .Z(n2189) );
  AND U4379 ( .A(n2190), .B(p_input[802]), .Z(o[802]) );
  AND U4380 ( .A(p_input[20802]), .B(p_input[10802]), .Z(n2190) );
  AND U4381 ( .A(n2191), .B(p_input[8029]), .Z(o[8029]) );
  AND U4382 ( .A(p_input[28029]), .B(p_input[18029]), .Z(n2191) );
  AND U4383 ( .A(n2192), .B(p_input[8028]), .Z(o[8028]) );
  AND U4384 ( .A(p_input[28028]), .B(p_input[18028]), .Z(n2192) );
  AND U4385 ( .A(n2193), .B(p_input[8027]), .Z(o[8027]) );
  AND U4386 ( .A(p_input[28027]), .B(p_input[18027]), .Z(n2193) );
  AND U4387 ( .A(n2194), .B(p_input[8026]), .Z(o[8026]) );
  AND U4388 ( .A(p_input[28026]), .B(p_input[18026]), .Z(n2194) );
  AND U4389 ( .A(n2195), .B(p_input[8025]), .Z(o[8025]) );
  AND U4390 ( .A(p_input[28025]), .B(p_input[18025]), .Z(n2195) );
  AND U4391 ( .A(n2196), .B(p_input[8024]), .Z(o[8024]) );
  AND U4392 ( .A(p_input[28024]), .B(p_input[18024]), .Z(n2196) );
  AND U4393 ( .A(n2197), .B(p_input[8023]), .Z(o[8023]) );
  AND U4394 ( .A(p_input[28023]), .B(p_input[18023]), .Z(n2197) );
  AND U4395 ( .A(n2198), .B(p_input[8022]), .Z(o[8022]) );
  AND U4396 ( .A(p_input[28022]), .B(p_input[18022]), .Z(n2198) );
  AND U4397 ( .A(n2199), .B(p_input[8021]), .Z(o[8021]) );
  AND U4398 ( .A(p_input[28021]), .B(p_input[18021]), .Z(n2199) );
  AND U4399 ( .A(n2200), .B(p_input[8020]), .Z(o[8020]) );
  AND U4400 ( .A(p_input[28020]), .B(p_input[18020]), .Z(n2200) );
  AND U4401 ( .A(n2201), .B(p_input[801]), .Z(o[801]) );
  AND U4402 ( .A(p_input[20801]), .B(p_input[10801]), .Z(n2201) );
  AND U4403 ( .A(n2202), .B(p_input[8019]), .Z(o[8019]) );
  AND U4404 ( .A(p_input[28019]), .B(p_input[18019]), .Z(n2202) );
  AND U4405 ( .A(n2203), .B(p_input[8018]), .Z(o[8018]) );
  AND U4406 ( .A(p_input[28018]), .B(p_input[18018]), .Z(n2203) );
  AND U4407 ( .A(n2204), .B(p_input[8017]), .Z(o[8017]) );
  AND U4408 ( .A(p_input[28017]), .B(p_input[18017]), .Z(n2204) );
  AND U4409 ( .A(n2205), .B(p_input[8016]), .Z(o[8016]) );
  AND U4410 ( .A(p_input[28016]), .B(p_input[18016]), .Z(n2205) );
  AND U4411 ( .A(n2206), .B(p_input[8015]), .Z(o[8015]) );
  AND U4412 ( .A(p_input[28015]), .B(p_input[18015]), .Z(n2206) );
  AND U4413 ( .A(n2207), .B(p_input[8014]), .Z(o[8014]) );
  AND U4414 ( .A(p_input[28014]), .B(p_input[18014]), .Z(n2207) );
  AND U4415 ( .A(n2208), .B(p_input[8013]), .Z(o[8013]) );
  AND U4416 ( .A(p_input[28013]), .B(p_input[18013]), .Z(n2208) );
  AND U4417 ( .A(n2209), .B(p_input[8012]), .Z(o[8012]) );
  AND U4418 ( .A(p_input[28012]), .B(p_input[18012]), .Z(n2209) );
  AND U4419 ( .A(n2210), .B(p_input[8011]), .Z(o[8011]) );
  AND U4420 ( .A(p_input[28011]), .B(p_input[18011]), .Z(n2210) );
  AND U4421 ( .A(n2211), .B(p_input[8010]), .Z(o[8010]) );
  AND U4422 ( .A(p_input[28010]), .B(p_input[18010]), .Z(n2211) );
  AND U4423 ( .A(n2212), .B(p_input[800]), .Z(o[800]) );
  AND U4424 ( .A(p_input[20800]), .B(p_input[10800]), .Z(n2212) );
  AND U4425 ( .A(n2213), .B(p_input[8009]), .Z(o[8009]) );
  AND U4426 ( .A(p_input[28009]), .B(p_input[18009]), .Z(n2213) );
  AND U4427 ( .A(n2214), .B(p_input[8008]), .Z(o[8008]) );
  AND U4428 ( .A(p_input[28008]), .B(p_input[18008]), .Z(n2214) );
  AND U4429 ( .A(n2215), .B(p_input[8007]), .Z(o[8007]) );
  AND U4430 ( .A(p_input[28007]), .B(p_input[18007]), .Z(n2215) );
  AND U4431 ( .A(n2216), .B(p_input[8006]), .Z(o[8006]) );
  AND U4432 ( .A(p_input[28006]), .B(p_input[18006]), .Z(n2216) );
  AND U4433 ( .A(n2217), .B(p_input[8005]), .Z(o[8005]) );
  AND U4434 ( .A(p_input[28005]), .B(p_input[18005]), .Z(n2217) );
  AND U4435 ( .A(n2218), .B(p_input[8004]), .Z(o[8004]) );
  AND U4436 ( .A(p_input[28004]), .B(p_input[18004]), .Z(n2218) );
  AND U4437 ( .A(n2219), .B(p_input[8003]), .Z(o[8003]) );
  AND U4438 ( .A(p_input[28003]), .B(p_input[18003]), .Z(n2219) );
  AND U4439 ( .A(n2220), .B(p_input[8002]), .Z(o[8002]) );
  AND U4440 ( .A(p_input[28002]), .B(p_input[18002]), .Z(n2220) );
  AND U4441 ( .A(n2221), .B(p_input[8001]), .Z(o[8001]) );
  AND U4442 ( .A(p_input[28001]), .B(p_input[18001]), .Z(n2221) );
  AND U4443 ( .A(n2222), .B(p_input[8000]), .Z(o[8000]) );
  AND U4444 ( .A(p_input[28000]), .B(p_input[18000]), .Z(n2222) );
  AND U4445 ( .A(n2223), .B(p_input[7]), .Z(o[7]) );
  AND U4446 ( .A(p_input[20007]), .B(p_input[10007]), .Z(n2223) );
  AND U4447 ( .A(n2224), .B(p_input[79]), .Z(o[79]) );
  AND U4448 ( .A(p_input[20079]), .B(p_input[10079]), .Z(n2224) );
  AND U4449 ( .A(n2225), .B(p_input[799]), .Z(o[799]) );
  AND U4450 ( .A(p_input[20799]), .B(p_input[10799]), .Z(n2225) );
  AND U4451 ( .A(n2226), .B(p_input[7999]), .Z(o[7999]) );
  AND U4452 ( .A(p_input[27999]), .B(p_input[17999]), .Z(n2226) );
  AND U4453 ( .A(n2227), .B(p_input[7998]), .Z(o[7998]) );
  AND U4454 ( .A(p_input[27998]), .B(p_input[17998]), .Z(n2227) );
  AND U4455 ( .A(n2228), .B(p_input[7997]), .Z(o[7997]) );
  AND U4456 ( .A(p_input[27997]), .B(p_input[17997]), .Z(n2228) );
  AND U4457 ( .A(n2229), .B(p_input[7996]), .Z(o[7996]) );
  AND U4458 ( .A(p_input[27996]), .B(p_input[17996]), .Z(n2229) );
  AND U4459 ( .A(n2230), .B(p_input[7995]), .Z(o[7995]) );
  AND U4460 ( .A(p_input[27995]), .B(p_input[17995]), .Z(n2230) );
  AND U4461 ( .A(n2231), .B(p_input[7994]), .Z(o[7994]) );
  AND U4462 ( .A(p_input[27994]), .B(p_input[17994]), .Z(n2231) );
  AND U4463 ( .A(n2232), .B(p_input[7993]), .Z(o[7993]) );
  AND U4464 ( .A(p_input[27993]), .B(p_input[17993]), .Z(n2232) );
  AND U4465 ( .A(n2233), .B(p_input[7992]), .Z(o[7992]) );
  AND U4466 ( .A(p_input[27992]), .B(p_input[17992]), .Z(n2233) );
  AND U4467 ( .A(n2234), .B(p_input[7991]), .Z(o[7991]) );
  AND U4468 ( .A(p_input[27991]), .B(p_input[17991]), .Z(n2234) );
  AND U4469 ( .A(n2235), .B(p_input[7990]), .Z(o[7990]) );
  AND U4470 ( .A(p_input[27990]), .B(p_input[17990]), .Z(n2235) );
  AND U4471 ( .A(n2236), .B(p_input[798]), .Z(o[798]) );
  AND U4472 ( .A(p_input[20798]), .B(p_input[10798]), .Z(n2236) );
  AND U4473 ( .A(n2237), .B(p_input[7989]), .Z(o[7989]) );
  AND U4474 ( .A(p_input[27989]), .B(p_input[17989]), .Z(n2237) );
  AND U4475 ( .A(n2238), .B(p_input[7988]), .Z(o[7988]) );
  AND U4476 ( .A(p_input[27988]), .B(p_input[17988]), .Z(n2238) );
  AND U4477 ( .A(n2239), .B(p_input[7987]), .Z(o[7987]) );
  AND U4478 ( .A(p_input[27987]), .B(p_input[17987]), .Z(n2239) );
  AND U4479 ( .A(n2240), .B(p_input[7986]), .Z(o[7986]) );
  AND U4480 ( .A(p_input[27986]), .B(p_input[17986]), .Z(n2240) );
  AND U4481 ( .A(n2241), .B(p_input[7985]), .Z(o[7985]) );
  AND U4482 ( .A(p_input[27985]), .B(p_input[17985]), .Z(n2241) );
  AND U4483 ( .A(n2242), .B(p_input[7984]), .Z(o[7984]) );
  AND U4484 ( .A(p_input[27984]), .B(p_input[17984]), .Z(n2242) );
  AND U4485 ( .A(n2243), .B(p_input[7983]), .Z(o[7983]) );
  AND U4486 ( .A(p_input[27983]), .B(p_input[17983]), .Z(n2243) );
  AND U4487 ( .A(n2244), .B(p_input[7982]), .Z(o[7982]) );
  AND U4488 ( .A(p_input[27982]), .B(p_input[17982]), .Z(n2244) );
  AND U4489 ( .A(n2245), .B(p_input[7981]), .Z(o[7981]) );
  AND U4490 ( .A(p_input[27981]), .B(p_input[17981]), .Z(n2245) );
  AND U4491 ( .A(n2246), .B(p_input[7980]), .Z(o[7980]) );
  AND U4492 ( .A(p_input[27980]), .B(p_input[17980]), .Z(n2246) );
  AND U4493 ( .A(n2247), .B(p_input[797]), .Z(o[797]) );
  AND U4494 ( .A(p_input[20797]), .B(p_input[10797]), .Z(n2247) );
  AND U4495 ( .A(n2248), .B(p_input[7979]), .Z(o[7979]) );
  AND U4496 ( .A(p_input[27979]), .B(p_input[17979]), .Z(n2248) );
  AND U4497 ( .A(n2249), .B(p_input[7978]), .Z(o[7978]) );
  AND U4498 ( .A(p_input[27978]), .B(p_input[17978]), .Z(n2249) );
  AND U4499 ( .A(n2250), .B(p_input[7977]), .Z(o[7977]) );
  AND U4500 ( .A(p_input[27977]), .B(p_input[17977]), .Z(n2250) );
  AND U4501 ( .A(n2251), .B(p_input[7976]), .Z(o[7976]) );
  AND U4502 ( .A(p_input[27976]), .B(p_input[17976]), .Z(n2251) );
  AND U4503 ( .A(n2252), .B(p_input[7975]), .Z(o[7975]) );
  AND U4504 ( .A(p_input[27975]), .B(p_input[17975]), .Z(n2252) );
  AND U4505 ( .A(n2253), .B(p_input[7974]), .Z(o[7974]) );
  AND U4506 ( .A(p_input[27974]), .B(p_input[17974]), .Z(n2253) );
  AND U4507 ( .A(n2254), .B(p_input[7973]), .Z(o[7973]) );
  AND U4508 ( .A(p_input[27973]), .B(p_input[17973]), .Z(n2254) );
  AND U4509 ( .A(n2255), .B(p_input[7972]), .Z(o[7972]) );
  AND U4510 ( .A(p_input[27972]), .B(p_input[17972]), .Z(n2255) );
  AND U4511 ( .A(n2256), .B(p_input[7971]), .Z(o[7971]) );
  AND U4512 ( .A(p_input[27971]), .B(p_input[17971]), .Z(n2256) );
  AND U4513 ( .A(n2257), .B(p_input[7970]), .Z(o[7970]) );
  AND U4514 ( .A(p_input[27970]), .B(p_input[17970]), .Z(n2257) );
  AND U4515 ( .A(n2258), .B(p_input[796]), .Z(o[796]) );
  AND U4516 ( .A(p_input[20796]), .B(p_input[10796]), .Z(n2258) );
  AND U4517 ( .A(n2259), .B(p_input[7969]), .Z(o[7969]) );
  AND U4518 ( .A(p_input[27969]), .B(p_input[17969]), .Z(n2259) );
  AND U4519 ( .A(n2260), .B(p_input[7968]), .Z(o[7968]) );
  AND U4520 ( .A(p_input[27968]), .B(p_input[17968]), .Z(n2260) );
  AND U4521 ( .A(n2261), .B(p_input[7967]), .Z(o[7967]) );
  AND U4522 ( .A(p_input[27967]), .B(p_input[17967]), .Z(n2261) );
  AND U4523 ( .A(n2262), .B(p_input[7966]), .Z(o[7966]) );
  AND U4524 ( .A(p_input[27966]), .B(p_input[17966]), .Z(n2262) );
  AND U4525 ( .A(n2263), .B(p_input[7965]), .Z(o[7965]) );
  AND U4526 ( .A(p_input[27965]), .B(p_input[17965]), .Z(n2263) );
  AND U4527 ( .A(n2264), .B(p_input[7964]), .Z(o[7964]) );
  AND U4528 ( .A(p_input[27964]), .B(p_input[17964]), .Z(n2264) );
  AND U4529 ( .A(n2265), .B(p_input[7963]), .Z(o[7963]) );
  AND U4530 ( .A(p_input[27963]), .B(p_input[17963]), .Z(n2265) );
  AND U4531 ( .A(n2266), .B(p_input[7962]), .Z(o[7962]) );
  AND U4532 ( .A(p_input[27962]), .B(p_input[17962]), .Z(n2266) );
  AND U4533 ( .A(n2267), .B(p_input[7961]), .Z(o[7961]) );
  AND U4534 ( .A(p_input[27961]), .B(p_input[17961]), .Z(n2267) );
  AND U4535 ( .A(n2268), .B(p_input[7960]), .Z(o[7960]) );
  AND U4536 ( .A(p_input[27960]), .B(p_input[17960]), .Z(n2268) );
  AND U4537 ( .A(n2269), .B(p_input[795]), .Z(o[795]) );
  AND U4538 ( .A(p_input[20795]), .B(p_input[10795]), .Z(n2269) );
  AND U4539 ( .A(n2270), .B(p_input[7959]), .Z(o[7959]) );
  AND U4540 ( .A(p_input[27959]), .B(p_input[17959]), .Z(n2270) );
  AND U4541 ( .A(n2271), .B(p_input[7958]), .Z(o[7958]) );
  AND U4542 ( .A(p_input[27958]), .B(p_input[17958]), .Z(n2271) );
  AND U4543 ( .A(n2272), .B(p_input[7957]), .Z(o[7957]) );
  AND U4544 ( .A(p_input[27957]), .B(p_input[17957]), .Z(n2272) );
  AND U4545 ( .A(n2273), .B(p_input[7956]), .Z(o[7956]) );
  AND U4546 ( .A(p_input[27956]), .B(p_input[17956]), .Z(n2273) );
  AND U4547 ( .A(n2274), .B(p_input[7955]), .Z(o[7955]) );
  AND U4548 ( .A(p_input[27955]), .B(p_input[17955]), .Z(n2274) );
  AND U4549 ( .A(n2275), .B(p_input[7954]), .Z(o[7954]) );
  AND U4550 ( .A(p_input[27954]), .B(p_input[17954]), .Z(n2275) );
  AND U4551 ( .A(n2276), .B(p_input[7953]), .Z(o[7953]) );
  AND U4552 ( .A(p_input[27953]), .B(p_input[17953]), .Z(n2276) );
  AND U4553 ( .A(n2277), .B(p_input[7952]), .Z(o[7952]) );
  AND U4554 ( .A(p_input[27952]), .B(p_input[17952]), .Z(n2277) );
  AND U4555 ( .A(n2278), .B(p_input[7951]), .Z(o[7951]) );
  AND U4556 ( .A(p_input[27951]), .B(p_input[17951]), .Z(n2278) );
  AND U4557 ( .A(n2279), .B(p_input[7950]), .Z(o[7950]) );
  AND U4558 ( .A(p_input[27950]), .B(p_input[17950]), .Z(n2279) );
  AND U4559 ( .A(n2280), .B(p_input[794]), .Z(o[794]) );
  AND U4560 ( .A(p_input[20794]), .B(p_input[10794]), .Z(n2280) );
  AND U4561 ( .A(n2281), .B(p_input[7949]), .Z(o[7949]) );
  AND U4562 ( .A(p_input[27949]), .B(p_input[17949]), .Z(n2281) );
  AND U4563 ( .A(n2282), .B(p_input[7948]), .Z(o[7948]) );
  AND U4564 ( .A(p_input[27948]), .B(p_input[17948]), .Z(n2282) );
  AND U4565 ( .A(n2283), .B(p_input[7947]), .Z(o[7947]) );
  AND U4566 ( .A(p_input[27947]), .B(p_input[17947]), .Z(n2283) );
  AND U4567 ( .A(n2284), .B(p_input[7946]), .Z(o[7946]) );
  AND U4568 ( .A(p_input[27946]), .B(p_input[17946]), .Z(n2284) );
  AND U4569 ( .A(n2285), .B(p_input[7945]), .Z(o[7945]) );
  AND U4570 ( .A(p_input[27945]), .B(p_input[17945]), .Z(n2285) );
  AND U4571 ( .A(n2286), .B(p_input[7944]), .Z(o[7944]) );
  AND U4572 ( .A(p_input[27944]), .B(p_input[17944]), .Z(n2286) );
  AND U4573 ( .A(n2287), .B(p_input[7943]), .Z(o[7943]) );
  AND U4574 ( .A(p_input[27943]), .B(p_input[17943]), .Z(n2287) );
  AND U4575 ( .A(n2288), .B(p_input[7942]), .Z(o[7942]) );
  AND U4576 ( .A(p_input[27942]), .B(p_input[17942]), .Z(n2288) );
  AND U4577 ( .A(n2289), .B(p_input[7941]), .Z(o[7941]) );
  AND U4578 ( .A(p_input[27941]), .B(p_input[17941]), .Z(n2289) );
  AND U4579 ( .A(n2290), .B(p_input[7940]), .Z(o[7940]) );
  AND U4580 ( .A(p_input[27940]), .B(p_input[17940]), .Z(n2290) );
  AND U4581 ( .A(n2291), .B(p_input[793]), .Z(o[793]) );
  AND U4582 ( .A(p_input[20793]), .B(p_input[10793]), .Z(n2291) );
  AND U4583 ( .A(n2292), .B(p_input[7939]), .Z(o[7939]) );
  AND U4584 ( .A(p_input[27939]), .B(p_input[17939]), .Z(n2292) );
  AND U4585 ( .A(n2293), .B(p_input[7938]), .Z(o[7938]) );
  AND U4586 ( .A(p_input[27938]), .B(p_input[17938]), .Z(n2293) );
  AND U4587 ( .A(n2294), .B(p_input[7937]), .Z(o[7937]) );
  AND U4588 ( .A(p_input[27937]), .B(p_input[17937]), .Z(n2294) );
  AND U4589 ( .A(n2295), .B(p_input[7936]), .Z(o[7936]) );
  AND U4590 ( .A(p_input[27936]), .B(p_input[17936]), .Z(n2295) );
  AND U4591 ( .A(n2296), .B(p_input[7935]), .Z(o[7935]) );
  AND U4592 ( .A(p_input[27935]), .B(p_input[17935]), .Z(n2296) );
  AND U4593 ( .A(n2297), .B(p_input[7934]), .Z(o[7934]) );
  AND U4594 ( .A(p_input[27934]), .B(p_input[17934]), .Z(n2297) );
  AND U4595 ( .A(n2298), .B(p_input[7933]), .Z(o[7933]) );
  AND U4596 ( .A(p_input[27933]), .B(p_input[17933]), .Z(n2298) );
  AND U4597 ( .A(n2299), .B(p_input[7932]), .Z(o[7932]) );
  AND U4598 ( .A(p_input[27932]), .B(p_input[17932]), .Z(n2299) );
  AND U4599 ( .A(n2300), .B(p_input[7931]), .Z(o[7931]) );
  AND U4600 ( .A(p_input[27931]), .B(p_input[17931]), .Z(n2300) );
  AND U4601 ( .A(n2301), .B(p_input[7930]), .Z(o[7930]) );
  AND U4602 ( .A(p_input[27930]), .B(p_input[17930]), .Z(n2301) );
  AND U4603 ( .A(n2302), .B(p_input[792]), .Z(o[792]) );
  AND U4604 ( .A(p_input[20792]), .B(p_input[10792]), .Z(n2302) );
  AND U4605 ( .A(n2303), .B(p_input[7929]), .Z(o[7929]) );
  AND U4606 ( .A(p_input[27929]), .B(p_input[17929]), .Z(n2303) );
  AND U4607 ( .A(n2304), .B(p_input[7928]), .Z(o[7928]) );
  AND U4608 ( .A(p_input[27928]), .B(p_input[17928]), .Z(n2304) );
  AND U4609 ( .A(n2305), .B(p_input[7927]), .Z(o[7927]) );
  AND U4610 ( .A(p_input[27927]), .B(p_input[17927]), .Z(n2305) );
  AND U4611 ( .A(n2306), .B(p_input[7926]), .Z(o[7926]) );
  AND U4612 ( .A(p_input[27926]), .B(p_input[17926]), .Z(n2306) );
  AND U4613 ( .A(n2307), .B(p_input[7925]), .Z(o[7925]) );
  AND U4614 ( .A(p_input[27925]), .B(p_input[17925]), .Z(n2307) );
  AND U4615 ( .A(n2308), .B(p_input[7924]), .Z(o[7924]) );
  AND U4616 ( .A(p_input[27924]), .B(p_input[17924]), .Z(n2308) );
  AND U4617 ( .A(n2309), .B(p_input[7923]), .Z(o[7923]) );
  AND U4618 ( .A(p_input[27923]), .B(p_input[17923]), .Z(n2309) );
  AND U4619 ( .A(n2310), .B(p_input[7922]), .Z(o[7922]) );
  AND U4620 ( .A(p_input[27922]), .B(p_input[17922]), .Z(n2310) );
  AND U4621 ( .A(n2311), .B(p_input[7921]), .Z(o[7921]) );
  AND U4622 ( .A(p_input[27921]), .B(p_input[17921]), .Z(n2311) );
  AND U4623 ( .A(n2312), .B(p_input[7920]), .Z(o[7920]) );
  AND U4624 ( .A(p_input[27920]), .B(p_input[17920]), .Z(n2312) );
  AND U4625 ( .A(n2313), .B(p_input[791]), .Z(o[791]) );
  AND U4626 ( .A(p_input[20791]), .B(p_input[10791]), .Z(n2313) );
  AND U4627 ( .A(n2314), .B(p_input[7919]), .Z(o[7919]) );
  AND U4628 ( .A(p_input[27919]), .B(p_input[17919]), .Z(n2314) );
  AND U4629 ( .A(n2315), .B(p_input[7918]), .Z(o[7918]) );
  AND U4630 ( .A(p_input[27918]), .B(p_input[17918]), .Z(n2315) );
  AND U4631 ( .A(n2316), .B(p_input[7917]), .Z(o[7917]) );
  AND U4632 ( .A(p_input[27917]), .B(p_input[17917]), .Z(n2316) );
  AND U4633 ( .A(n2317), .B(p_input[7916]), .Z(o[7916]) );
  AND U4634 ( .A(p_input[27916]), .B(p_input[17916]), .Z(n2317) );
  AND U4635 ( .A(n2318), .B(p_input[7915]), .Z(o[7915]) );
  AND U4636 ( .A(p_input[27915]), .B(p_input[17915]), .Z(n2318) );
  AND U4637 ( .A(n2319), .B(p_input[7914]), .Z(o[7914]) );
  AND U4638 ( .A(p_input[27914]), .B(p_input[17914]), .Z(n2319) );
  AND U4639 ( .A(n2320), .B(p_input[7913]), .Z(o[7913]) );
  AND U4640 ( .A(p_input[27913]), .B(p_input[17913]), .Z(n2320) );
  AND U4641 ( .A(n2321), .B(p_input[7912]), .Z(o[7912]) );
  AND U4642 ( .A(p_input[27912]), .B(p_input[17912]), .Z(n2321) );
  AND U4643 ( .A(n2322), .B(p_input[7911]), .Z(o[7911]) );
  AND U4644 ( .A(p_input[27911]), .B(p_input[17911]), .Z(n2322) );
  AND U4645 ( .A(n2323), .B(p_input[7910]), .Z(o[7910]) );
  AND U4646 ( .A(p_input[27910]), .B(p_input[17910]), .Z(n2323) );
  AND U4647 ( .A(n2324), .B(p_input[790]), .Z(o[790]) );
  AND U4648 ( .A(p_input[20790]), .B(p_input[10790]), .Z(n2324) );
  AND U4649 ( .A(n2325), .B(p_input[7909]), .Z(o[7909]) );
  AND U4650 ( .A(p_input[27909]), .B(p_input[17909]), .Z(n2325) );
  AND U4651 ( .A(n2326), .B(p_input[7908]), .Z(o[7908]) );
  AND U4652 ( .A(p_input[27908]), .B(p_input[17908]), .Z(n2326) );
  AND U4653 ( .A(n2327), .B(p_input[7907]), .Z(o[7907]) );
  AND U4654 ( .A(p_input[27907]), .B(p_input[17907]), .Z(n2327) );
  AND U4655 ( .A(n2328), .B(p_input[7906]), .Z(o[7906]) );
  AND U4656 ( .A(p_input[27906]), .B(p_input[17906]), .Z(n2328) );
  AND U4657 ( .A(n2329), .B(p_input[7905]), .Z(o[7905]) );
  AND U4658 ( .A(p_input[27905]), .B(p_input[17905]), .Z(n2329) );
  AND U4659 ( .A(n2330), .B(p_input[7904]), .Z(o[7904]) );
  AND U4660 ( .A(p_input[27904]), .B(p_input[17904]), .Z(n2330) );
  AND U4661 ( .A(n2331), .B(p_input[7903]), .Z(o[7903]) );
  AND U4662 ( .A(p_input[27903]), .B(p_input[17903]), .Z(n2331) );
  AND U4663 ( .A(n2332), .B(p_input[7902]), .Z(o[7902]) );
  AND U4664 ( .A(p_input[27902]), .B(p_input[17902]), .Z(n2332) );
  AND U4665 ( .A(n2333), .B(p_input[7901]), .Z(o[7901]) );
  AND U4666 ( .A(p_input[27901]), .B(p_input[17901]), .Z(n2333) );
  AND U4667 ( .A(n2334), .B(p_input[7900]), .Z(o[7900]) );
  AND U4668 ( .A(p_input[27900]), .B(p_input[17900]), .Z(n2334) );
  AND U4669 ( .A(n2335), .B(p_input[78]), .Z(o[78]) );
  AND U4670 ( .A(p_input[20078]), .B(p_input[10078]), .Z(n2335) );
  AND U4671 ( .A(n2336), .B(p_input[789]), .Z(o[789]) );
  AND U4672 ( .A(p_input[20789]), .B(p_input[10789]), .Z(n2336) );
  AND U4673 ( .A(n2337), .B(p_input[7899]), .Z(o[7899]) );
  AND U4674 ( .A(p_input[27899]), .B(p_input[17899]), .Z(n2337) );
  AND U4675 ( .A(n2338), .B(p_input[7898]), .Z(o[7898]) );
  AND U4676 ( .A(p_input[27898]), .B(p_input[17898]), .Z(n2338) );
  AND U4677 ( .A(n2339), .B(p_input[7897]), .Z(o[7897]) );
  AND U4678 ( .A(p_input[27897]), .B(p_input[17897]), .Z(n2339) );
  AND U4679 ( .A(n2340), .B(p_input[7896]), .Z(o[7896]) );
  AND U4680 ( .A(p_input[27896]), .B(p_input[17896]), .Z(n2340) );
  AND U4681 ( .A(n2341), .B(p_input[7895]), .Z(o[7895]) );
  AND U4682 ( .A(p_input[27895]), .B(p_input[17895]), .Z(n2341) );
  AND U4683 ( .A(n2342), .B(p_input[7894]), .Z(o[7894]) );
  AND U4684 ( .A(p_input[27894]), .B(p_input[17894]), .Z(n2342) );
  AND U4685 ( .A(n2343), .B(p_input[7893]), .Z(o[7893]) );
  AND U4686 ( .A(p_input[27893]), .B(p_input[17893]), .Z(n2343) );
  AND U4687 ( .A(n2344), .B(p_input[7892]), .Z(o[7892]) );
  AND U4688 ( .A(p_input[27892]), .B(p_input[17892]), .Z(n2344) );
  AND U4689 ( .A(n2345), .B(p_input[7891]), .Z(o[7891]) );
  AND U4690 ( .A(p_input[27891]), .B(p_input[17891]), .Z(n2345) );
  AND U4691 ( .A(n2346), .B(p_input[7890]), .Z(o[7890]) );
  AND U4692 ( .A(p_input[27890]), .B(p_input[17890]), .Z(n2346) );
  AND U4693 ( .A(n2347), .B(p_input[788]), .Z(o[788]) );
  AND U4694 ( .A(p_input[20788]), .B(p_input[10788]), .Z(n2347) );
  AND U4695 ( .A(n2348), .B(p_input[7889]), .Z(o[7889]) );
  AND U4696 ( .A(p_input[27889]), .B(p_input[17889]), .Z(n2348) );
  AND U4697 ( .A(n2349), .B(p_input[7888]), .Z(o[7888]) );
  AND U4698 ( .A(p_input[27888]), .B(p_input[17888]), .Z(n2349) );
  AND U4699 ( .A(n2350), .B(p_input[7887]), .Z(o[7887]) );
  AND U4700 ( .A(p_input[27887]), .B(p_input[17887]), .Z(n2350) );
  AND U4701 ( .A(n2351), .B(p_input[7886]), .Z(o[7886]) );
  AND U4702 ( .A(p_input[27886]), .B(p_input[17886]), .Z(n2351) );
  AND U4703 ( .A(n2352), .B(p_input[7885]), .Z(o[7885]) );
  AND U4704 ( .A(p_input[27885]), .B(p_input[17885]), .Z(n2352) );
  AND U4705 ( .A(n2353), .B(p_input[7884]), .Z(o[7884]) );
  AND U4706 ( .A(p_input[27884]), .B(p_input[17884]), .Z(n2353) );
  AND U4707 ( .A(n2354), .B(p_input[7883]), .Z(o[7883]) );
  AND U4708 ( .A(p_input[27883]), .B(p_input[17883]), .Z(n2354) );
  AND U4709 ( .A(n2355), .B(p_input[7882]), .Z(o[7882]) );
  AND U4710 ( .A(p_input[27882]), .B(p_input[17882]), .Z(n2355) );
  AND U4711 ( .A(n2356), .B(p_input[7881]), .Z(o[7881]) );
  AND U4712 ( .A(p_input[27881]), .B(p_input[17881]), .Z(n2356) );
  AND U4713 ( .A(n2357), .B(p_input[7880]), .Z(o[7880]) );
  AND U4714 ( .A(p_input[27880]), .B(p_input[17880]), .Z(n2357) );
  AND U4715 ( .A(n2358), .B(p_input[787]), .Z(o[787]) );
  AND U4716 ( .A(p_input[20787]), .B(p_input[10787]), .Z(n2358) );
  AND U4717 ( .A(n2359), .B(p_input[7879]), .Z(o[7879]) );
  AND U4718 ( .A(p_input[27879]), .B(p_input[17879]), .Z(n2359) );
  AND U4719 ( .A(n2360), .B(p_input[7878]), .Z(o[7878]) );
  AND U4720 ( .A(p_input[27878]), .B(p_input[17878]), .Z(n2360) );
  AND U4721 ( .A(n2361), .B(p_input[7877]), .Z(o[7877]) );
  AND U4722 ( .A(p_input[27877]), .B(p_input[17877]), .Z(n2361) );
  AND U4723 ( .A(n2362), .B(p_input[7876]), .Z(o[7876]) );
  AND U4724 ( .A(p_input[27876]), .B(p_input[17876]), .Z(n2362) );
  AND U4725 ( .A(n2363), .B(p_input[7875]), .Z(o[7875]) );
  AND U4726 ( .A(p_input[27875]), .B(p_input[17875]), .Z(n2363) );
  AND U4727 ( .A(n2364), .B(p_input[7874]), .Z(o[7874]) );
  AND U4728 ( .A(p_input[27874]), .B(p_input[17874]), .Z(n2364) );
  AND U4729 ( .A(n2365), .B(p_input[7873]), .Z(o[7873]) );
  AND U4730 ( .A(p_input[27873]), .B(p_input[17873]), .Z(n2365) );
  AND U4731 ( .A(n2366), .B(p_input[7872]), .Z(o[7872]) );
  AND U4732 ( .A(p_input[27872]), .B(p_input[17872]), .Z(n2366) );
  AND U4733 ( .A(n2367), .B(p_input[7871]), .Z(o[7871]) );
  AND U4734 ( .A(p_input[27871]), .B(p_input[17871]), .Z(n2367) );
  AND U4735 ( .A(n2368), .B(p_input[7870]), .Z(o[7870]) );
  AND U4736 ( .A(p_input[27870]), .B(p_input[17870]), .Z(n2368) );
  AND U4737 ( .A(n2369), .B(p_input[786]), .Z(o[786]) );
  AND U4738 ( .A(p_input[20786]), .B(p_input[10786]), .Z(n2369) );
  AND U4739 ( .A(n2370), .B(p_input[7869]), .Z(o[7869]) );
  AND U4740 ( .A(p_input[27869]), .B(p_input[17869]), .Z(n2370) );
  AND U4741 ( .A(n2371), .B(p_input[7868]), .Z(o[7868]) );
  AND U4742 ( .A(p_input[27868]), .B(p_input[17868]), .Z(n2371) );
  AND U4743 ( .A(n2372), .B(p_input[7867]), .Z(o[7867]) );
  AND U4744 ( .A(p_input[27867]), .B(p_input[17867]), .Z(n2372) );
  AND U4745 ( .A(n2373), .B(p_input[7866]), .Z(o[7866]) );
  AND U4746 ( .A(p_input[27866]), .B(p_input[17866]), .Z(n2373) );
  AND U4747 ( .A(n2374), .B(p_input[7865]), .Z(o[7865]) );
  AND U4748 ( .A(p_input[27865]), .B(p_input[17865]), .Z(n2374) );
  AND U4749 ( .A(n2375), .B(p_input[7864]), .Z(o[7864]) );
  AND U4750 ( .A(p_input[27864]), .B(p_input[17864]), .Z(n2375) );
  AND U4751 ( .A(n2376), .B(p_input[7863]), .Z(o[7863]) );
  AND U4752 ( .A(p_input[27863]), .B(p_input[17863]), .Z(n2376) );
  AND U4753 ( .A(n2377), .B(p_input[7862]), .Z(o[7862]) );
  AND U4754 ( .A(p_input[27862]), .B(p_input[17862]), .Z(n2377) );
  AND U4755 ( .A(n2378), .B(p_input[7861]), .Z(o[7861]) );
  AND U4756 ( .A(p_input[27861]), .B(p_input[17861]), .Z(n2378) );
  AND U4757 ( .A(n2379), .B(p_input[7860]), .Z(o[7860]) );
  AND U4758 ( .A(p_input[27860]), .B(p_input[17860]), .Z(n2379) );
  AND U4759 ( .A(n2380), .B(p_input[785]), .Z(o[785]) );
  AND U4760 ( .A(p_input[20785]), .B(p_input[10785]), .Z(n2380) );
  AND U4761 ( .A(n2381), .B(p_input[7859]), .Z(o[7859]) );
  AND U4762 ( .A(p_input[27859]), .B(p_input[17859]), .Z(n2381) );
  AND U4763 ( .A(n2382), .B(p_input[7858]), .Z(o[7858]) );
  AND U4764 ( .A(p_input[27858]), .B(p_input[17858]), .Z(n2382) );
  AND U4765 ( .A(n2383), .B(p_input[7857]), .Z(o[7857]) );
  AND U4766 ( .A(p_input[27857]), .B(p_input[17857]), .Z(n2383) );
  AND U4767 ( .A(n2384), .B(p_input[7856]), .Z(o[7856]) );
  AND U4768 ( .A(p_input[27856]), .B(p_input[17856]), .Z(n2384) );
  AND U4769 ( .A(n2385), .B(p_input[7855]), .Z(o[7855]) );
  AND U4770 ( .A(p_input[27855]), .B(p_input[17855]), .Z(n2385) );
  AND U4771 ( .A(n2386), .B(p_input[7854]), .Z(o[7854]) );
  AND U4772 ( .A(p_input[27854]), .B(p_input[17854]), .Z(n2386) );
  AND U4773 ( .A(n2387), .B(p_input[7853]), .Z(o[7853]) );
  AND U4774 ( .A(p_input[27853]), .B(p_input[17853]), .Z(n2387) );
  AND U4775 ( .A(n2388), .B(p_input[7852]), .Z(o[7852]) );
  AND U4776 ( .A(p_input[27852]), .B(p_input[17852]), .Z(n2388) );
  AND U4777 ( .A(n2389), .B(p_input[7851]), .Z(o[7851]) );
  AND U4778 ( .A(p_input[27851]), .B(p_input[17851]), .Z(n2389) );
  AND U4779 ( .A(n2390), .B(p_input[7850]), .Z(o[7850]) );
  AND U4780 ( .A(p_input[27850]), .B(p_input[17850]), .Z(n2390) );
  AND U4781 ( .A(n2391), .B(p_input[784]), .Z(o[784]) );
  AND U4782 ( .A(p_input[20784]), .B(p_input[10784]), .Z(n2391) );
  AND U4783 ( .A(n2392), .B(p_input[7849]), .Z(o[7849]) );
  AND U4784 ( .A(p_input[27849]), .B(p_input[17849]), .Z(n2392) );
  AND U4785 ( .A(n2393), .B(p_input[7848]), .Z(o[7848]) );
  AND U4786 ( .A(p_input[27848]), .B(p_input[17848]), .Z(n2393) );
  AND U4787 ( .A(n2394), .B(p_input[7847]), .Z(o[7847]) );
  AND U4788 ( .A(p_input[27847]), .B(p_input[17847]), .Z(n2394) );
  AND U4789 ( .A(n2395), .B(p_input[7846]), .Z(o[7846]) );
  AND U4790 ( .A(p_input[27846]), .B(p_input[17846]), .Z(n2395) );
  AND U4791 ( .A(n2396), .B(p_input[7845]), .Z(o[7845]) );
  AND U4792 ( .A(p_input[27845]), .B(p_input[17845]), .Z(n2396) );
  AND U4793 ( .A(n2397), .B(p_input[7844]), .Z(o[7844]) );
  AND U4794 ( .A(p_input[27844]), .B(p_input[17844]), .Z(n2397) );
  AND U4795 ( .A(n2398), .B(p_input[7843]), .Z(o[7843]) );
  AND U4796 ( .A(p_input[27843]), .B(p_input[17843]), .Z(n2398) );
  AND U4797 ( .A(n2399), .B(p_input[7842]), .Z(o[7842]) );
  AND U4798 ( .A(p_input[27842]), .B(p_input[17842]), .Z(n2399) );
  AND U4799 ( .A(n2400), .B(p_input[7841]), .Z(o[7841]) );
  AND U4800 ( .A(p_input[27841]), .B(p_input[17841]), .Z(n2400) );
  AND U4801 ( .A(n2401), .B(p_input[7840]), .Z(o[7840]) );
  AND U4802 ( .A(p_input[27840]), .B(p_input[17840]), .Z(n2401) );
  AND U4803 ( .A(n2402), .B(p_input[783]), .Z(o[783]) );
  AND U4804 ( .A(p_input[20783]), .B(p_input[10783]), .Z(n2402) );
  AND U4805 ( .A(n2403), .B(p_input[7839]), .Z(o[7839]) );
  AND U4806 ( .A(p_input[27839]), .B(p_input[17839]), .Z(n2403) );
  AND U4807 ( .A(n2404), .B(p_input[7838]), .Z(o[7838]) );
  AND U4808 ( .A(p_input[27838]), .B(p_input[17838]), .Z(n2404) );
  AND U4809 ( .A(n2405), .B(p_input[7837]), .Z(o[7837]) );
  AND U4810 ( .A(p_input[27837]), .B(p_input[17837]), .Z(n2405) );
  AND U4811 ( .A(n2406), .B(p_input[7836]), .Z(o[7836]) );
  AND U4812 ( .A(p_input[27836]), .B(p_input[17836]), .Z(n2406) );
  AND U4813 ( .A(n2407), .B(p_input[7835]), .Z(o[7835]) );
  AND U4814 ( .A(p_input[27835]), .B(p_input[17835]), .Z(n2407) );
  AND U4815 ( .A(n2408), .B(p_input[7834]), .Z(o[7834]) );
  AND U4816 ( .A(p_input[27834]), .B(p_input[17834]), .Z(n2408) );
  AND U4817 ( .A(n2409), .B(p_input[7833]), .Z(o[7833]) );
  AND U4818 ( .A(p_input[27833]), .B(p_input[17833]), .Z(n2409) );
  AND U4819 ( .A(n2410), .B(p_input[7832]), .Z(o[7832]) );
  AND U4820 ( .A(p_input[27832]), .B(p_input[17832]), .Z(n2410) );
  AND U4821 ( .A(n2411), .B(p_input[7831]), .Z(o[7831]) );
  AND U4822 ( .A(p_input[27831]), .B(p_input[17831]), .Z(n2411) );
  AND U4823 ( .A(n2412), .B(p_input[7830]), .Z(o[7830]) );
  AND U4824 ( .A(p_input[27830]), .B(p_input[17830]), .Z(n2412) );
  AND U4825 ( .A(n2413), .B(p_input[782]), .Z(o[782]) );
  AND U4826 ( .A(p_input[20782]), .B(p_input[10782]), .Z(n2413) );
  AND U4827 ( .A(n2414), .B(p_input[7829]), .Z(o[7829]) );
  AND U4828 ( .A(p_input[27829]), .B(p_input[17829]), .Z(n2414) );
  AND U4829 ( .A(n2415), .B(p_input[7828]), .Z(o[7828]) );
  AND U4830 ( .A(p_input[27828]), .B(p_input[17828]), .Z(n2415) );
  AND U4831 ( .A(n2416), .B(p_input[7827]), .Z(o[7827]) );
  AND U4832 ( .A(p_input[27827]), .B(p_input[17827]), .Z(n2416) );
  AND U4833 ( .A(n2417), .B(p_input[7826]), .Z(o[7826]) );
  AND U4834 ( .A(p_input[27826]), .B(p_input[17826]), .Z(n2417) );
  AND U4835 ( .A(n2418), .B(p_input[7825]), .Z(o[7825]) );
  AND U4836 ( .A(p_input[27825]), .B(p_input[17825]), .Z(n2418) );
  AND U4837 ( .A(n2419), .B(p_input[7824]), .Z(o[7824]) );
  AND U4838 ( .A(p_input[27824]), .B(p_input[17824]), .Z(n2419) );
  AND U4839 ( .A(n2420), .B(p_input[7823]), .Z(o[7823]) );
  AND U4840 ( .A(p_input[27823]), .B(p_input[17823]), .Z(n2420) );
  AND U4841 ( .A(n2421), .B(p_input[7822]), .Z(o[7822]) );
  AND U4842 ( .A(p_input[27822]), .B(p_input[17822]), .Z(n2421) );
  AND U4843 ( .A(n2422), .B(p_input[7821]), .Z(o[7821]) );
  AND U4844 ( .A(p_input[27821]), .B(p_input[17821]), .Z(n2422) );
  AND U4845 ( .A(n2423), .B(p_input[7820]), .Z(o[7820]) );
  AND U4846 ( .A(p_input[27820]), .B(p_input[17820]), .Z(n2423) );
  AND U4847 ( .A(n2424), .B(p_input[781]), .Z(o[781]) );
  AND U4848 ( .A(p_input[20781]), .B(p_input[10781]), .Z(n2424) );
  AND U4849 ( .A(n2425), .B(p_input[7819]), .Z(o[7819]) );
  AND U4850 ( .A(p_input[27819]), .B(p_input[17819]), .Z(n2425) );
  AND U4851 ( .A(n2426), .B(p_input[7818]), .Z(o[7818]) );
  AND U4852 ( .A(p_input[27818]), .B(p_input[17818]), .Z(n2426) );
  AND U4853 ( .A(n2427), .B(p_input[7817]), .Z(o[7817]) );
  AND U4854 ( .A(p_input[27817]), .B(p_input[17817]), .Z(n2427) );
  AND U4855 ( .A(n2428), .B(p_input[7816]), .Z(o[7816]) );
  AND U4856 ( .A(p_input[27816]), .B(p_input[17816]), .Z(n2428) );
  AND U4857 ( .A(n2429), .B(p_input[7815]), .Z(o[7815]) );
  AND U4858 ( .A(p_input[27815]), .B(p_input[17815]), .Z(n2429) );
  AND U4859 ( .A(n2430), .B(p_input[7814]), .Z(o[7814]) );
  AND U4860 ( .A(p_input[27814]), .B(p_input[17814]), .Z(n2430) );
  AND U4861 ( .A(n2431), .B(p_input[7813]), .Z(o[7813]) );
  AND U4862 ( .A(p_input[27813]), .B(p_input[17813]), .Z(n2431) );
  AND U4863 ( .A(n2432), .B(p_input[7812]), .Z(o[7812]) );
  AND U4864 ( .A(p_input[27812]), .B(p_input[17812]), .Z(n2432) );
  AND U4865 ( .A(n2433), .B(p_input[7811]), .Z(o[7811]) );
  AND U4866 ( .A(p_input[27811]), .B(p_input[17811]), .Z(n2433) );
  AND U4867 ( .A(n2434), .B(p_input[7810]), .Z(o[7810]) );
  AND U4868 ( .A(p_input[27810]), .B(p_input[17810]), .Z(n2434) );
  AND U4869 ( .A(n2435), .B(p_input[780]), .Z(o[780]) );
  AND U4870 ( .A(p_input[20780]), .B(p_input[10780]), .Z(n2435) );
  AND U4871 ( .A(n2436), .B(p_input[7809]), .Z(o[7809]) );
  AND U4872 ( .A(p_input[27809]), .B(p_input[17809]), .Z(n2436) );
  AND U4873 ( .A(n2437), .B(p_input[7808]), .Z(o[7808]) );
  AND U4874 ( .A(p_input[27808]), .B(p_input[17808]), .Z(n2437) );
  AND U4875 ( .A(n2438), .B(p_input[7807]), .Z(o[7807]) );
  AND U4876 ( .A(p_input[27807]), .B(p_input[17807]), .Z(n2438) );
  AND U4877 ( .A(n2439), .B(p_input[7806]), .Z(o[7806]) );
  AND U4878 ( .A(p_input[27806]), .B(p_input[17806]), .Z(n2439) );
  AND U4879 ( .A(n2440), .B(p_input[7805]), .Z(o[7805]) );
  AND U4880 ( .A(p_input[27805]), .B(p_input[17805]), .Z(n2440) );
  AND U4881 ( .A(n2441), .B(p_input[7804]), .Z(o[7804]) );
  AND U4882 ( .A(p_input[27804]), .B(p_input[17804]), .Z(n2441) );
  AND U4883 ( .A(n2442), .B(p_input[7803]), .Z(o[7803]) );
  AND U4884 ( .A(p_input[27803]), .B(p_input[17803]), .Z(n2442) );
  AND U4885 ( .A(n2443), .B(p_input[7802]), .Z(o[7802]) );
  AND U4886 ( .A(p_input[27802]), .B(p_input[17802]), .Z(n2443) );
  AND U4887 ( .A(n2444), .B(p_input[7801]), .Z(o[7801]) );
  AND U4888 ( .A(p_input[27801]), .B(p_input[17801]), .Z(n2444) );
  AND U4889 ( .A(n2445), .B(p_input[7800]), .Z(o[7800]) );
  AND U4890 ( .A(p_input[27800]), .B(p_input[17800]), .Z(n2445) );
  AND U4891 ( .A(n2446), .B(p_input[77]), .Z(o[77]) );
  AND U4892 ( .A(p_input[20077]), .B(p_input[10077]), .Z(n2446) );
  AND U4893 ( .A(n2447), .B(p_input[779]), .Z(o[779]) );
  AND U4894 ( .A(p_input[20779]), .B(p_input[10779]), .Z(n2447) );
  AND U4895 ( .A(n2448), .B(p_input[7799]), .Z(o[7799]) );
  AND U4896 ( .A(p_input[27799]), .B(p_input[17799]), .Z(n2448) );
  AND U4897 ( .A(n2449), .B(p_input[7798]), .Z(o[7798]) );
  AND U4898 ( .A(p_input[27798]), .B(p_input[17798]), .Z(n2449) );
  AND U4899 ( .A(n2450), .B(p_input[7797]), .Z(o[7797]) );
  AND U4900 ( .A(p_input[27797]), .B(p_input[17797]), .Z(n2450) );
  AND U4901 ( .A(n2451), .B(p_input[7796]), .Z(o[7796]) );
  AND U4902 ( .A(p_input[27796]), .B(p_input[17796]), .Z(n2451) );
  AND U4903 ( .A(n2452), .B(p_input[7795]), .Z(o[7795]) );
  AND U4904 ( .A(p_input[27795]), .B(p_input[17795]), .Z(n2452) );
  AND U4905 ( .A(n2453), .B(p_input[7794]), .Z(o[7794]) );
  AND U4906 ( .A(p_input[27794]), .B(p_input[17794]), .Z(n2453) );
  AND U4907 ( .A(n2454), .B(p_input[7793]), .Z(o[7793]) );
  AND U4908 ( .A(p_input[27793]), .B(p_input[17793]), .Z(n2454) );
  AND U4909 ( .A(n2455), .B(p_input[7792]), .Z(o[7792]) );
  AND U4910 ( .A(p_input[27792]), .B(p_input[17792]), .Z(n2455) );
  AND U4911 ( .A(n2456), .B(p_input[7791]), .Z(o[7791]) );
  AND U4912 ( .A(p_input[27791]), .B(p_input[17791]), .Z(n2456) );
  AND U4913 ( .A(n2457), .B(p_input[7790]), .Z(o[7790]) );
  AND U4914 ( .A(p_input[27790]), .B(p_input[17790]), .Z(n2457) );
  AND U4915 ( .A(n2458), .B(p_input[778]), .Z(o[778]) );
  AND U4916 ( .A(p_input[20778]), .B(p_input[10778]), .Z(n2458) );
  AND U4917 ( .A(n2459), .B(p_input[7789]), .Z(o[7789]) );
  AND U4918 ( .A(p_input[27789]), .B(p_input[17789]), .Z(n2459) );
  AND U4919 ( .A(n2460), .B(p_input[7788]), .Z(o[7788]) );
  AND U4920 ( .A(p_input[27788]), .B(p_input[17788]), .Z(n2460) );
  AND U4921 ( .A(n2461), .B(p_input[7787]), .Z(o[7787]) );
  AND U4922 ( .A(p_input[27787]), .B(p_input[17787]), .Z(n2461) );
  AND U4923 ( .A(n2462), .B(p_input[7786]), .Z(o[7786]) );
  AND U4924 ( .A(p_input[27786]), .B(p_input[17786]), .Z(n2462) );
  AND U4925 ( .A(n2463), .B(p_input[7785]), .Z(o[7785]) );
  AND U4926 ( .A(p_input[27785]), .B(p_input[17785]), .Z(n2463) );
  AND U4927 ( .A(n2464), .B(p_input[7784]), .Z(o[7784]) );
  AND U4928 ( .A(p_input[27784]), .B(p_input[17784]), .Z(n2464) );
  AND U4929 ( .A(n2465), .B(p_input[7783]), .Z(o[7783]) );
  AND U4930 ( .A(p_input[27783]), .B(p_input[17783]), .Z(n2465) );
  AND U4931 ( .A(n2466), .B(p_input[7782]), .Z(o[7782]) );
  AND U4932 ( .A(p_input[27782]), .B(p_input[17782]), .Z(n2466) );
  AND U4933 ( .A(n2467), .B(p_input[7781]), .Z(o[7781]) );
  AND U4934 ( .A(p_input[27781]), .B(p_input[17781]), .Z(n2467) );
  AND U4935 ( .A(n2468), .B(p_input[7780]), .Z(o[7780]) );
  AND U4936 ( .A(p_input[27780]), .B(p_input[17780]), .Z(n2468) );
  AND U4937 ( .A(n2469), .B(p_input[777]), .Z(o[777]) );
  AND U4938 ( .A(p_input[20777]), .B(p_input[10777]), .Z(n2469) );
  AND U4939 ( .A(n2470), .B(p_input[7779]), .Z(o[7779]) );
  AND U4940 ( .A(p_input[27779]), .B(p_input[17779]), .Z(n2470) );
  AND U4941 ( .A(n2471), .B(p_input[7778]), .Z(o[7778]) );
  AND U4942 ( .A(p_input[27778]), .B(p_input[17778]), .Z(n2471) );
  AND U4943 ( .A(n2472), .B(p_input[7777]), .Z(o[7777]) );
  AND U4944 ( .A(p_input[27777]), .B(p_input[17777]), .Z(n2472) );
  AND U4945 ( .A(n2473), .B(p_input[7776]), .Z(o[7776]) );
  AND U4946 ( .A(p_input[27776]), .B(p_input[17776]), .Z(n2473) );
  AND U4947 ( .A(n2474), .B(p_input[7775]), .Z(o[7775]) );
  AND U4948 ( .A(p_input[27775]), .B(p_input[17775]), .Z(n2474) );
  AND U4949 ( .A(n2475), .B(p_input[7774]), .Z(o[7774]) );
  AND U4950 ( .A(p_input[27774]), .B(p_input[17774]), .Z(n2475) );
  AND U4951 ( .A(n2476), .B(p_input[7773]), .Z(o[7773]) );
  AND U4952 ( .A(p_input[27773]), .B(p_input[17773]), .Z(n2476) );
  AND U4953 ( .A(n2477), .B(p_input[7772]), .Z(o[7772]) );
  AND U4954 ( .A(p_input[27772]), .B(p_input[17772]), .Z(n2477) );
  AND U4955 ( .A(n2478), .B(p_input[7771]), .Z(o[7771]) );
  AND U4956 ( .A(p_input[27771]), .B(p_input[17771]), .Z(n2478) );
  AND U4957 ( .A(n2479), .B(p_input[7770]), .Z(o[7770]) );
  AND U4958 ( .A(p_input[27770]), .B(p_input[17770]), .Z(n2479) );
  AND U4959 ( .A(n2480), .B(p_input[776]), .Z(o[776]) );
  AND U4960 ( .A(p_input[20776]), .B(p_input[10776]), .Z(n2480) );
  AND U4961 ( .A(n2481), .B(p_input[7769]), .Z(o[7769]) );
  AND U4962 ( .A(p_input[27769]), .B(p_input[17769]), .Z(n2481) );
  AND U4963 ( .A(n2482), .B(p_input[7768]), .Z(o[7768]) );
  AND U4964 ( .A(p_input[27768]), .B(p_input[17768]), .Z(n2482) );
  AND U4965 ( .A(n2483), .B(p_input[7767]), .Z(o[7767]) );
  AND U4966 ( .A(p_input[27767]), .B(p_input[17767]), .Z(n2483) );
  AND U4967 ( .A(n2484), .B(p_input[7766]), .Z(o[7766]) );
  AND U4968 ( .A(p_input[27766]), .B(p_input[17766]), .Z(n2484) );
  AND U4969 ( .A(n2485), .B(p_input[7765]), .Z(o[7765]) );
  AND U4970 ( .A(p_input[27765]), .B(p_input[17765]), .Z(n2485) );
  AND U4971 ( .A(n2486), .B(p_input[7764]), .Z(o[7764]) );
  AND U4972 ( .A(p_input[27764]), .B(p_input[17764]), .Z(n2486) );
  AND U4973 ( .A(n2487), .B(p_input[7763]), .Z(o[7763]) );
  AND U4974 ( .A(p_input[27763]), .B(p_input[17763]), .Z(n2487) );
  AND U4975 ( .A(n2488), .B(p_input[7762]), .Z(o[7762]) );
  AND U4976 ( .A(p_input[27762]), .B(p_input[17762]), .Z(n2488) );
  AND U4977 ( .A(n2489), .B(p_input[7761]), .Z(o[7761]) );
  AND U4978 ( .A(p_input[27761]), .B(p_input[17761]), .Z(n2489) );
  AND U4979 ( .A(n2490), .B(p_input[7760]), .Z(o[7760]) );
  AND U4980 ( .A(p_input[27760]), .B(p_input[17760]), .Z(n2490) );
  AND U4981 ( .A(n2491), .B(p_input[775]), .Z(o[775]) );
  AND U4982 ( .A(p_input[20775]), .B(p_input[10775]), .Z(n2491) );
  AND U4983 ( .A(n2492), .B(p_input[7759]), .Z(o[7759]) );
  AND U4984 ( .A(p_input[27759]), .B(p_input[17759]), .Z(n2492) );
  AND U4985 ( .A(n2493), .B(p_input[7758]), .Z(o[7758]) );
  AND U4986 ( .A(p_input[27758]), .B(p_input[17758]), .Z(n2493) );
  AND U4987 ( .A(n2494), .B(p_input[7757]), .Z(o[7757]) );
  AND U4988 ( .A(p_input[27757]), .B(p_input[17757]), .Z(n2494) );
  AND U4989 ( .A(n2495), .B(p_input[7756]), .Z(o[7756]) );
  AND U4990 ( .A(p_input[27756]), .B(p_input[17756]), .Z(n2495) );
  AND U4991 ( .A(n2496), .B(p_input[7755]), .Z(o[7755]) );
  AND U4992 ( .A(p_input[27755]), .B(p_input[17755]), .Z(n2496) );
  AND U4993 ( .A(n2497), .B(p_input[7754]), .Z(o[7754]) );
  AND U4994 ( .A(p_input[27754]), .B(p_input[17754]), .Z(n2497) );
  AND U4995 ( .A(n2498), .B(p_input[7753]), .Z(o[7753]) );
  AND U4996 ( .A(p_input[27753]), .B(p_input[17753]), .Z(n2498) );
  AND U4997 ( .A(n2499), .B(p_input[7752]), .Z(o[7752]) );
  AND U4998 ( .A(p_input[27752]), .B(p_input[17752]), .Z(n2499) );
  AND U4999 ( .A(n2500), .B(p_input[7751]), .Z(o[7751]) );
  AND U5000 ( .A(p_input[27751]), .B(p_input[17751]), .Z(n2500) );
  AND U5001 ( .A(n2501), .B(p_input[7750]), .Z(o[7750]) );
  AND U5002 ( .A(p_input[27750]), .B(p_input[17750]), .Z(n2501) );
  AND U5003 ( .A(n2502), .B(p_input[774]), .Z(o[774]) );
  AND U5004 ( .A(p_input[20774]), .B(p_input[10774]), .Z(n2502) );
  AND U5005 ( .A(n2503), .B(p_input[7749]), .Z(o[7749]) );
  AND U5006 ( .A(p_input[27749]), .B(p_input[17749]), .Z(n2503) );
  AND U5007 ( .A(n2504), .B(p_input[7748]), .Z(o[7748]) );
  AND U5008 ( .A(p_input[27748]), .B(p_input[17748]), .Z(n2504) );
  AND U5009 ( .A(n2505), .B(p_input[7747]), .Z(o[7747]) );
  AND U5010 ( .A(p_input[27747]), .B(p_input[17747]), .Z(n2505) );
  AND U5011 ( .A(n2506), .B(p_input[7746]), .Z(o[7746]) );
  AND U5012 ( .A(p_input[27746]), .B(p_input[17746]), .Z(n2506) );
  AND U5013 ( .A(n2507), .B(p_input[7745]), .Z(o[7745]) );
  AND U5014 ( .A(p_input[27745]), .B(p_input[17745]), .Z(n2507) );
  AND U5015 ( .A(n2508), .B(p_input[7744]), .Z(o[7744]) );
  AND U5016 ( .A(p_input[27744]), .B(p_input[17744]), .Z(n2508) );
  AND U5017 ( .A(n2509), .B(p_input[7743]), .Z(o[7743]) );
  AND U5018 ( .A(p_input[27743]), .B(p_input[17743]), .Z(n2509) );
  AND U5019 ( .A(n2510), .B(p_input[7742]), .Z(o[7742]) );
  AND U5020 ( .A(p_input[27742]), .B(p_input[17742]), .Z(n2510) );
  AND U5021 ( .A(n2511), .B(p_input[7741]), .Z(o[7741]) );
  AND U5022 ( .A(p_input[27741]), .B(p_input[17741]), .Z(n2511) );
  AND U5023 ( .A(n2512), .B(p_input[7740]), .Z(o[7740]) );
  AND U5024 ( .A(p_input[27740]), .B(p_input[17740]), .Z(n2512) );
  AND U5025 ( .A(n2513), .B(p_input[773]), .Z(o[773]) );
  AND U5026 ( .A(p_input[20773]), .B(p_input[10773]), .Z(n2513) );
  AND U5027 ( .A(n2514), .B(p_input[7739]), .Z(o[7739]) );
  AND U5028 ( .A(p_input[27739]), .B(p_input[17739]), .Z(n2514) );
  AND U5029 ( .A(n2515), .B(p_input[7738]), .Z(o[7738]) );
  AND U5030 ( .A(p_input[27738]), .B(p_input[17738]), .Z(n2515) );
  AND U5031 ( .A(n2516), .B(p_input[7737]), .Z(o[7737]) );
  AND U5032 ( .A(p_input[27737]), .B(p_input[17737]), .Z(n2516) );
  AND U5033 ( .A(n2517), .B(p_input[7736]), .Z(o[7736]) );
  AND U5034 ( .A(p_input[27736]), .B(p_input[17736]), .Z(n2517) );
  AND U5035 ( .A(n2518), .B(p_input[7735]), .Z(o[7735]) );
  AND U5036 ( .A(p_input[27735]), .B(p_input[17735]), .Z(n2518) );
  AND U5037 ( .A(n2519), .B(p_input[7734]), .Z(o[7734]) );
  AND U5038 ( .A(p_input[27734]), .B(p_input[17734]), .Z(n2519) );
  AND U5039 ( .A(n2520), .B(p_input[7733]), .Z(o[7733]) );
  AND U5040 ( .A(p_input[27733]), .B(p_input[17733]), .Z(n2520) );
  AND U5041 ( .A(n2521), .B(p_input[7732]), .Z(o[7732]) );
  AND U5042 ( .A(p_input[27732]), .B(p_input[17732]), .Z(n2521) );
  AND U5043 ( .A(n2522), .B(p_input[7731]), .Z(o[7731]) );
  AND U5044 ( .A(p_input[27731]), .B(p_input[17731]), .Z(n2522) );
  AND U5045 ( .A(n2523), .B(p_input[7730]), .Z(o[7730]) );
  AND U5046 ( .A(p_input[27730]), .B(p_input[17730]), .Z(n2523) );
  AND U5047 ( .A(n2524), .B(p_input[772]), .Z(o[772]) );
  AND U5048 ( .A(p_input[20772]), .B(p_input[10772]), .Z(n2524) );
  AND U5049 ( .A(n2525), .B(p_input[7729]), .Z(o[7729]) );
  AND U5050 ( .A(p_input[27729]), .B(p_input[17729]), .Z(n2525) );
  AND U5051 ( .A(n2526), .B(p_input[7728]), .Z(o[7728]) );
  AND U5052 ( .A(p_input[27728]), .B(p_input[17728]), .Z(n2526) );
  AND U5053 ( .A(n2527), .B(p_input[7727]), .Z(o[7727]) );
  AND U5054 ( .A(p_input[27727]), .B(p_input[17727]), .Z(n2527) );
  AND U5055 ( .A(n2528), .B(p_input[7726]), .Z(o[7726]) );
  AND U5056 ( .A(p_input[27726]), .B(p_input[17726]), .Z(n2528) );
  AND U5057 ( .A(n2529), .B(p_input[7725]), .Z(o[7725]) );
  AND U5058 ( .A(p_input[27725]), .B(p_input[17725]), .Z(n2529) );
  AND U5059 ( .A(n2530), .B(p_input[7724]), .Z(o[7724]) );
  AND U5060 ( .A(p_input[27724]), .B(p_input[17724]), .Z(n2530) );
  AND U5061 ( .A(n2531), .B(p_input[7723]), .Z(o[7723]) );
  AND U5062 ( .A(p_input[27723]), .B(p_input[17723]), .Z(n2531) );
  AND U5063 ( .A(n2532), .B(p_input[7722]), .Z(o[7722]) );
  AND U5064 ( .A(p_input[27722]), .B(p_input[17722]), .Z(n2532) );
  AND U5065 ( .A(n2533), .B(p_input[7721]), .Z(o[7721]) );
  AND U5066 ( .A(p_input[27721]), .B(p_input[17721]), .Z(n2533) );
  AND U5067 ( .A(n2534), .B(p_input[7720]), .Z(o[7720]) );
  AND U5068 ( .A(p_input[27720]), .B(p_input[17720]), .Z(n2534) );
  AND U5069 ( .A(n2535), .B(p_input[771]), .Z(o[771]) );
  AND U5070 ( .A(p_input[20771]), .B(p_input[10771]), .Z(n2535) );
  AND U5071 ( .A(n2536), .B(p_input[7719]), .Z(o[7719]) );
  AND U5072 ( .A(p_input[27719]), .B(p_input[17719]), .Z(n2536) );
  AND U5073 ( .A(n2537), .B(p_input[7718]), .Z(o[7718]) );
  AND U5074 ( .A(p_input[27718]), .B(p_input[17718]), .Z(n2537) );
  AND U5075 ( .A(n2538), .B(p_input[7717]), .Z(o[7717]) );
  AND U5076 ( .A(p_input[27717]), .B(p_input[17717]), .Z(n2538) );
  AND U5077 ( .A(n2539), .B(p_input[7716]), .Z(o[7716]) );
  AND U5078 ( .A(p_input[27716]), .B(p_input[17716]), .Z(n2539) );
  AND U5079 ( .A(n2540), .B(p_input[7715]), .Z(o[7715]) );
  AND U5080 ( .A(p_input[27715]), .B(p_input[17715]), .Z(n2540) );
  AND U5081 ( .A(n2541), .B(p_input[7714]), .Z(o[7714]) );
  AND U5082 ( .A(p_input[27714]), .B(p_input[17714]), .Z(n2541) );
  AND U5083 ( .A(n2542), .B(p_input[7713]), .Z(o[7713]) );
  AND U5084 ( .A(p_input[27713]), .B(p_input[17713]), .Z(n2542) );
  AND U5085 ( .A(n2543), .B(p_input[7712]), .Z(o[7712]) );
  AND U5086 ( .A(p_input[27712]), .B(p_input[17712]), .Z(n2543) );
  AND U5087 ( .A(n2544), .B(p_input[7711]), .Z(o[7711]) );
  AND U5088 ( .A(p_input[27711]), .B(p_input[17711]), .Z(n2544) );
  AND U5089 ( .A(n2545), .B(p_input[7710]), .Z(o[7710]) );
  AND U5090 ( .A(p_input[27710]), .B(p_input[17710]), .Z(n2545) );
  AND U5091 ( .A(n2546), .B(p_input[770]), .Z(o[770]) );
  AND U5092 ( .A(p_input[20770]), .B(p_input[10770]), .Z(n2546) );
  AND U5093 ( .A(n2547), .B(p_input[7709]), .Z(o[7709]) );
  AND U5094 ( .A(p_input[27709]), .B(p_input[17709]), .Z(n2547) );
  AND U5095 ( .A(n2548), .B(p_input[7708]), .Z(o[7708]) );
  AND U5096 ( .A(p_input[27708]), .B(p_input[17708]), .Z(n2548) );
  AND U5097 ( .A(n2549), .B(p_input[7707]), .Z(o[7707]) );
  AND U5098 ( .A(p_input[27707]), .B(p_input[17707]), .Z(n2549) );
  AND U5099 ( .A(n2550), .B(p_input[7706]), .Z(o[7706]) );
  AND U5100 ( .A(p_input[27706]), .B(p_input[17706]), .Z(n2550) );
  AND U5101 ( .A(n2551), .B(p_input[7705]), .Z(o[7705]) );
  AND U5102 ( .A(p_input[27705]), .B(p_input[17705]), .Z(n2551) );
  AND U5103 ( .A(n2552), .B(p_input[7704]), .Z(o[7704]) );
  AND U5104 ( .A(p_input[27704]), .B(p_input[17704]), .Z(n2552) );
  AND U5105 ( .A(n2553), .B(p_input[7703]), .Z(o[7703]) );
  AND U5106 ( .A(p_input[27703]), .B(p_input[17703]), .Z(n2553) );
  AND U5107 ( .A(n2554), .B(p_input[7702]), .Z(o[7702]) );
  AND U5108 ( .A(p_input[27702]), .B(p_input[17702]), .Z(n2554) );
  AND U5109 ( .A(n2555), .B(p_input[7701]), .Z(o[7701]) );
  AND U5110 ( .A(p_input[27701]), .B(p_input[17701]), .Z(n2555) );
  AND U5111 ( .A(n2556), .B(p_input[7700]), .Z(o[7700]) );
  AND U5112 ( .A(p_input[27700]), .B(p_input[17700]), .Z(n2556) );
  AND U5113 ( .A(n2557), .B(p_input[76]), .Z(o[76]) );
  AND U5114 ( .A(p_input[20076]), .B(p_input[10076]), .Z(n2557) );
  AND U5115 ( .A(n2558), .B(p_input[769]), .Z(o[769]) );
  AND U5116 ( .A(p_input[20769]), .B(p_input[10769]), .Z(n2558) );
  AND U5117 ( .A(n2559), .B(p_input[7699]), .Z(o[7699]) );
  AND U5118 ( .A(p_input[27699]), .B(p_input[17699]), .Z(n2559) );
  AND U5119 ( .A(n2560), .B(p_input[7698]), .Z(o[7698]) );
  AND U5120 ( .A(p_input[27698]), .B(p_input[17698]), .Z(n2560) );
  AND U5121 ( .A(n2561), .B(p_input[7697]), .Z(o[7697]) );
  AND U5122 ( .A(p_input[27697]), .B(p_input[17697]), .Z(n2561) );
  AND U5123 ( .A(n2562), .B(p_input[7696]), .Z(o[7696]) );
  AND U5124 ( .A(p_input[27696]), .B(p_input[17696]), .Z(n2562) );
  AND U5125 ( .A(n2563), .B(p_input[7695]), .Z(o[7695]) );
  AND U5126 ( .A(p_input[27695]), .B(p_input[17695]), .Z(n2563) );
  AND U5127 ( .A(n2564), .B(p_input[7694]), .Z(o[7694]) );
  AND U5128 ( .A(p_input[27694]), .B(p_input[17694]), .Z(n2564) );
  AND U5129 ( .A(n2565), .B(p_input[7693]), .Z(o[7693]) );
  AND U5130 ( .A(p_input[27693]), .B(p_input[17693]), .Z(n2565) );
  AND U5131 ( .A(n2566), .B(p_input[7692]), .Z(o[7692]) );
  AND U5132 ( .A(p_input[27692]), .B(p_input[17692]), .Z(n2566) );
  AND U5133 ( .A(n2567), .B(p_input[7691]), .Z(o[7691]) );
  AND U5134 ( .A(p_input[27691]), .B(p_input[17691]), .Z(n2567) );
  AND U5135 ( .A(n2568), .B(p_input[7690]), .Z(o[7690]) );
  AND U5136 ( .A(p_input[27690]), .B(p_input[17690]), .Z(n2568) );
  AND U5137 ( .A(n2569), .B(p_input[768]), .Z(o[768]) );
  AND U5138 ( .A(p_input[20768]), .B(p_input[10768]), .Z(n2569) );
  AND U5139 ( .A(n2570), .B(p_input[7689]), .Z(o[7689]) );
  AND U5140 ( .A(p_input[27689]), .B(p_input[17689]), .Z(n2570) );
  AND U5141 ( .A(n2571), .B(p_input[7688]), .Z(o[7688]) );
  AND U5142 ( .A(p_input[27688]), .B(p_input[17688]), .Z(n2571) );
  AND U5143 ( .A(n2572), .B(p_input[7687]), .Z(o[7687]) );
  AND U5144 ( .A(p_input[27687]), .B(p_input[17687]), .Z(n2572) );
  AND U5145 ( .A(n2573), .B(p_input[7686]), .Z(o[7686]) );
  AND U5146 ( .A(p_input[27686]), .B(p_input[17686]), .Z(n2573) );
  AND U5147 ( .A(n2574), .B(p_input[7685]), .Z(o[7685]) );
  AND U5148 ( .A(p_input[27685]), .B(p_input[17685]), .Z(n2574) );
  AND U5149 ( .A(n2575), .B(p_input[7684]), .Z(o[7684]) );
  AND U5150 ( .A(p_input[27684]), .B(p_input[17684]), .Z(n2575) );
  AND U5151 ( .A(n2576), .B(p_input[7683]), .Z(o[7683]) );
  AND U5152 ( .A(p_input[27683]), .B(p_input[17683]), .Z(n2576) );
  AND U5153 ( .A(n2577), .B(p_input[7682]), .Z(o[7682]) );
  AND U5154 ( .A(p_input[27682]), .B(p_input[17682]), .Z(n2577) );
  AND U5155 ( .A(n2578), .B(p_input[7681]), .Z(o[7681]) );
  AND U5156 ( .A(p_input[27681]), .B(p_input[17681]), .Z(n2578) );
  AND U5157 ( .A(n2579), .B(p_input[7680]), .Z(o[7680]) );
  AND U5158 ( .A(p_input[27680]), .B(p_input[17680]), .Z(n2579) );
  AND U5159 ( .A(n2580), .B(p_input[767]), .Z(o[767]) );
  AND U5160 ( .A(p_input[20767]), .B(p_input[10767]), .Z(n2580) );
  AND U5161 ( .A(n2581), .B(p_input[7679]), .Z(o[7679]) );
  AND U5162 ( .A(p_input[27679]), .B(p_input[17679]), .Z(n2581) );
  AND U5163 ( .A(n2582), .B(p_input[7678]), .Z(o[7678]) );
  AND U5164 ( .A(p_input[27678]), .B(p_input[17678]), .Z(n2582) );
  AND U5165 ( .A(n2583), .B(p_input[7677]), .Z(o[7677]) );
  AND U5166 ( .A(p_input[27677]), .B(p_input[17677]), .Z(n2583) );
  AND U5167 ( .A(n2584), .B(p_input[7676]), .Z(o[7676]) );
  AND U5168 ( .A(p_input[27676]), .B(p_input[17676]), .Z(n2584) );
  AND U5169 ( .A(n2585), .B(p_input[7675]), .Z(o[7675]) );
  AND U5170 ( .A(p_input[27675]), .B(p_input[17675]), .Z(n2585) );
  AND U5171 ( .A(n2586), .B(p_input[7674]), .Z(o[7674]) );
  AND U5172 ( .A(p_input[27674]), .B(p_input[17674]), .Z(n2586) );
  AND U5173 ( .A(n2587), .B(p_input[7673]), .Z(o[7673]) );
  AND U5174 ( .A(p_input[27673]), .B(p_input[17673]), .Z(n2587) );
  AND U5175 ( .A(n2588), .B(p_input[7672]), .Z(o[7672]) );
  AND U5176 ( .A(p_input[27672]), .B(p_input[17672]), .Z(n2588) );
  AND U5177 ( .A(n2589), .B(p_input[7671]), .Z(o[7671]) );
  AND U5178 ( .A(p_input[27671]), .B(p_input[17671]), .Z(n2589) );
  AND U5179 ( .A(n2590), .B(p_input[7670]), .Z(o[7670]) );
  AND U5180 ( .A(p_input[27670]), .B(p_input[17670]), .Z(n2590) );
  AND U5181 ( .A(n2591), .B(p_input[766]), .Z(o[766]) );
  AND U5182 ( .A(p_input[20766]), .B(p_input[10766]), .Z(n2591) );
  AND U5183 ( .A(n2592), .B(p_input[7669]), .Z(o[7669]) );
  AND U5184 ( .A(p_input[27669]), .B(p_input[17669]), .Z(n2592) );
  AND U5185 ( .A(n2593), .B(p_input[7668]), .Z(o[7668]) );
  AND U5186 ( .A(p_input[27668]), .B(p_input[17668]), .Z(n2593) );
  AND U5187 ( .A(n2594), .B(p_input[7667]), .Z(o[7667]) );
  AND U5188 ( .A(p_input[27667]), .B(p_input[17667]), .Z(n2594) );
  AND U5189 ( .A(n2595), .B(p_input[7666]), .Z(o[7666]) );
  AND U5190 ( .A(p_input[27666]), .B(p_input[17666]), .Z(n2595) );
  AND U5191 ( .A(n2596), .B(p_input[7665]), .Z(o[7665]) );
  AND U5192 ( .A(p_input[27665]), .B(p_input[17665]), .Z(n2596) );
  AND U5193 ( .A(n2597), .B(p_input[7664]), .Z(o[7664]) );
  AND U5194 ( .A(p_input[27664]), .B(p_input[17664]), .Z(n2597) );
  AND U5195 ( .A(n2598), .B(p_input[7663]), .Z(o[7663]) );
  AND U5196 ( .A(p_input[27663]), .B(p_input[17663]), .Z(n2598) );
  AND U5197 ( .A(n2599), .B(p_input[7662]), .Z(o[7662]) );
  AND U5198 ( .A(p_input[27662]), .B(p_input[17662]), .Z(n2599) );
  AND U5199 ( .A(n2600), .B(p_input[7661]), .Z(o[7661]) );
  AND U5200 ( .A(p_input[27661]), .B(p_input[17661]), .Z(n2600) );
  AND U5201 ( .A(n2601), .B(p_input[7660]), .Z(o[7660]) );
  AND U5202 ( .A(p_input[27660]), .B(p_input[17660]), .Z(n2601) );
  AND U5203 ( .A(n2602), .B(p_input[765]), .Z(o[765]) );
  AND U5204 ( .A(p_input[20765]), .B(p_input[10765]), .Z(n2602) );
  AND U5205 ( .A(n2603), .B(p_input[7659]), .Z(o[7659]) );
  AND U5206 ( .A(p_input[27659]), .B(p_input[17659]), .Z(n2603) );
  AND U5207 ( .A(n2604), .B(p_input[7658]), .Z(o[7658]) );
  AND U5208 ( .A(p_input[27658]), .B(p_input[17658]), .Z(n2604) );
  AND U5209 ( .A(n2605), .B(p_input[7657]), .Z(o[7657]) );
  AND U5210 ( .A(p_input[27657]), .B(p_input[17657]), .Z(n2605) );
  AND U5211 ( .A(n2606), .B(p_input[7656]), .Z(o[7656]) );
  AND U5212 ( .A(p_input[27656]), .B(p_input[17656]), .Z(n2606) );
  AND U5213 ( .A(n2607), .B(p_input[7655]), .Z(o[7655]) );
  AND U5214 ( .A(p_input[27655]), .B(p_input[17655]), .Z(n2607) );
  AND U5215 ( .A(n2608), .B(p_input[7654]), .Z(o[7654]) );
  AND U5216 ( .A(p_input[27654]), .B(p_input[17654]), .Z(n2608) );
  AND U5217 ( .A(n2609), .B(p_input[7653]), .Z(o[7653]) );
  AND U5218 ( .A(p_input[27653]), .B(p_input[17653]), .Z(n2609) );
  AND U5219 ( .A(n2610), .B(p_input[7652]), .Z(o[7652]) );
  AND U5220 ( .A(p_input[27652]), .B(p_input[17652]), .Z(n2610) );
  AND U5221 ( .A(n2611), .B(p_input[7651]), .Z(o[7651]) );
  AND U5222 ( .A(p_input[27651]), .B(p_input[17651]), .Z(n2611) );
  AND U5223 ( .A(n2612), .B(p_input[7650]), .Z(o[7650]) );
  AND U5224 ( .A(p_input[27650]), .B(p_input[17650]), .Z(n2612) );
  AND U5225 ( .A(n2613), .B(p_input[764]), .Z(o[764]) );
  AND U5226 ( .A(p_input[20764]), .B(p_input[10764]), .Z(n2613) );
  AND U5227 ( .A(n2614), .B(p_input[7649]), .Z(o[7649]) );
  AND U5228 ( .A(p_input[27649]), .B(p_input[17649]), .Z(n2614) );
  AND U5229 ( .A(n2615), .B(p_input[7648]), .Z(o[7648]) );
  AND U5230 ( .A(p_input[27648]), .B(p_input[17648]), .Z(n2615) );
  AND U5231 ( .A(n2616), .B(p_input[7647]), .Z(o[7647]) );
  AND U5232 ( .A(p_input[27647]), .B(p_input[17647]), .Z(n2616) );
  AND U5233 ( .A(n2617), .B(p_input[7646]), .Z(o[7646]) );
  AND U5234 ( .A(p_input[27646]), .B(p_input[17646]), .Z(n2617) );
  AND U5235 ( .A(n2618), .B(p_input[7645]), .Z(o[7645]) );
  AND U5236 ( .A(p_input[27645]), .B(p_input[17645]), .Z(n2618) );
  AND U5237 ( .A(n2619), .B(p_input[7644]), .Z(o[7644]) );
  AND U5238 ( .A(p_input[27644]), .B(p_input[17644]), .Z(n2619) );
  AND U5239 ( .A(n2620), .B(p_input[7643]), .Z(o[7643]) );
  AND U5240 ( .A(p_input[27643]), .B(p_input[17643]), .Z(n2620) );
  AND U5241 ( .A(n2621), .B(p_input[7642]), .Z(o[7642]) );
  AND U5242 ( .A(p_input[27642]), .B(p_input[17642]), .Z(n2621) );
  AND U5243 ( .A(n2622), .B(p_input[7641]), .Z(o[7641]) );
  AND U5244 ( .A(p_input[27641]), .B(p_input[17641]), .Z(n2622) );
  AND U5245 ( .A(n2623), .B(p_input[7640]), .Z(o[7640]) );
  AND U5246 ( .A(p_input[27640]), .B(p_input[17640]), .Z(n2623) );
  AND U5247 ( .A(n2624), .B(p_input[763]), .Z(o[763]) );
  AND U5248 ( .A(p_input[20763]), .B(p_input[10763]), .Z(n2624) );
  AND U5249 ( .A(n2625), .B(p_input[7639]), .Z(o[7639]) );
  AND U5250 ( .A(p_input[27639]), .B(p_input[17639]), .Z(n2625) );
  AND U5251 ( .A(n2626), .B(p_input[7638]), .Z(o[7638]) );
  AND U5252 ( .A(p_input[27638]), .B(p_input[17638]), .Z(n2626) );
  AND U5253 ( .A(n2627), .B(p_input[7637]), .Z(o[7637]) );
  AND U5254 ( .A(p_input[27637]), .B(p_input[17637]), .Z(n2627) );
  AND U5255 ( .A(n2628), .B(p_input[7636]), .Z(o[7636]) );
  AND U5256 ( .A(p_input[27636]), .B(p_input[17636]), .Z(n2628) );
  AND U5257 ( .A(n2629), .B(p_input[7635]), .Z(o[7635]) );
  AND U5258 ( .A(p_input[27635]), .B(p_input[17635]), .Z(n2629) );
  AND U5259 ( .A(n2630), .B(p_input[7634]), .Z(o[7634]) );
  AND U5260 ( .A(p_input[27634]), .B(p_input[17634]), .Z(n2630) );
  AND U5261 ( .A(n2631), .B(p_input[7633]), .Z(o[7633]) );
  AND U5262 ( .A(p_input[27633]), .B(p_input[17633]), .Z(n2631) );
  AND U5263 ( .A(n2632), .B(p_input[7632]), .Z(o[7632]) );
  AND U5264 ( .A(p_input[27632]), .B(p_input[17632]), .Z(n2632) );
  AND U5265 ( .A(n2633), .B(p_input[7631]), .Z(o[7631]) );
  AND U5266 ( .A(p_input[27631]), .B(p_input[17631]), .Z(n2633) );
  AND U5267 ( .A(n2634), .B(p_input[7630]), .Z(o[7630]) );
  AND U5268 ( .A(p_input[27630]), .B(p_input[17630]), .Z(n2634) );
  AND U5269 ( .A(n2635), .B(p_input[762]), .Z(o[762]) );
  AND U5270 ( .A(p_input[20762]), .B(p_input[10762]), .Z(n2635) );
  AND U5271 ( .A(n2636), .B(p_input[7629]), .Z(o[7629]) );
  AND U5272 ( .A(p_input[27629]), .B(p_input[17629]), .Z(n2636) );
  AND U5273 ( .A(n2637), .B(p_input[7628]), .Z(o[7628]) );
  AND U5274 ( .A(p_input[27628]), .B(p_input[17628]), .Z(n2637) );
  AND U5275 ( .A(n2638), .B(p_input[7627]), .Z(o[7627]) );
  AND U5276 ( .A(p_input[27627]), .B(p_input[17627]), .Z(n2638) );
  AND U5277 ( .A(n2639), .B(p_input[7626]), .Z(o[7626]) );
  AND U5278 ( .A(p_input[27626]), .B(p_input[17626]), .Z(n2639) );
  AND U5279 ( .A(n2640), .B(p_input[7625]), .Z(o[7625]) );
  AND U5280 ( .A(p_input[27625]), .B(p_input[17625]), .Z(n2640) );
  AND U5281 ( .A(n2641), .B(p_input[7624]), .Z(o[7624]) );
  AND U5282 ( .A(p_input[27624]), .B(p_input[17624]), .Z(n2641) );
  AND U5283 ( .A(n2642), .B(p_input[7623]), .Z(o[7623]) );
  AND U5284 ( .A(p_input[27623]), .B(p_input[17623]), .Z(n2642) );
  AND U5285 ( .A(n2643), .B(p_input[7622]), .Z(o[7622]) );
  AND U5286 ( .A(p_input[27622]), .B(p_input[17622]), .Z(n2643) );
  AND U5287 ( .A(n2644), .B(p_input[7621]), .Z(o[7621]) );
  AND U5288 ( .A(p_input[27621]), .B(p_input[17621]), .Z(n2644) );
  AND U5289 ( .A(n2645), .B(p_input[7620]), .Z(o[7620]) );
  AND U5290 ( .A(p_input[27620]), .B(p_input[17620]), .Z(n2645) );
  AND U5291 ( .A(n2646), .B(p_input[761]), .Z(o[761]) );
  AND U5292 ( .A(p_input[20761]), .B(p_input[10761]), .Z(n2646) );
  AND U5293 ( .A(n2647), .B(p_input[7619]), .Z(o[7619]) );
  AND U5294 ( .A(p_input[27619]), .B(p_input[17619]), .Z(n2647) );
  AND U5295 ( .A(n2648), .B(p_input[7618]), .Z(o[7618]) );
  AND U5296 ( .A(p_input[27618]), .B(p_input[17618]), .Z(n2648) );
  AND U5297 ( .A(n2649), .B(p_input[7617]), .Z(o[7617]) );
  AND U5298 ( .A(p_input[27617]), .B(p_input[17617]), .Z(n2649) );
  AND U5299 ( .A(n2650), .B(p_input[7616]), .Z(o[7616]) );
  AND U5300 ( .A(p_input[27616]), .B(p_input[17616]), .Z(n2650) );
  AND U5301 ( .A(n2651), .B(p_input[7615]), .Z(o[7615]) );
  AND U5302 ( .A(p_input[27615]), .B(p_input[17615]), .Z(n2651) );
  AND U5303 ( .A(n2652), .B(p_input[7614]), .Z(o[7614]) );
  AND U5304 ( .A(p_input[27614]), .B(p_input[17614]), .Z(n2652) );
  AND U5305 ( .A(n2653), .B(p_input[7613]), .Z(o[7613]) );
  AND U5306 ( .A(p_input[27613]), .B(p_input[17613]), .Z(n2653) );
  AND U5307 ( .A(n2654), .B(p_input[7612]), .Z(o[7612]) );
  AND U5308 ( .A(p_input[27612]), .B(p_input[17612]), .Z(n2654) );
  AND U5309 ( .A(n2655), .B(p_input[7611]), .Z(o[7611]) );
  AND U5310 ( .A(p_input[27611]), .B(p_input[17611]), .Z(n2655) );
  AND U5311 ( .A(n2656), .B(p_input[7610]), .Z(o[7610]) );
  AND U5312 ( .A(p_input[27610]), .B(p_input[17610]), .Z(n2656) );
  AND U5313 ( .A(n2657), .B(p_input[760]), .Z(o[760]) );
  AND U5314 ( .A(p_input[20760]), .B(p_input[10760]), .Z(n2657) );
  AND U5315 ( .A(n2658), .B(p_input[7609]), .Z(o[7609]) );
  AND U5316 ( .A(p_input[27609]), .B(p_input[17609]), .Z(n2658) );
  AND U5317 ( .A(n2659), .B(p_input[7608]), .Z(o[7608]) );
  AND U5318 ( .A(p_input[27608]), .B(p_input[17608]), .Z(n2659) );
  AND U5319 ( .A(n2660), .B(p_input[7607]), .Z(o[7607]) );
  AND U5320 ( .A(p_input[27607]), .B(p_input[17607]), .Z(n2660) );
  AND U5321 ( .A(n2661), .B(p_input[7606]), .Z(o[7606]) );
  AND U5322 ( .A(p_input[27606]), .B(p_input[17606]), .Z(n2661) );
  AND U5323 ( .A(n2662), .B(p_input[7605]), .Z(o[7605]) );
  AND U5324 ( .A(p_input[27605]), .B(p_input[17605]), .Z(n2662) );
  AND U5325 ( .A(n2663), .B(p_input[7604]), .Z(o[7604]) );
  AND U5326 ( .A(p_input[27604]), .B(p_input[17604]), .Z(n2663) );
  AND U5327 ( .A(n2664), .B(p_input[7603]), .Z(o[7603]) );
  AND U5328 ( .A(p_input[27603]), .B(p_input[17603]), .Z(n2664) );
  AND U5329 ( .A(n2665), .B(p_input[7602]), .Z(o[7602]) );
  AND U5330 ( .A(p_input[27602]), .B(p_input[17602]), .Z(n2665) );
  AND U5331 ( .A(n2666), .B(p_input[7601]), .Z(o[7601]) );
  AND U5332 ( .A(p_input[27601]), .B(p_input[17601]), .Z(n2666) );
  AND U5333 ( .A(n2667), .B(p_input[7600]), .Z(o[7600]) );
  AND U5334 ( .A(p_input[27600]), .B(p_input[17600]), .Z(n2667) );
  AND U5335 ( .A(n2668), .B(p_input[75]), .Z(o[75]) );
  AND U5336 ( .A(p_input[20075]), .B(p_input[10075]), .Z(n2668) );
  AND U5337 ( .A(n2669), .B(p_input[759]), .Z(o[759]) );
  AND U5338 ( .A(p_input[20759]), .B(p_input[10759]), .Z(n2669) );
  AND U5339 ( .A(n2670), .B(p_input[7599]), .Z(o[7599]) );
  AND U5340 ( .A(p_input[27599]), .B(p_input[17599]), .Z(n2670) );
  AND U5341 ( .A(n2671), .B(p_input[7598]), .Z(o[7598]) );
  AND U5342 ( .A(p_input[27598]), .B(p_input[17598]), .Z(n2671) );
  AND U5343 ( .A(n2672), .B(p_input[7597]), .Z(o[7597]) );
  AND U5344 ( .A(p_input[27597]), .B(p_input[17597]), .Z(n2672) );
  AND U5345 ( .A(n2673), .B(p_input[7596]), .Z(o[7596]) );
  AND U5346 ( .A(p_input[27596]), .B(p_input[17596]), .Z(n2673) );
  AND U5347 ( .A(n2674), .B(p_input[7595]), .Z(o[7595]) );
  AND U5348 ( .A(p_input[27595]), .B(p_input[17595]), .Z(n2674) );
  AND U5349 ( .A(n2675), .B(p_input[7594]), .Z(o[7594]) );
  AND U5350 ( .A(p_input[27594]), .B(p_input[17594]), .Z(n2675) );
  AND U5351 ( .A(n2676), .B(p_input[7593]), .Z(o[7593]) );
  AND U5352 ( .A(p_input[27593]), .B(p_input[17593]), .Z(n2676) );
  AND U5353 ( .A(n2677), .B(p_input[7592]), .Z(o[7592]) );
  AND U5354 ( .A(p_input[27592]), .B(p_input[17592]), .Z(n2677) );
  AND U5355 ( .A(n2678), .B(p_input[7591]), .Z(o[7591]) );
  AND U5356 ( .A(p_input[27591]), .B(p_input[17591]), .Z(n2678) );
  AND U5357 ( .A(n2679), .B(p_input[7590]), .Z(o[7590]) );
  AND U5358 ( .A(p_input[27590]), .B(p_input[17590]), .Z(n2679) );
  AND U5359 ( .A(n2680), .B(p_input[758]), .Z(o[758]) );
  AND U5360 ( .A(p_input[20758]), .B(p_input[10758]), .Z(n2680) );
  AND U5361 ( .A(n2681), .B(p_input[7589]), .Z(o[7589]) );
  AND U5362 ( .A(p_input[27589]), .B(p_input[17589]), .Z(n2681) );
  AND U5363 ( .A(n2682), .B(p_input[7588]), .Z(o[7588]) );
  AND U5364 ( .A(p_input[27588]), .B(p_input[17588]), .Z(n2682) );
  AND U5365 ( .A(n2683), .B(p_input[7587]), .Z(o[7587]) );
  AND U5366 ( .A(p_input[27587]), .B(p_input[17587]), .Z(n2683) );
  AND U5367 ( .A(n2684), .B(p_input[7586]), .Z(o[7586]) );
  AND U5368 ( .A(p_input[27586]), .B(p_input[17586]), .Z(n2684) );
  AND U5369 ( .A(n2685), .B(p_input[7585]), .Z(o[7585]) );
  AND U5370 ( .A(p_input[27585]), .B(p_input[17585]), .Z(n2685) );
  AND U5371 ( .A(n2686), .B(p_input[7584]), .Z(o[7584]) );
  AND U5372 ( .A(p_input[27584]), .B(p_input[17584]), .Z(n2686) );
  AND U5373 ( .A(n2687), .B(p_input[7583]), .Z(o[7583]) );
  AND U5374 ( .A(p_input[27583]), .B(p_input[17583]), .Z(n2687) );
  AND U5375 ( .A(n2688), .B(p_input[7582]), .Z(o[7582]) );
  AND U5376 ( .A(p_input[27582]), .B(p_input[17582]), .Z(n2688) );
  AND U5377 ( .A(n2689), .B(p_input[7581]), .Z(o[7581]) );
  AND U5378 ( .A(p_input[27581]), .B(p_input[17581]), .Z(n2689) );
  AND U5379 ( .A(n2690), .B(p_input[7580]), .Z(o[7580]) );
  AND U5380 ( .A(p_input[27580]), .B(p_input[17580]), .Z(n2690) );
  AND U5381 ( .A(n2691), .B(p_input[757]), .Z(o[757]) );
  AND U5382 ( .A(p_input[20757]), .B(p_input[10757]), .Z(n2691) );
  AND U5383 ( .A(n2692), .B(p_input[7579]), .Z(o[7579]) );
  AND U5384 ( .A(p_input[27579]), .B(p_input[17579]), .Z(n2692) );
  AND U5385 ( .A(n2693), .B(p_input[7578]), .Z(o[7578]) );
  AND U5386 ( .A(p_input[27578]), .B(p_input[17578]), .Z(n2693) );
  AND U5387 ( .A(n2694), .B(p_input[7577]), .Z(o[7577]) );
  AND U5388 ( .A(p_input[27577]), .B(p_input[17577]), .Z(n2694) );
  AND U5389 ( .A(n2695), .B(p_input[7576]), .Z(o[7576]) );
  AND U5390 ( .A(p_input[27576]), .B(p_input[17576]), .Z(n2695) );
  AND U5391 ( .A(n2696), .B(p_input[7575]), .Z(o[7575]) );
  AND U5392 ( .A(p_input[27575]), .B(p_input[17575]), .Z(n2696) );
  AND U5393 ( .A(n2697), .B(p_input[7574]), .Z(o[7574]) );
  AND U5394 ( .A(p_input[27574]), .B(p_input[17574]), .Z(n2697) );
  AND U5395 ( .A(n2698), .B(p_input[7573]), .Z(o[7573]) );
  AND U5396 ( .A(p_input[27573]), .B(p_input[17573]), .Z(n2698) );
  AND U5397 ( .A(n2699), .B(p_input[7572]), .Z(o[7572]) );
  AND U5398 ( .A(p_input[27572]), .B(p_input[17572]), .Z(n2699) );
  AND U5399 ( .A(n2700), .B(p_input[7571]), .Z(o[7571]) );
  AND U5400 ( .A(p_input[27571]), .B(p_input[17571]), .Z(n2700) );
  AND U5401 ( .A(n2701), .B(p_input[7570]), .Z(o[7570]) );
  AND U5402 ( .A(p_input[27570]), .B(p_input[17570]), .Z(n2701) );
  AND U5403 ( .A(n2702), .B(p_input[756]), .Z(o[756]) );
  AND U5404 ( .A(p_input[20756]), .B(p_input[10756]), .Z(n2702) );
  AND U5405 ( .A(n2703), .B(p_input[7569]), .Z(o[7569]) );
  AND U5406 ( .A(p_input[27569]), .B(p_input[17569]), .Z(n2703) );
  AND U5407 ( .A(n2704), .B(p_input[7568]), .Z(o[7568]) );
  AND U5408 ( .A(p_input[27568]), .B(p_input[17568]), .Z(n2704) );
  AND U5409 ( .A(n2705), .B(p_input[7567]), .Z(o[7567]) );
  AND U5410 ( .A(p_input[27567]), .B(p_input[17567]), .Z(n2705) );
  AND U5411 ( .A(n2706), .B(p_input[7566]), .Z(o[7566]) );
  AND U5412 ( .A(p_input[27566]), .B(p_input[17566]), .Z(n2706) );
  AND U5413 ( .A(n2707), .B(p_input[7565]), .Z(o[7565]) );
  AND U5414 ( .A(p_input[27565]), .B(p_input[17565]), .Z(n2707) );
  AND U5415 ( .A(n2708), .B(p_input[7564]), .Z(o[7564]) );
  AND U5416 ( .A(p_input[27564]), .B(p_input[17564]), .Z(n2708) );
  AND U5417 ( .A(n2709), .B(p_input[7563]), .Z(o[7563]) );
  AND U5418 ( .A(p_input[27563]), .B(p_input[17563]), .Z(n2709) );
  AND U5419 ( .A(n2710), .B(p_input[7562]), .Z(o[7562]) );
  AND U5420 ( .A(p_input[27562]), .B(p_input[17562]), .Z(n2710) );
  AND U5421 ( .A(n2711), .B(p_input[7561]), .Z(o[7561]) );
  AND U5422 ( .A(p_input[27561]), .B(p_input[17561]), .Z(n2711) );
  AND U5423 ( .A(n2712), .B(p_input[7560]), .Z(o[7560]) );
  AND U5424 ( .A(p_input[27560]), .B(p_input[17560]), .Z(n2712) );
  AND U5425 ( .A(n2713), .B(p_input[755]), .Z(o[755]) );
  AND U5426 ( .A(p_input[20755]), .B(p_input[10755]), .Z(n2713) );
  AND U5427 ( .A(n2714), .B(p_input[7559]), .Z(o[7559]) );
  AND U5428 ( .A(p_input[27559]), .B(p_input[17559]), .Z(n2714) );
  AND U5429 ( .A(n2715), .B(p_input[7558]), .Z(o[7558]) );
  AND U5430 ( .A(p_input[27558]), .B(p_input[17558]), .Z(n2715) );
  AND U5431 ( .A(n2716), .B(p_input[7557]), .Z(o[7557]) );
  AND U5432 ( .A(p_input[27557]), .B(p_input[17557]), .Z(n2716) );
  AND U5433 ( .A(n2717), .B(p_input[7556]), .Z(o[7556]) );
  AND U5434 ( .A(p_input[27556]), .B(p_input[17556]), .Z(n2717) );
  AND U5435 ( .A(n2718), .B(p_input[7555]), .Z(o[7555]) );
  AND U5436 ( .A(p_input[27555]), .B(p_input[17555]), .Z(n2718) );
  AND U5437 ( .A(n2719), .B(p_input[7554]), .Z(o[7554]) );
  AND U5438 ( .A(p_input[27554]), .B(p_input[17554]), .Z(n2719) );
  AND U5439 ( .A(n2720), .B(p_input[7553]), .Z(o[7553]) );
  AND U5440 ( .A(p_input[27553]), .B(p_input[17553]), .Z(n2720) );
  AND U5441 ( .A(n2721), .B(p_input[7552]), .Z(o[7552]) );
  AND U5442 ( .A(p_input[27552]), .B(p_input[17552]), .Z(n2721) );
  AND U5443 ( .A(n2722), .B(p_input[7551]), .Z(o[7551]) );
  AND U5444 ( .A(p_input[27551]), .B(p_input[17551]), .Z(n2722) );
  AND U5445 ( .A(n2723), .B(p_input[7550]), .Z(o[7550]) );
  AND U5446 ( .A(p_input[27550]), .B(p_input[17550]), .Z(n2723) );
  AND U5447 ( .A(n2724), .B(p_input[754]), .Z(o[754]) );
  AND U5448 ( .A(p_input[20754]), .B(p_input[10754]), .Z(n2724) );
  AND U5449 ( .A(n2725), .B(p_input[7549]), .Z(o[7549]) );
  AND U5450 ( .A(p_input[27549]), .B(p_input[17549]), .Z(n2725) );
  AND U5451 ( .A(n2726), .B(p_input[7548]), .Z(o[7548]) );
  AND U5452 ( .A(p_input[27548]), .B(p_input[17548]), .Z(n2726) );
  AND U5453 ( .A(n2727), .B(p_input[7547]), .Z(o[7547]) );
  AND U5454 ( .A(p_input[27547]), .B(p_input[17547]), .Z(n2727) );
  AND U5455 ( .A(n2728), .B(p_input[7546]), .Z(o[7546]) );
  AND U5456 ( .A(p_input[27546]), .B(p_input[17546]), .Z(n2728) );
  AND U5457 ( .A(n2729), .B(p_input[7545]), .Z(o[7545]) );
  AND U5458 ( .A(p_input[27545]), .B(p_input[17545]), .Z(n2729) );
  AND U5459 ( .A(n2730), .B(p_input[7544]), .Z(o[7544]) );
  AND U5460 ( .A(p_input[27544]), .B(p_input[17544]), .Z(n2730) );
  AND U5461 ( .A(n2731), .B(p_input[7543]), .Z(o[7543]) );
  AND U5462 ( .A(p_input[27543]), .B(p_input[17543]), .Z(n2731) );
  AND U5463 ( .A(n2732), .B(p_input[7542]), .Z(o[7542]) );
  AND U5464 ( .A(p_input[27542]), .B(p_input[17542]), .Z(n2732) );
  AND U5465 ( .A(n2733), .B(p_input[7541]), .Z(o[7541]) );
  AND U5466 ( .A(p_input[27541]), .B(p_input[17541]), .Z(n2733) );
  AND U5467 ( .A(n2734), .B(p_input[7540]), .Z(o[7540]) );
  AND U5468 ( .A(p_input[27540]), .B(p_input[17540]), .Z(n2734) );
  AND U5469 ( .A(n2735), .B(p_input[753]), .Z(o[753]) );
  AND U5470 ( .A(p_input[20753]), .B(p_input[10753]), .Z(n2735) );
  AND U5471 ( .A(n2736), .B(p_input[7539]), .Z(o[7539]) );
  AND U5472 ( .A(p_input[27539]), .B(p_input[17539]), .Z(n2736) );
  AND U5473 ( .A(n2737), .B(p_input[7538]), .Z(o[7538]) );
  AND U5474 ( .A(p_input[27538]), .B(p_input[17538]), .Z(n2737) );
  AND U5475 ( .A(n2738), .B(p_input[7537]), .Z(o[7537]) );
  AND U5476 ( .A(p_input[27537]), .B(p_input[17537]), .Z(n2738) );
  AND U5477 ( .A(n2739), .B(p_input[7536]), .Z(o[7536]) );
  AND U5478 ( .A(p_input[27536]), .B(p_input[17536]), .Z(n2739) );
  AND U5479 ( .A(n2740), .B(p_input[7535]), .Z(o[7535]) );
  AND U5480 ( .A(p_input[27535]), .B(p_input[17535]), .Z(n2740) );
  AND U5481 ( .A(n2741), .B(p_input[7534]), .Z(o[7534]) );
  AND U5482 ( .A(p_input[27534]), .B(p_input[17534]), .Z(n2741) );
  AND U5483 ( .A(n2742), .B(p_input[7533]), .Z(o[7533]) );
  AND U5484 ( .A(p_input[27533]), .B(p_input[17533]), .Z(n2742) );
  AND U5485 ( .A(n2743), .B(p_input[7532]), .Z(o[7532]) );
  AND U5486 ( .A(p_input[27532]), .B(p_input[17532]), .Z(n2743) );
  AND U5487 ( .A(n2744), .B(p_input[7531]), .Z(o[7531]) );
  AND U5488 ( .A(p_input[27531]), .B(p_input[17531]), .Z(n2744) );
  AND U5489 ( .A(n2745), .B(p_input[7530]), .Z(o[7530]) );
  AND U5490 ( .A(p_input[27530]), .B(p_input[17530]), .Z(n2745) );
  AND U5491 ( .A(n2746), .B(p_input[752]), .Z(o[752]) );
  AND U5492 ( .A(p_input[20752]), .B(p_input[10752]), .Z(n2746) );
  AND U5493 ( .A(n2747), .B(p_input[7529]), .Z(o[7529]) );
  AND U5494 ( .A(p_input[27529]), .B(p_input[17529]), .Z(n2747) );
  AND U5495 ( .A(n2748), .B(p_input[7528]), .Z(o[7528]) );
  AND U5496 ( .A(p_input[27528]), .B(p_input[17528]), .Z(n2748) );
  AND U5497 ( .A(n2749), .B(p_input[7527]), .Z(o[7527]) );
  AND U5498 ( .A(p_input[27527]), .B(p_input[17527]), .Z(n2749) );
  AND U5499 ( .A(n2750), .B(p_input[7526]), .Z(o[7526]) );
  AND U5500 ( .A(p_input[27526]), .B(p_input[17526]), .Z(n2750) );
  AND U5501 ( .A(n2751), .B(p_input[7525]), .Z(o[7525]) );
  AND U5502 ( .A(p_input[27525]), .B(p_input[17525]), .Z(n2751) );
  AND U5503 ( .A(n2752), .B(p_input[7524]), .Z(o[7524]) );
  AND U5504 ( .A(p_input[27524]), .B(p_input[17524]), .Z(n2752) );
  AND U5505 ( .A(n2753), .B(p_input[7523]), .Z(o[7523]) );
  AND U5506 ( .A(p_input[27523]), .B(p_input[17523]), .Z(n2753) );
  AND U5507 ( .A(n2754), .B(p_input[7522]), .Z(o[7522]) );
  AND U5508 ( .A(p_input[27522]), .B(p_input[17522]), .Z(n2754) );
  AND U5509 ( .A(n2755), .B(p_input[7521]), .Z(o[7521]) );
  AND U5510 ( .A(p_input[27521]), .B(p_input[17521]), .Z(n2755) );
  AND U5511 ( .A(n2756), .B(p_input[7520]), .Z(o[7520]) );
  AND U5512 ( .A(p_input[27520]), .B(p_input[17520]), .Z(n2756) );
  AND U5513 ( .A(n2757), .B(p_input[751]), .Z(o[751]) );
  AND U5514 ( .A(p_input[20751]), .B(p_input[10751]), .Z(n2757) );
  AND U5515 ( .A(n2758), .B(p_input[7519]), .Z(o[7519]) );
  AND U5516 ( .A(p_input[27519]), .B(p_input[17519]), .Z(n2758) );
  AND U5517 ( .A(n2759), .B(p_input[7518]), .Z(o[7518]) );
  AND U5518 ( .A(p_input[27518]), .B(p_input[17518]), .Z(n2759) );
  AND U5519 ( .A(n2760), .B(p_input[7517]), .Z(o[7517]) );
  AND U5520 ( .A(p_input[27517]), .B(p_input[17517]), .Z(n2760) );
  AND U5521 ( .A(n2761), .B(p_input[7516]), .Z(o[7516]) );
  AND U5522 ( .A(p_input[27516]), .B(p_input[17516]), .Z(n2761) );
  AND U5523 ( .A(n2762), .B(p_input[7515]), .Z(o[7515]) );
  AND U5524 ( .A(p_input[27515]), .B(p_input[17515]), .Z(n2762) );
  AND U5525 ( .A(n2763), .B(p_input[7514]), .Z(o[7514]) );
  AND U5526 ( .A(p_input[27514]), .B(p_input[17514]), .Z(n2763) );
  AND U5527 ( .A(n2764), .B(p_input[7513]), .Z(o[7513]) );
  AND U5528 ( .A(p_input[27513]), .B(p_input[17513]), .Z(n2764) );
  AND U5529 ( .A(n2765), .B(p_input[7512]), .Z(o[7512]) );
  AND U5530 ( .A(p_input[27512]), .B(p_input[17512]), .Z(n2765) );
  AND U5531 ( .A(n2766), .B(p_input[7511]), .Z(o[7511]) );
  AND U5532 ( .A(p_input[27511]), .B(p_input[17511]), .Z(n2766) );
  AND U5533 ( .A(n2767), .B(p_input[7510]), .Z(o[7510]) );
  AND U5534 ( .A(p_input[27510]), .B(p_input[17510]), .Z(n2767) );
  AND U5535 ( .A(n2768), .B(p_input[750]), .Z(o[750]) );
  AND U5536 ( .A(p_input[20750]), .B(p_input[10750]), .Z(n2768) );
  AND U5537 ( .A(n2769), .B(p_input[7509]), .Z(o[7509]) );
  AND U5538 ( .A(p_input[27509]), .B(p_input[17509]), .Z(n2769) );
  AND U5539 ( .A(n2770), .B(p_input[7508]), .Z(o[7508]) );
  AND U5540 ( .A(p_input[27508]), .B(p_input[17508]), .Z(n2770) );
  AND U5541 ( .A(n2771), .B(p_input[7507]), .Z(o[7507]) );
  AND U5542 ( .A(p_input[27507]), .B(p_input[17507]), .Z(n2771) );
  AND U5543 ( .A(n2772), .B(p_input[7506]), .Z(o[7506]) );
  AND U5544 ( .A(p_input[27506]), .B(p_input[17506]), .Z(n2772) );
  AND U5545 ( .A(n2773), .B(p_input[7505]), .Z(o[7505]) );
  AND U5546 ( .A(p_input[27505]), .B(p_input[17505]), .Z(n2773) );
  AND U5547 ( .A(n2774), .B(p_input[7504]), .Z(o[7504]) );
  AND U5548 ( .A(p_input[27504]), .B(p_input[17504]), .Z(n2774) );
  AND U5549 ( .A(n2775), .B(p_input[7503]), .Z(o[7503]) );
  AND U5550 ( .A(p_input[27503]), .B(p_input[17503]), .Z(n2775) );
  AND U5551 ( .A(n2776), .B(p_input[7502]), .Z(o[7502]) );
  AND U5552 ( .A(p_input[27502]), .B(p_input[17502]), .Z(n2776) );
  AND U5553 ( .A(n2777), .B(p_input[7501]), .Z(o[7501]) );
  AND U5554 ( .A(p_input[27501]), .B(p_input[17501]), .Z(n2777) );
  AND U5555 ( .A(n2778), .B(p_input[7500]), .Z(o[7500]) );
  AND U5556 ( .A(p_input[27500]), .B(p_input[17500]), .Z(n2778) );
  AND U5557 ( .A(n2779), .B(p_input[74]), .Z(o[74]) );
  AND U5558 ( .A(p_input[20074]), .B(p_input[10074]), .Z(n2779) );
  AND U5559 ( .A(n2780), .B(p_input[749]), .Z(o[749]) );
  AND U5560 ( .A(p_input[20749]), .B(p_input[10749]), .Z(n2780) );
  AND U5561 ( .A(n2781), .B(p_input[7499]), .Z(o[7499]) );
  AND U5562 ( .A(p_input[27499]), .B(p_input[17499]), .Z(n2781) );
  AND U5563 ( .A(n2782), .B(p_input[7498]), .Z(o[7498]) );
  AND U5564 ( .A(p_input[27498]), .B(p_input[17498]), .Z(n2782) );
  AND U5565 ( .A(n2783), .B(p_input[7497]), .Z(o[7497]) );
  AND U5566 ( .A(p_input[27497]), .B(p_input[17497]), .Z(n2783) );
  AND U5567 ( .A(n2784), .B(p_input[7496]), .Z(o[7496]) );
  AND U5568 ( .A(p_input[27496]), .B(p_input[17496]), .Z(n2784) );
  AND U5569 ( .A(n2785), .B(p_input[7495]), .Z(o[7495]) );
  AND U5570 ( .A(p_input[27495]), .B(p_input[17495]), .Z(n2785) );
  AND U5571 ( .A(n2786), .B(p_input[7494]), .Z(o[7494]) );
  AND U5572 ( .A(p_input[27494]), .B(p_input[17494]), .Z(n2786) );
  AND U5573 ( .A(n2787), .B(p_input[7493]), .Z(o[7493]) );
  AND U5574 ( .A(p_input[27493]), .B(p_input[17493]), .Z(n2787) );
  AND U5575 ( .A(n2788), .B(p_input[7492]), .Z(o[7492]) );
  AND U5576 ( .A(p_input[27492]), .B(p_input[17492]), .Z(n2788) );
  AND U5577 ( .A(n2789), .B(p_input[7491]), .Z(o[7491]) );
  AND U5578 ( .A(p_input[27491]), .B(p_input[17491]), .Z(n2789) );
  AND U5579 ( .A(n2790), .B(p_input[7490]), .Z(o[7490]) );
  AND U5580 ( .A(p_input[27490]), .B(p_input[17490]), .Z(n2790) );
  AND U5581 ( .A(n2791), .B(p_input[748]), .Z(o[748]) );
  AND U5582 ( .A(p_input[20748]), .B(p_input[10748]), .Z(n2791) );
  AND U5583 ( .A(n2792), .B(p_input[7489]), .Z(o[7489]) );
  AND U5584 ( .A(p_input[27489]), .B(p_input[17489]), .Z(n2792) );
  AND U5585 ( .A(n2793), .B(p_input[7488]), .Z(o[7488]) );
  AND U5586 ( .A(p_input[27488]), .B(p_input[17488]), .Z(n2793) );
  AND U5587 ( .A(n2794), .B(p_input[7487]), .Z(o[7487]) );
  AND U5588 ( .A(p_input[27487]), .B(p_input[17487]), .Z(n2794) );
  AND U5589 ( .A(n2795), .B(p_input[7486]), .Z(o[7486]) );
  AND U5590 ( .A(p_input[27486]), .B(p_input[17486]), .Z(n2795) );
  AND U5591 ( .A(n2796), .B(p_input[7485]), .Z(o[7485]) );
  AND U5592 ( .A(p_input[27485]), .B(p_input[17485]), .Z(n2796) );
  AND U5593 ( .A(n2797), .B(p_input[7484]), .Z(o[7484]) );
  AND U5594 ( .A(p_input[27484]), .B(p_input[17484]), .Z(n2797) );
  AND U5595 ( .A(n2798), .B(p_input[7483]), .Z(o[7483]) );
  AND U5596 ( .A(p_input[27483]), .B(p_input[17483]), .Z(n2798) );
  AND U5597 ( .A(n2799), .B(p_input[7482]), .Z(o[7482]) );
  AND U5598 ( .A(p_input[27482]), .B(p_input[17482]), .Z(n2799) );
  AND U5599 ( .A(n2800), .B(p_input[7481]), .Z(o[7481]) );
  AND U5600 ( .A(p_input[27481]), .B(p_input[17481]), .Z(n2800) );
  AND U5601 ( .A(n2801), .B(p_input[7480]), .Z(o[7480]) );
  AND U5602 ( .A(p_input[27480]), .B(p_input[17480]), .Z(n2801) );
  AND U5603 ( .A(n2802), .B(p_input[747]), .Z(o[747]) );
  AND U5604 ( .A(p_input[20747]), .B(p_input[10747]), .Z(n2802) );
  AND U5605 ( .A(n2803), .B(p_input[7479]), .Z(o[7479]) );
  AND U5606 ( .A(p_input[27479]), .B(p_input[17479]), .Z(n2803) );
  AND U5607 ( .A(n2804), .B(p_input[7478]), .Z(o[7478]) );
  AND U5608 ( .A(p_input[27478]), .B(p_input[17478]), .Z(n2804) );
  AND U5609 ( .A(n2805), .B(p_input[7477]), .Z(o[7477]) );
  AND U5610 ( .A(p_input[27477]), .B(p_input[17477]), .Z(n2805) );
  AND U5611 ( .A(n2806), .B(p_input[7476]), .Z(o[7476]) );
  AND U5612 ( .A(p_input[27476]), .B(p_input[17476]), .Z(n2806) );
  AND U5613 ( .A(n2807), .B(p_input[7475]), .Z(o[7475]) );
  AND U5614 ( .A(p_input[27475]), .B(p_input[17475]), .Z(n2807) );
  AND U5615 ( .A(n2808), .B(p_input[7474]), .Z(o[7474]) );
  AND U5616 ( .A(p_input[27474]), .B(p_input[17474]), .Z(n2808) );
  AND U5617 ( .A(n2809), .B(p_input[7473]), .Z(o[7473]) );
  AND U5618 ( .A(p_input[27473]), .B(p_input[17473]), .Z(n2809) );
  AND U5619 ( .A(n2810), .B(p_input[7472]), .Z(o[7472]) );
  AND U5620 ( .A(p_input[27472]), .B(p_input[17472]), .Z(n2810) );
  AND U5621 ( .A(n2811), .B(p_input[7471]), .Z(o[7471]) );
  AND U5622 ( .A(p_input[27471]), .B(p_input[17471]), .Z(n2811) );
  AND U5623 ( .A(n2812), .B(p_input[7470]), .Z(o[7470]) );
  AND U5624 ( .A(p_input[27470]), .B(p_input[17470]), .Z(n2812) );
  AND U5625 ( .A(n2813), .B(p_input[746]), .Z(o[746]) );
  AND U5626 ( .A(p_input[20746]), .B(p_input[10746]), .Z(n2813) );
  AND U5627 ( .A(n2814), .B(p_input[7469]), .Z(o[7469]) );
  AND U5628 ( .A(p_input[27469]), .B(p_input[17469]), .Z(n2814) );
  AND U5629 ( .A(n2815), .B(p_input[7468]), .Z(o[7468]) );
  AND U5630 ( .A(p_input[27468]), .B(p_input[17468]), .Z(n2815) );
  AND U5631 ( .A(n2816), .B(p_input[7467]), .Z(o[7467]) );
  AND U5632 ( .A(p_input[27467]), .B(p_input[17467]), .Z(n2816) );
  AND U5633 ( .A(n2817), .B(p_input[7466]), .Z(o[7466]) );
  AND U5634 ( .A(p_input[27466]), .B(p_input[17466]), .Z(n2817) );
  AND U5635 ( .A(n2818), .B(p_input[7465]), .Z(o[7465]) );
  AND U5636 ( .A(p_input[27465]), .B(p_input[17465]), .Z(n2818) );
  AND U5637 ( .A(n2819), .B(p_input[7464]), .Z(o[7464]) );
  AND U5638 ( .A(p_input[27464]), .B(p_input[17464]), .Z(n2819) );
  AND U5639 ( .A(n2820), .B(p_input[7463]), .Z(o[7463]) );
  AND U5640 ( .A(p_input[27463]), .B(p_input[17463]), .Z(n2820) );
  AND U5641 ( .A(n2821), .B(p_input[7462]), .Z(o[7462]) );
  AND U5642 ( .A(p_input[27462]), .B(p_input[17462]), .Z(n2821) );
  AND U5643 ( .A(n2822), .B(p_input[7461]), .Z(o[7461]) );
  AND U5644 ( .A(p_input[27461]), .B(p_input[17461]), .Z(n2822) );
  AND U5645 ( .A(n2823), .B(p_input[7460]), .Z(o[7460]) );
  AND U5646 ( .A(p_input[27460]), .B(p_input[17460]), .Z(n2823) );
  AND U5647 ( .A(n2824), .B(p_input[745]), .Z(o[745]) );
  AND U5648 ( .A(p_input[20745]), .B(p_input[10745]), .Z(n2824) );
  AND U5649 ( .A(n2825), .B(p_input[7459]), .Z(o[7459]) );
  AND U5650 ( .A(p_input[27459]), .B(p_input[17459]), .Z(n2825) );
  AND U5651 ( .A(n2826), .B(p_input[7458]), .Z(o[7458]) );
  AND U5652 ( .A(p_input[27458]), .B(p_input[17458]), .Z(n2826) );
  AND U5653 ( .A(n2827), .B(p_input[7457]), .Z(o[7457]) );
  AND U5654 ( .A(p_input[27457]), .B(p_input[17457]), .Z(n2827) );
  AND U5655 ( .A(n2828), .B(p_input[7456]), .Z(o[7456]) );
  AND U5656 ( .A(p_input[27456]), .B(p_input[17456]), .Z(n2828) );
  AND U5657 ( .A(n2829), .B(p_input[7455]), .Z(o[7455]) );
  AND U5658 ( .A(p_input[27455]), .B(p_input[17455]), .Z(n2829) );
  AND U5659 ( .A(n2830), .B(p_input[7454]), .Z(o[7454]) );
  AND U5660 ( .A(p_input[27454]), .B(p_input[17454]), .Z(n2830) );
  AND U5661 ( .A(n2831), .B(p_input[7453]), .Z(o[7453]) );
  AND U5662 ( .A(p_input[27453]), .B(p_input[17453]), .Z(n2831) );
  AND U5663 ( .A(n2832), .B(p_input[7452]), .Z(o[7452]) );
  AND U5664 ( .A(p_input[27452]), .B(p_input[17452]), .Z(n2832) );
  AND U5665 ( .A(n2833), .B(p_input[7451]), .Z(o[7451]) );
  AND U5666 ( .A(p_input[27451]), .B(p_input[17451]), .Z(n2833) );
  AND U5667 ( .A(n2834), .B(p_input[7450]), .Z(o[7450]) );
  AND U5668 ( .A(p_input[27450]), .B(p_input[17450]), .Z(n2834) );
  AND U5669 ( .A(n2835), .B(p_input[744]), .Z(o[744]) );
  AND U5670 ( .A(p_input[20744]), .B(p_input[10744]), .Z(n2835) );
  AND U5671 ( .A(n2836), .B(p_input[7449]), .Z(o[7449]) );
  AND U5672 ( .A(p_input[27449]), .B(p_input[17449]), .Z(n2836) );
  AND U5673 ( .A(n2837), .B(p_input[7448]), .Z(o[7448]) );
  AND U5674 ( .A(p_input[27448]), .B(p_input[17448]), .Z(n2837) );
  AND U5675 ( .A(n2838), .B(p_input[7447]), .Z(o[7447]) );
  AND U5676 ( .A(p_input[27447]), .B(p_input[17447]), .Z(n2838) );
  AND U5677 ( .A(n2839), .B(p_input[7446]), .Z(o[7446]) );
  AND U5678 ( .A(p_input[27446]), .B(p_input[17446]), .Z(n2839) );
  AND U5679 ( .A(n2840), .B(p_input[7445]), .Z(o[7445]) );
  AND U5680 ( .A(p_input[27445]), .B(p_input[17445]), .Z(n2840) );
  AND U5681 ( .A(n2841), .B(p_input[7444]), .Z(o[7444]) );
  AND U5682 ( .A(p_input[27444]), .B(p_input[17444]), .Z(n2841) );
  AND U5683 ( .A(n2842), .B(p_input[7443]), .Z(o[7443]) );
  AND U5684 ( .A(p_input[27443]), .B(p_input[17443]), .Z(n2842) );
  AND U5685 ( .A(n2843), .B(p_input[7442]), .Z(o[7442]) );
  AND U5686 ( .A(p_input[27442]), .B(p_input[17442]), .Z(n2843) );
  AND U5687 ( .A(n2844), .B(p_input[7441]), .Z(o[7441]) );
  AND U5688 ( .A(p_input[27441]), .B(p_input[17441]), .Z(n2844) );
  AND U5689 ( .A(n2845), .B(p_input[7440]), .Z(o[7440]) );
  AND U5690 ( .A(p_input[27440]), .B(p_input[17440]), .Z(n2845) );
  AND U5691 ( .A(n2846), .B(p_input[743]), .Z(o[743]) );
  AND U5692 ( .A(p_input[20743]), .B(p_input[10743]), .Z(n2846) );
  AND U5693 ( .A(n2847), .B(p_input[7439]), .Z(o[7439]) );
  AND U5694 ( .A(p_input[27439]), .B(p_input[17439]), .Z(n2847) );
  AND U5695 ( .A(n2848), .B(p_input[7438]), .Z(o[7438]) );
  AND U5696 ( .A(p_input[27438]), .B(p_input[17438]), .Z(n2848) );
  AND U5697 ( .A(n2849), .B(p_input[7437]), .Z(o[7437]) );
  AND U5698 ( .A(p_input[27437]), .B(p_input[17437]), .Z(n2849) );
  AND U5699 ( .A(n2850), .B(p_input[7436]), .Z(o[7436]) );
  AND U5700 ( .A(p_input[27436]), .B(p_input[17436]), .Z(n2850) );
  AND U5701 ( .A(n2851), .B(p_input[7435]), .Z(o[7435]) );
  AND U5702 ( .A(p_input[27435]), .B(p_input[17435]), .Z(n2851) );
  AND U5703 ( .A(n2852), .B(p_input[7434]), .Z(o[7434]) );
  AND U5704 ( .A(p_input[27434]), .B(p_input[17434]), .Z(n2852) );
  AND U5705 ( .A(n2853), .B(p_input[7433]), .Z(o[7433]) );
  AND U5706 ( .A(p_input[27433]), .B(p_input[17433]), .Z(n2853) );
  AND U5707 ( .A(n2854), .B(p_input[7432]), .Z(o[7432]) );
  AND U5708 ( .A(p_input[27432]), .B(p_input[17432]), .Z(n2854) );
  AND U5709 ( .A(n2855), .B(p_input[7431]), .Z(o[7431]) );
  AND U5710 ( .A(p_input[27431]), .B(p_input[17431]), .Z(n2855) );
  AND U5711 ( .A(n2856), .B(p_input[7430]), .Z(o[7430]) );
  AND U5712 ( .A(p_input[27430]), .B(p_input[17430]), .Z(n2856) );
  AND U5713 ( .A(n2857), .B(p_input[742]), .Z(o[742]) );
  AND U5714 ( .A(p_input[20742]), .B(p_input[10742]), .Z(n2857) );
  AND U5715 ( .A(n2858), .B(p_input[7429]), .Z(o[7429]) );
  AND U5716 ( .A(p_input[27429]), .B(p_input[17429]), .Z(n2858) );
  AND U5717 ( .A(n2859), .B(p_input[7428]), .Z(o[7428]) );
  AND U5718 ( .A(p_input[27428]), .B(p_input[17428]), .Z(n2859) );
  AND U5719 ( .A(n2860), .B(p_input[7427]), .Z(o[7427]) );
  AND U5720 ( .A(p_input[27427]), .B(p_input[17427]), .Z(n2860) );
  AND U5721 ( .A(n2861), .B(p_input[7426]), .Z(o[7426]) );
  AND U5722 ( .A(p_input[27426]), .B(p_input[17426]), .Z(n2861) );
  AND U5723 ( .A(n2862), .B(p_input[7425]), .Z(o[7425]) );
  AND U5724 ( .A(p_input[27425]), .B(p_input[17425]), .Z(n2862) );
  AND U5725 ( .A(n2863), .B(p_input[7424]), .Z(o[7424]) );
  AND U5726 ( .A(p_input[27424]), .B(p_input[17424]), .Z(n2863) );
  AND U5727 ( .A(n2864), .B(p_input[7423]), .Z(o[7423]) );
  AND U5728 ( .A(p_input[27423]), .B(p_input[17423]), .Z(n2864) );
  AND U5729 ( .A(n2865), .B(p_input[7422]), .Z(o[7422]) );
  AND U5730 ( .A(p_input[27422]), .B(p_input[17422]), .Z(n2865) );
  AND U5731 ( .A(n2866), .B(p_input[7421]), .Z(o[7421]) );
  AND U5732 ( .A(p_input[27421]), .B(p_input[17421]), .Z(n2866) );
  AND U5733 ( .A(n2867), .B(p_input[7420]), .Z(o[7420]) );
  AND U5734 ( .A(p_input[27420]), .B(p_input[17420]), .Z(n2867) );
  AND U5735 ( .A(n2868), .B(p_input[741]), .Z(o[741]) );
  AND U5736 ( .A(p_input[20741]), .B(p_input[10741]), .Z(n2868) );
  AND U5737 ( .A(n2869), .B(p_input[7419]), .Z(o[7419]) );
  AND U5738 ( .A(p_input[27419]), .B(p_input[17419]), .Z(n2869) );
  AND U5739 ( .A(n2870), .B(p_input[7418]), .Z(o[7418]) );
  AND U5740 ( .A(p_input[27418]), .B(p_input[17418]), .Z(n2870) );
  AND U5741 ( .A(n2871), .B(p_input[7417]), .Z(o[7417]) );
  AND U5742 ( .A(p_input[27417]), .B(p_input[17417]), .Z(n2871) );
  AND U5743 ( .A(n2872), .B(p_input[7416]), .Z(o[7416]) );
  AND U5744 ( .A(p_input[27416]), .B(p_input[17416]), .Z(n2872) );
  AND U5745 ( .A(n2873), .B(p_input[7415]), .Z(o[7415]) );
  AND U5746 ( .A(p_input[27415]), .B(p_input[17415]), .Z(n2873) );
  AND U5747 ( .A(n2874), .B(p_input[7414]), .Z(o[7414]) );
  AND U5748 ( .A(p_input[27414]), .B(p_input[17414]), .Z(n2874) );
  AND U5749 ( .A(n2875), .B(p_input[7413]), .Z(o[7413]) );
  AND U5750 ( .A(p_input[27413]), .B(p_input[17413]), .Z(n2875) );
  AND U5751 ( .A(n2876), .B(p_input[7412]), .Z(o[7412]) );
  AND U5752 ( .A(p_input[27412]), .B(p_input[17412]), .Z(n2876) );
  AND U5753 ( .A(n2877), .B(p_input[7411]), .Z(o[7411]) );
  AND U5754 ( .A(p_input[27411]), .B(p_input[17411]), .Z(n2877) );
  AND U5755 ( .A(n2878), .B(p_input[7410]), .Z(o[7410]) );
  AND U5756 ( .A(p_input[27410]), .B(p_input[17410]), .Z(n2878) );
  AND U5757 ( .A(n2879), .B(p_input[740]), .Z(o[740]) );
  AND U5758 ( .A(p_input[20740]), .B(p_input[10740]), .Z(n2879) );
  AND U5759 ( .A(n2880), .B(p_input[7409]), .Z(o[7409]) );
  AND U5760 ( .A(p_input[27409]), .B(p_input[17409]), .Z(n2880) );
  AND U5761 ( .A(n2881), .B(p_input[7408]), .Z(o[7408]) );
  AND U5762 ( .A(p_input[27408]), .B(p_input[17408]), .Z(n2881) );
  AND U5763 ( .A(n2882), .B(p_input[7407]), .Z(o[7407]) );
  AND U5764 ( .A(p_input[27407]), .B(p_input[17407]), .Z(n2882) );
  AND U5765 ( .A(n2883), .B(p_input[7406]), .Z(o[7406]) );
  AND U5766 ( .A(p_input[27406]), .B(p_input[17406]), .Z(n2883) );
  AND U5767 ( .A(n2884), .B(p_input[7405]), .Z(o[7405]) );
  AND U5768 ( .A(p_input[27405]), .B(p_input[17405]), .Z(n2884) );
  AND U5769 ( .A(n2885), .B(p_input[7404]), .Z(o[7404]) );
  AND U5770 ( .A(p_input[27404]), .B(p_input[17404]), .Z(n2885) );
  AND U5771 ( .A(n2886), .B(p_input[7403]), .Z(o[7403]) );
  AND U5772 ( .A(p_input[27403]), .B(p_input[17403]), .Z(n2886) );
  AND U5773 ( .A(n2887), .B(p_input[7402]), .Z(o[7402]) );
  AND U5774 ( .A(p_input[27402]), .B(p_input[17402]), .Z(n2887) );
  AND U5775 ( .A(n2888), .B(p_input[7401]), .Z(o[7401]) );
  AND U5776 ( .A(p_input[27401]), .B(p_input[17401]), .Z(n2888) );
  AND U5777 ( .A(n2889), .B(p_input[7400]), .Z(o[7400]) );
  AND U5778 ( .A(p_input[27400]), .B(p_input[17400]), .Z(n2889) );
  AND U5779 ( .A(n2890), .B(p_input[73]), .Z(o[73]) );
  AND U5780 ( .A(p_input[20073]), .B(p_input[10073]), .Z(n2890) );
  AND U5781 ( .A(n2891), .B(p_input[739]), .Z(o[739]) );
  AND U5782 ( .A(p_input[20739]), .B(p_input[10739]), .Z(n2891) );
  AND U5783 ( .A(n2892), .B(p_input[7399]), .Z(o[7399]) );
  AND U5784 ( .A(p_input[27399]), .B(p_input[17399]), .Z(n2892) );
  AND U5785 ( .A(n2893), .B(p_input[7398]), .Z(o[7398]) );
  AND U5786 ( .A(p_input[27398]), .B(p_input[17398]), .Z(n2893) );
  AND U5787 ( .A(n2894), .B(p_input[7397]), .Z(o[7397]) );
  AND U5788 ( .A(p_input[27397]), .B(p_input[17397]), .Z(n2894) );
  AND U5789 ( .A(n2895), .B(p_input[7396]), .Z(o[7396]) );
  AND U5790 ( .A(p_input[27396]), .B(p_input[17396]), .Z(n2895) );
  AND U5791 ( .A(n2896), .B(p_input[7395]), .Z(o[7395]) );
  AND U5792 ( .A(p_input[27395]), .B(p_input[17395]), .Z(n2896) );
  AND U5793 ( .A(n2897), .B(p_input[7394]), .Z(o[7394]) );
  AND U5794 ( .A(p_input[27394]), .B(p_input[17394]), .Z(n2897) );
  AND U5795 ( .A(n2898), .B(p_input[7393]), .Z(o[7393]) );
  AND U5796 ( .A(p_input[27393]), .B(p_input[17393]), .Z(n2898) );
  AND U5797 ( .A(n2899), .B(p_input[7392]), .Z(o[7392]) );
  AND U5798 ( .A(p_input[27392]), .B(p_input[17392]), .Z(n2899) );
  AND U5799 ( .A(n2900), .B(p_input[7391]), .Z(o[7391]) );
  AND U5800 ( .A(p_input[27391]), .B(p_input[17391]), .Z(n2900) );
  AND U5801 ( .A(n2901), .B(p_input[7390]), .Z(o[7390]) );
  AND U5802 ( .A(p_input[27390]), .B(p_input[17390]), .Z(n2901) );
  AND U5803 ( .A(n2902), .B(p_input[738]), .Z(o[738]) );
  AND U5804 ( .A(p_input[20738]), .B(p_input[10738]), .Z(n2902) );
  AND U5805 ( .A(n2903), .B(p_input[7389]), .Z(o[7389]) );
  AND U5806 ( .A(p_input[27389]), .B(p_input[17389]), .Z(n2903) );
  AND U5807 ( .A(n2904), .B(p_input[7388]), .Z(o[7388]) );
  AND U5808 ( .A(p_input[27388]), .B(p_input[17388]), .Z(n2904) );
  AND U5809 ( .A(n2905), .B(p_input[7387]), .Z(o[7387]) );
  AND U5810 ( .A(p_input[27387]), .B(p_input[17387]), .Z(n2905) );
  AND U5811 ( .A(n2906), .B(p_input[7386]), .Z(o[7386]) );
  AND U5812 ( .A(p_input[27386]), .B(p_input[17386]), .Z(n2906) );
  AND U5813 ( .A(n2907), .B(p_input[7385]), .Z(o[7385]) );
  AND U5814 ( .A(p_input[27385]), .B(p_input[17385]), .Z(n2907) );
  AND U5815 ( .A(n2908), .B(p_input[7384]), .Z(o[7384]) );
  AND U5816 ( .A(p_input[27384]), .B(p_input[17384]), .Z(n2908) );
  AND U5817 ( .A(n2909), .B(p_input[7383]), .Z(o[7383]) );
  AND U5818 ( .A(p_input[27383]), .B(p_input[17383]), .Z(n2909) );
  AND U5819 ( .A(n2910), .B(p_input[7382]), .Z(o[7382]) );
  AND U5820 ( .A(p_input[27382]), .B(p_input[17382]), .Z(n2910) );
  AND U5821 ( .A(n2911), .B(p_input[7381]), .Z(o[7381]) );
  AND U5822 ( .A(p_input[27381]), .B(p_input[17381]), .Z(n2911) );
  AND U5823 ( .A(n2912), .B(p_input[7380]), .Z(o[7380]) );
  AND U5824 ( .A(p_input[27380]), .B(p_input[17380]), .Z(n2912) );
  AND U5825 ( .A(n2913), .B(p_input[737]), .Z(o[737]) );
  AND U5826 ( .A(p_input[20737]), .B(p_input[10737]), .Z(n2913) );
  AND U5827 ( .A(n2914), .B(p_input[7379]), .Z(o[7379]) );
  AND U5828 ( .A(p_input[27379]), .B(p_input[17379]), .Z(n2914) );
  AND U5829 ( .A(n2915), .B(p_input[7378]), .Z(o[7378]) );
  AND U5830 ( .A(p_input[27378]), .B(p_input[17378]), .Z(n2915) );
  AND U5831 ( .A(n2916), .B(p_input[7377]), .Z(o[7377]) );
  AND U5832 ( .A(p_input[27377]), .B(p_input[17377]), .Z(n2916) );
  AND U5833 ( .A(n2917), .B(p_input[7376]), .Z(o[7376]) );
  AND U5834 ( .A(p_input[27376]), .B(p_input[17376]), .Z(n2917) );
  AND U5835 ( .A(n2918), .B(p_input[7375]), .Z(o[7375]) );
  AND U5836 ( .A(p_input[27375]), .B(p_input[17375]), .Z(n2918) );
  AND U5837 ( .A(n2919), .B(p_input[7374]), .Z(o[7374]) );
  AND U5838 ( .A(p_input[27374]), .B(p_input[17374]), .Z(n2919) );
  AND U5839 ( .A(n2920), .B(p_input[7373]), .Z(o[7373]) );
  AND U5840 ( .A(p_input[27373]), .B(p_input[17373]), .Z(n2920) );
  AND U5841 ( .A(n2921), .B(p_input[7372]), .Z(o[7372]) );
  AND U5842 ( .A(p_input[27372]), .B(p_input[17372]), .Z(n2921) );
  AND U5843 ( .A(n2922), .B(p_input[7371]), .Z(o[7371]) );
  AND U5844 ( .A(p_input[27371]), .B(p_input[17371]), .Z(n2922) );
  AND U5845 ( .A(n2923), .B(p_input[7370]), .Z(o[7370]) );
  AND U5846 ( .A(p_input[27370]), .B(p_input[17370]), .Z(n2923) );
  AND U5847 ( .A(n2924), .B(p_input[736]), .Z(o[736]) );
  AND U5848 ( .A(p_input[20736]), .B(p_input[10736]), .Z(n2924) );
  AND U5849 ( .A(n2925), .B(p_input[7369]), .Z(o[7369]) );
  AND U5850 ( .A(p_input[27369]), .B(p_input[17369]), .Z(n2925) );
  AND U5851 ( .A(n2926), .B(p_input[7368]), .Z(o[7368]) );
  AND U5852 ( .A(p_input[27368]), .B(p_input[17368]), .Z(n2926) );
  AND U5853 ( .A(n2927), .B(p_input[7367]), .Z(o[7367]) );
  AND U5854 ( .A(p_input[27367]), .B(p_input[17367]), .Z(n2927) );
  AND U5855 ( .A(n2928), .B(p_input[7366]), .Z(o[7366]) );
  AND U5856 ( .A(p_input[27366]), .B(p_input[17366]), .Z(n2928) );
  AND U5857 ( .A(n2929), .B(p_input[7365]), .Z(o[7365]) );
  AND U5858 ( .A(p_input[27365]), .B(p_input[17365]), .Z(n2929) );
  AND U5859 ( .A(n2930), .B(p_input[7364]), .Z(o[7364]) );
  AND U5860 ( .A(p_input[27364]), .B(p_input[17364]), .Z(n2930) );
  AND U5861 ( .A(n2931), .B(p_input[7363]), .Z(o[7363]) );
  AND U5862 ( .A(p_input[27363]), .B(p_input[17363]), .Z(n2931) );
  AND U5863 ( .A(n2932), .B(p_input[7362]), .Z(o[7362]) );
  AND U5864 ( .A(p_input[27362]), .B(p_input[17362]), .Z(n2932) );
  AND U5865 ( .A(n2933), .B(p_input[7361]), .Z(o[7361]) );
  AND U5866 ( .A(p_input[27361]), .B(p_input[17361]), .Z(n2933) );
  AND U5867 ( .A(n2934), .B(p_input[7360]), .Z(o[7360]) );
  AND U5868 ( .A(p_input[27360]), .B(p_input[17360]), .Z(n2934) );
  AND U5869 ( .A(n2935), .B(p_input[735]), .Z(o[735]) );
  AND U5870 ( .A(p_input[20735]), .B(p_input[10735]), .Z(n2935) );
  AND U5871 ( .A(n2936), .B(p_input[7359]), .Z(o[7359]) );
  AND U5872 ( .A(p_input[27359]), .B(p_input[17359]), .Z(n2936) );
  AND U5873 ( .A(n2937), .B(p_input[7358]), .Z(o[7358]) );
  AND U5874 ( .A(p_input[27358]), .B(p_input[17358]), .Z(n2937) );
  AND U5875 ( .A(n2938), .B(p_input[7357]), .Z(o[7357]) );
  AND U5876 ( .A(p_input[27357]), .B(p_input[17357]), .Z(n2938) );
  AND U5877 ( .A(n2939), .B(p_input[7356]), .Z(o[7356]) );
  AND U5878 ( .A(p_input[27356]), .B(p_input[17356]), .Z(n2939) );
  AND U5879 ( .A(n2940), .B(p_input[7355]), .Z(o[7355]) );
  AND U5880 ( .A(p_input[27355]), .B(p_input[17355]), .Z(n2940) );
  AND U5881 ( .A(n2941), .B(p_input[7354]), .Z(o[7354]) );
  AND U5882 ( .A(p_input[27354]), .B(p_input[17354]), .Z(n2941) );
  AND U5883 ( .A(n2942), .B(p_input[7353]), .Z(o[7353]) );
  AND U5884 ( .A(p_input[27353]), .B(p_input[17353]), .Z(n2942) );
  AND U5885 ( .A(n2943), .B(p_input[7352]), .Z(o[7352]) );
  AND U5886 ( .A(p_input[27352]), .B(p_input[17352]), .Z(n2943) );
  AND U5887 ( .A(n2944), .B(p_input[7351]), .Z(o[7351]) );
  AND U5888 ( .A(p_input[27351]), .B(p_input[17351]), .Z(n2944) );
  AND U5889 ( .A(n2945), .B(p_input[7350]), .Z(o[7350]) );
  AND U5890 ( .A(p_input[27350]), .B(p_input[17350]), .Z(n2945) );
  AND U5891 ( .A(n2946), .B(p_input[734]), .Z(o[734]) );
  AND U5892 ( .A(p_input[20734]), .B(p_input[10734]), .Z(n2946) );
  AND U5893 ( .A(n2947), .B(p_input[7349]), .Z(o[7349]) );
  AND U5894 ( .A(p_input[27349]), .B(p_input[17349]), .Z(n2947) );
  AND U5895 ( .A(n2948), .B(p_input[7348]), .Z(o[7348]) );
  AND U5896 ( .A(p_input[27348]), .B(p_input[17348]), .Z(n2948) );
  AND U5897 ( .A(n2949), .B(p_input[7347]), .Z(o[7347]) );
  AND U5898 ( .A(p_input[27347]), .B(p_input[17347]), .Z(n2949) );
  AND U5899 ( .A(n2950), .B(p_input[7346]), .Z(o[7346]) );
  AND U5900 ( .A(p_input[27346]), .B(p_input[17346]), .Z(n2950) );
  AND U5901 ( .A(n2951), .B(p_input[7345]), .Z(o[7345]) );
  AND U5902 ( .A(p_input[27345]), .B(p_input[17345]), .Z(n2951) );
  AND U5903 ( .A(n2952), .B(p_input[7344]), .Z(o[7344]) );
  AND U5904 ( .A(p_input[27344]), .B(p_input[17344]), .Z(n2952) );
  AND U5905 ( .A(n2953), .B(p_input[7343]), .Z(o[7343]) );
  AND U5906 ( .A(p_input[27343]), .B(p_input[17343]), .Z(n2953) );
  AND U5907 ( .A(n2954), .B(p_input[7342]), .Z(o[7342]) );
  AND U5908 ( .A(p_input[27342]), .B(p_input[17342]), .Z(n2954) );
  AND U5909 ( .A(n2955), .B(p_input[7341]), .Z(o[7341]) );
  AND U5910 ( .A(p_input[27341]), .B(p_input[17341]), .Z(n2955) );
  AND U5911 ( .A(n2956), .B(p_input[7340]), .Z(o[7340]) );
  AND U5912 ( .A(p_input[27340]), .B(p_input[17340]), .Z(n2956) );
  AND U5913 ( .A(n2957), .B(p_input[733]), .Z(o[733]) );
  AND U5914 ( .A(p_input[20733]), .B(p_input[10733]), .Z(n2957) );
  AND U5915 ( .A(n2958), .B(p_input[7339]), .Z(o[7339]) );
  AND U5916 ( .A(p_input[27339]), .B(p_input[17339]), .Z(n2958) );
  AND U5917 ( .A(n2959), .B(p_input[7338]), .Z(o[7338]) );
  AND U5918 ( .A(p_input[27338]), .B(p_input[17338]), .Z(n2959) );
  AND U5919 ( .A(n2960), .B(p_input[7337]), .Z(o[7337]) );
  AND U5920 ( .A(p_input[27337]), .B(p_input[17337]), .Z(n2960) );
  AND U5921 ( .A(n2961), .B(p_input[7336]), .Z(o[7336]) );
  AND U5922 ( .A(p_input[27336]), .B(p_input[17336]), .Z(n2961) );
  AND U5923 ( .A(n2962), .B(p_input[7335]), .Z(o[7335]) );
  AND U5924 ( .A(p_input[27335]), .B(p_input[17335]), .Z(n2962) );
  AND U5925 ( .A(n2963), .B(p_input[7334]), .Z(o[7334]) );
  AND U5926 ( .A(p_input[27334]), .B(p_input[17334]), .Z(n2963) );
  AND U5927 ( .A(n2964), .B(p_input[7333]), .Z(o[7333]) );
  AND U5928 ( .A(p_input[27333]), .B(p_input[17333]), .Z(n2964) );
  AND U5929 ( .A(n2965), .B(p_input[7332]), .Z(o[7332]) );
  AND U5930 ( .A(p_input[27332]), .B(p_input[17332]), .Z(n2965) );
  AND U5931 ( .A(n2966), .B(p_input[7331]), .Z(o[7331]) );
  AND U5932 ( .A(p_input[27331]), .B(p_input[17331]), .Z(n2966) );
  AND U5933 ( .A(n2967), .B(p_input[7330]), .Z(o[7330]) );
  AND U5934 ( .A(p_input[27330]), .B(p_input[17330]), .Z(n2967) );
  AND U5935 ( .A(n2968), .B(p_input[732]), .Z(o[732]) );
  AND U5936 ( .A(p_input[20732]), .B(p_input[10732]), .Z(n2968) );
  AND U5937 ( .A(n2969), .B(p_input[7329]), .Z(o[7329]) );
  AND U5938 ( .A(p_input[27329]), .B(p_input[17329]), .Z(n2969) );
  AND U5939 ( .A(n2970), .B(p_input[7328]), .Z(o[7328]) );
  AND U5940 ( .A(p_input[27328]), .B(p_input[17328]), .Z(n2970) );
  AND U5941 ( .A(n2971), .B(p_input[7327]), .Z(o[7327]) );
  AND U5942 ( .A(p_input[27327]), .B(p_input[17327]), .Z(n2971) );
  AND U5943 ( .A(n2972), .B(p_input[7326]), .Z(o[7326]) );
  AND U5944 ( .A(p_input[27326]), .B(p_input[17326]), .Z(n2972) );
  AND U5945 ( .A(n2973), .B(p_input[7325]), .Z(o[7325]) );
  AND U5946 ( .A(p_input[27325]), .B(p_input[17325]), .Z(n2973) );
  AND U5947 ( .A(n2974), .B(p_input[7324]), .Z(o[7324]) );
  AND U5948 ( .A(p_input[27324]), .B(p_input[17324]), .Z(n2974) );
  AND U5949 ( .A(n2975), .B(p_input[7323]), .Z(o[7323]) );
  AND U5950 ( .A(p_input[27323]), .B(p_input[17323]), .Z(n2975) );
  AND U5951 ( .A(n2976), .B(p_input[7322]), .Z(o[7322]) );
  AND U5952 ( .A(p_input[27322]), .B(p_input[17322]), .Z(n2976) );
  AND U5953 ( .A(n2977), .B(p_input[7321]), .Z(o[7321]) );
  AND U5954 ( .A(p_input[27321]), .B(p_input[17321]), .Z(n2977) );
  AND U5955 ( .A(n2978), .B(p_input[7320]), .Z(o[7320]) );
  AND U5956 ( .A(p_input[27320]), .B(p_input[17320]), .Z(n2978) );
  AND U5957 ( .A(n2979), .B(p_input[731]), .Z(o[731]) );
  AND U5958 ( .A(p_input[20731]), .B(p_input[10731]), .Z(n2979) );
  AND U5959 ( .A(n2980), .B(p_input[7319]), .Z(o[7319]) );
  AND U5960 ( .A(p_input[27319]), .B(p_input[17319]), .Z(n2980) );
  AND U5961 ( .A(n2981), .B(p_input[7318]), .Z(o[7318]) );
  AND U5962 ( .A(p_input[27318]), .B(p_input[17318]), .Z(n2981) );
  AND U5963 ( .A(n2982), .B(p_input[7317]), .Z(o[7317]) );
  AND U5964 ( .A(p_input[27317]), .B(p_input[17317]), .Z(n2982) );
  AND U5965 ( .A(n2983), .B(p_input[7316]), .Z(o[7316]) );
  AND U5966 ( .A(p_input[27316]), .B(p_input[17316]), .Z(n2983) );
  AND U5967 ( .A(n2984), .B(p_input[7315]), .Z(o[7315]) );
  AND U5968 ( .A(p_input[27315]), .B(p_input[17315]), .Z(n2984) );
  AND U5969 ( .A(n2985), .B(p_input[7314]), .Z(o[7314]) );
  AND U5970 ( .A(p_input[27314]), .B(p_input[17314]), .Z(n2985) );
  AND U5971 ( .A(n2986), .B(p_input[7313]), .Z(o[7313]) );
  AND U5972 ( .A(p_input[27313]), .B(p_input[17313]), .Z(n2986) );
  AND U5973 ( .A(n2987), .B(p_input[7312]), .Z(o[7312]) );
  AND U5974 ( .A(p_input[27312]), .B(p_input[17312]), .Z(n2987) );
  AND U5975 ( .A(n2988), .B(p_input[7311]), .Z(o[7311]) );
  AND U5976 ( .A(p_input[27311]), .B(p_input[17311]), .Z(n2988) );
  AND U5977 ( .A(n2989), .B(p_input[7310]), .Z(o[7310]) );
  AND U5978 ( .A(p_input[27310]), .B(p_input[17310]), .Z(n2989) );
  AND U5979 ( .A(n2990), .B(p_input[730]), .Z(o[730]) );
  AND U5980 ( .A(p_input[20730]), .B(p_input[10730]), .Z(n2990) );
  AND U5981 ( .A(n2991), .B(p_input[7309]), .Z(o[7309]) );
  AND U5982 ( .A(p_input[27309]), .B(p_input[17309]), .Z(n2991) );
  AND U5983 ( .A(n2992), .B(p_input[7308]), .Z(o[7308]) );
  AND U5984 ( .A(p_input[27308]), .B(p_input[17308]), .Z(n2992) );
  AND U5985 ( .A(n2993), .B(p_input[7307]), .Z(o[7307]) );
  AND U5986 ( .A(p_input[27307]), .B(p_input[17307]), .Z(n2993) );
  AND U5987 ( .A(n2994), .B(p_input[7306]), .Z(o[7306]) );
  AND U5988 ( .A(p_input[27306]), .B(p_input[17306]), .Z(n2994) );
  AND U5989 ( .A(n2995), .B(p_input[7305]), .Z(o[7305]) );
  AND U5990 ( .A(p_input[27305]), .B(p_input[17305]), .Z(n2995) );
  AND U5991 ( .A(n2996), .B(p_input[7304]), .Z(o[7304]) );
  AND U5992 ( .A(p_input[27304]), .B(p_input[17304]), .Z(n2996) );
  AND U5993 ( .A(n2997), .B(p_input[7303]), .Z(o[7303]) );
  AND U5994 ( .A(p_input[27303]), .B(p_input[17303]), .Z(n2997) );
  AND U5995 ( .A(n2998), .B(p_input[7302]), .Z(o[7302]) );
  AND U5996 ( .A(p_input[27302]), .B(p_input[17302]), .Z(n2998) );
  AND U5997 ( .A(n2999), .B(p_input[7301]), .Z(o[7301]) );
  AND U5998 ( .A(p_input[27301]), .B(p_input[17301]), .Z(n2999) );
  AND U5999 ( .A(n3000), .B(p_input[7300]), .Z(o[7300]) );
  AND U6000 ( .A(p_input[27300]), .B(p_input[17300]), .Z(n3000) );
  AND U6001 ( .A(n3001), .B(p_input[72]), .Z(o[72]) );
  AND U6002 ( .A(p_input[20072]), .B(p_input[10072]), .Z(n3001) );
  AND U6003 ( .A(n3002), .B(p_input[729]), .Z(o[729]) );
  AND U6004 ( .A(p_input[20729]), .B(p_input[10729]), .Z(n3002) );
  AND U6005 ( .A(n3003), .B(p_input[7299]), .Z(o[7299]) );
  AND U6006 ( .A(p_input[27299]), .B(p_input[17299]), .Z(n3003) );
  AND U6007 ( .A(n3004), .B(p_input[7298]), .Z(o[7298]) );
  AND U6008 ( .A(p_input[27298]), .B(p_input[17298]), .Z(n3004) );
  AND U6009 ( .A(n3005), .B(p_input[7297]), .Z(o[7297]) );
  AND U6010 ( .A(p_input[27297]), .B(p_input[17297]), .Z(n3005) );
  AND U6011 ( .A(n3006), .B(p_input[7296]), .Z(o[7296]) );
  AND U6012 ( .A(p_input[27296]), .B(p_input[17296]), .Z(n3006) );
  AND U6013 ( .A(n3007), .B(p_input[7295]), .Z(o[7295]) );
  AND U6014 ( .A(p_input[27295]), .B(p_input[17295]), .Z(n3007) );
  AND U6015 ( .A(n3008), .B(p_input[7294]), .Z(o[7294]) );
  AND U6016 ( .A(p_input[27294]), .B(p_input[17294]), .Z(n3008) );
  AND U6017 ( .A(n3009), .B(p_input[7293]), .Z(o[7293]) );
  AND U6018 ( .A(p_input[27293]), .B(p_input[17293]), .Z(n3009) );
  AND U6019 ( .A(n3010), .B(p_input[7292]), .Z(o[7292]) );
  AND U6020 ( .A(p_input[27292]), .B(p_input[17292]), .Z(n3010) );
  AND U6021 ( .A(n3011), .B(p_input[7291]), .Z(o[7291]) );
  AND U6022 ( .A(p_input[27291]), .B(p_input[17291]), .Z(n3011) );
  AND U6023 ( .A(n3012), .B(p_input[7290]), .Z(o[7290]) );
  AND U6024 ( .A(p_input[27290]), .B(p_input[17290]), .Z(n3012) );
  AND U6025 ( .A(n3013), .B(p_input[728]), .Z(o[728]) );
  AND U6026 ( .A(p_input[20728]), .B(p_input[10728]), .Z(n3013) );
  AND U6027 ( .A(n3014), .B(p_input[7289]), .Z(o[7289]) );
  AND U6028 ( .A(p_input[27289]), .B(p_input[17289]), .Z(n3014) );
  AND U6029 ( .A(n3015), .B(p_input[7288]), .Z(o[7288]) );
  AND U6030 ( .A(p_input[27288]), .B(p_input[17288]), .Z(n3015) );
  AND U6031 ( .A(n3016), .B(p_input[7287]), .Z(o[7287]) );
  AND U6032 ( .A(p_input[27287]), .B(p_input[17287]), .Z(n3016) );
  AND U6033 ( .A(n3017), .B(p_input[7286]), .Z(o[7286]) );
  AND U6034 ( .A(p_input[27286]), .B(p_input[17286]), .Z(n3017) );
  AND U6035 ( .A(n3018), .B(p_input[7285]), .Z(o[7285]) );
  AND U6036 ( .A(p_input[27285]), .B(p_input[17285]), .Z(n3018) );
  AND U6037 ( .A(n3019), .B(p_input[7284]), .Z(o[7284]) );
  AND U6038 ( .A(p_input[27284]), .B(p_input[17284]), .Z(n3019) );
  AND U6039 ( .A(n3020), .B(p_input[7283]), .Z(o[7283]) );
  AND U6040 ( .A(p_input[27283]), .B(p_input[17283]), .Z(n3020) );
  AND U6041 ( .A(n3021), .B(p_input[7282]), .Z(o[7282]) );
  AND U6042 ( .A(p_input[27282]), .B(p_input[17282]), .Z(n3021) );
  AND U6043 ( .A(n3022), .B(p_input[7281]), .Z(o[7281]) );
  AND U6044 ( .A(p_input[27281]), .B(p_input[17281]), .Z(n3022) );
  AND U6045 ( .A(n3023), .B(p_input[7280]), .Z(o[7280]) );
  AND U6046 ( .A(p_input[27280]), .B(p_input[17280]), .Z(n3023) );
  AND U6047 ( .A(n3024), .B(p_input[727]), .Z(o[727]) );
  AND U6048 ( .A(p_input[20727]), .B(p_input[10727]), .Z(n3024) );
  AND U6049 ( .A(n3025), .B(p_input[7279]), .Z(o[7279]) );
  AND U6050 ( .A(p_input[27279]), .B(p_input[17279]), .Z(n3025) );
  AND U6051 ( .A(n3026), .B(p_input[7278]), .Z(o[7278]) );
  AND U6052 ( .A(p_input[27278]), .B(p_input[17278]), .Z(n3026) );
  AND U6053 ( .A(n3027), .B(p_input[7277]), .Z(o[7277]) );
  AND U6054 ( .A(p_input[27277]), .B(p_input[17277]), .Z(n3027) );
  AND U6055 ( .A(n3028), .B(p_input[7276]), .Z(o[7276]) );
  AND U6056 ( .A(p_input[27276]), .B(p_input[17276]), .Z(n3028) );
  AND U6057 ( .A(n3029), .B(p_input[7275]), .Z(o[7275]) );
  AND U6058 ( .A(p_input[27275]), .B(p_input[17275]), .Z(n3029) );
  AND U6059 ( .A(n3030), .B(p_input[7274]), .Z(o[7274]) );
  AND U6060 ( .A(p_input[27274]), .B(p_input[17274]), .Z(n3030) );
  AND U6061 ( .A(n3031), .B(p_input[7273]), .Z(o[7273]) );
  AND U6062 ( .A(p_input[27273]), .B(p_input[17273]), .Z(n3031) );
  AND U6063 ( .A(n3032), .B(p_input[7272]), .Z(o[7272]) );
  AND U6064 ( .A(p_input[27272]), .B(p_input[17272]), .Z(n3032) );
  AND U6065 ( .A(n3033), .B(p_input[7271]), .Z(o[7271]) );
  AND U6066 ( .A(p_input[27271]), .B(p_input[17271]), .Z(n3033) );
  AND U6067 ( .A(n3034), .B(p_input[7270]), .Z(o[7270]) );
  AND U6068 ( .A(p_input[27270]), .B(p_input[17270]), .Z(n3034) );
  AND U6069 ( .A(n3035), .B(p_input[726]), .Z(o[726]) );
  AND U6070 ( .A(p_input[20726]), .B(p_input[10726]), .Z(n3035) );
  AND U6071 ( .A(n3036), .B(p_input[7269]), .Z(o[7269]) );
  AND U6072 ( .A(p_input[27269]), .B(p_input[17269]), .Z(n3036) );
  AND U6073 ( .A(n3037), .B(p_input[7268]), .Z(o[7268]) );
  AND U6074 ( .A(p_input[27268]), .B(p_input[17268]), .Z(n3037) );
  AND U6075 ( .A(n3038), .B(p_input[7267]), .Z(o[7267]) );
  AND U6076 ( .A(p_input[27267]), .B(p_input[17267]), .Z(n3038) );
  AND U6077 ( .A(n3039), .B(p_input[7266]), .Z(o[7266]) );
  AND U6078 ( .A(p_input[27266]), .B(p_input[17266]), .Z(n3039) );
  AND U6079 ( .A(n3040), .B(p_input[7265]), .Z(o[7265]) );
  AND U6080 ( .A(p_input[27265]), .B(p_input[17265]), .Z(n3040) );
  AND U6081 ( .A(n3041), .B(p_input[7264]), .Z(o[7264]) );
  AND U6082 ( .A(p_input[27264]), .B(p_input[17264]), .Z(n3041) );
  AND U6083 ( .A(n3042), .B(p_input[7263]), .Z(o[7263]) );
  AND U6084 ( .A(p_input[27263]), .B(p_input[17263]), .Z(n3042) );
  AND U6085 ( .A(n3043), .B(p_input[7262]), .Z(o[7262]) );
  AND U6086 ( .A(p_input[27262]), .B(p_input[17262]), .Z(n3043) );
  AND U6087 ( .A(n3044), .B(p_input[7261]), .Z(o[7261]) );
  AND U6088 ( .A(p_input[27261]), .B(p_input[17261]), .Z(n3044) );
  AND U6089 ( .A(n3045), .B(p_input[7260]), .Z(o[7260]) );
  AND U6090 ( .A(p_input[27260]), .B(p_input[17260]), .Z(n3045) );
  AND U6091 ( .A(n3046), .B(p_input[725]), .Z(o[725]) );
  AND U6092 ( .A(p_input[20725]), .B(p_input[10725]), .Z(n3046) );
  AND U6093 ( .A(n3047), .B(p_input[7259]), .Z(o[7259]) );
  AND U6094 ( .A(p_input[27259]), .B(p_input[17259]), .Z(n3047) );
  AND U6095 ( .A(n3048), .B(p_input[7258]), .Z(o[7258]) );
  AND U6096 ( .A(p_input[27258]), .B(p_input[17258]), .Z(n3048) );
  AND U6097 ( .A(n3049), .B(p_input[7257]), .Z(o[7257]) );
  AND U6098 ( .A(p_input[27257]), .B(p_input[17257]), .Z(n3049) );
  AND U6099 ( .A(n3050), .B(p_input[7256]), .Z(o[7256]) );
  AND U6100 ( .A(p_input[27256]), .B(p_input[17256]), .Z(n3050) );
  AND U6101 ( .A(n3051), .B(p_input[7255]), .Z(o[7255]) );
  AND U6102 ( .A(p_input[27255]), .B(p_input[17255]), .Z(n3051) );
  AND U6103 ( .A(n3052), .B(p_input[7254]), .Z(o[7254]) );
  AND U6104 ( .A(p_input[27254]), .B(p_input[17254]), .Z(n3052) );
  AND U6105 ( .A(n3053), .B(p_input[7253]), .Z(o[7253]) );
  AND U6106 ( .A(p_input[27253]), .B(p_input[17253]), .Z(n3053) );
  AND U6107 ( .A(n3054), .B(p_input[7252]), .Z(o[7252]) );
  AND U6108 ( .A(p_input[27252]), .B(p_input[17252]), .Z(n3054) );
  AND U6109 ( .A(n3055), .B(p_input[7251]), .Z(o[7251]) );
  AND U6110 ( .A(p_input[27251]), .B(p_input[17251]), .Z(n3055) );
  AND U6111 ( .A(n3056), .B(p_input[7250]), .Z(o[7250]) );
  AND U6112 ( .A(p_input[27250]), .B(p_input[17250]), .Z(n3056) );
  AND U6113 ( .A(n3057), .B(p_input[724]), .Z(o[724]) );
  AND U6114 ( .A(p_input[20724]), .B(p_input[10724]), .Z(n3057) );
  AND U6115 ( .A(n3058), .B(p_input[7249]), .Z(o[7249]) );
  AND U6116 ( .A(p_input[27249]), .B(p_input[17249]), .Z(n3058) );
  AND U6117 ( .A(n3059), .B(p_input[7248]), .Z(o[7248]) );
  AND U6118 ( .A(p_input[27248]), .B(p_input[17248]), .Z(n3059) );
  AND U6119 ( .A(n3060), .B(p_input[7247]), .Z(o[7247]) );
  AND U6120 ( .A(p_input[27247]), .B(p_input[17247]), .Z(n3060) );
  AND U6121 ( .A(n3061), .B(p_input[7246]), .Z(o[7246]) );
  AND U6122 ( .A(p_input[27246]), .B(p_input[17246]), .Z(n3061) );
  AND U6123 ( .A(n3062), .B(p_input[7245]), .Z(o[7245]) );
  AND U6124 ( .A(p_input[27245]), .B(p_input[17245]), .Z(n3062) );
  AND U6125 ( .A(n3063), .B(p_input[7244]), .Z(o[7244]) );
  AND U6126 ( .A(p_input[27244]), .B(p_input[17244]), .Z(n3063) );
  AND U6127 ( .A(n3064), .B(p_input[7243]), .Z(o[7243]) );
  AND U6128 ( .A(p_input[27243]), .B(p_input[17243]), .Z(n3064) );
  AND U6129 ( .A(n3065), .B(p_input[7242]), .Z(o[7242]) );
  AND U6130 ( .A(p_input[27242]), .B(p_input[17242]), .Z(n3065) );
  AND U6131 ( .A(n3066), .B(p_input[7241]), .Z(o[7241]) );
  AND U6132 ( .A(p_input[27241]), .B(p_input[17241]), .Z(n3066) );
  AND U6133 ( .A(n3067), .B(p_input[7240]), .Z(o[7240]) );
  AND U6134 ( .A(p_input[27240]), .B(p_input[17240]), .Z(n3067) );
  AND U6135 ( .A(n3068), .B(p_input[723]), .Z(o[723]) );
  AND U6136 ( .A(p_input[20723]), .B(p_input[10723]), .Z(n3068) );
  AND U6137 ( .A(n3069), .B(p_input[7239]), .Z(o[7239]) );
  AND U6138 ( .A(p_input[27239]), .B(p_input[17239]), .Z(n3069) );
  AND U6139 ( .A(n3070), .B(p_input[7238]), .Z(o[7238]) );
  AND U6140 ( .A(p_input[27238]), .B(p_input[17238]), .Z(n3070) );
  AND U6141 ( .A(n3071), .B(p_input[7237]), .Z(o[7237]) );
  AND U6142 ( .A(p_input[27237]), .B(p_input[17237]), .Z(n3071) );
  AND U6143 ( .A(n3072), .B(p_input[7236]), .Z(o[7236]) );
  AND U6144 ( .A(p_input[27236]), .B(p_input[17236]), .Z(n3072) );
  AND U6145 ( .A(n3073), .B(p_input[7235]), .Z(o[7235]) );
  AND U6146 ( .A(p_input[27235]), .B(p_input[17235]), .Z(n3073) );
  AND U6147 ( .A(n3074), .B(p_input[7234]), .Z(o[7234]) );
  AND U6148 ( .A(p_input[27234]), .B(p_input[17234]), .Z(n3074) );
  AND U6149 ( .A(n3075), .B(p_input[7233]), .Z(o[7233]) );
  AND U6150 ( .A(p_input[27233]), .B(p_input[17233]), .Z(n3075) );
  AND U6151 ( .A(n3076), .B(p_input[7232]), .Z(o[7232]) );
  AND U6152 ( .A(p_input[27232]), .B(p_input[17232]), .Z(n3076) );
  AND U6153 ( .A(n3077), .B(p_input[7231]), .Z(o[7231]) );
  AND U6154 ( .A(p_input[27231]), .B(p_input[17231]), .Z(n3077) );
  AND U6155 ( .A(n3078), .B(p_input[7230]), .Z(o[7230]) );
  AND U6156 ( .A(p_input[27230]), .B(p_input[17230]), .Z(n3078) );
  AND U6157 ( .A(n3079), .B(p_input[722]), .Z(o[722]) );
  AND U6158 ( .A(p_input[20722]), .B(p_input[10722]), .Z(n3079) );
  AND U6159 ( .A(n3080), .B(p_input[7229]), .Z(o[7229]) );
  AND U6160 ( .A(p_input[27229]), .B(p_input[17229]), .Z(n3080) );
  AND U6161 ( .A(n3081), .B(p_input[7228]), .Z(o[7228]) );
  AND U6162 ( .A(p_input[27228]), .B(p_input[17228]), .Z(n3081) );
  AND U6163 ( .A(n3082), .B(p_input[7227]), .Z(o[7227]) );
  AND U6164 ( .A(p_input[27227]), .B(p_input[17227]), .Z(n3082) );
  AND U6165 ( .A(n3083), .B(p_input[7226]), .Z(o[7226]) );
  AND U6166 ( .A(p_input[27226]), .B(p_input[17226]), .Z(n3083) );
  AND U6167 ( .A(n3084), .B(p_input[7225]), .Z(o[7225]) );
  AND U6168 ( .A(p_input[27225]), .B(p_input[17225]), .Z(n3084) );
  AND U6169 ( .A(n3085), .B(p_input[7224]), .Z(o[7224]) );
  AND U6170 ( .A(p_input[27224]), .B(p_input[17224]), .Z(n3085) );
  AND U6171 ( .A(n3086), .B(p_input[7223]), .Z(o[7223]) );
  AND U6172 ( .A(p_input[27223]), .B(p_input[17223]), .Z(n3086) );
  AND U6173 ( .A(n3087), .B(p_input[7222]), .Z(o[7222]) );
  AND U6174 ( .A(p_input[27222]), .B(p_input[17222]), .Z(n3087) );
  AND U6175 ( .A(n3088), .B(p_input[7221]), .Z(o[7221]) );
  AND U6176 ( .A(p_input[27221]), .B(p_input[17221]), .Z(n3088) );
  AND U6177 ( .A(n3089), .B(p_input[7220]), .Z(o[7220]) );
  AND U6178 ( .A(p_input[27220]), .B(p_input[17220]), .Z(n3089) );
  AND U6179 ( .A(n3090), .B(p_input[721]), .Z(o[721]) );
  AND U6180 ( .A(p_input[20721]), .B(p_input[10721]), .Z(n3090) );
  AND U6181 ( .A(n3091), .B(p_input[7219]), .Z(o[7219]) );
  AND U6182 ( .A(p_input[27219]), .B(p_input[17219]), .Z(n3091) );
  AND U6183 ( .A(n3092), .B(p_input[7218]), .Z(o[7218]) );
  AND U6184 ( .A(p_input[27218]), .B(p_input[17218]), .Z(n3092) );
  AND U6185 ( .A(n3093), .B(p_input[7217]), .Z(o[7217]) );
  AND U6186 ( .A(p_input[27217]), .B(p_input[17217]), .Z(n3093) );
  AND U6187 ( .A(n3094), .B(p_input[7216]), .Z(o[7216]) );
  AND U6188 ( .A(p_input[27216]), .B(p_input[17216]), .Z(n3094) );
  AND U6189 ( .A(n3095), .B(p_input[7215]), .Z(o[7215]) );
  AND U6190 ( .A(p_input[27215]), .B(p_input[17215]), .Z(n3095) );
  AND U6191 ( .A(n3096), .B(p_input[7214]), .Z(o[7214]) );
  AND U6192 ( .A(p_input[27214]), .B(p_input[17214]), .Z(n3096) );
  AND U6193 ( .A(n3097), .B(p_input[7213]), .Z(o[7213]) );
  AND U6194 ( .A(p_input[27213]), .B(p_input[17213]), .Z(n3097) );
  AND U6195 ( .A(n3098), .B(p_input[7212]), .Z(o[7212]) );
  AND U6196 ( .A(p_input[27212]), .B(p_input[17212]), .Z(n3098) );
  AND U6197 ( .A(n3099), .B(p_input[7211]), .Z(o[7211]) );
  AND U6198 ( .A(p_input[27211]), .B(p_input[17211]), .Z(n3099) );
  AND U6199 ( .A(n3100), .B(p_input[7210]), .Z(o[7210]) );
  AND U6200 ( .A(p_input[27210]), .B(p_input[17210]), .Z(n3100) );
  AND U6201 ( .A(n3101), .B(p_input[720]), .Z(o[720]) );
  AND U6202 ( .A(p_input[20720]), .B(p_input[10720]), .Z(n3101) );
  AND U6203 ( .A(n3102), .B(p_input[7209]), .Z(o[7209]) );
  AND U6204 ( .A(p_input[27209]), .B(p_input[17209]), .Z(n3102) );
  AND U6205 ( .A(n3103), .B(p_input[7208]), .Z(o[7208]) );
  AND U6206 ( .A(p_input[27208]), .B(p_input[17208]), .Z(n3103) );
  AND U6207 ( .A(n3104), .B(p_input[7207]), .Z(o[7207]) );
  AND U6208 ( .A(p_input[27207]), .B(p_input[17207]), .Z(n3104) );
  AND U6209 ( .A(n3105), .B(p_input[7206]), .Z(o[7206]) );
  AND U6210 ( .A(p_input[27206]), .B(p_input[17206]), .Z(n3105) );
  AND U6211 ( .A(n3106), .B(p_input[7205]), .Z(o[7205]) );
  AND U6212 ( .A(p_input[27205]), .B(p_input[17205]), .Z(n3106) );
  AND U6213 ( .A(n3107), .B(p_input[7204]), .Z(o[7204]) );
  AND U6214 ( .A(p_input[27204]), .B(p_input[17204]), .Z(n3107) );
  AND U6215 ( .A(n3108), .B(p_input[7203]), .Z(o[7203]) );
  AND U6216 ( .A(p_input[27203]), .B(p_input[17203]), .Z(n3108) );
  AND U6217 ( .A(n3109), .B(p_input[7202]), .Z(o[7202]) );
  AND U6218 ( .A(p_input[27202]), .B(p_input[17202]), .Z(n3109) );
  AND U6219 ( .A(n3110), .B(p_input[7201]), .Z(o[7201]) );
  AND U6220 ( .A(p_input[27201]), .B(p_input[17201]), .Z(n3110) );
  AND U6221 ( .A(n3111), .B(p_input[7200]), .Z(o[7200]) );
  AND U6222 ( .A(p_input[27200]), .B(p_input[17200]), .Z(n3111) );
  AND U6223 ( .A(n3112), .B(p_input[71]), .Z(o[71]) );
  AND U6224 ( .A(p_input[20071]), .B(p_input[10071]), .Z(n3112) );
  AND U6225 ( .A(n3113), .B(p_input[719]), .Z(o[719]) );
  AND U6226 ( .A(p_input[20719]), .B(p_input[10719]), .Z(n3113) );
  AND U6227 ( .A(n3114), .B(p_input[7199]), .Z(o[7199]) );
  AND U6228 ( .A(p_input[27199]), .B(p_input[17199]), .Z(n3114) );
  AND U6229 ( .A(n3115), .B(p_input[7198]), .Z(o[7198]) );
  AND U6230 ( .A(p_input[27198]), .B(p_input[17198]), .Z(n3115) );
  AND U6231 ( .A(n3116), .B(p_input[7197]), .Z(o[7197]) );
  AND U6232 ( .A(p_input[27197]), .B(p_input[17197]), .Z(n3116) );
  AND U6233 ( .A(n3117), .B(p_input[7196]), .Z(o[7196]) );
  AND U6234 ( .A(p_input[27196]), .B(p_input[17196]), .Z(n3117) );
  AND U6235 ( .A(n3118), .B(p_input[7195]), .Z(o[7195]) );
  AND U6236 ( .A(p_input[27195]), .B(p_input[17195]), .Z(n3118) );
  AND U6237 ( .A(n3119), .B(p_input[7194]), .Z(o[7194]) );
  AND U6238 ( .A(p_input[27194]), .B(p_input[17194]), .Z(n3119) );
  AND U6239 ( .A(n3120), .B(p_input[7193]), .Z(o[7193]) );
  AND U6240 ( .A(p_input[27193]), .B(p_input[17193]), .Z(n3120) );
  AND U6241 ( .A(n3121), .B(p_input[7192]), .Z(o[7192]) );
  AND U6242 ( .A(p_input[27192]), .B(p_input[17192]), .Z(n3121) );
  AND U6243 ( .A(n3122), .B(p_input[7191]), .Z(o[7191]) );
  AND U6244 ( .A(p_input[27191]), .B(p_input[17191]), .Z(n3122) );
  AND U6245 ( .A(n3123), .B(p_input[7190]), .Z(o[7190]) );
  AND U6246 ( .A(p_input[27190]), .B(p_input[17190]), .Z(n3123) );
  AND U6247 ( .A(n3124), .B(p_input[718]), .Z(o[718]) );
  AND U6248 ( .A(p_input[20718]), .B(p_input[10718]), .Z(n3124) );
  AND U6249 ( .A(n3125), .B(p_input[7189]), .Z(o[7189]) );
  AND U6250 ( .A(p_input[27189]), .B(p_input[17189]), .Z(n3125) );
  AND U6251 ( .A(n3126), .B(p_input[7188]), .Z(o[7188]) );
  AND U6252 ( .A(p_input[27188]), .B(p_input[17188]), .Z(n3126) );
  AND U6253 ( .A(n3127), .B(p_input[7187]), .Z(o[7187]) );
  AND U6254 ( .A(p_input[27187]), .B(p_input[17187]), .Z(n3127) );
  AND U6255 ( .A(n3128), .B(p_input[7186]), .Z(o[7186]) );
  AND U6256 ( .A(p_input[27186]), .B(p_input[17186]), .Z(n3128) );
  AND U6257 ( .A(n3129), .B(p_input[7185]), .Z(o[7185]) );
  AND U6258 ( .A(p_input[27185]), .B(p_input[17185]), .Z(n3129) );
  AND U6259 ( .A(n3130), .B(p_input[7184]), .Z(o[7184]) );
  AND U6260 ( .A(p_input[27184]), .B(p_input[17184]), .Z(n3130) );
  AND U6261 ( .A(n3131), .B(p_input[7183]), .Z(o[7183]) );
  AND U6262 ( .A(p_input[27183]), .B(p_input[17183]), .Z(n3131) );
  AND U6263 ( .A(n3132), .B(p_input[7182]), .Z(o[7182]) );
  AND U6264 ( .A(p_input[27182]), .B(p_input[17182]), .Z(n3132) );
  AND U6265 ( .A(n3133), .B(p_input[7181]), .Z(o[7181]) );
  AND U6266 ( .A(p_input[27181]), .B(p_input[17181]), .Z(n3133) );
  AND U6267 ( .A(n3134), .B(p_input[7180]), .Z(o[7180]) );
  AND U6268 ( .A(p_input[27180]), .B(p_input[17180]), .Z(n3134) );
  AND U6269 ( .A(n3135), .B(p_input[717]), .Z(o[717]) );
  AND U6270 ( .A(p_input[20717]), .B(p_input[10717]), .Z(n3135) );
  AND U6271 ( .A(n3136), .B(p_input[7179]), .Z(o[7179]) );
  AND U6272 ( .A(p_input[27179]), .B(p_input[17179]), .Z(n3136) );
  AND U6273 ( .A(n3137), .B(p_input[7178]), .Z(o[7178]) );
  AND U6274 ( .A(p_input[27178]), .B(p_input[17178]), .Z(n3137) );
  AND U6275 ( .A(n3138), .B(p_input[7177]), .Z(o[7177]) );
  AND U6276 ( .A(p_input[27177]), .B(p_input[17177]), .Z(n3138) );
  AND U6277 ( .A(n3139), .B(p_input[7176]), .Z(o[7176]) );
  AND U6278 ( .A(p_input[27176]), .B(p_input[17176]), .Z(n3139) );
  AND U6279 ( .A(n3140), .B(p_input[7175]), .Z(o[7175]) );
  AND U6280 ( .A(p_input[27175]), .B(p_input[17175]), .Z(n3140) );
  AND U6281 ( .A(n3141), .B(p_input[7174]), .Z(o[7174]) );
  AND U6282 ( .A(p_input[27174]), .B(p_input[17174]), .Z(n3141) );
  AND U6283 ( .A(n3142), .B(p_input[7173]), .Z(o[7173]) );
  AND U6284 ( .A(p_input[27173]), .B(p_input[17173]), .Z(n3142) );
  AND U6285 ( .A(n3143), .B(p_input[7172]), .Z(o[7172]) );
  AND U6286 ( .A(p_input[27172]), .B(p_input[17172]), .Z(n3143) );
  AND U6287 ( .A(n3144), .B(p_input[7171]), .Z(o[7171]) );
  AND U6288 ( .A(p_input[27171]), .B(p_input[17171]), .Z(n3144) );
  AND U6289 ( .A(n3145), .B(p_input[7170]), .Z(o[7170]) );
  AND U6290 ( .A(p_input[27170]), .B(p_input[17170]), .Z(n3145) );
  AND U6291 ( .A(n3146), .B(p_input[716]), .Z(o[716]) );
  AND U6292 ( .A(p_input[20716]), .B(p_input[10716]), .Z(n3146) );
  AND U6293 ( .A(n3147), .B(p_input[7169]), .Z(o[7169]) );
  AND U6294 ( .A(p_input[27169]), .B(p_input[17169]), .Z(n3147) );
  AND U6295 ( .A(n3148), .B(p_input[7168]), .Z(o[7168]) );
  AND U6296 ( .A(p_input[27168]), .B(p_input[17168]), .Z(n3148) );
  AND U6297 ( .A(n3149), .B(p_input[7167]), .Z(o[7167]) );
  AND U6298 ( .A(p_input[27167]), .B(p_input[17167]), .Z(n3149) );
  AND U6299 ( .A(n3150), .B(p_input[7166]), .Z(o[7166]) );
  AND U6300 ( .A(p_input[27166]), .B(p_input[17166]), .Z(n3150) );
  AND U6301 ( .A(n3151), .B(p_input[7165]), .Z(o[7165]) );
  AND U6302 ( .A(p_input[27165]), .B(p_input[17165]), .Z(n3151) );
  AND U6303 ( .A(n3152), .B(p_input[7164]), .Z(o[7164]) );
  AND U6304 ( .A(p_input[27164]), .B(p_input[17164]), .Z(n3152) );
  AND U6305 ( .A(n3153), .B(p_input[7163]), .Z(o[7163]) );
  AND U6306 ( .A(p_input[27163]), .B(p_input[17163]), .Z(n3153) );
  AND U6307 ( .A(n3154), .B(p_input[7162]), .Z(o[7162]) );
  AND U6308 ( .A(p_input[27162]), .B(p_input[17162]), .Z(n3154) );
  AND U6309 ( .A(n3155), .B(p_input[7161]), .Z(o[7161]) );
  AND U6310 ( .A(p_input[27161]), .B(p_input[17161]), .Z(n3155) );
  AND U6311 ( .A(n3156), .B(p_input[7160]), .Z(o[7160]) );
  AND U6312 ( .A(p_input[27160]), .B(p_input[17160]), .Z(n3156) );
  AND U6313 ( .A(n3157), .B(p_input[715]), .Z(o[715]) );
  AND U6314 ( .A(p_input[20715]), .B(p_input[10715]), .Z(n3157) );
  AND U6315 ( .A(n3158), .B(p_input[7159]), .Z(o[7159]) );
  AND U6316 ( .A(p_input[27159]), .B(p_input[17159]), .Z(n3158) );
  AND U6317 ( .A(n3159), .B(p_input[7158]), .Z(o[7158]) );
  AND U6318 ( .A(p_input[27158]), .B(p_input[17158]), .Z(n3159) );
  AND U6319 ( .A(n3160), .B(p_input[7157]), .Z(o[7157]) );
  AND U6320 ( .A(p_input[27157]), .B(p_input[17157]), .Z(n3160) );
  AND U6321 ( .A(n3161), .B(p_input[7156]), .Z(o[7156]) );
  AND U6322 ( .A(p_input[27156]), .B(p_input[17156]), .Z(n3161) );
  AND U6323 ( .A(n3162), .B(p_input[7155]), .Z(o[7155]) );
  AND U6324 ( .A(p_input[27155]), .B(p_input[17155]), .Z(n3162) );
  AND U6325 ( .A(n3163), .B(p_input[7154]), .Z(o[7154]) );
  AND U6326 ( .A(p_input[27154]), .B(p_input[17154]), .Z(n3163) );
  AND U6327 ( .A(n3164), .B(p_input[7153]), .Z(o[7153]) );
  AND U6328 ( .A(p_input[27153]), .B(p_input[17153]), .Z(n3164) );
  AND U6329 ( .A(n3165), .B(p_input[7152]), .Z(o[7152]) );
  AND U6330 ( .A(p_input[27152]), .B(p_input[17152]), .Z(n3165) );
  AND U6331 ( .A(n3166), .B(p_input[7151]), .Z(o[7151]) );
  AND U6332 ( .A(p_input[27151]), .B(p_input[17151]), .Z(n3166) );
  AND U6333 ( .A(n3167), .B(p_input[7150]), .Z(o[7150]) );
  AND U6334 ( .A(p_input[27150]), .B(p_input[17150]), .Z(n3167) );
  AND U6335 ( .A(n3168), .B(p_input[714]), .Z(o[714]) );
  AND U6336 ( .A(p_input[20714]), .B(p_input[10714]), .Z(n3168) );
  AND U6337 ( .A(n3169), .B(p_input[7149]), .Z(o[7149]) );
  AND U6338 ( .A(p_input[27149]), .B(p_input[17149]), .Z(n3169) );
  AND U6339 ( .A(n3170), .B(p_input[7148]), .Z(o[7148]) );
  AND U6340 ( .A(p_input[27148]), .B(p_input[17148]), .Z(n3170) );
  AND U6341 ( .A(n3171), .B(p_input[7147]), .Z(o[7147]) );
  AND U6342 ( .A(p_input[27147]), .B(p_input[17147]), .Z(n3171) );
  AND U6343 ( .A(n3172), .B(p_input[7146]), .Z(o[7146]) );
  AND U6344 ( .A(p_input[27146]), .B(p_input[17146]), .Z(n3172) );
  AND U6345 ( .A(n3173), .B(p_input[7145]), .Z(o[7145]) );
  AND U6346 ( .A(p_input[27145]), .B(p_input[17145]), .Z(n3173) );
  AND U6347 ( .A(n3174), .B(p_input[7144]), .Z(o[7144]) );
  AND U6348 ( .A(p_input[27144]), .B(p_input[17144]), .Z(n3174) );
  AND U6349 ( .A(n3175), .B(p_input[7143]), .Z(o[7143]) );
  AND U6350 ( .A(p_input[27143]), .B(p_input[17143]), .Z(n3175) );
  AND U6351 ( .A(n3176), .B(p_input[7142]), .Z(o[7142]) );
  AND U6352 ( .A(p_input[27142]), .B(p_input[17142]), .Z(n3176) );
  AND U6353 ( .A(n3177), .B(p_input[7141]), .Z(o[7141]) );
  AND U6354 ( .A(p_input[27141]), .B(p_input[17141]), .Z(n3177) );
  AND U6355 ( .A(n3178), .B(p_input[7140]), .Z(o[7140]) );
  AND U6356 ( .A(p_input[27140]), .B(p_input[17140]), .Z(n3178) );
  AND U6357 ( .A(n3179), .B(p_input[713]), .Z(o[713]) );
  AND U6358 ( .A(p_input[20713]), .B(p_input[10713]), .Z(n3179) );
  AND U6359 ( .A(n3180), .B(p_input[7139]), .Z(o[7139]) );
  AND U6360 ( .A(p_input[27139]), .B(p_input[17139]), .Z(n3180) );
  AND U6361 ( .A(n3181), .B(p_input[7138]), .Z(o[7138]) );
  AND U6362 ( .A(p_input[27138]), .B(p_input[17138]), .Z(n3181) );
  AND U6363 ( .A(n3182), .B(p_input[7137]), .Z(o[7137]) );
  AND U6364 ( .A(p_input[27137]), .B(p_input[17137]), .Z(n3182) );
  AND U6365 ( .A(n3183), .B(p_input[7136]), .Z(o[7136]) );
  AND U6366 ( .A(p_input[27136]), .B(p_input[17136]), .Z(n3183) );
  AND U6367 ( .A(n3184), .B(p_input[7135]), .Z(o[7135]) );
  AND U6368 ( .A(p_input[27135]), .B(p_input[17135]), .Z(n3184) );
  AND U6369 ( .A(n3185), .B(p_input[7134]), .Z(o[7134]) );
  AND U6370 ( .A(p_input[27134]), .B(p_input[17134]), .Z(n3185) );
  AND U6371 ( .A(n3186), .B(p_input[7133]), .Z(o[7133]) );
  AND U6372 ( .A(p_input[27133]), .B(p_input[17133]), .Z(n3186) );
  AND U6373 ( .A(n3187), .B(p_input[7132]), .Z(o[7132]) );
  AND U6374 ( .A(p_input[27132]), .B(p_input[17132]), .Z(n3187) );
  AND U6375 ( .A(n3188), .B(p_input[7131]), .Z(o[7131]) );
  AND U6376 ( .A(p_input[27131]), .B(p_input[17131]), .Z(n3188) );
  AND U6377 ( .A(n3189), .B(p_input[7130]), .Z(o[7130]) );
  AND U6378 ( .A(p_input[27130]), .B(p_input[17130]), .Z(n3189) );
  AND U6379 ( .A(n3190), .B(p_input[712]), .Z(o[712]) );
  AND U6380 ( .A(p_input[20712]), .B(p_input[10712]), .Z(n3190) );
  AND U6381 ( .A(n3191), .B(p_input[7129]), .Z(o[7129]) );
  AND U6382 ( .A(p_input[27129]), .B(p_input[17129]), .Z(n3191) );
  AND U6383 ( .A(n3192), .B(p_input[7128]), .Z(o[7128]) );
  AND U6384 ( .A(p_input[27128]), .B(p_input[17128]), .Z(n3192) );
  AND U6385 ( .A(n3193), .B(p_input[7127]), .Z(o[7127]) );
  AND U6386 ( .A(p_input[27127]), .B(p_input[17127]), .Z(n3193) );
  AND U6387 ( .A(n3194), .B(p_input[7126]), .Z(o[7126]) );
  AND U6388 ( .A(p_input[27126]), .B(p_input[17126]), .Z(n3194) );
  AND U6389 ( .A(n3195), .B(p_input[7125]), .Z(o[7125]) );
  AND U6390 ( .A(p_input[27125]), .B(p_input[17125]), .Z(n3195) );
  AND U6391 ( .A(n3196), .B(p_input[7124]), .Z(o[7124]) );
  AND U6392 ( .A(p_input[27124]), .B(p_input[17124]), .Z(n3196) );
  AND U6393 ( .A(n3197), .B(p_input[7123]), .Z(o[7123]) );
  AND U6394 ( .A(p_input[27123]), .B(p_input[17123]), .Z(n3197) );
  AND U6395 ( .A(n3198), .B(p_input[7122]), .Z(o[7122]) );
  AND U6396 ( .A(p_input[27122]), .B(p_input[17122]), .Z(n3198) );
  AND U6397 ( .A(n3199), .B(p_input[7121]), .Z(o[7121]) );
  AND U6398 ( .A(p_input[27121]), .B(p_input[17121]), .Z(n3199) );
  AND U6399 ( .A(n3200), .B(p_input[7120]), .Z(o[7120]) );
  AND U6400 ( .A(p_input[27120]), .B(p_input[17120]), .Z(n3200) );
  AND U6401 ( .A(n3201), .B(p_input[711]), .Z(o[711]) );
  AND U6402 ( .A(p_input[20711]), .B(p_input[10711]), .Z(n3201) );
  AND U6403 ( .A(n3202), .B(p_input[7119]), .Z(o[7119]) );
  AND U6404 ( .A(p_input[27119]), .B(p_input[17119]), .Z(n3202) );
  AND U6405 ( .A(n3203), .B(p_input[7118]), .Z(o[7118]) );
  AND U6406 ( .A(p_input[27118]), .B(p_input[17118]), .Z(n3203) );
  AND U6407 ( .A(n3204), .B(p_input[7117]), .Z(o[7117]) );
  AND U6408 ( .A(p_input[27117]), .B(p_input[17117]), .Z(n3204) );
  AND U6409 ( .A(n3205), .B(p_input[7116]), .Z(o[7116]) );
  AND U6410 ( .A(p_input[27116]), .B(p_input[17116]), .Z(n3205) );
  AND U6411 ( .A(n3206), .B(p_input[7115]), .Z(o[7115]) );
  AND U6412 ( .A(p_input[27115]), .B(p_input[17115]), .Z(n3206) );
  AND U6413 ( .A(n3207), .B(p_input[7114]), .Z(o[7114]) );
  AND U6414 ( .A(p_input[27114]), .B(p_input[17114]), .Z(n3207) );
  AND U6415 ( .A(n3208), .B(p_input[7113]), .Z(o[7113]) );
  AND U6416 ( .A(p_input[27113]), .B(p_input[17113]), .Z(n3208) );
  AND U6417 ( .A(n3209), .B(p_input[7112]), .Z(o[7112]) );
  AND U6418 ( .A(p_input[27112]), .B(p_input[17112]), .Z(n3209) );
  AND U6419 ( .A(n3210), .B(p_input[7111]), .Z(o[7111]) );
  AND U6420 ( .A(p_input[27111]), .B(p_input[17111]), .Z(n3210) );
  AND U6421 ( .A(n3211), .B(p_input[7110]), .Z(o[7110]) );
  AND U6422 ( .A(p_input[27110]), .B(p_input[17110]), .Z(n3211) );
  AND U6423 ( .A(n3212), .B(p_input[710]), .Z(o[710]) );
  AND U6424 ( .A(p_input[20710]), .B(p_input[10710]), .Z(n3212) );
  AND U6425 ( .A(n3213), .B(p_input[7109]), .Z(o[7109]) );
  AND U6426 ( .A(p_input[27109]), .B(p_input[17109]), .Z(n3213) );
  AND U6427 ( .A(n3214), .B(p_input[7108]), .Z(o[7108]) );
  AND U6428 ( .A(p_input[27108]), .B(p_input[17108]), .Z(n3214) );
  AND U6429 ( .A(n3215), .B(p_input[7107]), .Z(o[7107]) );
  AND U6430 ( .A(p_input[27107]), .B(p_input[17107]), .Z(n3215) );
  AND U6431 ( .A(n3216), .B(p_input[7106]), .Z(o[7106]) );
  AND U6432 ( .A(p_input[27106]), .B(p_input[17106]), .Z(n3216) );
  AND U6433 ( .A(n3217), .B(p_input[7105]), .Z(o[7105]) );
  AND U6434 ( .A(p_input[27105]), .B(p_input[17105]), .Z(n3217) );
  AND U6435 ( .A(n3218), .B(p_input[7104]), .Z(o[7104]) );
  AND U6436 ( .A(p_input[27104]), .B(p_input[17104]), .Z(n3218) );
  AND U6437 ( .A(n3219), .B(p_input[7103]), .Z(o[7103]) );
  AND U6438 ( .A(p_input[27103]), .B(p_input[17103]), .Z(n3219) );
  AND U6439 ( .A(n3220), .B(p_input[7102]), .Z(o[7102]) );
  AND U6440 ( .A(p_input[27102]), .B(p_input[17102]), .Z(n3220) );
  AND U6441 ( .A(n3221), .B(p_input[7101]), .Z(o[7101]) );
  AND U6442 ( .A(p_input[27101]), .B(p_input[17101]), .Z(n3221) );
  AND U6443 ( .A(n3222), .B(p_input[7100]), .Z(o[7100]) );
  AND U6444 ( .A(p_input[27100]), .B(p_input[17100]), .Z(n3222) );
  AND U6445 ( .A(n3223), .B(p_input[70]), .Z(o[70]) );
  AND U6446 ( .A(p_input[20070]), .B(p_input[10070]), .Z(n3223) );
  AND U6447 ( .A(n3224), .B(p_input[709]), .Z(o[709]) );
  AND U6448 ( .A(p_input[20709]), .B(p_input[10709]), .Z(n3224) );
  AND U6449 ( .A(n3225), .B(p_input[7099]), .Z(o[7099]) );
  AND U6450 ( .A(p_input[27099]), .B(p_input[17099]), .Z(n3225) );
  AND U6451 ( .A(n3226), .B(p_input[7098]), .Z(o[7098]) );
  AND U6452 ( .A(p_input[27098]), .B(p_input[17098]), .Z(n3226) );
  AND U6453 ( .A(n3227), .B(p_input[7097]), .Z(o[7097]) );
  AND U6454 ( .A(p_input[27097]), .B(p_input[17097]), .Z(n3227) );
  AND U6455 ( .A(n3228), .B(p_input[7096]), .Z(o[7096]) );
  AND U6456 ( .A(p_input[27096]), .B(p_input[17096]), .Z(n3228) );
  AND U6457 ( .A(n3229), .B(p_input[7095]), .Z(o[7095]) );
  AND U6458 ( .A(p_input[27095]), .B(p_input[17095]), .Z(n3229) );
  AND U6459 ( .A(n3230), .B(p_input[7094]), .Z(o[7094]) );
  AND U6460 ( .A(p_input[27094]), .B(p_input[17094]), .Z(n3230) );
  AND U6461 ( .A(n3231), .B(p_input[7093]), .Z(o[7093]) );
  AND U6462 ( .A(p_input[27093]), .B(p_input[17093]), .Z(n3231) );
  AND U6463 ( .A(n3232), .B(p_input[7092]), .Z(o[7092]) );
  AND U6464 ( .A(p_input[27092]), .B(p_input[17092]), .Z(n3232) );
  AND U6465 ( .A(n3233), .B(p_input[7091]), .Z(o[7091]) );
  AND U6466 ( .A(p_input[27091]), .B(p_input[17091]), .Z(n3233) );
  AND U6467 ( .A(n3234), .B(p_input[7090]), .Z(o[7090]) );
  AND U6468 ( .A(p_input[27090]), .B(p_input[17090]), .Z(n3234) );
  AND U6469 ( .A(n3235), .B(p_input[708]), .Z(o[708]) );
  AND U6470 ( .A(p_input[20708]), .B(p_input[10708]), .Z(n3235) );
  AND U6471 ( .A(n3236), .B(p_input[7089]), .Z(o[7089]) );
  AND U6472 ( .A(p_input[27089]), .B(p_input[17089]), .Z(n3236) );
  AND U6473 ( .A(n3237), .B(p_input[7088]), .Z(o[7088]) );
  AND U6474 ( .A(p_input[27088]), .B(p_input[17088]), .Z(n3237) );
  AND U6475 ( .A(n3238), .B(p_input[7087]), .Z(o[7087]) );
  AND U6476 ( .A(p_input[27087]), .B(p_input[17087]), .Z(n3238) );
  AND U6477 ( .A(n3239), .B(p_input[7086]), .Z(o[7086]) );
  AND U6478 ( .A(p_input[27086]), .B(p_input[17086]), .Z(n3239) );
  AND U6479 ( .A(n3240), .B(p_input[7085]), .Z(o[7085]) );
  AND U6480 ( .A(p_input[27085]), .B(p_input[17085]), .Z(n3240) );
  AND U6481 ( .A(n3241), .B(p_input[7084]), .Z(o[7084]) );
  AND U6482 ( .A(p_input[27084]), .B(p_input[17084]), .Z(n3241) );
  AND U6483 ( .A(n3242), .B(p_input[7083]), .Z(o[7083]) );
  AND U6484 ( .A(p_input[27083]), .B(p_input[17083]), .Z(n3242) );
  AND U6485 ( .A(n3243), .B(p_input[7082]), .Z(o[7082]) );
  AND U6486 ( .A(p_input[27082]), .B(p_input[17082]), .Z(n3243) );
  AND U6487 ( .A(n3244), .B(p_input[7081]), .Z(o[7081]) );
  AND U6488 ( .A(p_input[27081]), .B(p_input[17081]), .Z(n3244) );
  AND U6489 ( .A(n3245), .B(p_input[7080]), .Z(o[7080]) );
  AND U6490 ( .A(p_input[27080]), .B(p_input[17080]), .Z(n3245) );
  AND U6491 ( .A(n3246), .B(p_input[707]), .Z(o[707]) );
  AND U6492 ( .A(p_input[20707]), .B(p_input[10707]), .Z(n3246) );
  AND U6493 ( .A(n3247), .B(p_input[7079]), .Z(o[7079]) );
  AND U6494 ( .A(p_input[27079]), .B(p_input[17079]), .Z(n3247) );
  AND U6495 ( .A(n3248), .B(p_input[7078]), .Z(o[7078]) );
  AND U6496 ( .A(p_input[27078]), .B(p_input[17078]), .Z(n3248) );
  AND U6497 ( .A(n3249), .B(p_input[7077]), .Z(o[7077]) );
  AND U6498 ( .A(p_input[27077]), .B(p_input[17077]), .Z(n3249) );
  AND U6499 ( .A(n3250), .B(p_input[7076]), .Z(o[7076]) );
  AND U6500 ( .A(p_input[27076]), .B(p_input[17076]), .Z(n3250) );
  AND U6501 ( .A(n3251), .B(p_input[7075]), .Z(o[7075]) );
  AND U6502 ( .A(p_input[27075]), .B(p_input[17075]), .Z(n3251) );
  AND U6503 ( .A(n3252), .B(p_input[7074]), .Z(o[7074]) );
  AND U6504 ( .A(p_input[27074]), .B(p_input[17074]), .Z(n3252) );
  AND U6505 ( .A(n3253), .B(p_input[7073]), .Z(o[7073]) );
  AND U6506 ( .A(p_input[27073]), .B(p_input[17073]), .Z(n3253) );
  AND U6507 ( .A(n3254), .B(p_input[7072]), .Z(o[7072]) );
  AND U6508 ( .A(p_input[27072]), .B(p_input[17072]), .Z(n3254) );
  AND U6509 ( .A(n3255), .B(p_input[7071]), .Z(o[7071]) );
  AND U6510 ( .A(p_input[27071]), .B(p_input[17071]), .Z(n3255) );
  AND U6511 ( .A(n3256), .B(p_input[7070]), .Z(o[7070]) );
  AND U6512 ( .A(p_input[27070]), .B(p_input[17070]), .Z(n3256) );
  AND U6513 ( .A(n3257), .B(p_input[706]), .Z(o[706]) );
  AND U6514 ( .A(p_input[20706]), .B(p_input[10706]), .Z(n3257) );
  AND U6515 ( .A(n3258), .B(p_input[7069]), .Z(o[7069]) );
  AND U6516 ( .A(p_input[27069]), .B(p_input[17069]), .Z(n3258) );
  AND U6517 ( .A(n3259), .B(p_input[7068]), .Z(o[7068]) );
  AND U6518 ( .A(p_input[27068]), .B(p_input[17068]), .Z(n3259) );
  AND U6519 ( .A(n3260), .B(p_input[7067]), .Z(o[7067]) );
  AND U6520 ( .A(p_input[27067]), .B(p_input[17067]), .Z(n3260) );
  AND U6521 ( .A(n3261), .B(p_input[7066]), .Z(o[7066]) );
  AND U6522 ( .A(p_input[27066]), .B(p_input[17066]), .Z(n3261) );
  AND U6523 ( .A(n3262), .B(p_input[7065]), .Z(o[7065]) );
  AND U6524 ( .A(p_input[27065]), .B(p_input[17065]), .Z(n3262) );
  AND U6525 ( .A(n3263), .B(p_input[7064]), .Z(o[7064]) );
  AND U6526 ( .A(p_input[27064]), .B(p_input[17064]), .Z(n3263) );
  AND U6527 ( .A(n3264), .B(p_input[7063]), .Z(o[7063]) );
  AND U6528 ( .A(p_input[27063]), .B(p_input[17063]), .Z(n3264) );
  AND U6529 ( .A(n3265), .B(p_input[7062]), .Z(o[7062]) );
  AND U6530 ( .A(p_input[27062]), .B(p_input[17062]), .Z(n3265) );
  AND U6531 ( .A(n3266), .B(p_input[7061]), .Z(o[7061]) );
  AND U6532 ( .A(p_input[27061]), .B(p_input[17061]), .Z(n3266) );
  AND U6533 ( .A(n3267), .B(p_input[7060]), .Z(o[7060]) );
  AND U6534 ( .A(p_input[27060]), .B(p_input[17060]), .Z(n3267) );
  AND U6535 ( .A(n3268), .B(p_input[705]), .Z(o[705]) );
  AND U6536 ( .A(p_input[20705]), .B(p_input[10705]), .Z(n3268) );
  AND U6537 ( .A(n3269), .B(p_input[7059]), .Z(o[7059]) );
  AND U6538 ( .A(p_input[27059]), .B(p_input[17059]), .Z(n3269) );
  AND U6539 ( .A(n3270), .B(p_input[7058]), .Z(o[7058]) );
  AND U6540 ( .A(p_input[27058]), .B(p_input[17058]), .Z(n3270) );
  AND U6541 ( .A(n3271), .B(p_input[7057]), .Z(o[7057]) );
  AND U6542 ( .A(p_input[27057]), .B(p_input[17057]), .Z(n3271) );
  AND U6543 ( .A(n3272), .B(p_input[7056]), .Z(o[7056]) );
  AND U6544 ( .A(p_input[27056]), .B(p_input[17056]), .Z(n3272) );
  AND U6545 ( .A(n3273), .B(p_input[7055]), .Z(o[7055]) );
  AND U6546 ( .A(p_input[27055]), .B(p_input[17055]), .Z(n3273) );
  AND U6547 ( .A(n3274), .B(p_input[7054]), .Z(o[7054]) );
  AND U6548 ( .A(p_input[27054]), .B(p_input[17054]), .Z(n3274) );
  AND U6549 ( .A(n3275), .B(p_input[7053]), .Z(o[7053]) );
  AND U6550 ( .A(p_input[27053]), .B(p_input[17053]), .Z(n3275) );
  AND U6551 ( .A(n3276), .B(p_input[7052]), .Z(o[7052]) );
  AND U6552 ( .A(p_input[27052]), .B(p_input[17052]), .Z(n3276) );
  AND U6553 ( .A(n3277), .B(p_input[7051]), .Z(o[7051]) );
  AND U6554 ( .A(p_input[27051]), .B(p_input[17051]), .Z(n3277) );
  AND U6555 ( .A(n3278), .B(p_input[7050]), .Z(o[7050]) );
  AND U6556 ( .A(p_input[27050]), .B(p_input[17050]), .Z(n3278) );
  AND U6557 ( .A(n3279), .B(p_input[704]), .Z(o[704]) );
  AND U6558 ( .A(p_input[20704]), .B(p_input[10704]), .Z(n3279) );
  AND U6559 ( .A(n3280), .B(p_input[7049]), .Z(o[7049]) );
  AND U6560 ( .A(p_input[27049]), .B(p_input[17049]), .Z(n3280) );
  AND U6561 ( .A(n3281), .B(p_input[7048]), .Z(o[7048]) );
  AND U6562 ( .A(p_input[27048]), .B(p_input[17048]), .Z(n3281) );
  AND U6563 ( .A(n3282), .B(p_input[7047]), .Z(o[7047]) );
  AND U6564 ( .A(p_input[27047]), .B(p_input[17047]), .Z(n3282) );
  AND U6565 ( .A(n3283), .B(p_input[7046]), .Z(o[7046]) );
  AND U6566 ( .A(p_input[27046]), .B(p_input[17046]), .Z(n3283) );
  AND U6567 ( .A(n3284), .B(p_input[7045]), .Z(o[7045]) );
  AND U6568 ( .A(p_input[27045]), .B(p_input[17045]), .Z(n3284) );
  AND U6569 ( .A(n3285), .B(p_input[7044]), .Z(o[7044]) );
  AND U6570 ( .A(p_input[27044]), .B(p_input[17044]), .Z(n3285) );
  AND U6571 ( .A(n3286), .B(p_input[7043]), .Z(o[7043]) );
  AND U6572 ( .A(p_input[27043]), .B(p_input[17043]), .Z(n3286) );
  AND U6573 ( .A(n3287), .B(p_input[7042]), .Z(o[7042]) );
  AND U6574 ( .A(p_input[27042]), .B(p_input[17042]), .Z(n3287) );
  AND U6575 ( .A(n3288), .B(p_input[7041]), .Z(o[7041]) );
  AND U6576 ( .A(p_input[27041]), .B(p_input[17041]), .Z(n3288) );
  AND U6577 ( .A(n3289), .B(p_input[7040]), .Z(o[7040]) );
  AND U6578 ( .A(p_input[27040]), .B(p_input[17040]), .Z(n3289) );
  AND U6579 ( .A(n3290), .B(p_input[703]), .Z(o[703]) );
  AND U6580 ( .A(p_input[20703]), .B(p_input[10703]), .Z(n3290) );
  AND U6581 ( .A(n3291), .B(p_input[7039]), .Z(o[7039]) );
  AND U6582 ( .A(p_input[27039]), .B(p_input[17039]), .Z(n3291) );
  AND U6583 ( .A(n3292), .B(p_input[7038]), .Z(o[7038]) );
  AND U6584 ( .A(p_input[27038]), .B(p_input[17038]), .Z(n3292) );
  AND U6585 ( .A(n3293), .B(p_input[7037]), .Z(o[7037]) );
  AND U6586 ( .A(p_input[27037]), .B(p_input[17037]), .Z(n3293) );
  AND U6587 ( .A(n3294), .B(p_input[7036]), .Z(o[7036]) );
  AND U6588 ( .A(p_input[27036]), .B(p_input[17036]), .Z(n3294) );
  AND U6589 ( .A(n3295), .B(p_input[7035]), .Z(o[7035]) );
  AND U6590 ( .A(p_input[27035]), .B(p_input[17035]), .Z(n3295) );
  AND U6591 ( .A(n3296), .B(p_input[7034]), .Z(o[7034]) );
  AND U6592 ( .A(p_input[27034]), .B(p_input[17034]), .Z(n3296) );
  AND U6593 ( .A(n3297), .B(p_input[7033]), .Z(o[7033]) );
  AND U6594 ( .A(p_input[27033]), .B(p_input[17033]), .Z(n3297) );
  AND U6595 ( .A(n3298), .B(p_input[7032]), .Z(o[7032]) );
  AND U6596 ( .A(p_input[27032]), .B(p_input[17032]), .Z(n3298) );
  AND U6597 ( .A(n3299), .B(p_input[7031]), .Z(o[7031]) );
  AND U6598 ( .A(p_input[27031]), .B(p_input[17031]), .Z(n3299) );
  AND U6599 ( .A(n3300), .B(p_input[7030]), .Z(o[7030]) );
  AND U6600 ( .A(p_input[27030]), .B(p_input[17030]), .Z(n3300) );
  AND U6601 ( .A(n3301), .B(p_input[702]), .Z(o[702]) );
  AND U6602 ( .A(p_input[20702]), .B(p_input[10702]), .Z(n3301) );
  AND U6603 ( .A(n3302), .B(p_input[7029]), .Z(o[7029]) );
  AND U6604 ( .A(p_input[27029]), .B(p_input[17029]), .Z(n3302) );
  AND U6605 ( .A(n3303), .B(p_input[7028]), .Z(o[7028]) );
  AND U6606 ( .A(p_input[27028]), .B(p_input[17028]), .Z(n3303) );
  AND U6607 ( .A(n3304), .B(p_input[7027]), .Z(o[7027]) );
  AND U6608 ( .A(p_input[27027]), .B(p_input[17027]), .Z(n3304) );
  AND U6609 ( .A(n3305), .B(p_input[7026]), .Z(o[7026]) );
  AND U6610 ( .A(p_input[27026]), .B(p_input[17026]), .Z(n3305) );
  AND U6611 ( .A(n3306), .B(p_input[7025]), .Z(o[7025]) );
  AND U6612 ( .A(p_input[27025]), .B(p_input[17025]), .Z(n3306) );
  AND U6613 ( .A(n3307), .B(p_input[7024]), .Z(o[7024]) );
  AND U6614 ( .A(p_input[27024]), .B(p_input[17024]), .Z(n3307) );
  AND U6615 ( .A(n3308), .B(p_input[7023]), .Z(o[7023]) );
  AND U6616 ( .A(p_input[27023]), .B(p_input[17023]), .Z(n3308) );
  AND U6617 ( .A(n3309), .B(p_input[7022]), .Z(o[7022]) );
  AND U6618 ( .A(p_input[27022]), .B(p_input[17022]), .Z(n3309) );
  AND U6619 ( .A(n3310), .B(p_input[7021]), .Z(o[7021]) );
  AND U6620 ( .A(p_input[27021]), .B(p_input[17021]), .Z(n3310) );
  AND U6621 ( .A(n3311), .B(p_input[7020]), .Z(o[7020]) );
  AND U6622 ( .A(p_input[27020]), .B(p_input[17020]), .Z(n3311) );
  AND U6623 ( .A(n3312), .B(p_input[701]), .Z(o[701]) );
  AND U6624 ( .A(p_input[20701]), .B(p_input[10701]), .Z(n3312) );
  AND U6625 ( .A(n3313), .B(p_input[7019]), .Z(o[7019]) );
  AND U6626 ( .A(p_input[27019]), .B(p_input[17019]), .Z(n3313) );
  AND U6627 ( .A(n3314), .B(p_input[7018]), .Z(o[7018]) );
  AND U6628 ( .A(p_input[27018]), .B(p_input[17018]), .Z(n3314) );
  AND U6629 ( .A(n3315), .B(p_input[7017]), .Z(o[7017]) );
  AND U6630 ( .A(p_input[27017]), .B(p_input[17017]), .Z(n3315) );
  AND U6631 ( .A(n3316), .B(p_input[7016]), .Z(o[7016]) );
  AND U6632 ( .A(p_input[27016]), .B(p_input[17016]), .Z(n3316) );
  AND U6633 ( .A(n3317), .B(p_input[7015]), .Z(o[7015]) );
  AND U6634 ( .A(p_input[27015]), .B(p_input[17015]), .Z(n3317) );
  AND U6635 ( .A(n3318), .B(p_input[7014]), .Z(o[7014]) );
  AND U6636 ( .A(p_input[27014]), .B(p_input[17014]), .Z(n3318) );
  AND U6637 ( .A(n3319), .B(p_input[7013]), .Z(o[7013]) );
  AND U6638 ( .A(p_input[27013]), .B(p_input[17013]), .Z(n3319) );
  AND U6639 ( .A(n3320), .B(p_input[7012]), .Z(o[7012]) );
  AND U6640 ( .A(p_input[27012]), .B(p_input[17012]), .Z(n3320) );
  AND U6641 ( .A(n3321), .B(p_input[7011]), .Z(o[7011]) );
  AND U6642 ( .A(p_input[27011]), .B(p_input[17011]), .Z(n3321) );
  AND U6643 ( .A(n3322), .B(p_input[7010]), .Z(o[7010]) );
  AND U6644 ( .A(p_input[27010]), .B(p_input[17010]), .Z(n3322) );
  AND U6645 ( .A(n3323), .B(p_input[700]), .Z(o[700]) );
  AND U6646 ( .A(p_input[20700]), .B(p_input[10700]), .Z(n3323) );
  AND U6647 ( .A(n3324), .B(p_input[7009]), .Z(o[7009]) );
  AND U6648 ( .A(p_input[27009]), .B(p_input[17009]), .Z(n3324) );
  AND U6649 ( .A(n3325), .B(p_input[7008]), .Z(o[7008]) );
  AND U6650 ( .A(p_input[27008]), .B(p_input[17008]), .Z(n3325) );
  AND U6651 ( .A(n3326), .B(p_input[7007]), .Z(o[7007]) );
  AND U6652 ( .A(p_input[27007]), .B(p_input[17007]), .Z(n3326) );
  AND U6653 ( .A(n3327), .B(p_input[7006]), .Z(o[7006]) );
  AND U6654 ( .A(p_input[27006]), .B(p_input[17006]), .Z(n3327) );
  AND U6655 ( .A(n3328), .B(p_input[7005]), .Z(o[7005]) );
  AND U6656 ( .A(p_input[27005]), .B(p_input[17005]), .Z(n3328) );
  AND U6657 ( .A(n3329), .B(p_input[7004]), .Z(o[7004]) );
  AND U6658 ( .A(p_input[27004]), .B(p_input[17004]), .Z(n3329) );
  AND U6659 ( .A(n3330), .B(p_input[7003]), .Z(o[7003]) );
  AND U6660 ( .A(p_input[27003]), .B(p_input[17003]), .Z(n3330) );
  AND U6661 ( .A(n3331), .B(p_input[7002]), .Z(o[7002]) );
  AND U6662 ( .A(p_input[27002]), .B(p_input[17002]), .Z(n3331) );
  AND U6663 ( .A(n3332), .B(p_input[7001]), .Z(o[7001]) );
  AND U6664 ( .A(p_input[27001]), .B(p_input[17001]), .Z(n3332) );
  AND U6665 ( .A(n3333), .B(p_input[7000]), .Z(o[7000]) );
  AND U6666 ( .A(p_input[27000]), .B(p_input[17000]), .Z(n3333) );
  AND U6667 ( .A(n3334), .B(p_input[6]), .Z(o[6]) );
  AND U6668 ( .A(p_input[20006]), .B(p_input[10006]), .Z(n3334) );
  AND U6669 ( .A(n3335), .B(p_input[69]), .Z(o[69]) );
  AND U6670 ( .A(p_input[20069]), .B(p_input[10069]), .Z(n3335) );
  AND U6671 ( .A(n3336), .B(p_input[699]), .Z(o[699]) );
  AND U6672 ( .A(p_input[20699]), .B(p_input[10699]), .Z(n3336) );
  AND U6673 ( .A(n3337), .B(p_input[6999]), .Z(o[6999]) );
  AND U6674 ( .A(p_input[26999]), .B(p_input[16999]), .Z(n3337) );
  AND U6675 ( .A(n3338), .B(p_input[6998]), .Z(o[6998]) );
  AND U6676 ( .A(p_input[26998]), .B(p_input[16998]), .Z(n3338) );
  AND U6677 ( .A(n3339), .B(p_input[6997]), .Z(o[6997]) );
  AND U6678 ( .A(p_input[26997]), .B(p_input[16997]), .Z(n3339) );
  AND U6679 ( .A(n3340), .B(p_input[6996]), .Z(o[6996]) );
  AND U6680 ( .A(p_input[26996]), .B(p_input[16996]), .Z(n3340) );
  AND U6681 ( .A(n3341), .B(p_input[6995]), .Z(o[6995]) );
  AND U6682 ( .A(p_input[26995]), .B(p_input[16995]), .Z(n3341) );
  AND U6683 ( .A(n3342), .B(p_input[6994]), .Z(o[6994]) );
  AND U6684 ( .A(p_input[26994]), .B(p_input[16994]), .Z(n3342) );
  AND U6685 ( .A(n3343), .B(p_input[6993]), .Z(o[6993]) );
  AND U6686 ( .A(p_input[26993]), .B(p_input[16993]), .Z(n3343) );
  AND U6687 ( .A(n3344), .B(p_input[6992]), .Z(o[6992]) );
  AND U6688 ( .A(p_input[26992]), .B(p_input[16992]), .Z(n3344) );
  AND U6689 ( .A(n3345), .B(p_input[6991]), .Z(o[6991]) );
  AND U6690 ( .A(p_input[26991]), .B(p_input[16991]), .Z(n3345) );
  AND U6691 ( .A(n3346), .B(p_input[6990]), .Z(o[6990]) );
  AND U6692 ( .A(p_input[26990]), .B(p_input[16990]), .Z(n3346) );
  AND U6693 ( .A(n3347), .B(p_input[698]), .Z(o[698]) );
  AND U6694 ( .A(p_input[20698]), .B(p_input[10698]), .Z(n3347) );
  AND U6695 ( .A(n3348), .B(p_input[6989]), .Z(o[6989]) );
  AND U6696 ( .A(p_input[26989]), .B(p_input[16989]), .Z(n3348) );
  AND U6697 ( .A(n3349), .B(p_input[6988]), .Z(o[6988]) );
  AND U6698 ( .A(p_input[26988]), .B(p_input[16988]), .Z(n3349) );
  AND U6699 ( .A(n3350), .B(p_input[6987]), .Z(o[6987]) );
  AND U6700 ( .A(p_input[26987]), .B(p_input[16987]), .Z(n3350) );
  AND U6701 ( .A(n3351), .B(p_input[6986]), .Z(o[6986]) );
  AND U6702 ( .A(p_input[26986]), .B(p_input[16986]), .Z(n3351) );
  AND U6703 ( .A(n3352), .B(p_input[6985]), .Z(o[6985]) );
  AND U6704 ( .A(p_input[26985]), .B(p_input[16985]), .Z(n3352) );
  AND U6705 ( .A(n3353), .B(p_input[6984]), .Z(o[6984]) );
  AND U6706 ( .A(p_input[26984]), .B(p_input[16984]), .Z(n3353) );
  AND U6707 ( .A(n3354), .B(p_input[6983]), .Z(o[6983]) );
  AND U6708 ( .A(p_input[26983]), .B(p_input[16983]), .Z(n3354) );
  AND U6709 ( .A(n3355), .B(p_input[6982]), .Z(o[6982]) );
  AND U6710 ( .A(p_input[26982]), .B(p_input[16982]), .Z(n3355) );
  AND U6711 ( .A(n3356), .B(p_input[6981]), .Z(o[6981]) );
  AND U6712 ( .A(p_input[26981]), .B(p_input[16981]), .Z(n3356) );
  AND U6713 ( .A(n3357), .B(p_input[6980]), .Z(o[6980]) );
  AND U6714 ( .A(p_input[26980]), .B(p_input[16980]), .Z(n3357) );
  AND U6715 ( .A(n3358), .B(p_input[697]), .Z(o[697]) );
  AND U6716 ( .A(p_input[20697]), .B(p_input[10697]), .Z(n3358) );
  AND U6717 ( .A(n3359), .B(p_input[6979]), .Z(o[6979]) );
  AND U6718 ( .A(p_input[26979]), .B(p_input[16979]), .Z(n3359) );
  AND U6719 ( .A(n3360), .B(p_input[6978]), .Z(o[6978]) );
  AND U6720 ( .A(p_input[26978]), .B(p_input[16978]), .Z(n3360) );
  AND U6721 ( .A(n3361), .B(p_input[6977]), .Z(o[6977]) );
  AND U6722 ( .A(p_input[26977]), .B(p_input[16977]), .Z(n3361) );
  AND U6723 ( .A(n3362), .B(p_input[6976]), .Z(o[6976]) );
  AND U6724 ( .A(p_input[26976]), .B(p_input[16976]), .Z(n3362) );
  AND U6725 ( .A(n3363), .B(p_input[6975]), .Z(o[6975]) );
  AND U6726 ( .A(p_input[26975]), .B(p_input[16975]), .Z(n3363) );
  AND U6727 ( .A(n3364), .B(p_input[6974]), .Z(o[6974]) );
  AND U6728 ( .A(p_input[26974]), .B(p_input[16974]), .Z(n3364) );
  AND U6729 ( .A(n3365), .B(p_input[6973]), .Z(o[6973]) );
  AND U6730 ( .A(p_input[26973]), .B(p_input[16973]), .Z(n3365) );
  AND U6731 ( .A(n3366), .B(p_input[6972]), .Z(o[6972]) );
  AND U6732 ( .A(p_input[26972]), .B(p_input[16972]), .Z(n3366) );
  AND U6733 ( .A(n3367), .B(p_input[6971]), .Z(o[6971]) );
  AND U6734 ( .A(p_input[26971]), .B(p_input[16971]), .Z(n3367) );
  AND U6735 ( .A(n3368), .B(p_input[6970]), .Z(o[6970]) );
  AND U6736 ( .A(p_input[26970]), .B(p_input[16970]), .Z(n3368) );
  AND U6737 ( .A(n3369), .B(p_input[696]), .Z(o[696]) );
  AND U6738 ( .A(p_input[20696]), .B(p_input[10696]), .Z(n3369) );
  AND U6739 ( .A(n3370), .B(p_input[6969]), .Z(o[6969]) );
  AND U6740 ( .A(p_input[26969]), .B(p_input[16969]), .Z(n3370) );
  AND U6741 ( .A(n3371), .B(p_input[6968]), .Z(o[6968]) );
  AND U6742 ( .A(p_input[26968]), .B(p_input[16968]), .Z(n3371) );
  AND U6743 ( .A(n3372), .B(p_input[6967]), .Z(o[6967]) );
  AND U6744 ( .A(p_input[26967]), .B(p_input[16967]), .Z(n3372) );
  AND U6745 ( .A(n3373), .B(p_input[6966]), .Z(o[6966]) );
  AND U6746 ( .A(p_input[26966]), .B(p_input[16966]), .Z(n3373) );
  AND U6747 ( .A(n3374), .B(p_input[6965]), .Z(o[6965]) );
  AND U6748 ( .A(p_input[26965]), .B(p_input[16965]), .Z(n3374) );
  AND U6749 ( .A(n3375), .B(p_input[6964]), .Z(o[6964]) );
  AND U6750 ( .A(p_input[26964]), .B(p_input[16964]), .Z(n3375) );
  AND U6751 ( .A(n3376), .B(p_input[6963]), .Z(o[6963]) );
  AND U6752 ( .A(p_input[26963]), .B(p_input[16963]), .Z(n3376) );
  AND U6753 ( .A(n3377), .B(p_input[6962]), .Z(o[6962]) );
  AND U6754 ( .A(p_input[26962]), .B(p_input[16962]), .Z(n3377) );
  AND U6755 ( .A(n3378), .B(p_input[6961]), .Z(o[6961]) );
  AND U6756 ( .A(p_input[26961]), .B(p_input[16961]), .Z(n3378) );
  AND U6757 ( .A(n3379), .B(p_input[6960]), .Z(o[6960]) );
  AND U6758 ( .A(p_input[26960]), .B(p_input[16960]), .Z(n3379) );
  AND U6759 ( .A(n3380), .B(p_input[695]), .Z(o[695]) );
  AND U6760 ( .A(p_input[20695]), .B(p_input[10695]), .Z(n3380) );
  AND U6761 ( .A(n3381), .B(p_input[6959]), .Z(o[6959]) );
  AND U6762 ( .A(p_input[26959]), .B(p_input[16959]), .Z(n3381) );
  AND U6763 ( .A(n3382), .B(p_input[6958]), .Z(o[6958]) );
  AND U6764 ( .A(p_input[26958]), .B(p_input[16958]), .Z(n3382) );
  AND U6765 ( .A(n3383), .B(p_input[6957]), .Z(o[6957]) );
  AND U6766 ( .A(p_input[26957]), .B(p_input[16957]), .Z(n3383) );
  AND U6767 ( .A(n3384), .B(p_input[6956]), .Z(o[6956]) );
  AND U6768 ( .A(p_input[26956]), .B(p_input[16956]), .Z(n3384) );
  AND U6769 ( .A(n3385), .B(p_input[6955]), .Z(o[6955]) );
  AND U6770 ( .A(p_input[26955]), .B(p_input[16955]), .Z(n3385) );
  AND U6771 ( .A(n3386), .B(p_input[6954]), .Z(o[6954]) );
  AND U6772 ( .A(p_input[26954]), .B(p_input[16954]), .Z(n3386) );
  AND U6773 ( .A(n3387), .B(p_input[6953]), .Z(o[6953]) );
  AND U6774 ( .A(p_input[26953]), .B(p_input[16953]), .Z(n3387) );
  AND U6775 ( .A(n3388), .B(p_input[6952]), .Z(o[6952]) );
  AND U6776 ( .A(p_input[26952]), .B(p_input[16952]), .Z(n3388) );
  AND U6777 ( .A(n3389), .B(p_input[6951]), .Z(o[6951]) );
  AND U6778 ( .A(p_input[26951]), .B(p_input[16951]), .Z(n3389) );
  AND U6779 ( .A(n3390), .B(p_input[6950]), .Z(o[6950]) );
  AND U6780 ( .A(p_input[26950]), .B(p_input[16950]), .Z(n3390) );
  AND U6781 ( .A(n3391), .B(p_input[694]), .Z(o[694]) );
  AND U6782 ( .A(p_input[20694]), .B(p_input[10694]), .Z(n3391) );
  AND U6783 ( .A(n3392), .B(p_input[6949]), .Z(o[6949]) );
  AND U6784 ( .A(p_input[26949]), .B(p_input[16949]), .Z(n3392) );
  AND U6785 ( .A(n3393), .B(p_input[6948]), .Z(o[6948]) );
  AND U6786 ( .A(p_input[26948]), .B(p_input[16948]), .Z(n3393) );
  AND U6787 ( .A(n3394), .B(p_input[6947]), .Z(o[6947]) );
  AND U6788 ( .A(p_input[26947]), .B(p_input[16947]), .Z(n3394) );
  AND U6789 ( .A(n3395), .B(p_input[6946]), .Z(o[6946]) );
  AND U6790 ( .A(p_input[26946]), .B(p_input[16946]), .Z(n3395) );
  AND U6791 ( .A(n3396), .B(p_input[6945]), .Z(o[6945]) );
  AND U6792 ( .A(p_input[26945]), .B(p_input[16945]), .Z(n3396) );
  AND U6793 ( .A(n3397), .B(p_input[6944]), .Z(o[6944]) );
  AND U6794 ( .A(p_input[26944]), .B(p_input[16944]), .Z(n3397) );
  AND U6795 ( .A(n3398), .B(p_input[6943]), .Z(o[6943]) );
  AND U6796 ( .A(p_input[26943]), .B(p_input[16943]), .Z(n3398) );
  AND U6797 ( .A(n3399), .B(p_input[6942]), .Z(o[6942]) );
  AND U6798 ( .A(p_input[26942]), .B(p_input[16942]), .Z(n3399) );
  AND U6799 ( .A(n3400), .B(p_input[6941]), .Z(o[6941]) );
  AND U6800 ( .A(p_input[26941]), .B(p_input[16941]), .Z(n3400) );
  AND U6801 ( .A(n3401), .B(p_input[6940]), .Z(o[6940]) );
  AND U6802 ( .A(p_input[26940]), .B(p_input[16940]), .Z(n3401) );
  AND U6803 ( .A(n3402), .B(p_input[693]), .Z(o[693]) );
  AND U6804 ( .A(p_input[20693]), .B(p_input[10693]), .Z(n3402) );
  AND U6805 ( .A(n3403), .B(p_input[6939]), .Z(o[6939]) );
  AND U6806 ( .A(p_input[26939]), .B(p_input[16939]), .Z(n3403) );
  AND U6807 ( .A(n3404), .B(p_input[6938]), .Z(o[6938]) );
  AND U6808 ( .A(p_input[26938]), .B(p_input[16938]), .Z(n3404) );
  AND U6809 ( .A(n3405), .B(p_input[6937]), .Z(o[6937]) );
  AND U6810 ( .A(p_input[26937]), .B(p_input[16937]), .Z(n3405) );
  AND U6811 ( .A(n3406), .B(p_input[6936]), .Z(o[6936]) );
  AND U6812 ( .A(p_input[26936]), .B(p_input[16936]), .Z(n3406) );
  AND U6813 ( .A(n3407), .B(p_input[6935]), .Z(o[6935]) );
  AND U6814 ( .A(p_input[26935]), .B(p_input[16935]), .Z(n3407) );
  AND U6815 ( .A(n3408), .B(p_input[6934]), .Z(o[6934]) );
  AND U6816 ( .A(p_input[26934]), .B(p_input[16934]), .Z(n3408) );
  AND U6817 ( .A(n3409), .B(p_input[6933]), .Z(o[6933]) );
  AND U6818 ( .A(p_input[26933]), .B(p_input[16933]), .Z(n3409) );
  AND U6819 ( .A(n3410), .B(p_input[6932]), .Z(o[6932]) );
  AND U6820 ( .A(p_input[26932]), .B(p_input[16932]), .Z(n3410) );
  AND U6821 ( .A(n3411), .B(p_input[6931]), .Z(o[6931]) );
  AND U6822 ( .A(p_input[26931]), .B(p_input[16931]), .Z(n3411) );
  AND U6823 ( .A(n3412), .B(p_input[6930]), .Z(o[6930]) );
  AND U6824 ( .A(p_input[26930]), .B(p_input[16930]), .Z(n3412) );
  AND U6825 ( .A(n3413), .B(p_input[692]), .Z(o[692]) );
  AND U6826 ( .A(p_input[20692]), .B(p_input[10692]), .Z(n3413) );
  AND U6827 ( .A(n3414), .B(p_input[6929]), .Z(o[6929]) );
  AND U6828 ( .A(p_input[26929]), .B(p_input[16929]), .Z(n3414) );
  AND U6829 ( .A(n3415), .B(p_input[6928]), .Z(o[6928]) );
  AND U6830 ( .A(p_input[26928]), .B(p_input[16928]), .Z(n3415) );
  AND U6831 ( .A(n3416), .B(p_input[6927]), .Z(o[6927]) );
  AND U6832 ( .A(p_input[26927]), .B(p_input[16927]), .Z(n3416) );
  AND U6833 ( .A(n3417), .B(p_input[6926]), .Z(o[6926]) );
  AND U6834 ( .A(p_input[26926]), .B(p_input[16926]), .Z(n3417) );
  AND U6835 ( .A(n3418), .B(p_input[6925]), .Z(o[6925]) );
  AND U6836 ( .A(p_input[26925]), .B(p_input[16925]), .Z(n3418) );
  AND U6837 ( .A(n3419), .B(p_input[6924]), .Z(o[6924]) );
  AND U6838 ( .A(p_input[26924]), .B(p_input[16924]), .Z(n3419) );
  AND U6839 ( .A(n3420), .B(p_input[6923]), .Z(o[6923]) );
  AND U6840 ( .A(p_input[26923]), .B(p_input[16923]), .Z(n3420) );
  AND U6841 ( .A(n3421), .B(p_input[6922]), .Z(o[6922]) );
  AND U6842 ( .A(p_input[26922]), .B(p_input[16922]), .Z(n3421) );
  AND U6843 ( .A(n3422), .B(p_input[6921]), .Z(o[6921]) );
  AND U6844 ( .A(p_input[26921]), .B(p_input[16921]), .Z(n3422) );
  AND U6845 ( .A(n3423), .B(p_input[6920]), .Z(o[6920]) );
  AND U6846 ( .A(p_input[26920]), .B(p_input[16920]), .Z(n3423) );
  AND U6847 ( .A(n3424), .B(p_input[691]), .Z(o[691]) );
  AND U6848 ( .A(p_input[20691]), .B(p_input[10691]), .Z(n3424) );
  AND U6849 ( .A(n3425), .B(p_input[6919]), .Z(o[6919]) );
  AND U6850 ( .A(p_input[26919]), .B(p_input[16919]), .Z(n3425) );
  AND U6851 ( .A(n3426), .B(p_input[6918]), .Z(o[6918]) );
  AND U6852 ( .A(p_input[26918]), .B(p_input[16918]), .Z(n3426) );
  AND U6853 ( .A(n3427), .B(p_input[6917]), .Z(o[6917]) );
  AND U6854 ( .A(p_input[26917]), .B(p_input[16917]), .Z(n3427) );
  AND U6855 ( .A(n3428), .B(p_input[6916]), .Z(o[6916]) );
  AND U6856 ( .A(p_input[26916]), .B(p_input[16916]), .Z(n3428) );
  AND U6857 ( .A(n3429), .B(p_input[6915]), .Z(o[6915]) );
  AND U6858 ( .A(p_input[26915]), .B(p_input[16915]), .Z(n3429) );
  AND U6859 ( .A(n3430), .B(p_input[6914]), .Z(o[6914]) );
  AND U6860 ( .A(p_input[26914]), .B(p_input[16914]), .Z(n3430) );
  AND U6861 ( .A(n3431), .B(p_input[6913]), .Z(o[6913]) );
  AND U6862 ( .A(p_input[26913]), .B(p_input[16913]), .Z(n3431) );
  AND U6863 ( .A(n3432), .B(p_input[6912]), .Z(o[6912]) );
  AND U6864 ( .A(p_input[26912]), .B(p_input[16912]), .Z(n3432) );
  AND U6865 ( .A(n3433), .B(p_input[6911]), .Z(o[6911]) );
  AND U6866 ( .A(p_input[26911]), .B(p_input[16911]), .Z(n3433) );
  AND U6867 ( .A(n3434), .B(p_input[6910]), .Z(o[6910]) );
  AND U6868 ( .A(p_input[26910]), .B(p_input[16910]), .Z(n3434) );
  AND U6869 ( .A(n3435), .B(p_input[690]), .Z(o[690]) );
  AND U6870 ( .A(p_input[20690]), .B(p_input[10690]), .Z(n3435) );
  AND U6871 ( .A(n3436), .B(p_input[6909]), .Z(o[6909]) );
  AND U6872 ( .A(p_input[26909]), .B(p_input[16909]), .Z(n3436) );
  AND U6873 ( .A(n3437), .B(p_input[6908]), .Z(o[6908]) );
  AND U6874 ( .A(p_input[26908]), .B(p_input[16908]), .Z(n3437) );
  AND U6875 ( .A(n3438), .B(p_input[6907]), .Z(o[6907]) );
  AND U6876 ( .A(p_input[26907]), .B(p_input[16907]), .Z(n3438) );
  AND U6877 ( .A(n3439), .B(p_input[6906]), .Z(o[6906]) );
  AND U6878 ( .A(p_input[26906]), .B(p_input[16906]), .Z(n3439) );
  AND U6879 ( .A(n3440), .B(p_input[6905]), .Z(o[6905]) );
  AND U6880 ( .A(p_input[26905]), .B(p_input[16905]), .Z(n3440) );
  AND U6881 ( .A(n3441), .B(p_input[6904]), .Z(o[6904]) );
  AND U6882 ( .A(p_input[26904]), .B(p_input[16904]), .Z(n3441) );
  AND U6883 ( .A(n3442), .B(p_input[6903]), .Z(o[6903]) );
  AND U6884 ( .A(p_input[26903]), .B(p_input[16903]), .Z(n3442) );
  AND U6885 ( .A(n3443), .B(p_input[6902]), .Z(o[6902]) );
  AND U6886 ( .A(p_input[26902]), .B(p_input[16902]), .Z(n3443) );
  AND U6887 ( .A(n3444), .B(p_input[6901]), .Z(o[6901]) );
  AND U6888 ( .A(p_input[26901]), .B(p_input[16901]), .Z(n3444) );
  AND U6889 ( .A(n3445), .B(p_input[6900]), .Z(o[6900]) );
  AND U6890 ( .A(p_input[26900]), .B(p_input[16900]), .Z(n3445) );
  AND U6891 ( .A(n3446), .B(p_input[68]), .Z(o[68]) );
  AND U6892 ( .A(p_input[20068]), .B(p_input[10068]), .Z(n3446) );
  AND U6893 ( .A(n3447), .B(p_input[689]), .Z(o[689]) );
  AND U6894 ( .A(p_input[20689]), .B(p_input[10689]), .Z(n3447) );
  AND U6895 ( .A(n3448), .B(p_input[6899]), .Z(o[6899]) );
  AND U6896 ( .A(p_input[26899]), .B(p_input[16899]), .Z(n3448) );
  AND U6897 ( .A(n3449), .B(p_input[6898]), .Z(o[6898]) );
  AND U6898 ( .A(p_input[26898]), .B(p_input[16898]), .Z(n3449) );
  AND U6899 ( .A(n3450), .B(p_input[6897]), .Z(o[6897]) );
  AND U6900 ( .A(p_input[26897]), .B(p_input[16897]), .Z(n3450) );
  AND U6901 ( .A(n3451), .B(p_input[6896]), .Z(o[6896]) );
  AND U6902 ( .A(p_input[26896]), .B(p_input[16896]), .Z(n3451) );
  AND U6903 ( .A(n3452), .B(p_input[6895]), .Z(o[6895]) );
  AND U6904 ( .A(p_input[26895]), .B(p_input[16895]), .Z(n3452) );
  AND U6905 ( .A(n3453), .B(p_input[6894]), .Z(o[6894]) );
  AND U6906 ( .A(p_input[26894]), .B(p_input[16894]), .Z(n3453) );
  AND U6907 ( .A(n3454), .B(p_input[6893]), .Z(o[6893]) );
  AND U6908 ( .A(p_input[26893]), .B(p_input[16893]), .Z(n3454) );
  AND U6909 ( .A(n3455), .B(p_input[6892]), .Z(o[6892]) );
  AND U6910 ( .A(p_input[26892]), .B(p_input[16892]), .Z(n3455) );
  AND U6911 ( .A(n3456), .B(p_input[6891]), .Z(o[6891]) );
  AND U6912 ( .A(p_input[26891]), .B(p_input[16891]), .Z(n3456) );
  AND U6913 ( .A(n3457), .B(p_input[6890]), .Z(o[6890]) );
  AND U6914 ( .A(p_input[26890]), .B(p_input[16890]), .Z(n3457) );
  AND U6915 ( .A(n3458), .B(p_input[688]), .Z(o[688]) );
  AND U6916 ( .A(p_input[20688]), .B(p_input[10688]), .Z(n3458) );
  AND U6917 ( .A(n3459), .B(p_input[6889]), .Z(o[6889]) );
  AND U6918 ( .A(p_input[26889]), .B(p_input[16889]), .Z(n3459) );
  AND U6919 ( .A(n3460), .B(p_input[6888]), .Z(o[6888]) );
  AND U6920 ( .A(p_input[26888]), .B(p_input[16888]), .Z(n3460) );
  AND U6921 ( .A(n3461), .B(p_input[6887]), .Z(o[6887]) );
  AND U6922 ( .A(p_input[26887]), .B(p_input[16887]), .Z(n3461) );
  AND U6923 ( .A(n3462), .B(p_input[6886]), .Z(o[6886]) );
  AND U6924 ( .A(p_input[26886]), .B(p_input[16886]), .Z(n3462) );
  AND U6925 ( .A(n3463), .B(p_input[6885]), .Z(o[6885]) );
  AND U6926 ( .A(p_input[26885]), .B(p_input[16885]), .Z(n3463) );
  AND U6927 ( .A(n3464), .B(p_input[6884]), .Z(o[6884]) );
  AND U6928 ( .A(p_input[26884]), .B(p_input[16884]), .Z(n3464) );
  AND U6929 ( .A(n3465), .B(p_input[6883]), .Z(o[6883]) );
  AND U6930 ( .A(p_input[26883]), .B(p_input[16883]), .Z(n3465) );
  AND U6931 ( .A(n3466), .B(p_input[6882]), .Z(o[6882]) );
  AND U6932 ( .A(p_input[26882]), .B(p_input[16882]), .Z(n3466) );
  AND U6933 ( .A(n3467), .B(p_input[6881]), .Z(o[6881]) );
  AND U6934 ( .A(p_input[26881]), .B(p_input[16881]), .Z(n3467) );
  AND U6935 ( .A(n3468), .B(p_input[6880]), .Z(o[6880]) );
  AND U6936 ( .A(p_input[26880]), .B(p_input[16880]), .Z(n3468) );
  AND U6937 ( .A(n3469), .B(p_input[687]), .Z(o[687]) );
  AND U6938 ( .A(p_input[20687]), .B(p_input[10687]), .Z(n3469) );
  AND U6939 ( .A(n3470), .B(p_input[6879]), .Z(o[6879]) );
  AND U6940 ( .A(p_input[26879]), .B(p_input[16879]), .Z(n3470) );
  AND U6941 ( .A(n3471), .B(p_input[6878]), .Z(o[6878]) );
  AND U6942 ( .A(p_input[26878]), .B(p_input[16878]), .Z(n3471) );
  AND U6943 ( .A(n3472), .B(p_input[6877]), .Z(o[6877]) );
  AND U6944 ( .A(p_input[26877]), .B(p_input[16877]), .Z(n3472) );
  AND U6945 ( .A(n3473), .B(p_input[6876]), .Z(o[6876]) );
  AND U6946 ( .A(p_input[26876]), .B(p_input[16876]), .Z(n3473) );
  AND U6947 ( .A(n3474), .B(p_input[6875]), .Z(o[6875]) );
  AND U6948 ( .A(p_input[26875]), .B(p_input[16875]), .Z(n3474) );
  AND U6949 ( .A(n3475), .B(p_input[6874]), .Z(o[6874]) );
  AND U6950 ( .A(p_input[26874]), .B(p_input[16874]), .Z(n3475) );
  AND U6951 ( .A(n3476), .B(p_input[6873]), .Z(o[6873]) );
  AND U6952 ( .A(p_input[26873]), .B(p_input[16873]), .Z(n3476) );
  AND U6953 ( .A(n3477), .B(p_input[6872]), .Z(o[6872]) );
  AND U6954 ( .A(p_input[26872]), .B(p_input[16872]), .Z(n3477) );
  AND U6955 ( .A(n3478), .B(p_input[6871]), .Z(o[6871]) );
  AND U6956 ( .A(p_input[26871]), .B(p_input[16871]), .Z(n3478) );
  AND U6957 ( .A(n3479), .B(p_input[6870]), .Z(o[6870]) );
  AND U6958 ( .A(p_input[26870]), .B(p_input[16870]), .Z(n3479) );
  AND U6959 ( .A(n3480), .B(p_input[686]), .Z(o[686]) );
  AND U6960 ( .A(p_input[20686]), .B(p_input[10686]), .Z(n3480) );
  AND U6961 ( .A(n3481), .B(p_input[6869]), .Z(o[6869]) );
  AND U6962 ( .A(p_input[26869]), .B(p_input[16869]), .Z(n3481) );
  AND U6963 ( .A(n3482), .B(p_input[6868]), .Z(o[6868]) );
  AND U6964 ( .A(p_input[26868]), .B(p_input[16868]), .Z(n3482) );
  AND U6965 ( .A(n3483), .B(p_input[6867]), .Z(o[6867]) );
  AND U6966 ( .A(p_input[26867]), .B(p_input[16867]), .Z(n3483) );
  AND U6967 ( .A(n3484), .B(p_input[6866]), .Z(o[6866]) );
  AND U6968 ( .A(p_input[26866]), .B(p_input[16866]), .Z(n3484) );
  AND U6969 ( .A(n3485), .B(p_input[6865]), .Z(o[6865]) );
  AND U6970 ( .A(p_input[26865]), .B(p_input[16865]), .Z(n3485) );
  AND U6971 ( .A(n3486), .B(p_input[6864]), .Z(o[6864]) );
  AND U6972 ( .A(p_input[26864]), .B(p_input[16864]), .Z(n3486) );
  AND U6973 ( .A(n3487), .B(p_input[6863]), .Z(o[6863]) );
  AND U6974 ( .A(p_input[26863]), .B(p_input[16863]), .Z(n3487) );
  AND U6975 ( .A(n3488), .B(p_input[6862]), .Z(o[6862]) );
  AND U6976 ( .A(p_input[26862]), .B(p_input[16862]), .Z(n3488) );
  AND U6977 ( .A(n3489), .B(p_input[6861]), .Z(o[6861]) );
  AND U6978 ( .A(p_input[26861]), .B(p_input[16861]), .Z(n3489) );
  AND U6979 ( .A(n3490), .B(p_input[6860]), .Z(o[6860]) );
  AND U6980 ( .A(p_input[26860]), .B(p_input[16860]), .Z(n3490) );
  AND U6981 ( .A(n3491), .B(p_input[685]), .Z(o[685]) );
  AND U6982 ( .A(p_input[20685]), .B(p_input[10685]), .Z(n3491) );
  AND U6983 ( .A(n3492), .B(p_input[6859]), .Z(o[6859]) );
  AND U6984 ( .A(p_input[26859]), .B(p_input[16859]), .Z(n3492) );
  AND U6985 ( .A(n3493), .B(p_input[6858]), .Z(o[6858]) );
  AND U6986 ( .A(p_input[26858]), .B(p_input[16858]), .Z(n3493) );
  AND U6987 ( .A(n3494), .B(p_input[6857]), .Z(o[6857]) );
  AND U6988 ( .A(p_input[26857]), .B(p_input[16857]), .Z(n3494) );
  AND U6989 ( .A(n3495), .B(p_input[6856]), .Z(o[6856]) );
  AND U6990 ( .A(p_input[26856]), .B(p_input[16856]), .Z(n3495) );
  AND U6991 ( .A(n3496), .B(p_input[6855]), .Z(o[6855]) );
  AND U6992 ( .A(p_input[26855]), .B(p_input[16855]), .Z(n3496) );
  AND U6993 ( .A(n3497), .B(p_input[6854]), .Z(o[6854]) );
  AND U6994 ( .A(p_input[26854]), .B(p_input[16854]), .Z(n3497) );
  AND U6995 ( .A(n3498), .B(p_input[6853]), .Z(o[6853]) );
  AND U6996 ( .A(p_input[26853]), .B(p_input[16853]), .Z(n3498) );
  AND U6997 ( .A(n3499), .B(p_input[6852]), .Z(o[6852]) );
  AND U6998 ( .A(p_input[26852]), .B(p_input[16852]), .Z(n3499) );
  AND U6999 ( .A(n3500), .B(p_input[6851]), .Z(o[6851]) );
  AND U7000 ( .A(p_input[26851]), .B(p_input[16851]), .Z(n3500) );
  AND U7001 ( .A(n3501), .B(p_input[6850]), .Z(o[6850]) );
  AND U7002 ( .A(p_input[26850]), .B(p_input[16850]), .Z(n3501) );
  AND U7003 ( .A(n3502), .B(p_input[684]), .Z(o[684]) );
  AND U7004 ( .A(p_input[20684]), .B(p_input[10684]), .Z(n3502) );
  AND U7005 ( .A(n3503), .B(p_input[6849]), .Z(o[6849]) );
  AND U7006 ( .A(p_input[26849]), .B(p_input[16849]), .Z(n3503) );
  AND U7007 ( .A(n3504), .B(p_input[6848]), .Z(o[6848]) );
  AND U7008 ( .A(p_input[26848]), .B(p_input[16848]), .Z(n3504) );
  AND U7009 ( .A(n3505), .B(p_input[6847]), .Z(o[6847]) );
  AND U7010 ( .A(p_input[26847]), .B(p_input[16847]), .Z(n3505) );
  AND U7011 ( .A(n3506), .B(p_input[6846]), .Z(o[6846]) );
  AND U7012 ( .A(p_input[26846]), .B(p_input[16846]), .Z(n3506) );
  AND U7013 ( .A(n3507), .B(p_input[6845]), .Z(o[6845]) );
  AND U7014 ( .A(p_input[26845]), .B(p_input[16845]), .Z(n3507) );
  AND U7015 ( .A(n3508), .B(p_input[6844]), .Z(o[6844]) );
  AND U7016 ( .A(p_input[26844]), .B(p_input[16844]), .Z(n3508) );
  AND U7017 ( .A(n3509), .B(p_input[6843]), .Z(o[6843]) );
  AND U7018 ( .A(p_input[26843]), .B(p_input[16843]), .Z(n3509) );
  AND U7019 ( .A(n3510), .B(p_input[6842]), .Z(o[6842]) );
  AND U7020 ( .A(p_input[26842]), .B(p_input[16842]), .Z(n3510) );
  AND U7021 ( .A(n3511), .B(p_input[6841]), .Z(o[6841]) );
  AND U7022 ( .A(p_input[26841]), .B(p_input[16841]), .Z(n3511) );
  AND U7023 ( .A(n3512), .B(p_input[6840]), .Z(o[6840]) );
  AND U7024 ( .A(p_input[26840]), .B(p_input[16840]), .Z(n3512) );
  AND U7025 ( .A(n3513), .B(p_input[683]), .Z(o[683]) );
  AND U7026 ( .A(p_input[20683]), .B(p_input[10683]), .Z(n3513) );
  AND U7027 ( .A(n3514), .B(p_input[6839]), .Z(o[6839]) );
  AND U7028 ( .A(p_input[26839]), .B(p_input[16839]), .Z(n3514) );
  AND U7029 ( .A(n3515), .B(p_input[6838]), .Z(o[6838]) );
  AND U7030 ( .A(p_input[26838]), .B(p_input[16838]), .Z(n3515) );
  AND U7031 ( .A(n3516), .B(p_input[6837]), .Z(o[6837]) );
  AND U7032 ( .A(p_input[26837]), .B(p_input[16837]), .Z(n3516) );
  AND U7033 ( .A(n3517), .B(p_input[6836]), .Z(o[6836]) );
  AND U7034 ( .A(p_input[26836]), .B(p_input[16836]), .Z(n3517) );
  AND U7035 ( .A(n3518), .B(p_input[6835]), .Z(o[6835]) );
  AND U7036 ( .A(p_input[26835]), .B(p_input[16835]), .Z(n3518) );
  AND U7037 ( .A(n3519), .B(p_input[6834]), .Z(o[6834]) );
  AND U7038 ( .A(p_input[26834]), .B(p_input[16834]), .Z(n3519) );
  AND U7039 ( .A(n3520), .B(p_input[6833]), .Z(o[6833]) );
  AND U7040 ( .A(p_input[26833]), .B(p_input[16833]), .Z(n3520) );
  AND U7041 ( .A(n3521), .B(p_input[6832]), .Z(o[6832]) );
  AND U7042 ( .A(p_input[26832]), .B(p_input[16832]), .Z(n3521) );
  AND U7043 ( .A(n3522), .B(p_input[6831]), .Z(o[6831]) );
  AND U7044 ( .A(p_input[26831]), .B(p_input[16831]), .Z(n3522) );
  AND U7045 ( .A(n3523), .B(p_input[6830]), .Z(o[6830]) );
  AND U7046 ( .A(p_input[26830]), .B(p_input[16830]), .Z(n3523) );
  AND U7047 ( .A(n3524), .B(p_input[682]), .Z(o[682]) );
  AND U7048 ( .A(p_input[20682]), .B(p_input[10682]), .Z(n3524) );
  AND U7049 ( .A(n3525), .B(p_input[6829]), .Z(o[6829]) );
  AND U7050 ( .A(p_input[26829]), .B(p_input[16829]), .Z(n3525) );
  AND U7051 ( .A(n3526), .B(p_input[6828]), .Z(o[6828]) );
  AND U7052 ( .A(p_input[26828]), .B(p_input[16828]), .Z(n3526) );
  AND U7053 ( .A(n3527), .B(p_input[6827]), .Z(o[6827]) );
  AND U7054 ( .A(p_input[26827]), .B(p_input[16827]), .Z(n3527) );
  AND U7055 ( .A(n3528), .B(p_input[6826]), .Z(o[6826]) );
  AND U7056 ( .A(p_input[26826]), .B(p_input[16826]), .Z(n3528) );
  AND U7057 ( .A(n3529), .B(p_input[6825]), .Z(o[6825]) );
  AND U7058 ( .A(p_input[26825]), .B(p_input[16825]), .Z(n3529) );
  AND U7059 ( .A(n3530), .B(p_input[6824]), .Z(o[6824]) );
  AND U7060 ( .A(p_input[26824]), .B(p_input[16824]), .Z(n3530) );
  AND U7061 ( .A(n3531), .B(p_input[6823]), .Z(o[6823]) );
  AND U7062 ( .A(p_input[26823]), .B(p_input[16823]), .Z(n3531) );
  AND U7063 ( .A(n3532), .B(p_input[6822]), .Z(o[6822]) );
  AND U7064 ( .A(p_input[26822]), .B(p_input[16822]), .Z(n3532) );
  AND U7065 ( .A(n3533), .B(p_input[6821]), .Z(o[6821]) );
  AND U7066 ( .A(p_input[26821]), .B(p_input[16821]), .Z(n3533) );
  AND U7067 ( .A(n3534), .B(p_input[6820]), .Z(o[6820]) );
  AND U7068 ( .A(p_input[26820]), .B(p_input[16820]), .Z(n3534) );
  AND U7069 ( .A(n3535), .B(p_input[681]), .Z(o[681]) );
  AND U7070 ( .A(p_input[20681]), .B(p_input[10681]), .Z(n3535) );
  AND U7071 ( .A(n3536), .B(p_input[6819]), .Z(o[6819]) );
  AND U7072 ( .A(p_input[26819]), .B(p_input[16819]), .Z(n3536) );
  AND U7073 ( .A(n3537), .B(p_input[6818]), .Z(o[6818]) );
  AND U7074 ( .A(p_input[26818]), .B(p_input[16818]), .Z(n3537) );
  AND U7075 ( .A(n3538), .B(p_input[6817]), .Z(o[6817]) );
  AND U7076 ( .A(p_input[26817]), .B(p_input[16817]), .Z(n3538) );
  AND U7077 ( .A(n3539), .B(p_input[6816]), .Z(o[6816]) );
  AND U7078 ( .A(p_input[26816]), .B(p_input[16816]), .Z(n3539) );
  AND U7079 ( .A(n3540), .B(p_input[6815]), .Z(o[6815]) );
  AND U7080 ( .A(p_input[26815]), .B(p_input[16815]), .Z(n3540) );
  AND U7081 ( .A(n3541), .B(p_input[6814]), .Z(o[6814]) );
  AND U7082 ( .A(p_input[26814]), .B(p_input[16814]), .Z(n3541) );
  AND U7083 ( .A(n3542), .B(p_input[6813]), .Z(o[6813]) );
  AND U7084 ( .A(p_input[26813]), .B(p_input[16813]), .Z(n3542) );
  AND U7085 ( .A(n3543), .B(p_input[6812]), .Z(o[6812]) );
  AND U7086 ( .A(p_input[26812]), .B(p_input[16812]), .Z(n3543) );
  AND U7087 ( .A(n3544), .B(p_input[6811]), .Z(o[6811]) );
  AND U7088 ( .A(p_input[26811]), .B(p_input[16811]), .Z(n3544) );
  AND U7089 ( .A(n3545), .B(p_input[6810]), .Z(o[6810]) );
  AND U7090 ( .A(p_input[26810]), .B(p_input[16810]), .Z(n3545) );
  AND U7091 ( .A(n3546), .B(p_input[680]), .Z(o[680]) );
  AND U7092 ( .A(p_input[20680]), .B(p_input[10680]), .Z(n3546) );
  AND U7093 ( .A(n3547), .B(p_input[6809]), .Z(o[6809]) );
  AND U7094 ( .A(p_input[26809]), .B(p_input[16809]), .Z(n3547) );
  AND U7095 ( .A(n3548), .B(p_input[6808]), .Z(o[6808]) );
  AND U7096 ( .A(p_input[26808]), .B(p_input[16808]), .Z(n3548) );
  AND U7097 ( .A(n3549), .B(p_input[6807]), .Z(o[6807]) );
  AND U7098 ( .A(p_input[26807]), .B(p_input[16807]), .Z(n3549) );
  AND U7099 ( .A(n3550), .B(p_input[6806]), .Z(o[6806]) );
  AND U7100 ( .A(p_input[26806]), .B(p_input[16806]), .Z(n3550) );
  AND U7101 ( .A(n3551), .B(p_input[6805]), .Z(o[6805]) );
  AND U7102 ( .A(p_input[26805]), .B(p_input[16805]), .Z(n3551) );
  AND U7103 ( .A(n3552), .B(p_input[6804]), .Z(o[6804]) );
  AND U7104 ( .A(p_input[26804]), .B(p_input[16804]), .Z(n3552) );
  AND U7105 ( .A(n3553), .B(p_input[6803]), .Z(o[6803]) );
  AND U7106 ( .A(p_input[26803]), .B(p_input[16803]), .Z(n3553) );
  AND U7107 ( .A(n3554), .B(p_input[6802]), .Z(o[6802]) );
  AND U7108 ( .A(p_input[26802]), .B(p_input[16802]), .Z(n3554) );
  AND U7109 ( .A(n3555), .B(p_input[6801]), .Z(o[6801]) );
  AND U7110 ( .A(p_input[26801]), .B(p_input[16801]), .Z(n3555) );
  AND U7111 ( .A(n3556), .B(p_input[6800]), .Z(o[6800]) );
  AND U7112 ( .A(p_input[26800]), .B(p_input[16800]), .Z(n3556) );
  AND U7113 ( .A(n3557), .B(p_input[67]), .Z(o[67]) );
  AND U7114 ( .A(p_input[20067]), .B(p_input[10067]), .Z(n3557) );
  AND U7115 ( .A(n3558), .B(p_input[679]), .Z(o[679]) );
  AND U7116 ( .A(p_input[20679]), .B(p_input[10679]), .Z(n3558) );
  AND U7117 ( .A(n3559), .B(p_input[6799]), .Z(o[6799]) );
  AND U7118 ( .A(p_input[26799]), .B(p_input[16799]), .Z(n3559) );
  AND U7119 ( .A(n3560), .B(p_input[6798]), .Z(o[6798]) );
  AND U7120 ( .A(p_input[26798]), .B(p_input[16798]), .Z(n3560) );
  AND U7121 ( .A(n3561), .B(p_input[6797]), .Z(o[6797]) );
  AND U7122 ( .A(p_input[26797]), .B(p_input[16797]), .Z(n3561) );
  AND U7123 ( .A(n3562), .B(p_input[6796]), .Z(o[6796]) );
  AND U7124 ( .A(p_input[26796]), .B(p_input[16796]), .Z(n3562) );
  AND U7125 ( .A(n3563), .B(p_input[6795]), .Z(o[6795]) );
  AND U7126 ( .A(p_input[26795]), .B(p_input[16795]), .Z(n3563) );
  AND U7127 ( .A(n3564), .B(p_input[6794]), .Z(o[6794]) );
  AND U7128 ( .A(p_input[26794]), .B(p_input[16794]), .Z(n3564) );
  AND U7129 ( .A(n3565), .B(p_input[6793]), .Z(o[6793]) );
  AND U7130 ( .A(p_input[26793]), .B(p_input[16793]), .Z(n3565) );
  AND U7131 ( .A(n3566), .B(p_input[6792]), .Z(o[6792]) );
  AND U7132 ( .A(p_input[26792]), .B(p_input[16792]), .Z(n3566) );
  AND U7133 ( .A(n3567), .B(p_input[6791]), .Z(o[6791]) );
  AND U7134 ( .A(p_input[26791]), .B(p_input[16791]), .Z(n3567) );
  AND U7135 ( .A(n3568), .B(p_input[6790]), .Z(o[6790]) );
  AND U7136 ( .A(p_input[26790]), .B(p_input[16790]), .Z(n3568) );
  AND U7137 ( .A(n3569), .B(p_input[678]), .Z(o[678]) );
  AND U7138 ( .A(p_input[20678]), .B(p_input[10678]), .Z(n3569) );
  AND U7139 ( .A(n3570), .B(p_input[6789]), .Z(o[6789]) );
  AND U7140 ( .A(p_input[26789]), .B(p_input[16789]), .Z(n3570) );
  AND U7141 ( .A(n3571), .B(p_input[6788]), .Z(o[6788]) );
  AND U7142 ( .A(p_input[26788]), .B(p_input[16788]), .Z(n3571) );
  AND U7143 ( .A(n3572), .B(p_input[6787]), .Z(o[6787]) );
  AND U7144 ( .A(p_input[26787]), .B(p_input[16787]), .Z(n3572) );
  AND U7145 ( .A(n3573), .B(p_input[6786]), .Z(o[6786]) );
  AND U7146 ( .A(p_input[26786]), .B(p_input[16786]), .Z(n3573) );
  AND U7147 ( .A(n3574), .B(p_input[6785]), .Z(o[6785]) );
  AND U7148 ( .A(p_input[26785]), .B(p_input[16785]), .Z(n3574) );
  AND U7149 ( .A(n3575), .B(p_input[6784]), .Z(o[6784]) );
  AND U7150 ( .A(p_input[26784]), .B(p_input[16784]), .Z(n3575) );
  AND U7151 ( .A(n3576), .B(p_input[6783]), .Z(o[6783]) );
  AND U7152 ( .A(p_input[26783]), .B(p_input[16783]), .Z(n3576) );
  AND U7153 ( .A(n3577), .B(p_input[6782]), .Z(o[6782]) );
  AND U7154 ( .A(p_input[26782]), .B(p_input[16782]), .Z(n3577) );
  AND U7155 ( .A(n3578), .B(p_input[6781]), .Z(o[6781]) );
  AND U7156 ( .A(p_input[26781]), .B(p_input[16781]), .Z(n3578) );
  AND U7157 ( .A(n3579), .B(p_input[6780]), .Z(o[6780]) );
  AND U7158 ( .A(p_input[26780]), .B(p_input[16780]), .Z(n3579) );
  AND U7159 ( .A(n3580), .B(p_input[677]), .Z(o[677]) );
  AND U7160 ( .A(p_input[20677]), .B(p_input[10677]), .Z(n3580) );
  AND U7161 ( .A(n3581), .B(p_input[6779]), .Z(o[6779]) );
  AND U7162 ( .A(p_input[26779]), .B(p_input[16779]), .Z(n3581) );
  AND U7163 ( .A(n3582), .B(p_input[6778]), .Z(o[6778]) );
  AND U7164 ( .A(p_input[26778]), .B(p_input[16778]), .Z(n3582) );
  AND U7165 ( .A(n3583), .B(p_input[6777]), .Z(o[6777]) );
  AND U7166 ( .A(p_input[26777]), .B(p_input[16777]), .Z(n3583) );
  AND U7167 ( .A(n3584), .B(p_input[6776]), .Z(o[6776]) );
  AND U7168 ( .A(p_input[26776]), .B(p_input[16776]), .Z(n3584) );
  AND U7169 ( .A(n3585), .B(p_input[6775]), .Z(o[6775]) );
  AND U7170 ( .A(p_input[26775]), .B(p_input[16775]), .Z(n3585) );
  AND U7171 ( .A(n3586), .B(p_input[6774]), .Z(o[6774]) );
  AND U7172 ( .A(p_input[26774]), .B(p_input[16774]), .Z(n3586) );
  AND U7173 ( .A(n3587), .B(p_input[6773]), .Z(o[6773]) );
  AND U7174 ( .A(p_input[26773]), .B(p_input[16773]), .Z(n3587) );
  AND U7175 ( .A(n3588), .B(p_input[6772]), .Z(o[6772]) );
  AND U7176 ( .A(p_input[26772]), .B(p_input[16772]), .Z(n3588) );
  AND U7177 ( .A(n3589), .B(p_input[6771]), .Z(o[6771]) );
  AND U7178 ( .A(p_input[26771]), .B(p_input[16771]), .Z(n3589) );
  AND U7179 ( .A(n3590), .B(p_input[6770]), .Z(o[6770]) );
  AND U7180 ( .A(p_input[26770]), .B(p_input[16770]), .Z(n3590) );
  AND U7181 ( .A(n3591), .B(p_input[676]), .Z(o[676]) );
  AND U7182 ( .A(p_input[20676]), .B(p_input[10676]), .Z(n3591) );
  AND U7183 ( .A(n3592), .B(p_input[6769]), .Z(o[6769]) );
  AND U7184 ( .A(p_input[26769]), .B(p_input[16769]), .Z(n3592) );
  AND U7185 ( .A(n3593), .B(p_input[6768]), .Z(o[6768]) );
  AND U7186 ( .A(p_input[26768]), .B(p_input[16768]), .Z(n3593) );
  AND U7187 ( .A(n3594), .B(p_input[6767]), .Z(o[6767]) );
  AND U7188 ( .A(p_input[26767]), .B(p_input[16767]), .Z(n3594) );
  AND U7189 ( .A(n3595), .B(p_input[6766]), .Z(o[6766]) );
  AND U7190 ( .A(p_input[26766]), .B(p_input[16766]), .Z(n3595) );
  AND U7191 ( .A(n3596), .B(p_input[6765]), .Z(o[6765]) );
  AND U7192 ( .A(p_input[26765]), .B(p_input[16765]), .Z(n3596) );
  AND U7193 ( .A(n3597), .B(p_input[6764]), .Z(o[6764]) );
  AND U7194 ( .A(p_input[26764]), .B(p_input[16764]), .Z(n3597) );
  AND U7195 ( .A(n3598), .B(p_input[6763]), .Z(o[6763]) );
  AND U7196 ( .A(p_input[26763]), .B(p_input[16763]), .Z(n3598) );
  AND U7197 ( .A(n3599), .B(p_input[6762]), .Z(o[6762]) );
  AND U7198 ( .A(p_input[26762]), .B(p_input[16762]), .Z(n3599) );
  AND U7199 ( .A(n3600), .B(p_input[6761]), .Z(o[6761]) );
  AND U7200 ( .A(p_input[26761]), .B(p_input[16761]), .Z(n3600) );
  AND U7201 ( .A(n3601), .B(p_input[6760]), .Z(o[6760]) );
  AND U7202 ( .A(p_input[26760]), .B(p_input[16760]), .Z(n3601) );
  AND U7203 ( .A(n3602), .B(p_input[675]), .Z(o[675]) );
  AND U7204 ( .A(p_input[20675]), .B(p_input[10675]), .Z(n3602) );
  AND U7205 ( .A(n3603), .B(p_input[6759]), .Z(o[6759]) );
  AND U7206 ( .A(p_input[26759]), .B(p_input[16759]), .Z(n3603) );
  AND U7207 ( .A(n3604), .B(p_input[6758]), .Z(o[6758]) );
  AND U7208 ( .A(p_input[26758]), .B(p_input[16758]), .Z(n3604) );
  AND U7209 ( .A(n3605), .B(p_input[6757]), .Z(o[6757]) );
  AND U7210 ( .A(p_input[26757]), .B(p_input[16757]), .Z(n3605) );
  AND U7211 ( .A(n3606), .B(p_input[6756]), .Z(o[6756]) );
  AND U7212 ( .A(p_input[26756]), .B(p_input[16756]), .Z(n3606) );
  AND U7213 ( .A(n3607), .B(p_input[6755]), .Z(o[6755]) );
  AND U7214 ( .A(p_input[26755]), .B(p_input[16755]), .Z(n3607) );
  AND U7215 ( .A(n3608), .B(p_input[6754]), .Z(o[6754]) );
  AND U7216 ( .A(p_input[26754]), .B(p_input[16754]), .Z(n3608) );
  AND U7217 ( .A(n3609), .B(p_input[6753]), .Z(o[6753]) );
  AND U7218 ( .A(p_input[26753]), .B(p_input[16753]), .Z(n3609) );
  AND U7219 ( .A(n3610), .B(p_input[6752]), .Z(o[6752]) );
  AND U7220 ( .A(p_input[26752]), .B(p_input[16752]), .Z(n3610) );
  AND U7221 ( .A(n3611), .B(p_input[6751]), .Z(o[6751]) );
  AND U7222 ( .A(p_input[26751]), .B(p_input[16751]), .Z(n3611) );
  AND U7223 ( .A(n3612), .B(p_input[6750]), .Z(o[6750]) );
  AND U7224 ( .A(p_input[26750]), .B(p_input[16750]), .Z(n3612) );
  AND U7225 ( .A(n3613), .B(p_input[674]), .Z(o[674]) );
  AND U7226 ( .A(p_input[20674]), .B(p_input[10674]), .Z(n3613) );
  AND U7227 ( .A(n3614), .B(p_input[6749]), .Z(o[6749]) );
  AND U7228 ( .A(p_input[26749]), .B(p_input[16749]), .Z(n3614) );
  AND U7229 ( .A(n3615), .B(p_input[6748]), .Z(o[6748]) );
  AND U7230 ( .A(p_input[26748]), .B(p_input[16748]), .Z(n3615) );
  AND U7231 ( .A(n3616), .B(p_input[6747]), .Z(o[6747]) );
  AND U7232 ( .A(p_input[26747]), .B(p_input[16747]), .Z(n3616) );
  AND U7233 ( .A(n3617), .B(p_input[6746]), .Z(o[6746]) );
  AND U7234 ( .A(p_input[26746]), .B(p_input[16746]), .Z(n3617) );
  AND U7235 ( .A(n3618), .B(p_input[6745]), .Z(o[6745]) );
  AND U7236 ( .A(p_input[26745]), .B(p_input[16745]), .Z(n3618) );
  AND U7237 ( .A(n3619), .B(p_input[6744]), .Z(o[6744]) );
  AND U7238 ( .A(p_input[26744]), .B(p_input[16744]), .Z(n3619) );
  AND U7239 ( .A(n3620), .B(p_input[6743]), .Z(o[6743]) );
  AND U7240 ( .A(p_input[26743]), .B(p_input[16743]), .Z(n3620) );
  AND U7241 ( .A(n3621), .B(p_input[6742]), .Z(o[6742]) );
  AND U7242 ( .A(p_input[26742]), .B(p_input[16742]), .Z(n3621) );
  AND U7243 ( .A(n3622), .B(p_input[6741]), .Z(o[6741]) );
  AND U7244 ( .A(p_input[26741]), .B(p_input[16741]), .Z(n3622) );
  AND U7245 ( .A(n3623), .B(p_input[6740]), .Z(o[6740]) );
  AND U7246 ( .A(p_input[26740]), .B(p_input[16740]), .Z(n3623) );
  AND U7247 ( .A(n3624), .B(p_input[673]), .Z(o[673]) );
  AND U7248 ( .A(p_input[20673]), .B(p_input[10673]), .Z(n3624) );
  AND U7249 ( .A(n3625), .B(p_input[6739]), .Z(o[6739]) );
  AND U7250 ( .A(p_input[26739]), .B(p_input[16739]), .Z(n3625) );
  AND U7251 ( .A(n3626), .B(p_input[6738]), .Z(o[6738]) );
  AND U7252 ( .A(p_input[26738]), .B(p_input[16738]), .Z(n3626) );
  AND U7253 ( .A(n3627), .B(p_input[6737]), .Z(o[6737]) );
  AND U7254 ( .A(p_input[26737]), .B(p_input[16737]), .Z(n3627) );
  AND U7255 ( .A(n3628), .B(p_input[6736]), .Z(o[6736]) );
  AND U7256 ( .A(p_input[26736]), .B(p_input[16736]), .Z(n3628) );
  AND U7257 ( .A(n3629), .B(p_input[6735]), .Z(o[6735]) );
  AND U7258 ( .A(p_input[26735]), .B(p_input[16735]), .Z(n3629) );
  AND U7259 ( .A(n3630), .B(p_input[6734]), .Z(o[6734]) );
  AND U7260 ( .A(p_input[26734]), .B(p_input[16734]), .Z(n3630) );
  AND U7261 ( .A(n3631), .B(p_input[6733]), .Z(o[6733]) );
  AND U7262 ( .A(p_input[26733]), .B(p_input[16733]), .Z(n3631) );
  AND U7263 ( .A(n3632), .B(p_input[6732]), .Z(o[6732]) );
  AND U7264 ( .A(p_input[26732]), .B(p_input[16732]), .Z(n3632) );
  AND U7265 ( .A(n3633), .B(p_input[6731]), .Z(o[6731]) );
  AND U7266 ( .A(p_input[26731]), .B(p_input[16731]), .Z(n3633) );
  AND U7267 ( .A(n3634), .B(p_input[6730]), .Z(o[6730]) );
  AND U7268 ( .A(p_input[26730]), .B(p_input[16730]), .Z(n3634) );
  AND U7269 ( .A(n3635), .B(p_input[672]), .Z(o[672]) );
  AND U7270 ( .A(p_input[20672]), .B(p_input[10672]), .Z(n3635) );
  AND U7271 ( .A(n3636), .B(p_input[6729]), .Z(o[6729]) );
  AND U7272 ( .A(p_input[26729]), .B(p_input[16729]), .Z(n3636) );
  AND U7273 ( .A(n3637), .B(p_input[6728]), .Z(o[6728]) );
  AND U7274 ( .A(p_input[26728]), .B(p_input[16728]), .Z(n3637) );
  AND U7275 ( .A(n3638), .B(p_input[6727]), .Z(o[6727]) );
  AND U7276 ( .A(p_input[26727]), .B(p_input[16727]), .Z(n3638) );
  AND U7277 ( .A(n3639), .B(p_input[6726]), .Z(o[6726]) );
  AND U7278 ( .A(p_input[26726]), .B(p_input[16726]), .Z(n3639) );
  AND U7279 ( .A(n3640), .B(p_input[6725]), .Z(o[6725]) );
  AND U7280 ( .A(p_input[26725]), .B(p_input[16725]), .Z(n3640) );
  AND U7281 ( .A(n3641), .B(p_input[6724]), .Z(o[6724]) );
  AND U7282 ( .A(p_input[26724]), .B(p_input[16724]), .Z(n3641) );
  AND U7283 ( .A(n3642), .B(p_input[6723]), .Z(o[6723]) );
  AND U7284 ( .A(p_input[26723]), .B(p_input[16723]), .Z(n3642) );
  AND U7285 ( .A(n3643), .B(p_input[6722]), .Z(o[6722]) );
  AND U7286 ( .A(p_input[26722]), .B(p_input[16722]), .Z(n3643) );
  AND U7287 ( .A(n3644), .B(p_input[6721]), .Z(o[6721]) );
  AND U7288 ( .A(p_input[26721]), .B(p_input[16721]), .Z(n3644) );
  AND U7289 ( .A(n3645), .B(p_input[6720]), .Z(o[6720]) );
  AND U7290 ( .A(p_input[26720]), .B(p_input[16720]), .Z(n3645) );
  AND U7291 ( .A(n3646), .B(p_input[671]), .Z(o[671]) );
  AND U7292 ( .A(p_input[20671]), .B(p_input[10671]), .Z(n3646) );
  AND U7293 ( .A(n3647), .B(p_input[6719]), .Z(o[6719]) );
  AND U7294 ( .A(p_input[26719]), .B(p_input[16719]), .Z(n3647) );
  AND U7295 ( .A(n3648), .B(p_input[6718]), .Z(o[6718]) );
  AND U7296 ( .A(p_input[26718]), .B(p_input[16718]), .Z(n3648) );
  AND U7297 ( .A(n3649), .B(p_input[6717]), .Z(o[6717]) );
  AND U7298 ( .A(p_input[26717]), .B(p_input[16717]), .Z(n3649) );
  AND U7299 ( .A(n3650), .B(p_input[6716]), .Z(o[6716]) );
  AND U7300 ( .A(p_input[26716]), .B(p_input[16716]), .Z(n3650) );
  AND U7301 ( .A(n3651), .B(p_input[6715]), .Z(o[6715]) );
  AND U7302 ( .A(p_input[26715]), .B(p_input[16715]), .Z(n3651) );
  AND U7303 ( .A(n3652), .B(p_input[6714]), .Z(o[6714]) );
  AND U7304 ( .A(p_input[26714]), .B(p_input[16714]), .Z(n3652) );
  AND U7305 ( .A(n3653), .B(p_input[6713]), .Z(o[6713]) );
  AND U7306 ( .A(p_input[26713]), .B(p_input[16713]), .Z(n3653) );
  AND U7307 ( .A(n3654), .B(p_input[6712]), .Z(o[6712]) );
  AND U7308 ( .A(p_input[26712]), .B(p_input[16712]), .Z(n3654) );
  AND U7309 ( .A(n3655), .B(p_input[6711]), .Z(o[6711]) );
  AND U7310 ( .A(p_input[26711]), .B(p_input[16711]), .Z(n3655) );
  AND U7311 ( .A(n3656), .B(p_input[6710]), .Z(o[6710]) );
  AND U7312 ( .A(p_input[26710]), .B(p_input[16710]), .Z(n3656) );
  AND U7313 ( .A(n3657), .B(p_input[670]), .Z(o[670]) );
  AND U7314 ( .A(p_input[20670]), .B(p_input[10670]), .Z(n3657) );
  AND U7315 ( .A(n3658), .B(p_input[6709]), .Z(o[6709]) );
  AND U7316 ( .A(p_input[26709]), .B(p_input[16709]), .Z(n3658) );
  AND U7317 ( .A(n3659), .B(p_input[6708]), .Z(o[6708]) );
  AND U7318 ( .A(p_input[26708]), .B(p_input[16708]), .Z(n3659) );
  AND U7319 ( .A(n3660), .B(p_input[6707]), .Z(o[6707]) );
  AND U7320 ( .A(p_input[26707]), .B(p_input[16707]), .Z(n3660) );
  AND U7321 ( .A(n3661), .B(p_input[6706]), .Z(o[6706]) );
  AND U7322 ( .A(p_input[26706]), .B(p_input[16706]), .Z(n3661) );
  AND U7323 ( .A(n3662), .B(p_input[6705]), .Z(o[6705]) );
  AND U7324 ( .A(p_input[26705]), .B(p_input[16705]), .Z(n3662) );
  AND U7325 ( .A(n3663), .B(p_input[6704]), .Z(o[6704]) );
  AND U7326 ( .A(p_input[26704]), .B(p_input[16704]), .Z(n3663) );
  AND U7327 ( .A(n3664), .B(p_input[6703]), .Z(o[6703]) );
  AND U7328 ( .A(p_input[26703]), .B(p_input[16703]), .Z(n3664) );
  AND U7329 ( .A(n3665), .B(p_input[6702]), .Z(o[6702]) );
  AND U7330 ( .A(p_input[26702]), .B(p_input[16702]), .Z(n3665) );
  AND U7331 ( .A(n3666), .B(p_input[6701]), .Z(o[6701]) );
  AND U7332 ( .A(p_input[26701]), .B(p_input[16701]), .Z(n3666) );
  AND U7333 ( .A(n3667), .B(p_input[6700]), .Z(o[6700]) );
  AND U7334 ( .A(p_input[26700]), .B(p_input[16700]), .Z(n3667) );
  AND U7335 ( .A(n3668), .B(p_input[66]), .Z(o[66]) );
  AND U7336 ( .A(p_input[20066]), .B(p_input[10066]), .Z(n3668) );
  AND U7337 ( .A(n3669), .B(p_input[669]), .Z(o[669]) );
  AND U7338 ( .A(p_input[20669]), .B(p_input[10669]), .Z(n3669) );
  AND U7339 ( .A(n3670), .B(p_input[6699]), .Z(o[6699]) );
  AND U7340 ( .A(p_input[26699]), .B(p_input[16699]), .Z(n3670) );
  AND U7341 ( .A(n3671), .B(p_input[6698]), .Z(o[6698]) );
  AND U7342 ( .A(p_input[26698]), .B(p_input[16698]), .Z(n3671) );
  AND U7343 ( .A(n3672), .B(p_input[6697]), .Z(o[6697]) );
  AND U7344 ( .A(p_input[26697]), .B(p_input[16697]), .Z(n3672) );
  AND U7345 ( .A(n3673), .B(p_input[6696]), .Z(o[6696]) );
  AND U7346 ( .A(p_input[26696]), .B(p_input[16696]), .Z(n3673) );
  AND U7347 ( .A(n3674), .B(p_input[6695]), .Z(o[6695]) );
  AND U7348 ( .A(p_input[26695]), .B(p_input[16695]), .Z(n3674) );
  AND U7349 ( .A(n3675), .B(p_input[6694]), .Z(o[6694]) );
  AND U7350 ( .A(p_input[26694]), .B(p_input[16694]), .Z(n3675) );
  AND U7351 ( .A(n3676), .B(p_input[6693]), .Z(o[6693]) );
  AND U7352 ( .A(p_input[26693]), .B(p_input[16693]), .Z(n3676) );
  AND U7353 ( .A(n3677), .B(p_input[6692]), .Z(o[6692]) );
  AND U7354 ( .A(p_input[26692]), .B(p_input[16692]), .Z(n3677) );
  AND U7355 ( .A(n3678), .B(p_input[6691]), .Z(o[6691]) );
  AND U7356 ( .A(p_input[26691]), .B(p_input[16691]), .Z(n3678) );
  AND U7357 ( .A(n3679), .B(p_input[6690]), .Z(o[6690]) );
  AND U7358 ( .A(p_input[26690]), .B(p_input[16690]), .Z(n3679) );
  AND U7359 ( .A(n3680), .B(p_input[668]), .Z(o[668]) );
  AND U7360 ( .A(p_input[20668]), .B(p_input[10668]), .Z(n3680) );
  AND U7361 ( .A(n3681), .B(p_input[6689]), .Z(o[6689]) );
  AND U7362 ( .A(p_input[26689]), .B(p_input[16689]), .Z(n3681) );
  AND U7363 ( .A(n3682), .B(p_input[6688]), .Z(o[6688]) );
  AND U7364 ( .A(p_input[26688]), .B(p_input[16688]), .Z(n3682) );
  AND U7365 ( .A(n3683), .B(p_input[6687]), .Z(o[6687]) );
  AND U7366 ( .A(p_input[26687]), .B(p_input[16687]), .Z(n3683) );
  AND U7367 ( .A(n3684), .B(p_input[6686]), .Z(o[6686]) );
  AND U7368 ( .A(p_input[26686]), .B(p_input[16686]), .Z(n3684) );
  AND U7369 ( .A(n3685), .B(p_input[6685]), .Z(o[6685]) );
  AND U7370 ( .A(p_input[26685]), .B(p_input[16685]), .Z(n3685) );
  AND U7371 ( .A(n3686), .B(p_input[6684]), .Z(o[6684]) );
  AND U7372 ( .A(p_input[26684]), .B(p_input[16684]), .Z(n3686) );
  AND U7373 ( .A(n3687), .B(p_input[6683]), .Z(o[6683]) );
  AND U7374 ( .A(p_input[26683]), .B(p_input[16683]), .Z(n3687) );
  AND U7375 ( .A(n3688), .B(p_input[6682]), .Z(o[6682]) );
  AND U7376 ( .A(p_input[26682]), .B(p_input[16682]), .Z(n3688) );
  AND U7377 ( .A(n3689), .B(p_input[6681]), .Z(o[6681]) );
  AND U7378 ( .A(p_input[26681]), .B(p_input[16681]), .Z(n3689) );
  AND U7379 ( .A(n3690), .B(p_input[6680]), .Z(o[6680]) );
  AND U7380 ( .A(p_input[26680]), .B(p_input[16680]), .Z(n3690) );
  AND U7381 ( .A(n3691), .B(p_input[667]), .Z(o[667]) );
  AND U7382 ( .A(p_input[20667]), .B(p_input[10667]), .Z(n3691) );
  AND U7383 ( .A(n3692), .B(p_input[6679]), .Z(o[6679]) );
  AND U7384 ( .A(p_input[26679]), .B(p_input[16679]), .Z(n3692) );
  AND U7385 ( .A(n3693), .B(p_input[6678]), .Z(o[6678]) );
  AND U7386 ( .A(p_input[26678]), .B(p_input[16678]), .Z(n3693) );
  AND U7387 ( .A(n3694), .B(p_input[6677]), .Z(o[6677]) );
  AND U7388 ( .A(p_input[26677]), .B(p_input[16677]), .Z(n3694) );
  AND U7389 ( .A(n3695), .B(p_input[6676]), .Z(o[6676]) );
  AND U7390 ( .A(p_input[26676]), .B(p_input[16676]), .Z(n3695) );
  AND U7391 ( .A(n3696), .B(p_input[6675]), .Z(o[6675]) );
  AND U7392 ( .A(p_input[26675]), .B(p_input[16675]), .Z(n3696) );
  AND U7393 ( .A(n3697), .B(p_input[6674]), .Z(o[6674]) );
  AND U7394 ( .A(p_input[26674]), .B(p_input[16674]), .Z(n3697) );
  AND U7395 ( .A(n3698), .B(p_input[6673]), .Z(o[6673]) );
  AND U7396 ( .A(p_input[26673]), .B(p_input[16673]), .Z(n3698) );
  AND U7397 ( .A(n3699), .B(p_input[6672]), .Z(o[6672]) );
  AND U7398 ( .A(p_input[26672]), .B(p_input[16672]), .Z(n3699) );
  AND U7399 ( .A(n3700), .B(p_input[6671]), .Z(o[6671]) );
  AND U7400 ( .A(p_input[26671]), .B(p_input[16671]), .Z(n3700) );
  AND U7401 ( .A(n3701), .B(p_input[6670]), .Z(o[6670]) );
  AND U7402 ( .A(p_input[26670]), .B(p_input[16670]), .Z(n3701) );
  AND U7403 ( .A(n3702), .B(p_input[666]), .Z(o[666]) );
  AND U7404 ( .A(p_input[20666]), .B(p_input[10666]), .Z(n3702) );
  AND U7405 ( .A(n3703), .B(p_input[6669]), .Z(o[6669]) );
  AND U7406 ( .A(p_input[26669]), .B(p_input[16669]), .Z(n3703) );
  AND U7407 ( .A(n3704), .B(p_input[6668]), .Z(o[6668]) );
  AND U7408 ( .A(p_input[26668]), .B(p_input[16668]), .Z(n3704) );
  AND U7409 ( .A(n3705), .B(p_input[6667]), .Z(o[6667]) );
  AND U7410 ( .A(p_input[26667]), .B(p_input[16667]), .Z(n3705) );
  AND U7411 ( .A(n3706), .B(p_input[6666]), .Z(o[6666]) );
  AND U7412 ( .A(p_input[26666]), .B(p_input[16666]), .Z(n3706) );
  AND U7413 ( .A(n3707), .B(p_input[6665]), .Z(o[6665]) );
  AND U7414 ( .A(p_input[26665]), .B(p_input[16665]), .Z(n3707) );
  AND U7415 ( .A(n3708), .B(p_input[6664]), .Z(o[6664]) );
  AND U7416 ( .A(p_input[26664]), .B(p_input[16664]), .Z(n3708) );
  AND U7417 ( .A(n3709), .B(p_input[6663]), .Z(o[6663]) );
  AND U7418 ( .A(p_input[26663]), .B(p_input[16663]), .Z(n3709) );
  AND U7419 ( .A(n3710), .B(p_input[6662]), .Z(o[6662]) );
  AND U7420 ( .A(p_input[26662]), .B(p_input[16662]), .Z(n3710) );
  AND U7421 ( .A(n3711), .B(p_input[6661]), .Z(o[6661]) );
  AND U7422 ( .A(p_input[26661]), .B(p_input[16661]), .Z(n3711) );
  AND U7423 ( .A(n3712), .B(p_input[6660]), .Z(o[6660]) );
  AND U7424 ( .A(p_input[26660]), .B(p_input[16660]), .Z(n3712) );
  AND U7425 ( .A(n3713), .B(p_input[665]), .Z(o[665]) );
  AND U7426 ( .A(p_input[20665]), .B(p_input[10665]), .Z(n3713) );
  AND U7427 ( .A(n3714), .B(p_input[6659]), .Z(o[6659]) );
  AND U7428 ( .A(p_input[26659]), .B(p_input[16659]), .Z(n3714) );
  AND U7429 ( .A(n3715), .B(p_input[6658]), .Z(o[6658]) );
  AND U7430 ( .A(p_input[26658]), .B(p_input[16658]), .Z(n3715) );
  AND U7431 ( .A(n3716), .B(p_input[6657]), .Z(o[6657]) );
  AND U7432 ( .A(p_input[26657]), .B(p_input[16657]), .Z(n3716) );
  AND U7433 ( .A(n3717), .B(p_input[6656]), .Z(o[6656]) );
  AND U7434 ( .A(p_input[26656]), .B(p_input[16656]), .Z(n3717) );
  AND U7435 ( .A(n3718), .B(p_input[6655]), .Z(o[6655]) );
  AND U7436 ( .A(p_input[26655]), .B(p_input[16655]), .Z(n3718) );
  AND U7437 ( .A(n3719), .B(p_input[6654]), .Z(o[6654]) );
  AND U7438 ( .A(p_input[26654]), .B(p_input[16654]), .Z(n3719) );
  AND U7439 ( .A(n3720), .B(p_input[6653]), .Z(o[6653]) );
  AND U7440 ( .A(p_input[26653]), .B(p_input[16653]), .Z(n3720) );
  AND U7441 ( .A(n3721), .B(p_input[6652]), .Z(o[6652]) );
  AND U7442 ( .A(p_input[26652]), .B(p_input[16652]), .Z(n3721) );
  AND U7443 ( .A(n3722), .B(p_input[6651]), .Z(o[6651]) );
  AND U7444 ( .A(p_input[26651]), .B(p_input[16651]), .Z(n3722) );
  AND U7445 ( .A(n3723), .B(p_input[6650]), .Z(o[6650]) );
  AND U7446 ( .A(p_input[26650]), .B(p_input[16650]), .Z(n3723) );
  AND U7447 ( .A(n3724), .B(p_input[664]), .Z(o[664]) );
  AND U7448 ( .A(p_input[20664]), .B(p_input[10664]), .Z(n3724) );
  AND U7449 ( .A(n3725), .B(p_input[6649]), .Z(o[6649]) );
  AND U7450 ( .A(p_input[26649]), .B(p_input[16649]), .Z(n3725) );
  AND U7451 ( .A(n3726), .B(p_input[6648]), .Z(o[6648]) );
  AND U7452 ( .A(p_input[26648]), .B(p_input[16648]), .Z(n3726) );
  AND U7453 ( .A(n3727), .B(p_input[6647]), .Z(o[6647]) );
  AND U7454 ( .A(p_input[26647]), .B(p_input[16647]), .Z(n3727) );
  AND U7455 ( .A(n3728), .B(p_input[6646]), .Z(o[6646]) );
  AND U7456 ( .A(p_input[26646]), .B(p_input[16646]), .Z(n3728) );
  AND U7457 ( .A(n3729), .B(p_input[6645]), .Z(o[6645]) );
  AND U7458 ( .A(p_input[26645]), .B(p_input[16645]), .Z(n3729) );
  AND U7459 ( .A(n3730), .B(p_input[6644]), .Z(o[6644]) );
  AND U7460 ( .A(p_input[26644]), .B(p_input[16644]), .Z(n3730) );
  AND U7461 ( .A(n3731), .B(p_input[6643]), .Z(o[6643]) );
  AND U7462 ( .A(p_input[26643]), .B(p_input[16643]), .Z(n3731) );
  AND U7463 ( .A(n3732), .B(p_input[6642]), .Z(o[6642]) );
  AND U7464 ( .A(p_input[26642]), .B(p_input[16642]), .Z(n3732) );
  AND U7465 ( .A(n3733), .B(p_input[6641]), .Z(o[6641]) );
  AND U7466 ( .A(p_input[26641]), .B(p_input[16641]), .Z(n3733) );
  AND U7467 ( .A(n3734), .B(p_input[6640]), .Z(o[6640]) );
  AND U7468 ( .A(p_input[26640]), .B(p_input[16640]), .Z(n3734) );
  AND U7469 ( .A(n3735), .B(p_input[663]), .Z(o[663]) );
  AND U7470 ( .A(p_input[20663]), .B(p_input[10663]), .Z(n3735) );
  AND U7471 ( .A(n3736), .B(p_input[6639]), .Z(o[6639]) );
  AND U7472 ( .A(p_input[26639]), .B(p_input[16639]), .Z(n3736) );
  AND U7473 ( .A(n3737), .B(p_input[6638]), .Z(o[6638]) );
  AND U7474 ( .A(p_input[26638]), .B(p_input[16638]), .Z(n3737) );
  AND U7475 ( .A(n3738), .B(p_input[6637]), .Z(o[6637]) );
  AND U7476 ( .A(p_input[26637]), .B(p_input[16637]), .Z(n3738) );
  AND U7477 ( .A(n3739), .B(p_input[6636]), .Z(o[6636]) );
  AND U7478 ( .A(p_input[26636]), .B(p_input[16636]), .Z(n3739) );
  AND U7479 ( .A(n3740), .B(p_input[6635]), .Z(o[6635]) );
  AND U7480 ( .A(p_input[26635]), .B(p_input[16635]), .Z(n3740) );
  AND U7481 ( .A(n3741), .B(p_input[6634]), .Z(o[6634]) );
  AND U7482 ( .A(p_input[26634]), .B(p_input[16634]), .Z(n3741) );
  AND U7483 ( .A(n3742), .B(p_input[6633]), .Z(o[6633]) );
  AND U7484 ( .A(p_input[26633]), .B(p_input[16633]), .Z(n3742) );
  AND U7485 ( .A(n3743), .B(p_input[6632]), .Z(o[6632]) );
  AND U7486 ( .A(p_input[26632]), .B(p_input[16632]), .Z(n3743) );
  AND U7487 ( .A(n3744), .B(p_input[6631]), .Z(o[6631]) );
  AND U7488 ( .A(p_input[26631]), .B(p_input[16631]), .Z(n3744) );
  AND U7489 ( .A(n3745), .B(p_input[6630]), .Z(o[6630]) );
  AND U7490 ( .A(p_input[26630]), .B(p_input[16630]), .Z(n3745) );
  AND U7491 ( .A(n3746), .B(p_input[662]), .Z(o[662]) );
  AND U7492 ( .A(p_input[20662]), .B(p_input[10662]), .Z(n3746) );
  AND U7493 ( .A(n3747), .B(p_input[6629]), .Z(o[6629]) );
  AND U7494 ( .A(p_input[26629]), .B(p_input[16629]), .Z(n3747) );
  AND U7495 ( .A(n3748), .B(p_input[6628]), .Z(o[6628]) );
  AND U7496 ( .A(p_input[26628]), .B(p_input[16628]), .Z(n3748) );
  AND U7497 ( .A(n3749), .B(p_input[6627]), .Z(o[6627]) );
  AND U7498 ( .A(p_input[26627]), .B(p_input[16627]), .Z(n3749) );
  AND U7499 ( .A(n3750), .B(p_input[6626]), .Z(o[6626]) );
  AND U7500 ( .A(p_input[26626]), .B(p_input[16626]), .Z(n3750) );
  AND U7501 ( .A(n3751), .B(p_input[6625]), .Z(o[6625]) );
  AND U7502 ( .A(p_input[26625]), .B(p_input[16625]), .Z(n3751) );
  AND U7503 ( .A(n3752), .B(p_input[6624]), .Z(o[6624]) );
  AND U7504 ( .A(p_input[26624]), .B(p_input[16624]), .Z(n3752) );
  AND U7505 ( .A(n3753), .B(p_input[6623]), .Z(o[6623]) );
  AND U7506 ( .A(p_input[26623]), .B(p_input[16623]), .Z(n3753) );
  AND U7507 ( .A(n3754), .B(p_input[6622]), .Z(o[6622]) );
  AND U7508 ( .A(p_input[26622]), .B(p_input[16622]), .Z(n3754) );
  AND U7509 ( .A(n3755), .B(p_input[6621]), .Z(o[6621]) );
  AND U7510 ( .A(p_input[26621]), .B(p_input[16621]), .Z(n3755) );
  AND U7511 ( .A(n3756), .B(p_input[6620]), .Z(o[6620]) );
  AND U7512 ( .A(p_input[26620]), .B(p_input[16620]), .Z(n3756) );
  AND U7513 ( .A(n3757), .B(p_input[661]), .Z(o[661]) );
  AND U7514 ( .A(p_input[20661]), .B(p_input[10661]), .Z(n3757) );
  AND U7515 ( .A(n3758), .B(p_input[6619]), .Z(o[6619]) );
  AND U7516 ( .A(p_input[26619]), .B(p_input[16619]), .Z(n3758) );
  AND U7517 ( .A(n3759), .B(p_input[6618]), .Z(o[6618]) );
  AND U7518 ( .A(p_input[26618]), .B(p_input[16618]), .Z(n3759) );
  AND U7519 ( .A(n3760), .B(p_input[6617]), .Z(o[6617]) );
  AND U7520 ( .A(p_input[26617]), .B(p_input[16617]), .Z(n3760) );
  AND U7521 ( .A(n3761), .B(p_input[6616]), .Z(o[6616]) );
  AND U7522 ( .A(p_input[26616]), .B(p_input[16616]), .Z(n3761) );
  AND U7523 ( .A(n3762), .B(p_input[6615]), .Z(o[6615]) );
  AND U7524 ( .A(p_input[26615]), .B(p_input[16615]), .Z(n3762) );
  AND U7525 ( .A(n3763), .B(p_input[6614]), .Z(o[6614]) );
  AND U7526 ( .A(p_input[26614]), .B(p_input[16614]), .Z(n3763) );
  AND U7527 ( .A(n3764), .B(p_input[6613]), .Z(o[6613]) );
  AND U7528 ( .A(p_input[26613]), .B(p_input[16613]), .Z(n3764) );
  AND U7529 ( .A(n3765), .B(p_input[6612]), .Z(o[6612]) );
  AND U7530 ( .A(p_input[26612]), .B(p_input[16612]), .Z(n3765) );
  AND U7531 ( .A(n3766), .B(p_input[6611]), .Z(o[6611]) );
  AND U7532 ( .A(p_input[26611]), .B(p_input[16611]), .Z(n3766) );
  AND U7533 ( .A(n3767), .B(p_input[6610]), .Z(o[6610]) );
  AND U7534 ( .A(p_input[26610]), .B(p_input[16610]), .Z(n3767) );
  AND U7535 ( .A(n3768), .B(p_input[660]), .Z(o[660]) );
  AND U7536 ( .A(p_input[20660]), .B(p_input[10660]), .Z(n3768) );
  AND U7537 ( .A(n3769), .B(p_input[6609]), .Z(o[6609]) );
  AND U7538 ( .A(p_input[26609]), .B(p_input[16609]), .Z(n3769) );
  AND U7539 ( .A(n3770), .B(p_input[6608]), .Z(o[6608]) );
  AND U7540 ( .A(p_input[26608]), .B(p_input[16608]), .Z(n3770) );
  AND U7541 ( .A(n3771), .B(p_input[6607]), .Z(o[6607]) );
  AND U7542 ( .A(p_input[26607]), .B(p_input[16607]), .Z(n3771) );
  AND U7543 ( .A(n3772), .B(p_input[6606]), .Z(o[6606]) );
  AND U7544 ( .A(p_input[26606]), .B(p_input[16606]), .Z(n3772) );
  AND U7545 ( .A(n3773), .B(p_input[6605]), .Z(o[6605]) );
  AND U7546 ( .A(p_input[26605]), .B(p_input[16605]), .Z(n3773) );
  AND U7547 ( .A(n3774), .B(p_input[6604]), .Z(o[6604]) );
  AND U7548 ( .A(p_input[26604]), .B(p_input[16604]), .Z(n3774) );
  AND U7549 ( .A(n3775), .B(p_input[6603]), .Z(o[6603]) );
  AND U7550 ( .A(p_input[26603]), .B(p_input[16603]), .Z(n3775) );
  AND U7551 ( .A(n3776), .B(p_input[6602]), .Z(o[6602]) );
  AND U7552 ( .A(p_input[26602]), .B(p_input[16602]), .Z(n3776) );
  AND U7553 ( .A(n3777), .B(p_input[6601]), .Z(o[6601]) );
  AND U7554 ( .A(p_input[26601]), .B(p_input[16601]), .Z(n3777) );
  AND U7555 ( .A(n3778), .B(p_input[6600]), .Z(o[6600]) );
  AND U7556 ( .A(p_input[26600]), .B(p_input[16600]), .Z(n3778) );
  AND U7557 ( .A(n3779), .B(p_input[65]), .Z(o[65]) );
  AND U7558 ( .A(p_input[20065]), .B(p_input[10065]), .Z(n3779) );
  AND U7559 ( .A(n3780), .B(p_input[659]), .Z(o[659]) );
  AND U7560 ( .A(p_input[20659]), .B(p_input[10659]), .Z(n3780) );
  AND U7561 ( .A(n3781), .B(p_input[6599]), .Z(o[6599]) );
  AND U7562 ( .A(p_input[26599]), .B(p_input[16599]), .Z(n3781) );
  AND U7563 ( .A(n3782), .B(p_input[6598]), .Z(o[6598]) );
  AND U7564 ( .A(p_input[26598]), .B(p_input[16598]), .Z(n3782) );
  AND U7565 ( .A(n3783), .B(p_input[6597]), .Z(o[6597]) );
  AND U7566 ( .A(p_input[26597]), .B(p_input[16597]), .Z(n3783) );
  AND U7567 ( .A(n3784), .B(p_input[6596]), .Z(o[6596]) );
  AND U7568 ( .A(p_input[26596]), .B(p_input[16596]), .Z(n3784) );
  AND U7569 ( .A(n3785), .B(p_input[6595]), .Z(o[6595]) );
  AND U7570 ( .A(p_input[26595]), .B(p_input[16595]), .Z(n3785) );
  AND U7571 ( .A(n3786), .B(p_input[6594]), .Z(o[6594]) );
  AND U7572 ( .A(p_input[26594]), .B(p_input[16594]), .Z(n3786) );
  AND U7573 ( .A(n3787), .B(p_input[6593]), .Z(o[6593]) );
  AND U7574 ( .A(p_input[26593]), .B(p_input[16593]), .Z(n3787) );
  AND U7575 ( .A(n3788), .B(p_input[6592]), .Z(o[6592]) );
  AND U7576 ( .A(p_input[26592]), .B(p_input[16592]), .Z(n3788) );
  AND U7577 ( .A(n3789), .B(p_input[6591]), .Z(o[6591]) );
  AND U7578 ( .A(p_input[26591]), .B(p_input[16591]), .Z(n3789) );
  AND U7579 ( .A(n3790), .B(p_input[6590]), .Z(o[6590]) );
  AND U7580 ( .A(p_input[26590]), .B(p_input[16590]), .Z(n3790) );
  AND U7581 ( .A(n3791), .B(p_input[658]), .Z(o[658]) );
  AND U7582 ( .A(p_input[20658]), .B(p_input[10658]), .Z(n3791) );
  AND U7583 ( .A(n3792), .B(p_input[6589]), .Z(o[6589]) );
  AND U7584 ( .A(p_input[26589]), .B(p_input[16589]), .Z(n3792) );
  AND U7585 ( .A(n3793), .B(p_input[6588]), .Z(o[6588]) );
  AND U7586 ( .A(p_input[26588]), .B(p_input[16588]), .Z(n3793) );
  AND U7587 ( .A(n3794), .B(p_input[6587]), .Z(o[6587]) );
  AND U7588 ( .A(p_input[26587]), .B(p_input[16587]), .Z(n3794) );
  AND U7589 ( .A(n3795), .B(p_input[6586]), .Z(o[6586]) );
  AND U7590 ( .A(p_input[26586]), .B(p_input[16586]), .Z(n3795) );
  AND U7591 ( .A(n3796), .B(p_input[6585]), .Z(o[6585]) );
  AND U7592 ( .A(p_input[26585]), .B(p_input[16585]), .Z(n3796) );
  AND U7593 ( .A(n3797), .B(p_input[6584]), .Z(o[6584]) );
  AND U7594 ( .A(p_input[26584]), .B(p_input[16584]), .Z(n3797) );
  AND U7595 ( .A(n3798), .B(p_input[6583]), .Z(o[6583]) );
  AND U7596 ( .A(p_input[26583]), .B(p_input[16583]), .Z(n3798) );
  AND U7597 ( .A(n3799), .B(p_input[6582]), .Z(o[6582]) );
  AND U7598 ( .A(p_input[26582]), .B(p_input[16582]), .Z(n3799) );
  AND U7599 ( .A(n3800), .B(p_input[6581]), .Z(o[6581]) );
  AND U7600 ( .A(p_input[26581]), .B(p_input[16581]), .Z(n3800) );
  AND U7601 ( .A(n3801), .B(p_input[6580]), .Z(o[6580]) );
  AND U7602 ( .A(p_input[26580]), .B(p_input[16580]), .Z(n3801) );
  AND U7603 ( .A(n3802), .B(p_input[657]), .Z(o[657]) );
  AND U7604 ( .A(p_input[20657]), .B(p_input[10657]), .Z(n3802) );
  AND U7605 ( .A(n3803), .B(p_input[6579]), .Z(o[6579]) );
  AND U7606 ( .A(p_input[26579]), .B(p_input[16579]), .Z(n3803) );
  AND U7607 ( .A(n3804), .B(p_input[6578]), .Z(o[6578]) );
  AND U7608 ( .A(p_input[26578]), .B(p_input[16578]), .Z(n3804) );
  AND U7609 ( .A(n3805), .B(p_input[6577]), .Z(o[6577]) );
  AND U7610 ( .A(p_input[26577]), .B(p_input[16577]), .Z(n3805) );
  AND U7611 ( .A(n3806), .B(p_input[6576]), .Z(o[6576]) );
  AND U7612 ( .A(p_input[26576]), .B(p_input[16576]), .Z(n3806) );
  AND U7613 ( .A(n3807), .B(p_input[6575]), .Z(o[6575]) );
  AND U7614 ( .A(p_input[26575]), .B(p_input[16575]), .Z(n3807) );
  AND U7615 ( .A(n3808), .B(p_input[6574]), .Z(o[6574]) );
  AND U7616 ( .A(p_input[26574]), .B(p_input[16574]), .Z(n3808) );
  AND U7617 ( .A(n3809), .B(p_input[6573]), .Z(o[6573]) );
  AND U7618 ( .A(p_input[26573]), .B(p_input[16573]), .Z(n3809) );
  AND U7619 ( .A(n3810), .B(p_input[6572]), .Z(o[6572]) );
  AND U7620 ( .A(p_input[26572]), .B(p_input[16572]), .Z(n3810) );
  AND U7621 ( .A(n3811), .B(p_input[6571]), .Z(o[6571]) );
  AND U7622 ( .A(p_input[26571]), .B(p_input[16571]), .Z(n3811) );
  AND U7623 ( .A(n3812), .B(p_input[6570]), .Z(o[6570]) );
  AND U7624 ( .A(p_input[26570]), .B(p_input[16570]), .Z(n3812) );
  AND U7625 ( .A(n3813), .B(p_input[656]), .Z(o[656]) );
  AND U7626 ( .A(p_input[20656]), .B(p_input[10656]), .Z(n3813) );
  AND U7627 ( .A(n3814), .B(p_input[6569]), .Z(o[6569]) );
  AND U7628 ( .A(p_input[26569]), .B(p_input[16569]), .Z(n3814) );
  AND U7629 ( .A(n3815), .B(p_input[6568]), .Z(o[6568]) );
  AND U7630 ( .A(p_input[26568]), .B(p_input[16568]), .Z(n3815) );
  AND U7631 ( .A(n3816), .B(p_input[6567]), .Z(o[6567]) );
  AND U7632 ( .A(p_input[26567]), .B(p_input[16567]), .Z(n3816) );
  AND U7633 ( .A(n3817), .B(p_input[6566]), .Z(o[6566]) );
  AND U7634 ( .A(p_input[26566]), .B(p_input[16566]), .Z(n3817) );
  AND U7635 ( .A(n3818), .B(p_input[6565]), .Z(o[6565]) );
  AND U7636 ( .A(p_input[26565]), .B(p_input[16565]), .Z(n3818) );
  AND U7637 ( .A(n3819), .B(p_input[6564]), .Z(o[6564]) );
  AND U7638 ( .A(p_input[26564]), .B(p_input[16564]), .Z(n3819) );
  AND U7639 ( .A(n3820), .B(p_input[6563]), .Z(o[6563]) );
  AND U7640 ( .A(p_input[26563]), .B(p_input[16563]), .Z(n3820) );
  AND U7641 ( .A(n3821), .B(p_input[6562]), .Z(o[6562]) );
  AND U7642 ( .A(p_input[26562]), .B(p_input[16562]), .Z(n3821) );
  AND U7643 ( .A(n3822), .B(p_input[6561]), .Z(o[6561]) );
  AND U7644 ( .A(p_input[26561]), .B(p_input[16561]), .Z(n3822) );
  AND U7645 ( .A(n3823), .B(p_input[6560]), .Z(o[6560]) );
  AND U7646 ( .A(p_input[26560]), .B(p_input[16560]), .Z(n3823) );
  AND U7647 ( .A(n3824), .B(p_input[655]), .Z(o[655]) );
  AND U7648 ( .A(p_input[20655]), .B(p_input[10655]), .Z(n3824) );
  AND U7649 ( .A(n3825), .B(p_input[6559]), .Z(o[6559]) );
  AND U7650 ( .A(p_input[26559]), .B(p_input[16559]), .Z(n3825) );
  AND U7651 ( .A(n3826), .B(p_input[6558]), .Z(o[6558]) );
  AND U7652 ( .A(p_input[26558]), .B(p_input[16558]), .Z(n3826) );
  AND U7653 ( .A(n3827), .B(p_input[6557]), .Z(o[6557]) );
  AND U7654 ( .A(p_input[26557]), .B(p_input[16557]), .Z(n3827) );
  AND U7655 ( .A(n3828), .B(p_input[6556]), .Z(o[6556]) );
  AND U7656 ( .A(p_input[26556]), .B(p_input[16556]), .Z(n3828) );
  AND U7657 ( .A(n3829), .B(p_input[6555]), .Z(o[6555]) );
  AND U7658 ( .A(p_input[26555]), .B(p_input[16555]), .Z(n3829) );
  AND U7659 ( .A(n3830), .B(p_input[6554]), .Z(o[6554]) );
  AND U7660 ( .A(p_input[26554]), .B(p_input[16554]), .Z(n3830) );
  AND U7661 ( .A(n3831), .B(p_input[6553]), .Z(o[6553]) );
  AND U7662 ( .A(p_input[26553]), .B(p_input[16553]), .Z(n3831) );
  AND U7663 ( .A(n3832), .B(p_input[6552]), .Z(o[6552]) );
  AND U7664 ( .A(p_input[26552]), .B(p_input[16552]), .Z(n3832) );
  AND U7665 ( .A(n3833), .B(p_input[6551]), .Z(o[6551]) );
  AND U7666 ( .A(p_input[26551]), .B(p_input[16551]), .Z(n3833) );
  AND U7667 ( .A(n3834), .B(p_input[6550]), .Z(o[6550]) );
  AND U7668 ( .A(p_input[26550]), .B(p_input[16550]), .Z(n3834) );
  AND U7669 ( .A(n3835), .B(p_input[654]), .Z(o[654]) );
  AND U7670 ( .A(p_input[20654]), .B(p_input[10654]), .Z(n3835) );
  AND U7671 ( .A(n3836), .B(p_input[6549]), .Z(o[6549]) );
  AND U7672 ( .A(p_input[26549]), .B(p_input[16549]), .Z(n3836) );
  AND U7673 ( .A(n3837), .B(p_input[6548]), .Z(o[6548]) );
  AND U7674 ( .A(p_input[26548]), .B(p_input[16548]), .Z(n3837) );
  AND U7675 ( .A(n3838), .B(p_input[6547]), .Z(o[6547]) );
  AND U7676 ( .A(p_input[26547]), .B(p_input[16547]), .Z(n3838) );
  AND U7677 ( .A(n3839), .B(p_input[6546]), .Z(o[6546]) );
  AND U7678 ( .A(p_input[26546]), .B(p_input[16546]), .Z(n3839) );
  AND U7679 ( .A(n3840), .B(p_input[6545]), .Z(o[6545]) );
  AND U7680 ( .A(p_input[26545]), .B(p_input[16545]), .Z(n3840) );
  AND U7681 ( .A(n3841), .B(p_input[6544]), .Z(o[6544]) );
  AND U7682 ( .A(p_input[26544]), .B(p_input[16544]), .Z(n3841) );
  AND U7683 ( .A(n3842), .B(p_input[6543]), .Z(o[6543]) );
  AND U7684 ( .A(p_input[26543]), .B(p_input[16543]), .Z(n3842) );
  AND U7685 ( .A(n3843), .B(p_input[6542]), .Z(o[6542]) );
  AND U7686 ( .A(p_input[26542]), .B(p_input[16542]), .Z(n3843) );
  AND U7687 ( .A(n3844), .B(p_input[6541]), .Z(o[6541]) );
  AND U7688 ( .A(p_input[26541]), .B(p_input[16541]), .Z(n3844) );
  AND U7689 ( .A(n3845), .B(p_input[6540]), .Z(o[6540]) );
  AND U7690 ( .A(p_input[26540]), .B(p_input[16540]), .Z(n3845) );
  AND U7691 ( .A(n3846), .B(p_input[653]), .Z(o[653]) );
  AND U7692 ( .A(p_input[20653]), .B(p_input[10653]), .Z(n3846) );
  AND U7693 ( .A(n3847), .B(p_input[6539]), .Z(o[6539]) );
  AND U7694 ( .A(p_input[26539]), .B(p_input[16539]), .Z(n3847) );
  AND U7695 ( .A(n3848), .B(p_input[6538]), .Z(o[6538]) );
  AND U7696 ( .A(p_input[26538]), .B(p_input[16538]), .Z(n3848) );
  AND U7697 ( .A(n3849), .B(p_input[6537]), .Z(o[6537]) );
  AND U7698 ( .A(p_input[26537]), .B(p_input[16537]), .Z(n3849) );
  AND U7699 ( .A(n3850), .B(p_input[6536]), .Z(o[6536]) );
  AND U7700 ( .A(p_input[26536]), .B(p_input[16536]), .Z(n3850) );
  AND U7701 ( .A(n3851), .B(p_input[6535]), .Z(o[6535]) );
  AND U7702 ( .A(p_input[26535]), .B(p_input[16535]), .Z(n3851) );
  AND U7703 ( .A(n3852), .B(p_input[6534]), .Z(o[6534]) );
  AND U7704 ( .A(p_input[26534]), .B(p_input[16534]), .Z(n3852) );
  AND U7705 ( .A(n3853), .B(p_input[6533]), .Z(o[6533]) );
  AND U7706 ( .A(p_input[26533]), .B(p_input[16533]), .Z(n3853) );
  AND U7707 ( .A(n3854), .B(p_input[6532]), .Z(o[6532]) );
  AND U7708 ( .A(p_input[26532]), .B(p_input[16532]), .Z(n3854) );
  AND U7709 ( .A(n3855), .B(p_input[6531]), .Z(o[6531]) );
  AND U7710 ( .A(p_input[26531]), .B(p_input[16531]), .Z(n3855) );
  AND U7711 ( .A(n3856), .B(p_input[6530]), .Z(o[6530]) );
  AND U7712 ( .A(p_input[26530]), .B(p_input[16530]), .Z(n3856) );
  AND U7713 ( .A(n3857), .B(p_input[652]), .Z(o[652]) );
  AND U7714 ( .A(p_input[20652]), .B(p_input[10652]), .Z(n3857) );
  AND U7715 ( .A(n3858), .B(p_input[6529]), .Z(o[6529]) );
  AND U7716 ( .A(p_input[26529]), .B(p_input[16529]), .Z(n3858) );
  AND U7717 ( .A(n3859), .B(p_input[6528]), .Z(o[6528]) );
  AND U7718 ( .A(p_input[26528]), .B(p_input[16528]), .Z(n3859) );
  AND U7719 ( .A(n3860), .B(p_input[6527]), .Z(o[6527]) );
  AND U7720 ( .A(p_input[26527]), .B(p_input[16527]), .Z(n3860) );
  AND U7721 ( .A(n3861), .B(p_input[6526]), .Z(o[6526]) );
  AND U7722 ( .A(p_input[26526]), .B(p_input[16526]), .Z(n3861) );
  AND U7723 ( .A(n3862), .B(p_input[6525]), .Z(o[6525]) );
  AND U7724 ( .A(p_input[26525]), .B(p_input[16525]), .Z(n3862) );
  AND U7725 ( .A(n3863), .B(p_input[6524]), .Z(o[6524]) );
  AND U7726 ( .A(p_input[26524]), .B(p_input[16524]), .Z(n3863) );
  AND U7727 ( .A(n3864), .B(p_input[6523]), .Z(o[6523]) );
  AND U7728 ( .A(p_input[26523]), .B(p_input[16523]), .Z(n3864) );
  AND U7729 ( .A(n3865), .B(p_input[6522]), .Z(o[6522]) );
  AND U7730 ( .A(p_input[26522]), .B(p_input[16522]), .Z(n3865) );
  AND U7731 ( .A(n3866), .B(p_input[6521]), .Z(o[6521]) );
  AND U7732 ( .A(p_input[26521]), .B(p_input[16521]), .Z(n3866) );
  AND U7733 ( .A(n3867), .B(p_input[6520]), .Z(o[6520]) );
  AND U7734 ( .A(p_input[26520]), .B(p_input[16520]), .Z(n3867) );
  AND U7735 ( .A(n3868), .B(p_input[651]), .Z(o[651]) );
  AND U7736 ( .A(p_input[20651]), .B(p_input[10651]), .Z(n3868) );
  AND U7737 ( .A(n3869), .B(p_input[6519]), .Z(o[6519]) );
  AND U7738 ( .A(p_input[26519]), .B(p_input[16519]), .Z(n3869) );
  AND U7739 ( .A(n3870), .B(p_input[6518]), .Z(o[6518]) );
  AND U7740 ( .A(p_input[26518]), .B(p_input[16518]), .Z(n3870) );
  AND U7741 ( .A(n3871), .B(p_input[6517]), .Z(o[6517]) );
  AND U7742 ( .A(p_input[26517]), .B(p_input[16517]), .Z(n3871) );
  AND U7743 ( .A(n3872), .B(p_input[6516]), .Z(o[6516]) );
  AND U7744 ( .A(p_input[26516]), .B(p_input[16516]), .Z(n3872) );
  AND U7745 ( .A(n3873), .B(p_input[6515]), .Z(o[6515]) );
  AND U7746 ( .A(p_input[26515]), .B(p_input[16515]), .Z(n3873) );
  AND U7747 ( .A(n3874), .B(p_input[6514]), .Z(o[6514]) );
  AND U7748 ( .A(p_input[26514]), .B(p_input[16514]), .Z(n3874) );
  AND U7749 ( .A(n3875), .B(p_input[6513]), .Z(o[6513]) );
  AND U7750 ( .A(p_input[26513]), .B(p_input[16513]), .Z(n3875) );
  AND U7751 ( .A(n3876), .B(p_input[6512]), .Z(o[6512]) );
  AND U7752 ( .A(p_input[26512]), .B(p_input[16512]), .Z(n3876) );
  AND U7753 ( .A(n3877), .B(p_input[6511]), .Z(o[6511]) );
  AND U7754 ( .A(p_input[26511]), .B(p_input[16511]), .Z(n3877) );
  AND U7755 ( .A(n3878), .B(p_input[6510]), .Z(o[6510]) );
  AND U7756 ( .A(p_input[26510]), .B(p_input[16510]), .Z(n3878) );
  AND U7757 ( .A(n3879), .B(p_input[650]), .Z(o[650]) );
  AND U7758 ( .A(p_input[20650]), .B(p_input[10650]), .Z(n3879) );
  AND U7759 ( .A(n3880), .B(p_input[6509]), .Z(o[6509]) );
  AND U7760 ( .A(p_input[26509]), .B(p_input[16509]), .Z(n3880) );
  AND U7761 ( .A(n3881), .B(p_input[6508]), .Z(o[6508]) );
  AND U7762 ( .A(p_input[26508]), .B(p_input[16508]), .Z(n3881) );
  AND U7763 ( .A(n3882), .B(p_input[6507]), .Z(o[6507]) );
  AND U7764 ( .A(p_input[26507]), .B(p_input[16507]), .Z(n3882) );
  AND U7765 ( .A(n3883), .B(p_input[6506]), .Z(o[6506]) );
  AND U7766 ( .A(p_input[26506]), .B(p_input[16506]), .Z(n3883) );
  AND U7767 ( .A(n3884), .B(p_input[6505]), .Z(o[6505]) );
  AND U7768 ( .A(p_input[26505]), .B(p_input[16505]), .Z(n3884) );
  AND U7769 ( .A(n3885), .B(p_input[6504]), .Z(o[6504]) );
  AND U7770 ( .A(p_input[26504]), .B(p_input[16504]), .Z(n3885) );
  AND U7771 ( .A(n3886), .B(p_input[6503]), .Z(o[6503]) );
  AND U7772 ( .A(p_input[26503]), .B(p_input[16503]), .Z(n3886) );
  AND U7773 ( .A(n3887), .B(p_input[6502]), .Z(o[6502]) );
  AND U7774 ( .A(p_input[26502]), .B(p_input[16502]), .Z(n3887) );
  AND U7775 ( .A(n3888), .B(p_input[6501]), .Z(o[6501]) );
  AND U7776 ( .A(p_input[26501]), .B(p_input[16501]), .Z(n3888) );
  AND U7777 ( .A(n3889), .B(p_input[6500]), .Z(o[6500]) );
  AND U7778 ( .A(p_input[26500]), .B(p_input[16500]), .Z(n3889) );
  AND U7779 ( .A(n3890), .B(p_input[64]), .Z(o[64]) );
  AND U7780 ( .A(p_input[20064]), .B(p_input[10064]), .Z(n3890) );
  AND U7781 ( .A(n3891), .B(p_input[649]), .Z(o[649]) );
  AND U7782 ( .A(p_input[20649]), .B(p_input[10649]), .Z(n3891) );
  AND U7783 ( .A(n3892), .B(p_input[6499]), .Z(o[6499]) );
  AND U7784 ( .A(p_input[26499]), .B(p_input[16499]), .Z(n3892) );
  AND U7785 ( .A(n3893), .B(p_input[6498]), .Z(o[6498]) );
  AND U7786 ( .A(p_input[26498]), .B(p_input[16498]), .Z(n3893) );
  AND U7787 ( .A(n3894), .B(p_input[6497]), .Z(o[6497]) );
  AND U7788 ( .A(p_input[26497]), .B(p_input[16497]), .Z(n3894) );
  AND U7789 ( .A(n3895), .B(p_input[6496]), .Z(o[6496]) );
  AND U7790 ( .A(p_input[26496]), .B(p_input[16496]), .Z(n3895) );
  AND U7791 ( .A(n3896), .B(p_input[6495]), .Z(o[6495]) );
  AND U7792 ( .A(p_input[26495]), .B(p_input[16495]), .Z(n3896) );
  AND U7793 ( .A(n3897), .B(p_input[6494]), .Z(o[6494]) );
  AND U7794 ( .A(p_input[26494]), .B(p_input[16494]), .Z(n3897) );
  AND U7795 ( .A(n3898), .B(p_input[6493]), .Z(o[6493]) );
  AND U7796 ( .A(p_input[26493]), .B(p_input[16493]), .Z(n3898) );
  AND U7797 ( .A(n3899), .B(p_input[6492]), .Z(o[6492]) );
  AND U7798 ( .A(p_input[26492]), .B(p_input[16492]), .Z(n3899) );
  AND U7799 ( .A(n3900), .B(p_input[6491]), .Z(o[6491]) );
  AND U7800 ( .A(p_input[26491]), .B(p_input[16491]), .Z(n3900) );
  AND U7801 ( .A(n3901), .B(p_input[6490]), .Z(o[6490]) );
  AND U7802 ( .A(p_input[26490]), .B(p_input[16490]), .Z(n3901) );
  AND U7803 ( .A(n3902), .B(p_input[648]), .Z(o[648]) );
  AND U7804 ( .A(p_input[20648]), .B(p_input[10648]), .Z(n3902) );
  AND U7805 ( .A(n3903), .B(p_input[6489]), .Z(o[6489]) );
  AND U7806 ( .A(p_input[26489]), .B(p_input[16489]), .Z(n3903) );
  AND U7807 ( .A(n3904), .B(p_input[6488]), .Z(o[6488]) );
  AND U7808 ( .A(p_input[26488]), .B(p_input[16488]), .Z(n3904) );
  AND U7809 ( .A(n3905), .B(p_input[6487]), .Z(o[6487]) );
  AND U7810 ( .A(p_input[26487]), .B(p_input[16487]), .Z(n3905) );
  AND U7811 ( .A(n3906), .B(p_input[6486]), .Z(o[6486]) );
  AND U7812 ( .A(p_input[26486]), .B(p_input[16486]), .Z(n3906) );
  AND U7813 ( .A(n3907), .B(p_input[6485]), .Z(o[6485]) );
  AND U7814 ( .A(p_input[26485]), .B(p_input[16485]), .Z(n3907) );
  AND U7815 ( .A(n3908), .B(p_input[6484]), .Z(o[6484]) );
  AND U7816 ( .A(p_input[26484]), .B(p_input[16484]), .Z(n3908) );
  AND U7817 ( .A(n3909), .B(p_input[6483]), .Z(o[6483]) );
  AND U7818 ( .A(p_input[26483]), .B(p_input[16483]), .Z(n3909) );
  AND U7819 ( .A(n3910), .B(p_input[6482]), .Z(o[6482]) );
  AND U7820 ( .A(p_input[26482]), .B(p_input[16482]), .Z(n3910) );
  AND U7821 ( .A(n3911), .B(p_input[6481]), .Z(o[6481]) );
  AND U7822 ( .A(p_input[26481]), .B(p_input[16481]), .Z(n3911) );
  AND U7823 ( .A(n3912), .B(p_input[6480]), .Z(o[6480]) );
  AND U7824 ( .A(p_input[26480]), .B(p_input[16480]), .Z(n3912) );
  AND U7825 ( .A(n3913), .B(p_input[647]), .Z(o[647]) );
  AND U7826 ( .A(p_input[20647]), .B(p_input[10647]), .Z(n3913) );
  AND U7827 ( .A(n3914), .B(p_input[6479]), .Z(o[6479]) );
  AND U7828 ( .A(p_input[26479]), .B(p_input[16479]), .Z(n3914) );
  AND U7829 ( .A(n3915), .B(p_input[6478]), .Z(o[6478]) );
  AND U7830 ( .A(p_input[26478]), .B(p_input[16478]), .Z(n3915) );
  AND U7831 ( .A(n3916), .B(p_input[6477]), .Z(o[6477]) );
  AND U7832 ( .A(p_input[26477]), .B(p_input[16477]), .Z(n3916) );
  AND U7833 ( .A(n3917), .B(p_input[6476]), .Z(o[6476]) );
  AND U7834 ( .A(p_input[26476]), .B(p_input[16476]), .Z(n3917) );
  AND U7835 ( .A(n3918), .B(p_input[6475]), .Z(o[6475]) );
  AND U7836 ( .A(p_input[26475]), .B(p_input[16475]), .Z(n3918) );
  AND U7837 ( .A(n3919), .B(p_input[6474]), .Z(o[6474]) );
  AND U7838 ( .A(p_input[26474]), .B(p_input[16474]), .Z(n3919) );
  AND U7839 ( .A(n3920), .B(p_input[6473]), .Z(o[6473]) );
  AND U7840 ( .A(p_input[26473]), .B(p_input[16473]), .Z(n3920) );
  AND U7841 ( .A(n3921), .B(p_input[6472]), .Z(o[6472]) );
  AND U7842 ( .A(p_input[26472]), .B(p_input[16472]), .Z(n3921) );
  AND U7843 ( .A(n3922), .B(p_input[6471]), .Z(o[6471]) );
  AND U7844 ( .A(p_input[26471]), .B(p_input[16471]), .Z(n3922) );
  AND U7845 ( .A(n3923), .B(p_input[6470]), .Z(o[6470]) );
  AND U7846 ( .A(p_input[26470]), .B(p_input[16470]), .Z(n3923) );
  AND U7847 ( .A(n3924), .B(p_input[646]), .Z(o[646]) );
  AND U7848 ( .A(p_input[20646]), .B(p_input[10646]), .Z(n3924) );
  AND U7849 ( .A(n3925), .B(p_input[6469]), .Z(o[6469]) );
  AND U7850 ( .A(p_input[26469]), .B(p_input[16469]), .Z(n3925) );
  AND U7851 ( .A(n3926), .B(p_input[6468]), .Z(o[6468]) );
  AND U7852 ( .A(p_input[26468]), .B(p_input[16468]), .Z(n3926) );
  AND U7853 ( .A(n3927), .B(p_input[6467]), .Z(o[6467]) );
  AND U7854 ( .A(p_input[26467]), .B(p_input[16467]), .Z(n3927) );
  AND U7855 ( .A(n3928), .B(p_input[6466]), .Z(o[6466]) );
  AND U7856 ( .A(p_input[26466]), .B(p_input[16466]), .Z(n3928) );
  AND U7857 ( .A(n3929), .B(p_input[6465]), .Z(o[6465]) );
  AND U7858 ( .A(p_input[26465]), .B(p_input[16465]), .Z(n3929) );
  AND U7859 ( .A(n3930), .B(p_input[6464]), .Z(o[6464]) );
  AND U7860 ( .A(p_input[26464]), .B(p_input[16464]), .Z(n3930) );
  AND U7861 ( .A(n3931), .B(p_input[6463]), .Z(o[6463]) );
  AND U7862 ( .A(p_input[26463]), .B(p_input[16463]), .Z(n3931) );
  AND U7863 ( .A(n3932), .B(p_input[6462]), .Z(o[6462]) );
  AND U7864 ( .A(p_input[26462]), .B(p_input[16462]), .Z(n3932) );
  AND U7865 ( .A(n3933), .B(p_input[6461]), .Z(o[6461]) );
  AND U7866 ( .A(p_input[26461]), .B(p_input[16461]), .Z(n3933) );
  AND U7867 ( .A(n3934), .B(p_input[6460]), .Z(o[6460]) );
  AND U7868 ( .A(p_input[26460]), .B(p_input[16460]), .Z(n3934) );
  AND U7869 ( .A(n3935), .B(p_input[645]), .Z(o[645]) );
  AND U7870 ( .A(p_input[20645]), .B(p_input[10645]), .Z(n3935) );
  AND U7871 ( .A(n3936), .B(p_input[6459]), .Z(o[6459]) );
  AND U7872 ( .A(p_input[26459]), .B(p_input[16459]), .Z(n3936) );
  AND U7873 ( .A(n3937), .B(p_input[6458]), .Z(o[6458]) );
  AND U7874 ( .A(p_input[26458]), .B(p_input[16458]), .Z(n3937) );
  AND U7875 ( .A(n3938), .B(p_input[6457]), .Z(o[6457]) );
  AND U7876 ( .A(p_input[26457]), .B(p_input[16457]), .Z(n3938) );
  AND U7877 ( .A(n3939), .B(p_input[6456]), .Z(o[6456]) );
  AND U7878 ( .A(p_input[26456]), .B(p_input[16456]), .Z(n3939) );
  AND U7879 ( .A(n3940), .B(p_input[6455]), .Z(o[6455]) );
  AND U7880 ( .A(p_input[26455]), .B(p_input[16455]), .Z(n3940) );
  AND U7881 ( .A(n3941), .B(p_input[6454]), .Z(o[6454]) );
  AND U7882 ( .A(p_input[26454]), .B(p_input[16454]), .Z(n3941) );
  AND U7883 ( .A(n3942), .B(p_input[6453]), .Z(o[6453]) );
  AND U7884 ( .A(p_input[26453]), .B(p_input[16453]), .Z(n3942) );
  AND U7885 ( .A(n3943), .B(p_input[6452]), .Z(o[6452]) );
  AND U7886 ( .A(p_input[26452]), .B(p_input[16452]), .Z(n3943) );
  AND U7887 ( .A(n3944), .B(p_input[6451]), .Z(o[6451]) );
  AND U7888 ( .A(p_input[26451]), .B(p_input[16451]), .Z(n3944) );
  AND U7889 ( .A(n3945), .B(p_input[6450]), .Z(o[6450]) );
  AND U7890 ( .A(p_input[26450]), .B(p_input[16450]), .Z(n3945) );
  AND U7891 ( .A(n3946), .B(p_input[644]), .Z(o[644]) );
  AND U7892 ( .A(p_input[20644]), .B(p_input[10644]), .Z(n3946) );
  AND U7893 ( .A(n3947), .B(p_input[6449]), .Z(o[6449]) );
  AND U7894 ( .A(p_input[26449]), .B(p_input[16449]), .Z(n3947) );
  AND U7895 ( .A(n3948), .B(p_input[6448]), .Z(o[6448]) );
  AND U7896 ( .A(p_input[26448]), .B(p_input[16448]), .Z(n3948) );
  AND U7897 ( .A(n3949), .B(p_input[6447]), .Z(o[6447]) );
  AND U7898 ( .A(p_input[26447]), .B(p_input[16447]), .Z(n3949) );
  AND U7899 ( .A(n3950), .B(p_input[6446]), .Z(o[6446]) );
  AND U7900 ( .A(p_input[26446]), .B(p_input[16446]), .Z(n3950) );
  AND U7901 ( .A(n3951), .B(p_input[6445]), .Z(o[6445]) );
  AND U7902 ( .A(p_input[26445]), .B(p_input[16445]), .Z(n3951) );
  AND U7903 ( .A(n3952), .B(p_input[6444]), .Z(o[6444]) );
  AND U7904 ( .A(p_input[26444]), .B(p_input[16444]), .Z(n3952) );
  AND U7905 ( .A(n3953), .B(p_input[6443]), .Z(o[6443]) );
  AND U7906 ( .A(p_input[26443]), .B(p_input[16443]), .Z(n3953) );
  AND U7907 ( .A(n3954), .B(p_input[6442]), .Z(o[6442]) );
  AND U7908 ( .A(p_input[26442]), .B(p_input[16442]), .Z(n3954) );
  AND U7909 ( .A(n3955), .B(p_input[6441]), .Z(o[6441]) );
  AND U7910 ( .A(p_input[26441]), .B(p_input[16441]), .Z(n3955) );
  AND U7911 ( .A(n3956), .B(p_input[6440]), .Z(o[6440]) );
  AND U7912 ( .A(p_input[26440]), .B(p_input[16440]), .Z(n3956) );
  AND U7913 ( .A(n3957), .B(p_input[643]), .Z(o[643]) );
  AND U7914 ( .A(p_input[20643]), .B(p_input[10643]), .Z(n3957) );
  AND U7915 ( .A(n3958), .B(p_input[6439]), .Z(o[6439]) );
  AND U7916 ( .A(p_input[26439]), .B(p_input[16439]), .Z(n3958) );
  AND U7917 ( .A(n3959), .B(p_input[6438]), .Z(o[6438]) );
  AND U7918 ( .A(p_input[26438]), .B(p_input[16438]), .Z(n3959) );
  AND U7919 ( .A(n3960), .B(p_input[6437]), .Z(o[6437]) );
  AND U7920 ( .A(p_input[26437]), .B(p_input[16437]), .Z(n3960) );
  AND U7921 ( .A(n3961), .B(p_input[6436]), .Z(o[6436]) );
  AND U7922 ( .A(p_input[26436]), .B(p_input[16436]), .Z(n3961) );
  AND U7923 ( .A(n3962), .B(p_input[6435]), .Z(o[6435]) );
  AND U7924 ( .A(p_input[26435]), .B(p_input[16435]), .Z(n3962) );
  AND U7925 ( .A(n3963), .B(p_input[6434]), .Z(o[6434]) );
  AND U7926 ( .A(p_input[26434]), .B(p_input[16434]), .Z(n3963) );
  AND U7927 ( .A(n3964), .B(p_input[6433]), .Z(o[6433]) );
  AND U7928 ( .A(p_input[26433]), .B(p_input[16433]), .Z(n3964) );
  AND U7929 ( .A(n3965), .B(p_input[6432]), .Z(o[6432]) );
  AND U7930 ( .A(p_input[26432]), .B(p_input[16432]), .Z(n3965) );
  AND U7931 ( .A(n3966), .B(p_input[6431]), .Z(o[6431]) );
  AND U7932 ( .A(p_input[26431]), .B(p_input[16431]), .Z(n3966) );
  AND U7933 ( .A(n3967), .B(p_input[6430]), .Z(o[6430]) );
  AND U7934 ( .A(p_input[26430]), .B(p_input[16430]), .Z(n3967) );
  AND U7935 ( .A(n3968), .B(p_input[642]), .Z(o[642]) );
  AND U7936 ( .A(p_input[20642]), .B(p_input[10642]), .Z(n3968) );
  AND U7937 ( .A(n3969), .B(p_input[6429]), .Z(o[6429]) );
  AND U7938 ( .A(p_input[26429]), .B(p_input[16429]), .Z(n3969) );
  AND U7939 ( .A(n3970), .B(p_input[6428]), .Z(o[6428]) );
  AND U7940 ( .A(p_input[26428]), .B(p_input[16428]), .Z(n3970) );
  AND U7941 ( .A(n3971), .B(p_input[6427]), .Z(o[6427]) );
  AND U7942 ( .A(p_input[26427]), .B(p_input[16427]), .Z(n3971) );
  AND U7943 ( .A(n3972), .B(p_input[6426]), .Z(o[6426]) );
  AND U7944 ( .A(p_input[26426]), .B(p_input[16426]), .Z(n3972) );
  AND U7945 ( .A(n3973), .B(p_input[6425]), .Z(o[6425]) );
  AND U7946 ( .A(p_input[26425]), .B(p_input[16425]), .Z(n3973) );
  AND U7947 ( .A(n3974), .B(p_input[6424]), .Z(o[6424]) );
  AND U7948 ( .A(p_input[26424]), .B(p_input[16424]), .Z(n3974) );
  AND U7949 ( .A(n3975), .B(p_input[6423]), .Z(o[6423]) );
  AND U7950 ( .A(p_input[26423]), .B(p_input[16423]), .Z(n3975) );
  AND U7951 ( .A(n3976), .B(p_input[6422]), .Z(o[6422]) );
  AND U7952 ( .A(p_input[26422]), .B(p_input[16422]), .Z(n3976) );
  AND U7953 ( .A(n3977), .B(p_input[6421]), .Z(o[6421]) );
  AND U7954 ( .A(p_input[26421]), .B(p_input[16421]), .Z(n3977) );
  AND U7955 ( .A(n3978), .B(p_input[6420]), .Z(o[6420]) );
  AND U7956 ( .A(p_input[26420]), .B(p_input[16420]), .Z(n3978) );
  AND U7957 ( .A(n3979), .B(p_input[641]), .Z(o[641]) );
  AND U7958 ( .A(p_input[20641]), .B(p_input[10641]), .Z(n3979) );
  AND U7959 ( .A(n3980), .B(p_input[6419]), .Z(o[6419]) );
  AND U7960 ( .A(p_input[26419]), .B(p_input[16419]), .Z(n3980) );
  AND U7961 ( .A(n3981), .B(p_input[6418]), .Z(o[6418]) );
  AND U7962 ( .A(p_input[26418]), .B(p_input[16418]), .Z(n3981) );
  AND U7963 ( .A(n3982), .B(p_input[6417]), .Z(o[6417]) );
  AND U7964 ( .A(p_input[26417]), .B(p_input[16417]), .Z(n3982) );
  AND U7965 ( .A(n3983), .B(p_input[6416]), .Z(o[6416]) );
  AND U7966 ( .A(p_input[26416]), .B(p_input[16416]), .Z(n3983) );
  AND U7967 ( .A(n3984), .B(p_input[6415]), .Z(o[6415]) );
  AND U7968 ( .A(p_input[26415]), .B(p_input[16415]), .Z(n3984) );
  AND U7969 ( .A(n3985), .B(p_input[6414]), .Z(o[6414]) );
  AND U7970 ( .A(p_input[26414]), .B(p_input[16414]), .Z(n3985) );
  AND U7971 ( .A(n3986), .B(p_input[6413]), .Z(o[6413]) );
  AND U7972 ( .A(p_input[26413]), .B(p_input[16413]), .Z(n3986) );
  AND U7973 ( .A(n3987), .B(p_input[6412]), .Z(o[6412]) );
  AND U7974 ( .A(p_input[26412]), .B(p_input[16412]), .Z(n3987) );
  AND U7975 ( .A(n3988), .B(p_input[6411]), .Z(o[6411]) );
  AND U7976 ( .A(p_input[26411]), .B(p_input[16411]), .Z(n3988) );
  AND U7977 ( .A(n3989), .B(p_input[6410]), .Z(o[6410]) );
  AND U7978 ( .A(p_input[26410]), .B(p_input[16410]), .Z(n3989) );
  AND U7979 ( .A(n3990), .B(p_input[640]), .Z(o[640]) );
  AND U7980 ( .A(p_input[20640]), .B(p_input[10640]), .Z(n3990) );
  AND U7981 ( .A(n3991), .B(p_input[6409]), .Z(o[6409]) );
  AND U7982 ( .A(p_input[26409]), .B(p_input[16409]), .Z(n3991) );
  AND U7983 ( .A(n3992), .B(p_input[6408]), .Z(o[6408]) );
  AND U7984 ( .A(p_input[26408]), .B(p_input[16408]), .Z(n3992) );
  AND U7985 ( .A(n3993), .B(p_input[6407]), .Z(o[6407]) );
  AND U7986 ( .A(p_input[26407]), .B(p_input[16407]), .Z(n3993) );
  AND U7987 ( .A(n3994), .B(p_input[6406]), .Z(o[6406]) );
  AND U7988 ( .A(p_input[26406]), .B(p_input[16406]), .Z(n3994) );
  AND U7989 ( .A(n3995), .B(p_input[6405]), .Z(o[6405]) );
  AND U7990 ( .A(p_input[26405]), .B(p_input[16405]), .Z(n3995) );
  AND U7991 ( .A(n3996), .B(p_input[6404]), .Z(o[6404]) );
  AND U7992 ( .A(p_input[26404]), .B(p_input[16404]), .Z(n3996) );
  AND U7993 ( .A(n3997), .B(p_input[6403]), .Z(o[6403]) );
  AND U7994 ( .A(p_input[26403]), .B(p_input[16403]), .Z(n3997) );
  AND U7995 ( .A(n3998), .B(p_input[6402]), .Z(o[6402]) );
  AND U7996 ( .A(p_input[26402]), .B(p_input[16402]), .Z(n3998) );
  AND U7997 ( .A(n3999), .B(p_input[6401]), .Z(o[6401]) );
  AND U7998 ( .A(p_input[26401]), .B(p_input[16401]), .Z(n3999) );
  AND U7999 ( .A(n4000), .B(p_input[6400]), .Z(o[6400]) );
  AND U8000 ( .A(p_input[26400]), .B(p_input[16400]), .Z(n4000) );
  AND U8001 ( .A(n4001), .B(p_input[63]), .Z(o[63]) );
  AND U8002 ( .A(p_input[20063]), .B(p_input[10063]), .Z(n4001) );
  AND U8003 ( .A(n4002), .B(p_input[639]), .Z(o[639]) );
  AND U8004 ( .A(p_input[20639]), .B(p_input[10639]), .Z(n4002) );
  AND U8005 ( .A(n4003), .B(p_input[6399]), .Z(o[6399]) );
  AND U8006 ( .A(p_input[26399]), .B(p_input[16399]), .Z(n4003) );
  AND U8007 ( .A(n4004), .B(p_input[6398]), .Z(o[6398]) );
  AND U8008 ( .A(p_input[26398]), .B(p_input[16398]), .Z(n4004) );
  AND U8009 ( .A(n4005), .B(p_input[6397]), .Z(o[6397]) );
  AND U8010 ( .A(p_input[26397]), .B(p_input[16397]), .Z(n4005) );
  AND U8011 ( .A(n4006), .B(p_input[6396]), .Z(o[6396]) );
  AND U8012 ( .A(p_input[26396]), .B(p_input[16396]), .Z(n4006) );
  AND U8013 ( .A(n4007), .B(p_input[6395]), .Z(o[6395]) );
  AND U8014 ( .A(p_input[26395]), .B(p_input[16395]), .Z(n4007) );
  AND U8015 ( .A(n4008), .B(p_input[6394]), .Z(o[6394]) );
  AND U8016 ( .A(p_input[26394]), .B(p_input[16394]), .Z(n4008) );
  AND U8017 ( .A(n4009), .B(p_input[6393]), .Z(o[6393]) );
  AND U8018 ( .A(p_input[26393]), .B(p_input[16393]), .Z(n4009) );
  AND U8019 ( .A(n4010), .B(p_input[6392]), .Z(o[6392]) );
  AND U8020 ( .A(p_input[26392]), .B(p_input[16392]), .Z(n4010) );
  AND U8021 ( .A(n4011), .B(p_input[6391]), .Z(o[6391]) );
  AND U8022 ( .A(p_input[26391]), .B(p_input[16391]), .Z(n4011) );
  AND U8023 ( .A(n4012), .B(p_input[6390]), .Z(o[6390]) );
  AND U8024 ( .A(p_input[26390]), .B(p_input[16390]), .Z(n4012) );
  AND U8025 ( .A(n4013), .B(p_input[638]), .Z(o[638]) );
  AND U8026 ( .A(p_input[20638]), .B(p_input[10638]), .Z(n4013) );
  AND U8027 ( .A(n4014), .B(p_input[6389]), .Z(o[6389]) );
  AND U8028 ( .A(p_input[26389]), .B(p_input[16389]), .Z(n4014) );
  AND U8029 ( .A(n4015), .B(p_input[6388]), .Z(o[6388]) );
  AND U8030 ( .A(p_input[26388]), .B(p_input[16388]), .Z(n4015) );
  AND U8031 ( .A(n4016), .B(p_input[6387]), .Z(o[6387]) );
  AND U8032 ( .A(p_input[26387]), .B(p_input[16387]), .Z(n4016) );
  AND U8033 ( .A(n4017), .B(p_input[6386]), .Z(o[6386]) );
  AND U8034 ( .A(p_input[26386]), .B(p_input[16386]), .Z(n4017) );
  AND U8035 ( .A(n4018), .B(p_input[6385]), .Z(o[6385]) );
  AND U8036 ( .A(p_input[26385]), .B(p_input[16385]), .Z(n4018) );
  AND U8037 ( .A(n4019), .B(p_input[6384]), .Z(o[6384]) );
  AND U8038 ( .A(p_input[26384]), .B(p_input[16384]), .Z(n4019) );
  AND U8039 ( .A(n4020), .B(p_input[6383]), .Z(o[6383]) );
  AND U8040 ( .A(p_input[26383]), .B(p_input[16383]), .Z(n4020) );
  AND U8041 ( .A(n4021), .B(p_input[6382]), .Z(o[6382]) );
  AND U8042 ( .A(p_input[26382]), .B(p_input[16382]), .Z(n4021) );
  AND U8043 ( .A(n4022), .B(p_input[6381]), .Z(o[6381]) );
  AND U8044 ( .A(p_input[26381]), .B(p_input[16381]), .Z(n4022) );
  AND U8045 ( .A(n4023), .B(p_input[6380]), .Z(o[6380]) );
  AND U8046 ( .A(p_input[26380]), .B(p_input[16380]), .Z(n4023) );
  AND U8047 ( .A(n4024), .B(p_input[637]), .Z(o[637]) );
  AND U8048 ( .A(p_input[20637]), .B(p_input[10637]), .Z(n4024) );
  AND U8049 ( .A(n4025), .B(p_input[6379]), .Z(o[6379]) );
  AND U8050 ( .A(p_input[26379]), .B(p_input[16379]), .Z(n4025) );
  AND U8051 ( .A(n4026), .B(p_input[6378]), .Z(o[6378]) );
  AND U8052 ( .A(p_input[26378]), .B(p_input[16378]), .Z(n4026) );
  AND U8053 ( .A(n4027), .B(p_input[6377]), .Z(o[6377]) );
  AND U8054 ( .A(p_input[26377]), .B(p_input[16377]), .Z(n4027) );
  AND U8055 ( .A(n4028), .B(p_input[6376]), .Z(o[6376]) );
  AND U8056 ( .A(p_input[26376]), .B(p_input[16376]), .Z(n4028) );
  AND U8057 ( .A(n4029), .B(p_input[6375]), .Z(o[6375]) );
  AND U8058 ( .A(p_input[26375]), .B(p_input[16375]), .Z(n4029) );
  AND U8059 ( .A(n4030), .B(p_input[6374]), .Z(o[6374]) );
  AND U8060 ( .A(p_input[26374]), .B(p_input[16374]), .Z(n4030) );
  AND U8061 ( .A(n4031), .B(p_input[6373]), .Z(o[6373]) );
  AND U8062 ( .A(p_input[26373]), .B(p_input[16373]), .Z(n4031) );
  AND U8063 ( .A(n4032), .B(p_input[6372]), .Z(o[6372]) );
  AND U8064 ( .A(p_input[26372]), .B(p_input[16372]), .Z(n4032) );
  AND U8065 ( .A(n4033), .B(p_input[6371]), .Z(o[6371]) );
  AND U8066 ( .A(p_input[26371]), .B(p_input[16371]), .Z(n4033) );
  AND U8067 ( .A(n4034), .B(p_input[6370]), .Z(o[6370]) );
  AND U8068 ( .A(p_input[26370]), .B(p_input[16370]), .Z(n4034) );
  AND U8069 ( .A(n4035), .B(p_input[636]), .Z(o[636]) );
  AND U8070 ( .A(p_input[20636]), .B(p_input[10636]), .Z(n4035) );
  AND U8071 ( .A(n4036), .B(p_input[6369]), .Z(o[6369]) );
  AND U8072 ( .A(p_input[26369]), .B(p_input[16369]), .Z(n4036) );
  AND U8073 ( .A(n4037), .B(p_input[6368]), .Z(o[6368]) );
  AND U8074 ( .A(p_input[26368]), .B(p_input[16368]), .Z(n4037) );
  AND U8075 ( .A(n4038), .B(p_input[6367]), .Z(o[6367]) );
  AND U8076 ( .A(p_input[26367]), .B(p_input[16367]), .Z(n4038) );
  AND U8077 ( .A(n4039), .B(p_input[6366]), .Z(o[6366]) );
  AND U8078 ( .A(p_input[26366]), .B(p_input[16366]), .Z(n4039) );
  AND U8079 ( .A(n4040), .B(p_input[6365]), .Z(o[6365]) );
  AND U8080 ( .A(p_input[26365]), .B(p_input[16365]), .Z(n4040) );
  AND U8081 ( .A(n4041), .B(p_input[6364]), .Z(o[6364]) );
  AND U8082 ( .A(p_input[26364]), .B(p_input[16364]), .Z(n4041) );
  AND U8083 ( .A(n4042), .B(p_input[6363]), .Z(o[6363]) );
  AND U8084 ( .A(p_input[26363]), .B(p_input[16363]), .Z(n4042) );
  AND U8085 ( .A(n4043), .B(p_input[6362]), .Z(o[6362]) );
  AND U8086 ( .A(p_input[26362]), .B(p_input[16362]), .Z(n4043) );
  AND U8087 ( .A(n4044), .B(p_input[6361]), .Z(o[6361]) );
  AND U8088 ( .A(p_input[26361]), .B(p_input[16361]), .Z(n4044) );
  AND U8089 ( .A(n4045), .B(p_input[6360]), .Z(o[6360]) );
  AND U8090 ( .A(p_input[26360]), .B(p_input[16360]), .Z(n4045) );
  AND U8091 ( .A(n4046), .B(p_input[635]), .Z(o[635]) );
  AND U8092 ( .A(p_input[20635]), .B(p_input[10635]), .Z(n4046) );
  AND U8093 ( .A(n4047), .B(p_input[6359]), .Z(o[6359]) );
  AND U8094 ( .A(p_input[26359]), .B(p_input[16359]), .Z(n4047) );
  AND U8095 ( .A(n4048), .B(p_input[6358]), .Z(o[6358]) );
  AND U8096 ( .A(p_input[26358]), .B(p_input[16358]), .Z(n4048) );
  AND U8097 ( .A(n4049), .B(p_input[6357]), .Z(o[6357]) );
  AND U8098 ( .A(p_input[26357]), .B(p_input[16357]), .Z(n4049) );
  AND U8099 ( .A(n4050), .B(p_input[6356]), .Z(o[6356]) );
  AND U8100 ( .A(p_input[26356]), .B(p_input[16356]), .Z(n4050) );
  AND U8101 ( .A(n4051), .B(p_input[6355]), .Z(o[6355]) );
  AND U8102 ( .A(p_input[26355]), .B(p_input[16355]), .Z(n4051) );
  AND U8103 ( .A(n4052), .B(p_input[6354]), .Z(o[6354]) );
  AND U8104 ( .A(p_input[26354]), .B(p_input[16354]), .Z(n4052) );
  AND U8105 ( .A(n4053), .B(p_input[6353]), .Z(o[6353]) );
  AND U8106 ( .A(p_input[26353]), .B(p_input[16353]), .Z(n4053) );
  AND U8107 ( .A(n4054), .B(p_input[6352]), .Z(o[6352]) );
  AND U8108 ( .A(p_input[26352]), .B(p_input[16352]), .Z(n4054) );
  AND U8109 ( .A(n4055), .B(p_input[6351]), .Z(o[6351]) );
  AND U8110 ( .A(p_input[26351]), .B(p_input[16351]), .Z(n4055) );
  AND U8111 ( .A(n4056), .B(p_input[6350]), .Z(o[6350]) );
  AND U8112 ( .A(p_input[26350]), .B(p_input[16350]), .Z(n4056) );
  AND U8113 ( .A(n4057), .B(p_input[634]), .Z(o[634]) );
  AND U8114 ( .A(p_input[20634]), .B(p_input[10634]), .Z(n4057) );
  AND U8115 ( .A(n4058), .B(p_input[6349]), .Z(o[6349]) );
  AND U8116 ( .A(p_input[26349]), .B(p_input[16349]), .Z(n4058) );
  AND U8117 ( .A(n4059), .B(p_input[6348]), .Z(o[6348]) );
  AND U8118 ( .A(p_input[26348]), .B(p_input[16348]), .Z(n4059) );
  AND U8119 ( .A(n4060), .B(p_input[6347]), .Z(o[6347]) );
  AND U8120 ( .A(p_input[26347]), .B(p_input[16347]), .Z(n4060) );
  AND U8121 ( .A(n4061), .B(p_input[6346]), .Z(o[6346]) );
  AND U8122 ( .A(p_input[26346]), .B(p_input[16346]), .Z(n4061) );
  AND U8123 ( .A(n4062), .B(p_input[6345]), .Z(o[6345]) );
  AND U8124 ( .A(p_input[26345]), .B(p_input[16345]), .Z(n4062) );
  AND U8125 ( .A(n4063), .B(p_input[6344]), .Z(o[6344]) );
  AND U8126 ( .A(p_input[26344]), .B(p_input[16344]), .Z(n4063) );
  AND U8127 ( .A(n4064), .B(p_input[6343]), .Z(o[6343]) );
  AND U8128 ( .A(p_input[26343]), .B(p_input[16343]), .Z(n4064) );
  AND U8129 ( .A(n4065), .B(p_input[6342]), .Z(o[6342]) );
  AND U8130 ( .A(p_input[26342]), .B(p_input[16342]), .Z(n4065) );
  AND U8131 ( .A(n4066), .B(p_input[6341]), .Z(o[6341]) );
  AND U8132 ( .A(p_input[26341]), .B(p_input[16341]), .Z(n4066) );
  AND U8133 ( .A(n4067), .B(p_input[6340]), .Z(o[6340]) );
  AND U8134 ( .A(p_input[26340]), .B(p_input[16340]), .Z(n4067) );
  AND U8135 ( .A(n4068), .B(p_input[633]), .Z(o[633]) );
  AND U8136 ( .A(p_input[20633]), .B(p_input[10633]), .Z(n4068) );
  AND U8137 ( .A(n4069), .B(p_input[6339]), .Z(o[6339]) );
  AND U8138 ( .A(p_input[26339]), .B(p_input[16339]), .Z(n4069) );
  AND U8139 ( .A(n4070), .B(p_input[6338]), .Z(o[6338]) );
  AND U8140 ( .A(p_input[26338]), .B(p_input[16338]), .Z(n4070) );
  AND U8141 ( .A(n4071), .B(p_input[6337]), .Z(o[6337]) );
  AND U8142 ( .A(p_input[26337]), .B(p_input[16337]), .Z(n4071) );
  AND U8143 ( .A(n4072), .B(p_input[6336]), .Z(o[6336]) );
  AND U8144 ( .A(p_input[26336]), .B(p_input[16336]), .Z(n4072) );
  AND U8145 ( .A(n4073), .B(p_input[6335]), .Z(o[6335]) );
  AND U8146 ( .A(p_input[26335]), .B(p_input[16335]), .Z(n4073) );
  AND U8147 ( .A(n4074), .B(p_input[6334]), .Z(o[6334]) );
  AND U8148 ( .A(p_input[26334]), .B(p_input[16334]), .Z(n4074) );
  AND U8149 ( .A(n4075), .B(p_input[6333]), .Z(o[6333]) );
  AND U8150 ( .A(p_input[26333]), .B(p_input[16333]), .Z(n4075) );
  AND U8151 ( .A(n4076), .B(p_input[6332]), .Z(o[6332]) );
  AND U8152 ( .A(p_input[26332]), .B(p_input[16332]), .Z(n4076) );
  AND U8153 ( .A(n4077), .B(p_input[6331]), .Z(o[6331]) );
  AND U8154 ( .A(p_input[26331]), .B(p_input[16331]), .Z(n4077) );
  AND U8155 ( .A(n4078), .B(p_input[6330]), .Z(o[6330]) );
  AND U8156 ( .A(p_input[26330]), .B(p_input[16330]), .Z(n4078) );
  AND U8157 ( .A(n4079), .B(p_input[632]), .Z(o[632]) );
  AND U8158 ( .A(p_input[20632]), .B(p_input[10632]), .Z(n4079) );
  AND U8159 ( .A(n4080), .B(p_input[6329]), .Z(o[6329]) );
  AND U8160 ( .A(p_input[26329]), .B(p_input[16329]), .Z(n4080) );
  AND U8161 ( .A(n4081), .B(p_input[6328]), .Z(o[6328]) );
  AND U8162 ( .A(p_input[26328]), .B(p_input[16328]), .Z(n4081) );
  AND U8163 ( .A(n4082), .B(p_input[6327]), .Z(o[6327]) );
  AND U8164 ( .A(p_input[26327]), .B(p_input[16327]), .Z(n4082) );
  AND U8165 ( .A(n4083), .B(p_input[6326]), .Z(o[6326]) );
  AND U8166 ( .A(p_input[26326]), .B(p_input[16326]), .Z(n4083) );
  AND U8167 ( .A(n4084), .B(p_input[6325]), .Z(o[6325]) );
  AND U8168 ( .A(p_input[26325]), .B(p_input[16325]), .Z(n4084) );
  AND U8169 ( .A(n4085), .B(p_input[6324]), .Z(o[6324]) );
  AND U8170 ( .A(p_input[26324]), .B(p_input[16324]), .Z(n4085) );
  AND U8171 ( .A(n4086), .B(p_input[6323]), .Z(o[6323]) );
  AND U8172 ( .A(p_input[26323]), .B(p_input[16323]), .Z(n4086) );
  AND U8173 ( .A(n4087), .B(p_input[6322]), .Z(o[6322]) );
  AND U8174 ( .A(p_input[26322]), .B(p_input[16322]), .Z(n4087) );
  AND U8175 ( .A(n4088), .B(p_input[6321]), .Z(o[6321]) );
  AND U8176 ( .A(p_input[26321]), .B(p_input[16321]), .Z(n4088) );
  AND U8177 ( .A(n4089), .B(p_input[6320]), .Z(o[6320]) );
  AND U8178 ( .A(p_input[26320]), .B(p_input[16320]), .Z(n4089) );
  AND U8179 ( .A(n4090), .B(p_input[631]), .Z(o[631]) );
  AND U8180 ( .A(p_input[20631]), .B(p_input[10631]), .Z(n4090) );
  AND U8181 ( .A(n4091), .B(p_input[6319]), .Z(o[6319]) );
  AND U8182 ( .A(p_input[26319]), .B(p_input[16319]), .Z(n4091) );
  AND U8183 ( .A(n4092), .B(p_input[6318]), .Z(o[6318]) );
  AND U8184 ( .A(p_input[26318]), .B(p_input[16318]), .Z(n4092) );
  AND U8185 ( .A(n4093), .B(p_input[6317]), .Z(o[6317]) );
  AND U8186 ( .A(p_input[26317]), .B(p_input[16317]), .Z(n4093) );
  AND U8187 ( .A(n4094), .B(p_input[6316]), .Z(o[6316]) );
  AND U8188 ( .A(p_input[26316]), .B(p_input[16316]), .Z(n4094) );
  AND U8189 ( .A(n4095), .B(p_input[6315]), .Z(o[6315]) );
  AND U8190 ( .A(p_input[26315]), .B(p_input[16315]), .Z(n4095) );
  AND U8191 ( .A(n4096), .B(p_input[6314]), .Z(o[6314]) );
  AND U8192 ( .A(p_input[26314]), .B(p_input[16314]), .Z(n4096) );
  AND U8193 ( .A(n4097), .B(p_input[6313]), .Z(o[6313]) );
  AND U8194 ( .A(p_input[26313]), .B(p_input[16313]), .Z(n4097) );
  AND U8195 ( .A(n4098), .B(p_input[6312]), .Z(o[6312]) );
  AND U8196 ( .A(p_input[26312]), .B(p_input[16312]), .Z(n4098) );
  AND U8197 ( .A(n4099), .B(p_input[6311]), .Z(o[6311]) );
  AND U8198 ( .A(p_input[26311]), .B(p_input[16311]), .Z(n4099) );
  AND U8199 ( .A(n4100), .B(p_input[6310]), .Z(o[6310]) );
  AND U8200 ( .A(p_input[26310]), .B(p_input[16310]), .Z(n4100) );
  AND U8201 ( .A(n4101), .B(p_input[630]), .Z(o[630]) );
  AND U8202 ( .A(p_input[20630]), .B(p_input[10630]), .Z(n4101) );
  AND U8203 ( .A(n4102), .B(p_input[6309]), .Z(o[6309]) );
  AND U8204 ( .A(p_input[26309]), .B(p_input[16309]), .Z(n4102) );
  AND U8205 ( .A(n4103), .B(p_input[6308]), .Z(o[6308]) );
  AND U8206 ( .A(p_input[26308]), .B(p_input[16308]), .Z(n4103) );
  AND U8207 ( .A(n4104), .B(p_input[6307]), .Z(o[6307]) );
  AND U8208 ( .A(p_input[26307]), .B(p_input[16307]), .Z(n4104) );
  AND U8209 ( .A(n4105), .B(p_input[6306]), .Z(o[6306]) );
  AND U8210 ( .A(p_input[26306]), .B(p_input[16306]), .Z(n4105) );
  AND U8211 ( .A(n4106), .B(p_input[6305]), .Z(o[6305]) );
  AND U8212 ( .A(p_input[26305]), .B(p_input[16305]), .Z(n4106) );
  AND U8213 ( .A(n4107), .B(p_input[6304]), .Z(o[6304]) );
  AND U8214 ( .A(p_input[26304]), .B(p_input[16304]), .Z(n4107) );
  AND U8215 ( .A(n4108), .B(p_input[6303]), .Z(o[6303]) );
  AND U8216 ( .A(p_input[26303]), .B(p_input[16303]), .Z(n4108) );
  AND U8217 ( .A(n4109), .B(p_input[6302]), .Z(o[6302]) );
  AND U8218 ( .A(p_input[26302]), .B(p_input[16302]), .Z(n4109) );
  AND U8219 ( .A(n4110), .B(p_input[6301]), .Z(o[6301]) );
  AND U8220 ( .A(p_input[26301]), .B(p_input[16301]), .Z(n4110) );
  AND U8221 ( .A(n4111), .B(p_input[6300]), .Z(o[6300]) );
  AND U8222 ( .A(p_input[26300]), .B(p_input[16300]), .Z(n4111) );
  AND U8223 ( .A(n4112), .B(p_input[62]), .Z(o[62]) );
  AND U8224 ( .A(p_input[20062]), .B(p_input[10062]), .Z(n4112) );
  AND U8225 ( .A(n4113), .B(p_input[629]), .Z(o[629]) );
  AND U8226 ( .A(p_input[20629]), .B(p_input[10629]), .Z(n4113) );
  AND U8227 ( .A(n4114), .B(p_input[6299]), .Z(o[6299]) );
  AND U8228 ( .A(p_input[26299]), .B(p_input[16299]), .Z(n4114) );
  AND U8229 ( .A(n4115), .B(p_input[6298]), .Z(o[6298]) );
  AND U8230 ( .A(p_input[26298]), .B(p_input[16298]), .Z(n4115) );
  AND U8231 ( .A(n4116), .B(p_input[6297]), .Z(o[6297]) );
  AND U8232 ( .A(p_input[26297]), .B(p_input[16297]), .Z(n4116) );
  AND U8233 ( .A(n4117), .B(p_input[6296]), .Z(o[6296]) );
  AND U8234 ( .A(p_input[26296]), .B(p_input[16296]), .Z(n4117) );
  AND U8235 ( .A(n4118), .B(p_input[6295]), .Z(o[6295]) );
  AND U8236 ( .A(p_input[26295]), .B(p_input[16295]), .Z(n4118) );
  AND U8237 ( .A(n4119), .B(p_input[6294]), .Z(o[6294]) );
  AND U8238 ( .A(p_input[26294]), .B(p_input[16294]), .Z(n4119) );
  AND U8239 ( .A(n4120), .B(p_input[6293]), .Z(o[6293]) );
  AND U8240 ( .A(p_input[26293]), .B(p_input[16293]), .Z(n4120) );
  AND U8241 ( .A(n4121), .B(p_input[6292]), .Z(o[6292]) );
  AND U8242 ( .A(p_input[26292]), .B(p_input[16292]), .Z(n4121) );
  AND U8243 ( .A(n4122), .B(p_input[6291]), .Z(o[6291]) );
  AND U8244 ( .A(p_input[26291]), .B(p_input[16291]), .Z(n4122) );
  AND U8245 ( .A(n4123), .B(p_input[6290]), .Z(o[6290]) );
  AND U8246 ( .A(p_input[26290]), .B(p_input[16290]), .Z(n4123) );
  AND U8247 ( .A(n4124), .B(p_input[628]), .Z(o[628]) );
  AND U8248 ( .A(p_input[20628]), .B(p_input[10628]), .Z(n4124) );
  AND U8249 ( .A(n4125), .B(p_input[6289]), .Z(o[6289]) );
  AND U8250 ( .A(p_input[26289]), .B(p_input[16289]), .Z(n4125) );
  AND U8251 ( .A(n4126), .B(p_input[6288]), .Z(o[6288]) );
  AND U8252 ( .A(p_input[26288]), .B(p_input[16288]), .Z(n4126) );
  AND U8253 ( .A(n4127), .B(p_input[6287]), .Z(o[6287]) );
  AND U8254 ( .A(p_input[26287]), .B(p_input[16287]), .Z(n4127) );
  AND U8255 ( .A(n4128), .B(p_input[6286]), .Z(o[6286]) );
  AND U8256 ( .A(p_input[26286]), .B(p_input[16286]), .Z(n4128) );
  AND U8257 ( .A(n4129), .B(p_input[6285]), .Z(o[6285]) );
  AND U8258 ( .A(p_input[26285]), .B(p_input[16285]), .Z(n4129) );
  AND U8259 ( .A(n4130), .B(p_input[6284]), .Z(o[6284]) );
  AND U8260 ( .A(p_input[26284]), .B(p_input[16284]), .Z(n4130) );
  AND U8261 ( .A(n4131), .B(p_input[6283]), .Z(o[6283]) );
  AND U8262 ( .A(p_input[26283]), .B(p_input[16283]), .Z(n4131) );
  AND U8263 ( .A(n4132), .B(p_input[6282]), .Z(o[6282]) );
  AND U8264 ( .A(p_input[26282]), .B(p_input[16282]), .Z(n4132) );
  AND U8265 ( .A(n4133), .B(p_input[6281]), .Z(o[6281]) );
  AND U8266 ( .A(p_input[26281]), .B(p_input[16281]), .Z(n4133) );
  AND U8267 ( .A(n4134), .B(p_input[6280]), .Z(o[6280]) );
  AND U8268 ( .A(p_input[26280]), .B(p_input[16280]), .Z(n4134) );
  AND U8269 ( .A(n4135), .B(p_input[627]), .Z(o[627]) );
  AND U8270 ( .A(p_input[20627]), .B(p_input[10627]), .Z(n4135) );
  AND U8271 ( .A(n4136), .B(p_input[6279]), .Z(o[6279]) );
  AND U8272 ( .A(p_input[26279]), .B(p_input[16279]), .Z(n4136) );
  AND U8273 ( .A(n4137), .B(p_input[6278]), .Z(o[6278]) );
  AND U8274 ( .A(p_input[26278]), .B(p_input[16278]), .Z(n4137) );
  AND U8275 ( .A(n4138), .B(p_input[6277]), .Z(o[6277]) );
  AND U8276 ( .A(p_input[26277]), .B(p_input[16277]), .Z(n4138) );
  AND U8277 ( .A(n4139), .B(p_input[6276]), .Z(o[6276]) );
  AND U8278 ( .A(p_input[26276]), .B(p_input[16276]), .Z(n4139) );
  AND U8279 ( .A(n4140), .B(p_input[6275]), .Z(o[6275]) );
  AND U8280 ( .A(p_input[26275]), .B(p_input[16275]), .Z(n4140) );
  AND U8281 ( .A(n4141), .B(p_input[6274]), .Z(o[6274]) );
  AND U8282 ( .A(p_input[26274]), .B(p_input[16274]), .Z(n4141) );
  AND U8283 ( .A(n4142), .B(p_input[6273]), .Z(o[6273]) );
  AND U8284 ( .A(p_input[26273]), .B(p_input[16273]), .Z(n4142) );
  AND U8285 ( .A(n4143), .B(p_input[6272]), .Z(o[6272]) );
  AND U8286 ( .A(p_input[26272]), .B(p_input[16272]), .Z(n4143) );
  AND U8287 ( .A(n4144), .B(p_input[6271]), .Z(o[6271]) );
  AND U8288 ( .A(p_input[26271]), .B(p_input[16271]), .Z(n4144) );
  AND U8289 ( .A(n4145), .B(p_input[6270]), .Z(o[6270]) );
  AND U8290 ( .A(p_input[26270]), .B(p_input[16270]), .Z(n4145) );
  AND U8291 ( .A(n4146), .B(p_input[626]), .Z(o[626]) );
  AND U8292 ( .A(p_input[20626]), .B(p_input[10626]), .Z(n4146) );
  AND U8293 ( .A(n4147), .B(p_input[6269]), .Z(o[6269]) );
  AND U8294 ( .A(p_input[26269]), .B(p_input[16269]), .Z(n4147) );
  AND U8295 ( .A(n4148), .B(p_input[6268]), .Z(o[6268]) );
  AND U8296 ( .A(p_input[26268]), .B(p_input[16268]), .Z(n4148) );
  AND U8297 ( .A(n4149), .B(p_input[6267]), .Z(o[6267]) );
  AND U8298 ( .A(p_input[26267]), .B(p_input[16267]), .Z(n4149) );
  AND U8299 ( .A(n4150), .B(p_input[6266]), .Z(o[6266]) );
  AND U8300 ( .A(p_input[26266]), .B(p_input[16266]), .Z(n4150) );
  AND U8301 ( .A(n4151), .B(p_input[6265]), .Z(o[6265]) );
  AND U8302 ( .A(p_input[26265]), .B(p_input[16265]), .Z(n4151) );
  AND U8303 ( .A(n4152), .B(p_input[6264]), .Z(o[6264]) );
  AND U8304 ( .A(p_input[26264]), .B(p_input[16264]), .Z(n4152) );
  AND U8305 ( .A(n4153), .B(p_input[6263]), .Z(o[6263]) );
  AND U8306 ( .A(p_input[26263]), .B(p_input[16263]), .Z(n4153) );
  AND U8307 ( .A(n4154), .B(p_input[6262]), .Z(o[6262]) );
  AND U8308 ( .A(p_input[26262]), .B(p_input[16262]), .Z(n4154) );
  AND U8309 ( .A(n4155), .B(p_input[6261]), .Z(o[6261]) );
  AND U8310 ( .A(p_input[26261]), .B(p_input[16261]), .Z(n4155) );
  AND U8311 ( .A(n4156), .B(p_input[6260]), .Z(o[6260]) );
  AND U8312 ( .A(p_input[26260]), .B(p_input[16260]), .Z(n4156) );
  AND U8313 ( .A(n4157), .B(p_input[625]), .Z(o[625]) );
  AND U8314 ( .A(p_input[20625]), .B(p_input[10625]), .Z(n4157) );
  AND U8315 ( .A(n4158), .B(p_input[6259]), .Z(o[6259]) );
  AND U8316 ( .A(p_input[26259]), .B(p_input[16259]), .Z(n4158) );
  AND U8317 ( .A(n4159), .B(p_input[6258]), .Z(o[6258]) );
  AND U8318 ( .A(p_input[26258]), .B(p_input[16258]), .Z(n4159) );
  AND U8319 ( .A(n4160), .B(p_input[6257]), .Z(o[6257]) );
  AND U8320 ( .A(p_input[26257]), .B(p_input[16257]), .Z(n4160) );
  AND U8321 ( .A(n4161), .B(p_input[6256]), .Z(o[6256]) );
  AND U8322 ( .A(p_input[26256]), .B(p_input[16256]), .Z(n4161) );
  AND U8323 ( .A(n4162), .B(p_input[6255]), .Z(o[6255]) );
  AND U8324 ( .A(p_input[26255]), .B(p_input[16255]), .Z(n4162) );
  AND U8325 ( .A(n4163), .B(p_input[6254]), .Z(o[6254]) );
  AND U8326 ( .A(p_input[26254]), .B(p_input[16254]), .Z(n4163) );
  AND U8327 ( .A(n4164), .B(p_input[6253]), .Z(o[6253]) );
  AND U8328 ( .A(p_input[26253]), .B(p_input[16253]), .Z(n4164) );
  AND U8329 ( .A(n4165), .B(p_input[6252]), .Z(o[6252]) );
  AND U8330 ( .A(p_input[26252]), .B(p_input[16252]), .Z(n4165) );
  AND U8331 ( .A(n4166), .B(p_input[6251]), .Z(o[6251]) );
  AND U8332 ( .A(p_input[26251]), .B(p_input[16251]), .Z(n4166) );
  AND U8333 ( .A(n4167), .B(p_input[6250]), .Z(o[6250]) );
  AND U8334 ( .A(p_input[26250]), .B(p_input[16250]), .Z(n4167) );
  AND U8335 ( .A(n4168), .B(p_input[624]), .Z(o[624]) );
  AND U8336 ( .A(p_input[20624]), .B(p_input[10624]), .Z(n4168) );
  AND U8337 ( .A(n4169), .B(p_input[6249]), .Z(o[6249]) );
  AND U8338 ( .A(p_input[26249]), .B(p_input[16249]), .Z(n4169) );
  AND U8339 ( .A(n4170), .B(p_input[6248]), .Z(o[6248]) );
  AND U8340 ( .A(p_input[26248]), .B(p_input[16248]), .Z(n4170) );
  AND U8341 ( .A(n4171), .B(p_input[6247]), .Z(o[6247]) );
  AND U8342 ( .A(p_input[26247]), .B(p_input[16247]), .Z(n4171) );
  AND U8343 ( .A(n4172), .B(p_input[6246]), .Z(o[6246]) );
  AND U8344 ( .A(p_input[26246]), .B(p_input[16246]), .Z(n4172) );
  AND U8345 ( .A(n4173), .B(p_input[6245]), .Z(o[6245]) );
  AND U8346 ( .A(p_input[26245]), .B(p_input[16245]), .Z(n4173) );
  AND U8347 ( .A(n4174), .B(p_input[6244]), .Z(o[6244]) );
  AND U8348 ( .A(p_input[26244]), .B(p_input[16244]), .Z(n4174) );
  AND U8349 ( .A(n4175), .B(p_input[6243]), .Z(o[6243]) );
  AND U8350 ( .A(p_input[26243]), .B(p_input[16243]), .Z(n4175) );
  AND U8351 ( .A(n4176), .B(p_input[6242]), .Z(o[6242]) );
  AND U8352 ( .A(p_input[26242]), .B(p_input[16242]), .Z(n4176) );
  AND U8353 ( .A(n4177), .B(p_input[6241]), .Z(o[6241]) );
  AND U8354 ( .A(p_input[26241]), .B(p_input[16241]), .Z(n4177) );
  AND U8355 ( .A(n4178), .B(p_input[6240]), .Z(o[6240]) );
  AND U8356 ( .A(p_input[26240]), .B(p_input[16240]), .Z(n4178) );
  AND U8357 ( .A(n4179), .B(p_input[623]), .Z(o[623]) );
  AND U8358 ( .A(p_input[20623]), .B(p_input[10623]), .Z(n4179) );
  AND U8359 ( .A(n4180), .B(p_input[6239]), .Z(o[6239]) );
  AND U8360 ( .A(p_input[26239]), .B(p_input[16239]), .Z(n4180) );
  AND U8361 ( .A(n4181), .B(p_input[6238]), .Z(o[6238]) );
  AND U8362 ( .A(p_input[26238]), .B(p_input[16238]), .Z(n4181) );
  AND U8363 ( .A(n4182), .B(p_input[6237]), .Z(o[6237]) );
  AND U8364 ( .A(p_input[26237]), .B(p_input[16237]), .Z(n4182) );
  AND U8365 ( .A(n4183), .B(p_input[6236]), .Z(o[6236]) );
  AND U8366 ( .A(p_input[26236]), .B(p_input[16236]), .Z(n4183) );
  AND U8367 ( .A(n4184), .B(p_input[6235]), .Z(o[6235]) );
  AND U8368 ( .A(p_input[26235]), .B(p_input[16235]), .Z(n4184) );
  AND U8369 ( .A(n4185), .B(p_input[6234]), .Z(o[6234]) );
  AND U8370 ( .A(p_input[26234]), .B(p_input[16234]), .Z(n4185) );
  AND U8371 ( .A(n4186), .B(p_input[6233]), .Z(o[6233]) );
  AND U8372 ( .A(p_input[26233]), .B(p_input[16233]), .Z(n4186) );
  AND U8373 ( .A(n4187), .B(p_input[6232]), .Z(o[6232]) );
  AND U8374 ( .A(p_input[26232]), .B(p_input[16232]), .Z(n4187) );
  AND U8375 ( .A(n4188), .B(p_input[6231]), .Z(o[6231]) );
  AND U8376 ( .A(p_input[26231]), .B(p_input[16231]), .Z(n4188) );
  AND U8377 ( .A(n4189), .B(p_input[6230]), .Z(o[6230]) );
  AND U8378 ( .A(p_input[26230]), .B(p_input[16230]), .Z(n4189) );
  AND U8379 ( .A(n4190), .B(p_input[622]), .Z(o[622]) );
  AND U8380 ( .A(p_input[20622]), .B(p_input[10622]), .Z(n4190) );
  AND U8381 ( .A(n4191), .B(p_input[6229]), .Z(o[6229]) );
  AND U8382 ( .A(p_input[26229]), .B(p_input[16229]), .Z(n4191) );
  AND U8383 ( .A(n4192), .B(p_input[6228]), .Z(o[6228]) );
  AND U8384 ( .A(p_input[26228]), .B(p_input[16228]), .Z(n4192) );
  AND U8385 ( .A(n4193), .B(p_input[6227]), .Z(o[6227]) );
  AND U8386 ( .A(p_input[26227]), .B(p_input[16227]), .Z(n4193) );
  AND U8387 ( .A(n4194), .B(p_input[6226]), .Z(o[6226]) );
  AND U8388 ( .A(p_input[26226]), .B(p_input[16226]), .Z(n4194) );
  AND U8389 ( .A(n4195), .B(p_input[6225]), .Z(o[6225]) );
  AND U8390 ( .A(p_input[26225]), .B(p_input[16225]), .Z(n4195) );
  AND U8391 ( .A(n4196), .B(p_input[6224]), .Z(o[6224]) );
  AND U8392 ( .A(p_input[26224]), .B(p_input[16224]), .Z(n4196) );
  AND U8393 ( .A(n4197), .B(p_input[6223]), .Z(o[6223]) );
  AND U8394 ( .A(p_input[26223]), .B(p_input[16223]), .Z(n4197) );
  AND U8395 ( .A(n4198), .B(p_input[6222]), .Z(o[6222]) );
  AND U8396 ( .A(p_input[26222]), .B(p_input[16222]), .Z(n4198) );
  AND U8397 ( .A(n4199), .B(p_input[6221]), .Z(o[6221]) );
  AND U8398 ( .A(p_input[26221]), .B(p_input[16221]), .Z(n4199) );
  AND U8399 ( .A(n4200), .B(p_input[6220]), .Z(o[6220]) );
  AND U8400 ( .A(p_input[26220]), .B(p_input[16220]), .Z(n4200) );
  AND U8401 ( .A(n4201), .B(p_input[621]), .Z(o[621]) );
  AND U8402 ( .A(p_input[20621]), .B(p_input[10621]), .Z(n4201) );
  AND U8403 ( .A(n4202), .B(p_input[6219]), .Z(o[6219]) );
  AND U8404 ( .A(p_input[26219]), .B(p_input[16219]), .Z(n4202) );
  AND U8405 ( .A(n4203), .B(p_input[6218]), .Z(o[6218]) );
  AND U8406 ( .A(p_input[26218]), .B(p_input[16218]), .Z(n4203) );
  AND U8407 ( .A(n4204), .B(p_input[6217]), .Z(o[6217]) );
  AND U8408 ( .A(p_input[26217]), .B(p_input[16217]), .Z(n4204) );
  AND U8409 ( .A(n4205), .B(p_input[6216]), .Z(o[6216]) );
  AND U8410 ( .A(p_input[26216]), .B(p_input[16216]), .Z(n4205) );
  AND U8411 ( .A(n4206), .B(p_input[6215]), .Z(o[6215]) );
  AND U8412 ( .A(p_input[26215]), .B(p_input[16215]), .Z(n4206) );
  AND U8413 ( .A(n4207), .B(p_input[6214]), .Z(o[6214]) );
  AND U8414 ( .A(p_input[26214]), .B(p_input[16214]), .Z(n4207) );
  AND U8415 ( .A(n4208), .B(p_input[6213]), .Z(o[6213]) );
  AND U8416 ( .A(p_input[26213]), .B(p_input[16213]), .Z(n4208) );
  AND U8417 ( .A(n4209), .B(p_input[6212]), .Z(o[6212]) );
  AND U8418 ( .A(p_input[26212]), .B(p_input[16212]), .Z(n4209) );
  AND U8419 ( .A(n4210), .B(p_input[6211]), .Z(o[6211]) );
  AND U8420 ( .A(p_input[26211]), .B(p_input[16211]), .Z(n4210) );
  AND U8421 ( .A(n4211), .B(p_input[6210]), .Z(o[6210]) );
  AND U8422 ( .A(p_input[26210]), .B(p_input[16210]), .Z(n4211) );
  AND U8423 ( .A(n4212), .B(p_input[620]), .Z(o[620]) );
  AND U8424 ( .A(p_input[20620]), .B(p_input[10620]), .Z(n4212) );
  AND U8425 ( .A(n4213), .B(p_input[6209]), .Z(o[6209]) );
  AND U8426 ( .A(p_input[26209]), .B(p_input[16209]), .Z(n4213) );
  AND U8427 ( .A(n4214), .B(p_input[6208]), .Z(o[6208]) );
  AND U8428 ( .A(p_input[26208]), .B(p_input[16208]), .Z(n4214) );
  AND U8429 ( .A(n4215), .B(p_input[6207]), .Z(o[6207]) );
  AND U8430 ( .A(p_input[26207]), .B(p_input[16207]), .Z(n4215) );
  AND U8431 ( .A(n4216), .B(p_input[6206]), .Z(o[6206]) );
  AND U8432 ( .A(p_input[26206]), .B(p_input[16206]), .Z(n4216) );
  AND U8433 ( .A(n4217), .B(p_input[6205]), .Z(o[6205]) );
  AND U8434 ( .A(p_input[26205]), .B(p_input[16205]), .Z(n4217) );
  AND U8435 ( .A(n4218), .B(p_input[6204]), .Z(o[6204]) );
  AND U8436 ( .A(p_input[26204]), .B(p_input[16204]), .Z(n4218) );
  AND U8437 ( .A(n4219), .B(p_input[6203]), .Z(o[6203]) );
  AND U8438 ( .A(p_input[26203]), .B(p_input[16203]), .Z(n4219) );
  AND U8439 ( .A(n4220), .B(p_input[6202]), .Z(o[6202]) );
  AND U8440 ( .A(p_input[26202]), .B(p_input[16202]), .Z(n4220) );
  AND U8441 ( .A(n4221), .B(p_input[6201]), .Z(o[6201]) );
  AND U8442 ( .A(p_input[26201]), .B(p_input[16201]), .Z(n4221) );
  AND U8443 ( .A(n4222), .B(p_input[6200]), .Z(o[6200]) );
  AND U8444 ( .A(p_input[26200]), .B(p_input[16200]), .Z(n4222) );
  AND U8445 ( .A(n4223), .B(p_input[61]), .Z(o[61]) );
  AND U8446 ( .A(p_input[20061]), .B(p_input[10061]), .Z(n4223) );
  AND U8447 ( .A(n4224), .B(p_input[619]), .Z(o[619]) );
  AND U8448 ( .A(p_input[20619]), .B(p_input[10619]), .Z(n4224) );
  AND U8449 ( .A(n4225), .B(p_input[6199]), .Z(o[6199]) );
  AND U8450 ( .A(p_input[26199]), .B(p_input[16199]), .Z(n4225) );
  AND U8451 ( .A(n4226), .B(p_input[6198]), .Z(o[6198]) );
  AND U8452 ( .A(p_input[26198]), .B(p_input[16198]), .Z(n4226) );
  AND U8453 ( .A(n4227), .B(p_input[6197]), .Z(o[6197]) );
  AND U8454 ( .A(p_input[26197]), .B(p_input[16197]), .Z(n4227) );
  AND U8455 ( .A(n4228), .B(p_input[6196]), .Z(o[6196]) );
  AND U8456 ( .A(p_input[26196]), .B(p_input[16196]), .Z(n4228) );
  AND U8457 ( .A(n4229), .B(p_input[6195]), .Z(o[6195]) );
  AND U8458 ( .A(p_input[26195]), .B(p_input[16195]), .Z(n4229) );
  AND U8459 ( .A(n4230), .B(p_input[6194]), .Z(o[6194]) );
  AND U8460 ( .A(p_input[26194]), .B(p_input[16194]), .Z(n4230) );
  AND U8461 ( .A(n4231), .B(p_input[6193]), .Z(o[6193]) );
  AND U8462 ( .A(p_input[26193]), .B(p_input[16193]), .Z(n4231) );
  AND U8463 ( .A(n4232), .B(p_input[6192]), .Z(o[6192]) );
  AND U8464 ( .A(p_input[26192]), .B(p_input[16192]), .Z(n4232) );
  AND U8465 ( .A(n4233), .B(p_input[6191]), .Z(o[6191]) );
  AND U8466 ( .A(p_input[26191]), .B(p_input[16191]), .Z(n4233) );
  AND U8467 ( .A(n4234), .B(p_input[6190]), .Z(o[6190]) );
  AND U8468 ( .A(p_input[26190]), .B(p_input[16190]), .Z(n4234) );
  AND U8469 ( .A(n4235), .B(p_input[618]), .Z(o[618]) );
  AND U8470 ( .A(p_input[20618]), .B(p_input[10618]), .Z(n4235) );
  AND U8471 ( .A(n4236), .B(p_input[6189]), .Z(o[6189]) );
  AND U8472 ( .A(p_input[26189]), .B(p_input[16189]), .Z(n4236) );
  AND U8473 ( .A(n4237), .B(p_input[6188]), .Z(o[6188]) );
  AND U8474 ( .A(p_input[26188]), .B(p_input[16188]), .Z(n4237) );
  AND U8475 ( .A(n4238), .B(p_input[6187]), .Z(o[6187]) );
  AND U8476 ( .A(p_input[26187]), .B(p_input[16187]), .Z(n4238) );
  AND U8477 ( .A(n4239), .B(p_input[6186]), .Z(o[6186]) );
  AND U8478 ( .A(p_input[26186]), .B(p_input[16186]), .Z(n4239) );
  AND U8479 ( .A(n4240), .B(p_input[6185]), .Z(o[6185]) );
  AND U8480 ( .A(p_input[26185]), .B(p_input[16185]), .Z(n4240) );
  AND U8481 ( .A(n4241), .B(p_input[6184]), .Z(o[6184]) );
  AND U8482 ( .A(p_input[26184]), .B(p_input[16184]), .Z(n4241) );
  AND U8483 ( .A(n4242), .B(p_input[6183]), .Z(o[6183]) );
  AND U8484 ( .A(p_input[26183]), .B(p_input[16183]), .Z(n4242) );
  AND U8485 ( .A(n4243), .B(p_input[6182]), .Z(o[6182]) );
  AND U8486 ( .A(p_input[26182]), .B(p_input[16182]), .Z(n4243) );
  AND U8487 ( .A(n4244), .B(p_input[6181]), .Z(o[6181]) );
  AND U8488 ( .A(p_input[26181]), .B(p_input[16181]), .Z(n4244) );
  AND U8489 ( .A(n4245), .B(p_input[6180]), .Z(o[6180]) );
  AND U8490 ( .A(p_input[26180]), .B(p_input[16180]), .Z(n4245) );
  AND U8491 ( .A(n4246), .B(p_input[617]), .Z(o[617]) );
  AND U8492 ( .A(p_input[20617]), .B(p_input[10617]), .Z(n4246) );
  AND U8493 ( .A(n4247), .B(p_input[6179]), .Z(o[6179]) );
  AND U8494 ( .A(p_input[26179]), .B(p_input[16179]), .Z(n4247) );
  AND U8495 ( .A(n4248), .B(p_input[6178]), .Z(o[6178]) );
  AND U8496 ( .A(p_input[26178]), .B(p_input[16178]), .Z(n4248) );
  AND U8497 ( .A(n4249), .B(p_input[6177]), .Z(o[6177]) );
  AND U8498 ( .A(p_input[26177]), .B(p_input[16177]), .Z(n4249) );
  AND U8499 ( .A(n4250), .B(p_input[6176]), .Z(o[6176]) );
  AND U8500 ( .A(p_input[26176]), .B(p_input[16176]), .Z(n4250) );
  AND U8501 ( .A(n4251), .B(p_input[6175]), .Z(o[6175]) );
  AND U8502 ( .A(p_input[26175]), .B(p_input[16175]), .Z(n4251) );
  AND U8503 ( .A(n4252), .B(p_input[6174]), .Z(o[6174]) );
  AND U8504 ( .A(p_input[26174]), .B(p_input[16174]), .Z(n4252) );
  AND U8505 ( .A(n4253), .B(p_input[6173]), .Z(o[6173]) );
  AND U8506 ( .A(p_input[26173]), .B(p_input[16173]), .Z(n4253) );
  AND U8507 ( .A(n4254), .B(p_input[6172]), .Z(o[6172]) );
  AND U8508 ( .A(p_input[26172]), .B(p_input[16172]), .Z(n4254) );
  AND U8509 ( .A(n4255), .B(p_input[6171]), .Z(o[6171]) );
  AND U8510 ( .A(p_input[26171]), .B(p_input[16171]), .Z(n4255) );
  AND U8511 ( .A(n4256), .B(p_input[6170]), .Z(o[6170]) );
  AND U8512 ( .A(p_input[26170]), .B(p_input[16170]), .Z(n4256) );
  AND U8513 ( .A(n4257), .B(p_input[616]), .Z(o[616]) );
  AND U8514 ( .A(p_input[20616]), .B(p_input[10616]), .Z(n4257) );
  AND U8515 ( .A(n4258), .B(p_input[6169]), .Z(o[6169]) );
  AND U8516 ( .A(p_input[26169]), .B(p_input[16169]), .Z(n4258) );
  AND U8517 ( .A(n4259), .B(p_input[6168]), .Z(o[6168]) );
  AND U8518 ( .A(p_input[26168]), .B(p_input[16168]), .Z(n4259) );
  AND U8519 ( .A(n4260), .B(p_input[6167]), .Z(o[6167]) );
  AND U8520 ( .A(p_input[26167]), .B(p_input[16167]), .Z(n4260) );
  AND U8521 ( .A(n4261), .B(p_input[6166]), .Z(o[6166]) );
  AND U8522 ( .A(p_input[26166]), .B(p_input[16166]), .Z(n4261) );
  AND U8523 ( .A(n4262), .B(p_input[6165]), .Z(o[6165]) );
  AND U8524 ( .A(p_input[26165]), .B(p_input[16165]), .Z(n4262) );
  AND U8525 ( .A(n4263), .B(p_input[6164]), .Z(o[6164]) );
  AND U8526 ( .A(p_input[26164]), .B(p_input[16164]), .Z(n4263) );
  AND U8527 ( .A(n4264), .B(p_input[6163]), .Z(o[6163]) );
  AND U8528 ( .A(p_input[26163]), .B(p_input[16163]), .Z(n4264) );
  AND U8529 ( .A(n4265), .B(p_input[6162]), .Z(o[6162]) );
  AND U8530 ( .A(p_input[26162]), .B(p_input[16162]), .Z(n4265) );
  AND U8531 ( .A(n4266), .B(p_input[6161]), .Z(o[6161]) );
  AND U8532 ( .A(p_input[26161]), .B(p_input[16161]), .Z(n4266) );
  AND U8533 ( .A(n4267), .B(p_input[6160]), .Z(o[6160]) );
  AND U8534 ( .A(p_input[26160]), .B(p_input[16160]), .Z(n4267) );
  AND U8535 ( .A(n4268), .B(p_input[615]), .Z(o[615]) );
  AND U8536 ( .A(p_input[20615]), .B(p_input[10615]), .Z(n4268) );
  AND U8537 ( .A(n4269), .B(p_input[6159]), .Z(o[6159]) );
  AND U8538 ( .A(p_input[26159]), .B(p_input[16159]), .Z(n4269) );
  AND U8539 ( .A(n4270), .B(p_input[6158]), .Z(o[6158]) );
  AND U8540 ( .A(p_input[26158]), .B(p_input[16158]), .Z(n4270) );
  AND U8541 ( .A(n4271), .B(p_input[6157]), .Z(o[6157]) );
  AND U8542 ( .A(p_input[26157]), .B(p_input[16157]), .Z(n4271) );
  AND U8543 ( .A(n4272), .B(p_input[6156]), .Z(o[6156]) );
  AND U8544 ( .A(p_input[26156]), .B(p_input[16156]), .Z(n4272) );
  AND U8545 ( .A(n4273), .B(p_input[6155]), .Z(o[6155]) );
  AND U8546 ( .A(p_input[26155]), .B(p_input[16155]), .Z(n4273) );
  AND U8547 ( .A(n4274), .B(p_input[6154]), .Z(o[6154]) );
  AND U8548 ( .A(p_input[26154]), .B(p_input[16154]), .Z(n4274) );
  AND U8549 ( .A(n4275), .B(p_input[6153]), .Z(o[6153]) );
  AND U8550 ( .A(p_input[26153]), .B(p_input[16153]), .Z(n4275) );
  AND U8551 ( .A(n4276), .B(p_input[6152]), .Z(o[6152]) );
  AND U8552 ( .A(p_input[26152]), .B(p_input[16152]), .Z(n4276) );
  AND U8553 ( .A(n4277), .B(p_input[6151]), .Z(o[6151]) );
  AND U8554 ( .A(p_input[26151]), .B(p_input[16151]), .Z(n4277) );
  AND U8555 ( .A(n4278), .B(p_input[6150]), .Z(o[6150]) );
  AND U8556 ( .A(p_input[26150]), .B(p_input[16150]), .Z(n4278) );
  AND U8557 ( .A(n4279), .B(p_input[614]), .Z(o[614]) );
  AND U8558 ( .A(p_input[20614]), .B(p_input[10614]), .Z(n4279) );
  AND U8559 ( .A(n4280), .B(p_input[6149]), .Z(o[6149]) );
  AND U8560 ( .A(p_input[26149]), .B(p_input[16149]), .Z(n4280) );
  AND U8561 ( .A(n4281), .B(p_input[6148]), .Z(o[6148]) );
  AND U8562 ( .A(p_input[26148]), .B(p_input[16148]), .Z(n4281) );
  AND U8563 ( .A(n4282), .B(p_input[6147]), .Z(o[6147]) );
  AND U8564 ( .A(p_input[26147]), .B(p_input[16147]), .Z(n4282) );
  AND U8565 ( .A(n4283), .B(p_input[6146]), .Z(o[6146]) );
  AND U8566 ( .A(p_input[26146]), .B(p_input[16146]), .Z(n4283) );
  AND U8567 ( .A(n4284), .B(p_input[6145]), .Z(o[6145]) );
  AND U8568 ( .A(p_input[26145]), .B(p_input[16145]), .Z(n4284) );
  AND U8569 ( .A(n4285), .B(p_input[6144]), .Z(o[6144]) );
  AND U8570 ( .A(p_input[26144]), .B(p_input[16144]), .Z(n4285) );
  AND U8571 ( .A(n4286), .B(p_input[6143]), .Z(o[6143]) );
  AND U8572 ( .A(p_input[26143]), .B(p_input[16143]), .Z(n4286) );
  AND U8573 ( .A(n4287), .B(p_input[6142]), .Z(o[6142]) );
  AND U8574 ( .A(p_input[26142]), .B(p_input[16142]), .Z(n4287) );
  AND U8575 ( .A(n4288), .B(p_input[6141]), .Z(o[6141]) );
  AND U8576 ( .A(p_input[26141]), .B(p_input[16141]), .Z(n4288) );
  AND U8577 ( .A(n4289), .B(p_input[6140]), .Z(o[6140]) );
  AND U8578 ( .A(p_input[26140]), .B(p_input[16140]), .Z(n4289) );
  AND U8579 ( .A(n4290), .B(p_input[613]), .Z(o[613]) );
  AND U8580 ( .A(p_input[20613]), .B(p_input[10613]), .Z(n4290) );
  AND U8581 ( .A(n4291), .B(p_input[6139]), .Z(o[6139]) );
  AND U8582 ( .A(p_input[26139]), .B(p_input[16139]), .Z(n4291) );
  AND U8583 ( .A(n4292), .B(p_input[6138]), .Z(o[6138]) );
  AND U8584 ( .A(p_input[26138]), .B(p_input[16138]), .Z(n4292) );
  AND U8585 ( .A(n4293), .B(p_input[6137]), .Z(o[6137]) );
  AND U8586 ( .A(p_input[26137]), .B(p_input[16137]), .Z(n4293) );
  AND U8587 ( .A(n4294), .B(p_input[6136]), .Z(o[6136]) );
  AND U8588 ( .A(p_input[26136]), .B(p_input[16136]), .Z(n4294) );
  AND U8589 ( .A(n4295), .B(p_input[6135]), .Z(o[6135]) );
  AND U8590 ( .A(p_input[26135]), .B(p_input[16135]), .Z(n4295) );
  AND U8591 ( .A(n4296), .B(p_input[6134]), .Z(o[6134]) );
  AND U8592 ( .A(p_input[26134]), .B(p_input[16134]), .Z(n4296) );
  AND U8593 ( .A(n4297), .B(p_input[6133]), .Z(o[6133]) );
  AND U8594 ( .A(p_input[26133]), .B(p_input[16133]), .Z(n4297) );
  AND U8595 ( .A(n4298), .B(p_input[6132]), .Z(o[6132]) );
  AND U8596 ( .A(p_input[26132]), .B(p_input[16132]), .Z(n4298) );
  AND U8597 ( .A(n4299), .B(p_input[6131]), .Z(o[6131]) );
  AND U8598 ( .A(p_input[26131]), .B(p_input[16131]), .Z(n4299) );
  AND U8599 ( .A(n4300), .B(p_input[6130]), .Z(o[6130]) );
  AND U8600 ( .A(p_input[26130]), .B(p_input[16130]), .Z(n4300) );
  AND U8601 ( .A(n4301), .B(p_input[612]), .Z(o[612]) );
  AND U8602 ( .A(p_input[20612]), .B(p_input[10612]), .Z(n4301) );
  AND U8603 ( .A(n4302), .B(p_input[6129]), .Z(o[6129]) );
  AND U8604 ( .A(p_input[26129]), .B(p_input[16129]), .Z(n4302) );
  AND U8605 ( .A(n4303), .B(p_input[6128]), .Z(o[6128]) );
  AND U8606 ( .A(p_input[26128]), .B(p_input[16128]), .Z(n4303) );
  AND U8607 ( .A(n4304), .B(p_input[6127]), .Z(o[6127]) );
  AND U8608 ( .A(p_input[26127]), .B(p_input[16127]), .Z(n4304) );
  AND U8609 ( .A(n4305), .B(p_input[6126]), .Z(o[6126]) );
  AND U8610 ( .A(p_input[26126]), .B(p_input[16126]), .Z(n4305) );
  AND U8611 ( .A(n4306), .B(p_input[6125]), .Z(o[6125]) );
  AND U8612 ( .A(p_input[26125]), .B(p_input[16125]), .Z(n4306) );
  AND U8613 ( .A(n4307), .B(p_input[6124]), .Z(o[6124]) );
  AND U8614 ( .A(p_input[26124]), .B(p_input[16124]), .Z(n4307) );
  AND U8615 ( .A(n4308), .B(p_input[6123]), .Z(o[6123]) );
  AND U8616 ( .A(p_input[26123]), .B(p_input[16123]), .Z(n4308) );
  AND U8617 ( .A(n4309), .B(p_input[6122]), .Z(o[6122]) );
  AND U8618 ( .A(p_input[26122]), .B(p_input[16122]), .Z(n4309) );
  AND U8619 ( .A(n4310), .B(p_input[6121]), .Z(o[6121]) );
  AND U8620 ( .A(p_input[26121]), .B(p_input[16121]), .Z(n4310) );
  AND U8621 ( .A(n4311), .B(p_input[6120]), .Z(o[6120]) );
  AND U8622 ( .A(p_input[26120]), .B(p_input[16120]), .Z(n4311) );
  AND U8623 ( .A(n4312), .B(p_input[611]), .Z(o[611]) );
  AND U8624 ( .A(p_input[20611]), .B(p_input[10611]), .Z(n4312) );
  AND U8625 ( .A(n4313), .B(p_input[6119]), .Z(o[6119]) );
  AND U8626 ( .A(p_input[26119]), .B(p_input[16119]), .Z(n4313) );
  AND U8627 ( .A(n4314), .B(p_input[6118]), .Z(o[6118]) );
  AND U8628 ( .A(p_input[26118]), .B(p_input[16118]), .Z(n4314) );
  AND U8629 ( .A(n4315), .B(p_input[6117]), .Z(o[6117]) );
  AND U8630 ( .A(p_input[26117]), .B(p_input[16117]), .Z(n4315) );
  AND U8631 ( .A(n4316), .B(p_input[6116]), .Z(o[6116]) );
  AND U8632 ( .A(p_input[26116]), .B(p_input[16116]), .Z(n4316) );
  AND U8633 ( .A(n4317), .B(p_input[6115]), .Z(o[6115]) );
  AND U8634 ( .A(p_input[26115]), .B(p_input[16115]), .Z(n4317) );
  AND U8635 ( .A(n4318), .B(p_input[6114]), .Z(o[6114]) );
  AND U8636 ( .A(p_input[26114]), .B(p_input[16114]), .Z(n4318) );
  AND U8637 ( .A(n4319), .B(p_input[6113]), .Z(o[6113]) );
  AND U8638 ( .A(p_input[26113]), .B(p_input[16113]), .Z(n4319) );
  AND U8639 ( .A(n4320), .B(p_input[6112]), .Z(o[6112]) );
  AND U8640 ( .A(p_input[26112]), .B(p_input[16112]), .Z(n4320) );
  AND U8641 ( .A(n4321), .B(p_input[6111]), .Z(o[6111]) );
  AND U8642 ( .A(p_input[26111]), .B(p_input[16111]), .Z(n4321) );
  AND U8643 ( .A(n4322), .B(p_input[6110]), .Z(o[6110]) );
  AND U8644 ( .A(p_input[26110]), .B(p_input[16110]), .Z(n4322) );
  AND U8645 ( .A(n4323), .B(p_input[610]), .Z(o[610]) );
  AND U8646 ( .A(p_input[20610]), .B(p_input[10610]), .Z(n4323) );
  AND U8647 ( .A(n4324), .B(p_input[6109]), .Z(o[6109]) );
  AND U8648 ( .A(p_input[26109]), .B(p_input[16109]), .Z(n4324) );
  AND U8649 ( .A(n4325), .B(p_input[6108]), .Z(o[6108]) );
  AND U8650 ( .A(p_input[26108]), .B(p_input[16108]), .Z(n4325) );
  AND U8651 ( .A(n4326), .B(p_input[6107]), .Z(o[6107]) );
  AND U8652 ( .A(p_input[26107]), .B(p_input[16107]), .Z(n4326) );
  AND U8653 ( .A(n4327), .B(p_input[6106]), .Z(o[6106]) );
  AND U8654 ( .A(p_input[26106]), .B(p_input[16106]), .Z(n4327) );
  AND U8655 ( .A(n4328), .B(p_input[6105]), .Z(o[6105]) );
  AND U8656 ( .A(p_input[26105]), .B(p_input[16105]), .Z(n4328) );
  AND U8657 ( .A(n4329), .B(p_input[6104]), .Z(o[6104]) );
  AND U8658 ( .A(p_input[26104]), .B(p_input[16104]), .Z(n4329) );
  AND U8659 ( .A(n4330), .B(p_input[6103]), .Z(o[6103]) );
  AND U8660 ( .A(p_input[26103]), .B(p_input[16103]), .Z(n4330) );
  AND U8661 ( .A(n4331), .B(p_input[6102]), .Z(o[6102]) );
  AND U8662 ( .A(p_input[26102]), .B(p_input[16102]), .Z(n4331) );
  AND U8663 ( .A(n4332), .B(p_input[6101]), .Z(o[6101]) );
  AND U8664 ( .A(p_input[26101]), .B(p_input[16101]), .Z(n4332) );
  AND U8665 ( .A(n4333), .B(p_input[6100]), .Z(o[6100]) );
  AND U8666 ( .A(p_input[26100]), .B(p_input[16100]), .Z(n4333) );
  AND U8667 ( .A(n4334), .B(p_input[60]), .Z(o[60]) );
  AND U8668 ( .A(p_input[20060]), .B(p_input[10060]), .Z(n4334) );
  AND U8669 ( .A(n4335), .B(p_input[609]), .Z(o[609]) );
  AND U8670 ( .A(p_input[20609]), .B(p_input[10609]), .Z(n4335) );
  AND U8671 ( .A(n4336), .B(p_input[6099]), .Z(o[6099]) );
  AND U8672 ( .A(p_input[26099]), .B(p_input[16099]), .Z(n4336) );
  AND U8673 ( .A(n4337), .B(p_input[6098]), .Z(o[6098]) );
  AND U8674 ( .A(p_input[26098]), .B(p_input[16098]), .Z(n4337) );
  AND U8675 ( .A(n4338), .B(p_input[6097]), .Z(o[6097]) );
  AND U8676 ( .A(p_input[26097]), .B(p_input[16097]), .Z(n4338) );
  AND U8677 ( .A(n4339), .B(p_input[6096]), .Z(o[6096]) );
  AND U8678 ( .A(p_input[26096]), .B(p_input[16096]), .Z(n4339) );
  AND U8679 ( .A(n4340), .B(p_input[6095]), .Z(o[6095]) );
  AND U8680 ( .A(p_input[26095]), .B(p_input[16095]), .Z(n4340) );
  AND U8681 ( .A(n4341), .B(p_input[6094]), .Z(o[6094]) );
  AND U8682 ( .A(p_input[26094]), .B(p_input[16094]), .Z(n4341) );
  AND U8683 ( .A(n4342), .B(p_input[6093]), .Z(o[6093]) );
  AND U8684 ( .A(p_input[26093]), .B(p_input[16093]), .Z(n4342) );
  AND U8685 ( .A(n4343), .B(p_input[6092]), .Z(o[6092]) );
  AND U8686 ( .A(p_input[26092]), .B(p_input[16092]), .Z(n4343) );
  AND U8687 ( .A(n4344), .B(p_input[6091]), .Z(o[6091]) );
  AND U8688 ( .A(p_input[26091]), .B(p_input[16091]), .Z(n4344) );
  AND U8689 ( .A(n4345), .B(p_input[6090]), .Z(o[6090]) );
  AND U8690 ( .A(p_input[26090]), .B(p_input[16090]), .Z(n4345) );
  AND U8691 ( .A(n4346), .B(p_input[608]), .Z(o[608]) );
  AND U8692 ( .A(p_input[20608]), .B(p_input[10608]), .Z(n4346) );
  AND U8693 ( .A(n4347), .B(p_input[6089]), .Z(o[6089]) );
  AND U8694 ( .A(p_input[26089]), .B(p_input[16089]), .Z(n4347) );
  AND U8695 ( .A(n4348), .B(p_input[6088]), .Z(o[6088]) );
  AND U8696 ( .A(p_input[26088]), .B(p_input[16088]), .Z(n4348) );
  AND U8697 ( .A(n4349), .B(p_input[6087]), .Z(o[6087]) );
  AND U8698 ( .A(p_input[26087]), .B(p_input[16087]), .Z(n4349) );
  AND U8699 ( .A(n4350), .B(p_input[6086]), .Z(o[6086]) );
  AND U8700 ( .A(p_input[26086]), .B(p_input[16086]), .Z(n4350) );
  AND U8701 ( .A(n4351), .B(p_input[6085]), .Z(o[6085]) );
  AND U8702 ( .A(p_input[26085]), .B(p_input[16085]), .Z(n4351) );
  AND U8703 ( .A(n4352), .B(p_input[6084]), .Z(o[6084]) );
  AND U8704 ( .A(p_input[26084]), .B(p_input[16084]), .Z(n4352) );
  AND U8705 ( .A(n4353), .B(p_input[6083]), .Z(o[6083]) );
  AND U8706 ( .A(p_input[26083]), .B(p_input[16083]), .Z(n4353) );
  AND U8707 ( .A(n4354), .B(p_input[6082]), .Z(o[6082]) );
  AND U8708 ( .A(p_input[26082]), .B(p_input[16082]), .Z(n4354) );
  AND U8709 ( .A(n4355), .B(p_input[6081]), .Z(o[6081]) );
  AND U8710 ( .A(p_input[26081]), .B(p_input[16081]), .Z(n4355) );
  AND U8711 ( .A(n4356), .B(p_input[6080]), .Z(o[6080]) );
  AND U8712 ( .A(p_input[26080]), .B(p_input[16080]), .Z(n4356) );
  AND U8713 ( .A(n4357), .B(p_input[607]), .Z(o[607]) );
  AND U8714 ( .A(p_input[20607]), .B(p_input[10607]), .Z(n4357) );
  AND U8715 ( .A(n4358), .B(p_input[6079]), .Z(o[6079]) );
  AND U8716 ( .A(p_input[26079]), .B(p_input[16079]), .Z(n4358) );
  AND U8717 ( .A(n4359), .B(p_input[6078]), .Z(o[6078]) );
  AND U8718 ( .A(p_input[26078]), .B(p_input[16078]), .Z(n4359) );
  AND U8719 ( .A(n4360), .B(p_input[6077]), .Z(o[6077]) );
  AND U8720 ( .A(p_input[26077]), .B(p_input[16077]), .Z(n4360) );
  AND U8721 ( .A(n4361), .B(p_input[6076]), .Z(o[6076]) );
  AND U8722 ( .A(p_input[26076]), .B(p_input[16076]), .Z(n4361) );
  AND U8723 ( .A(n4362), .B(p_input[6075]), .Z(o[6075]) );
  AND U8724 ( .A(p_input[26075]), .B(p_input[16075]), .Z(n4362) );
  AND U8725 ( .A(n4363), .B(p_input[6074]), .Z(o[6074]) );
  AND U8726 ( .A(p_input[26074]), .B(p_input[16074]), .Z(n4363) );
  AND U8727 ( .A(n4364), .B(p_input[6073]), .Z(o[6073]) );
  AND U8728 ( .A(p_input[26073]), .B(p_input[16073]), .Z(n4364) );
  AND U8729 ( .A(n4365), .B(p_input[6072]), .Z(o[6072]) );
  AND U8730 ( .A(p_input[26072]), .B(p_input[16072]), .Z(n4365) );
  AND U8731 ( .A(n4366), .B(p_input[6071]), .Z(o[6071]) );
  AND U8732 ( .A(p_input[26071]), .B(p_input[16071]), .Z(n4366) );
  AND U8733 ( .A(n4367), .B(p_input[6070]), .Z(o[6070]) );
  AND U8734 ( .A(p_input[26070]), .B(p_input[16070]), .Z(n4367) );
  AND U8735 ( .A(n4368), .B(p_input[606]), .Z(o[606]) );
  AND U8736 ( .A(p_input[20606]), .B(p_input[10606]), .Z(n4368) );
  AND U8737 ( .A(n4369), .B(p_input[6069]), .Z(o[6069]) );
  AND U8738 ( .A(p_input[26069]), .B(p_input[16069]), .Z(n4369) );
  AND U8739 ( .A(n4370), .B(p_input[6068]), .Z(o[6068]) );
  AND U8740 ( .A(p_input[26068]), .B(p_input[16068]), .Z(n4370) );
  AND U8741 ( .A(n4371), .B(p_input[6067]), .Z(o[6067]) );
  AND U8742 ( .A(p_input[26067]), .B(p_input[16067]), .Z(n4371) );
  AND U8743 ( .A(n4372), .B(p_input[6066]), .Z(o[6066]) );
  AND U8744 ( .A(p_input[26066]), .B(p_input[16066]), .Z(n4372) );
  AND U8745 ( .A(n4373), .B(p_input[6065]), .Z(o[6065]) );
  AND U8746 ( .A(p_input[26065]), .B(p_input[16065]), .Z(n4373) );
  AND U8747 ( .A(n4374), .B(p_input[6064]), .Z(o[6064]) );
  AND U8748 ( .A(p_input[26064]), .B(p_input[16064]), .Z(n4374) );
  AND U8749 ( .A(n4375), .B(p_input[6063]), .Z(o[6063]) );
  AND U8750 ( .A(p_input[26063]), .B(p_input[16063]), .Z(n4375) );
  AND U8751 ( .A(n4376), .B(p_input[6062]), .Z(o[6062]) );
  AND U8752 ( .A(p_input[26062]), .B(p_input[16062]), .Z(n4376) );
  AND U8753 ( .A(n4377), .B(p_input[6061]), .Z(o[6061]) );
  AND U8754 ( .A(p_input[26061]), .B(p_input[16061]), .Z(n4377) );
  AND U8755 ( .A(n4378), .B(p_input[6060]), .Z(o[6060]) );
  AND U8756 ( .A(p_input[26060]), .B(p_input[16060]), .Z(n4378) );
  AND U8757 ( .A(n4379), .B(p_input[605]), .Z(o[605]) );
  AND U8758 ( .A(p_input[20605]), .B(p_input[10605]), .Z(n4379) );
  AND U8759 ( .A(n4380), .B(p_input[6059]), .Z(o[6059]) );
  AND U8760 ( .A(p_input[26059]), .B(p_input[16059]), .Z(n4380) );
  AND U8761 ( .A(n4381), .B(p_input[6058]), .Z(o[6058]) );
  AND U8762 ( .A(p_input[26058]), .B(p_input[16058]), .Z(n4381) );
  AND U8763 ( .A(n4382), .B(p_input[6057]), .Z(o[6057]) );
  AND U8764 ( .A(p_input[26057]), .B(p_input[16057]), .Z(n4382) );
  AND U8765 ( .A(n4383), .B(p_input[6056]), .Z(o[6056]) );
  AND U8766 ( .A(p_input[26056]), .B(p_input[16056]), .Z(n4383) );
  AND U8767 ( .A(n4384), .B(p_input[6055]), .Z(o[6055]) );
  AND U8768 ( .A(p_input[26055]), .B(p_input[16055]), .Z(n4384) );
  AND U8769 ( .A(n4385), .B(p_input[6054]), .Z(o[6054]) );
  AND U8770 ( .A(p_input[26054]), .B(p_input[16054]), .Z(n4385) );
  AND U8771 ( .A(n4386), .B(p_input[6053]), .Z(o[6053]) );
  AND U8772 ( .A(p_input[26053]), .B(p_input[16053]), .Z(n4386) );
  AND U8773 ( .A(n4387), .B(p_input[6052]), .Z(o[6052]) );
  AND U8774 ( .A(p_input[26052]), .B(p_input[16052]), .Z(n4387) );
  AND U8775 ( .A(n4388), .B(p_input[6051]), .Z(o[6051]) );
  AND U8776 ( .A(p_input[26051]), .B(p_input[16051]), .Z(n4388) );
  AND U8777 ( .A(n4389), .B(p_input[6050]), .Z(o[6050]) );
  AND U8778 ( .A(p_input[26050]), .B(p_input[16050]), .Z(n4389) );
  AND U8779 ( .A(n4390), .B(p_input[604]), .Z(o[604]) );
  AND U8780 ( .A(p_input[20604]), .B(p_input[10604]), .Z(n4390) );
  AND U8781 ( .A(n4391), .B(p_input[6049]), .Z(o[6049]) );
  AND U8782 ( .A(p_input[26049]), .B(p_input[16049]), .Z(n4391) );
  AND U8783 ( .A(n4392), .B(p_input[6048]), .Z(o[6048]) );
  AND U8784 ( .A(p_input[26048]), .B(p_input[16048]), .Z(n4392) );
  AND U8785 ( .A(n4393), .B(p_input[6047]), .Z(o[6047]) );
  AND U8786 ( .A(p_input[26047]), .B(p_input[16047]), .Z(n4393) );
  AND U8787 ( .A(n4394), .B(p_input[6046]), .Z(o[6046]) );
  AND U8788 ( .A(p_input[26046]), .B(p_input[16046]), .Z(n4394) );
  AND U8789 ( .A(n4395), .B(p_input[6045]), .Z(o[6045]) );
  AND U8790 ( .A(p_input[26045]), .B(p_input[16045]), .Z(n4395) );
  AND U8791 ( .A(n4396), .B(p_input[6044]), .Z(o[6044]) );
  AND U8792 ( .A(p_input[26044]), .B(p_input[16044]), .Z(n4396) );
  AND U8793 ( .A(n4397), .B(p_input[6043]), .Z(o[6043]) );
  AND U8794 ( .A(p_input[26043]), .B(p_input[16043]), .Z(n4397) );
  AND U8795 ( .A(n4398), .B(p_input[6042]), .Z(o[6042]) );
  AND U8796 ( .A(p_input[26042]), .B(p_input[16042]), .Z(n4398) );
  AND U8797 ( .A(n4399), .B(p_input[6041]), .Z(o[6041]) );
  AND U8798 ( .A(p_input[26041]), .B(p_input[16041]), .Z(n4399) );
  AND U8799 ( .A(n4400), .B(p_input[6040]), .Z(o[6040]) );
  AND U8800 ( .A(p_input[26040]), .B(p_input[16040]), .Z(n4400) );
  AND U8801 ( .A(n4401), .B(p_input[603]), .Z(o[603]) );
  AND U8802 ( .A(p_input[20603]), .B(p_input[10603]), .Z(n4401) );
  AND U8803 ( .A(n4402), .B(p_input[6039]), .Z(o[6039]) );
  AND U8804 ( .A(p_input[26039]), .B(p_input[16039]), .Z(n4402) );
  AND U8805 ( .A(n4403), .B(p_input[6038]), .Z(o[6038]) );
  AND U8806 ( .A(p_input[26038]), .B(p_input[16038]), .Z(n4403) );
  AND U8807 ( .A(n4404), .B(p_input[6037]), .Z(o[6037]) );
  AND U8808 ( .A(p_input[26037]), .B(p_input[16037]), .Z(n4404) );
  AND U8809 ( .A(n4405), .B(p_input[6036]), .Z(o[6036]) );
  AND U8810 ( .A(p_input[26036]), .B(p_input[16036]), .Z(n4405) );
  AND U8811 ( .A(n4406), .B(p_input[6035]), .Z(o[6035]) );
  AND U8812 ( .A(p_input[26035]), .B(p_input[16035]), .Z(n4406) );
  AND U8813 ( .A(n4407), .B(p_input[6034]), .Z(o[6034]) );
  AND U8814 ( .A(p_input[26034]), .B(p_input[16034]), .Z(n4407) );
  AND U8815 ( .A(n4408), .B(p_input[6033]), .Z(o[6033]) );
  AND U8816 ( .A(p_input[26033]), .B(p_input[16033]), .Z(n4408) );
  AND U8817 ( .A(n4409), .B(p_input[6032]), .Z(o[6032]) );
  AND U8818 ( .A(p_input[26032]), .B(p_input[16032]), .Z(n4409) );
  AND U8819 ( .A(n4410), .B(p_input[6031]), .Z(o[6031]) );
  AND U8820 ( .A(p_input[26031]), .B(p_input[16031]), .Z(n4410) );
  AND U8821 ( .A(n4411), .B(p_input[6030]), .Z(o[6030]) );
  AND U8822 ( .A(p_input[26030]), .B(p_input[16030]), .Z(n4411) );
  AND U8823 ( .A(n4412), .B(p_input[602]), .Z(o[602]) );
  AND U8824 ( .A(p_input[20602]), .B(p_input[10602]), .Z(n4412) );
  AND U8825 ( .A(n4413), .B(p_input[6029]), .Z(o[6029]) );
  AND U8826 ( .A(p_input[26029]), .B(p_input[16029]), .Z(n4413) );
  AND U8827 ( .A(n4414), .B(p_input[6028]), .Z(o[6028]) );
  AND U8828 ( .A(p_input[26028]), .B(p_input[16028]), .Z(n4414) );
  AND U8829 ( .A(n4415), .B(p_input[6027]), .Z(o[6027]) );
  AND U8830 ( .A(p_input[26027]), .B(p_input[16027]), .Z(n4415) );
  AND U8831 ( .A(n4416), .B(p_input[6026]), .Z(o[6026]) );
  AND U8832 ( .A(p_input[26026]), .B(p_input[16026]), .Z(n4416) );
  AND U8833 ( .A(n4417), .B(p_input[6025]), .Z(o[6025]) );
  AND U8834 ( .A(p_input[26025]), .B(p_input[16025]), .Z(n4417) );
  AND U8835 ( .A(n4418), .B(p_input[6024]), .Z(o[6024]) );
  AND U8836 ( .A(p_input[26024]), .B(p_input[16024]), .Z(n4418) );
  AND U8837 ( .A(n4419), .B(p_input[6023]), .Z(o[6023]) );
  AND U8838 ( .A(p_input[26023]), .B(p_input[16023]), .Z(n4419) );
  AND U8839 ( .A(n4420), .B(p_input[6022]), .Z(o[6022]) );
  AND U8840 ( .A(p_input[26022]), .B(p_input[16022]), .Z(n4420) );
  AND U8841 ( .A(n4421), .B(p_input[6021]), .Z(o[6021]) );
  AND U8842 ( .A(p_input[26021]), .B(p_input[16021]), .Z(n4421) );
  AND U8843 ( .A(n4422), .B(p_input[6020]), .Z(o[6020]) );
  AND U8844 ( .A(p_input[26020]), .B(p_input[16020]), .Z(n4422) );
  AND U8845 ( .A(n4423), .B(p_input[601]), .Z(o[601]) );
  AND U8846 ( .A(p_input[20601]), .B(p_input[10601]), .Z(n4423) );
  AND U8847 ( .A(n4424), .B(p_input[6019]), .Z(o[6019]) );
  AND U8848 ( .A(p_input[26019]), .B(p_input[16019]), .Z(n4424) );
  AND U8849 ( .A(n4425), .B(p_input[6018]), .Z(o[6018]) );
  AND U8850 ( .A(p_input[26018]), .B(p_input[16018]), .Z(n4425) );
  AND U8851 ( .A(n4426), .B(p_input[6017]), .Z(o[6017]) );
  AND U8852 ( .A(p_input[26017]), .B(p_input[16017]), .Z(n4426) );
  AND U8853 ( .A(n4427), .B(p_input[6016]), .Z(o[6016]) );
  AND U8854 ( .A(p_input[26016]), .B(p_input[16016]), .Z(n4427) );
  AND U8855 ( .A(n4428), .B(p_input[6015]), .Z(o[6015]) );
  AND U8856 ( .A(p_input[26015]), .B(p_input[16015]), .Z(n4428) );
  AND U8857 ( .A(n4429), .B(p_input[6014]), .Z(o[6014]) );
  AND U8858 ( .A(p_input[26014]), .B(p_input[16014]), .Z(n4429) );
  AND U8859 ( .A(n4430), .B(p_input[6013]), .Z(o[6013]) );
  AND U8860 ( .A(p_input[26013]), .B(p_input[16013]), .Z(n4430) );
  AND U8861 ( .A(n4431), .B(p_input[6012]), .Z(o[6012]) );
  AND U8862 ( .A(p_input[26012]), .B(p_input[16012]), .Z(n4431) );
  AND U8863 ( .A(n4432), .B(p_input[6011]), .Z(o[6011]) );
  AND U8864 ( .A(p_input[26011]), .B(p_input[16011]), .Z(n4432) );
  AND U8865 ( .A(n4433), .B(p_input[6010]), .Z(o[6010]) );
  AND U8866 ( .A(p_input[26010]), .B(p_input[16010]), .Z(n4433) );
  AND U8867 ( .A(n4434), .B(p_input[600]), .Z(o[600]) );
  AND U8868 ( .A(p_input[20600]), .B(p_input[10600]), .Z(n4434) );
  AND U8869 ( .A(n4435), .B(p_input[6009]), .Z(o[6009]) );
  AND U8870 ( .A(p_input[26009]), .B(p_input[16009]), .Z(n4435) );
  AND U8871 ( .A(n4436), .B(p_input[6008]), .Z(o[6008]) );
  AND U8872 ( .A(p_input[26008]), .B(p_input[16008]), .Z(n4436) );
  AND U8873 ( .A(n4437), .B(p_input[6007]), .Z(o[6007]) );
  AND U8874 ( .A(p_input[26007]), .B(p_input[16007]), .Z(n4437) );
  AND U8875 ( .A(n4438), .B(p_input[6006]), .Z(o[6006]) );
  AND U8876 ( .A(p_input[26006]), .B(p_input[16006]), .Z(n4438) );
  AND U8877 ( .A(n4439), .B(p_input[6005]), .Z(o[6005]) );
  AND U8878 ( .A(p_input[26005]), .B(p_input[16005]), .Z(n4439) );
  AND U8879 ( .A(n4440), .B(p_input[6004]), .Z(o[6004]) );
  AND U8880 ( .A(p_input[26004]), .B(p_input[16004]), .Z(n4440) );
  AND U8881 ( .A(n4441), .B(p_input[6003]), .Z(o[6003]) );
  AND U8882 ( .A(p_input[26003]), .B(p_input[16003]), .Z(n4441) );
  AND U8883 ( .A(n4442), .B(p_input[6002]), .Z(o[6002]) );
  AND U8884 ( .A(p_input[26002]), .B(p_input[16002]), .Z(n4442) );
  AND U8885 ( .A(n4443), .B(p_input[6001]), .Z(o[6001]) );
  AND U8886 ( .A(p_input[26001]), .B(p_input[16001]), .Z(n4443) );
  AND U8887 ( .A(n4444), .B(p_input[6000]), .Z(o[6000]) );
  AND U8888 ( .A(p_input[26000]), .B(p_input[16000]), .Z(n4444) );
  AND U8889 ( .A(n4445), .B(p_input[5]), .Z(o[5]) );
  AND U8890 ( .A(p_input[20005]), .B(p_input[10005]), .Z(n4445) );
  AND U8891 ( .A(n4446), .B(p_input[59]), .Z(o[59]) );
  AND U8892 ( .A(p_input[20059]), .B(p_input[10059]), .Z(n4446) );
  AND U8893 ( .A(n4447), .B(p_input[599]), .Z(o[599]) );
  AND U8894 ( .A(p_input[20599]), .B(p_input[10599]), .Z(n4447) );
  AND U8895 ( .A(n4448), .B(p_input[5999]), .Z(o[5999]) );
  AND U8896 ( .A(p_input[25999]), .B(p_input[15999]), .Z(n4448) );
  AND U8897 ( .A(n4449), .B(p_input[5998]), .Z(o[5998]) );
  AND U8898 ( .A(p_input[25998]), .B(p_input[15998]), .Z(n4449) );
  AND U8899 ( .A(n4450), .B(p_input[5997]), .Z(o[5997]) );
  AND U8900 ( .A(p_input[25997]), .B(p_input[15997]), .Z(n4450) );
  AND U8901 ( .A(n4451), .B(p_input[5996]), .Z(o[5996]) );
  AND U8902 ( .A(p_input[25996]), .B(p_input[15996]), .Z(n4451) );
  AND U8903 ( .A(n4452), .B(p_input[5995]), .Z(o[5995]) );
  AND U8904 ( .A(p_input[25995]), .B(p_input[15995]), .Z(n4452) );
  AND U8905 ( .A(n4453), .B(p_input[5994]), .Z(o[5994]) );
  AND U8906 ( .A(p_input[25994]), .B(p_input[15994]), .Z(n4453) );
  AND U8907 ( .A(n4454), .B(p_input[5993]), .Z(o[5993]) );
  AND U8908 ( .A(p_input[25993]), .B(p_input[15993]), .Z(n4454) );
  AND U8909 ( .A(n4455), .B(p_input[5992]), .Z(o[5992]) );
  AND U8910 ( .A(p_input[25992]), .B(p_input[15992]), .Z(n4455) );
  AND U8911 ( .A(n4456), .B(p_input[5991]), .Z(o[5991]) );
  AND U8912 ( .A(p_input[25991]), .B(p_input[15991]), .Z(n4456) );
  AND U8913 ( .A(n4457), .B(p_input[5990]), .Z(o[5990]) );
  AND U8914 ( .A(p_input[25990]), .B(p_input[15990]), .Z(n4457) );
  AND U8915 ( .A(n4458), .B(p_input[598]), .Z(o[598]) );
  AND U8916 ( .A(p_input[20598]), .B(p_input[10598]), .Z(n4458) );
  AND U8917 ( .A(n4459), .B(p_input[5989]), .Z(o[5989]) );
  AND U8918 ( .A(p_input[25989]), .B(p_input[15989]), .Z(n4459) );
  AND U8919 ( .A(n4460), .B(p_input[5988]), .Z(o[5988]) );
  AND U8920 ( .A(p_input[25988]), .B(p_input[15988]), .Z(n4460) );
  AND U8921 ( .A(n4461), .B(p_input[5987]), .Z(o[5987]) );
  AND U8922 ( .A(p_input[25987]), .B(p_input[15987]), .Z(n4461) );
  AND U8923 ( .A(n4462), .B(p_input[5986]), .Z(o[5986]) );
  AND U8924 ( .A(p_input[25986]), .B(p_input[15986]), .Z(n4462) );
  AND U8925 ( .A(n4463), .B(p_input[5985]), .Z(o[5985]) );
  AND U8926 ( .A(p_input[25985]), .B(p_input[15985]), .Z(n4463) );
  AND U8927 ( .A(n4464), .B(p_input[5984]), .Z(o[5984]) );
  AND U8928 ( .A(p_input[25984]), .B(p_input[15984]), .Z(n4464) );
  AND U8929 ( .A(n4465), .B(p_input[5983]), .Z(o[5983]) );
  AND U8930 ( .A(p_input[25983]), .B(p_input[15983]), .Z(n4465) );
  AND U8931 ( .A(n4466), .B(p_input[5982]), .Z(o[5982]) );
  AND U8932 ( .A(p_input[25982]), .B(p_input[15982]), .Z(n4466) );
  AND U8933 ( .A(n4467), .B(p_input[5981]), .Z(o[5981]) );
  AND U8934 ( .A(p_input[25981]), .B(p_input[15981]), .Z(n4467) );
  AND U8935 ( .A(n4468), .B(p_input[5980]), .Z(o[5980]) );
  AND U8936 ( .A(p_input[25980]), .B(p_input[15980]), .Z(n4468) );
  AND U8937 ( .A(n4469), .B(p_input[597]), .Z(o[597]) );
  AND U8938 ( .A(p_input[20597]), .B(p_input[10597]), .Z(n4469) );
  AND U8939 ( .A(n4470), .B(p_input[5979]), .Z(o[5979]) );
  AND U8940 ( .A(p_input[25979]), .B(p_input[15979]), .Z(n4470) );
  AND U8941 ( .A(n4471), .B(p_input[5978]), .Z(o[5978]) );
  AND U8942 ( .A(p_input[25978]), .B(p_input[15978]), .Z(n4471) );
  AND U8943 ( .A(n4472), .B(p_input[5977]), .Z(o[5977]) );
  AND U8944 ( .A(p_input[25977]), .B(p_input[15977]), .Z(n4472) );
  AND U8945 ( .A(n4473), .B(p_input[5976]), .Z(o[5976]) );
  AND U8946 ( .A(p_input[25976]), .B(p_input[15976]), .Z(n4473) );
  AND U8947 ( .A(n4474), .B(p_input[5975]), .Z(o[5975]) );
  AND U8948 ( .A(p_input[25975]), .B(p_input[15975]), .Z(n4474) );
  AND U8949 ( .A(n4475), .B(p_input[5974]), .Z(o[5974]) );
  AND U8950 ( .A(p_input[25974]), .B(p_input[15974]), .Z(n4475) );
  AND U8951 ( .A(n4476), .B(p_input[5973]), .Z(o[5973]) );
  AND U8952 ( .A(p_input[25973]), .B(p_input[15973]), .Z(n4476) );
  AND U8953 ( .A(n4477), .B(p_input[5972]), .Z(o[5972]) );
  AND U8954 ( .A(p_input[25972]), .B(p_input[15972]), .Z(n4477) );
  AND U8955 ( .A(n4478), .B(p_input[5971]), .Z(o[5971]) );
  AND U8956 ( .A(p_input[25971]), .B(p_input[15971]), .Z(n4478) );
  AND U8957 ( .A(n4479), .B(p_input[5970]), .Z(o[5970]) );
  AND U8958 ( .A(p_input[25970]), .B(p_input[15970]), .Z(n4479) );
  AND U8959 ( .A(n4480), .B(p_input[596]), .Z(o[596]) );
  AND U8960 ( .A(p_input[20596]), .B(p_input[10596]), .Z(n4480) );
  AND U8961 ( .A(n4481), .B(p_input[5969]), .Z(o[5969]) );
  AND U8962 ( .A(p_input[25969]), .B(p_input[15969]), .Z(n4481) );
  AND U8963 ( .A(n4482), .B(p_input[5968]), .Z(o[5968]) );
  AND U8964 ( .A(p_input[25968]), .B(p_input[15968]), .Z(n4482) );
  AND U8965 ( .A(n4483), .B(p_input[5967]), .Z(o[5967]) );
  AND U8966 ( .A(p_input[25967]), .B(p_input[15967]), .Z(n4483) );
  AND U8967 ( .A(n4484), .B(p_input[5966]), .Z(o[5966]) );
  AND U8968 ( .A(p_input[25966]), .B(p_input[15966]), .Z(n4484) );
  AND U8969 ( .A(n4485), .B(p_input[5965]), .Z(o[5965]) );
  AND U8970 ( .A(p_input[25965]), .B(p_input[15965]), .Z(n4485) );
  AND U8971 ( .A(n4486), .B(p_input[5964]), .Z(o[5964]) );
  AND U8972 ( .A(p_input[25964]), .B(p_input[15964]), .Z(n4486) );
  AND U8973 ( .A(n4487), .B(p_input[5963]), .Z(o[5963]) );
  AND U8974 ( .A(p_input[25963]), .B(p_input[15963]), .Z(n4487) );
  AND U8975 ( .A(n4488), .B(p_input[5962]), .Z(o[5962]) );
  AND U8976 ( .A(p_input[25962]), .B(p_input[15962]), .Z(n4488) );
  AND U8977 ( .A(n4489), .B(p_input[5961]), .Z(o[5961]) );
  AND U8978 ( .A(p_input[25961]), .B(p_input[15961]), .Z(n4489) );
  AND U8979 ( .A(n4490), .B(p_input[5960]), .Z(o[5960]) );
  AND U8980 ( .A(p_input[25960]), .B(p_input[15960]), .Z(n4490) );
  AND U8981 ( .A(n4491), .B(p_input[595]), .Z(o[595]) );
  AND U8982 ( .A(p_input[20595]), .B(p_input[10595]), .Z(n4491) );
  AND U8983 ( .A(n4492), .B(p_input[5959]), .Z(o[5959]) );
  AND U8984 ( .A(p_input[25959]), .B(p_input[15959]), .Z(n4492) );
  AND U8985 ( .A(n4493), .B(p_input[5958]), .Z(o[5958]) );
  AND U8986 ( .A(p_input[25958]), .B(p_input[15958]), .Z(n4493) );
  AND U8987 ( .A(n4494), .B(p_input[5957]), .Z(o[5957]) );
  AND U8988 ( .A(p_input[25957]), .B(p_input[15957]), .Z(n4494) );
  AND U8989 ( .A(n4495), .B(p_input[5956]), .Z(o[5956]) );
  AND U8990 ( .A(p_input[25956]), .B(p_input[15956]), .Z(n4495) );
  AND U8991 ( .A(n4496), .B(p_input[5955]), .Z(o[5955]) );
  AND U8992 ( .A(p_input[25955]), .B(p_input[15955]), .Z(n4496) );
  AND U8993 ( .A(n4497), .B(p_input[5954]), .Z(o[5954]) );
  AND U8994 ( .A(p_input[25954]), .B(p_input[15954]), .Z(n4497) );
  AND U8995 ( .A(n4498), .B(p_input[5953]), .Z(o[5953]) );
  AND U8996 ( .A(p_input[25953]), .B(p_input[15953]), .Z(n4498) );
  AND U8997 ( .A(n4499), .B(p_input[5952]), .Z(o[5952]) );
  AND U8998 ( .A(p_input[25952]), .B(p_input[15952]), .Z(n4499) );
  AND U8999 ( .A(n4500), .B(p_input[5951]), .Z(o[5951]) );
  AND U9000 ( .A(p_input[25951]), .B(p_input[15951]), .Z(n4500) );
  AND U9001 ( .A(n4501), .B(p_input[5950]), .Z(o[5950]) );
  AND U9002 ( .A(p_input[25950]), .B(p_input[15950]), .Z(n4501) );
  AND U9003 ( .A(n4502), .B(p_input[594]), .Z(o[594]) );
  AND U9004 ( .A(p_input[20594]), .B(p_input[10594]), .Z(n4502) );
  AND U9005 ( .A(n4503), .B(p_input[5949]), .Z(o[5949]) );
  AND U9006 ( .A(p_input[25949]), .B(p_input[15949]), .Z(n4503) );
  AND U9007 ( .A(n4504), .B(p_input[5948]), .Z(o[5948]) );
  AND U9008 ( .A(p_input[25948]), .B(p_input[15948]), .Z(n4504) );
  AND U9009 ( .A(n4505), .B(p_input[5947]), .Z(o[5947]) );
  AND U9010 ( .A(p_input[25947]), .B(p_input[15947]), .Z(n4505) );
  AND U9011 ( .A(n4506), .B(p_input[5946]), .Z(o[5946]) );
  AND U9012 ( .A(p_input[25946]), .B(p_input[15946]), .Z(n4506) );
  AND U9013 ( .A(n4507), .B(p_input[5945]), .Z(o[5945]) );
  AND U9014 ( .A(p_input[25945]), .B(p_input[15945]), .Z(n4507) );
  AND U9015 ( .A(n4508), .B(p_input[5944]), .Z(o[5944]) );
  AND U9016 ( .A(p_input[25944]), .B(p_input[15944]), .Z(n4508) );
  AND U9017 ( .A(n4509), .B(p_input[5943]), .Z(o[5943]) );
  AND U9018 ( .A(p_input[25943]), .B(p_input[15943]), .Z(n4509) );
  AND U9019 ( .A(n4510), .B(p_input[5942]), .Z(o[5942]) );
  AND U9020 ( .A(p_input[25942]), .B(p_input[15942]), .Z(n4510) );
  AND U9021 ( .A(n4511), .B(p_input[5941]), .Z(o[5941]) );
  AND U9022 ( .A(p_input[25941]), .B(p_input[15941]), .Z(n4511) );
  AND U9023 ( .A(n4512), .B(p_input[5940]), .Z(o[5940]) );
  AND U9024 ( .A(p_input[25940]), .B(p_input[15940]), .Z(n4512) );
  AND U9025 ( .A(n4513), .B(p_input[593]), .Z(o[593]) );
  AND U9026 ( .A(p_input[20593]), .B(p_input[10593]), .Z(n4513) );
  AND U9027 ( .A(n4514), .B(p_input[5939]), .Z(o[5939]) );
  AND U9028 ( .A(p_input[25939]), .B(p_input[15939]), .Z(n4514) );
  AND U9029 ( .A(n4515), .B(p_input[5938]), .Z(o[5938]) );
  AND U9030 ( .A(p_input[25938]), .B(p_input[15938]), .Z(n4515) );
  AND U9031 ( .A(n4516), .B(p_input[5937]), .Z(o[5937]) );
  AND U9032 ( .A(p_input[25937]), .B(p_input[15937]), .Z(n4516) );
  AND U9033 ( .A(n4517), .B(p_input[5936]), .Z(o[5936]) );
  AND U9034 ( .A(p_input[25936]), .B(p_input[15936]), .Z(n4517) );
  AND U9035 ( .A(n4518), .B(p_input[5935]), .Z(o[5935]) );
  AND U9036 ( .A(p_input[25935]), .B(p_input[15935]), .Z(n4518) );
  AND U9037 ( .A(n4519), .B(p_input[5934]), .Z(o[5934]) );
  AND U9038 ( .A(p_input[25934]), .B(p_input[15934]), .Z(n4519) );
  AND U9039 ( .A(n4520), .B(p_input[5933]), .Z(o[5933]) );
  AND U9040 ( .A(p_input[25933]), .B(p_input[15933]), .Z(n4520) );
  AND U9041 ( .A(n4521), .B(p_input[5932]), .Z(o[5932]) );
  AND U9042 ( .A(p_input[25932]), .B(p_input[15932]), .Z(n4521) );
  AND U9043 ( .A(n4522), .B(p_input[5931]), .Z(o[5931]) );
  AND U9044 ( .A(p_input[25931]), .B(p_input[15931]), .Z(n4522) );
  AND U9045 ( .A(n4523), .B(p_input[5930]), .Z(o[5930]) );
  AND U9046 ( .A(p_input[25930]), .B(p_input[15930]), .Z(n4523) );
  AND U9047 ( .A(n4524), .B(p_input[592]), .Z(o[592]) );
  AND U9048 ( .A(p_input[20592]), .B(p_input[10592]), .Z(n4524) );
  AND U9049 ( .A(n4525), .B(p_input[5929]), .Z(o[5929]) );
  AND U9050 ( .A(p_input[25929]), .B(p_input[15929]), .Z(n4525) );
  AND U9051 ( .A(n4526), .B(p_input[5928]), .Z(o[5928]) );
  AND U9052 ( .A(p_input[25928]), .B(p_input[15928]), .Z(n4526) );
  AND U9053 ( .A(n4527), .B(p_input[5927]), .Z(o[5927]) );
  AND U9054 ( .A(p_input[25927]), .B(p_input[15927]), .Z(n4527) );
  AND U9055 ( .A(n4528), .B(p_input[5926]), .Z(o[5926]) );
  AND U9056 ( .A(p_input[25926]), .B(p_input[15926]), .Z(n4528) );
  AND U9057 ( .A(n4529), .B(p_input[5925]), .Z(o[5925]) );
  AND U9058 ( .A(p_input[25925]), .B(p_input[15925]), .Z(n4529) );
  AND U9059 ( .A(n4530), .B(p_input[5924]), .Z(o[5924]) );
  AND U9060 ( .A(p_input[25924]), .B(p_input[15924]), .Z(n4530) );
  AND U9061 ( .A(n4531), .B(p_input[5923]), .Z(o[5923]) );
  AND U9062 ( .A(p_input[25923]), .B(p_input[15923]), .Z(n4531) );
  AND U9063 ( .A(n4532), .B(p_input[5922]), .Z(o[5922]) );
  AND U9064 ( .A(p_input[25922]), .B(p_input[15922]), .Z(n4532) );
  AND U9065 ( .A(n4533), .B(p_input[5921]), .Z(o[5921]) );
  AND U9066 ( .A(p_input[25921]), .B(p_input[15921]), .Z(n4533) );
  AND U9067 ( .A(n4534), .B(p_input[5920]), .Z(o[5920]) );
  AND U9068 ( .A(p_input[25920]), .B(p_input[15920]), .Z(n4534) );
  AND U9069 ( .A(n4535), .B(p_input[591]), .Z(o[591]) );
  AND U9070 ( .A(p_input[20591]), .B(p_input[10591]), .Z(n4535) );
  AND U9071 ( .A(n4536), .B(p_input[5919]), .Z(o[5919]) );
  AND U9072 ( .A(p_input[25919]), .B(p_input[15919]), .Z(n4536) );
  AND U9073 ( .A(n4537), .B(p_input[5918]), .Z(o[5918]) );
  AND U9074 ( .A(p_input[25918]), .B(p_input[15918]), .Z(n4537) );
  AND U9075 ( .A(n4538), .B(p_input[5917]), .Z(o[5917]) );
  AND U9076 ( .A(p_input[25917]), .B(p_input[15917]), .Z(n4538) );
  AND U9077 ( .A(n4539), .B(p_input[5916]), .Z(o[5916]) );
  AND U9078 ( .A(p_input[25916]), .B(p_input[15916]), .Z(n4539) );
  AND U9079 ( .A(n4540), .B(p_input[5915]), .Z(o[5915]) );
  AND U9080 ( .A(p_input[25915]), .B(p_input[15915]), .Z(n4540) );
  AND U9081 ( .A(n4541), .B(p_input[5914]), .Z(o[5914]) );
  AND U9082 ( .A(p_input[25914]), .B(p_input[15914]), .Z(n4541) );
  AND U9083 ( .A(n4542), .B(p_input[5913]), .Z(o[5913]) );
  AND U9084 ( .A(p_input[25913]), .B(p_input[15913]), .Z(n4542) );
  AND U9085 ( .A(n4543), .B(p_input[5912]), .Z(o[5912]) );
  AND U9086 ( .A(p_input[25912]), .B(p_input[15912]), .Z(n4543) );
  AND U9087 ( .A(n4544), .B(p_input[5911]), .Z(o[5911]) );
  AND U9088 ( .A(p_input[25911]), .B(p_input[15911]), .Z(n4544) );
  AND U9089 ( .A(n4545), .B(p_input[5910]), .Z(o[5910]) );
  AND U9090 ( .A(p_input[25910]), .B(p_input[15910]), .Z(n4545) );
  AND U9091 ( .A(n4546), .B(p_input[590]), .Z(o[590]) );
  AND U9092 ( .A(p_input[20590]), .B(p_input[10590]), .Z(n4546) );
  AND U9093 ( .A(n4547), .B(p_input[5909]), .Z(o[5909]) );
  AND U9094 ( .A(p_input[25909]), .B(p_input[15909]), .Z(n4547) );
  AND U9095 ( .A(n4548), .B(p_input[5908]), .Z(o[5908]) );
  AND U9096 ( .A(p_input[25908]), .B(p_input[15908]), .Z(n4548) );
  AND U9097 ( .A(n4549), .B(p_input[5907]), .Z(o[5907]) );
  AND U9098 ( .A(p_input[25907]), .B(p_input[15907]), .Z(n4549) );
  AND U9099 ( .A(n4550), .B(p_input[5906]), .Z(o[5906]) );
  AND U9100 ( .A(p_input[25906]), .B(p_input[15906]), .Z(n4550) );
  AND U9101 ( .A(n4551), .B(p_input[5905]), .Z(o[5905]) );
  AND U9102 ( .A(p_input[25905]), .B(p_input[15905]), .Z(n4551) );
  AND U9103 ( .A(n4552), .B(p_input[5904]), .Z(o[5904]) );
  AND U9104 ( .A(p_input[25904]), .B(p_input[15904]), .Z(n4552) );
  AND U9105 ( .A(n4553), .B(p_input[5903]), .Z(o[5903]) );
  AND U9106 ( .A(p_input[25903]), .B(p_input[15903]), .Z(n4553) );
  AND U9107 ( .A(n4554), .B(p_input[5902]), .Z(o[5902]) );
  AND U9108 ( .A(p_input[25902]), .B(p_input[15902]), .Z(n4554) );
  AND U9109 ( .A(n4555), .B(p_input[5901]), .Z(o[5901]) );
  AND U9110 ( .A(p_input[25901]), .B(p_input[15901]), .Z(n4555) );
  AND U9111 ( .A(n4556), .B(p_input[5900]), .Z(o[5900]) );
  AND U9112 ( .A(p_input[25900]), .B(p_input[15900]), .Z(n4556) );
  AND U9113 ( .A(n4557), .B(p_input[58]), .Z(o[58]) );
  AND U9114 ( .A(p_input[20058]), .B(p_input[10058]), .Z(n4557) );
  AND U9115 ( .A(n4558), .B(p_input[589]), .Z(o[589]) );
  AND U9116 ( .A(p_input[20589]), .B(p_input[10589]), .Z(n4558) );
  AND U9117 ( .A(n4559), .B(p_input[5899]), .Z(o[5899]) );
  AND U9118 ( .A(p_input[25899]), .B(p_input[15899]), .Z(n4559) );
  AND U9119 ( .A(n4560), .B(p_input[5898]), .Z(o[5898]) );
  AND U9120 ( .A(p_input[25898]), .B(p_input[15898]), .Z(n4560) );
  AND U9121 ( .A(n4561), .B(p_input[5897]), .Z(o[5897]) );
  AND U9122 ( .A(p_input[25897]), .B(p_input[15897]), .Z(n4561) );
  AND U9123 ( .A(n4562), .B(p_input[5896]), .Z(o[5896]) );
  AND U9124 ( .A(p_input[25896]), .B(p_input[15896]), .Z(n4562) );
  AND U9125 ( .A(n4563), .B(p_input[5895]), .Z(o[5895]) );
  AND U9126 ( .A(p_input[25895]), .B(p_input[15895]), .Z(n4563) );
  AND U9127 ( .A(n4564), .B(p_input[5894]), .Z(o[5894]) );
  AND U9128 ( .A(p_input[25894]), .B(p_input[15894]), .Z(n4564) );
  AND U9129 ( .A(n4565), .B(p_input[5893]), .Z(o[5893]) );
  AND U9130 ( .A(p_input[25893]), .B(p_input[15893]), .Z(n4565) );
  AND U9131 ( .A(n4566), .B(p_input[5892]), .Z(o[5892]) );
  AND U9132 ( .A(p_input[25892]), .B(p_input[15892]), .Z(n4566) );
  AND U9133 ( .A(n4567), .B(p_input[5891]), .Z(o[5891]) );
  AND U9134 ( .A(p_input[25891]), .B(p_input[15891]), .Z(n4567) );
  AND U9135 ( .A(n4568), .B(p_input[5890]), .Z(o[5890]) );
  AND U9136 ( .A(p_input[25890]), .B(p_input[15890]), .Z(n4568) );
  AND U9137 ( .A(n4569), .B(p_input[588]), .Z(o[588]) );
  AND U9138 ( .A(p_input[20588]), .B(p_input[10588]), .Z(n4569) );
  AND U9139 ( .A(n4570), .B(p_input[5889]), .Z(o[5889]) );
  AND U9140 ( .A(p_input[25889]), .B(p_input[15889]), .Z(n4570) );
  AND U9141 ( .A(n4571), .B(p_input[5888]), .Z(o[5888]) );
  AND U9142 ( .A(p_input[25888]), .B(p_input[15888]), .Z(n4571) );
  AND U9143 ( .A(n4572), .B(p_input[5887]), .Z(o[5887]) );
  AND U9144 ( .A(p_input[25887]), .B(p_input[15887]), .Z(n4572) );
  AND U9145 ( .A(n4573), .B(p_input[5886]), .Z(o[5886]) );
  AND U9146 ( .A(p_input[25886]), .B(p_input[15886]), .Z(n4573) );
  AND U9147 ( .A(n4574), .B(p_input[5885]), .Z(o[5885]) );
  AND U9148 ( .A(p_input[25885]), .B(p_input[15885]), .Z(n4574) );
  AND U9149 ( .A(n4575), .B(p_input[5884]), .Z(o[5884]) );
  AND U9150 ( .A(p_input[25884]), .B(p_input[15884]), .Z(n4575) );
  AND U9151 ( .A(n4576), .B(p_input[5883]), .Z(o[5883]) );
  AND U9152 ( .A(p_input[25883]), .B(p_input[15883]), .Z(n4576) );
  AND U9153 ( .A(n4577), .B(p_input[5882]), .Z(o[5882]) );
  AND U9154 ( .A(p_input[25882]), .B(p_input[15882]), .Z(n4577) );
  AND U9155 ( .A(n4578), .B(p_input[5881]), .Z(o[5881]) );
  AND U9156 ( .A(p_input[25881]), .B(p_input[15881]), .Z(n4578) );
  AND U9157 ( .A(n4579), .B(p_input[5880]), .Z(o[5880]) );
  AND U9158 ( .A(p_input[25880]), .B(p_input[15880]), .Z(n4579) );
  AND U9159 ( .A(n4580), .B(p_input[587]), .Z(o[587]) );
  AND U9160 ( .A(p_input[20587]), .B(p_input[10587]), .Z(n4580) );
  AND U9161 ( .A(n4581), .B(p_input[5879]), .Z(o[5879]) );
  AND U9162 ( .A(p_input[25879]), .B(p_input[15879]), .Z(n4581) );
  AND U9163 ( .A(n4582), .B(p_input[5878]), .Z(o[5878]) );
  AND U9164 ( .A(p_input[25878]), .B(p_input[15878]), .Z(n4582) );
  AND U9165 ( .A(n4583), .B(p_input[5877]), .Z(o[5877]) );
  AND U9166 ( .A(p_input[25877]), .B(p_input[15877]), .Z(n4583) );
  AND U9167 ( .A(n4584), .B(p_input[5876]), .Z(o[5876]) );
  AND U9168 ( .A(p_input[25876]), .B(p_input[15876]), .Z(n4584) );
  AND U9169 ( .A(n4585), .B(p_input[5875]), .Z(o[5875]) );
  AND U9170 ( .A(p_input[25875]), .B(p_input[15875]), .Z(n4585) );
  AND U9171 ( .A(n4586), .B(p_input[5874]), .Z(o[5874]) );
  AND U9172 ( .A(p_input[25874]), .B(p_input[15874]), .Z(n4586) );
  AND U9173 ( .A(n4587), .B(p_input[5873]), .Z(o[5873]) );
  AND U9174 ( .A(p_input[25873]), .B(p_input[15873]), .Z(n4587) );
  AND U9175 ( .A(n4588), .B(p_input[5872]), .Z(o[5872]) );
  AND U9176 ( .A(p_input[25872]), .B(p_input[15872]), .Z(n4588) );
  AND U9177 ( .A(n4589), .B(p_input[5871]), .Z(o[5871]) );
  AND U9178 ( .A(p_input[25871]), .B(p_input[15871]), .Z(n4589) );
  AND U9179 ( .A(n4590), .B(p_input[5870]), .Z(o[5870]) );
  AND U9180 ( .A(p_input[25870]), .B(p_input[15870]), .Z(n4590) );
  AND U9181 ( .A(n4591), .B(p_input[586]), .Z(o[586]) );
  AND U9182 ( .A(p_input[20586]), .B(p_input[10586]), .Z(n4591) );
  AND U9183 ( .A(n4592), .B(p_input[5869]), .Z(o[5869]) );
  AND U9184 ( .A(p_input[25869]), .B(p_input[15869]), .Z(n4592) );
  AND U9185 ( .A(n4593), .B(p_input[5868]), .Z(o[5868]) );
  AND U9186 ( .A(p_input[25868]), .B(p_input[15868]), .Z(n4593) );
  AND U9187 ( .A(n4594), .B(p_input[5867]), .Z(o[5867]) );
  AND U9188 ( .A(p_input[25867]), .B(p_input[15867]), .Z(n4594) );
  AND U9189 ( .A(n4595), .B(p_input[5866]), .Z(o[5866]) );
  AND U9190 ( .A(p_input[25866]), .B(p_input[15866]), .Z(n4595) );
  AND U9191 ( .A(n4596), .B(p_input[5865]), .Z(o[5865]) );
  AND U9192 ( .A(p_input[25865]), .B(p_input[15865]), .Z(n4596) );
  AND U9193 ( .A(n4597), .B(p_input[5864]), .Z(o[5864]) );
  AND U9194 ( .A(p_input[25864]), .B(p_input[15864]), .Z(n4597) );
  AND U9195 ( .A(n4598), .B(p_input[5863]), .Z(o[5863]) );
  AND U9196 ( .A(p_input[25863]), .B(p_input[15863]), .Z(n4598) );
  AND U9197 ( .A(n4599), .B(p_input[5862]), .Z(o[5862]) );
  AND U9198 ( .A(p_input[25862]), .B(p_input[15862]), .Z(n4599) );
  AND U9199 ( .A(n4600), .B(p_input[5861]), .Z(o[5861]) );
  AND U9200 ( .A(p_input[25861]), .B(p_input[15861]), .Z(n4600) );
  AND U9201 ( .A(n4601), .B(p_input[5860]), .Z(o[5860]) );
  AND U9202 ( .A(p_input[25860]), .B(p_input[15860]), .Z(n4601) );
  AND U9203 ( .A(n4602), .B(p_input[585]), .Z(o[585]) );
  AND U9204 ( .A(p_input[20585]), .B(p_input[10585]), .Z(n4602) );
  AND U9205 ( .A(n4603), .B(p_input[5859]), .Z(o[5859]) );
  AND U9206 ( .A(p_input[25859]), .B(p_input[15859]), .Z(n4603) );
  AND U9207 ( .A(n4604), .B(p_input[5858]), .Z(o[5858]) );
  AND U9208 ( .A(p_input[25858]), .B(p_input[15858]), .Z(n4604) );
  AND U9209 ( .A(n4605), .B(p_input[5857]), .Z(o[5857]) );
  AND U9210 ( .A(p_input[25857]), .B(p_input[15857]), .Z(n4605) );
  AND U9211 ( .A(n4606), .B(p_input[5856]), .Z(o[5856]) );
  AND U9212 ( .A(p_input[25856]), .B(p_input[15856]), .Z(n4606) );
  AND U9213 ( .A(n4607), .B(p_input[5855]), .Z(o[5855]) );
  AND U9214 ( .A(p_input[25855]), .B(p_input[15855]), .Z(n4607) );
  AND U9215 ( .A(n4608), .B(p_input[5854]), .Z(o[5854]) );
  AND U9216 ( .A(p_input[25854]), .B(p_input[15854]), .Z(n4608) );
  AND U9217 ( .A(n4609), .B(p_input[5853]), .Z(o[5853]) );
  AND U9218 ( .A(p_input[25853]), .B(p_input[15853]), .Z(n4609) );
  AND U9219 ( .A(n4610), .B(p_input[5852]), .Z(o[5852]) );
  AND U9220 ( .A(p_input[25852]), .B(p_input[15852]), .Z(n4610) );
  AND U9221 ( .A(n4611), .B(p_input[5851]), .Z(o[5851]) );
  AND U9222 ( .A(p_input[25851]), .B(p_input[15851]), .Z(n4611) );
  AND U9223 ( .A(n4612), .B(p_input[5850]), .Z(o[5850]) );
  AND U9224 ( .A(p_input[25850]), .B(p_input[15850]), .Z(n4612) );
  AND U9225 ( .A(n4613), .B(p_input[584]), .Z(o[584]) );
  AND U9226 ( .A(p_input[20584]), .B(p_input[10584]), .Z(n4613) );
  AND U9227 ( .A(n4614), .B(p_input[5849]), .Z(o[5849]) );
  AND U9228 ( .A(p_input[25849]), .B(p_input[15849]), .Z(n4614) );
  AND U9229 ( .A(n4615), .B(p_input[5848]), .Z(o[5848]) );
  AND U9230 ( .A(p_input[25848]), .B(p_input[15848]), .Z(n4615) );
  AND U9231 ( .A(n4616), .B(p_input[5847]), .Z(o[5847]) );
  AND U9232 ( .A(p_input[25847]), .B(p_input[15847]), .Z(n4616) );
  AND U9233 ( .A(n4617), .B(p_input[5846]), .Z(o[5846]) );
  AND U9234 ( .A(p_input[25846]), .B(p_input[15846]), .Z(n4617) );
  AND U9235 ( .A(n4618), .B(p_input[5845]), .Z(o[5845]) );
  AND U9236 ( .A(p_input[25845]), .B(p_input[15845]), .Z(n4618) );
  AND U9237 ( .A(n4619), .B(p_input[5844]), .Z(o[5844]) );
  AND U9238 ( .A(p_input[25844]), .B(p_input[15844]), .Z(n4619) );
  AND U9239 ( .A(n4620), .B(p_input[5843]), .Z(o[5843]) );
  AND U9240 ( .A(p_input[25843]), .B(p_input[15843]), .Z(n4620) );
  AND U9241 ( .A(n4621), .B(p_input[5842]), .Z(o[5842]) );
  AND U9242 ( .A(p_input[25842]), .B(p_input[15842]), .Z(n4621) );
  AND U9243 ( .A(n4622), .B(p_input[5841]), .Z(o[5841]) );
  AND U9244 ( .A(p_input[25841]), .B(p_input[15841]), .Z(n4622) );
  AND U9245 ( .A(n4623), .B(p_input[5840]), .Z(o[5840]) );
  AND U9246 ( .A(p_input[25840]), .B(p_input[15840]), .Z(n4623) );
  AND U9247 ( .A(n4624), .B(p_input[583]), .Z(o[583]) );
  AND U9248 ( .A(p_input[20583]), .B(p_input[10583]), .Z(n4624) );
  AND U9249 ( .A(n4625), .B(p_input[5839]), .Z(o[5839]) );
  AND U9250 ( .A(p_input[25839]), .B(p_input[15839]), .Z(n4625) );
  AND U9251 ( .A(n4626), .B(p_input[5838]), .Z(o[5838]) );
  AND U9252 ( .A(p_input[25838]), .B(p_input[15838]), .Z(n4626) );
  AND U9253 ( .A(n4627), .B(p_input[5837]), .Z(o[5837]) );
  AND U9254 ( .A(p_input[25837]), .B(p_input[15837]), .Z(n4627) );
  AND U9255 ( .A(n4628), .B(p_input[5836]), .Z(o[5836]) );
  AND U9256 ( .A(p_input[25836]), .B(p_input[15836]), .Z(n4628) );
  AND U9257 ( .A(n4629), .B(p_input[5835]), .Z(o[5835]) );
  AND U9258 ( .A(p_input[25835]), .B(p_input[15835]), .Z(n4629) );
  AND U9259 ( .A(n4630), .B(p_input[5834]), .Z(o[5834]) );
  AND U9260 ( .A(p_input[25834]), .B(p_input[15834]), .Z(n4630) );
  AND U9261 ( .A(n4631), .B(p_input[5833]), .Z(o[5833]) );
  AND U9262 ( .A(p_input[25833]), .B(p_input[15833]), .Z(n4631) );
  AND U9263 ( .A(n4632), .B(p_input[5832]), .Z(o[5832]) );
  AND U9264 ( .A(p_input[25832]), .B(p_input[15832]), .Z(n4632) );
  AND U9265 ( .A(n4633), .B(p_input[5831]), .Z(o[5831]) );
  AND U9266 ( .A(p_input[25831]), .B(p_input[15831]), .Z(n4633) );
  AND U9267 ( .A(n4634), .B(p_input[5830]), .Z(o[5830]) );
  AND U9268 ( .A(p_input[25830]), .B(p_input[15830]), .Z(n4634) );
  AND U9269 ( .A(n4635), .B(p_input[582]), .Z(o[582]) );
  AND U9270 ( .A(p_input[20582]), .B(p_input[10582]), .Z(n4635) );
  AND U9271 ( .A(n4636), .B(p_input[5829]), .Z(o[5829]) );
  AND U9272 ( .A(p_input[25829]), .B(p_input[15829]), .Z(n4636) );
  AND U9273 ( .A(n4637), .B(p_input[5828]), .Z(o[5828]) );
  AND U9274 ( .A(p_input[25828]), .B(p_input[15828]), .Z(n4637) );
  AND U9275 ( .A(n4638), .B(p_input[5827]), .Z(o[5827]) );
  AND U9276 ( .A(p_input[25827]), .B(p_input[15827]), .Z(n4638) );
  AND U9277 ( .A(n4639), .B(p_input[5826]), .Z(o[5826]) );
  AND U9278 ( .A(p_input[25826]), .B(p_input[15826]), .Z(n4639) );
  AND U9279 ( .A(n4640), .B(p_input[5825]), .Z(o[5825]) );
  AND U9280 ( .A(p_input[25825]), .B(p_input[15825]), .Z(n4640) );
  AND U9281 ( .A(n4641), .B(p_input[5824]), .Z(o[5824]) );
  AND U9282 ( .A(p_input[25824]), .B(p_input[15824]), .Z(n4641) );
  AND U9283 ( .A(n4642), .B(p_input[5823]), .Z(o[5823]) );
  AND U9284 ( .A(p_input[25823]), .B(p_input[15823]), .Z(n4642) );
  AND U9285 ( .A(n4643), .B(p_input[5822]), .Z(o[5822]) );
  AND U9286 ( .A(p_input[25822]), .B(p_input[15822]), .Z(n4643) );
  AND U9287 ( .A(n4644), .B(p_input[5821]), .Z(o[5821]) );
  AND U9288 ( .A(p_input[25821]), .B(p_input[15821]), .Z(n4644) );
  AND U9289 ( .A(n4645), .B(p_input[5820]), .Z(o[5820]) );
  AND U9290 ( .A(p_input[25820]), .B(p_input[15820]), .Z(n4645) );
  AND U9291 ( .A(n4646), .B(p_input[581]), .Z(o[581]) );
  AND U9292 ( .A(p_input[20581]), .B(p_input[10581]), .Z(n4646) );
  AND U9293 ( .A(n4647), .B(p_input[5819]), .Z(o[5819]) );
  AND U9294 ( .A(p_input[25819]), .B(p_input[15819]), .Z(n4647) );
  AND U9295 ( .A(n4648), .B(p_input[5818]), .Z(o[5818]) );
  AND U9296 ( .A(p_input[25818]), .B(p_input[15818]), .Z(n4648) );
  AND U9297 ( .A(n4649), .B(p_input[5817]), .Z(o[5817]) );
  AND U9298 ( .A(p_input[25817]), .B(p_input[15817]), .Z(n4649) );
  AND U9299 ( .A(n4650), .B(p_input[5816]), .Z(o[5816]) );
  AND U9300 ( .A(p_input[25816]), .B(p_input[15816]), .Z(n4650) );
  AND U9301 ( .A(n4651), .B(p_input[5815]), .Z(o[5815]) );
  AND U9302 ( .A(p_input[25815]), .B(p_input[15815]), .Z(n4651) );
  AND U9303 ( .A(n4652), .B(p_input[5814]), .Z(o[5814]) );
  AND U9304 ( .A(p_input[25814]), .B(p_input[15814]), .Z(n4652) );
  AND U9305 ( .A(n4653), .B(p_input[5813]), .Z(o[5813]) );
  AND U9306 ( .A(p_input[25813]), .B(p_input[15813]), .Z(n4653) );
  AND U9307 ( .A(n4654), .B(p_input[5812]), .Z(o[5812]) );
  AND U9308 ( .A(p_input[25812]), .B(p_input[15812]), .Z(n4654) );
  AND U9309 ( .A(n4655), .B(p_input[5811]), .Z(o[5811]) );
  AND U9310 ( .A(p_input[25811]), .B(p_input[15811]), .Z(n4655) );
  AND U9311 ( .A(n4656), .B(p_input[5810]), .Z(o[5810]) );
  AND U9312 ( .A(p_input[25810]), .B(p_input[15810]), .Z(n4656) );
  AND U9313 ( .A(n4657), .B(p_input[580]), .Z(o[580]) );
  AND U9314 ( .A(p_input[20580]), .B(p_input[10580]), .Z(n4657) );
  AND U9315 ( .A(n4658), .B(p_input[5809]), .Z(o[5809]) );
  AND U9316 ( .A(p_input[25809]), .B(p_input[15809]), .Z(n4658) );
  AND U9317 ( .A(n4659), .B(p_input[5808]), .Z(o[5808]) );
  AND U9318 ( .A(p_input[25808]), .B(p_input[15808]), .Z(n4659) );
  AND U9319 ( .A(n4660), .B(p_input[5807]), .Z(o[5807]) );
  AND U9320 ( .A(p_input[25807]), .B(p_input[15807]), .Z(n4660) );
  AND U9321 ( .A(n4661), .B(p_input[5806]), .Z(o[5806]) );
  AND U9322 ( .A(p_input[25806]), .B(p_input[15806]), .Z(n4661) );
  AND U9323 ( .A(n4662), .B(p_input[5805]), .Z(o[5805]) );
  AND U9324 ( .A(p_input[25805]), .B(p_input[15805]), .Z(n4662) );
  AND U9325 ( .A(n4663), .B(p_input[5804]), .Z(o[5804]) );
  AND U9326 ( .A(p_input[25804]), .B(p_input[15804]), .Z(n4663) );
  AND U9327 ( .A(n4664), .B(p_input[5803]), .Z(o[5803]) );
  AND U9328 ( .A(p_input[25803]), .B(p_input[15803]), .Z(n4664) );
  AND U9329 ( .A(n4665), .B(p_input[5802]), .Z(o[5802]) );
  AND U9330 ( .A(p_input[25802]), .B(p_input[15802]), .Z(n4665) );
  AND U9331 ( .A(n4666), .B(p_input[5801]), .Z(o[5801]) );
  AND U9332 ( .A(p_input[25801]), .B(p_input[15801]), .Z(n4666) );
  AND U9333 ( .A(n4667), .B(p_input[5800]), .Z(o[5800]) );
  AND U9334 ( .A(p_input[25800]), .B(p_input[15800]), .Z(n4667) );
  AND U9335 ( .A(n4668), .B(p_input[57]), .Z(o[57]) );
  AND U9336 ( .A(p_input[20057]), .B(p_input[10057]), .Z(n4668) );
  AND U9337 ( .A(n4669), .B(p_input[579]), .Z(o[579]) );
  AND U9338 ( .A(p_input[20579]), .B(p_input[10579]), .Z(n4669) );
  AND U9339 ( .A(n4670), .B(p_input[5799]), .Z(o[5799]) );
  AND U9340 ( .A(p_input[25799]), .B(p_input[15799]), .Z(n4670) );
  AND U9341 ( .A(n4671), .B(p_input[5798]), .Z(o[5798]) );
  AND U9342 ( .A(p_input[25798]), .B(p_input[15798]), .Z(n4671) );
  AND U9343 ( .A(n4672), .B(p_input[5797]), .Z(o[5797]) );
  AND U9344 ( .A(p_input[25797]), .B(p_input[15797]), .Z(n4672) );
  AND U9345 ( .A(n4673), .B(p_input[5796]), .Z(o[5796]) );
  AND U9346 ( .A(p_input[25796]), .B(p_input[15796]), .Z(n4673) );
  AND U9347 ( .A(n4674), .B(p_input[5795]), .Z(o[5795]) );
  AND U9348 ( .A(p_input[25795]), .B(p_input[15795]), .Z(n4674) );
  AND U9349 ( .A(n4675), .B(p_input[5794]), .Z(o[5794]) );
  AND U9350 ( .A(p_input[25794]), .B(p_input[15794]), .Z(n4675) );
  AND U9351 ( .A(n4676), .B(p_input[5793]), .Z(o[5793]) );
  AND U9352 ( .A(p_input[25793]), .B(p_input[15793]), .Z(n4676) );
  AND U9353 ( .A(n4677), .B(p_input[5792]), .Z(o[5792]) );
  AND U9354 ( .A(p_input[25792]), .B(p_input[15792]), .Z(n4677) );
  AND U9355 ( .A(n4678), .B(p_input[5791]), .Z(o[5791]) );
  AND U9356 ( .A(p_input[25791]), .B(p_input[15791]), .Z(n4678) );
  AND U9357 ( .A(n4679), .B(p_input[5790]), .Z(o[5790]) );
  AND U9358 ( .A(p_input[25790]), .B(p_input[15790]), .Z(n4679) );
  AND U9359 ( .A(n4680), .B(p_input[578]), .Z(o[578]) );
  AND U9360 ( .A(p_input[20578]), .B(p_input[10578]), .Z(n4680) );
  AND U9361 ( .A(n4681), .B(p_input[5789]), .Z(o[5789]) );
  AND U9362 ( .A(p_input[25789]), .B(p_input[15789]), .Z(n4681) );
  AND U9363 ( .A(n4682), .B(p_input[5788]), .Z(o[5788]) );
  AND U9364 ( .A(p_input[25788]), .B(p_input[15788]), .Z(n4682) );
  AND U9365 ( .A(n4683), .B(p_input[5787]), .Z(o[5787]) );
  AND U9366 ( .A(p_input[25787]), .B(p_input[15787]), .Z(n4683) );
  AND U9367 ( .A(n4684), .B(p_input[5786]), .Z(o[5786]) );
  AND U9368 ( .A(p_input[25786]), .B(p_input[15786]), .Z(n4684) );
  AND U9369 ( .A(n4685), .B(p_input[5785]), .Z(o[5785]) );
  AND U9370 ( .A(p_input[25785]), .B(p_input[15785]), .Z(n4685) );
  AND U9371 ( .A(n4686), .B(p_input[5784]), .Z(o[5784]) );
  AND U9372 ( .A(p_input[25784]), .B(p_input[15784]), .Z(n4686) );
  AND U9373 ( .A(n4687), .B(p_input[5783]), .Z(o[5783]) );
  AND U9374 ( .A(p_input[25783]), .B(p_input[15783]), .Z(n4687) );
  AND U9375 ( .A(n4688), .B(p_input[5782]), .Z(o[5782]) );
  AND U9376 ( .A(p_input[25782]), .B(p_input[15782]), .Z(n4688) );
  AND U9377 ( .A(n4689), .B(p_input[5781]), .Z(o[5781]) );
  AND U9378 ( .A(p_input[25781]), .B(p_input[15781]), .Z(n4689) );
  AND U9379 ( .A(n4690), .B(p_input[5780]), .Z(o[5780]) );
  AND U9380 ( .A(p_input[25780]), .B(p_input[15780]), .Z(n4690) );
  AND U9381 ( .A(n4691), .B(p_input[577]), .Z(o[577]) );
  AND U9382 ( .A(p_input[20577]), .B(p_input[10577]), .Z(n4691) );
  AND U9383 ( .A(n4692), .B(p_input[5779]), .Z(o[5779]) );
  AND U9384 ( .A(p_input[25779]), .B(p_input[15779]), .Z(n4692) );
  AND U9385 ( .A(n4693), .B(p_input[5778]), .Z(o[5778]) );
  AND U9386 ( .A(p_input[25778]), .B(p_input[15778]), .Z(n4693) );
  AND U9387 ( .A(n4694), .B(p_input[5777]), .Z(o[5777]) );
  AND U9388 ( .A(p_input[25777]), .B(p_input[15777]), .Z(n4694) );
  AND U9389 ( .A(n4695), .B(p_input[5776]), .Z(o[5776]) );
  AND U9390 ( .A(p_input[25776]), .B(p_input[15776]), .Z(n4695) );
  AND U9391 ( .A(n4696), .B(p_input[5775]), .Z(o[5775]) );
  AND U9392 ( .A(p_input[25775]), .B(p_input[15775]), .Z(n4696) );
  AND U9393 ( .A(n4697), .B(p_input[5774]), .Z(o[5774]) );
  AND U9394 ( .A(p_input[25774]), .B(p_input[15774]), .Z(n4697) );
  AND U9395 ( .A(n4698), .B(p_input[5773]), .Z(o[5773]) );
  AND U9396 ( .A(p_input[25773]), .B(p_input[15773]), .Z(n4698) );
  AND U9397 ( .A(n4699), .B(p_input[5772]), .Z(o[5772]) );
  AND U9398 ( .A(p_input[25772]), .B(p_input[15772]), .Z(n4699) );
  AND U9399 ( .A(n4700), .B(p_input[5771]), .Z(o[5771]) );
  AND U9400 ( .A(p_input[25771]), .B(p_input[15771]), .Z(n4700) );
  AND U9401 ( .A(n4701), .B(p_input[5770]), .Z(o[5770]) );
  AND U9402 ( .A(p_input[25770]), .B(p_input[15770]), .Z(n4701) );
  AND U9403 ( .A(n4702), .B(p_input[576]), .Z(o[576]) );
  AND U9404 ( .A(p_input[20576]), .B(p_input[10576]), .Z(n4702) );
  AND U9405 ( .A(n4703), .B(p_input[5769]), .Z(o[5769]) );
  AND U9406 ( .A(p_input[25769]), .B(p_input[15769]), .Z(n4703) );
  AND U9407 ( .A(n4704), .B(p_input[5768]), .Z(o[5768]) );
  AND U9408 ( .A(p_input[25768]), .B(p_input[15768]), .Z(n4704) );
  AND U9409 ( .A(n4705), .B(p_input[5767]), .Z(o[5767]) );
  AND U9410 ( .A(p_input[25767]), .B(p_input[15767]), .Z(n4705) );
  AND U9411 ( .A(n4706), .B(p_input[5766]), .Z(o[5766]) );
  AND U9412 ( .A(p_input[25766]), .B(p_input[15766]), .Z(n4706) );
  AND U9413 ( .A(n4707), .B(p_input[5765]), .Z(o[5765]) );
  AND U9414 ( .A(p_input[25765]), .B(p_input[15765]), .Z(n4707) );
  AND U9415 ( .A(n4708), .B(p_input[5764]), .Z(o[5764]) );
  AND U9416 ( .A(p_input[25764]), .B(p_input[15764]), .Z(n4708) );
  AND U9417 ( .A(n4709), .B(p_input[5763]), .Z(o[5763]) );
  AND U9418 ( .A(p_input[25763]), .B(p_input[15763]), .Z(n4709) );
  AND U9419 ( .A(n4710), .B(p_input[5762]), .Z(o[5762]) );
  AND U9420 ( .A(p_input[25762]), .B(p_input[15762]), .Z(n4710) );
  AND U9421 ( .A(n4711), .B(p_input[5761]), .Z(o[5761]) );
  AND U9422 ( .A(p_input[25761]), .B(p_input[15761]), .Z(n4711) );
  AND U9423 ( .A(n4712), .B(p_input[5760]), .Z(o[5760]) );
  AND U9424 ( .A(p_input[25760]), .B(p_input[15760]), .Z(n4712) );
  AND U9425 ( .A(n4713), .B(p_input[575]), .Z(o[575]) );
  AND U9426 ( .A(p_input[20575]), .B(p_input[10575]), .Z(n4713) );
  AND U9427 ( .A(n4714), .B(p_input[5759]), .Z(o[5759]) );
  AND U9428 ( .A(p_input[25759]), .B(p_input[15759]), .Z(n4714) );
  AND U9429 ( .A(n4715), .B(p_input[5758]), .Z(o[5758]) );
  AND U9430 ( .A(p_input[25758]), .B(p_input[15758]), .Z(n4715) );
  AND U9431 ( .A(n4716), .B(p_input[5757]), .Z(o[5757]) );
  AND U9432 ( .A(p_input[25757]), .B(p_input[15757]), .Z(n4716) );
  AND U9433 ( .A(n4717), .B(p_input[5756]), .Z(o[5756]) );
  AND U9434 ( .A(p_input[25756]), .B(p_input[15756]), .Z(n4717) );
  AND U9435 ( .A(n4718), .B(p_input[5755]), .Z(o[5755]) );
  AND U9436 ( .A(p_input[25755]), .B(p_input[15755]), .Z(n4718) );
  AND U9437 ( .A(n4719), .B(p_input[5754]), .Z(o[5754]) );
  AND U9438 ( .A(p_input[25754]), .B(p_input[15754]), .Z(n4719) );
  AND U9439 ( .A(n4720), .B(p_input[5753]), .Z(o[5753]) );
  AND U9440 ( .A(p_input[25753]), .B(p_input[15753]), .Z(n4720) );
  AND U9441 ( .A(n4721), .B(p_input[5752]), .Z(o[5752]) );
  AND U9442 ( .A(p_input[25752]), .B(p_input[15752]), .Z(n4721) );
  AND U9443 ( .A(n4722), .B(p_input[5751]), .Z(o[5751]) );
  AND U9444 ( .A(p_input[25751]), .B(p_input[15751]), .Z(n4722) );
  AND U9445 ( .A(n4723), .B(p_input[5750]), .Z(o[5750]) );
  AND U9446 ( .A(p_input[25750]), .B(p_input[15750]), .Z(n4723) );
  AND U9447 ( .A(n4724), .B(p_input[574]), .Z(o[574]) );
  AND U9448 ( .A(p_input[20574]), .B(p_input[10574]), .Z(n4724) );
  AND U9449 ( .A(n4725), .B(p_input[5749]), .Z(o[5749]) );
  AND U9450 ( .A(p_input[25749]), .B(p_input[15749]), .Z(n4725) );
  AND U9451 ( .A(n4726), .B(p_input[5748]), .Z(o[5748]) );
  AND U9452 ( .A(p_input[25748]), .B(p_input[15748]), .Z(n4726) );
  AND U9453 ( .A(n4727), .B(p_input[5747]), .Z(o[5747]) );
  AND U9454 ( .A(p_input[25747]), .B(p_input[15747]), .Z(n4727) );
  AND U9455 ( .A(n4728), .B(p_input[5746]), .Z(o[5746]) );
  AND U9456 ( .A(p_input[25746]), .B(p_input[15746]), .Z(n4728) );
  AND U9457 ( .A(n4729), .B(p_input[5745]), .Z(o[5745]) );
  AND U9458 ( .A(p_input[25745]), .B(p_input[15745]), .Z(n4729) );
  AND U9459 ( .A(n4730), .B(p_input[5744]), .Z(o[5744]) );
  AND U9460 ( .A(p_input[25744]), .B(p_input[15744]), .Z(n4730) );
  AND U9461 ( .A(n4731), .B(p_input[5743]), .Z(o[5743]) );
  AND U9462 ( .A(p_input[25743]), .B(p_input[15743]), .Z(n4731) );
  AND U9463 ( .A(n4732), .B(p_input[5742]), .Z(o[5742]) );
  AND U9464 ( .A(p_input[25742]), .B(p_input[15742]), .Z(n4732) );
  AND U9465 ( .A(n4733), .B(p_input[5741]), .Z(o[5741]) );
  AND U9466 ( .A(p_input[25741]), .B(p_input[15741]), .Z(n4733) );
  AND U9467 ( .A(n4734), .B(p_input[5740]), .Z(o[5740]) );
  AND U9468 ( .A(p_input[25740]), .B(p_input[15740]), .Z(n4734) );
  AND U9469 ( .A(n4735), .B(p_input[573]), .Z(o[573]) );
  AND U9470 ( .A(p_input[20573]), .B(p_input[10573]), .Z(n4735) );
  AND U9471 ( .A(n4736), .B(p_input[5739]), .Z(o[5739]) );
  AND U9472 ( .A(p_input[25739]), .B(p_input[15739]), .Z(n4736) );
  AND U9473 ( .A(n4737), .B(p_input[5738]), .Z(o[5738]) );
  AND U9474 ( .A(p_input[25738]), .B(p_input[15738]), .Z(n4737) );
  AND U9475 ( .A(n4738), .B(p_input[5737]), .Z(o[5737]) );
  AND U9476 ( .A(p_input[25737]), .B(p_input[15737]), .Z(n4738) );
  AND U9477 ( .A(n4739), .B(p_input[5736]), .Z(o[5736]) );
  AND U9478 ( .A(p_input[25736]), .B(p_input[15736]), .Z(n4739) );
  AND U9479 ( .A(n4740), .B(p_input[5735]), .Z(o[5735]) );
  AND U9480 ( .A(p_input[25735]), .B(p_input[15735]), .Z(n4740) );
  AND U9481 ( .A(n4741), .B(p_input[5734]), .Z(o[5734]) );
  AND U9482 ( .A(p_input[25734]), .B(p_input[15734]), .Z(n4741) );
  AND U9483 ( .A(n4742), .B(p_input[5733]), .Z(o[5733]) );
  AND U9484 ( .A(p_input[25733]), .B(p_input[15733]), .Z(n4742) );
  AND U9485 ( .A(n4743), .B(p_input[5732]), .Z(o[5732]) );
  AND U9486 ( .A(p_input[25732]), .B(p_input[15732]), .Z(n4743) );
  AND U9487 ( .A(n4744), .B(p_input[5731]), .Z(o[5731]) );
  AND U9488 ( .A(p_input[25731]), .B(p_input[15731]), .Z(n4744) );
  AND U9489 ( .A(n4745), .B(p_input[5730]), .Z(o[5730]) );
  AND U9490 ( .A(p_input[25730]), .B(p_input[15730]), .Z(n4745) );
  AND U9491 ( .A(n4746), .B(p_input[572]), .Z(o[572]) );
  AND U9492 ( .A(p_input[20572]), .B(p_input[10572]), .Z(n4746) );
  AND U9493 ( .A(n4747), .B(p_input[5729]), .Z(o[5729]) );
  AND U9494 ( .A(p_input[25729]), .B(p_input[15729]), .Z(n4747) );
  AND U9495 ( .A(n4748), .B(p_input[5728]), .Z(o[5728]) );
  AND U9496 ( .A(p_input[25728]), .B(p_input[15728]), .Z(n4748) );
  AND U9497 ( .A(n4749), .B(p_input[5727]), .Z(o[5727]) );
  AND U9498 ( .A(p_input[25727]), .B(p_input[15727]), .Z(n4749) );
  AND U9499 ( .A(n4750), .B(p_input[5726]), .Z(o[5726]) );
  AND U9500 ( .A(p_input[25726]), .B(p_input[15726]), .Z(n4750) );
  AND U9501 ( .A(n4751), .B(p_input[5725]), .Z(o[5725]) );
  AND U9502 ( .A(p_input[25725]), .B(p_input[15725]), .Z(n4751) );
  AND U9503 ( .A(n4752), .B(p_input[5724]), .Z(o[5724]) );
  AND U9504 ( .A(p_input[25724]), .B(p_input[15724]), .Z(n4752) );
  AND U9505 ( .A(n4753), .B(p_input[5723]), .Z(o[5723]) );
  AND U9506 ( .A(p_input[25723]), .B(p_input[15723]), .Z(n4753) );
  AND U9507 ( .A(n4754), .B(p_input[5722]), .Z(o[5722]) );
  AND U9508 ( .A(p_input[25722]), .B(p_input[15722]), .Z(n4754) );
  AND U9509 ( .A(n4755), .B(p_input[5721]), .Z(o[5721]) );
  AND U9510 ( .A(p_input[25721]), .B(p_input[15721]), .Z(n4755) );
  AND U9511 ( .A(n4756), .B(p_input[5720]), .Z(o[5720]) );
  AND U9512 ( .A(p_input[25720]), .B(p_input[15720]), .Z(n4756) );
  AND U9513 ( .A(n4757), .B(p_input[571]), .Z(o[571]) );
  AND U9514 ( .A(p_input[20571]), .B(p_input[10571]), .Z(n4757) );
  AND U9515 ( .A(n4758), .B(p_input[5719]), .Z(o[5719]) );
  AND U9516 ( .A(p_input[25719]), .B(p_input[15719]), .Z(n4758) );
  AND U9517 ( .A(n4759), .B(p_input[5718]), .Z(o[5718]) );
  AND U9518 ( .A(p_input[25718]), .B(p_input[15718]), .Z(n4759) );
  AND U9519 ( .A(n4760), .B(p_input[5717]), .Z(o[5717]) );
  AND U9520 ( .A(p_input[25717]), .B(p_input[15717]), .Z(n4760) );
  AND U9521 ( .A(n4761), .B(p_input[5716]), .Z(o[5716]) );
  AND U9522 ( .A(p_input[25716]), .B(p_input[15716]), .Z(n4761) );
  AND U9523 ( .A(n4762), .B(p_input[5715]), .Z(o[5715]) );
  AND U9524 ( .A(p_input[25715]), .B(p_input[15715]), .Z(n4762) );
  AND U9525 ( .A(n4763), .B(p_input[5714]), .Z(o[5714]) );
  AND U9526 ( .A(p_input[25714]), .B(p_input[15714]), .Z(n4763) );
  AND U9527 ( .A(n4764), .B(p_input[5713]), .Z(o[5713]) );
  AND U9528 ( .A(p_input[25713]), .B(p_input[15713]), .Z(n4764) );
  AND U9529 ( .A(n4765), .B(p_input[5712]), .Z(o[5712]) );
  AND U9530 ( .A(p_input[25712]), .B(p_input[15712]), .Z(n4765) );
  AND U9531 ( .A(n4766), .B(p_input[5711]), .Z(o[5711]) );
  AND U9532 ( .A(p_input[25711]), .B(p_input[15711]), .Z(n4766) );
  AND U9533 ( .A(n4767), .B(p_input[5710]), .Z(o[5710]) );
  AND U9534 ( .A(p_input[25710]), .B(p_input[15710]), .Z(n4767) );
  AND U9535 ( .A(n4768), .B(p_input[570]), .Z(o[570]) );
  AND U9536 ( .A(p_input[20570]), .B(p_input[10570]), .Z(n4768) );
  AND U9537 ( .A(n4769), .B(p_input[5709]), .Z(o[5709]) );
  AND U9538 ( .A(p_input[25709]), .B(p_input[15709]), .Z(n4769) );
  AND U9539 ( .A(n4770), .B(p_input[5708]), .Z(o[5708]) );
  AND U9540 ( .A(p_input[25708]), .B(p_input[15708]), .Z(n4770) );
  AND U9541 ( .A(n4771), .B(p_input[5707]), .Z(o[5707]) );
  AND U9542 ( .A(p_input[25707]), .B(p_input[15707]), .Z(n4771) );
  AND U9543 ( .A(n4772), .B(p_input[5706]), .Z(o[5706]) );
  AND U9544 ( .A(p_input[25706]), .B(p_input[15706]), .Z(n4772) );
  AND U9545 ( .A(n4773), .B(p_input[5705]), .Z(o[5705]) );
  AND U9546 ( .A(p_input[25705]), .B(p_input[15705]), .Z(n4773) );
  AND U9547 ( .A(n4774), .B(p_input[5704]), .Z(o[5704]) );
  AND U9548 ( .A(p_input[25704]), .B(p_input[15704]), .Z(n4774) );
  AND U9549 ( .A(n4775), .B(p_input[5703]), .Z(o[5703]) );
  AND U9550 ( .A(p_input[25703]), .B(p_input[15703]), .Z(n4775) );
  AND U9551 ( .A(n4776), .B(p_input[5702]), .Z(o[5702]) );
  AND U9552 ( .A(p_input[25702]), .B(p_input[15702]), .Z(n4776) );
  AND U9553 ( .A(n4777), .B(p_input[5701]), .Z(o[5701]) );
  AND U9554 ( .A(p_input[25701]), .B(p_input[15701]), .Z(n4777) );
  AND U9555 ( .A(n4778), .B(p_input[5700]), .Z(o[5700]) );
  AND U9556 ( .A(p_input[25700]), .B(p_input[15700]), .Z(n4778) );
  AND U9557 ( .A(n4779), .B(p_input[56]), .Z(o[56]) );
  AND U9558 ( .A(p_input[20056]), .B(p_input[10056]), .Z(n4779) );
  AND U9559 ( .A(n4780), .B(p_input[569]), .Z(o[569]) );
  AND U9560 ( .A(p_input[20569]), .B(p_input[10569]), .Z(n4780) );
  AND U9561 ( .A(n4781), .B(p_input[5699]), .Z(o[5699]) );
  AND U9562 ( .A(p_input[25699]), .B(p_input[15699]), .Z(n4781) );
  AND U9563 ( .A(n4782), .B(p_input[5698]), .Z(o[5698]) );
  AND U9564 ( .A(p_input[25698]), .B(p_input[15698]), .Z(n4782) );
  AND U9565 ( .A(n4783), .B(p_input[5697]), .Z(o[5697]) );
  AND U9566 ( .A(p_input[25697]), .B(p_input[15697]), .Z(n4783) );
  AND U9567 ( .A(n4784), .B(p_input[5696]), .Z(o[5696]) );
  AND U9568 ( .A(p_input[25696]), .B(p_input[15696]), .Z(n4784) );
  AND U9569 ( .A(n4785), .B(p_input[5695]), .Z(o[5695]) );
  AND U9570 ( .A(p_input[25695]), .B(p_input[15695]), .Z(n4785) );
  AND U9571 ( .A(n4786), .B(p_input[5694]), .Z(o[5694]) );
  AND U9572 ( .A(p_input[25694]), .B(p_input[15694]), .Z(n4786) );
  AND U9573 ( .A(n4787), .B(p_input[5693]), .Z(o[5693]) );
  AND U9574 ( .A(p_input[25693]), .B(p_input[15693]), .Z(n4787) );
  AND U9575 ( .A(n4788), .B(p_input[5692]), .Z(o[5692]) );
  AND U9576 ( .A(p_input[25692]), .B(p_input[15692]), .Z(n4788) );
  AND U9577 ( .A(n4789), .B(p_input[5691]), .Z(o[5691]) );
  AND U9578 ( .A(p_input[25691]), .B(p_input[15691]), .Z(n4789) );
  AND U9579 ( .A(n4790), .B(p_input[5690]), .Z(o[5690]) );
  AND U9580 ( .A(p_input[25690]), .B(p_input[15690]), .Z(n4790) );
  AND U9581 ( .A(n4791), .B(p_input[568]), .Z(o[568]) );
  AND U9582 ( .A(p_input[20568]), .B(p_input[10568]), .Z(n4791) );
  AND U9583 ( .A(n4792), .B(p_input[5689]), .Z(o[5689]) );
  AND U9584 ( .A(p_input[25689]), .B(p_input[15689]), .Z(n4792) );
  AND U9585 ( .A(n4793), .B(p_input[5688]), .Z(o[5688]) );
  AND U9586 ( .A(p_input[25688]), .B(p_input[15688]), .Z(n4793) );
  AND U9587 ( .A(n4794), .B(p_input[5687]), .Z(o[5687]) );
  AND U9588 ( .A(p_input[25687]), .B(p_input[15687]), .Z(n4794) );
  AND U9589 ( .A(n4795), .B(p_input[5686]), .Z(o[5686]) );
  AND U9590 ( .A(p_input[25686]), .B(p_input[15686]), .Z(n4795) );
  AND U9591 ( .A(n4796), .B(p_input[5685]), .Z(o[5685]) );
  AND U9592 ( .A(p_input[25685]), .B(p_input[15685]), .Z(n4796) );
  AND U9593 ( .A(n4797), .B(p_input[5684]), .Z(o[5684]) );
  AND U9594 ( .A(p_input[25684]), .B(p_input[15684]), .Z(n4797) );
  AND U9595 ( .A(n4798), .B(p_input[5683]), .Z(o[5683]) );
  AND U9596 ( .A(p_input[25683]), .B(p_input[15683]), .Z(n4798) );
  AND U9597 ( .A(n4799), .B(p_input[5682]), .Z(o[5682]) );
  AND U9598 ( .A(p_input[25682]), .B(p_input[15682]), .Z(n4799) );
  AND U9599 ( .A(n4800), .B(p_input[5681]), .Z(o[5681]) );
  AND U9600 ( .A(p_input[25681]), .B(p_input[15681]), .Z(n4800) );
  AND U9601 ( .A(n4801), .B(p_input[5680]), .Z(o[5680]) );
  AND U9602 ( .A(p_input[25680]), .B(p_input[15680]), .Z(n4801) );
  AND U9603 ( .A(n4802), .B(p_input[567]), .Z(o[567]) );
  AND U9604 ( .A(p_input[20567]), .B(p_input[10567]), .Z(n4802) );
  AND U9605 ( .A(n4803), .B(p_input[5679]), .Z(o[5679]) );
  AND U9606 ( .A(p_input[25679]), .B(p_input[15679]), .Z(n4803) );
  AND U9607 ( .A(n4804), .B(p_input[5678]), .Z(o[5678]) );
  AND U9608 ( .A(p_input[25678]), .B(p_input[15678]), .Z(n4804) );
  AND U9609 ( .A(n4805), .B(p_input[5677]), .Z(o[5677]) );
  AND U9610 ( .A(p_input[25677]), .B(p_input[15677]), .Z(n4805) );
  AND U9611 ( .A(n4806), .B(p_input[5676]), .Z(o[5676]) );
  AND U9612 ( .A(p_input[25676]), .B(p_input[15676]), .Z(n4806) );
  AND U9613 ( .A(n4807), .B(p_input[5675]), .Z(o[5675]) );
  AND U9614 ( .A(p_input[25675]), .B(p_input[15675]), .Z(n4807) );
  AND U9615 ( .A(n4808), .B(p_input[5674]), .Z(o[5674]) );
  AND U9616 ( .A(p_input[25674]), .B(p_input[15674]), .Z(n4808) );
  AND U9617 ( .A(n4809), .B(p_input[5673]), .Z(o[5673]) );
  AND U9618 ( .A(p_input[25673]), .B(p_input[15673]), .Z(n4809) );
  AND U9619 ( .A(n4810), .B(p_input[5672]), .Z(o[5672]) );
  AND U9620 ( .A(p_input[25672]), .B(p_input[15672]), .Z(n4810) );
  AND U9621 ( .A(n4811), .B(p_input[5671]), .Z(o[5671]) );
  AND U9622 ( .A(p_input[25671]), .B(p_input[15671]), .Z(n4811) );
  AND U9623 ( .A(n4812), .B(p_input[5670]), .Z(o[5670]) );
  AND U9624 ( .A(p_input[25670]), .B(p_input[15670]), .Z(n4812) );
  AND U9625 ( .A(n4813), .B(p_input[566]), .Z(o[566]) );
  AND U9626 ( .A(p_input[20566]), .B(p_input[10566]), .Z(n4813) );
  AND U9627 ( .A(n4814), .B(p_input[5669]), .Z(o[5669]) );
  AND U9628 ( .A(p_input[25669]), .B(p_input[15669]), .Z(n4814) );
  AND U9629 ( .A(n4815), .B(p_input[5668]), .Z(o[5668]) );
  AND U9630 ( .A(p_input[25668]), .B(p_input[15668]), .Z(n4815) );
  AND U9631 ( .A(n4816), .B(p_input[5667]), .Z(o[5667]) );
  AND U9632 ( .A(p_input[25667]), .B(p_input[15667]), .Z(n4816) );
  AND U9633 ( .A(n4817), .B(p_input[5666]), .Z(o[5666]) );
  AND U9634 ( .A(p_input[25666]), .B(p_input[15666]), .Z(n4817) );
  AND U9635 ( .A(n4818), .B(p_input[5665]), .Z(o[5665]) );
  AND U9636 ( .A(p_input[25665]), .B(p_input[15665]), .Z(n4818) );
  AND U9637 ( .A(n4819), .B(p_input[5664]), .Z(o[5664]) );
  AND U9638 ( .A(p_input[25664]), .B(p_input[15664]), .Z(n4819) );
  AND U9639 ( .A(n4820), .B(p_input[5663]), .Z(o[5663]) );
  AND U9640 ( .A(p_input[25663]), .B(p_input[15663]), .Z(n4820) );
  AND U9641 ( .A(n4821), .B(p_input[5662]), .Z(o[5662]) );
  AND U9642 ( .A(p_input[25662]), .B(p_input[15662]), .Z(n4821) );
  AND U9643 ( .A(n4822), .B(p_input[5661]), .Z(o[5661]) );
  AND U9644 ( .A(p_input[25661]), .B(p_input[15661]), .Z(n4822) );
  AND U9645 ( .A(n4823), .B(p_input[5660]), .Z(o[5660]) );
  AND U9646 ( .A(p_input[25660]), .B(p_input[15660]), .Z(n4823) );
  AND U9647 ( .A(n4824), .B(p_input[565]), .Z(o[565]) );
  AND U9648 ( .A(p_input[20565]), .B(p_input[10565]), .Z(n4824) );
  AND U9649 ( .A(n4825), .B(p_input[5659]), .Z(o[5659]) );
  AND U9650 ( .A(p_input[25659]), .B(p_input[15659]), .Z(n4825) );
  AND U9651 ( .A(n4826), .B(p_input[5658]), .Z(o[5658]) );
  AND U9652 ( .A(p_input[25658]), .B(p_input[15658]), .Z(n4826) );
  AND U9653 ( .A(n4827), .B(p_input[5657]), .Z(o[5657]) );
  AND U9654 ( .A(p_input[25657]), .B(p_input[15657]), .Z(n4827) );
  AND U9655 ( .A(n4828), .B(p_input[5656]), .Z(o[5656]) );
  AND U9656 ( .A(p_input[25656]), .B(p_input[15656]), .Z(n4828) );
  AND U9657 ( .A(n4829), .B(p_input[5655]), .Z(o[5655]) );
  AND U9658 ( .A(p_input[25655]), .B(p_input[15655]), .Z(n4829) );
  AND U9659 ( .A(n4830), .B(p_input[5654]), .Z(o[5654]) );
  AND U9660 ( .A(p_input[25654]), .B(p_input[15654]), .Z(n4830) );
  AND U9661 ( .A(n4831), .B(p_input[5653]), .Z(o[5653]) );
  AND U9662 ( .A(p_input[25653]), .B(p_input[15653]), .Z(n4831) );
  AND U9663 ( .A(n4832), .B(p_input[5652]), .Z(o[5652]) );
  AND U9664 ( .A(p_input[25652]), .B(p_input[15652]), .Z(n4832) );
  AND U9665 ( .A(n4833), .B(p_input[5651]), .Z(o[5651]) );
  AND U9666 ( .A(p_input[25651]), .B(p_input[15651]), .Z(n4833) );
  AND U9667 ( .A(n4834), .B(p_input[5650]), .Z(o[5650]) );
  AND U9668 ( .A(p_input[25650]), .B(p_input[15650]), .Z(n4834) );
  AND U9669 ( .A(n4835), .B(p_input[564]), .Z(o[564]) );
  AND U9670 ( .A(p_input[20564]), .B(p_input[10564]), .Z(n4835) );
  AND U9671 ( .A(n4836), .B(p_input[5649]), .Z(o[5649]) );
  AND U9672 ( .A(p_input[25649]), .B(p_input[15649]), .Z(n4836) );
  AND U9673 ( .A(n4837), .B(p_input[5648]), .Z(o[5648]) );
  AND U9674 ( .A(p_input[25648]), .B(p_input[15648]), .Z(n4837) );
  AND U9675 ( .A(n4838), .B(p_input[5647]), .Z(o[5647]) );
  AND U9676 ( .A(p_input[25647]), .B(p_input[15647]), .Z(n4838) );
  AND U9677 ( .A(n4839), .B(p_input[5646]), .Z(o[5646]) );
  AND U9678 ( .A(p_input[25646]), .B(p_input[15646]), .Z(n4839) );
  AND U9679 ( .A(n4840), .B(p_input[5645]), .Z(o[5645]) );
  AND U9680 ( .A(p_input[25645]), .B(p_input[15645]), .Z(n4840) );
  AND U9681 ( .A(n4841), .B(p_input[5644]), .Z(o[5644]) );
  AND U9682 ( .A(p_input[25644]), .B(p_input[15644]), .Z(n4841) );
  AND U9683 ( .A(n4842), .B(p_input[5643]), .Z(o[5643]) );
  AND U9684 ( .A(p_input[25643]), .B(p_input[15643]), .Z(n4842) );
  AND U9685 ( .A(n4843), .B(p_input[5642]), .Z(o[5642]) );
  AND U9686 ( .A(p_input[25642]), .B(p_input[15642]), .Z(n4843) );
  AND U9687 ( .A(n4844), .B(p_input[5641]), .Z(o[5641]) );
  AND U9688 ( .A(p_input[25641]), .B(p_input[15641]), .Z(n4844) );
  AND U9689 ( .A(n4845), .B(p_input[5640]), .Z(o[5640]) );
  AND U9690 ( .A(p_input[25640]), .B(p_input[15640]), .Z(n4845) );
  AND U9691 ( .A(n4846), .B(p_input[563]), .Z(o[563]) );
  AND U9692 ( .A(p_input[20563]), .B(p_input[10563]), .Z(n4846) );
  AND U9693 ( .A(n4847), .B(p_input[5639]), .Z(o[5639]) );
  AND U9694 ( .A(p_input[25639]), .B(p_input[15639]), .Z(n4847) );
  AND U9695 ( .A(n4848), .B(p_input[5638]), .Z(o[5638]) );
  AND U9696 ( .A(p_input[25638]), .B(p_input[15638]), .Z(n4848) );
  AND U9697 ( .A(n4849), .B(p_input[5637]), .Z(o[5637]) );
  AND U9698 ( .A(p_input[25637]), .B(p_input[15637]), .Z(n4849) );
  AND U9699 ( .A(n4850), .B(p_input[5636]), .Z(o[5636]) );
  AND U9700 ( .A(p_input[25636]), .B(p_input[15636]), .Z(n4850) );
  AND U9701 ( .A(n4851), .B(p_input[5635]), .Z(o[5635]) );
  AND U9702 ( .A(p_input[25635]), .B(p_input[15635]), .Z(n4851) );
  AND U9703 ( .A(n4852), .B(p_input[5634]), .Z(o[5634]) );
  AND U9704 ( .A(p_input[25634]), .B(p_input[15634]), .Z(n4852) );
  AND U9705 ( .A(n4853), .B(p_input[5633]), .Z(o[5633]) );
  AND U9706 ( .A(p_input[25633]), .B(p_input[15633]), .Z(n4853) );
  AND U9707 ( .A(n4854), .B(p_input[5632]), .Z(o[5632]) );
  AND U9708 ( .A(p_input[25632]), .B(p_input[15632]), .Z(n4854) );
  AND U9709 ( .A(n4855), .B(p_input[5631]), .Z(o[5631]) );
  AND U9710 ( .A(p_input[25631]), .B(p_input[15631]), .Z(n4855) );
  AND U9711 ( .A(n4856), .B(p_input[5630]), .Z(o[5630]) );
  AND U9712 ( .A(p_input[25630]), .B(p_input[15630]), .Z(n4856) );
  AND U9713 ( .A(n4857), .B(p_input[562]), .Z(o[562]) );
  AND U9714 ( .A(p_input[20562]), .B(p_input[10562]), .Z(n4857) );
  AND U9715 ( .A(n4858), .B(p_input[5629]), .Z(o[5629]) );
  AND U9716 ( .A(p_input[25629]), .B(p_input[15629]), .Z(n4858) );
  AND U9717 ( .A(n4859), .B(p_input[5628]), .Z(o[5628]) );
  AND U9718 ( .A(p_input[25628]), .B(p_input[15628]), .Z(n4859) );
  AND U9719 ( .A(n4860), .B(p_input[5627]), .Z(o[5627]) );
  AND U9720 ( .A(p_input[25627]), .B(p_input[15627]), .Z(n4860) );
  AND U9721 ( .A(n4861), .B(p_input[5626]), .Z(o[5626]) );
  AND U9722 ( .A(p_input[25626]), .B(p_input[15626]), .Z(n4861) );
  AND U9723 ( .A(n4862), .B(p_input[5625]), .Z(o[5625]) );
  AND U9724 ( .A(p_input[25625]), .B(p_input[15625]), .Z(n4862) );
  AND U9725 ( .A(n4863), .B(p_input[5624]), .Z(o[5624]) );
  AND U9726 ( .A(p_input[25624]), .B(p_input[15624]), .Z(n4863) );
  AND U9727 ( .A(n4864), .B(p_input[5623]), .Z(o[5623]) );
  AND U9728 ( .A(p_input[25623]), .B(p_input[15623]), .Z(n4864) );
  AND U9729 ( .A(n4865), .B(p_input[5622]), .Z(o[5622]) );
  AND U9730 ( .A(p_input[25622]), .B(p_input[15622]), .Z(n4865) );
  AND U9731 ( .A(n4866), .B(p_input[5621]), .Z(o[5621]) );
  AND U9732 ( .A(p_input[25621]), .B(p_input[15621]), .Z(n4866) );
  AND U9733 ( .A(n4867), .B(p_input[5620]), .Z(o[5620]) );
  AND U9734 ( .A(p_input[25620]), .B(p_input[15620]), .Z(n4867) );
  AND U9735 ( .A(n4868), .B(p_input[561]), .Z(o[561]) );
  AND U9736 ( .A(p_input[20561]), .B(p_input[10561]), .Z(n4868) );
  AND U9737 ( .A(n4869), .B(p_input[5619]), .Z(o[5619]) );
  AND U9738 ( .A(p_input[25619]), .B(p_input[15619]), .Z(n4869) );
  AND U9739 ( .A(n4870), .B(p_input[5618]), .Z(o[5618]) );
  AND U9740 ( .A(p_input[25618]), .B(p_input[15618]), .Z(n4870) );
  AND U9741 ( .A(n4871), .B(p_input[5617]), .Z(o[5617]) );
  AND U9742 ( .A(p_input[25617]), .B(p_input[15617]), .Z(n4871) );
  AND U9743 ( .A(n4872), .B(p_input[5616]), .Z(o[5616]) );
  AND U9744 ( .A(p_input[25616]), .B(p_input[15616]), .Z(n4872) );
  AND U9745 ( .A(n4873), .B(p_input[5615]), .Z(o[5615]) );
  AND U9746 ( .A(p_input[25615]), .B(p_input[15615]), .Z(n4873) );
  AND U9747 ( .A(n4874), .B(p_input[5614]), .Z(o[5614]) );
  AND U9748 ( .A(p_input[25614]), .B(p_input[15614]), .Z(n4874) );
  AND U9749 ( .A(n4875), .B(p_input[5613]), .Z(o[5613]) );
  AND U9750 ( .A(p_input[25613]), .B(p_input[15613]), .Z(n4875) );
  AND U9751 ( .A(n4876), .B(p_input[5612]), .Z(o[5612]) );
  AND U9752 ( .A(p_input[25612]), .B(p_input[15612]), .Z(n4876) );
  AND U9753 ( .A(n4877), .B(p_input[5611]), .Z(o[5611]) );
  AND U9754 ( .A(p_input[25611]), .B(p_input[15611]), .Z(n4877) );
  AND U9755 ( .A(n4878), .B(p_input[5610]), .Z(o[5610]) );
  AND U9756 ( .A(p_input[25610]), .B(p_input[15610]), .Z(n4878) );
  AND U9757 ( .A(n4879), .B(p_input[560]), .Z(o[560]) );
  AND U9758 ( .A(p_input[20560]), .B(p_input[10560]), .Z(n4879) );
  AND U9759 ( .A(n4880), .B(p_input[5609]), .Z(o[5609]) );
  AND U9760 ( .A(p_input[25609]), .B(p_input[15609]), .Z(n4880) );
  AND U9761 ( .A(n4881), .B(p_input[5608]), .Z(o[5608]) );
  AND U9762 ( .A(p_input[25608]), .B(p_input[15608]), .Z(n4881) );
  AND U9763 ( .A(n4882), .B(p_input[5607]), .Z(o[5607]) );
  AND U9764 ( .A(p_input[25607]), .B(p_input[15607]), .Z(n4882) );
  AND U9765 ( .A(n4883), .B(p_input[5606]), .Z(o[5606]) );
  AND U9766 ( .A(p_input[25606]), .B(p_input[15606]), .Z(n4883) );
  AND U9767 ( .A(n4884), .B(p_input[5605]), .Z(o[5605]) );
  AND U9768 ( .A(p_input[25605]), .B(p_input[15605]), .Z(n4884) );
  AND U9769 ( .A(n4885), .B(p_input[5604]), .Z(o[5604]) );
  AND U9770 ( .A(p_input[25604]), .B(p_input[15604]), .Z(n4885) );
  AND U9771 ( .A(n4886), .B(p_input[5603]), .Z(o[5603]) );
  AND U9772 ( .A(p_input[25603]), .B(p_input[15603]), .Z(n4886) );
  AND U9773 ( .A(n4887), .B(p_input[5602]), .Z(o[5602]) );
  AND U9774 ( .A(p_input[25602]), .B(p_input[15602]), .Z(n4887) );
  AND U9775 ( .A(n4888), .B(p_input[5601]), .Z(o[5601]) );
  AND U9776 ( .A(p_input[25601]), .B(p_input[15601]), .Z(n4888) );
  AND U9777 ( .A(n4889), .B(p_input[5600]), .Z(o[5600]) );
  AND U9778 ( .A(p_input[25600]), .B(p_input[15600]), .Z(n4889) );
  AND U9779 ( .A(n4890), .B(p_input[55]), .Z(o[55]) );
  AND U9780 ( .A(p_input[20055]), .B(p_input[10055]), .Z(n4890) );
  AND U9781 ( .A(n4891), .B(p_input[559]), .Z(o[559]) );
  AND U9782 ( .A(p_input[20559]), .B(p_input[10559]), .Z(n4891) );
  AND U9783 ( .A(n4892), .B(p_input[5599]), .Z(o[5599]) );
  AND U9784 ( .A(p_input[25599]), .B(p_input[15599]), .Z(n4892) );
  AND U9785 ( .A(n4893), .B(p_input[5598]), .Z(o[5598]) );
  AND U9786 ( .A(p_input[25598]), .B(p_input[15598]), .Z(n4893) );
  AND U9787 ( .A(n4894), .B(p_input[5597]), .Z(o[5597]) );
  AND U9788 ( .A(p_input[25597]), .B(p_input[15597]), .Z(n4894) );
  AND U9789 ( .A(n4895), .B(p_input[5596]), .Z(o[5596]) );
  AND U9790 ( .A(p_input[25596]), .B(p_input[15596]), .Z(n4895) );
  AND U9791 ( .A(n4896), .B(p_input[5595]), .Z(o[5595]) );
  AND U9792 ( .A(p_input[25595]), .B(p_input[15595]), .Z(n4896) );
  AND U9793 ( .A(n4897), .B(p_input[5594]), .Z(o[5594]) );
  AND U9794 ( .A(p_input[25594]), .B(p_input[15594]), .Z(n4897) );
  AND U9795 ( .A(n4898), .B(p_input[5593]), .Z(o[5593]) );
  AND U9796 ( .A(p_input[25593]), .B(p_input[15593]), .Z(n4898) );
  AND U9797 ( .A(n4899), .B(p_input[5592]), .Z(o[5592]) );
  AND U9798 ( .A(p_input[25592]), .B(p_input[15592]), .Z(n4899) );
  AND U9799 ( .A(n4900), .B(p_input[5591]), .Z(o[5591]) );
  AND U9800 ( .A(p_input[25591]), .B(p_input[15591]), .Z(n4900) );
  AND U9801 ( .A(n4901), .B(p_input[5590]), .Z(o[5590]) );
  AND U9802 ( .A(p_input[25590]), .B(p_input[15590]), .Z(n4901) );
  AND U9803 ( .A(n4902), .B(p_input[558]), .Z(o[558]) );
  AND U9804 ( .A(p_input[20558]), .B(p_input[10558]), .Z(n4902) );
  AND U9805 ( .A(n4903), .B(p_input[5589]), .Z(o[5589]) );
  AND U9806 ( .A(p_input[25589]), .B(p_input[15589]), .Z(n4903) );
  AND U9807 ( .A(n4904), .B(p_input[5588]), .Z(o[5588]) );
  AND U9808 ( .A(p_input[25588]), .B(p_input[15588]), .Z(n4904) );
  AND U9809 ( .A(n4905), .B(p_input[5587]), .Z(o[5587]) );
  AND U9810 ( .A(p_input[25587]), .B(p_input[15587]), .Z(n4905) );
  AND U9811 ( .A(n4906), .B(p_input[5586]), .Z(o[5586]) );
  AND U9812 ( .A(p_input[25586]), .B(p_input[15586]), .Z(n4906) );
  AND U9813 ( .A(n4907), .B(p_input[5585]), .Z(o[5585]) );
  AND U9814 ( .A(p_input[25585]), .B(p_input[15585]), .Z(n4907) );
  AND U9815 ( .A(n4908), .B(p_input[5584]), .Z(o[5584]) );
  AND U9816 ( .A(p_input[25584]), .B(p_input[15584]), .Z(n4908) );
  AND U9817 ( .A(n4909), .B(p_input[5583]), .Z(o[5583]) );
  AND U9818 ( .A(p_input[25583]), .B(p_input[15583]), .Z(n4909) );
  AND U9819 ( .A(n4910), .B(p_input[5582]), .Z(o[5582]) );
  AND U9820 ( .A(p_input[25582]), .B(p_input[15582]), .Z(n4910) );
  AND U9821 ( .A(n4911), .B(p_input[5581]), .Z(o[5581]) );
  AND U9822 ( .A(p_input[25581]), .B(p_input[15581]), .Z(n4911) );
  AND U9823 ( .A(n4912), .B(p_input[5580]), .Z(o[5580]) );
  AND U9824 ( .A(p_input[25580]), .B(p_input[15580]), .Z(n4912) );
  AND U9825 ( .A(n4913), .B(p_input[557]), .Z(o[557]) );
  AND U9826 ( .A(p_input[20557]), .B(p_input[10557]), .Z(n4913) );
  AND U9827 ( .A(n4914), .B(p_input[5579]), .Z(o[5579]) );
  AND U9828 ( .A(p_input[25579]), .B(p_input[15579]), .Z(n4914) );
  AND U9829 ( .A(n4915), .B(p_input[5578]), .Z(o[5578]) );
  AND U9830 ( .A(p_input[25578]), .B(p_input[15578]), .Z(n4915) );
  AND U9831 ( .A(n4916), .B(p_input[5577]), .Z(o[5577]) );
  AND U9832 ( .A(p_input[25577]), .B(p_input[15577]), .Z(n4916) );
  AND U9833 ( .A(n4917), .B(p_input[5576]), .Z(o[5576]) );
  AND U9834 ( .A(p_input[25576]), .B(p_input[15576]), .Z(n4917) );
  AND U9835 ( .A(n4918), .B(p_input[5575]), .Z(o[5575]) );
  AND U9836 ( .A(p_input[25575]), .B(p_input[15575]), .Z(n4918) );
  AND U9837 ( .A(n4919), .B(p_input[5574]), .Z(o[5574]) );
  AND U9838 ( .A(p_input[25574]), .B(p_input[15574]), .Z(n4919) );
  AND U9839 ( .A(n4920), .B(p_input[5573]), .Z(o[5573]) );
  AND U9840 ( .A(p_input[25573]), .B(p_input[15573]), .Z(n4920) );
  AND U9841 ( .A(n4921), .B(p_input[5572]), .Z(o[5572]) );
  AND U9842 ( .A(p_input[25572]), .B(p_input[15572]), .Z(n4921) );
  AND U9843 ( .A(n4922), .B(p_input[5571]), .Z(o[5571]) );
  AND U9844 ( .A(p_input[25571]), .B(p_input[15571]), .Z(n4922) );
  AND U9845 ( .A(n4923), .B(p_input[5570]), .Z(o[5570]) );
  AND U9846 ( .A(p_input[25570]), .B(p_input[15570]), .Z(n4923) );
  AND U9847 ( .A(n4924), .B(p_input[556]), .Z(o[556]) );
  AND U9848 ( .A(p_input[20556]), .B(p_input[10556]), .Z(n4924) );
  AND U9849 ( .A(n4925), .B(p_input[5569]), .Z(o[5569]) );
  AND U9850 ( .A(p_input[25569]), .B(p_input[15569]), .Z(n4925) );
  AND U9851 ( .A(n4926), .B(p_input[5568]), .Z(o[5568]) );
  AND U9852 ( .A(p_input[25568]), .B(p_input[15568]), .Z(n4926) );
  AND U9853 ( .A(n4927), .B(p_input[5567]), .Z(o[5567]) );
  AND U9854 ( .A(p_input[25567]), .B(p_input[15567]), .Z(n4927) );
  AND U9855 ( .A(n4928), .B(p_input[5566]), .Z(o[5566]) );
  AND U9856 ( .A(p_input[25566]), .B(p_input[15566]), .Z(n4928) );
  AND U9857 ( .A(n4929), .B(p_input[5565]), .Z(o[5565]) );
  AND U9858 ( .A(p_input[25565]), .B(p_input[15565]), .Z(n4929) );
  AND U9859 ( .A(n4930), .B(p_input[5564]), .Z(o[5564]) );
  AND U9860 ( .A(p_input[25564]), .B(p_input[15564]), .Z(n4930) );
  AND U9861 ( .A(n4931), .B(p_input[5563]), .Z(o[5563]) );
  AND U9862 ( .A(p_input[25563]), .B(p_input[15563]), .Z(n4931) );
  AND U9863 ( .A(n4932), .B(p_input[5562]), .Z(o[5562]) );
  AND U9864 ( .A(p_input[25562]), .B(p_input[15562]), .Z(n4932) );
  AND U9865 ( .A(n4933), .B(p_input[5561]), .Z(o[5561]) );
  AND U9866 ( .A(p_input[25561]), .B(p_input[15561]), .Z(n4933) );
  AND U9867 ( .A(n4934), .B(p_input[5560]), .Z(o[5560]) );
  AND U9868 ( .A(p_input[25560]), .B(p_input[15560]), .Z(n4934) );
  AND U9869 ( .A(n4935), .B(p_input[555]), .Z(o[555]) );
  AND U9870 ( .A(p_input[20555]), .B(p_input[10555]), .Z(n4935) );
  AND U9871 ( .A(n4936), .B(p_input[5559]), .Z(o[5559]) );
  AND U9872 ( .A(p_input[25559]), .B(p_input[15559]), .Z(n4936) );
  AND U9873 ( .A(n4937), .B(p_input[5558]), .Z(o[5558]) );
  AND U9874 ( .A(p_input[25558]), .B(p_input[15558]), .Z(n4937) );
  AND U9875 ( .A(n4938), .B(p_input[5557]), .Z(o[5557]) );
  AND U9876 ( .A(p_input[25557]), .B(p_input[15557]), .Z(n4938) );
  AND U9877 ( .A(n4939), .B(p_input[5556]), .Z(o[5556]) );
  AND U9878 ( .A(p_input[25556]), .B(p_input[15556]), .Z(n4939) );
  AND U9879 ( .A(n4940), .B(p_input[5555]), .Z(o[5555]) );
  AND U9880 ( .A(p_input[25555]), .B(p_input[15555]), .Z(n4940) );
  AND U9881 ( .A(n4941), .B(p_input[5554]), .Z(o[5554]) );
  AND U9882 ( .A(p_input[25554]), .B(p_input[15554]), .Z(n4941) );
  AND U9883 ( .A(n4942), .B(p_input[5553]), .Z(o[5553]) );
  AND U9884 ( .A(p_input[25553]), .B(p_input[15553]), .Z(n4942) );
  AND U9885 ( .A(n4943), .B(p_input[5552]), .Z(o[5552]) );
  AND U9886 ( .A(p_input[25552]), .B(p_input[15552]), .Z(n4943) );
  AND U9887 ( .A(n4944), .B(p_input[5551]), .Z(o[5551]) );
  AND U9888 ( .A(p_input[25551]), .B(p_input[15551]), .Z(n4944) );
  AND U9889 ( .A(n4945), .B(p_input[5550]), .Z(o[5550]) );
  AND U9890 ( .A(p_input[25550]), .B(p_input[15550]), .Z(n4945) );
  AND U9891 ( .A(n4946), .B(p_input[554]), .Z(o[554]) );
  AND U9892 ( .A(p_input[20554]), .B(p_input[10554]), .Z(n4946) );
  AND U9893 ( .A(n4947), .B(p_input[5549]), .Z(o[5549]) );
  AND U9894 ( .A(p_input[25549]), .B(p_input[15549]), .Z(n4947) );
  AND U9895 ( .A(n4948), .B(p_input[5548]), .Z(o[5548]) );
  AND U9896 ( .A(p_input[25548]), .B(p_input[15548]), .Z(n4948) );
  AND U9897 ( .A(n4949), .B(p_input[5547]), .Z(o[5547]) );
  AND U9898 ( .A(p_input[25547]), .B(p_input[15547]), .Z(n4949) );
  AND U9899 ( .A(n4950), .B(p_input[5546]), .Z(o[5546]) );
  AND U9900 ( .A(p_input[25546]), .B(p_input[15546]), .Z(n4950) );
  AND U9901 ( .A(n4951), .B(p_input[5545]), .Z(o[5545]) );
  AND U9902 ( .A(p_input[25545]), .B(p_input[15545]), .Z(n4951) );
  AND U9903 ( .A(n4952), .B(p_input[5544]), .Z(o[5544]) );
  AND U9904 ( .A(p_input[25544]), .B(p_input[15544]), .Z(n4952) );
  AND U9905 ( .A(n4953), .B(p_input[5543]), .Z(o[5543]) );
  AND U9906 ( .A(p_input[25543]), .B(p_input[15543]), .Z(n4953) );
  AND U9907 ( .A(n4954), .B(p_input[5542]), .Z(o[5542]) );
  AND U9908 ( .A(p_input[25542]), .B(p_input[15542]), .Z(n4954) );
  AND U9909 ( .A(n4955), .B(p_input[5541]), .Z(o[5541]) );
  AND U9910 ( .A(p_input[25541]), .B(p_input[15541]), .Z(n4955) );
  AND U9911 ( .A(n4956), .B(p_input[5540]), .Z(o[5540]) );
  AND U9912 ( .A(p_input[25540]), .B(p_input[15540]), .Z(n4956) );
  AND U9913 ( .A(n4957), .B(p_input[553]), .Z(o[553]) );
  AND U9914 ( .A(p_input[20553]), .B(p_input[10553]), .Z(n4957) );
  AND U9915 ( .A(n4958), .B(p_input[5539]), .Z(o[5539]) );
  AND U9916 ( .A(p_input[25539]), .B(p_input[15539]), .Z(n4958) );
  AND U9917 ( .A(n4959), .B(p_input[5538]), .Z(o[5538]) );
  AND U9918 ( .A(p_input[25538]), .B(p_input[15538]), .Z(n4959) );
  AND U9919 ( .A(n4960), .B(p_input[5537]), .Z(o[5537]) );
  AND U9920 ( .A(p_input[25537]), .B(p_input[15537]), .Z(n4960) );
  AND U9921 ( .A(n4961), .B(p_input[5536]), .Z(o[5536]) );
  AND U9922 ( .A(p_input[25536]), .B(p_input[15536]), .Z(n4961) );
  AND U9923 ( .A(n4962), .B(p_input[5535]), .Z(o[5535]) );
  AND U9924 ( .A(p_input[25535]), .B(p_input[15535]), .Z(n4962) );
  AND U9925 ( .A(n4963), .B(p_input[5534]), .Z(o[5534]) );
  AND U9926 ( .A(p_input[25534]), .B(p_input[15534]), .Z(n4963) );
  AND U9927 ( .A(n4964), .B(p_input[5533]), .Z(o[5533]) );
  AND U9928 ( .A(p_input[25533]), .B(p_input[15533]), .Z(n4964) );
  AND U9929 ( .A(n4965), .B(p_input[5532]), .Z(o[5532]) );
  AND U9930 ( .A(p_input[25532]), .B(p_input[15532]), .Z(n4965) );
  AND U9931 ( .A(n4966), .B(p_input[5531]), .Z(o[5531]) );
  AND U9932 ( .A(p_input[25531]), .B(p_input[15531]), .Z(n4966) );
  AND U9933 ( .A(n4967), .B(p_input[5530]), .Z(o[5530]) );
  AND U9934 ( .A(p_input[25530]), .B(p_input[15530]), .Z(n4967) );
  AND U9935 ( .A(n4968), .B(p_input[552]), .Z(o[552]) );
  AND U9936 ( .A(p_input[20552]), .B(p_input[10552]), .Z(n4968) );
  AND U9937 ( .A(n4969), .B(p_input[5529]), .Z(o[5529]) );
  AND U9938 ( .A(p_input[25529]), .B(p_input[15529]), .Z(n4969) );
  AND U9939 ( .A(n4970), .B(p_input[5528]), .Z(o[5528]) );
  AND U9940 ( .A(p_input[25528]), .B(p_input[15528]), .Z(n4970) );
  AND U9941 ( .A(n4971), .B(p_input[5527]), .Z(o[5527]) );
  AND U9942 ( .A(p_input[25527]), .B(p_input[15527]), .Z(n4971) );
  AND U9943 ( .A(n4972), .B(p_input[5526]), .Z(o[5526]) );
  AND U9944 ( .A(p_input[25526]), .B(p_input[15526]), .Z(n4972) );
  AND U9945 ( .A(n4973), .B(p_input[5525]), .Z(o[5525]) );
  AND U9946 ( .A(p_input[25525]), .B(p_input[15525]), .Z(n4973) );
  AND U9947 ( .A(n4974), .B(p_input[5524]), .Z(o[5524]) );
  AND U9948 ( .A(p_input[25524]), .B(p_input[15524]), .Z(n4974) );
  AND U9949 ( .A(n4975), .B(p_input[5523]), .Z(o[5523]) );
  AND U9950 ( .A(p_input[25523]), .B(p_input[15523]), .Z(n4975) );
  AND U9951 ( .A(n4976), .B(p_input[5522]), .Z(o[5522]) );
  AND U9952 ( .A(p_input[25522]), .B(p_input[15522]), .Z(n4976) );
  AND U9953 ( .A(n4977), .B(p_input[5521]), .Z(o[5521]) );
  AND U9954 ( .A(p_input[25521]), .B(p_input[15521]), .Z(n4977) );
  AND U9955 ( .A(n4978), .B(p_input[5520]), .Z(o[5520]) );
  AND U9956 ( .A(p_input[25520]), .B(p_input[15520]), .Z(n4978) );
  AND U9957 ( .A(n4979), .B(p_input[551]), .Z(o[551]) );
  AND U9958 ( .A(p_input[20551]), .B(p_input[10551]), .Z(n4979) );
  AND U9959 ( .A(n4980), .B(p_input[5519]), .Z(o[5519]) );
  AND U9960 ( .A(p_input[25519]), .B(p_input[15519]), .Z(n4980) );
  AND U9961 ( .A(n4981), .B(p_input[5518]), .Z(o[5518]) );
  AND U9962 ( .A(p_input[25518]), .B(p_input[15518]), .Z(n4981) );
  AND U9963 ( .A(n4982), .B(p_input[5517]), .Z(o[5517]) );
  AND U9964 ( .A(p_input[25517]), .B(p_input[15517]), .Z(n4982) );
  AND U9965 ( .A(n4983), .B(p_input[5516]), .Z(o[5516]) );
  AND U9966 ( .A(p_input[25516]), .B(p_input[15516]), .Z(n4983) );
  AND U9967 ( .A(n4984), .B(p_input[5515]), .Z(o[5515]) );
  AND U9968 ( .A(p_input[25515]), .B(p_input[15515]), .Z(n4984) );
  AND U9969 ( .A(n4985), .B(p_input[5514]), .Z(o[5514]) );
  AND U9970 ( .A(p_input[25514]), .B(p_input[15514]), .Z(n4985) );
  AND U9971 ( .A(n4986), .B(p_input[5513]), .Z(o[5513]) );
  AND U9972 ( .A(p_input[25513]), .B(p_input[15513]), .Z(n4986) );
  AND U9973 ( .A(n4987), .B(p_input[5512]), .Z(o[5512]) );
  AND U9974 ( .A(p_input[25512]), .B(p_input[15512]), .Z(n4987) );
  AND U9975 ( .A(n4988), .B(p_input[5511]), .Z(o[5511]) );
  AND U9976 ( .A(p_input[25511]), .B(p_input[15511]), .Z(n4988) );
  AND U9977 ( .A(n4989), .B(p_input[5510]), .Z(o[5510]) );
  AND U9978 ( .A(p_input[25510]), .B(p_input[15510]), .Z(n4989) );
  AND U9979 ( .A(n4990), .B(p_input[550]), .Z(o[550]) );
  AND U9980 ( .A(p_input[20550]), .B(p_input[10550]), .Z(n4990) );
  AND U9981 ( .A(n4991), .B(p_input[5509]), .Z(o[5509]) );
  AND U9982 ( .A(p_input[25509]), .B(p_input[15509]), .Z(n4991) );
  AND U9983 ( .A(n4992), .B(p_input[5508]), .Z(o[5508]) );
  AND U9984 ( .A(p_input[25508]), .B(p_input[15508]), .Z(n4992) );
  AND U9985 ( .A(n4993), .B(p_input[5507]), .Z(o[5507]) );
  AND U9986 ( .A(p_input[25507]), .B(p_input[15507]), .Z(n4993) );
  AND U9987 ( .A(n4994), .B(p_input[5506]), .Z(o[5506]) );
  AND U9988 ( .A(p_input[25506]), .B(p_input[15506]), .Z(n4994) );
  AND U9989 ( .A(n4995), .B(p_input[5505]), .Z(o[5505]) );
  AND U9990 ( .A(p_input[25505]), .B(p_input[15505]), .Z(n4995) );
  AND U9991 ( .A(n4996), .B(p_input[5504]), .Z(o[5504]) );
  AND U9992 ( .A(p_input[25504]), .B(p_input[15504]), .Z(n4996) );
  AND U9993 ( .A(n4997), .B(p_input[5503]), .Z(o[5503]) );
  AND U9994 ( .A(p_input[25503]), .B(p_input[15503]), .Z(n4997) );
  AND U9995 ( .A(n4998), .B(p_input[5502]), .Z(o[5502]) );
  AND U9996 ( .A(p_input[25502]), .B(p_input[15502]), .Z(n4998) );
  AND U9997 ( .A(n4999), .B(p_input[5501]), .Z(o[5501]) );
  AND U9998 ( .A(p_input[25501]), .B(p_input[15501]), .Z(n4999) );
  AND U9999 ( .A(n5000), .B(p_input[5500]), .Z(o[5500]) );
  AND U10000 ( .A(p_input[25500]), .B(p_input[15500]), .Z(n5000) );
  AND U10001 ( .A(n5001), .B(p_input[54]), .Z(o[54]) );
  AND U10002 ( .A(p_input[20054]), .B(p_input[10054]), .Z(n5001) );
  AND U10003 ( .A(n5002), .B(p_input[549]), .Z(o[549]) );
  AND U10004 ( .A(p_input[20549]), .B(p_input[10549]), .Z(n5002) );
  AND U10005 ( .A(n5003), .B(p_input[5499]), .Z(o[5499]) );
  AND U10006 ( .A(p_input[25499]), .B(p_input[15499]), .Z(n5003) );
  AND U10007 ( .A(n5004), .B(p_input[5498]), .Z(o[5498]) );
  AND U10008 ( .A(p_input[25498]), .B(p_input[15498]), .Z(n5004) );
  AND U10009 ( .A(n5005), .B(p_input[5497]), .Z(o[5497]) );
  AND U10010 ( .A(p_input[25497]), .B(p_input[15497]), .Z(n5005) );
  AND U10011 ( .A(n5006), .B(p_input[5496]), .Z(o[5496]) );
  AND U10012 ( .A(p_input[25496]), .B(p_input[15496]), .Z(n5006) );
  AND U10013 ( .A(n5007), .B(p_input[5495]), .Z(o[5495]) );
  AND U10014 ( .A(p_input[25495]), .B(p_input[15495]), .Z(n5007) );
  AND U10015 ( .A(n5008), .B(p_input[5494]), .Z(o[5494]) );
  AND U10016 ( .A(p_input[25494]), .B(p_input[15494]), .Z(n5008) );
  AND U10017 ( .A(n5009), .B(p_input[5493]), .Z(o[5493]) );
  AND U10018 ( .A(p_input[25493]), .B(p_input[15493]), .Z(n5009) );
  AND U10019 ( .A(n5010), .B(p_input[5492]), .Z(o[5492]) );
  AND U10020 ( .A(p_input[25492]), .B(p_input[15492]), .Z(n5010) );
  AND U10021 ( .A(n5011), .B(p_input[5491]), .Z(o[5491]) );
  AND U10022 ( .A(p_input[25491]), .B(p_input[15491]), .Z(n5011) );
  AND U10023 ( .A(n5012), .B(p_input[5490]), .Z(o[5490]) );
  AND U10024 ( .A(p_input[25490]), .B(p_input[15490]), .Z(n5012) );
  AND U10025 ( .A(n5013), .B(p_input[548]), .Z(o[548]) );
  AND U10026 ( .A(p_input[20548]), .B(p_input[10548]), .Z(n5013) );
  AND U10027 ( .A(n5014), .B(p_input[5489]), .Z(o[5489]) );
  AND U10028 ( .A(p_input[25489]), .B(p_input[15489]), .Z(n5014) );
  AND U10029 ( .A(n5015), .B(p_input[5488]), .Z(o[5488]) );
  AND U10030 ( .A(p_input[25488]), .B(p_input[15488]), .Z(n5015) );
  AND U10031 ( .A(n5016), .B(p_input[5487]), .Z(o[5487]) );
  AND U10032 ( .A(p_input[25487]), .B(p_input[15487]), .Z(n5016) );
  AND U10033 ( .A(n5017), .B(p_input[5486]), .Z(o[5486]) );
  AND U10034 ( .A(p_input[25486]), .B(p_input[15486]), .Z(n5017) );
  AND U10035 ( .A(n5018), .B(p_input[5485]), .Z(o[5485]) );
  AND U10036 ( .A(p_input[25485]), .B(p_input[15485]), .Z(n5018) );
  AND U10037 ( .A(n5019), .B(p_input[5484]), .Z(o[5484]) );
  AND U10038 ( .A(p_input[25484]), .B(p_input[15484]), .Z(n5019) );
  AND U10039 ( .A(n5020), .B(p_input[5483]), .Z(o[5483]) );
  AND U10040 ( .A(p_input[25483]), .B(p_input[15483]), .Z(n5020) );
  AND U10041 ( .A(n5021), .B(p_input[5482]), .Z(o[5482]) );
  AND U10042 ( .A(p_input[25482]), .B(p_input[15482]), .Z(n5021) );
  AND U10043 ( .A(n5022), .B(p_input[5481]), .Z(o[5481]) );
  AND U10044 ( .A(p_input[25481]), .B(p_input[15481]), .Z(n5022) );
  AND U10045 ( .A(n5023), .B(p_input[5480]), .Z(o[5480]) );
  AND U10046 ( .A(p_input[25480]), .B(p_input[15480]), .Z(n5023) );
  AND U10047 ( .A(n5024), .B(p_input[547]), .Z(o[547]) );
  AND U10048 ( .A(p_input[20547]), .B(p_input[10547]), .Z(n5024) );
  AND U10049 ( .A(n5025), .B(p_input[5479]), .Z(o[5479]) );
  AND U10050 ( .A(p_input[25479]), .B(p_input[15479]), .Z(n5025) );
  AND U10051 ( .A(n5026), .B(p_input[5478]), .Z(o[5478]) );
  AND U10052 ( .A(p_input[25478]), .B(p_input[15478]), .Z(n5026) );
  AND U10053 ( .A(n5027), .B(p_input[5477]), .Z(o[5477]) );
  AND U10054 ( .A(p_input[25477]), .B(p_input[15477]), .Z(n5027) );
  AND U10055 ( .A(n5028), .B(p_input[5476]), .Z(o[5476]) );
  AND U10056 ( .A(p_input[25476]), .B(p_input[15476]), .Z(n5028) );
  AND U10057 ( .A(n5029), .B(p_input[5475]), .Z(o[5475]) );
  AND U10058 ( .A(p_input[25475]), .B(p_input[15475]), .Z(n5029) );
  AND U10059 ( .A(n5030), .B(p_input[5474]), .Z(o[5474]) );
  AND U10060 ( .A(p_input[25474]), .B(p_input[15474]), .Z(n5030) );
  AND U10061 ( .A(n5031), .B(p_input[5473]), .Z(o[5473]) );
  AND U10062 ( .A(p_input[25473]), .B(p_input[15473]), .Z(n5031) );
  AND U10063 ( .A(n5032), .B(p_input[5472]), .Z(o[5472]) );
  AND U10064 ( .A(p_input[25472]), .B(p_input[15472]), .Z(n5032) );
  AND U10065 ( .A(n5033), .B(p_input[5471]), .Z(o[5471]) );
  AND U10066 ( .A(p_input[25471]), .B(p_input[15471]), .Z(n5033) );
  AND U10067 ( .A(n5034), .B(p_input[5470]), .Z(o[5470]) );
  AND U10068 ( .A(p_input[25470]), .B(p_input[15470]), .Z(n5034) );
  AND U10069 ( .A(n5035), .B(p_input[546]), .Z(o[546]) );
  AND U10070 ( .A(p_input[20546]), .B(p_input[10546]), .Z(n5035) );
  AND U10071 ( .A(n5036), .B(p_input[5469]), .Z(o[5469]) );
  AND U10072 ( .A(p_input[25469]), .B(p_input[15469]), .Z(n5036) );
  AND U10073 ( .A(n5037), .B(p_input[5468]), .Z(o[5468]) );
  AND U10074 ( .A(p_input[25468]), .B(p_input[15468]), .Z(n5037) );
  AND U10075 ( .A(n5038), .B(p_input[5467]), .Z(o[5467]) );
  AND U10076 ( .A(p_input[25467]), .B(p_input[15467]), .Z(n5038) );
  AND U10077 ( .A(n5039), .B(p_input[5466]), .Z(o[5466]) );
  AND U10078 ( .A(p_input[25466]), .B(p_input[15466]), .Z(n5039) );
  AND U10079 ( .A(n5040), .B(p_input[5465]), .Z(o[5465]) );
  AND U10080 ( .A(p_input[25465]), .B(p_input[15465]), .Z(n5040) );
  AND U10081 ( .A(n5041), .B(p_input[5464]), .Z(o[5464]) );
  AND U10082 ( .A(p_input[25464]), .B(p_input[15464]), .Z(n5041) );
  AND U10083 ( .A(n5042), .B(p_input[5463]), .Z(o[5463]) );
  AND U10084 ( .A(p_input[25463]), .B(p_input[15463]), .Z(n5042) );
  AND U10085 ( .A(n5043), .B(p_input[5462]), .Z(o[5462]) );
  AND U10086 ( .A(p_input[25462]), .B(p_input[15462]), .Z(n5043) );
  AND U10087 ( .A(n5044), .B(p_input[5461]), .Z(o[5461]) );
  AND U10088 ( .A(p_input[25461]), .B(p_input[15461]), .Z(n5044) );
  AND U10089 ( .A(n5045), .B(p_input[5460]), .Z(o[5460]) );
  AND U10090 ( .A(p_input[25460]), .B(p_input[15460]), .Z(n5045) );
  AND U10091 ( .A(n5046), .B(p_input[545]), .Z(o[545]) );
  AND U10092 ( .A(p_input[20545]), .B(p_input[10545]), .Z(n5046) );
  AND U10093 ( .A(n5047), .B(p_input[5459]), .Z(o[5459]) );
  AND U10094 ( .A(p_input[25459]), .B(p_input[15459]), .Z(n5047) );
  AND U10095 ( .A(n5048), .B(p_input[5458]), .Z(o[5458]) );
  AND U10096 ( .A(p_input[25458]), .B(p_input[15458]), .Z(n5048) );
  AND U10097 ( .A(n5049), .B(p_input[5457]), .Z(o[5457]) );
  AND U10098 ( .A(p_input[25457]), .B(p_input[15457]), .Z(n5049) );
  AND U10099 ( .A(n5050), .B(p_input[5456]), .Z(o[5456]) );
  AND U10100 ( .A(p_input[25456]), .B(p_input[15456]), .Z(n5050) );
  AND U10101 ( .A(n5051), .B(p_input[5455]), .Z(o[5455]) );
  AND U10102 ( .A(p_input[25455]), .B(p_input[15455]), .Z(n5051) );
  AND U10103 ( .A(n5052), .B(p_input[5454]), .Z(o[5454]) );
  AND U10104 ( .A(p_input[25454]), .B(p_input[15454]), .Z(n5052) );
  AND U10105 ( .A(n5053), .B(p_input[5453]), .Z(o[5453]) );
  AND U10106 ( .A(p_input[25453]), .B(p_input[15453]), .Z(n5053) );
  AND U10107 ( .A(n5054), .B(p_input[5452]), .Z(o[5452]) );
  AND U10108 ( .A(p_input[25452]), .B(p_input[15452]), .Z(n5054) );
  AND U10109 ( .A(n5055), .B(p_input[5451]), .Z(o[5451]) );
  AND U10110 ( .A(p_input[25451]), .B(p_input[15451]), .Z(n5055) );
  AND U10111 ( .A(n5056), .B(p_input[5450]), .Z(o[5450]) );
  AND U10112 ( .A(p_input[25450]), .B(p_input[15450]), .Z(n5056) );
  AND U10113 ( .A(n5057), .B(p_input[544]), .Z(o[544]) );
  AND U10114 ( .A(p_input[20544]), .B(p_input[10544]), .Z(n5057) );
  AND U10115 ( .A(n5058), .B(p_input[5449]), .Z(o[5449]) );
  AND U10116 ( .A(p_input[25449]), .B(p_input[15449]), .Z(n5058) );
  AND U10117 ( .A(n5059), .B(p_input[5448]), .Z(o[5448]) );
  AND U10118 ( .A(p_input[25448]), .B(p_input[15448]), .Z(n5059) );
  AND U10119 ( .A(n5060), .B(p_input[5447]), .Z(o[5447]) );
  AND U10120 ( .A(p_input[25447]), .B(p_input[15447]), .Z(n5060) );
  AND U10121 ( .A(n5061), .B(p_input[5446]), .Z(o[5446]) );
  AND U10122 ( .A(p_input[25446]), .B(p_input[15446]), .Z(n5061) );
  AND U10123 ( .A(n5062), .B(p_input[5445]), .Z(o[5445]) );
  AND U10124 ( .A(p_input[25445]), .B(p_input[15445]), .Z(n5062) );
  AND U10125 ( .A(n5063), .B(p_input[5444]), .Z(o[5444]) );
  AND U10126 ( .A(p_input[25444]), .B(p_input[15444]), .Z(n5063) );
  AND U10127 ( .A(n5064), .B(p_input[5443]), .Z(o[5443]) );
  AND U10128 ( .A(p_input[25443]), .B(p_input[15443]), .Z(n5064) );
  AND U10129 ( .A(n5065), .B(p_input[5442]), .Z(o[5442]) );
  AND U10130 ( .A(p_input[25442]), .B(p_input[15442]), .Z(n5065) );
  AND U10131 ( .A(n5066), .B(p_input[5441]), .Z(o[5441]) );
  AND U10132 ( .A(p_input[25441]), .B(p_input[15441]), .Z(n5066) );
  AND U10133 ( .A(n5067), .B(p_input[5440]), .Z(o[5440]) );
  AND U10134 ( .A(p_input[25440]), .B(p_input[15440]), .Z(n5067) );
  AND U10135 ( .A(n5068), .B(p_input[543]), .Z(o[543]) );
  AND U10136 ( .A(p_input[20543]), .B(p_input[10543]), .Z(n5068) );
  AND U10137 ( .A(n5069), .B(p_input[5439]), .Z(o[5439]) );
  AND U10138 ( .A(p_input[25439]), .B(p_input[15439]), .Z(n5069) );
  AND U10139 ( .A(n5070), .B(p_input[5438]), .Z(o[5438]) );
  AND U10140 ( .A(p_input[25438]), .B(p_input[15438]), .Z(n5070) );
  AND U10141 ( .A(n5071), .B(p_input[5437]), .Z(o[5437]) );
  AND U10142 ( .A(p_input[25437]), .B(p_input[15437]), .Z(n5071) );
  AND U10143 ( .A(n5072), .B(p_input[5436]), .Z(o[5436]) );
  AND U10144 ( .A(p_input[25436]), .B(p_input[15436]), .Z(n5072) );
  AND U10145 ( .A(n5073), .B(p_input[5435]), .Z(o[5435]) );
  AND U10146 ( .A(p_input[25435]), .B(p_input[15435]), .Z(n5073) );
  AND U10147 ( .A(n5074), .B(p_input[5434]), .Z(o[5434]) );
  AND U10148 ( .A(p_input[25434]), .B(p_input[15434]), .Z(n5074) );
  AND U10149 ( .A(n5075), .B(p_input[5433]), .Z(o[5433]) );
  AND U10150 ( .A(p_input[25433]), .B(p_input[15433]), .Z(n5075) );
  AND U10151 ( .A(n5076), .B(p_input[5432]), .Z(o[5432]) );
  AND U10152 ( .A(p_input[25432]), .B(p_input[15432]), .Z(n5076) );
  AND U10153 ( .A(n5077), .B(p_input[5431]), .Z(o[5431]) );
  AND U10154 ( .A(p_input[25431]), .B(p_input[15431]), .Z(n5077) );
  AND U10155 ( .A(n5078), .B(p_input[5430]), .Z(o[5430]) );
  AND U10156 ( .A(p_input[25430]), .B(p_input[15430]), .Z(n5078) );
  AND U10157 ( .A(n5079), .B(p_input[542]), .Z(o[542]) );
  AND U10158 ( .A(p_input[20542]), .B(p_input[10542]), .Z(n5079) );
  AND U10159 ( .A(n5080), .B(p_input[5429]), .Z(o[5429]) );
  AND U10160 ( .A(p_input[25429]), .B(p_input[15429]), .Z(n5080) );
  AND U10161 ( .A(n5081), .B(p_input[5428]), .Z(o[5428]) );
  AND U10162 ( .A(p_input[25428]), .B(p_input[15428]), .Z(n5081) );
  AND U10163 ( .A(n5082), .B(p_input[5427]), .Z(o[5427]) );
  AND U10164 ( .A(p_input[25427]), .B(p_input[15427]), .Z(n5082) );
  AND U10165 ( .A(n5083), .B(p_input[5426]), .Z(o[5426]) );
  AND U10166 ( .A(p_input[25426]), .B(p_input[15426]), .Z(n5083) );
  AND U10167 ( .A(n5084), .B(p_input[5425]), .Z(o[5425]) );
  AND U10168 ( .A(p_input[25425]), .B(p_input[15425]), .Z(n5084) );
  AND U10169 ( .A(n5085), .B(p_input[5424]), .Z(o[5424]) );
  AND U10170 ( .A(p_input[25424]), .B(p_input[15424]), .Z(n5085) );
  AND U10171 ( .A(n5086), .B(p_input[5423]), .Z(o[5423]) );
  AND U10172 ( .A(p_input[25423]), .B(p_input[15423]), .Z(n5086) );
  AND U10173 ( .A(n5087), .B(p_input[5422]), .Z(o[5422]) );
  AND U10174 ( .A(p_input[25422]), .B(p_input[15422]), .Z(n5087) );
  AND U10175 ( .A(n5088), .B(p_input[5421]), .Z(o[5421]) );
  AND U10176 ( .A(p_input[25421]), .B(p_input[15421]), .Z(n5088) );
  AND U10177 ( .A(n5089), .B(p_input[5420]), .Z(o[5420]) );
  AND U10178 ( .A(p_input[25420]), .B(p_input[15420]), .Z(n5089) );
  AND U10179 ( .A(n5090), .B(p_input[541]), .Z(o[541]) );
  AND U10180 ( .A(p_input[20541]), .B(p_input[10541]), .Z(n5090) );
  AND U10181 ( .A(n5091), .B(p_input[5419]), .Z(o[5419]) );
  AND U10182 ( .A(p_input[25419]), .B(p_input[15419]), .Z(n5091) );
  AND U10183 ( .A(n5092), .B(p_input[5418]), .Z(o[5418]) );
  AND U10184 ( .A(p_input[25418]), .B(p_input[15418]), .Z(n5092) );
  AND U10185 ( .A(n5093), .B(p_input[5417]), .Z(o[5417]) );
  AND U10186 ( .A(p_input[25417]), .B(p_input[15417]), .Z(n5093) );
  AND U10187 ( .A(n5094), .B(p_input[5416]), .Z(o[5416]) );
  AND U10188 ( .A(p_input[25416]), .B(p_input[15416]), .Z(n5094) );
  AND U10189 ( .A(n5095), .B(p_input[5415]), .Z(o[5415]) );
  AND U10190 ( .A(p_input[25415]), .B(p_input[15415]), .Z(n5095) );
  AND U10191 ( .A(n5096), .B(p_input[5414]), .Z(o[5414]) );
  AND U10192 ( .A(p_input[25414]), .B(p_input[15414]), .Z(n5096) );
  AND U10193 ( .A(n5097), .B(p_input[5413]), .Z(o[5413]) );
  AND U10194 ( .A(p_input[25413]), .B(p_input[15413]), .Z(n5097) );
  AND U10195 ( .A(n5098), .B(p_input[5412]), .Z(o[5412]) );
  AND U10196 ( .A(p_input[25412]), .B(p_input[15412]), .Z(n5098) );
  AND U10197 ( .A(n5099), .B(p_input[5411]), .Z(o[5411]) );
  AND U10198 ( .A(p_input[25411]), .B(p_input[15411]), .Z(n5099) );
  AND U10199 ( .A(n5100), .B(p_input[5410]), .Z(o[5410]) );
  AND U10200 ( .A(p_input[25410]), .B(p_input[15410]), .Z(n5100) );
  AND U10201 ( .A(n5101), .B(p_input[540]), .Z(o[540]) );
  AND U10202 ( .A(p_input[20540]), .B(p_input[10540]), .Z(n5101) );
  AND U10203 ( .A(n5102), .B(p_input[5409]), .Z(o[5409]) );
  AND U10204 ( .A(p_input[25409]), .B(p_input[15409]), .Z(n5102) );
  AND U10205 ( .A(n5103), .B(p_input[5408]), .Z(o[5408]) );
  AND U10206 ( .A(p_input[25408]), .B(p_input[15408]), .Z(n5103) );
  AND U10207 ( .A(n5104), .B(p_input[5407]), .Z(o[5407]) );
  AND U10208 ( .A(p_input[25407]), .B(p_input[15407]), .Z(n5104) );
  AND U10209 ( .A(n5105), .B(p_input[5406]), .Z(o[5406]) );
  AND U10210 ( .A(p_input[25406]), .B(p_input[15406]), .Z(n5105) );
  AND U10211 ( .A(n5106), .B(p_input[5405]), .Z(o[5405]) );
  AND U10212 ( .A(p_input[25405]), .B(p_input[15405]), .Z(n5106) );
  AND U10213 ( .A(n5107), .B(p_input[5404]), .Z(o[5404]) );
  AND U10214 ( .A(p_input[25404]), .B(p_input[15404]), .Z(n5107) );
  AND U10215 ( .A(n5108), .B(p_input[5403]), .Z(o[5403]) );
  AND U10216 ( .A(p_input[25403]), .B(p_input[15403]), .Z(n5108) );
  AND U10217 ( .A(n5109), .B(p_input[5402]), .Z(o[5402]) );
  AND U10218 ( .A(p_input[25402]), .B(p_input[15402]), .Z(n5109) );
  AND U10219 ( .A(n5110), .B(p_input[5401]), .Z(o[5401]) );
  AND U10220 ( .A(p_input[25401]), .B(p_input[15401]), .Z(n5110) );
  AND U10221 ( .A(n5111), .B(p_input[5400]), .Z(o[5400]) );
  AND U10222 ( .A(p_input[25400]), .B(p_input[15400]), .Z(n5111) );
  AND U10223 ( .A(n5112), .B(p_input[53]), .Z(o[53]) );
  AND U10224 ( .A(p_input[20053]), .B(p_input[10053]), .Z(n5112) );
  AND U10225 ( .A(n5113), .B(p_input[539]), .Z(o[539]) );
  AND U10226 ( .A(p_input[20539]), .B(p_input[10539]), .Z(n5113) );
  AND U10227 ( .A(n5114), .B(p_input[5399]), .Z(o[5399]) );
  AND U10228 ( .A(p_input[25399]), .B(p_input[15399]), .Z(n5114) );
  AND U10229 ( .A(n5115), .B(p_input[5398]), .Z(o[5398]) );
  AND U10230 ( .A(p_input[25398]), .B(p_input[15398]), .Z(n5115) );
  AND U10231 ( .A(n5116), .B(p_input[5397]), .Z(o[5397]) );
  AND U10232 ( .A(p_input[25397]), .B(p_input[15397]), .Z(n5116) );
  AND U10233 ( .A(n5117), .B(p_input[5396]), .Z(o[5396]) );
  AND U10234 ( .A(p_input[25396]), .B(p_input[15396]), .Z(n5117) );
  AND U10235 ( .A(n5118), .B(p_input[5395]), .Z(o[5395]) );
  AND U10236 ( .A(p_input[25395]), .B(p_input[15395]), .Z(n5118) );
  AND U10237 ( .A(n5119), .B(p_input[5394]), .Z(o[5394]) );
  AND U10238 ( .A(p_input[25394]), .B(p_input[15394]), .Z(n5119) );
  AND U10239 ( .A(n5120), .B(p_input[5393]), .Z(o[5393]) );
  AND U10240 ( .A(p_input[25393]), .B(p_input[15393]), .Z(n5120) );
  AND U10241 ( .A(n5121), .B(p_input[5392]), .Z(o[5392]) );
  AND U10242 ( .A(p_input[25392]), .B(p_input[15392]), .Z(n5121) );
  AND U10243 ( .A(n5122), .B(p_input[5391]), .Z(o[5391]) );
  AND U10244 ( .A(p_input[25391]), .B(p_input[15391]), .Z(n5122) );
  AND U10245 ( .A(n5123), .B(p_input[5390]), .Z(o[5390]) );
  AND U10246 ( .A(p_input[25390]), .B(p_input[15390]), .Z(n5123) );
  AND U10247 ( .A(n5124), .B(p_input[538]), .Z(o[538]) );
  AND U10248 ( .A(p_input[20538]), .B(p_input[10538]), .Z(n5124) );
  AND U10249 ( .A(n5125), .B(p_input[5389]), .Z(o[5389]) );
  AND U10250 ( .A(p_input[25389]), .B(p_input[15389]), .Z(n5125) );
  AND U10251 ( .A(n5126), .B(p_input[5388]), .Z(o[5388]) );
  AND U10252 ( .A(p_input[25388]), .B(p_input[15388]), .Z(n5126) );
  AND U10253 ( .A(n5127), .B(p_input[5387]), .Z(o[5387]) );
  AND U10254 ( .A(p_input[25387]), .B(p_input[15387]), .Z(n5127) );
  AND U10255 ( .A(n5128), .B(p_input[5386]), .Z(o[5386]) );
  AND U10256 ( .A(p_input[25386]), .B(p_input[15386]), .Z(n5128) );
  AND U10257 ( .A(n5129), .B(p_input[5385]), .Z(o[5385]) );
  AND U10258 ( .A(p_input[25385]), .B(p_input[15385]), .Z(n5129) );
  AND U10259 ( .A(n5130), .B(p_input[5384]), .Z(o[5384]) );
  AND U10260 ( .A(p_input[25384]), .B(p_input[15384]), .Z(n5130) );
  AND U10261 ( .A(n5131), .B(p_input[5383]), .Z(o[5383]) );
  AND U10262 ( .A(p_input[25383]), .B(p_input[15383]), .Z(n5131) );
  AND U10263 ( .A(n5132), .B(p_input[5382]), .Z(o[5382]) );
  AND U10264 ( .A(p_input[25382]), .B(p_input[15382]), .Z(n5132) );
  AND U10265 ( .A(n5133), .B(p_input[5381]), .Z(o[5381]) );
  AND U10266 ( .A(p_input[25381]), .B(p_input[15381]), .Z(n5133) );
  AND U10267 ( .A(n5134), .B(p_input[5380]), .Z(o[5380]) );
  AND U10268 ( .A(p_input[25380]), .B(p_input[15380]), .Z(n5134) );
  AND U10269 ( .A(n5135), .B(p_input[537]), .Z(o[537]) );
  AND U10270 ( .A(p_input[20537]), .B(p_input[10537]), .Z(n5135) );
  AND U10271 ( .A(n5136), .B(p_input[5379]), .Z(o[5379]) );
  AND U10272 ( .A(p_input[25379]), .B(p_input[15379]), .Z(n5136) );
  AND U10273 ( .A(n5137), .B(p_input[5378]), .Z(o[5378]) );
  AND U10274 ( .A(p_input[25378]), .B(p_input[15378]), .Z(n5137) );
  AND U10275 ( .A(n5138), .B(p_input[5377]), .Z(o[5377]) );
  AND U10276 ( .A(p_input[25377]), .B(p_input[15377]), .Z(n5138) );
  AND U10277 ( .A(n5139), .B(p_input[5376]), .Z(o[5376]) );
  AND U10278 ( .A(p_input[25376]), .B(p_input[15376]), .Z(n5139) );
  AND U10279 ( .A(n5140), .B(p_input[5375]), .Z(o[5375]) );
  AND U10280 ( .A(p_input[25375]), .B(p_input[15375]), .Z(n5140) );
  AND U10281 ( .A(n5141), .B(p_input[5374]), .Z(o[5374]) );
  AND U10282 ( .A(p_input[25374]), .B(p_input[15374]), .Z(n5141) );
  AND U10283 ( .A(n5142), .B(p_input[5373]), .Z(o[5373]) );
  AND U10284 ( .A(p_input[25373]), .B(p_input[15373]), .Z(n5142) );
  AND U10285 ( .A(n5143), .B(p_input[5372]), .Z(o[5372]) );
  AND U10286 ( .A(p_input[25372]), .B(p_input[15372]), .Z(n5143) );
  AND U10287 ( .A(n5144), .B(p_input[5371]), .Z(o[5371]) );
  AND U10288 ( .A(p_input[25371]), .B(p_input[15371]), .Z(n5144) );
  AND U10289 ( .A(n5145), .B(p_input[5370]), .Z(o[5370]) );
  AND U10290 ( .A(p_input[25370]), .B(p_input[15370]), .Z(n5145) );
  AND U10291 ( .A(n5146), .B(p_input[536]), .Z(o[536]) );
  AND U10292 ( .A(p_input[20536]), .B(p_input[10536]), .Z(n5146) );
  AND U10293 ( .A(n5147), .B(p_input[5369]), .Z(o[5369]) );
  AND U10294 ( .A(p_input[25369]), .B(p_input[15369]), .Z(n5147) );
  AND U10295 ( .A(n5148), .B(p_input[5368]), .Z(o[5368]) );
  AND U10296 ( .A(p_input[25368]), .B(p_input[15368]), .Z(n5148) );
  AND U10297 ( .A(n5149), .B(p_input[5367]), .Z(o[5367]) );
  AND U10298 ( .A(p_input[25367]), .B(p_input[15367]), .Z(n5149) );
  AND U10299 ( .A(n5150), .B(p_input[5366]), .Z(o[5366]) );
  AND U10300 ( .A(p_input[25366]), .B(p_input[15366]), .Z(n5150) );
  AND U10301 ( .A(n5151), .B(p_input[5365]), .Z(o[5365]) );
  AND U10302 ( .A(p_input[25365]), .B(p_input[15365]), .Z(n5151) );
  AND U10303 ( .A(n5152), .B(p_input[5364]), .Z(o[5364]) );
  AND U10304 ( .A(p_input[25364]), .B(p_input[15364]), .Z(n5152) );
  AND U10305 ( .A(n5153), .B(p_input[5363]), .Z(o[5363]) );
  AND U10306 ( .A(p_input[25363]), .B(p_input[15363]), .Z(n5153) );
  AND U10307 ( .A(n5154), .B(p_input[5362]), .Z(o[5362]) );
  AND U10308 ( .A(p_input[25362]), .B(p_input[15362]), .Z(n5154) );
  AND U10309 ( .A(n5155), .B(p_input[5361]), .Z(o[5361]) );
  AND U10310 ( .A(p_input[25361]), .B(p_input[15361]), .Z(n5155) );
  AND U10311 ( .A(n5156), .B(p_input[5360]), .Z(o[5360]) );
  AND U10312 ( .A(p_input[25360]), .B(p_input[15360]), .Z(n5156) );
  AND U10313 ( .A(n5157), .B(p_input[535]), .Z(o[535]) );
  AND U10314 ( .A(p_input[20535]), .B(p_input[10535]), .Z(n5157) );
  AND U10315 ( .A(n5158), .B(p_input[5359]), .Z(o[5359]) );
  AND U10316 ( .A(p_input[25359]), .B(p_input[15359]), .Z(n5158) );
  AND U10317 ( .A(n5159), .B(p_input[5358]), .Z(o[5358]) );
  AND U10318 ( .A(p_input[25358]), .B(p_input[15358]), .Z(n5159) );
  AND U10319 ( .A(n5160), .B(p_input[5357]), .Z(o[5357]) );
  AND U10320 ( .A(p_input[25357]), .B(p_input[15357]), .Z(n5160) );
  AND U10321 ( .A(n5161), .B(p_input[5356]), .Z(o[5356]) );
  AND U10322 ( .A(p_input[25356]), .B(p_input[15356]), .Z(n5161) );
  AND U10323 ( .A(n5162), .B(p_input[5355]), .Z(o[5355]) );
  AND U10324 ( .A(p_input[25355]), .B(p_input[15355]), .Z(n5162) );
  AND U10325 ( .A(n5163), .B(p_input[5354]), .Z(o[5354]) );
  AND U10326 ( .A(p_input[25354]), .B(p_input[15354]), .Z(n5163) );
  AND U10327 ( .A(n5164), .B(p_input[5353]), .Z(o[5353]) );
  AND U10328 ( .A(p_input[25353]), .B(p_input[15353]), .Z(n5164) );
  AND U10329 ( .A(n5165), .B(p_input[5352]), .Z(o[5352]) );
  AND U10330 ( .A(p_input[25352]), .B(p_input[15352]), .Z(n5165) );
  AND U10331 ( .A(n5166), .B(p_input[5351]), .Z(o[5351]) );
  AND U10332 ( .A(p_input[25351]), .B(p_input[15351]), .Z(n5166) );
  AND U10333 ( .A(n5167), .B(p_input[5350]), .Z(o[5350]) );
  AND U10334 ( .A(p_input[25350]), .B(p_input[15350]), .Z(n5167) );
  AND U10335 ( .A(n5168), .B(p_input[534]), .Z(o[534]) );
  AND U10336 ( .A(p_input[20534]), .B(p_input[10534]), .Z(n5168) );
  AND U10337 ( .A(n5169), .B(p_input[5349]), .Z(o[5349]) );
  AND U10338 ( .A(p_input[25349]), .B(p_input[15349]), .Z(n5169) );
  AND U10339 ( .A(n5170), .B(p_input[5348]), .Z(o[5348]) );
  AND U10340 ( .A(p_input[25348]), .B(p_input[15348]), .Z(n5170) );
  AND U10341 ( .A(n5171), .B(p_input[5347]), .Z(o[5347]) );
  AND U10342 ( .A(p_input[25347]), .B(p_input[15347]), .Z(n5171) );
  AND U10343 ( .A(n5172), .B(p_input[5346]), .Z(o[5346]) );
  AND U10344 ( .A(p_input[25346]), .B(p_input[15346]), .Z(n5172) );
  AND U10345 ( .A(n5173), .B(p_input[5345]), .Z(o[5345]) );
  AND U10346 ( .A(p_input[25345]), .B(p_input[15345]), .Z(n5173) );
  AND U10347 ( .A(n5174), .B(p_input[5344]), .Z(o[5344]) );
  AND U10348 ( .A(p_input[25344]), .B(p_input[15344]), .Z(n5174) );
  AND U10349 ( .A(n5175), .B(p_input[5343]), .Z(o[5343]) );
  AND U10350 ( .A(p_input[25343]), .B(p_input[15343]), .Z(n5175) );
  AND U10351 ( .A(n5176), .B(p_input[5342]), .Z(o[5342]) );
  AND U10352 ( .A(p_input[25342]), .B(p_input[15342]), .Z(n5176) );
  AND U10353 ( .A(n5177), .B(p_input[5341]), .Z(o[5341]) );
  AND U10354 ( .A(p_input[25341]), .B(p_input[15341]), .Z(n5177) );
  AND U10355 ( .A(n5178), .B(p_input[5340]), .Z(o[5340]) );
  AND U10356 ( .A(p_input[25340]), .B(p_input[15340]), .Z(n5178) );
  AND U10357 ( .A(n5179), .B(p_input[533]), .Z(o[533]) );
  AND U10358 ( .A(p_input[20533]), .B(p_input[10533]), .Z(n5179) );
  AND U10359 ( .A(n5180), .B(p_input[5339]), .Z(o[5339]) );
  AND U10360 ( .A(p_input[25339]), .B(p_input[15339]), .Z(n5180) );
  AND U10361 ( .A(n5181), .B(p_input[5338]), .Z(o[5338]) );
  AND U10362 ( .A(p_input[25338]), .B(p_input[15338]), .Z(n5181) );
  AND U10363 ( .A(n5182), .B(p_input[5337]), .Z(o[5337]) );
  AND U10364 ( .A(p_input[25337]), .B(p_input[15337]), .Z(n5182) );
  AND U10365 ( .A(n5183), .B(p_input[5336]), .Z(o[5336]) );
  AND U10366 ( .A(p_input[25336]), .B(p_input[15336]), .Z(n5183) );
  AND U10367 ( .A(n5184), .B(p_input[5335]), .Z(o[5335]) );
  AND U10368 ( .A(p_input[25335]), .B(p_input[15335]), .Z(n5184) );
  AND U10369 ( .A(n5185), .B(p_input[5334]), .Z(o[5334]) );
  AND U10370 ( .A(p_input[25334]), .B(p_input[15334]), .Z(n5185) );
  AND U10371 ( .A(n5186), .B(p_input[5333]), .Z(o[5333]) );
  AND U10372 ( .A(p_input[25333]), .B(p_input[15333]), .Z(n5186) );
  AND U10373 ( .A(n5187), .B(p_input[5332]), .Z(o[5332]) );
  AND U10374 ( .A(p_input[25332]), .B(p_input[15332]), .Z(n5187) );
  AND U10375 ( .A(n5188), .B(p_input[5331]), .Z(o[5331]) );
  AND U10376 ( .A(p_input[25331]), .B(p_input[15331]), .Z(n5188) );
  AND U10377 ( .A(n5189), .B(p_input[5330]), .Z(o[5330]) );
  AND U10378 ( .A(p_input[25330]), .B(p_input[15330]), .Z(n5189) );
  AND U10379 ( .A(n5190), .B(p_input[532]), .Z(o[532]) );
  AND U10380 ( .A(p_input[20532]), .B(p_input[10532]), .Z(n5190) );
  AND U10381 ( .A(n5191), .B(p_input[5329]), .Z(o[5329]) );
  AND U10382 ( .A(p_input[25329]), .B(p_input[15329]), .Z(n5191) );
  AND U10383 ( .A(n5192), .B(p_input[5328]), .Z(o[5328]) );
  AND U10384 ( .A(p_input[25328]), .B(p_input[15328]), .Z(n5192) );
  AND U10385 ( .A(n5193), .B(p_input[5327]), .Z(o[5327]) );
  AND U10386 ( .A(p_input[25327]), .B(p_input[15327]), .Z(n5193) );
  AND U10387 ( .A(n5194), .B(p_input[5326]), .Z(o[5326]) );
  AND U10388 ( .A(p_input[25326]), .B(p_input[15326]), .Z(n5194) );
  AND U10389 ( .A(n5195), .B(p_input[5325]), .Z(o[5325]) );
  AND U10390 ( .A(p_input[25325]), .B(p_input[15325]), .Z(n5195) );
  AND U10391 ( .A(n5196), .B(p_input[5324]), .Z(o[5324]) );
  AND U10392 ( .A(p_input[25324]), .B(p_input[15324]), .Z(n5196) );
  AND U10393 ( .A(n5197), .B(p_input[5323]), .Z(o[5323]) );
  AND U10394 ( .A(p_input[25323]), .B(p_input[15323]), .Z(n5197) );
  AND U10395 ( .A(n5198), .B(p_input[5322]), .Z(o[5322]) );
  AND U10396 ( .A(p_input[25322]), .B(p_input[15322]), .Z(n5198) );
  AND U10397 ( .A(n5199), .B(p_input[5321]), .Z(o[5321]) );
  AND U10398 ( .A(p_input[25321]), .B(p_input[15321]), .Z(n5199) );
  AND U10399 ( .A(n5200), .B(p_input[5320]), .Z(o[5320]) );
  AND U10400 ( .A(p_input[25320]), .B(p_input[15320]), .Z(n5200) );
  AND U10401 ( .A(n5201), .B(p_input[531]), .Z(o[531]) );
  AND U10402 ( .A(p_input[20531]), .B(p_input[10531]), .Z(n5201) );
  AND U10403 ( .A(n5202), .B(p_input[5319]), .Z(o[5319]) );
  AND U10404 ( .A(p_input[25319]), .B(p_input[15319]), .Z(n5202) );
  AND U10405 ( .A(n5203), .B(p_input[5318]), .Z(o[5318]) );
  AND U10406 ( .A(p_input[25318]), .B(p_input[15318]), .Z(n5203) );
  AND U10407 ( .A(n5204), .B(p_input[5317]), .Z(o[5317]) );
  AND U10408 ( .A(p_input[25317]), .B(p_input[15317]), .Z(n5204) );
  AND U10409 ( .A(n5205), .B(p_input[5316]), .Z(o[5316]) );
  AND U10410 ( .A(p_input[25316]), .B(p_input[15316]), .Z(n5205) );
  AND U10411 ( .A(n5206), .B(p_input[5315]), .Z(o[5315]) );
  AND U10412 ( .A(p_input[25315]), .B(p_input[15315]), .Z(n5206) );
  AND U10413 ( .A(n5207), .B(p_input[5314]), .Z(o[5314]) );
  AND U10414 ( .A(p_input[25314]), .B(p_input[15314]), .Z(n5207) );
  AND U10415 ( .A(n5208), .B(p_input[5313]), .Z(o[5313]) );
  AND U10416 ( .A(p_input[25313]), .B(p_input[15313]), .Z(n5208) );
  AND U10417 ( .A(n5209), .B(p_input[5312]), .Z(o[5312]) );
  AND U10418 ( .A(p_input[25312]), .B(p_input[15312]), .Z(n5209) );
  AND U10419 ( .A(n5210), .B(p_input[5311]), .Z(o[5311]) );
  AND U10420 ( .A(p_input[25311]), .B(p_input[15311]), .Z(n5210) );
  AND U10421 ( .A(n5211), .B(p_input[5310]), .Z(o[5310]) );
  AND U10422 ( .A(p_input[25310]), .B(p_input[15310]), .Z(n5211) );
  AND U10423 ( .A(n5212), .B(p_input[530]), .Z(o[530]) );
  AND U10424 ( .A(p_input[20530]), .B(p_input[10530]), .Z(n5212) );
  AND U10425 ( .A(n5213), .B(p_input[5309]), .Z(o[5309]) );
  AND U10426 ( .A(p_input[25309]), .B(p_input[15309]), .Z(n5213) );
  AND U10427 ( .A(n5214), .B(p_input[5308]), .Z(o[5308]) );
  AND U10428 ( .A(p_input[25308]), .B(p_input[15308]), .Z(n5214) );
  AND U10429 ( .A(n5215), .B(p_input[5307]), .Z(o[5307]) );
  AND U10430 ( .A(p_input[25307]), .B(p_input[15307]), .Z(n5215) );
  AND U10431 ( .A(n5216), .B(p_input[5306]), .Z(o[5306]) );
  AND U10432 ( .A(p_input[25306]), .B(p_input[15306]), .Z(n5216) );
  AND U10433 ( .A(n5217), .B(p_input[5305]), .Z(o[5305]) );
  AND U10434 ( .A(p_input[25305]), .B(p_input[15305]), .Z(n5217) );
  AND U10435 ( .A(n5218), .B(p_input[5304]), .Z(o[5304]) );
  AND U10436 ( .A(p_input[25304]), .B(p_input[15304]), .Z(n5218) );
  AND U10437 ( .A(n5219), .B(p_input[5303]), .Z(o[5303]) );
  AND U10438 ( .A(p_input[25303]), .B(p_input[15303]), .Z(n5219) );
  AND U10439 ( .A(n5220), .B(p_input[5302]), .Z(o[5302]) );
  AND U10440 ( .A(p_input[25302]), .B(p_input[15302]), .Z(n5220) );
  AND U10441 ( .A(n5221), .B(p_input[5301]), .Z(o[5301]) );
  AND U10442 ( .A(p_input[25301]), .B(p_input[15301]), .Z(n5221) );
  AND U10443 ( .A(n5222), .B(p_input[5300]), .Z(o[5300]) );
  AND U10444 ( .A(p_input[25300]), .B(p_input[15300]), .Z(n5222) );
  AND U10445 ( .A(n5223), .B(p_input[52]), .Z(o[52]) );
  AND U10446 ( .A(p_input[20052]), .B(p_input[10052]), .Z(n5223) );
  AND U10447 ( .A(n5224), .B(p_input[529]), .Z(o[529]) );
  AND U10448 ( .A(p_input[20529]), .B(p_input[10529]), .Z(n5224) );
  AND U10449 ( .A(n5225), .B(p_input[5299]), .Z(o[5299]) );
  AND U10450 ( .A(p_input[25299]), .B(p_input[15299]), .Z(n5225) );
  AND U10451 ( .A(n5226), .B(p_input[5298]), .Z(o[5298]) );
  AND U10452 ( .A(p_input[25298]), .B(p_input[15298]), .Z(n5226) );
  AND U10453 ( .A(n5227), .B(p_input[5297]), .Z(o[5297]) );
  AND U10454 ( .A(p_input[25297]), .B(p_input[15297]), .Z(n5227) );
  AND U10455 ( .A(n5228), .B(p_input[5296]), .Z(o[5296]) );
  AND U10456 ( .A(p_input[25296]), .B(p_input[15296]), .Z(n5228) );
  AND U10457 ( .A(n5229), .B(p_input[5295]), .Z(o[5295]) );
  AND U10458 ( .A(p_input[25295]), .B(p_input[15295]), .Z(n5229) );
  AND U10459 ( .A(n5230), .B(p_input[5294]), .Z(o[5294]) );
  AND U10460 ( .A(p_input[25294]), .B(p_input[15294]), .Z(n5230) );
  AND U10461 ( .A(n5231), .B(p_input[5293]), .Z(o[5293]) );
  AND U10462 ( .A(p_input[25293]), .B(p_input[15293]), .Z(n5231) );
  AND U10463 ( .A(n5232), .B(p_input[5292]), .Z(o[5292]) );
  AND U10464 ( .A(p_input[25292]), .B(p_input[15292]), .Z(n5232) );
  AND U10465 ( .A(n5233), .B(p_input[5291]), .Z(o[5291]) );
  AND U10466 ( .A(p_input[25291]), .B(p_input[15291]), .Z(n5233) );
  AND U10467 ( .A(n5234), .B(p_input[5290]), .Z(o[5290]) );
  AND U10468 ( .A(p_input[25290]), .B(p_input[15290]), .Z(n5234) );
  AND U10469 ( .A(n5235), .B(p_input[528]), .Z(o[528]) );
  AND U10470 ( .A(p_input[20528]), .B(p_input[10528]), .Z(n5235) );
  AND U10471 ( .A(n5236), .B(p_input[5289]), .Z(o[5289]) );
  AND U10472 ( .A(p_input[25289]), .B(p_input[15289]), .Z(n5236) );
  AND U10473 ( .A(n5237), .B(p_input[5288]), .Z(o[5288]) );
  AND U10474 ( .A(p_input[25288]), .B(p_input[15288]), .Z(n5237) );
  AND U10475 ( .A(n5238), .B(p_input[5287]), .Z(o[5287]) );
  AND U10476 ( .A(p_input[25287]), .B(p_input[15287]), .Z(n5238) );
  AND U10477 ( .A(n5239), .B(p_input[5286]), .Z(o[5286]) );
  AND U10478 ( .A(p_input[25286]), .B(p_input[15286]), .Z(n5239) );
  AND U10479 ( .A(n5240), .B(p_input[5285]), .Z(o[5285]) );
  AND U10480 ( .A(p_input[25285]), .B(p_input[15285]), .Z(n5240) );
  AND U10481 ( .A(n5241), .B(p_input[5284]), .Z(o[5284]) );
  AND U10482 ( .A(p_input[25284]), .B(p_input[15284]), .Z(n5241) );
  AND U10483 ( .A(n5242), .B(p_input[5283]), .Z(o[5283]) );
  AND U10484 ( .A(p_input[25283]), .B(p_input[15283]), .Z(n5242) );
  AND U10485 ( .A(n5243), .B(p_input[5282]), .Z(o[5282]) );
  AND U10486 ( .A(p_input[25282]), .B(p_input[15282]), .Z(n5243) );
  AND U10487 ( .A(n5244), .B(p_input[5281]), .Z(o[5281]) );
  AND U10488 ( .A(p_input[25281]), .B(p_input[15281]), .Z(n5244) );
  AND U10489 ( .A(n5245), .B(p_input[5280]), .Z(o[5280]) );
  AND U10490 ( .A(p_input[25280]), .B(p_input[15280]), .Z(n5245) );
  AND U10491 ( .A(n5246), .B(p_input[527]), .Z(o[527]) );
  AND U10492 ( .A(p_input[20527]), .B(p_input[10527]), .Z(n5246) );
  AND U10493 ( .A(n5247), .B(p_input[5279]), .Z(o[5279]) );
  AND U10494 ( .A(p_input[25279]), .B(p_input[15279]), .Z(n5247) );
  AND U10495 ( .A(n5248), .B(p_input[5278]), .Z(o[5278]) );
  AND U10496 ( .A(p_input[25278]), .B(p_input[15278]), .Z(n5248) );
  AND U10497 ( .A(n5249), .B(p_input[5277]), .Z(o[5277]) );
  AND U10498 ( .A(p_input[25277]), .B(p_input[15277]), .Z(n5249) );
  AND U10499 ( .A(n5250), .B(p_input[5276]), .Z(o[5276]) );
  AND U10500 ( .A(p_input[25276]), .B(p_input[15276]), .Z(n5250) );
  AND U10501 ( .A(n5251), .B(p_input[5275]), .Z(o[5275]) );
  AND U10502 ( .A(p_input[25275]), .B(p_input[15275]), .Z(n5251) );
  AND U10503 ( .A(n5252), .B(p_input[5274]), .Z(o[5274]) );
  AND U10504 ( .A(p_input[25274]), .B(p_input[15274]), .Z(n5252) );
  AND U10505 ( .A(n5253), .B(p_input[5273]), .Z(o[5273]) );
  AND U10506 ( .A(p_input[25273]), .B(p_input[15273]), .Z(n5253) );
  AND U10507 ( .A(n5254), .B(p_input[5272]), .Z(o[5272]) );
  AND U10508 ( .A(p_input[25272]), .B(p_input[15272]), .Z(n5254) );
  AND U10509 ( .A(n5255), .B(p_input[5271]), .Z(o[5271]) );
  AND U10510 ( .A(p_input[25271]), .B(p_input[15271]), .Z(n5255) );
  AND U10511 ( .A(n5256), .B(p_input[5270]), .Z(o[5270]) );
  AND U10512 ( .A(p_input[25270]), .B(p_input[15270]), .Z(n5256) );
  AND U10513 ( .A(n5257), .B(p_input[526]), .Z(o[526]) );
  AND U10514 ( .A(p_input[20526]), .B(p_input[10526]), .Z(n5257) );
  AND U10515 ( .A(n5258), .B(p_input[5269]), .Z(o[5269]) );
  AND U10516 ( .A(p_input[25269]), .B(p_input[15269]), .Z(n5258) );
  AND U10517 ( .A(n5259), .B(p_input[5268]), .Z(o[5268]) );
  AND U10518 ( .A(p_input[25268]), .B(p_input[15268]), .Z(n5259) );
  AND U10519 ( .A(n5260), .B(p_input[5267]), .Z(o[5267]) );
  AND U10520 ( .A(p_input[25267]), .B(p_input[15267]), .Z(n5260) );
  AND U10521 ( .A(n5261), .B(p_input[5266]), .Z(o[5266]) );
  AND U10522 ( .A(p_input[25266]), .B(p_input[15266]), .Z(n5261) );
  AND U10523 ( .A(n5262), .B(p_input[5265]), .Z(o[5265]) );
  AND U10524 ( .A(p_input[25265]), .B(p_input[15265]), .Z(n5262) );
  AND U10525 ( .A(n5263), .B(p_input[5264]), .Z(o[5264]) );
  AND U10526 ( .A(p_input[25264]), .B(p_input[15264]), .Z(n5263) );
  AND U10527 ( .A(n5264), .B(p_input[5263]), .Z(o[5263]) );
  AND U10528 ( .A(p_input[25263]), .B(p_input[15263]), .Z(n5264) );
  AND U10529 ( .A(n5265), .B(p_input[5262]), .Z(o[5262]) );
  AND U10530 ( .A(p_input[25262]), .B(p_input[15262]), .Z(n5265) );
  AND U10531 ( .A(n5266), .B(p_input[5261]), .Z(o[5261]) );
  AND U10532 ( .A(p_input[25261]), .B(p_input[15261]), .Z(n5266) );
  AND U10533 ( .A(n5267), .B(p_input[5260]), .Z(o[5260]) );
  AND U10534 ( .A(p_input[25260]), .B(p_input[15260]), .Z(n5267) );
  AND U10535 ( .A(n5268), .B(p_input[525]), .Z(o[525]) );
  AND U10536 ( .A(p_input[20525]), .B(p_input[10525]), .Z(n5268) );
  AND U10537 ( .A(n5269), .B(p_input[5259]), .Z(o[5259]) );
  AND U10538 ( .A(p_input[25259]), .B(p_input[15259]), .Z(n5269) );
  AND U10539 ( .A(n5270), .B(p_input[5258]), .Z(o[5258]) );
  AND U10540 ( .A(p_input[25258]), .B(p_input[15258]), .Z(n5270) );
  AND U10541 ( .A(n5271), .B(p_input[5257]), .Z(o[5257]) );
  AND U10542 ( .A(p_input[25257]), .B(p_input[15257]), .Z(n5271) );
  AND U10543 ( .A(n5272), .B(p_input[5256]), .Z(o[5256]) );
  AND U10544 ( .A(p_input[25256]), .B(p_input[15256]), .Z(n5272) );
  AND U10545 ( .A(n5273), .B(p_input[5255]), .Z(o[5255]) );
  AND U10546 ( .A(p_input[25255]), .B(p_input[15255]), .Z(n5273) );
  AND U10547 ( .A(n5274), .B(p_input[5254]), .Z(o[5254]) );
  AND U10548 ( .A(p_input[25254]), .B(p_input[15254]), .Z(n5274) );
  AND U10549 ( .A(n5275), .B(p_input[5253]), .Z(o[5253]) );
  AND U10550 ( .A(p_input[25253]), .B(p_input[15253]), .Z(n5275) );
  AND U10551 ( .A(n5276), .B(p_input[5252]), .Z(o[5252]) );
  AND U10552 ( .A(p_input[25252]), .B(p_input[15252]), .Z(n5276) );
  AND U10553 ( .A(n5277), .B(p_input[5251]), .Z(o[5251]) );
  AND U10554 ( .A(p_input[25251]), .B(p_input[15251]), .Z(n5277) );
  AND U10555 ( .A(n5278), .B(p_input[5250]), .Z(o[5250]) );
  AND U10556 ( .A(p_input[25250]), .B(p_input[15250]), .Z(n5278) );
  AND U10557 ( .A(n5279), .B(p_input[524]), .Z(o[524]) );
  AND U10558 ( .A(p_input[20524]), .B(p_input[10524]), .Z(n5279) );
  AND U10559 ( .A(n5280), .B(p_input[5249]), .Z(o[5249]) );
  AND U10560 ( .A(p_input[25249]), .B(p_input[15249]), .Z(n5280) );
  AND U10561 ( .A(n5281), .B(p_input[5248]), .Z(o[5248]) );
  AND U10562 ( .A(p_input[25248]), .B(p_input[15248]), .Z(n5281) );
  AND U10563 ( .A(n5282), .B(p_input[5247]), .Z(o[5247]) );
  AND U10564 ( .A(p_input[25247]), .B(p_input[15247]), .Z(n5282) );
  AND U10565 ( .A(n5283), .B(p_input[5246]), .Z(o[5246]) );
  AND U10566 ( .A(p_input[25246]), .B(p_input[15246]), .Z(n5283) );
  AND U10567 ( .A(n5284), .B(p_input[5245]), .Z(o[5245]) );
  AND U10568 ( .A(p_input[25245]), .B(p_input[15245]), .Z(n5284) );
  AND U10569 ( .A(n5285), .B(p_input[5244]), .Z(o[5244]) );
  AND U10570 ( .A(p_input[25244]), .B(p_input[15244]), .Z(n5285) );
  AND U10571 ( .A(n5286), .B(p_input[5243]), .Z(o[5243]) );
  AND U10572 ( .A(p_input[25243]), .B(p_input[15243]), .Z(n5286) );
  AND U10573 ( .A(n5287), .B(p_input[5242]), .Z(o[5242]) );
  AND U10574 ( .A(p_input[25242]), .B(p_input[15242]), .Z(n5287) );
  AND U10575 ( .A(n5288), .B(p_input[5241]), .Z(o[5241]) );
  AND U10576 ( .A(p_input[25241]), .B(p_input[15241]), .Z(n5288) );
  AND U10577 ( .A(n5289), .B(p_input[5240]), .Z(o[5240]) );
  AND U10578 ( .A(p_input[25240]), .B(p_input[15240]), .Z(n5289) );
  AND U10579 ( .A(n5290), .B(p_input[523]), .Z(o[523]) );
  AND U10580 ( .A(p_input[20523]), .B(p_input[10523]), .Z(n5290) );
  AND U10581 ( .A(n5291), .B(p_input[5239]), .Z(o[5239]) );
  AND U10582 ( .A(p_input[25239]), .B(p_input[15239]), .Z(n5291) );
  AND U10583 ( .A(n5292), .B(p_input[5238]), .Z(o[5238]) );
  AND U10584 ( .A(p_input[25238]), .B(p_input[15238]), .Z(n5292) );
  AND U10585 ( .A(n5293), .B(p_input[5237]), .Z(o[5237]) );
  AND U10586 ( .A(p_input[25237]), .B(p_input[15237]), .Z(n5293) );
  AND U10587 ( .A(n5294), .B(p_input[5236]), .Z(o[5236]) );
  AND U10588 ( .A(p_input[25236]), .B(p_input[15236]), .Z(n5294) );
  AND U10589 ( .A(n5295), .B(p_input[5235]), .Z(o[5235]) );
  AND U10590 ( .A(p_input[25235]), .B(p_input[15235]), .Z(n5295) );
  AND U10591 ( .A(n5296), .B(p_input[5234]), .Z(o[5234]) );
  AND U10592 ( .A(p_input[25234]), .B(p_input[15234]), .Z(n5296) );
  AND U10593 ( .A(n5297), .B(p_input[5233]), .Z(o[5233]) );
  AND U10594 ( .A(p_input[25233]), .B(p_input[15233]), .Z(n5297) );
  AND U10595 ( .A(n5298), .B(p_input[5232]), .Z(o[5232]) );
  AND U10596 ( .A(p_input[25232]), .B(p_input[15232]), .Z(n5298) );
  AND U10597 ( .A(n5299), .B(p_input[5231]), .Z(o[5231]) );
  AND U10598 ( .A(p_input[25231]), .B(p_input[15231]), .Z(n5299) );
  AND U10599 ( .A(n5300), .B(p_input[5230]), .Z(o[5230]) );
  AND U10600 ( .A(p_input[25230]), .B(p_input[15230]), .Z(n5300) );
  AND U10601 ( .A(n5301), .B(p_input[522]), .Z(o[522]) );
  AND U10602 ( .A(p_input[20522]), .B(p_input[10522]), .Z(n5301) );
  AND U10603 ( .A(n5302), .B(p_input[5229]), .Z(o[5229]) );
  AND U10604 ( .A(p_input[25229]), .B(p_input[15229]), .Z(n5302) );
  AND U10605 ( .A(n5303), .B(p_input[5228]), .Z(o[5228]) );
  AND U10606 ( .A(p_input[25228]), .B(p_input[15228]), .Z(n5303) );
  AND U10607 ( .A(n5304), .B(p_input[5227]), .Z(o[5227]) );
  AND U10608 ( .A(p_input[25227]), .B(p_input[15227]), .Z(n5304) );
  AND U10609 ( .A(n5305), .B(p_input[5226]), .Z(o[5226]) );
  AND U10610 ( .A(p_input[25226]), .B(p_input[15226]), .Z(n5305) );
  AND U10611 ( .A(n5306), .B(p_input[5225]), .Z(o[5225]) );
  AND U10612 ( .A(p_input[25225]), .B(p_input[15225]), .Z(n5306) );
  AND U10613 ( .A(n5307), .B(p_input[5224]), .Z(o[5224]) );
  AND U10614 ( .A(p_input[25224]), .B(p_input[15224]), .Z(n5307) );
  AND U10615 ( .A(n5308), .B(p_input[5223]), .Z(o[5223]) );
  AND U10616 ( .A(p_input[25223]), .B(p_input[15223]), .Z(n5308) );
  AND U10617 ( .A(n5309), .B(p_input[5222]), .Z(o[5222]) );
  AND U10618 ( .A(p_input[25222]), .B(p_input[15222]), .Z(n5309) );
  AND U10619 ( .A(n5310), .B(p_input[5221]), .Z(o[5221]) );
  AND U10620 ( .A(p_input[25221]), .B(p_input[15221]), .Z(n5310) );
  AND U10621 ( .A(n5311), .B(p_input[5220]), .Z(o[5220]) );
  AND U10622 ( .A(p_input[25220]), .B(p_input[15220]), .Z(n5311) );
  AND U10623 ( .A(n5312), .B(p_input[521]), .Z(o[521]) );
  AND U10624 ( .A(p_input[20521]), .B(p_input[10521]), .Z(n5312) );
  AND U10625 ( .A(n5313), .B(p_input[5219]), .Z(o[5219]) );
  AND U10626 ( .A(p_input[25219]), .B(p_input[15219]), .Z(n5313) );
  AND U10627 ( .A(n5314), .B(p_input[5218]), .Z(o[5218]) );
  AND U10628 ( .A(p_input[25218]), .B(p_input[15218]), .Z(n5314) );
  AND U10629 ( .A(n5315), .B(p_input[5217]), .Z(o[5217]) );
  AND U10630 ( .A(p_input[25217]), .B(p_input[15217]), .Z(n5315) );
  AND U10631 ( .A(n5316), .B(p_input[5216]), .Z(o[5216]) );
  AND U10632 ( .A(p_input[25216]), .B(p_input[15216]), .Z(n5316) );
  AND U10633 ( .A(n5317), .B(p_input[5215]), .Z(o[5215]) );
  AND U10634 ( .A(p_input[25215]), .B(p_input[15215]), .Z(n5317) );
  AND U10635 ( .A(n5318), .B(p_input[5214]), .Z(o[5214]) );
  AND U10636 ( .A(p_input[25214]), .B(p_input[15214]), .Z(n5318) );
  AND U10637 ( .A(n5319), .B(p_input[5213]), .Z(o[5213]) );
  AND U10638 ( .A(p_input[25213]), .B(p_input[15213]), .Z(n5319) );
  AND U10639 ( .A(n5320), .B(p_input[5212]), .Z(o[5212]) );
  AND U10640 ( .A(p_input[25212]), .B(p_input[15212]), .Z(n5320) );
  AND U10641 ( .A(n5321), .B(p_input[5211]), .Z(o[5211]) );
  AND U10642 ( .A(p_input[25211]), .B(p_input[15211]), .Z(n5321) );
  AND U10643 ( .A(n5322), .B(p_input[5210]), .Z(o[5210]) );
  AND U10644 ( .A(p_input[25210]), .B(p_input[15210]), .Z(n5322) );
  AND U10645 ( .A(n5323), .B(p_input[520]), .Z(o[520]) );
  AND U10646 ( .A(p_input[20520]), .B(p_input[10520]), .Z(n5323) );
  AND U10647 ( .A(n5324), .B(p_input[5209]), .Z(o[5209]) );
  AND U10648 ( .A(p_input[25209]), .B(p_input[15209]), .Z(n5324) );
  AND U10649 ( .A(n5325), .B(p_input[5208]), .Z(o[5208]) );
  AND U10650 ( .A(p_input[25208]), .B(p_input[15208]), .Z(n5325) );
  AND U10651 ( .A(n5326), .B(p_input[5207]), .Z(o[5207]) );
  AND U10652 ( .A(p_input[25207]), .B(p_input[15207]), .Z(n5326) );
  AND U10653 ( .A(n5327), .B(p_input[5206]), .Z(o[5206]) );
  AND U10654 ( .A(p_input[25206]), .B(p_input[15206]), .Z(n5327) );
  AND U10655 ( .A(n5328), .B(p_input[5205]), .Z(o[5205]) );
  AND U10656 ( .A(p_input[25205]), .B(p_input[15205]), .Z(n5328) );
  AND U10657 ( .A(n5329), .B(p_input[5204]), .Z(o[5204]) );
  AND U10658 ( .A(p_input[25204]), .B(p_input[15204]), .Z(n5329) );
  AND U10659 ( .A(n5330), .B(p_input[5203]), .Z(o[5203]) );
  AND U10660 ( .A(p_input[25203]), .B(p_input[15203]), .Z(n5330) );
  AND U10661 ( .A(n5331), .B(p_input[5202]), .Z(o[5202]) );
  AND U10662 ( .A(p_input[25202]), .B(p_input[15202]), .Z(n5331) );
  AND U10663 ( .A(n5332), .B(p_input[5201]), .Z(o[5201]) );
  AND U10664 ( .A(p_input[25201]), .B(p_input[15201]), .Z(n5332) );
  AND U10665 ( .A(n5333), .B(p_input[5200]), .Z(o[5200]) );
  AND U10666 ( .A(p_input[25200]), .B(p_input[15200]), .Z(n5333) );
  AND U10667 ( .A(n5334), .B(p_input[51]), .Z(o[51]) );
  AND U10668 ( .A(p_input[20051]), .B(p_input[10051]), .Z(n5334) );
  AND U10669 ( .A(n5335), .B(p_input[519]), .Z(o[519]) );
  AND U10670 ( .A(p_input[20519]), .B(p_input[10519]), .Z(n5335) );
  AND U10671 ( .A(n5336), .B(p_input[5199]), .Z(o[5199]) );
  AND U10672 ( .A(p_input[25199]), .B(p_input[15199]), .Z(n5336) );
  AND U10673 ( .A(n5337), .B(p_input[5198]), .Z(o[5198]) );
  AND U10674 ( .A(p_input[25198]), .B(p_input[15198]), .Z(n5337) );
  AND U10675 ( .A(n5338), .B(p_input[5197]), .Z(o[5197]) );
  AND U10676 ( .A(p_input[25197]), .B(p_input[15197]), .Z(n5338) );
  AND U10677 ( .A(n5339), .B(p_input[5196]), .Z(o[5196]) );
  AND U10678 ( .A(p_input[25196]), .B(p_input[15196]), .Z(n5339) );
  AND U10679 ( .A(n5340), .B(p_input[5195]), .Z(o[5195]) );
  AND U10680 ( .A(p_input[25195]), .B(p_input[15195]), .Z(n5340) );
  AND U10681 ( .A(n5341), .B(p_input[5194]), .Z(o[5194]) );
  AND U10682 ( .A(p_input[25194]), .B(p_input[15194]), .Z(n5341) );
  AND U10683 ( .A(n5342), .B(p_input[5193]), .Z(o[5193]) );
  AND U10684 ( .A(p_input[25193]), .B(p_input[15193]), .Z(n5342) );
  AND U10685 ( .A(n5343), .B(p_input[5192]), .Z(o[5192]) );
  AND U10686 ( .A(p_input[25192]), .B(p_input[15192]), .Z(n5343) );
  AND U10687 ( .A(n5344), .B(p_input[5191]), .Z(o[5191]) );
  AND U10688 ( .A(p_input[25191]), .B(p_input[15191]), .Z(n5344) );
  AND U10689 ( .A(n5345), .B(p_input[5190]), .Z(o[5190]) );
  AND U10690 ( .A(p_input[25190]), .B(p_input[15190]), .Z(n5345) );
  AND U10691 ( .A(n5346), .B(p_input[518]), .Z(o[518]) );
  AND U10692 ( .A(p_input[20518]), .B(p_input[10518]), .Z(n5346) );
  AND U10693 ( .A(n5347), .B(p_input[5189]), .Z(o[5189]) );
  AND U10694 ( .A(p_input[25189]), .B(p_input[15189]), .Z(n5347) );
  AND U10695 ( .A(n5348), .B(p_input[5188]), .Z(o[5188]) );
  AND U10696 ( .A(p_input[25188]), .B(p_input[15188]), .Z(n5348) );
  AND U10697 ( .A(n5349), .B(p_input[5187]), .Z(o[5187]) );
  AND U10698 ( .A(p_input[25187]), .B(p_input[15187]), .Z(n5349) );
  AND U10699 ( .A(n5350), .B(p_input[5186]), .Z(o[5186]) );
  AND U10700 ( .A(p_input[25186]), .B(p_input[15186]), .Z(n5350) );
  AND U10701 ( .A(n5351), .B(p_input[5185]), .Z(o[5185]) );
  AND U10702 ( .A(p_input[25185]), .B(p_input[15185]), .Z(n5351) );
  AND U10703 ( .A(n5352), .B(p_input[5184]), .Z(o[5184]) );
  AND U10704 ( .A(p_input[25184]), .B(p_input[15184]), .Z(n5352) );
  AND U10705 ( .A(n5353), .B(p_input[5183]), .Z(o[5183]) );
  AND U10706 ( .A(p_input[25183]), .B(p_input[15183]), .Z(n5353) );
  AND U10707 ( .A(n5354), .B(p_input[5182]), .Z(o[5182]) );
  AND U10708 ( .A(p_input[25182]), .B(p_input[15182]), .Z(n5354) );
  AND U10709 ( .A(n5355), .B(p_input[5181]), .Z(o[5181]) );
  AND U10710 ( .A(p_input[25181]), .B(p_input[15181]), .Z(n5355) );
  AND U10711 ( .A(n5356), .B(p_input[5180]), .Z(o[5180]) );
  AND U10712 ( .A(p_input[25180]), .B(p_input[15180]), .Z(n5356) );
  AND U10713 ( .A(n5357), .B(p_input[517]), .Z(o[517]) );
  AND U10714 ( .A(p_input[20517]), .B(p_input[10517]), .Z(n5357) );
  AND U10715 ( .A(n5358), .B(p_input[5179]), .Z(o[5179]) );
  AND U10716 ( .A(p_input[25179]), .B(p_input[15179]), .Z(n5358) );
  AND U10717 ( .A(n5359), .B(p_input[5178]), .Z(o[5178]) );
  AND U10718 ( .A(p_input[25178]), .B(p_input[15178]), .Z(n5359) );
  AND U10719 ( .A(n5360), .B(p_input[5177]), .Z(o[5177]) );
  AND U10720 ( .A(p_input[25177]), .B(p_input[15177]), .Z(n5360) );
  AND U10721 ( .A(n5361), .B(p_input[5176]), .Z(o[5176]) );
  AND U10722 ( .A(p_input[25176]), .B(p_input[15176]), .Z(n5361) );
  AND U10723 ( .A(n5362), .B(p_input[5175]), .Z(o[5175]) );
  AND U10724 ( .A(p_input[25175]), .B(p_input[15175]), .Z(n5362) );
  AND U10725 ( .A(n5363), .B(p_input[5174]), .Z(o[5174]) );
  AND U10726 ( .A(p_input[25174]), .B(p_input[15174]), .Z(n5363) );
  AND U10727 ( .A(n5364), .B(p_input[5173]), .Z(o[5173]) );
  AND U10728 ( .A(p_input[25173]), .B(p_input[15173]), .Z(n5364) );
  AND U10729 ( .A(n5365), .B(p_input[5172]), .Z(o[5172]) );
  AND U10730 ( .A(p_input[25172]), .B(p_input[15172]), .Z(n5365) );
  AND U10731 ( .A(n5366), .B(p_input[5171]), .Z(o[5171]) );
  AND U10732 ( .A(p_input[25171]), .B(p_input[15171]), .Z(n5366) );
  AND U10733 ( .A(n5367), .B(p_input[5170]), .Z(o[5170]) );
  AND U10734 ( .A(p_input[25170]), .B(p_input[15170]), .Z(n5367) );
  AND U10735 ( .A(n5368), .B(p_input[516]), .Z(o[516]) );
  AND U10736 ( .A(p_input[20516]), .B(p_input[10516]), .Z(n5368) );
  AND U10737 ( .A(n5369), .B(p_input[5169]), .Z(o[5169]) );
  AND U10738 ( .A(p_input[25169]), .B(p_input[15169]), .Z(n5369) );
  AND U10739 ( .A(n5370), .B(p_input[5168]), .Z(o[5168]) );
  AND U10740 ( .A(p_input[25168]), .B(p_input[15168]), .Z(n5370) );
  AND U10741 ( .A(n5371), .B(p_input[5167]), .Z(o[5167]) );
  AND U10742 ( .A(p_input[25167]), .B(p_input[15167]), .Z(n5371) );
  AND U10743 ( .A(n5372), .B(p_input[5166]), .Z(o[5166]) );
  AND U10744 ( .A(p_input[25166]), .B(p_input[15166]), .Z(n5372) );
  AND U10745 ( .A(n5373), .B(p_input[5165]), .Z(o[5165]) );
  AND U10746 ( .A(p_input[25165]), .B(p_input[15165]), .Z(n5373) );
  AND U10747 ( .A(n5374), .B(p_input[5164]), .Z(o[5164]) );
  AND U10748 ( .A(p_input[25164]), .B(p_input[15164]), .Z(n5374) );
  AND U10749 ( .A(n5375), .B(p_input[5163]), .Z(o[5163]) );
  AND U10750 ( .A(p_input[25163]), .B(p_input[15163]), .Z(n5375) );
  AND U10751 ( .A(n5376), .B(p_input[5162]), .Z(o[5162]) );
  AND U10752 ( .A(p_input[25162]), .B(p_input[15162]), .Z(n5376) );
  AND U10753 ( .A(n5377), .B(p_input[5161]), .Z(o[5161]) );
  AND U10754 ( .A(p_input[25161]), .B(p_input[15161]), .Z(n5377) );
  AND U10755 ( .A(n5378), .B(p_input[5160]), .Z(o[5160]) );
  AND U10756 ( .A(p_input[25160]), .B(p_input[15160]), .Z(n5378) );
  AND U10757 ( .A(n5379), .B(p_input[515]), .Z(o[515]) );
  AND U10758 ( .A(p_input[20515]), .B(p_input[10515]), .Z(n5379) );
  AND U10759 ( .A(n5380), .B(p_input[5159]), .Z(o[5159]) );
  AND U10760 ( .A(p_input[25159]), .B(p_input[15159]), .Z(n5380) );
  AND U10761 ( .A(n5381), .B(p_input[5158]), .Z(o[5158]) );
  AND U10762 ( .A(p_input[25158]), .B(p_input[15158]), .Z(n5381) );
  AND U10763 ( .A(n5382), .B(p_input[5157]), .Z(o[5157]) );
  AND U10764 ( .A(p_input[25157]), .B(p_input[15157]), .Z(n5382) );
  AND U10765 ( .A(n5383), .B(p_input[5156]), .Z(o[5156]) );
  AND U10766 ( .A(p_input[25156]), .B(p_input[15156]), .Z(n5383) );
  AND U10767 ( .A(n5384), .B(p_input[5155]), .Z(o[5155]) );
  AND U10768 ( .A(p_input[25155]), .B(p_input[15155]), .Z(n5384) );
  AND U10769 ( .A(n5385), .B(p_input[5154]), .Z(o[5154]) );
  AND U10770 ( .A(p_input[25154]), .B(p_input[15154]), .Z(n5385) );
  AND U10771 ( .A(n5386), .B(p_input[5153]), .Z(o[5153]) );
  AND U10772 ( .A(p_input[25153]), .B(p_input[15153]), .Z(n5386) );
  AND U10773 ( .A(n5387), .B(p_input[5152]), .Z(o[5152]) );
  AND U10774 ( .A(p_input[25152]), .B(p_input[15152]), .Z(n5387) );
  AND U10775 ( .A(n5388), .B(p_input[5151]), .Z(o[5151]) );
  AND U10776 ( .A(p_input[25151]), .B(p_input[15151]), .Z(n5388) );
  AND U10777 ( .A(n5389), .B(p_input[5150]), .Z(o[5150]) );
  AND U10778 ( .A(p_input[25150]), .B(p_input[15150]), .Z(n5389) );
  AND U10779 ( .A(n5390), .B(p_input[514]), .Z(o[514]) );
  AND U10780 ( .A(p_input[20514]), .B(p_input[10514]), .Z(n5390) );
  AND U10781 ( .A(n5391), .B(p_input[5149]), .Z(o[5149]) );
  AND U10782 ( .A(p_input[25149]), .B(p_input[15149]), .Z(n5391) );
  AND U10783 ( .A(n5392), .B(p_input[5148]), .Z(o[5148]) );
  AND U10784 ( .A(p_input[25148]), .B(p_input[15148]), .Z(n5392) );
  AND U10785 ( .A(n5393), .B(p_input[5147]), .Z(o[5147]) );
  AND U10786 ( .A(p_input[25147]), .B(p_input[15147]), .Z(n5393) );
  AND U10787 ( .A(n5394), .B(p_input[5146]), .Z(o[5146]) );
  AND U10788 ( .A(p_input[25146]), .B(p_input[15146]), .Z(n5394) );
  AND U10789 ( .A(n5395), .B(p_input[5145]), .Z(o[5145]) );
  AND U10790 ( .A(p_input[25145]), .B(p_input[15145]), .Z(n5395) );
  AND U10791 ( .A(n5396), .B(p_input[5144]), .Z(o[5144]) );
  AND U10792 ( .A(p_input[25144]), .B(p_input[15144]), .Z(n5396) );
  AND U10793 ( .A(n5397), .B(p_input[5143]), .Z(o[5143]) );
  AND U10794 ( .A(p_input[25143]), .B(p_input[15143]), .Z(n5397) );
  AND U10795 ( .A(n5398), .B(p_input[5142]), .Z(o[5142]) );
  AND U10796 ( .A(p_input[25142]), .B(p_input[15142]), .Z(n5398) );
  AND U10797 ( .A(n5399), .B(p_input[5141]), .Z(o[5141]) );
  AND U10798 ( .A(p_input[25141]), .B(p_input[15141]), .Z(n5399) );
  AND U10799 ( .A(n5400), .B(p_input[5140]), .Z(o[5140]) );
  AND U10800 ( .A(p_input[25140]), .B(p_input[15140]), .Z(n5400) );
  AND U10801 ( .A(n5401), .B(p_input[513]), .Z(o[513]) );
  AND U10802 ( .A(p_input[20513]), .B(p_input[10513]), .Z(n5401) );
  AND U10803 ( .A(n5402), .B(p_input[5139]), .Z(o[5139]) );
  AND U10804 ( .A(p_input[25139]), .B(p_input[15139]), .Z(n5402) );
  AND U10805 ( .A(n5403), .B(p_input[5138]), .Z(o[5138]) );
  AND U10806 ( .A(p_input[25138]), .B(p_input[15138]), .Z(n5403) );
  AND U10807 ( .A(n5404), .B(p_input[5137]), .Z(o[5137]) );
  AND U10808 ( .A(p_input[25137]), .B(p_input[15137]), .Z(n5404) );
  AND U10809 ( .A(n5405), .B(p_input[5136]), .Z(o[5136]) );
  AND U10810 ( .A(p_input[25136]), .B(p_input[15136]), .Z(n5405) );
  AND U10811 ( .A(n5406), .B(p_input[5135]), .Z(o[5135]) );
  AND U10812 ( .A(p_input[25135]), .B(p_input[15135]), .Z(n5406) );
  AND U10813 ( .A(n5407), .B(p_input[5134]), .Z(o[5134]) );
  AND U10814 ( .A(p_input[25134]), .B(p_input[15134]), .Z(n5407) );
  AND U10815 ( .A(n5408), .B(p_input[5133]), .Z(o[5133]) );
  AND U10816 ( .A(p_input[25133]), .B(p_input[15133]), .Z(n5408) );
  AND U10817 ( .A(n5409), .B(p_input[5132]), .Z(o[5132]) );
  AND U10818 ( .A(p_input[25132]), .B(p_input[15132]), .Z(n5409) );
  AND U10819 ( .A(n5410), .B(p_input[5131]), .Z(o[5131]) );
  AND U10820 ( .A(p_input[25131]), .B(p_input[15131]), .Z(n5410) );
  AND U10821 ( .A(n5411), .B(p_input[5130]), .Z(o[5130]) );
  AND U10822 ( .A(p_input[25130]), .B(p_input[15130]), .Z(n5411) );
  AND U10823 ( .A(n5412), .B(p_input[512]), .Z(o[512]) );
  AND U10824 ( .A(p_input[20512]), .B(p_input[10512]), .Z(n5412) );
  AND U10825 ( .A(n5413), .B(p_input[5129]), .Z(o[5129]) );
  AND U10826 ( .A(p_input[25129]), .B(p_input[15129]), .Z(n5413) );
  AND U10827 ( .A(n5414), .B(p_input[5128]), .Z(o[5128]) );
  AND U10828 ( .A(p_input[25128]), .B(p_input[15128]), .Z(n5414) );
  AND U10829 ( .A(n5415), .B(p_input[5127]), .Z(o[5127]) );
  AND U10830 ( .A(p_input[25127]), .B(p_input[15127]), .Z(n5415) );
  AND U10831 ( .A(n5416), .B(p_input[5126]), .Z(o[5126]) );
  AND U10832 ( .A(p_input[25126]), .B(p_input[15126]), .Z(n5416) );
  AND U10833 ( .A(n5417), .B(p_input[5125]), .Z(o[5125]) );
  AND U10834 ( .A(p_input[25125]), .B(p_input[15125]), .Z(n5417) );
  AND U10835 ( .A(n5418), .B(p_input[5124]), .Z(o[5124]) );
  AND U10836 ( .A(p_input[25124]), .B(p_input[15124]), .Z(n5418) );
  AND U10837 ( .A(n5419), .B(p_input[5123]), .Z(o[5123]) );
  AND U10838 ( .A(p_input[25123]), .B(p_input[15123]), .Z(n5419) );
  AND U10839 ( .A(n5420), .B(p_input[5122]), .Z(o[5122]) );
  AND U10840 ( .A(p_input[25122]), .B(p_input[15122]), .Z(n5420) );
  AND U10841 ( .A(n5421), .B(p_input[5121]), .Z(o[5121]) );
  AND U10842 ( .A(p_input[25121]), .B(p_input[15121]), .Z(n5421) );
  AND U10843 ( .A(n5422), .B(p_input[5120]), .Z(o[5120]) );
  AND U10844 ( .A(p_input[25120]), .B(p_input[15120]), .Z(n5422) );
  AND U10845 ( .A(n5423), .B(p_input[511]), .Z(o[511]) );
  AND U10846 ( .A(p_input[20511]), .B(p_input[10511]), .Z(n5423) );
  AND U10847 ( .A(n5424), .B(p_input[5119]), .Z(o[5119]) );
  AND U10848 ( .A(p_input[25119]), .B(p_input[15119]), .Z(n5424) );
  AND U10849 ( .A(n5425), .B(p_input[5118]), .Z(o[5118]) );
  AND U10850 ( .A(p_input[25118]), .B(p_input[15118]), .Z(n5425) );
  AND U10851 ( .A(n5426), .B(p_input[5117]), .Z(o[5117]) );
  AND U10852 ( .A(p_input[25117]), .B(p_input[15117]), .Z(n5426) );
  AND U10853 ( .A(n5427), .B(p_input[5116]), .Z(o[5116]) );
  AND U10854 ( .A(p_input[25116]), .B(p_input[15116]), .Z(n5427) );
  AND U10855 ( .A(n5428), .B(p_input[5115]), .Z(o[5115]) );
  AND U10856 ( .A(p_input[25115]), .B(p_input[15115]), .Z(n5428) );
  AND U10857 ( .A(n5429), .B(p_input[5114]), .Z(o[5114]) );
  AND U10858 ( .A(p_input[25114]), .B(p_input[15114]), .Z(n5429) );
  AND U10859 ( .A(n5430), .B(p_input[5113]), .Z(o[5113]) );
  AND U10860 ( .A(p_input[25113]), .B(p_input[15113]), .Z(n5430) );
  AND U10861 ( .A(n5431), .B(p_input[5112]), .Z(o[5112]) );
  AND U10862 ( .A(p_input[25112]), .B(p_input[15112]), .Z(n5431) );
  AND U10863 ( .A(n5432), .B(p_input[5111]), .Z(o[5111]) );
  AND U10864 ( .A(p_input[25111]), .B(p_input[15111]), .Z(n5432) );
  AND U10865 ( .A(n5433), .B(p_input[5110]), .Z(o[5110]) );
  AND U10866 ( .A(p_input[25110]), .B(p_input[15110]), .Z(n5433) );
  AND U10867 ( .A(n5434), .B(p_input[510]), .Z(o[510]) );
  AND U10868 ( .A(p_input[20510]), .B(p_input[10510]), .Z(n5434) );
  AND U10869 ( .A(n5435), .B(p_input[5109]), .Z(o[5109]) );
  AND U10870 ( .A(p_input[25109]), .B(p_input[15109]), .Z(n5435) );
  AND U10871 ( .A(n5436), .B(p_input[5108]), .Z(o[5108]) );
  AND U10872 ( .A(p_input[25108]), .B(p_input[15108]), .Z(n5436) );
  AND U10873 ( .A(n5437), .B(p_input[5107]), .Z(o[5107]) );
  AND U10874 ( .A(p_input[25107]), .B(p_input[15107]), .Z(n5437) );
  AND U10875 ( .A(n5438), .B(p_input[5106]), .Z(o[5106]) );
  AND U10876 ( .A(p_input[25106]), .B(p_input[15106]), .Z(n5438) );
  AND U10877 ( .A(n5439), .B(p_input[5105]), .Z(o[5105]) );
  AND U10878 ( .A(p_input[25105]), .B(p_input[15105]), .Z(n5439) );
  AND U10879 ( .A(n5440), .B(p_input[5104]), .Z(o[5104]) );
  AND U10880 ( .A(p_input[25104]), .B(p_input[15104]), .Z(n5440) );
  AND U10881 ( .A(n5441), .B(p_input[5103]), .Z(o[5103]) );
  AND U10882 ( .A(p_input[25103]), .B(p_input[15103]), .Z(n5441) );
  AND U10883 ( .A(n5442), .B(p_input[5102]), .Z(o[5102]) );
  AND U10884 ( .A(p_input[25102]), .B(p_input[15102]), .Z(n5442) );
  AND U10885 ( .A(n5443), .B(p_input[5101]), .Z(o[5101]) );
  AND U10886 ( .A(p_input[25101]), .B(p_input[15101]), .Z(n5443) );
  AND U10887 ( .A(n5444), .B(p_input[5100]), .Z(o[5100]) );
  AND U10888 ( .A(p_input[25100]), .B(p_input[15100]), .Z(n5444) );
  AND U10889 ( .A(n5445), .B(p_input[50]), .Z(o[50]) );
  AND U10890 ( .A(p_input[20050]), .B(p_input[10050]), .Z(n5445) );
  AND U10891 ( .A(n5446), .B(p_input[509]), .Z(o[509]) );
  AND U10892 ( .A(p_input[20509]), .B(p_input[10509]), .Z(n5446) );
  AND U10893 ( .A(n5447), .B(p_input[5099]), .Z(o[5099]) );
  AND U10894 ( .A(p_input[25099]), .B(p_input[15099]), .Z(n5447) );
  AND U10895 ( .A(n5448), .B(p_input[5098]), .Z(o[5098]) );
  AND U10896 ( .A(p_input[25098]), .B(p_input[15098]), .Z(n5448) );
  AND U10897 ( .A(n5449), .B(p_input[5097]), .Z(o[5097]) );
  AND U10898 ( .A(p_input[25097]), .B(p_input[15097]), .Z(n5449) );
  AND U10899 ( .A(n5450), .B(p_input[5096]), .Z(o[5096]) );
  AND U10900 ( .A(p_input[25096]), .B(p_input[15096]), .Z(n5450) );
  AND U10901 ( .A(n5451), .B(p_input[5095]), .Z(o[5095]) );
  AND U10902 ( .A(p_input[25095]), .B(p_input[15095]), .Z(n5451) );
  AND U10903 ( .A(n5452), .B(p_input[5094]), .Z(o[5094]) );
  AND U10904 ( .A(p_input[25094]), .B(p_input[15094]), .Z(n5452) );
  AND U10905 ( .A(n5453), .B(p_input[5093]), .Z(o[5093]) );
  AND U10906 ( .A(p_input[25093]), .B(p_input[15093]), .Z(n5453) );
  AND U10907 ( .A(n5454), .B(p_input[5092]), .Z(o[5092]) );
  AND U10908 ( .A(p_input[25092]), .B(p_input[15092]), .Z(n5454) );
  AND U10909 ( .A(n5455), .B(p_input[5091]), .Z(o[5091]) );
  AND U10910 ( .A(p_input[25091]), .B(p_input[15091]), .Z(n5455) );
  AND U10911 ( .A(n5456), .B(p_input[5090]), .Z(o[5090]) );
  AND U10912 ( .A(p_input[25090]), .B(p_input[15090]), .Z(n5456) );
  AND U10913 ( .A(n5457), .B(p_input[508]), .Z(o[508]) );
  AND U10914 ( .A(p_input[20508]), .B(p_input[10508]), .Z(n5457) );
  AND U10915 ( .A(n5458), .B(p_input[5089]), .Z(o[5089]) );
  AND U10916 ( .A(p_input[25089]), .B(p_input[15089]), .Z(n5458) );
  AND U10917 ( .A(n5459), .B(p_input[5088]), .Z(o[5088]) );
  AND U10918 ( .A(p_input[25088]), .B(p_input[15088]), .Z(n5459) );
  AND U10919 ( .A(n5460), .B(p_input[5087]), .Z(o[5087]) );
  AND U10920 ( .A(p_input[25087]), .B(p_input[15087]), .Z(n5460) );
  AND U10921 ( .A(n5461), .B(p_input[5086]), .Z(o[5086]) );
  AND U10922 ( .A(p_input[25086]), .B(p_input[15086]), .Z(n5461) );
  AND U10923 ( .A(n5462), .B(p_input[5085]), .Z(o[5085]) );
  AND U10924 ( .A(p_input[25085]), .B(p_input[15085]), .Z(n5462) );
  AND U10925 ( .A(n5463), .B(p_input[5084]), .Z(o[5084]) );
  AND U10926 ( .A(p_input[25084]), .B(p_input[15084]), .Z(n5463) );
  AND U10927 ( .A(n5464), .B(p_input[5083]), .Z(o[5083]) );
  AND U10928 ( .A(p_input[25083]), .B(p_input[15083]), .Z(n5464) );
  AND U10929 ( .A(n5465), .B(p_input[5082]), .Z(o[5082]) );
  AND U10930 ( .A(p_input[25082]), .B(p_input[15082]), .Z(n5465) );
  AND U10931 ( .A(n5466), .B(p_input[5081]), .Z(o[5081]) );
  AND U10932 ( .A(p_input[25081]), .B(p_input[15081]), .Z(n5466) );
  AND U10933 ( .A(n5467), .B(p_input[5080]), .Z(o[5080]) );
  AND U10934 ( .A(p_input[25080]), .B(p_input[15080]), .Z(n5467) );
  AND U10935 ( .A(n5468), .B(p_input[507]), .Z(o[507]) );
  AND U10936 ( .A(p_input[20507]), .B(p_input[10507]), .Z(n5468) );
  AND U10937 ( .A(n5469), .B(p_input[5079]), .Z(o[5079]) );
  AND U10938 ( .A(p_input[25079]), .B(p_input[15079]), .Z(n5469) );
  AND U10939 ( .A(n5470), .B(p_input[5078]), .Z(o[5078]) );
  AND U10940 ( .A(p_input[25078]), .B(p_input[15078]), .Z(n5470) );
  AND U10941 ( .A(n5471), .B(p_input[5077]), .Z(o[5077]) );
  AND U10942 ( .A(p_input[25077]), .B(p_input[15077]), .Z(n5471) );
  AND U10943 ( .A(n5472), .B(p_input[5076]), .Z(o[5076]) );
  AND U10944 ( .A(p_input[25076]), .B(p_input[15076]), .Z(n5472) );
  AND U10945 ( .A(n5473), .B(p_input[5075]), .Z(o[5075]) );
  AND U10946 ( .A(p_input[25075]), .B(p_input[15075]), .Z(n5473) );
  AND U10947 ( .A(n5474), .B(p_input[5074]), .Z(o[5074]) );
  AND U10948 ( .A(p_input[25074]), .B(p_input[15074]), .Z(n5474) );
  AND U10949 ( .A(n5475), .B(p_input[5073]), .Z(o[5073]) );
  AND U10950 ( .A(p_input[25073]), .B(p_input[15073]), .Z(n5475) );
  AND U10951 ( .A(n5476), .B(p_input[5072]), .Z(o[5072]) );
  AND U10952 ( .A(p_input[25072]), .B(p_input[15072]), .Z(n5476) );
  AND U10953 ( .A(n5477), .B(p_input[5071]), .Z(o[5071]) );
  AND U10954 ( .A(p_input[25071]), .B(p_input[15071]), .Z(n5477) );
  AND U10955 ( .A(n5478), .B(p_input[5070]), .Z(o[5070]) );
  AND U10956 ( .A(p_input[25070]), .B(p_input[15070]), .Z(n5478) );
  AND U10957 ( .A(n5479), .B(p_input[506]), .Z(o[506]) );
  AND U10958 ( .A(p_input[20506]), .B(p_input[10506]), .Z(n5479) );
  AND U10959 ( .A(n5480), .B(p_input[5069]), .Z(o[5069]) );
  AND U10960 ( .A(p_input[25069]), .B(p_input[15069]), .Z(n5480) );
  AND U10961 ( .A(n5481), .B(p_input[5068]), .Z(o[5068]) );
  AND U10962 ( .A(p_input[25068]), .B(p_input[15068]), .Z(n5481) );
  AND U10963 ( .A(n5482), .B(p_input[5067]), .Z(o[5067]) );
  AND U10964 ( .A(p_input[25067]), .B(p_input[15067]), .Z(n5482) );
  AND U10965 ( .A(n5483), .B(p_input[5066]), .Z(o[5066]) );
  AND U10966 ( .A(p_input[25066]), .B(p_input[15066]), .Z(n5483) );
  AND U10967 ( .A(n5484), .B(p_input[5065]), .Z(o[5065]) );
  AND U10968 ( .A(p_input[25065]), .B(p_input[15065]), .Z(n5484) );
  AND U10969 ( .A(n5485), .B(p_input[5064]), .Z(o[5064]) );
  AND U10970 ( .A(p_input[25064]), .B(p_input[15064]), .Z(n5485) );
  AND U10971 ( .A(n5486), .B(p_input[5063]), .Z(o[5063]) );
  AND U10972 ( .A(p_input[25063]), .B(p_input[15063]), .Z(n5486) );
  AND U10973 ( .A(n5487), .B(p_input[5062]), .Z(o[5062]) );
  AND U10974 ( .A(p_input[25062]), .B(p_input[15062]), .Z(n5487) );
  AND U10975 ( .A(n5488), .B(p_input[5061]), .Z(o[5061]) );
  AND U10976 ( .A(p_input[25061]), .B(p_input[15061]), .Z(n5488) );
  AND U10977 ( .A(n5489), .B(p_input[5060]), .Z(o[5060]) );
  AND U10978 ( .A(p_input[25060]), .B(p_input[15060]), .Z(n5489) );
  AND U10979 ( .A(n5490), .B(p_input[505]), .Z(o[505]) );
  AND U10980 ( .A(p_input[20505]), .B(p_input[10505]), .Z(n5490) );
  AND U10981 ( .A(n5491), .B(p_input[5059]), .Z(o[5059]) );
  AND U10982 ( .A(p_input[25059]), .B(p_input[15059]), .Z(n5491) );
  AND U10983 ( .A(n5492), .B(p_input[5058]), .Z(o[5058]) );
  AND U10984 ( .A(p_input[25058]), .B(p_input[15058]), .Z(n5492) );
  AND U10985 ( .A(n5493), .B(p_input[5057]), .Z(o[5057]) );
  AND U10986 ( .A(p_input[25057]), .B(p_input[15057]), .Z(n5493) );
  AND U10987 ( .A(n5494), .B(p_input[5056]), .Z(o[5056]) );
  AND U10988 ( .A(p_input[25056]), .B(p_input[15056]), .Z(n5494) );
  AND U10989 ( .A(n5495), .B(p_input[5055]), .Z(o[5055]) );
  AND U10990 ( .A(p_input[25055]), .B(p_input[15055]), .Z(n5495) );
  AND U10991 ( .A(n5496), .B(p_input[5054]), .Z(o[5054]) );
  AND U10992 ( .A(p_input[25054]), .B(p_input[15054]), .Z(n5496) );
  AND U10993 ( .A(n5497), .B(p_input[5053]), .Z(o[5053]) );
  AND U10994 ( .A(p_input[25053]), .B(p_input[15053]), .Z(n5497) );
  AND U10995 ( .A(n5498), .B(p_input[5052]), .Z(o[5052]) );
  AND U10996 ( .A(p_input[25052]), .B(p_input[15052]), .Z(n5498) );
  AND U10997 ( .A(n5499), .B(p_input[5051]), .Z(o[5051]) );
  AND U10998 ( .A(p_input[25051]), .B(p_input[15051]), .Z(n5499) );
  AND U10999 ( .A(n5500), .B(p_input[5050]), .Z(o[5050]) );
  AND U11000 ( .A(p_input[25050]), .B(p_input[15050]), .Z(n5500) );
  AND U11001 ( .A(n5501), .B(p_input[504]), .Z(o[504]) );
  AND U11002 ( .A(p_input[20504]), .B(p_input[10504]), .Z(n5501) );
  AND U11003 ( .A(n5502), .B(p_input[5049]), .Z(o[5049]) );
  AND U11004 ( .A(p_input[25049]), .B(p_input[15049]), .Z(n5502) );
  AND U11005 ( .A(n5503), .B(p_input[5048]), .Z(o[5048]) );
  AND U11006 ( .A(p_input[25048]), .B(p_input[15048]), .Z(n5503) );
  AND U11007 ( .A(n5504), .B(p_input[5047]), .Z(o[5047]) );
  AND U11008 ( .A(p_input[25047]), .B(p_input[15047]), .Z(n5504) );
  AND U11009 ( .A(n5505), .B(p_input[5046]), .Z(o[5046]) );
  AND U11010 ( .A(p_input[25046]), .B(p_input[15046]), .Z(n5505) );
  AND U11011 ( .A(n5506), .B(p_input[5045]), .Z(o[5045]) );
  AND U11012 ( .A(p_input[25045]), .B(p_input[15045]), .Z(n5506) );
  AND U11013 ( .A(n5507), .B(p_input[5044]), .Z(o[5044]) );
  AND U11014 ( .A(p_input[25044]), .B(p_input[15044]), .Z(n5507) );
  AND U11015 ( .A(n5508), .B(p_input[5043]), .Z(o[5043]) );
  AND U11016 ( .A(p_input[25043]), .B(p_input[15043]), .Z(n5508) );
  AND U11017 ( .A(n5509), .B(p_input[5042]), .Z(o[5042]) );
  AND U11018 ( .A(p_input[25042]), .B(p_input[15042]), .Z(n5509) );
  AND U11019 ( .A(n5510), .B(p_input[5041]), .Z(o[5041]) );
  AND U11020 ( .A(p_input[25041]), .B(p_input[15041]), .Z(n5510) );
  AND U11021 ( .A(n5511), .B(p_input[5040]), .Z(o[5040]) );
  AND U11022 ( .A(p_input[25040]), .B(p_input[15040]), .Z(n5511) );
  AND U11023 ( .A(n5512), .B(p_input[503]), .Z(o[503]) );
  AND U11024 ( .A(p_input[20503]), .B(p_input[10503]), .Z(n5512) );
  AND U11025 ( .A(n5513), .B(p_input[5039]), .Z(o[5039]) );
  AND U11026 ( .A(p_input[25039]), .B(p_input[15039]), .Z(n5513) );
  AND U11027 ( .A(n5514), .B(p_input[5038]), .Z(o[5038]) );
  AND U11028 ( .A(p_input[25038]), .B(p_input[15038]), .Z(n5514) );
  AND U11029 ( .A(n5515), .B(p_input[5037]), .Z(o[5037]) );
  AND U11030 ( .A(p_input[25037]), .B(p_input[15037]), .Z(n5515) );
  AND U11031 ( .A(n5516), .B(p_input[5036]), .Z(o[5036]) );
  AND U11032 ( .A(p_input[25036]), .B(p_input[15036]), .Z(n5516) );
  AND U11033 ( .A(n5517), .B(p_input[5035]), .Z(o[5035]) );
  AND U11034 ( .A(p_input[25035]), .B(p_input[15035]), .Z(n5517) );
  AND U11035 ( .A(n5518), .B(p_input[5034]), .Z(o[5034]) );
  AND U11036 ( .A(p_input[25034]), .B(p_input[15034]), .Z(n5518) );
  AND U11037 ( .A(n5519), .B(p_input[5033]), .Z(o[5033]) );
  AND U11038 ( .A(p_input[25033]), .B(p_input[15033]), .Z(n5519) );
  AND U11039 ( .A(n5520), .B(p_input[5032]), .Z(o[5032]) );
  AND U11040 ( .A(p_input[25032]), .B(p_input[15032]), .Z(n5520) );
  AND U11041 ( .A(n5521), .B(p_input[5031]), .Z(o[5031]) );
  AND U11042 ( .A(p_input[25031]), .B(p_input[15031]), .Z(n5521) );
  AND U11043 ( .A(n5522), .B(p_input[5030]), .Z(o[5030]) );
  AND U11044 ( .A(p_input[25030]), .B(p_input[15030]), .Z(n5522) );
  AND U11045 ( .A(n5523), .B(p_input[502]), .Z(o[502]) );
  AND U11046 ( .A(p_input[20502]), .B(p_input[10502]), .Z(n5523) );
  AND U11047 ( .A(n5524), .B(p_input[5029]), .Z(o[5029]) );
  AND U11048 ( .A(p_input[25029]), .B(p_input[15029]), .Z(n5524) );
  AND U11049 ( .A(n5525), .B(p_input[5028]), .Z(o[5028]) );
  AND U11050 ( .A(p_input[25028]), .B(p_input[15028]), .Z(n5525) );
  AND U11051 ( .A(n5526), .B(p_input[5027]), .Z(o[5027]) );
  AND U11052 ( .A(p_input[25027]), .B(p_input[15027]), .Z(n5526) );
  AND U11053 ( .A(n5527), .B(p_input[5026]), .Z(o[5026]) );
  AND U11054 ( .A(p_input[25026]), .B(p_input[15026]), .Z(n5527) );
  AND U11055 ( .A(n5528), .B(p_input[5025]), .Z(o[5025]) );
  AND U11056 ( .A(p_input[25025]), .B(p_input[15025]), .Z(n5528) );
  AND U11057 ( .A(n5529), .B(p_input[5024]), .Z(o[5024]) );
  AND U11058 ( .A(p_input[25024]), .B(p_input[15024]), .Z(n5529) );
  AND U11059 ( .A(n5530), .B(p_input[5023]), .Z(o[5023]) );
  AND U11060 ( .A(p_input[25023]), .B(p_input[15023]), .Z(n5530) );
  AND U11061 ( .A(n5531), .B(p_input[5022]), .Z(o[5022]) );
  AND U11062 ( .A(p_input[25022]), .B(p_input[15022]), .Z(n5531) );
  AND U11063 ( .A(n5532), .B(p_input[5021]), .Z(o[5021]) );
  AND U11064 ( .A(p_input[25021]), .B(p_input[15021]), .Z(n5532) );
  AND U11065 ( .A(n5533), .B(p_input[5020]), .Z(o[5020]) );
  AND U11066 ( .A(p_input[25020]), .B(p_input[15020]), .Z(n5533) );
  AND U11067 ( .A(n5534), .B(p_input[501]), .Z(o[501]) );
  AND U11068 ( .A(p_input[20501]), .B(p_input[10501]), .Z(n5534) );
  AND U11069 ( .A(n5535), .B(p_input[5019]), .Z(o[5019]) );
  AND U11070 ( .A(p_input[25019]), .B(p_input[15019]), .Z(n5535) );
  AND U11071 ( .A(n5536), .B(p_input[5018]), .Z(o[5018]) );
  AND U11072 ( .A(p_input[25018]), .B(p_input[15018]), .Z(n5536) );
  AND U11073 ( .A(n5537), .B(p_input[5017]), .Z(o[5017]) );
  AND U11074 ( .A(p_input[25017]), .B(p_input[15017]), .Z(n5537) );
  AND U11075 ( .A(n5538), .B(p_input[5016]), .Z(o[5016]) );
  AND U11076 ( .A(p_input[25016]), .B(p_input[15016]), .Z(n5538) );
  AND U11077 ( .A(n5539), .B(p_input[5015]), .Z(o[5015]) );
  AND U11078 ( .A(p_input[25015]), .B(p_input[15015]), .Z(n5539) );
  AND U11079 ( .A(n5540), .B(p_input[5014]), .Z(o[5014]) );
  AND U11080 ( .A(p_input[25014]), .B(p_input[15014]), .Z(n5540) );
  AND U11081 ( .A(n5541), .B(p_input[5013]), .Z(o[5013]) );
  AND U11082 ( .A(p_input[25013]), .B(p_input[15013]), .Z(n5541) );
  AND U11083 ( .A(n5542), .B(p_input[5012]), .Z(o[5012]) );
  AND U11084 ( .A(p_input[25012]), .B(p_input[15012]), .Z(n5542) );
  AND U11085 ( .A(n5543), .B(p_input[5011]), .Z(o[5011]) );
  AND U11086 ( .A(p_input[25011]), .B(p_input[15011]), .Z(n5543) );
  AND U11087 ( .A(n5544), .B(p_input[5010]), .Z(o[5010]) );
  AND U11088 ( .A(p_input[25010]), .B(p_input[15010]), .Z(n5544) );
  AND U11089 ( .A(n5545), .B(p_input[500]), .Z(o[500]) );
  AND U11090 ( .A(p_input[20500]), .B(p_input[10500]), .Z(n5545) );
  AND U11091 ( .A(n5546), .B(p_input[5009]), .Z(o[5009]) );
  AND U11092 ( .A(p_input[25009]), .B(p_input[15009]), .Z(n5546) );
  AND U11093 ( .A(n5547), .B(p_input[5008]), .Z(o[5008]) );
  AND U11094 ( .A(p_input[25008]), .B(p_input[15008]), .Z(n5547) );
  AND U11095 ( .A(n5548), .B(p_input[5007]), .Z(o[5007]) );
  AND U11096 ( .A(p_input[25007]), .B(p_input[15007]), .Z(n5548) );
  AND U11097 ( .A(n5549), .B(p_input[5006]), .Z(o[5006]) );
  AND U11098 ( .A(p_input[25006]), .B(p_input[15006]), .Z(n5549) );
  AND U11099 ( .A(n5550), .B(p_input[5005]), .Z(o[5005]) );
  AND U11100 ( .A(p_input[25005]), .B(p_input[15005]), .Z(n5550) );
  AND U11101 ( .A(n5551), .B(p_input[5004]), .Z(o[5004]) );
  AND U11102 ( .A(p_input[25004]), .B(p_input[15004]), .Z(n5551) );
  AND U11103 ( .A(n5552), .B(p_input[5003]), .Z(o[5003]) );
  AND U11104 ( .A(p_input[25003]), .B(p_input[15003]), .Z(n5552) );
  AND U11105 ( .A(n5553), .B(p_input[5002]), .Z(o[5002]) );
  AND U11106 ( .A(p_input[25002]), .B(p_input[15002]), .Z(n5553) );
  AND U11107 ( .A(n5554), .B(p_input[5001]), .Z(o[5001]) );
  AND U11108 ( .A(p_input[25001]), .B(p_input[15001]), .Z(n5554) );
  AND U11109 ( .A(n5555), .B(p_input[5000]), .Z(o[5000]) );
  AND U11110 ( .A(p_input[25000]), .B(p_input[15000]), .Z(n5555) );
  AND U11111 ( .A(n5556), .B(p_input[4]), .Z(o[4]) );
  AND U11112 ( .A(p_input[20004]), .B(p_input[10004]), .Z(n5556) );
  AND U11113 ( .A(n5557), .B(p_input[49]), .Z(o[49]) );
  AND U11114 ( .A(p_input[20049]), .B(p_input[10049]), .Z(n5557) );
  AND U11115 ( .A(n5558), .B(p_input[499]), .Z(o[499]) );
  AND U11116 ( .A(p_input[20499]), .B(p_input[10499]), .Z(n5558) );
  AND U11117 ( .A(n5559), .B(p_input[4999]), .Z(o[4999]) );
  AND U11118 ( .A(p_input[24999]), .B(p_input[14999]), .Z(n5559) );
  AND U11119 ( .A(n5560), .B(p_input[4998]), .Z(o[4998]) );
  AND U11120 ( .A(p_input[24998]), .B(p_input[14998]), .Z(n5560) );
  AND U11121 ( .A(n5561), .B(p_input[4997]), .Z(o[4997]) );
  AND U11122 ( .A(p_input[24997]), .B(p_input[14997]), .Z(n5561) );
  AND U11123 ( .A(n5562), .B(p_input[4996]), .Z(o[4996]) );
  AND U11124 ( .A(p_input[24996]), .B(p_input[14996]), .Z(n5562) );
  AND U11125 ( .A(n5563), .B(p_input[4995]), .Z(o[4995]) );
  AND U11126 ( .A(p_input[24995]), .B(p_input[14995]), .Z(n5563) );
  AND U11127 ( .A(n5564), .B(p_input[4994]), .Z(o[4994]) );
  AND U11128 ( .A(p_input[24994]), .B(p_input[14994]), .Z(n5564) );
  AND U11129 ( .A(n5565), .B(p_input[4993]), .Z(o[4993]) );
  AND U11130 ( .A(p_input[24993]), .B(p_input[14993]), .Z(n5565) );
  AND U11131 ( .A(n5566), .B(p_input[4992]), .Z(o[4992]) );
  AND U11132 ( .A(p_input[24992]), .B(p_input[14992]), .Z(n5566) );
  AND U11133 ( .A(n5567), .B(p_input[4991]), .Z(o[4991]) );
  AND U11134 ( .A(p_input[24991]), .B(p_input[14991]), .Z(n5567) );
  AND U11135 ( .A(n5568), .B(p_input[4990]), .Z(o[4990]) );
  AND U11136 ( .A(p_input[24990]), .B(p_input[14990]), .Z(n5568) );
  AND U11137 ( .A(n5569), .B(p_input[498]), .Z(o[498]) );
  AND U11138 ( .A(p_input[20498]), .B(p_input[10498]), .Z(n5569) );
  AND U11139 ( .A(n5570), .B(p_input[4989]), .Z(o[4989]) );
  AND U11140 ( .A(p_input[24989]), .B(p_input[14989]), .Z(n5570) );
  AND U11141 ( .A(n5571), .B(p_input[4988]), .Z(o[4988]) );
  AND U11142 ( .A(p_input[24988]), .B(p_input[14988]), .Z(n5571) );
  AND U11143 ( .A(n5572), .B(p_input[4987]), .Z(o[4987]) );
  AND U11144 ( .A(p_input[24987]), .B(p_input[14987]), .Z(n5572) );
  AND U11145 ( .A(n5573), .B(p_input[4986]), .Z(o[4986]) );
  AND U11146 ( .A(p_input[24986]), .B(p_input[14986]), .Z(n5573) );
  AND U11147 ( .A(n5574), .B(p_input[4985]), .Z(o[4985]) );
  AND U11148 ( .A(p_input[24985]), .B(p_input[14985]), .Z(n5574) );
  AND U11149 ( .A(n5575), .B(p_input[4984]), .Z(o[4984]) );
  AND U11150 ( .A(p_input[24984]), .B(p_input[14984]), .Z(n5575) );
  AND U11151 ( .A(n5576), .B(p_input[4983]), .Z(o[4983]) );
  AND U11152 ( .A(p_input[24983]), .B(p_input[14983]), .Z(n5576) );
  AND U11153 ( .A(n5577), .B(p_input[4982]), .Z(o[4982]) );
  AND U11154 ( .A(p_input[24982]), .B(p_input[14982]), .Z(n5577) );
  AND U11155 ( .A(n5578), .B(p_input[4981]), .Z(o[4981]) );
  AND U11156 ( .A(p_input[24981]), .B(p_input[14981]), .Z(n5578) );
  AND U11157 ( .A(n5579), .B(p_input[4980]), .Z(o[4980]) );
  AND U11158 ( .A(p_input[24980]), .B(p_input[14980]), .Z(n5579) );
  AND U11159 ( .A(n5580), .B(p_input[497]), .Z(o[497]) );
  AND U11160 ( .A(p_input[20497]), .B(p_input[10497]), .Z(n5580) );
  AND U11161 ( .A(n5581), .B(p_input[4979]), .Z(o[4979]) );
  AND U11162 ( .A(p_input[24979]), .B(p_input[14979]), .Z(n5581) );
  AND U11163 ( .A(n5582), .B(p_input[4978]), .Z(o[4978]) );
  AND U11164 ( .A(p_input[24978]), .B(p_input[14978]), .Z(n5582) );
  AND U11165 ( .A(n5583), .B(p_input[4977]), .Z(o[4977]) );
  AND U11166 ( .A(p_input[24977]), .B(p_input[14977]), .Z(n5583) );
  AND U11167 ( .A(n5584), .B(p_input[4976]), .Z(o[4976]) );
  AND U11168 ( .A(p_input[24976]), .B(p_input[14976]), .Z(n5584) );
  AND U11169 ( .A(n5585), .B(p_input[4975]), .Z(o[4975]) );
  AND U11170 ( .A(p_input[24975]), .B(p_input[14975]), .Z(n5585) );
  AND U11171 ( .A(n5586), .B(p_input[4974]), .Z(o[4974]) );
  AND U11172 ( .A(p_input[24974]), .B(p_input[14974]), .Z(n5586) );
  AND U11173 ( .A(n5587), .B(p_input[4973]), .Z(o[4973]) );
  AND U11174 ( .A(p_input[24973]), .B(p_input[14973]), .Z(n5587) );
  AND U11175 ( .A(n5588), .B(p_input[4972]), .Z(o[4972]) );
  AND U11176 ( .A(p_input[24972]), .B(p_input[14972]), .Z(n5588) );
  AND U11177 ( .A(n5589), .B(p_input[4971]), .Z(o[4971]) );
  AND U11178 ( .A(p_input[24971]), .B(p_input[14971]), .Z(n5589) );
  AND U11179 ( .A(n5590), .B(p_input[4970]), .Z(o[4970]) );
  AND U11180 ( .A(p_input[24970]), .B(p_input[14970]), .Z(n5590) );
  AND U11181 ( .A(n5591), .B(p_input[496]), .Z(o[496]) );
  AND U11182 ( .A(p_input[20496]), .B(p_input[10496]), .Z(n5591) );
  AND U11183 ( .A(n5592), .B(p_input[4969]), .Z(o[4969]) );
  AND U11184 ( .A(p_input[24969]), .B(p_input[14969]), .Z(n5592) );
  AND U11185 ( .A(n5593), .B(p_input[4968]), .Z(o[4968]) );
  AND U11186 ( .A(p_input[24968]), .B(p_input[14968]), .Z(n5593) );
  AND U11187 ( .A(n5594), .B(p_input[4967]), .Z(o[4967]) );
  AND U11188 ( .A(p_input[24967]), .B(p_input[14967]), .Z(n5594) );
  AND U11189 ( .A(n5595), .B(p_input[4966]), .Z(o[4966]) );
  AND U11190 ( .A(p_input[24966]), .B(p_input[14966]), .Z(n5595) );
  AND U11191 ( .A(n5596), .B(p_input[4965]), .Z(o[4965]) );
  AND U11192 ( .A(p_input[24965]), .B(p_input[14965]), .Z(n5596) );
  AND U11193 ( .A(n5597), .B(p_input[4964]), .Z(o[4964]) );
  AND U11194 ( .A(p_input[24964]), .B(p_input[14964]), .Z(n5597) );
  AND U11195 ( .A(n5598), .B(p_input[4963]), .Z(o[4963]) );
  AND U11196 ( .A(p_input[24963]), .B(p_input[14963]), .Z(n5598) );
  AND U11197 ( .A(n5599), .B(p_input[4962]), .Z(o[4962]) );
  AND U11198 ( .A(p_input[24962]), .B(p_input[14962]), .Z(n5599) );
  AND U11199 ( .A(n5600), .B(p_input[4961]), .Z(o[4961]) );
  AND U11200 ( .A(p_input[24961]), .B(p_input[14961]), .Z(n5600) );
  AND U11201 ( .A(n5601), .B(p_input[4960]), .Z(o[4960]) );
  AND U11202 ( .A(p_input[24960]), .B(p_input[14960]), .Z(n5601) );
  AND U11203 ( .A(n5602), .B(p_input[495]), .Z(o[495]) );
  AND U11204 ( .A(p_input[20495]), .B(p_input[10495]), .Z(n5602) );
  AND U11205 ( .A(n5603), .B(p_input[4959]), .Z(o[4959]) );
  AND U11206 ( .A(p_input[24959]), .B(p_input[14959]), .Z(n5603) );
  AND U11207 ( .A(n5604), .B(p_input[4958]), .Z(o[4958]) );
  AND U11208 ( .A(p_input[24958]), .B(p_input[14958]), .Z(n5604) );
  AND U11209 ( .A(n5605), .B(p_input[4957]), .Z(o[4957]) );
  AND U11210 ( .A(p_input[24957]), .B(p_input[14957]), .Z(n5605) );
  AND U11211 ( .A(n5606), .B(p_input[4956]), .Z(o[4956]) );
  AND U11212 ( .A(p_input[24956]), .B(p_input[14956]), .Z(n5606) );
  AND U11213 ( .A(n5607), .B(p_input[4955]), .Z(o[4955]) );
  AND U11214 ( .A(p_input[24955]), .B(p_input[14955]), .Z(n5607) );
  AND U11215 ( .A(n5608), .B(p_input[4954]), .Z(o[4954]) );
  AND U11216 ( .A(p_input[24954]), .B(p_input[14954]), .Z(n5608) );
  AND U11217 ( .A(n5609), .B(p_input[4953]), .Z(o[4953]) );
  AND U11218 ( .A(p_input[24953]), .B(p_input[14953]), .Z(n5609) );
  AND U11219 ( .A(n5610), .B(p_input[4952]), .Z(o[4952]) );
  AND U11220 ( .A(p_input[24952]), .B(p_input[14952]), .Z(n5610) );
  AND U11221 ( .A(n5611), .B(p_input[4951]), .Z(o[4951]) );
  AND U11222 ( .A(p_input[24951]), .B(p_input[14951]), .Z(n5611) );
  AND U11223 ( .A(n5612), .B(p_input[4950]), .Z(o[4950]) );
  AND U11224 ( .A(p_input[24950]), .B(p_input[14950]), .Z(n5612) );
  AND U11225 ( .A(n5613), .B(p_input[494]), .Z(o[494]) );
  AND U11226 ( .A(p_input[20494]), .B(p_input[10494]), .Z(n5613) );
  AND U11227 ( .A(n5614), .B(p_input[4949]), .Z(o[4949]) );
  AND U11228 ( .A(p_input[24949]), .B(p_input[14949]), .Z(n5614) );
  AND U11229 ( .A(n5615), .B(p_input[4948]), .Z(o[4948]) );
  AND U11230 ( .A(p_input[24948]), .B(p_input[14948]), .Z(n5615) );
  AND U11231 ( .A(n5616), .B(p_input[4947]), .Z(o[4947]) );
  AND U11232 ( .A(p_input[24947]), .B(p_input[14947]), .Z(n5616) );
  AND U11233 ( .A(n5617), .B(p_input[4946]), .Z(o[4946]) );
  AND U11234 ( .A(p_input[24946]), .B(p_input[14946]), .Z(n5617) );
  AND U11235 ( .A(n5618), .B(p_input[4945]), .Z(o[4945]) );
  AND U11236 ( .A(p_input[24945]), .B(p_input[14945]), .Z(n5618) );
  AND U11237 ( .A(n5619), .B(p_input[4944]), .Z(o[4944]) );
  AND U11238 ( .A(p_input[24944]), .B(p_input[14944]), .Z(n5619) );
  AND U11239 ( .A(n5620), .B(p_input[4943]), .Z(o[4943]) );
  AND U11240 ( .A(p_input[24943]), .B(p_input[14943]), .Z(n5620) );
  AND U11241 ( .A(n5621), .B(p_input[4942]), .Z(o[4942]) );
  AND U11242 ( .A(p_input[24942]), .B(p_input[14942]), .Z(n5621) );
  AND U11243 ( .A(n5622), .B(p_input[4941]), .Z(o[4941]) );
  AND U11244 ( .A(p_input[24941]), .B(p_input[14941]), .Z(n5622) );
  AND U11245 ( .A(n5623), .B(p_input[4940]), .Z(o[4940]) );
  AND U11246 ( .A(p_input[24940]), .B(p_input[14940]), .Z(n5623) );
  AND U11247 ( .A(n5624), .B(p_input[493]), .Z(o[493]) );
  AND U11248 ( .A(p_input[20493]), .B(p_input[10493]), .Z(n5624) );
  AND U11249 ( .A(n5625), .B(p_input[4939]), .Z(o[4939]) );
  AND U11250 ( .A(p_input[24939]), .B(p_input[14939]), .Z(n5625) );
  AND U11251 ( .A(n5626), .B(p_input[4938]), .Z(o[4938]) );
  AND U11252 ( .A(p_input[24938]), .B(p_input[14938]), .Z(n5626) );
  AND U11253 ( .A(n5627), .B(p_input[4937]), .Z(o[4937]) );
  AND U11254 ( .A(p_input[24937]), .B(p_input[14937]), .Z(n5627) );
  AND U11255 ( .A(n5628), .B(p_input[4936]), .Z(o[4936]) );
  AND U11256 ( .A(p_input[24936]), .B(p_input[14936]), .Z(n5628) );
  AND U11257 ( .A(n5629), .B(p_input[4935]), .Z(o[4935]) );
  AND U11258 ( .A(p_input[24935]), .B(p_input[14935]), .Z(n5629) );
  AND U11259 ( .A(n5630), .B(p_input[4934]), .Z(o[4934]) );
  AND U11260 ( .A(p_input[24934]), .B(p_input[14934]), .Z(n5630) );
  AND U11261 ( .A(n5631), .B(p_input[4933]), .Z(o[4933]) );
  AND U11262 ( .A(p_input[24933]), .B(p_input[14933]), .Z(n5631) );
  AND U11263 ( .A(n5632), .B(p_input[4932]), .Z(o[4932]) );
  AND U11264 ( .A(p_input[24932]), .B(p_input[14932]), .Z(n5632) );
  AND U11265 ( .A(n5633), .B(p_input[4931]), .Z(o[4931]) );
  AND U11266 ( .A(p_input[24931]), .B(p_input[14931]), .Z(n5633) );
  AND U11267 ( .A(n5634), .B(p_input[4930]), .Z(o[4930]) );
  AND U11268 ( .A(p_input[24930]), .B(p_input[14930]), .Z(n5634) );
  AND U11269 ( .A(n5635), .B(p_input[492]), .Z(o[492]) );
  AND U11270 ( .A(p_input[20492]), .B(p_input[10492]), .Z(n5635) );
  AND U11271 ( .A(n5636), .B(p_input[4929]), .Z(o[4929]) );
  AND U11272 ( .A(p_input[24929]), .B(p_input[14929]), .Z(n5636) );
  AND U11273 ( .A(n5637), .B(p_input[4928]), .Z(o[4928]) );
  AND U11274 ( .A(p_input[24928]), .B(p_input[14928]), .Z(n5637) );
  AND U11275 ( .A(n5638), .B(p_input[4927]), .Z(o[4927]) );
  AND U11276 ( .A(p_input[24927]), .B(p_input[14927]), .Z(n5638) );
  AND U11277 ( .A(n5639), .B(p_input[4926]), .Z(o[4926]) );
  AND U11278 ( .A(p_input[24926]), .B(p_input[14926]), .Z(n5639) );
  AND U11279 ( .A(n5640), .B(p_input[4925]), .Z(o[4925]) );
  AND U11280 ( .A(p_input[24925]), .B(p_input[14925]), .Z(n5640) );
  AND U11281 ( .A(n5641), .B(p_input[4924]), .Z(o[4924]) );
  AND U11282 ( .A(p_input[24924]), .B(p_input[14924]), .Z(n5641) );
  AND U11283 ( .A(n5642), .B(p_input[4923]), .Z(o[4923]) );
  AND U11284 ( .A(p_input[24923]), .B(p_input[14923]), .Z(n5642) );
  AND U11285 ( .A(n5643), .B(p_input[4922]), .Z(o[4922]) );
  AND U11286 ( .A(p_input[24922]), .B(p_input[14922]), .Z(n5643) );
  AND U11287 ( .A(n5644), .B(p_input[4921]), .Z(o[4921]) );
  AND U11288 ( .A(p_input[24921]), .B(p_input[14921]), .Z(n5644) );
  AND U11289 ( .A(n5645), .B(p_input[4920]), .Z(o[4920]) );
  AND U11290 ( .A(p_input[24920]), .B(p_input[14920]), .Z(n5645) );
  AND U11291 ( .A(n5646), .B(p_input[491]), .Z(o[491]) );
  AND U11292 ( .A(p_input[20491]), .B(p_input[10491]), .Z(n5646) );
  AND U11293 ( .A(n5647), .B(p_input[4919]), .Z(o[4919]) );
  AND U11294 ( .A(p_input[24919]), .B(p_input[14919]), .Z(n5647) );
  AND U11295 ( .A(n5648), .B(p_input[4918]), .Z(o[4918]) );
  AND U11296 ( .A(p_input[24918]), .B(p_input[14918]), .Z(n5648) );
  AND U11297 ( .A(n5649), .B(p_input[4917]), .Z(o[4917]) );
  AND U11298 ( .A(p_input[24917]), .B(p_input[14917]), .Z(n5649) );
  AND U11299 ( .A(n5650), .B(p_input[4916]), .Z(o[4916]) );
  AND U11300 ( .A(p_input[24916]), .B(p_input[14916]), .Z(n5650) );
  AND U11301 ( .A(n5651), .B(p_input[4915]), .Z(o[4915]) );
  AND U11302 ( .A(p_input[24915]), .B(p_input[14915]), .Z(n5651) );
  AND U11303 ( .A(n5652), .B(p_input[4914]), .Z(o[4914]) );
  AND U11304 ( .A(p_input[24914]), .B(p_input[14914]), .Z(n5652) );
  AND U11305 ( .A(n5653), .B(p_input[4913]), .Z(o[4913]) );
  AND U11306 ( .A(p_input[24913]), .B(p_input[14913]), .Z(n5653) );
  AND U11307 ( .A(n5654), .B(p_input[4912]), .Z(o[4912]) );
  AND U11308 ( .A(p_input[24912]), .B(p_input[14912]), .Z(n5654) );
  AND U11309 ( .A(n5655), .B(p_input[4911]), .Z(o[4911]) );
  AND U11310 ( .A(p_input[24911]), .B(p_input[14911]), .Z(n5655) );
  AND U11311 ( .A(n5656), .B(p_input[4910]), .Z(o[4910]) );
  AND U11312 ( .A(p_input[24910]), .B(p_input[14910]), .Z(n5656) );
  AND U11313 ( .A(n5657), .B(p_input[490]), .Z(o[490]) );
  AND U11314 ( .A(p_input[20490]), .B(p_input[10490]), .Z(n5657) );
  AND U11315 ( .A(n5658), .B(p_input[4909]), .Z(o[4909]) );
  AND U11316 ( .A(p_input[24909]), .B(p_input[14909]), .Z(n5658) );
  AND U11317 ( .A(n5659), .B(p_input[4908]), .Z(o[4908]) );
  AND U11318 ( .A(p_input[24908]), .B(p_input[14908]), .Z(n5659) );
  AND U11319 ( .A(n5660), .B(p_input[4907]), .Z(o[4907]) );
  AND U11320 ( .A(p_input[24907]), .B(p_input[14907]), .Z(n5660) );
  AND U11321 ( .A(n5661), .B(p_input[4906]), .Z(o[4906]) );
  AND U11322 ( .A(p_input[24906]), .B(p_input[14906]), .Z(n5661) );
  AND U11323 ( .A(n5662), .B(p_input[4905]), .Z(o[4905]) );
  AND U11324 ( .A(p_input[24905]), .B(p_input[14905]), .Z(n5662) );
  AND U11325 ( .A(n5663), .B(p_input[4904]), .Z(o[4904]) );
  AND U11326 ( .A(p_input[24904]), .B(p_input[14904]), .Z(n5663) );
  AND U11327 ( .A(n5664), .B(p_input[4903]), .Z(o[4903]) );
  AND U11328 ( .A(p_input[24903]), .B(p_input[14903]), .Z(n5664) );
  AND U11329 ( .A(n5665), .B(p_input[4902]), .Z(o[4902]) );
  AND U11330 ( .A(p_input[24902]), .B(p_input[14902]), .Z(n5665) );
  AND U11331 ( .A(n5666), .B(p_input[4901]), .Z(o[4901]) );
  AND U11332 ( .A(p_input[24901]), .B(p_input[14901]), .Z(n5666) );
  AND U11333 ( .A(n5667), .B(p_input[4900]), .Z(o[4900]) );
  AND U11334 ( .A(p_input[24900]), .B(p_input[14900]), .Z(n5667) );
  AND U11335 ( .A(n5668), .B(p_input[48]), .Z(o[48]) );
  AND U11336 ( .A(p_input[20048]), .B(p_input[10048]), .Z(n5668) );
  AND U11337 ( .A(n5669), .B(p_input[489]), .Z(o[489]) );
  AND U11338 ( .A(p_input[20489]), .B(p_input[10489]), .Z(n5669) );
  AND U11339 ( .A(n5670), .B(p_input[4899]), .Z(o[4899]) );
  AND U11340 ( .A(p_input[24899]), .B(p_input[14899]), .Z(n5670) );
  AND U11341 ( .A(n5671), .B(p_input[4898]), .Z(o[4898]) );
  AND U11342 ( .A(p_input[24898]), .B(p_input[14898]), .Z(n5671) );
  AND U11343 ( .A(n5672), .B(p_input[4897]), .Z(o[4897]) );
  AND U11344 ( .A(p_input[24897]), .B(p_input[14897]), .Z(n5672) );
  AND U11345 ( .A(n5673), .B(p_input[4896]), .Z(o[4896]) );
  AND U11346 ( .A(p_input[24896]), .B(p_input[14896]), .Z(n5673) );
  AND U11347 ( .A(n5674), .B(p_input[4895]), .Z(o[4895]) );
  AND U11348 ( .A(p_input[24895]), .B(p_input[14895]), .Z(n5674) );
  AND U11349 ( .A(n5675), .B(p_input[4894]), .Z(o[4894]) );
  AND U11350 ( .A(p_input[24894]), .B(p_input[14894]), .Z(n5675) );
  AND U11351 ( .A(n5676), .B(p_input[4893]), .Z(o[4893]) );
  AND U11352 ( .A(p_input[24893]), .B(p_input[14893]), .Z(n5676) );
  AND U11353 ( .A(n5677), .B(p_input[4892]), .Z(o[4892]) );
  AND U11354 ( .A(p_input[24892]), .B(p_input[14892]), .Z(n5677) );
  AND U11355 ( .A(n5678), .B(p_input[4891]), .Z(o[4891]) );
  AND U11356 ( .A(p_input[24891]), .B(p_input[14891]), .Z(n5678) );
  AND U11357 ( .A(n5679), .B(p_input[4890]), .Z(o[4890]) );
  AND U11358 ( .A(p_input[24890]), .B(p_input[14890]), .Z(n5679) );
  AND U11359 ( .A(n5680), .B(p_input[488]), .Z(o[488]) );
  AND U11360 ( .A(p_input[20488]), .B(p_input[10488]), .Z(n5680) );
  AND U11361 ( .A(n5681), .B(p_input[4889]), .Z(o[4889]) );
  AND U11362 ( .A(p_input[24889]), .B(p_input[14889]), .Z(n5681) );
  AND U11363 ( .A(n5682), .B(p_input[4888]), .Z(o[4888]) );
  AND U11364 ( .A(p_input[24888]), .B(p_input[14888]), .Z(n5682) );
  AND U11365 ( .A(n5683), .B(p_input[4887]), .Z(o[4887]) );
  AND U11366 ( .A(p_input[24887]), .B(p_input[14887]), .Z(n5683) );
  AND U11367 ( .A(n5684), .B(p_input[4886]), .Z(o[4886]) );
  AND U11368 ( .A(p_input[24886]), .B(p_input[14886]), .Z(n5684) );
  AND U11369 ( .A(n5685), .B(p_input[4885]), .Z(o[4885]) );
  AND U11370 ( .A(p_input[24885]), .B(p_input[14885]), .Z(n5685) );
  AND U11371 ( .A(n5686), .B(p_input[4884]), .Z(o[4884]) );
  AND U11372 ( .A(p_input[24884]), .B(p_input[14884]), .Z(n5686) );
  AND U11373 ( .A(n5687), .B(p_input[4883]), .Z(o[4883]) );
  AND U11374 ( .A(p_input[24883]), .B(p_input[14883]), .Z(n5687) );
  AND U11375 ( .A(n5688), .B(p_input[4882]), .Z(o[4882]) );
  AND U11376 ( .A(p_input[24882]), .B(p_input[14882]), .Z(n5688) );
  AND U11377 ( .A(n5689), .B(p_input[4881]), .Z(o[4881]) );
  AND U11378 ( .A(p_input[24881]), .B(p_input[14881]), .Z(n5689) );
  AND U11379 ( .A(n5690), .B(p_input[4880]), .Z(o[4880]) );
  AND U11380 ( .A(p_input[24880]), .B(p_input[14880]), .Z(n5690) );
  AND U11381 ( .A(n5691), .B(p_input[487]), .Z(o[487]) );
  AND U11382 ( .A(p_input[20487]), .B(p_input[10487]), .Z(n5691) );
  AND U11383 ( .A(n5692), .B(p_input[4879]), .Z(o[4879]) );
  AND U11384 ( .A(p_input[24879]), .B(p_input[14879]), .Z(n5692) );
  AND U11385 ( .A(n5693), .B(p_input[4878]), .Z(o[4878]) );
  AND U11386 ( .A(p_input[24878]), .B(p_input[14878]), .Z(n5693) );
  AND U11387 ( .A(n5694), .B(p_input[4877]), .Z(o[4877]) );
  AND U11388 ( .A(p_input[24877]), .B(p_input[14877]), .Z(n5694) );
  AND U11389 ( .A(n5695), .B(p_input[4876]), .Z(o[4876]) );
  AND U11390 ( .A(p_input[24876]), .B(p_input[14876]), .Z(n5695) );
  AND U11391 ( .A(n5696), .B(p_input[4875]), .Z(o[4875]) );
  AND U11392 ( .A(p_input[24875]), .B(p_input[14875]), .Z(n5696) );
  AND U11393 ( .A(n5697), .B(p_input[4874]), .Z(o[4874]) );
  AND U11394 ( .A(p_input[24874]), .B(p_input[14874]), .Z(n5697) );
  AND U11395 ( .A(n5698), .B(p_input[4873]), .Z(o[4873]) );
  AND U11396 ( .A(p_input[24873]), .B(p_input[14873]), .Z(n5698) );
  AND U11397 ( .A(n5699), .B(p_input[4872]), .Z(o[4872]) );
  AND U11398 ( .A(p_input[24872]), .B(p_input[14872]), .Z(n5699) );
  AND U11399 ( .A(n5700), .B(p_input[4871]), .Z(o[4871]) );
  AND U11400 ( .A(p_input[24871]), .B(p_input[14871]), .Z(n5700) );
  AND U11401 ( .A(n5701), .B(p_input[4870]), .Z(o[4870]) );
  AND U11402 ( .A(p_input[24870]), .B(p_input[14870]), .Z(n5701) );
  AND U11403 ( .A(n5702), .B(p_input[486]), .Z(o[486]) );
  AND U11404 ( .A(p_input[20486]), .B(p_input[10486]), .Z(n5702) );
  AND U11405 ( .A(n5703), .B(p_input[4869]), .Z(o[4869]) );
  AND U11406 ( .A(p_input[24869]), .B(p_input[14869]), .Z(n5703) );
  AND U11407 ( .A(n5704), .B(p_input[4868]), .Z(o[4868]) );
  AND U11408 ( .A(p_input[24868]), .B(p_input[14868]), .Z(n5704) );
  AND U11409 ( .A(n5705), .B(p_input[4867]), .Z(o[4867]) );
  AND U11410 ( .A(p_input[24867]), .B(p_input[14867]), .Z(n5705) );
  AND U11411 ( .A(n5706), .B(p_input[4866]), .Z(o[4866]) );
  AND U11412 ( .A(p_input[24866]), .B(p_input[14866]), .Z(n5706) );
  AND U11413 ( .A(n5707), .B(p_input[4865]), .Z(o[4865]) );
  AND U11414 ( .A(p_input[24865]), .B(p_input[14865]), .Z(n5707) );
  AND U11415 ( .A(n5708), .B(p_input[4864]), .Z(o[4864]) );
  AND U11416 ( .A(p_input[24864]), .B(p_input[14864]), .Z(n5708) );
  AND U11417 ( .A(n5709), .B(p_input[4863]), .Z(o[4863]) );
  AND U11418 ( .A(p_input[24863]), .B(p_input[14863]), .Z(n5709) );
  AND U11419 ( .A(n5710), .B(p_input[4862]), .Z(o[4862]) );
  AND U11420 ( .A(p_input[24862]), .B(p_input[14862]), .Z(n5710) );
  AND U11421 ( .A(n5711), .B(p_input[4861]), .Z(o[4861]) );
  AND U11422 ( .A(p_input[24861]), .B(p_input[14861]), .Z(n5711) );
  AND U11423 ( .A(n5712), .B(p_input[4860]), .Z(o[4860]) );
  AND U11424 ( .A(p_input[24860]), .B(p_input[14860]), .Z(n5712) );
  AND U11425 ( .A(n5713), .B(p_input[485]), .Z(o[485]) );
  AND U11426 ( .A(p_input[20485]), .B(p_input[10485]), .Z(n5713) );
  AND U11427 ( .A(n5714), .B(p_input[4859]), .Z(o[4859]) );
  AND U11428 ( .A(p_input[24859]), .B(p_input[14859]), .Z(n5714) );
  AND U11429 ( .A(n5715), .B(p_input[4858]), .Z(o[4858]) );
  AND U11430 ( .A(p_input[24858]), .B(p_input[14858]), .Z(n5715) );
  AND U11431 ( .A(n5716), .B(p_input[4857]), .Z(o[4857]) );
  AND U11432 ( .A(p_input[24857]), .B(p_input[14857]), .Z(n5716) );
  AND U11433 ( .A(n5717), .B(p_input[4856]), .Z(o[4856]) );
  AND U11434 ( .A(p_input[24856]), .B(p_input[14856]), .Z(n5717) );
  AND U11435 ( .A(n5718), .B(p_input[4855]), .Z(o[4855]) );
  AND U11436 ( .A(p_input[24855]), .B(p_input[14855]), .Z(n5718) );
  AND U11437 ( .A(n5719), .B(p_input[4854]), .Z(o[4854]) );
  AND U11438 ( .A(p_input[24854]), .B(p_input[14854]), .Z(n5719) );
  AND U11439 ( .A(n5720), .B(p_input[4853]), .Z(o[4853]) );
  AND U11440 ( .A(p_input[24853]), .B(p_input[14853]), .Z(n5720) );
  AND U11441 ( .A(n5721), .B(p_input[4852]), .Z(o[4852]) );
  AND U11442 ( .A(p_input[24852]), .B(p_input[14852]), .Z(n5721) );
  AND U11443 ( .A(n5722), .B(p_input[4851]), .Z(o[4851]) );
  AND U11444 ( .A(p_input[24851]), .B(p_input[14851]), .Z(n5722) );
  AND U11445 ( .A(n5723), .B(p_input[4850]), .Z(o[4850]) );
  AND U11446 ( .A(p_input[24850]), .B(p_input[14850]), .Z(n5723) );
  AND U11447 ( .A(n5724), .B(p_input[484]), .Z(o[484]) );
  AND U11448 ( .A(p_input[20484]), .B(p_input[10484]), .Z(n5724) );
  AND U11449 ( .A(n5725), .B(p_input[4849]), .Z(o[4849]) );
  AND U11450 ( .A(p_input[24849]), .B(p_input[14849]), .Z(n5725) );
  AND U11451 ( .A(n5726), .B(p_input[4848]), .Z(o[4848]) );
  AND U11452 ( .A(p_input[24848]), .B(p_input[14848]), .Z(n5726) );
  AND U11453 ( .A(n5727), .B(p_input[4847]), .Z(o[4847]) );
  AND U11454 ( .A(p_input[24847]), .B(p_input[14847]), .Z(n5727) );
  AND U11455 ( .A(n5728), .B(p_input[4846]), .Z(o[4846]) );
  AND U11456 ( .A(p_input[24846]), .B(p_input[14846]), .Z(n5728) );
  AND U11457 ( .A(n5729), .B(p_input[4845]), .Z(o[4845]) );
  AND U11458 ( .A(p_input[24845]), .B(p_input[14845]), .Z(n5729) );
  AND U11459 ( .A(n5730), .B(p_input[4844]), .Z(o[4844]) );
  AND U11460 ( .A(p_input[24844]), .B(p_input[14844]), .Z(n5730) );
  AND U11461 ( .A(n5731), .B(p_input[4843]), .Z(o[4843]) );
  AND U11462 ( .A(p_input[24843]), .B(p_input[14843]), .Z(n5731) );
  AND U11463 ( .A(n5732), .B(p_input[4842]), .Z(o[4842]) );
  AND U11464 ( .A(p_input[24842]), .B(p_input[14842]), .Z(n5732) );
  AND U11465 ( .A(n5733), .B(p_input[4841]), .Z(o[4841]) );
  AND U11466 ( .A(p_input[24841]), .B(p_input[14841]), .Z(n5733) );
  AND U11467 ( .A(n5734), .B(p_input[4840]), .Z(o[4840]) );
  AND U11468 ( .A(p_input[24840]), .B(p_input[14840]), .Z(n5734) );
  AND U11469 ( .A(n5735), .B(p_input[483]), .Z(o[483]) );
  AND U11470 ( .A(p_input[20483]), .B(p_input[10483]), .Z(n5735) );
  AND U11471 ( .A(n5736), .B(p_input[4839]), .Z(o[4839]) );
  AND U11472 ( .A(p_input[24839]), .B(p_input[14839]), .Z(n5736) );
  AND U11473 ( .A(n5737), .B(p_input[4838]), .Z(o[4838]) );
  AND U11474 ( .A(p_input[24838]), .B(p_input[14838]), .Z(n5737) );
  AND U11475 ( .A(n5738), .B(p_input[4837]), .Z(o[4837]) );
  AND U11476 ( .A(p_input[24837]), .B(p_input[14837]), .Z(n5738) );
  AND U11477 ( .A(n5739), .B(p_input[4836]), .Z(o[4836]) );
  AND U11478 ( .A(p_input[24836]), .B(p_input[14836]), .Z(n5739) );
  AND U11479 ( .A(n5740), .B(p_input[4835]), .Z(o[4835]) );
  AND U11480 ( .A(p_input[24835]), .B(p_input[14835]), .Z(n5740) );
  AND U11481 ( .A(n5741), .B(p_input[4834]), .Z(o[4834]) );
  AND U11482 ( .A(p_input[24834]), .B(p_input[14834]), .Z(n5741) );
  AND U11483 ( .A(n5742), .B(p_input[4833]), .Z(o[4833]) );
  AND U11484 ( .A(p_input[24833]), .B(p_input[14833]), .Z(n5742) );
  AND U11485 ( .A(n5743), .B(p_input[4832]), .Z(o[4832]) );
  AND U11486 ( .A(p_input[24832]), .B(p_input[14832]), .Z(n5743) );
  AND U11487 ( .A(n5744), .B(p_input[4831]), .Z(o[4831]) );
  AND U11488 ( .A(p_input[24831]), .B(p_input[14831]), .Z(n5744) );
  AND U11489 ( .A(n5745), .B(p_input[4830]), .Z(o[4830]) );
  AND U11490 ( .A(p_input[24830]), .B(p_input[14830]), .Z(n5745) );
  AND U11491 ( .A(n5746), .B(p_input[482]), .Z(o[482]) );
  AND U11492 ( .A(p_input[20482]), .B(p_input[10482]), .Z(n5746) );
  AND U11493 ( .A(n5747), .B(p_input[4829]), .Z(o[4829]) );
  AND U11494 ( .A(p_input[24829]), .B(p_input[14829]), .Z(n5747) );
  AND U11495 ( .A(n5748), .B(p_input[4828]), .Z(o[4828]) );
  AND U11496 ( .A(p_input[24828]), .B(p_input[14828]), .Z(n5748) );
  AND U11497 ( .A(n5749), .B(p_input[4827]), .Z(o[4827]) );
  AND U11498 ( .A(p_input[24827]), .B(p_input[14827]), .Z(n5749) );
  AND U11499 ( .A(n5750), .B(p_input[4826]), .Z(o[4826]) );
  AND U11500 ( .A(p_input[24826]), .B(p_input[14826]), .Z(n5750) );
  AND U11501 ( .A(n5751), .B(p_input[4825]), .Z(o[4825]) );
  AND U11502 ( .A(p_input[24825]), .B(p_input[14825]), .Z(n5751) );
  AND U11503 ( .A(n5752), .B(p_input[4824]), .Z(o[4824]) );
  AND U11504 ( .A(p_input[24824]), .B(p_input[14824]), .Z(n5752) );
  AND U11505 ( .A(n5753), .B(p_input[4823]), .Z(o[4823]) );
  AND U11506 ( .A(p_input[24823]), .B(p_input[14823]), .Z(n5753) );
  AND U11507 ( .A(n5754), .B(p_input[4822]), .Z(o[4822]) );
  AND U11508 ( .A(p_input[24822]), .B(p_input[14822]), .Z(n5754) );
  AND U11509 ( .A(n5755), .B(p_input[4821]), .Z(o[4821]) );
  AND U11510 ( .A(p_input[24821]), .B(p_input[14821]), .Z(n5755) );
  AND U11511 ( .A(n5756), .B(p_input[4820]), .Z(o[4820]) );
  AND U11512 ( .A(p_input[24820]), .B(p_input[14820]), .Z(n5756) );
  AND U11513 ( .A(n5757), .B(p_input[481]), .Z(o[481]) );
  AND U11514 ( .A(p_input[20481]), .B(p_input[10481]), .Z(n5757) );
  AND U11515 ( .A(n5758), .B(p_input[4819]), .Z(o[4819]) );
  AND U11516 ( .A(p_input[24819]), .B(p_input[14819]), .Z(n5758) );
  AND U11517 ( .A(n5759), .B(p_input[4818]), .Z(o[4818]) );
  AND U11518 ( .A(p_input[24818]), .B(p_input[14818]), .Z(n5759) );
  AND U11519 ( .A(n5760), .B(p_input[4817]), .Z(o[4817]) );
  AND U11520 ( .A(p_input[24817]), .B(p_input[14817]), .Z(n5760) );
  AND U11521 ( .A(n5761), .B(p_input[4816]), .Z(o[4816]) );
  AND U11522 ( .A(p_input[24816]), .B(p_input[14816]), .Z(n5761) );
  AND U11523 ( .A(n5762), .B(p_input[4815]), .Z(o[4815]) );
  AND U11524 ( .A(p_input[24815]), .B(p_input[14815]), .Z(n5762) );
  AND U11525 ( .A(n5763), .B(p_input[4814]), .Z(o[4814]) );
  AND U11526 ( .A(p_input[24814]), .B(p_input[14814]), .Z(n5763) );
  AND U11527 ( .A(n5764), .B(p_input[4813]), .Z(o[4813]) );
  AND U11528 ( .A(p_input[24813]), .B(p_input[14813]), .Z(n5764) );
  AND U11529 ( .A(n5765), .B(p_input[4812]), .Z(o[4812]) );
  AND U11530 ( .A(p_input[24812]), .B(p_input[14812]), .Z(n5765) );
  AND U11531 ( .A(n5766), .B(p_input[4811]), .Z(o[4811]) );
  AND U11532 ( .A(p_input[24811]), .B(p_input[14811]), .Z(n5766) );
  AND U11533 ( .A(n5767), .B(p_input[4810]), .Z(o[4810]) );
  AND U11534 ( .A(p_input[24810]), .B(p_input[14810]), .Z(n5767) );
  AND U11535 ( .A(n5768), .B(p_input[480]), .Z(o[480]) );
  AND U11536 ( .A(p_input[20480]), .B(p_input[10480]), .Z(n5768) );
  AND U11537 ( .A(n5769), .B(p_input[4809]), .Z(o[4809]) );
  AND U11538 ( .A(p_input[24809]), .B(p_input[14809]), .Z(n5769) );
  AND U11539 ( .A(n5770), .B(p_input[4808]), .Z(o[4808]) );
  AND U11540 ( .A(p_input[24808]), .B(p_input[14808]), .Z(n5770) );
  AND U11541 ( .A(n5771), .B(p_input[4807]), .Z(o[4807]) );
  AND U11542 ( .A(p_input[24807]), .B(p_input[14807]), .Z(n5771) );
  AND U11543 ( .A(n5772), .B(p_input[4806]), .Z(o[4806]) );
  AND U11544 ( .A(p_input[24806]), .B(p_input[14806]), .Z(n5772) );
  AND U11545 ( .A(n5773), .B(p_input[4805]), .Z(o[4805]) );
  AND U11546 ( .A(p_input[24805]), .B(p_input[14805]), .Z(n5773) );
  AND U11547 ( .A(n5774), .B(p_input[4804]), .Z(o[4804]) );
  AND U11548 ( .A(p_input[24804]), .B(p_input[14804]), .Z(n5774) );
  AND U11549 ( .A(n5775), .B(p_input[4803]), .Z(o[4803]) );
  AND U11550 ( .A(p_input[24803]), .B(p_input[14803]), .Z(n5775) );
  AND U11551 ( .A(n5776), .B(p_input[4802]), .Z(o[4802]) );
  AND U11552 ( .A(p_input[24802]), .B(p_input[14802]), .Z(n5776) );
  AND U11553 ( .A(n5777), .B(p_input[4801]), .Z(o[4801]) );
  AND U11554 ( .A(p_input[24801]), .B(p_input[14801]), .Z(n5777) );
  AND U11555 ( .A(n5778), .B(p_input[4800]), .Z(o[4800]) );
  AND U11556 ( .A(p_input[24800]), .B(p_input[14800]), .Z(n5778) );
  AND U11557 ( .A(n5779), .B(p_input[47]), .Z(o[47]) );
  AND U11558 ( .A(p_input[20047]), .B(p_input[10047]), .Z(n5779) );
  AND U11559 ( .A(n5780), .B(p_input[479]), .Z(o[479]) );
  AND U11560 ( .A(p_input[20479]), .B(p_input[10479]), .Z(n5780) );
  AND U11561 ( .A(n5781), .B(p_input[4799]), .Z(o[4799]) );
  AND U11562 ( .A(p_input[24799]), .B(p_input[14799]), .Z(n5781) );
  AND U11563 ( .A(n5782), .B(p_input[4798]), .Z(o[4798]) );
  AND U11564 ( .A(p_input[24798]), .B(p_input[14798]), .Z(n5782) );
  AND U11565 ( .A(n5783), .B(p_input[4797]), .Z(o[4797]) );
  AND U11566 ( .A(p_input[24797]), .B(p_input[14797]), .Z(n5783) );
  AND U11567 ( .A(n5784), .B(p_input[4796]), .Z(o[4796]) );
  AND U11568 ( .A(p_input[24796]), .B(p_input[14796]), .Z(n5784) );
  AND U11569 ( .A(n5785), .B(p_input[4795]), .Z(o[4795]) );
  AND U11570 ( .A(p_input[24795]), .B(p_input[14795]), .Z(n5785) );
  AND U11571 ( .A(n5786), .B(p_input[4794]), .Z(o[4794]) );
  AND U11572 ( .A(p_input[24794]), .B(p_input[14794]), .Z(n5786) );
  AND U11573 ( .A(n5787), .B(p_input[4793]), .Z(o[4793]) );
  AND U11574 ( .A(p_input[24793]), .B(p_input[14793]), .Z(n5787) );
  AND U11575 ( .A(n5788), .B(p_input[4792]), .Z(o[4792]) );
  AND U11576 ( .A(p_input[24792]), .B(p_input[14792]), .Z(n5788) );
  AND U11577 ( .A(n5789), .B(p_input[4791]), .Z(o[4791]) );
  AND U11578 ( .A(p_input[24791]), .B(p_input[14791]), .Z(n5789) );
  AND U11579 ( .A(n5790), .B(p_input[4790]), .Z(o[4790]) );
  AND U11580 ( .A(p_input[24790]), .B(p_input[14790]), .Z(n5790) );
  AND U11581 ( .A(n5791), .B(p_input[478]), .Z(o[478]) );
  AND U11582 ( .A(p_input[20478]), .B(p_input[10478]), .Z(n5791) );
  AND U11583 ( .A(n5792), .B(p_input[4789]), .Z(o[4789]) );
  AND U11584 ( .A(p_input[24789]), .B(p_input[14789]), .Z(n5792) );
  AND U11585 ( .A(n5793), .B(p_input[4788]), .Z(o[4788]) );
  AND U11586 ( .A(p_input[24788]), .B(p_input[14788]), .Z(n5793) );
  AND U11587 ( .A(n5794), .B(p_input[4787]), .Z(o[4787]) );
  AND U11588 ( .A(p_input[24787]), .B(p_input[14787]), .Z(n5794) );
  AND U11589 ( .A(n5795), .B(p_input[4786]), .Z(o[4786]) );
  AND U11590 ( .A(p_input[24786]), .B(p_input[14786]), .Z(n5795) );
  AND U11591 ( .A(n5796), .B(p_input[4785]), .Z(o[4785]) );
  AND U11592 ( .A(p_input[24785]), .B(p_input[14785]), .Z(n5796) );
  AND U11593 ( .A(n5797), .B(p_input[4784]), .Z(o[4784]) );
  AND U11594 ( .A(p_input[24784]), .B(p_input[14784]), .Z(n5797) );
  AND U11595 ( .A(n5798), .B(p_input[4783]), .Z(o[4783]) );
  AND U11596 ( .A(p_input[24783]), .B(p_input[14783]), .Z(n5798) );
  AND U11597 ( .A(n5799), .B(p_input[4782]), .Z(o[4782]) );
  AND U11598 ( .A(p_input[24782]), .B(p_input[14782]), .Z(n5799) );
  AND U11599 ( .A(n5800), .B(p_input[4781]), .Z(o[4781]) );
  AND U11600 ( .A(p_input[24781]), .B(p_input[14781]), .Z(n5800) );
  AND U11601 ( .A(n5801), .B(p_input[4780]), .Z(o[4780]) );
  AND U11602 ( .A(p_input[24780]), .B(p_input[14780]), .Z(n5801) );
  AND U11603 ( .A(n5802), .B(p_input[477]), .Z(o[477]) );
  AND U11604 ( .A(p_input[20477]), .B(p_input[10477]), .Z(n5802) );
  AND U11605 ( .A(n5803), .B(p_input[4779]), .Z(o[4779]) );
  AND U11606 ( .A(p_input[24779]), .B(p_input[14779]), .Z(n5803) );
  AND U11607 ( .A(n5804), .B(p_input[4778]), .Z(o[4778]) );
  AND U11608 ( .A(p_input[24778]), .B(p_input[14778]), .Z(n5804) );
  AND U11609 ( .A(n5805), .B(p_input[4777]), .Z(o[4777]) );
  AND U11610 ( .A(p_input[24777]), .B(p_input[14777]), .Z(n5805) );
  AND U11611 ( .A(n5806), .B(p_input[4776]), .Z(o[4776]) );
  AND U11612 ( .A(p_input[24776]), .B(p_input[14776]), .Z(n5806) );
  AND U11613 ( .A(n5807), .B(p_input[4775]), .Z(o[4775]) );
  AND U11614 ( .A(p_input[24775]), .B(p_input[14775]), .Z(n5807) );
  AND U11615 ( .A(n5808), .B(p_input[4774]), .Z(o[4774]) );
  AND U11616 ( .A(p_input[24774]), .B(p_input[14774]), .Z(n5808) );
  AND U11617 ( .A(n5809), .B(p_input[4773]), .Z(o[4773]) );
  AND U11618 ( .A(p_input[24773]), .B(p_input[14773]), .Z(n5809) );
  AND U11619 ( .A(n5810), .B(p_input[4772]), .Z(o[4772]) );
  AND U11620 ( .A(p_input[24772]), .B(p_input[14772]), .Z(n5810) );
  AND U11621 ( .A(n5811), .B(p_input[4771]), .Z(o[4771]) );
  AND U11622 ( .A(p_input[24771]), .B(p_input[14771]), .Z(n5811) );
  AND U11623 ( .A(n5812), .B(p_input[4770]), .Z(o[4770]) );
  AND U11624 ( .A(p_input[24770]), .B(p_input[14770]), .Z(n5812) );
  AND U11625 ( .A(n5813), .B(p_input[476]), .Z(o[476]) );
  AND U11626 ( .A(p_input[20476]), .B(p_input[10476]), .Z(n5813) );
  AND U11627 ( .A(n5814), .B(p_input[4769]), .Z(o[4769]) );
  AND U11628 ( .A(p_input[24769]), .B(p_input[14769]), .Z(n5814) );
  AND U11629 ( .A(n5815), .B(p_input[4768]), .Z(o[4768]) );
  AND U11630 ( .A(p_input[24768]), .B(p_input[14768]), .Z(n5815) );
  AND U11631 ( .A(n5816), .B(p_input[4767]), .Z(o[4767]) );
  AND U11632 ( .A(p_input[24767]), .B(p_input[14767]), .Z(n5816) );
  AND U11633 ( .A(n5817), .B(p_input[4766]), .Z(o[4766]) );
  AND U11634 ( .A(p_input[24766]), .B(p_input[14766]), .Z(n5817) );
  AND U11635 ( .A(n5818), .B(p_input[4765]), .Z(o[4765]) );
  AND U11636 ( .A(p_input[24765]), .B(p_input[14765]), .Z(n5818) );
  AND U11637 ( .A(n5819), .B(p_input[4764]), .Z(o[4764]) );
  AND U11638 ( .A(p_input[24764]), .B(p_input[14764]), .Z(n5819) );
  AND U11639 ( .A(n5820), .B(p_input[4763]), .Z(o[4763]) );
  AND U11640 ( .A(p_input[24763]), .B(p_input[14763]), .Z(n5820) );
  AND U11641 ( .A(n5821), .B(p_input[4762]), .Z(o[4762]) );
  AND U11642 ( .A(p_input[24762]), .B(p_input[14762]), .Z(n5821) );
  AND U11643 ( .A(n5822), .B(p_input[4761]), .Z(o[4761]) );
  AND U11644 ( .A(p_input[24761]), .B(p_input[14761]), .Z(n5822) );
  AND U11645 ( .A(n5823), .B(p_input[4760]), .Z(o[4760]) );
  AND U11646 ( .A(p_input[24760]), .B(p_input[14760]), .Z(n5823) );
  AND U11647 ( .A(n5824), .B(p_input[475]), .Z(o[475]) );
  AND U11648 ( .A(p_input[20475]), .B(p_input[10475]), .Z(n5824) );
  AND U11649 ( .A(n5825), .B(p_input[4759]), .Z(o[4759]) );
  AND U11650 ( .A(p_input[24759]), .B(p_input[14759]), .Z(n5825) );
  AND U11651 ( .A(n5826), .B(p_input[4758]), .Z(o[4758]) );
  AND U11652 ( .A(p_input[24758]), .B(p_input[14758]), .Z(n5826) );
  AND U11653 ( .A(n5827), .B(p_input[4757]), .Z(o[4757]) );
  AND U11654 ( .A(p_input[24757]), .B(p_input[14757]), .Z(n5827) );
  AND U11655 ( .A(n5828), .B(p_input[4756]), .Z(o[4756]) );
  AND U11656 ( .A(p_input[24756]), .B(p_input[14756]), .Z(n5828) );
  AND U11657 ( .A(n5829), .B(p_input[4755]), .Z(o[4755]) );
  AND U11658 ( .A(p_input[24755]), .B(p_input[14755]), .Z(n5829) );
  AND U11659 ( .A(n5830), .B(p_input[4754]), .Z(o[4754]) );
  AND U11660 ( .A(p_input[24754]), .B(p_input[14754]), .Z(n5830) );
  AND U11661 ( .A(n5831), .B(p_input[4753]), .Z(o[4753]) );
  AND U11662 ( .A(p_input[24753]), .B(p_input[14753]), .Z(n5831) );
  AND U11663 ( .A(n5832), .B(p_input[4752]), .Z(o[4752]) );
  AND U11664 ( .A(p_input[24752]), .B(p_input[14752]), .Z(n5832) );
  AND U11665 ( .A(n5833), .B(p_input[4751]), .Z(o[4751]) );
  AND U11666 ( .A(p_input[24751]), .B(p_input[14751]), .Z(n5833) );
  AND U11667 ( .A(n5834), .B(p_input[4750]), .Z(o[4750]) );
  AND U11668 ( .A(p_input[24750]), .B(p_input[14750]), .Z(n5834) );
  AND U11669 ( .A(n5835), .B(p_input[474]), .Z(o[474]) );
  AND U11670 ( .A(p_input[20474]), .B(p_input[10474]), .Z(n5835) );
  AND U11671 ( .A(n5836), .B(p_input[4749]), .Z(o[4749]) );
  AND U11672 ( .A(p_input[24749]), .B(p_input[14749]), .Z(n5836) );
  AND U11673 ( .A(n5837), .B(p_input[4748]), .Z(o[4748]) );
  AND U11674 ( .A(p_input[24748]), .B(p_input[14748]), .Z(n5837) );
  AND U11675 ( .A(n5838), .B(p_input[4747]), .Z(o[4747]) );
  AND U11676 ( .A(p_input[24747]), .B(p_input[14747]), .Z(n5838) );
  AND U11677 ( .A(n5839), .B(p_input[4746]), .Z(o[4746]) );
  AND U11678 ( .A(p_input[24746]), .B(p_input[14746]), .Z(n5839) );
  AND U11679 ( .A(n5840), .B(p_input[4745]), .Z(o[4745]) );
  AND U11680 ( .A(p_input[24745]), .B(p_input[14745]), .Z(n5840) );
  AND U11681 ( .A(n5841), .B(p_input[4744]), .Z(o[4744]) );
  AND U11682 ( .A(p_input[24744]), .B(p_input[14744]), .Z(n5841) );
  AND U11683 ( .A(n5842), .B(p_input[4743]), .Z(o[4743]) );
  AND U11684 ( .A(p_input[24743]), .B(p_input[14743]), .Z(n5842) );
  AND U11685 ( .A(n5843), .B(p_input[4742]), .Z(o[4742]) );
  AND U11686 ( .A(p_input[24742]), .B(p_input[14742]), .Z(n5843) );
  AND U11687 ( .A(n5844), .B(p_input[4741]), .Z(o[4741]) );
  AND U11688 ( .A(p_input[24741]), .B(p_input[14741]), .Z(n5844) );
  AND U11689 ( .A(n5845), .B(p_input[4740]), .Z(o[4740]) );
  AND U11690 ( .A(p_input[24740]), .B(p_input[14740]), .Z(n5845) );
  AND U11691 ( .A(n5846), .B(p_input[473]), .Z(o[473]) );
  AND U11692 ( .A(p_input[20473]), .B(p_input[10473]), .Z(n5846) );
  AND U11693 ( .A(n5847), .B(p_input[4739]), .Z(o[4739]) );
  AND U11694 ( .A(p_input[24739]), .B(p_input[14739]), .Z(n5847) );
  AND U11695 ( .A(n5848), .B(p_input[4738]), .Z(o[4738]) );
  AND U11696 ( .A(p_input[24738]), .B(p_input[14738]), .Z(n5848) );
  AND U11697 ( .A(n5849), .B(p_input[4737]), .Z(o[4737]) );
  AND U11698 ( .A(p_input[24737]), .B(p_input[14737]), .Z(n5849) );
  AND U11699 ( .A(n5850), .B(p_input[4736]), .Z(o[4736]) );
  AND U11700 ( .A(p_input[24736]), .B(p_input[14736]), .Z(n5850) );
  AND U11701 ( .A(n5851), .B(p_input[4735]), .Z(o[4735]) );
  AND U11702 ( .A(p_input[24735]), .B(p_input[14735]), .Z(n5851) );
  AND U11703 ( .A(n5852), .B(p_input[4734]), .Z(o[4734]) );
  AND U11704 ( .A(p_input[24734]), .B(p_input[14734]), .Z(n5852) );
  AND U11705 ( .A(n5853), .B(p_input[4733]), .Z(o[4733]) );
  AND U11706 ( .A(p_input[24733]), .B(p_input[14733]), .Z(n5853) );
  AND U11707 ( .A(n5854), .B(p_input[4732]), .Z(o[4732]) );
  AND U11708 ( .A(p_input[24732]), .B(p_input[14732]), .Z(n5854) );
  AND U11709 ( .A(n5855), .B(p_input[4731]), .Z(o[4731]) );
  AND U11710 ( .A(p_input[24731]), .B(p_input[14731]), .Z(n5855) );
  AND U11711 ( .A(n5856), .B(p_input[4730]), .Z(o[4730]) );
  AND U11712 ( .A(p_input[24730]), .B(p_input[14730]), .Z(n5856) );
  AND U11713 ( .A(n5857), .B(p_input[472]), .Z(o[472]) );
  AND U11714 ( .A(p_input[20472]), .B(p_input[10472]), .Z(n5857) );
  AND U11715 ( .A(n5858), .B(p_input[4729]), .Z(o[4729]) );
  AND U11716 ( .A(p_input[24729]), .B(p_input[14729]), .Z(n5858) );
  AND U11717 ( .A(n5859), .B(p_input[4728]), .Z(o[4728]) );
  AND U11718 ( .A(p_input[24728]), .B(p_input[14728]), .Z(n5859) );
  AND U11719 ( .A(n5860), .B(p_input[4727]), .Z(o[4727]) );
  AND U11720 ( .A(p_input[24727]), .B(p_input[14727]), .Z(n5860) );
  AND U11721 ( .A(n5861), .B(p_input[4726]), .Z(o[4726]) );
  AND U11722 ( .A(p_input[24726]), .B(p_input[14726]), .Z(n5861) );
  AND U11723 ( .A(n5862), .B(p_input[4725]), .Z(o[4725]) );
  AND U11724 ( .A(p_input[24725]), .B(p_input[14725]), .Z(n5862) );
  AND U11725 ( .A(n5863), .B(p_input[4724]), .Z(o[4724]) );
  AND U11726 ( .A(p_input[24724]), .B(p_input[14724]), .Z(n5863) );
  AND U11727 ( .A(n5864), .B(p_input[4723]), .Z(o[4723]) );
  AND U11728 ( .A(p_input[24723]), .B(p_input[14723]), .Z(n5864) );
  AND U11729 ( .A(n5865), .B(p_input[4722]), .Z(o[4722]) );
  AND U11730 ( .A(p_input[24722]), .B(p_input[14722]), .Z(n5865) );
  AND U11731 ( .A(n5866), .B(p_input[4721]), .Z(o[4721]) );
  AND U11732 ( .A(p_input[24721]), .B(p_input[14721]), .Z(n5866) );
  AND U11733 ( .A(n5867), .B(p_input[4720]), .Z(o[4720]) );
  AND U11734 ( .A(p_input[24720]), .B(p_input[14720]), .Z(n5867) );
  AND U11735 ( .A(n5868), .B(p_input[471]), .Z(o[471]) );
  AND U11736 ( .A(p_input[20471]), .B(p_input[10471]), .Z(n5868) );
  AND U11737 ( .A(n5869), .B(p_input[4719]), .Z(o[4719]) );
  AND U11738 ( .A(p_input[24719]), .B(p_input[14719]), .Z(n5869) );
  AND U11739 ( .A(n5870), .B(p_input[4718]), .Z(o[4718]) );
  AND U11740 ( .A(p_input[24718]), .B(p_input[14718]), .Z(n5870) );
  AND U11741 ( .A(n5871), .B(p_input[4717]), .Z(o[4717]) );
  AND U11742 ( .A(p_input[24717]), .B(p_input[14717]), .Z(n5871) );
  AND U11743 ( .A(n5872), .B(p_input[4716]), .Z(o[4716]) );
  AND U11744 ( .A(p_input[24716]), .B(p_input[14716]), .Z(n5872) );
  AND U11745 ( .A(n5873), .B(p_input[4715]), .Z(o[4715]) );
  AND U11746 ( .A(p_input[24715]), .B(p_input[14715]), .Z(n5873) );
  AND U11747 ( .A(n5874), .B(p_input[4714]), .Z(o[4714]) );
  AND U11748 ( .A(p_input[24714]), .B(p_input[14714]), .Z(n5874) );
  AND U11749 ( .A(n5875), .B(p_input[4713]), .Z(o[4713]) );
  AND U11750 ( .A(p_input[24713]), .B(p_input[14713]), .Z(n5875) );
  AND U11751 ( .A(n5876), .B(p_input[4712]), .Z(o[4712]) );
  AND U11752 ( .A(p_input[24712]), .B(p_input[14712]), .Z(n5876) );
  AND U11753 ( .A(n5877), .B(p_input[4711]), .Z(o[4711]) );
  AND U11754 ( .A(p_input[24711]), .B(p_input[14711]), .Z(n5877) );
  AND U11755 ( .A(n5878), .B(p_input[4710]), .Z(o[4710]) );
  AND U11756 ( .A(p_input[24710]), .B(p_input[14710]), .Z(n5878) );
  AND U11757 ( .A(n5879), .B(p_input[470]), .Z(o[470]) );
  AND U11758 ( .A(p_input[20470]), .B(p_input[10470]), .Z(n5879) );
  AND U11759 ( .A(n5880), .B(p_input[4709]), .Z(o[4709]) );
  AND U11760 ( .A(p_input[24709]), .B(p_input[14709]), .Z(n5880) );
  AND U11761 ( .A(n5881), .B(p_input[4708]), .Z(o[4708]) );
  AND U11762 ( .A(p_input[24708]), .B(p_input[14708]), .Z(n5881) );
  AND U11763 ( .A(n5882), .B(p_input[4707]), .Z(o[4707]) );
  AND U11764 ( .A(p_input[24707]), .B(p_input[14707]), .Z(n5882) );
  AND U11765 ( .A(n5883), .B(p_input[4706]), .Z(o[4706]) );
  AND U11766 ( .A(p_input[24706]), .B(p_input[14706]), .Z(n5883) );
  AND U11767 ( .A(n5884), .B(p_input[4705]), .Z(o[4705]) );
  AND U11768 ( .A(p_input[24705]), .B(p_input[14705]), .Z(n5884) );
  AND U11769 ( .A(n5885), .B(p_input[4704]), .Z(o[4704]) );
  AND U11770 ( .A(p_input[24704]), .B(p_input[14704]), .Z(n5885) );
  AND U11771 ( .A(n5886), .B(p_input[4703]), .Z(o[4703]) );
  AND U11772 ( .A(p_input[24703]), .B(p_input[14703]), .Z(n5886) );
  AND U11773 ( .A(n5887), .B(p_input[4702]), .Z(o[4702]) );
  AND U11774 ( .A(p_input[24702]), .B(p_input[14702]), .Z(n5887) );
  AND U11775 ( .A(n5888), .B(p_input[4701]), .Z(o[4701]) );
  AND U11776 ( .A(p_input[24701]), .B(p_input[14701]), .Z(n5888) );
  AND U11777 ( .A(n5889), .B(p_input[4700]), .Z(o[4700]) );
  AND U11778 ( .A(p_input[24700]), .B(p_input[14700]), .Z(n5889) );
  AND U11779 ( .A(n5890), .B(p_input[46]), .Z(o[46]) );
  AND U11780 ( .A(p_input[20046]), .B(p_input[10046]), .Z(n5890) );
  AND U11781 ( .A(n5891), .B(p_input[469]), .Z(o[469]) );
  AND U11782 ( .A(p_input[20469]), .B(p_input[10469]), .Z(n5891) );
  AND U11783 ( .A(n5892), .B(p_input[4699]), .Z(o[4699]) );
  AND U11784 ( .A(p_input[24699]), .B(p_input[14699]), .Z(n5892) );
  AND U11785 ( .A(n5893), .B(p_input[4698]), .Z(o[4698]) );
  AND U11786 ( .A(p_input[24698]), .B(p_input[14698]), .Z(n5893) );
  AND U11787 ( .A(n5894), .B(p_input[4697]), .Z(o[4697]) );
  AND U11788 ( .A(p_input[24697]), .B(p_input[14697]), .Z(n5894) );
  AND U11789 ( .A(n5895), .B(p_input[4696]), .Z(o[4696]) );
  AND U11790 ( .A(p_input[24696]), .B(p_input[14696]), .Z(n5895) );
  AND U11791 ( .A(n5896), .B(p_input[4695]), .Z(o[4695]) );
  AND U11792 ( .A(p_input[24695]), .B(p_input[14695]), .Z(n5896) );
  AND U11793 ( .A(n5897), .B(p_input[4694]), .Z(o[4694]) );
  AND U11794 ( .A(p_input[24694]), .B(p_input[14694]), .Z(n5897) );
  AND U11795 ( .A(n5898), .B(p_input[4693]), .Z(o[4693]) );
  AND U11796 ( .A(p_input[24693]), .B(p_input[14693]), .Z(n5898) );
  AND U11797 ( .A(n5899), .B(p_input[4692]), .Z(o[4692]) );
  AND U11798 ( .A(p_input[24692]), .B(p_input[14692]), .Z(n5899) );
  AND U11799 ( .A(n5900), .B(p_input[4691]), .Z(o[4691]) );
  AND U11800 ( .A(p_input[24691]), .B(p_input[14691]), .Z(n5900) );
  AND U11801 ( .A(n5901), .B(p_input[4690]), .Z(o[4690]) );
  AND U11802 ( .A(p_input[24690]), .B(p_input[14690]), .Z(n5901) );
  AND U11803 ( .A(n5902), .B(p_input[468]), .Z(o[468]) );
  AND U11804 ( .A(p_input[20468]), .B(p_input[10468]), .Z(n5902) );
  AND U11805 ( .A(n5903), .B(p_input[4689]), .Z(o[4689]) );
  AND U11806 ( .A(p_input[24689]), .B(p_input[14689]), .Z(n5903) );
  AND U11807 ( .A(n5904), .B(p_input[4688]), .Z(o[4688]) );
  AND U11808 ( .A(p_input[24688]), .B(p_input[14688]), .Z(n5904) );
  AND U11809 ( .A(n5905), .B(p_input[4687]), .Z(o[4687]) );
  AND U11810 ( .A(p_input[24687]), .B(p_input[14687]), .Z(n5905) );
  AND U11811 ( .A(n5906), .B(p_input[4686]), .Z(o[4686]) );
  AND U11812 ( .A(p_input[24686]), .B(p_input[14686]), .Z(n5906) );
  AND U11813 ( .A(n5907), .B(p_input[4685]), .Z(o[4685]) );
  AND U11814 ( .A(p_input[24685]), .B(p_input[14685]), .Z(n5907) );
  AND U11815 ( .A(n5908), .B(p_input[4684]), .Z(o[4684]) );
  AND U11816 ( .A(p_input[24684]), .B(p_input[14684]), .Z(n5908) );
  AND U11817 ( .A(n5909), .B(p_input[4683]), .Z(o[4683]) );
  AND U11818 ( .A(p_input[24683]), .B(p_input[14683]), .Z(n5909) );
  AND U11819 ( .A(n5910), .B(p_input[4682]), .Z(o[4682]) );
  AND U11820 ( .A(p_input[24682]), .B(p_input[14682]), .Z(n5910) );
  AND U11821 ( .A(n5911), .B(p_input[4681]), .Z(o[4681]) );
  AND U11822 ( .A(p_input[24681]), .B(p_input[14681]), .Z(n5911) );
  AND U11823 ( .A(n5912), .B(p_input[4680]), .Z(o[4680]) );
  AND U11824 ( .A(p_input[24680]), .B(p_input[14680]), .Z(n5912) );
  AND U11825 ( .A(n5913), .B(p_input[467]), .Z(o[467]) );
  AND U11826 ( .A(p_input[20467]), .B(p_input[10467]), .Z(n5913) );
  AND U11827 ( .A(n5914), .B(p_input[4679]), .Z(o[4679]) );
  AND U11828 ( .A(p_input[24679]), .B(p_input[14679]), .Z(n5914) );
  AND U11829 ( .A(n5915), .B(p_input[4678]), .Z(o[4678]) );
  AND U11830 ( .A(p_input[24678]), .B(p_input[14678]), .Z(n5915) );
  AND U11831 ( .A(n5916), .B(p_input[4677]), .Z(o[4677]) );
  AND U11832 ( .A(p_input[24677]), .B(p_input[14677]), .Z(n5916) );
  AND U11833 ( .A(n5917), .B(p_input[4676]), .Z(o[4676]) );
  AND U11834 ( .A(p_input[24676]), .B(p_input[14676]), .Z(n5917) );
  AND U11835 ( .A(n5918), .B(p_input[4675]), .Z(o[4675]) );
  AND U11836 ( .A(p_input[24675]), .B(p_input[14675]), .Z(n5918) );
  AND U11837 ( .A(n5919), .B(p_input[4674]), .Z(o[4674]) );
  AND U11838 ( .A(p_input[24674]), .B(p_input[14674]), .Z(n5919) );
  AND U11839 ( .A(n5920), .B(p_input[4673]), .Z(o[4673]) );
  AND U11840 ( .A(p_input[24673]), .B(p_input[14673]), .Z(n5920) );
  AND U11841 ( .A(n5921), .B(p_input[4672]), .Z(o[4672]) );
  AND U11842 ( .A(p_input[24672]), .B(p_input[14672]), .Z(n5921) );
  AND U11843 ( .A(n5922), .B(p_input[4671]), .Z(o[4671]) );
  AND U11844 ( .A(p_input[24671]), .B(p_input[14671]), .Z(n5922) );
  AND U11845 ( .A(n5923), .B(p_input[4670]), .Z(o[4670]) );
  AND U11846 ( .A(p_input[24670]), .B(p_input[14670]), .Z(n5923) );
  AND U11847 ( .A(n5924), .B(p_input[466]), .Z(o[466]) );
  AND U11848 ( .A(p_input[20466]), .B(p_input[10466]), .Z(n5924) );
  AND U11849 ( .A(n5925), .B(p_input[4669]), .Z(o[4669]) );
  AND U11850 ( .A(p_input[24669]), .B(p_input[14669]), .Z(n5925) );
  AND U11851 ( .A(n5926), .B(p_input[4668]), .Z(o[4668]) );
  AND U11852 ( .A(p_input[24668]), .B(p_input[14668]), .Z(n5926) );
  AND U11853 ( .A(n5927), .B(p_input[4667]), .Z(o[4667]) );
  AND U11854 ( .A(p_input[24667]), .B(p_input[14667]), .Z(n5927) );
  AND U11855 ( .A(n5928), .B(p_input[4666]), .Z(o[4666]) );
  AND U11856 ( .A(p_input[24666]), .B(p_input[14666]), .Z(n5928) );
  AND U11857 ( .A(n5929), .B(p_input[4665]), .Z(o[4665]) );
  AND U11858 ( .A(p_input[24665]), .B(p_input[14665]), .Z(n5929) );
  AND U11859 ( .A(n5930), .B(p_input[4664]), .Z(o[4664]) );
  AND U11860 ( .A(p_input[24664]), .B(p_input[14664]), .Z(n5930) );
  AND U11861 ( .A(n5931), .B(p_input[4663]), .Z(o[4663]) );
  AND U11862 ( .A(p_input[24663]), .B(p_input[14663]), .Z(n5931) );
  AND U11863 ( .A(n5932), .B(p_input[4662]), .Z(o[4662]) );
  AND U11864 ( .A(p_input[24662]), .B(p_input[14662]), .Z(n5932) );
  AND U11865 ( .A(n5933), .B(p_input[4661]), .Z(o[4661]) );
  AND U11866 ( .A(p_input[24661]), .B(p_input[14661]), .Z(n5933) );
  AND U11867 ( .A(n5934), .B(p_input[4660]), .Z(o[4660]) );
  AND U11868 ( .A(p_input[24660]), .B(p_input[14660]), .Z(n5934) );
  AND U11869 ( .A(n5935), .B(p_input[465]), .Z(o[465]) );
  AND U11870 ( .A(p_input[20465]), .B(p_input[10465]), .Z(n5935) );
  AND U11871 ( .A(n5936), .B(p_input[4659]), .Z(o[4659]) );
  AND U11872 ( .A(p_input[24659]), .B(p_input[14659]), .Z(n5936) );
  AND U11873 ( .A(n5937), .B(p_input[4658]), .Z(o[4658]) );
  AND U11874 ( .A(p_input[24658]), .B(p_input[14658]), .Z(n5937) );
  AND U11875 ( .A(n5938), .B(p_input[4657]), .Z(o[4657]) );
  AND U11876 ( .A(p_input[24657]), .B(p_input[14657]), .Z(n5938) );
  AND U11877 ( .A(n5939), .B(p_input[4656]), .Z(o[4656]) );
  AND U11878 ( .A(p_input[24656]), .B(p_input[14656]), .Z(n5939) );
  AND U11879 ( .A(n5940), .B(p_input[4655]), .Z(o[4655]) );
  AND U11880 ( .A(p_input[24655]), .B(p_input[14655]), .Z(n5940) );
  AND U11881 ( .A(n5941), .B(p_input[4654]), .Z(o[4654]) );
  AND U11882 ( .A(p_input[24654]), .B(p_input[14654]), .Z(n5941) );
  AND U11883 ( .A(n5942), .B(p_input[4653]), .Z(o[4653]) );
  AND U11884 ( .A(p_input[24653]), .B(p_input[14653]), .Z(n5942) );
  AND U11885 ( .A(n5943), .B(p_input[4652]), .Z(o[4652]) );
  AND U11886 ( .A(p_input[24652]), .B(p_input[14652]), .Z(n5943) );
  AND U11887 ( .A(n5944), .B(p_input[4651]), .Z(o[4651]) );
  AND U11888 ( .A(p_input[24651]), .B(p_input[14651]), .Z(n5944) );
  AND U11889 ( .A(n5945), .B(p_input[4650]), .Z(o[4650]) );
  AND U11890 ( .A(p_input[24650]), .B(p_input[14650]), .Z(n5945) );
  AND U11891 ( .A(n5946), .B(p_input[464]), .Z(o[464]) );
  AND U11892 ( .A(p_input[20464]), .B(p_input[10464]), .Z(n5946) );
  AND U11893 ( .A(n5947), .B(p_input[4649]), .Z(o[4649]) );
  AND U11894 ( .A(p_input[24649]), .B(p_input[14649]), .Z(n5947) );
  AND U11895 ( .A(n5948), .B(p_input[4648]), .Z(o[4648]) );
  AND U11896 ( .A(p_input[24648]), .B(p_input[14648]), .Z(n5948) );
  AND U11897 ( .A(n5949), .B(p_input[4647]), .Z(o[4647]) );
  AND U11898 ( .A(p_input[24647]), .B(p_input[14647]), .Z(n5949) );
  AND U11899 ( .A(n5950), .B(p_input[4646]), .Z(o[4646]) );
  AND U11900 ( .A(p_input[24646]), .B(p_input[14646]), .Z(n5950) );
  AND U11901 ( .A(n5951), .B(p_input[4645]), .Z(o[4645]) );
  AND U11902 ( .A(p_input[24645]), .B(p_input[14645]), .Z(n5951) );
  AND U11903 ( .A(n5952), .B(p_input[4644]), .Z(o[4644]) );
  AND U11904 ( .A(p_input[24644]), .B(p_input[14644]), .Z(n5952) );
  AND U11905 ( .A(n5953), .B(p_input[4643]), .Z(o[4643]) );
  AND U11906 ( .A(p_input[24643]), .B(p_input[14643]), .Z(n5953) );
  AND U11907 ( .A(n5954), .B(p_input[4642]), .Z(o[4642]) );
  AND U11908 ( .A(p_input[24642]), .B(p_input[14642]), .Z(n5954) );
  AND U11909 ( .A(n5955), .B(p_input[4641]), .Z(o[4641]) );
  AND U11910 ( .A(p_input[24641]), .B(p_input[14641]), .Z(n5955) );
  AND U11911 ( .A(n5956), .B(p_input[4640]), .Z(o[4640]) );
  AND U11912 ( .A(p_input[24640]), .B(p_input[14640]), .Z(n5956) );
  AND U11913 ( .A(n5957), .B(p_input[463]), .Z(o[463]) );
  AND U11914 ( .A(p_input[20463]), .B(p_input[10463]), .Z(n5957) );
  AND U11915 ( .A(n5958), .B(p_input[4639]), .Z(o[4639]) );
  AND U11916 ( .A(p_input[24639]), .B(p_input[14639]), .Z(n5958) );
  AND U11917 ( .A(n5959), .B(p_input[4638]), .Z(o[4638]) );
  AND U11918 ( .A(p_input[24638]), .B(p_input[14638]), .Z(n5959) );
  AND U11919 ( .A(n5960), .B(p_input[4637]), .Z(o[4637]) );
  AND U11920 ( .A(p_input[24637]), .B(p_input[14637]), .Z(n5960) );
  AND U11921 ( .A(n5961), .B(p_input[4636]), .Z(o[4636]) );
  AND U11922 ( .A(p_input[24636]), .B(p_input[14636]), .Z(n5961) );
  AND U11923 ( .A(n5962), .B(p_input[4635]), .Z(o[4635]) );
  AND U11924 ( .A(p_input[24635]), .B(p_input[14635]), .Z(n5962) );
  AND U11925 ( .A(n5963), .B(p_input[4634]), .Z(o[4634]) );
  AND U11926 ( .A(p_input[24634]), .B(p_input[14634]), .Z(n5963) );
  AND U11927 ( .A(n5964), .B(p_input[4633]), .Z(o[4633]) );
  AND U11928 ( .A(p_input[24633]), .B(p_input[14633]), .Z(n5964) );
  AND U11929 ( .A(n5965), .B(p_input[4632]), .Z(o[4632]) );
  AND U11930 ( .A(p_input[24632]), .B(p_input[14632]), .Z(n5965) );
  AND U11931 ( .A(n5966), .B(p_input[4631]), .Z(o[4631]) );
  AND U11932 ( .A(p_input[24631]), .B(p_input[14631]), .Z(n5966) );
  AND U11933 ( .A(n5967), .B(p_input[4630]), .Z(o[4630]) );
  AND U11934 ( .A(p_input[24630]), .B(p_input[14630]), .Z(n5967) );
  AND U11935 ( .A(n5968), .B(p_input[462]), .Z(o[462]) );
  AND U11936 ( .A(p_input[20462]), .B(p_input[10462]), .Z(n5968) );
  AND U11937 ( .A(n5969), .B(p_input[4629]), .Z(o[4629]) );
  AND U11938 ( .A(p_input[24629]), .B(p_input[14629]), .Z(n5969) );
  AND U11939 ( .A(n5970), .B(p_input[4628]), .Z(o[4628]) );
  AND U11940 ( .A(p_input[24628]), .B(p_input[14628]), .Z(n5970) );
  AND U11941 ( .A(n5971), .B(p_input[4627]), .Z(o[4627]) );
  AND U11942 ( .A(p_input[24627]), .B(p_input[14627]), .Z(n5971) );
  AND U11943 ( .A(n5972), .B(p_input[4626]), .Z(o[4626]) );
  AND U11944 ( .A(p_input[24626]), .B(p_input[14626]), .Z(n5972) );
  AND U11945 ( .A(n5973), .B(p_input[4625]), .Z(o[4625]) );
  AND U11946 ( .A(p_input[24625]), .B(p_input[14625]), .Z(n5973) );
  AND U11947 ( .A(n5974), .B(p_input[4624]), .Z(o[4624]) );
  AND U11948 ( .A(p_input[24624]), .B(p_input[14624]), .Z(n5974) );
  AND U11949 ( .A(n5975), .B(p_input[4623]), .Z(o[4623]) );
  AND U11950 ( .A(p_input[24623]), .B(p_input[14623]), .Z(n5975) );
  AND U11951 ( .A(n5976), .B(p_input[4622]), .Z(o[4622]) );
  AND U11952 ( .A(p_input[24622]), .B(p_input[14622]), .Z(n5976) );
  AND U11953 ( .A(n5977), .B(p_input[4621]), .Z(o[4621]) );
  AND U11954 ( .A(p_input[24621]), .B(p_input[14621]), .Z(n5977) );
  AND U11955 ( .A(n5978), .B(p_input[4620]), .Z(o[4620]) );
  AND U11956 ( .A(p_input[24620]), .B(p_input[14620]), .Z(n5978) );
  AND U11957 ( .A(n5979), .B(p_input[461]), .Z(o[461]) );
  AND U11958 ( .A(p_input[20461]), .B(p_input[10461]), .Z(n5979) );
  AND U11959 ( .A(n5980), .B(p_input[4619]), .Z(o[4619]) );
  AND U11960 ( .A(p_input[24619]), .B(p_input[14619]), .Z(n5980) );
  AND U11961 ( .A(n5981), .B(p_input[4618]), .Z(o[4618]) );
  AND U11962 ( .A(p_input[24618]), .B(p_input[14618]), .Z(n5981) );
  AND U11963 ( .A(n5982), .B(p_input[4617]), .Z(o[4617]) );
  AND U11964 ( .A(p_input[24617]), .B(p_input[14617]), .Z(n5982) );
  AND U11965 ( .A(n5983), .B(p_input[4616]), .Z(o[4616]) );
  AND U11966 ( .A(p_input[24616]), .B(p_input[14616]), .Z(n5983) );
  AND U11967 ( .A(n5984), .B(p_input[4615]), .Z(o[4615]) );
  AND U11968 ( .A(p_input[24615]), .B(p_input[14615]), .Z(n5984) );
  AND U11969 ( .A(n5985), .B(p_input[4614]), .Z(o[4614]) );
  AND U11970 ( .A(p_input[24614]), .B(p_input[14614]), .Z(n5985) );
  AND U11971 ( .A(n5986), .B(p_input[4613]), .Z(o[4613]) );
  AND U11972 ( .A(p_input[24613]), .B(p_input[14613]), .Z(n5986) );
  AND U11973 ( .A(n5987), .B(p_input[4612]), .Z(o[4612]) );
  AND U11974 ( .A(p_input[24612]), .B(p_input[14612]), .Z(n5987) );
  AND U11975 ( .A(n5988), .B(p_input[4611]), .Z(o[4611]) );
  AND U11976 ( .A(p_input[24611]), .B(p_input[14611]), .Z(n5988) );
  AND U11977 ( .A(n5989), .B(p_input[4610]), .Z(o[4610]) );
  AND U11978 ( .A(p_input[24610]), .B(p_input[14610]), .Z(n5989) );
  AND U11979 ( .A(n5990), .B(p_input[460]), .Z(o[460]) );
  AND U11980 ( .A(p_input[20460]), .B(p_input[10460]), .Z(n5990) );
  AND U11981 ( .A(n5991), .B(p_input[4609]), .Z(o[4609]) );
  AND U11982 ( .A(p_input[24609]), .B(p_input[14609]), .Z(n5991) );
  AND U11983 ( .A(n5992), .B(p_input[4608]), .Z(o[4608]) );
  AND U11984 ( .A(p_input[24608]), .B(p_input[14608]), .Z(n5992) );
  AND U11985 ( .A(n5993), .B(p_input[4607]), .Z(o[4607]) );
  AND U11986 ( .A(p_input[24607]), .B(p_input[14607]), .Z(n5993) );
  AND U11987 ( .A(n5994), .B(p_input[4606]), .Z(o[4606]) );
  AND U11988 ( .A(p_input[24606]), .B(p_input[14606]), .Z(n5994) );
  AND U11989 ( .A(n5995), .B(p_input[4605]), .Z(o[4605]) );
  AND U11990 ( .A(p_input[24605]), .B(p_input[14605]), .Z(n5995) );
  AND U11991 ( .A(n5996), .B(p_input[4604]), .Z(o[4604]) );
  AND U11992 ( .A(p_input[24604]), .B(p_input[14604]), .Z(n5996) );
  AND U11993 ( .A(n5997), .B(p_input[4603]), .Z(o[4603]) );
  AND U11994 ( .A(p_input[24603]), .B(p_input[14603]), .Z(n5997) );
  AND U11995 ( .A(n5998), .B(p_input[4602]), .Z(o[4602]) );
  AND U11996 ( .A(p_input[24602]), .B(p_input[14602]), .Z(n5998) );
  AND U11997 ( .A(n5999), .B(p_input[4601]), .Z(o[4601]) );
  AND U11998 ( .A(p_input[24601]), .B(p_input[14601]), .Z(n5999) );
  AND U11999 ( .A(n6000), .B(p_input[4600]), .Z(o[4600]) );
  AND U12000 ( .A(p_input[24600]), .B(p_input[14600]), .Z(n6000) );
  AND U12001 ( .A(n6001), .B(p_input[45]), .Z(o[45]) );
  AND U12002 ( .A(p_input[20045]), .B(p_input[10045]), .Z(n6001) );
  AND U12003 ( .A(n6002), .B(p_input[459]), .Z(o[459]) );
  AND U12004 ( .A(p_input[20459]), .B(p_input[10459]), .Z(n6002) );
  AND U12005 ( .A(n6003), .B(p_input[4599]), .Z(o[4599]) );
  AND U12006 ( .A(p_input[24599]), .B(p_input[14599]), .Z(n6003) );
  AND U12007 ( .A(n6004), .B(p_input[4598]), .Z(o[4598]) );
  AND U12008 ( .A(p_input[24598]), .B(p_input[14598]), .Z(n6004) );
  AND U12009 ( .A(n6005), .B(p_input[4597]), .Z(o[4597]) );
  AND U12010 ( .A(p_input[24597]), .B(p_input[14597]), .Z(n6005) );
  AND U12011 ( .A(n6006), .B(p_input[4596]), .Z(o[4596]) );
  AND U12012 ( .A(p_input[24596]), .B(p_input[14596]), .Z(n6006) );
  AND U12013 ( .A(n6007), .B(p_input[4595]), .Z(o[4595]) );
  AND U12014 ( .A(p_input[24595]), .B(p_input[14595]), .Z(n6007) );
  AND U12015 ( .A(n6008), .B(p_input[4594]), .Z(o[4594]) );
  AND U12016 ( .A(p_input[24594]), .B(p_input[14594]), .Z(n6008) );
  AND U12017 ( .A(n6009), .B(p_input[4593]), .Z(o[4593]) );
  AND U12018 ( .A(p_input[24593]), .B(p_input[14593]), .Z(n6009) );
  AND U12019 ( .A(n6010), .B(p_input[4592]), .Z(o[4592]) );
  AND U12020 ( .A(p_input[24592]), .B(p_input[14592]), .Z(n6010) );
  AND U12021 ( .A(n6011), .B(p_input[4591]), .Z(o[4591]) );
  AND U12022 ( .A(p_input[24591]), .B(p_input[14591]), .Z(n6011) );
  AND U12023 ( .A(n6012), .B(p_input[4590]), .Z(o[4590]) );
  AND U12024 ( .A(p_input[24590]), .B(p_input[14590]), .Z(n6012) );
  AND U12025 ( .A(n6013), .B(p_input[458]), .Z(o[458]) );
  AND U12026 ( .A(p_input[20458]), .B(p_input[10458]), .Z(n6013) );
  AND U12027 ( .A(n6014), .B(p_input[4589]), .Z(o[4589]) );
  AND U12028 ( .A(p_input[24589]), .B(p_input[14589]), .Z(n6014) );
  AND U12029 ( .A(n6015), .B(p_input[4588]), .Z(o[4588]) );
  AND U12030 ( .A(p_input[24588]), .B(p_input[14588]), .Z(n6015) );
  AND U12031 ( .A(n6016), .B(p_input[4587]), .Z(o[4587]) );
  AND U12032 ( .A(p_input[24587]), .B(p_input[14587]), .Z(n6016) );
  AND U12033 ( .A(n6017), .B(p_input[4586]), .Z(o[4586]) );
  AND U12034 ( .A(p_input[24586]), .B(p_input[14586]), .Z(n6017) );
  AND U12035 ( .A(n6018), .B(p_input[4585]), .Z(o[4585]) );
  AND U12036 ( .A(p_input[24585]), .B(p_input[14585]), .Z(n6018) );
  AND U12037 ( .A(n6019), .B(p_input[4584]), .Z(o[4584]) );
  AND U12038 ( .A(p_input[24584]), .B(p_input[14584]), .Z(n6019) );
  AND U12039 ( .A(n6020), .B(p_input[4583]), .Z(o[4583]) );
  AND U12040 ( .A(p_input[24583]), .B(p_input[14583]), .Z(n6020) );
  AND U12041 ( .A(n6021), .B(p_input[4582]), .Z(o[4582]) );
  AND U12042 ( .A(p_input[24582]), .B(p_input[14582]), .Z(n6021) );
  AND U12043 ( .A(n6022), .B(p_input[4581]), .Z(o[4581]) );
  AND U12044 ( .A(p_input[24581]), .B(p_input[14581]), .Z(n6022) );
  AND U12045 ( .A(n6023), .B(p_input[4580]), .Z(o[4580]) );
  AND U12046 ( .A(p_input[24580]), .B(p_input[14580]), .Z(n6023) );
  AND U12047 ( .A(n6024), .B(p_input[457]), .Z(o[457]) );
  AND U12048 ( .A(p_input[20457]), .B(p_input[10457]), .Z(n6024) );
  AND U12049 ( .A(n6025), .B(p_input[4579]), .Z(o[4579]) );
  AND U12050 ( .A(p_input[24579]), .B(p_input[14579]), .Z(n6025) );
  AND U12051 ( .A(n6026), .B(p_input[4578]), .Z(o[4578]) );
  AND U12052 ( .A(p_input[24578]), .B(p_input[14578]), .Z(n6026) );
  AND U12053 ( .A(n6027), .B(p_input[4577]), .Z(o[4577]) );
  AND U12054 ( .A(p_input[24577]), .B(p_input[14577]), .Z(n6027) );
  AND U12055 ( .A(n6028), .B(p_input[4576]), .Z(o[4576]) );
  AND U12056 ( .A(p_input[24576]), .B(p_input[14576]), .Z(n6028) );
  AND U12057 ( .A(n6029), .B(p_input[4575]), .Z(o[4575]) );
  AND U12058 ( .A(p_input[24575]), .B(p_input[14575]), .Z(n6029) );
  AND U12059 ( .A(n6030), .B(p_input[4574]), .Z(o[4574]) );
  AND U12060 ( .A(p_input[24574]), .B(p_input[14574]), .Z(n6030) );
  AND U12061 ( .A(n6031), .B(p_input[4573]), .Z(o[4573]) );
  AND U12062 ( .A(p_input[24573]), .B(p_input[14573]), .Z(n6031) );
  AND U12063 ( .A(n6032), .B(p_input[4572]), .Z(o[4572]) );
  AND U12064 ( .A(p_input[24572]), .B(p_input[14572]), .Z(n6032) );
  AND U12065 ( .A(n6033), .B(p_input[4571]), .Z(o[4571]) );
  AND U12066 ( .A(p_input[24571]), .B(p_input[14571]), .Z(n6033) );
  AND U12067 ( .A(n6034), .B(p_input[4570]), .Z(o[4570]) );
  AND U12068 ( .A(p_input[24570]), .B(p_input[14570]), .Z(n6034) );
  AND U12069 ( .A(n6035), .B(p_input[456]), .Z(o[456]) );
  AND U12070 ( .A(p_input[20456]), .B(p_input[10456]), .Z(n6035) );
  AND U12071 ( .A(n6036), .B(p_input[4569]), .Z(o[4569]) );
  AND U12072 ( .A(p_input[24569]), .B(p_input[14569]), .Z(n6036) );
  AND U12073 ( .A(n6037), .B(p_input[4568]), .Z(o[4568]) );
  AND U12074 ( .A(p_input[24568]), .B(p_input[14568]), .Z(n6037) );
  AND U12075 ( .A(n6038), .B(p_input[4567]), .Z(o[4567]) );
  AND U12076 ( .A(p_input[24567]), .B(p_input[14567]), .Z(n6038) );
  AND U12077 ( .A(n6039), .B(p_input[4566]), .Z(o[4566]) );
  AND U12078 ( .A(p_input[24566]), .B(p_input[14566]), .Z(n6039) );
  AND U12079 ( .A(n6040), .B(p_input[4565]), .Z(o[4565]) );
  AND U12080 ( .A(p_input[24565]), .B(p_input[14565]), .Z(n6040) );
  AND U12081 ( .A(n6041), .B(p_input[4564]), .Z(o[4564]) );
  AND U12082 ( .A(p_input[24564]), .B(p_input[14564]), .Z(n6041) );
  AND U12083 ( .A(n6042), .B(p_input[4563]), .Z(o[4563]) );
  AND U12084 ( .A(p_input[24563]), .B(p_input[14563]), .Z(n6042) );
  AND U12085 ( .A(n6043), .B(p_input[4562]), .Z(o[4562]) );
  AND U12086 ( .A(p_input[24562]), .B(p_input[14562]), .Z(n6043) );
  AND U12087 ( .A(n6044), .B(p_input[4561]), .Z(o[4561]) );
  AND U12088 ( .A(p_input[24561]), .B(p_input[14561]), .Z(n6044) );
  AND U12089 ( .A(n6045), .B(p_input[4560]), .Z(o[4560]) );
  AND U12090 ( .A(p_input[24560]), .B(p_input[14560]), .Z(n6045) );
  AND U12091 ( .A(n6046), .B(p_input[455]), .Z(o[455]) );
  AND U12092 ( .A(p_input[20455]), .B(p_input[10455]), .Z(n6046) );
  AND U12093 ( .A(n6047), .B(p_input[4559]), .Z(o[4559]) );
  AND U12094 ( .A(p_input[24559]), .B(p_input[14559]), .Z(n6047) );
  AND U12095 ( .A(n6048), .B(p_input[4558]), .Z(o[4558]) );
  AND U12096 ( .A(p_input[24558]), .B(p_input[14558]), .Z(n6048) );
  AND U12097 ( .A(n6049), .B(p_input[4557]), .Z(o[4557]) );
  AND U12098 ( .A(p_input[24557]), .B(p_input[14557]), .Z(n6049) );
  AND U12099 ( .A(n6050), .B(p_input[4556]), .Z(o[4556]) );
  AND U12100 ( .A(p_input[24556]), .B(p_input[14556]), .Z(n6050) );
  AND U12101 ( .A(n6051), .B(p_input[4555]), .Z(o[4555]) );
  AND U12102 ( .A(p_input[24555]), .B(p_input[14555]), .Z(n6051) );
  AND U12103 ( .A(n6052), .B(p_input[4554]), .Z(o[4554]) );
  AND U12104 ( .A(p_input[24554]), .B(p_input[14554]), .Z(n6052) );
  AND U12105 ( .A(n6053), .B(p_input[4553]), .Z(o[4553]) );
  AND U12106 ( .A(p_input[24553]), .B(p_input[14553]), .Z(n6053) );
  AND U12107 ( .A(n6054), .B(p_input[4552]), .Z(o[4552]) );
  AND U12108 ( .A(p_input[24552]), .B(p_input[14552]), .Z(n6054) );
  AND U12109 ( .A(n6055), .B(p_input[4551]), .Z(o[4551]) );
  AND U12110 ( .A(p_input[24551]), .B(p_input[14551]), .Z(n6055) );
  AND U12111 ( .A(n6056), .B(p_input[4550]), .Z(o[4550]) );
  AND U12112 ( .A(p_input[24550]), .B(p_input[14550]), .Z(n6056) );
  AND U12113 ( .A(n6057), .B(p_input[454]), .Z(o[454]) );
  AND U12114 ( .A(p_input[20454]), .B(p_input[10454]), .Z(n6057) );
  AND U12115 ( .A(n6058), .B(p_input[4549]), .Z(o[4549]) );
  AND U12116 ( .A(p_input[24549]), .B(p_input[14549]), .Z(n6058) );
  AND U12117 ( .A(n6059), .B(p_input[4548]), .Z(o[4548]) );
  AND U12118 ( .A(p_input[24548]), .B(p_input[14548]), .Z(n6059) );
  AND U12119 ( .A(n6060), .B(p_input[4547]), .Z(o[4547]) );
  AND U12120 ( .A(p_input[24547]), .B(p_input[14547]), .Z(n6060) );
  AND U12121 ( .A(n6061), .B(p_input[4546]), .Z(o[4546]) );
  AND U12122 ( .A(p_input[24546]), .B(p_input[14546]), .Z(n6061) );
  AND U12123 ( .A(n6062), .B(p_input[4545]), .Z(o[4545]) );
  AND U12124 ( .A(p_input[24545]), .B(p_input[14545]), .Z(n6062) );
  AND U12125 ( .A(n6063), .B(p_input[4544]), .Z(o[4544]) );
  AND U12126 ( .A(p_input[24544]), .B(p_input[14544]), .Z(n6063) );
  AND U12127 ( .A(n6064), .B(p_input[4543]), .Z(o[4543]) );
  AND U12128 ( .A(p_input[24543]), .B(p_input[14543]), .Z(n6064) );
  AND U12129 ( .A(n6065), .B(p_input[4542]), .Z(o[4542]) );
  AND U12130 ( .A(p_input[24542]), .B(p_input[14542]), .Z(n6065) );
  AND U12131 ( .A(n6066), .B(p_input[4541]), .Z(o[4541]) );
  AND U12132 ( .A(p_input[24541]), .B(p_input[14541]), .Z(n6066) );
  AND U12133 ( .A(n6067), .B(p_input[4540]), .Z(o[4540]) );
  AND U12134 ( .A(p_input[24540]), .B(p_input[14540]), .Z(n6067) );
  AND U12135 ( .A(n6068), .B(p_input[453]), .Z(o[453]) );
  AND U12136 ( .A(p_input[20453]), .B(p_input[10453]), .Z(n6068) );
  AND U12137 ( .A(n6069), .B(p_input[4539]), .Z(o[4539]) );
  AND U12138 ( .A(p_input[24539]), .B(p_input[14539]), .Z(n6069) );
  AND U12139 ( .A(n6070), .B(p_input[4538]), .Z(o[4538]) );
  AND U12140 ( .A(p_input[24538]), .B(p_input[14538]), .Z(n6070) );
  AND U12141 ( .A(n6071), .B(p_input[4537]), .Z(o[4537]) );
  AND U12142 ( .A(p_input[24537]), .B(p_input[14537]), .Z(n6071) );
  AND U12143 ( .A(n6072), .B(p_input[4536]), .Z(o[4536]) );
  AND U12144 ( .A(p_input[24536]), .B(p_input[14536]), .Z(n6072) );
  AND U12145 ( .A(n6073), .B(p_input[4535]), .Z(o[4535]) );
  AND U12146 ( .A(p_input[24535]), .B(p_input[14535]), .Z(n6073) );
  AND U12147 ( .A(n6074), .B(p_input[4534]), .Z(o[4534]) );
  AND U12148 ( .A(p_input[24534]), .B(p_input[14534]), .Z(n6074) );
  AND U12149 ( .A(n6075), .B(p_input[4533]), .Z(o[4533]) );
  AND U12150 ( .A(p_input[24533]), .B(p_input[14533]), .Z(n6075) );
  AND U12151 ( .A(n6076), .B(p_input[4532]), .Z(o[4532]) );
  AND U12152 ( .A(p_input[24532]), .B(p_input[14532]), .Z(n6076) );
  AND U12153 ( .A(n6077), .B(p_input[4531]), .Z(o[4531]) );
  AND U12154 ( .A(p_input[24531]), .B(p_input[14531]), .Z(n6077) );
  AND U12155 ( .A(n6078), .B(p_input[4530]), .Z(o[4530]) );
  AND U12156 ( .A(p_input[24530]), .B(p_input[14530]), .Z(n6078) );
  AND U12157 ( .A(n6079), .B(p_input[452]), .Z(o[452]) );
  AND U12158 ( .A(p_input[20452]), .B(p_input[10452]), .Z(n6079) );
  AND U12159 ( .A(n6080), .B(p_input[4529]), .Z(o[4529]) );
  AND U12160 ( .A(p_input[24529]), .B(p_input[14529]), .Z(n6080) );
  AND U12161 ( .A(n6081), .B(p_input[4528]), .Z(o[4528]) );
  AND U12162 ( .A(p_input[24528]), .B(p_input[14528]), .Z(n6081) );
  AND U12163 ( .A(n6082), .B(p_input[4527]), .Z(o[4527]) );
  AND U12164 ( .A(p_input[24527]), .B(p_input[14527]), .Z(n6082) );
  AND U12165 ( .A(n6083), .B(p_input[4526]), .Z(o[4526]) );
  AND U12166 ( .A(p_input[24526]), .B(p_input[14526]), .Z(n6083) );
  AND U12167 ( .A(n6084), .B(p_input[4525]), .Z(o[4525]) );
  AND U12168 ( .A(p_input[24525]), .B(p_input[14525]), .Z(n6084) );
  AND U12169 ( .A(n6085), .B(p_input[4524]), .Z(o[4524]) );
  AND U12170 ( .A(p_input[24524]), .B(p_input[14524]), .Z(n6085) );
  AND U12171 ( .A(n6086), .B(p_input[4523]), .Z(o[4523]) );
  AND U12172 ( .A(p_input[24523]), .B(p_input[14523]), .Z(n6086) );
  AND U12173 ( .A(n6087), .B(p_input[4522]), .Z(o[4522]) );
  AND U12174 ( .A(p_input[24522]), .B(p_input[14522]), .Z(n6087) );
  AND U12175 ( .A(n6088), .B(p_input[4521]), .Z(o[4521]) );
  AND U12176 ( .A(p_input[24521]), .B(p_input[14521]), .Z(n6088) );
  AND U12177 ( .A(n6089), .B(p_input[4520]), .Z(o[4520]) );
  AND U12178 ( .A(p_input[24520]), .B(p_input[14520]), .Z(n6089) );
  AND U12179 ( .A(n6090), .B(p_input[451]), .Z(o[451]) );
  AND U12180 ( .A(p_input[20451]), .B(p_input[10451]), .Z(n6090) );
  AND U12181 ( .A(n6091), .B(p_input[4519]), .Z(o[4519]) );
  AND U12182 ( .A(p_input[24519]), .B(p_input[14519]), .Z(n6091) );
  AND U12183 ( .A(n6092), .B(p_input[4518]), .Z(o[4518]) );
  AND U12184 ( .A(p_input[24518]), .B(p_input[14518]), .Z(n6092) );
  AND U12185 ( .A(n6093), .B(p_input[4517]), .Z(o[4517]) );
  AND U12186 ( .A(p_input[24517]), .B(p_input[14517]), .Z(n6093) );
  AND U12187 ( .A(n6094), .B(p_input[4516]), .Z(o[4516]) );
  AND U12188 ( .A(p_input[24516]), .B(p_input[14516]), .Z(n6094) );
  AND U12189 ( .A(n6095), .B(p_input[4515]), .Z(o[4515]) );
  AND U12190 ( .A(p_input[24515]), .B(p_input[14515]), .Z(n6095) );
  AND U12191 ( .A(n6096), .B(p_input[4514]), .Z(o[4514]) );
  AND U12192 ( .A(p_input[24514]), .B(p_input[14514]), .Z(n6096) );
  AND U12193 ( .A(n6097), .B(p_input[4513]), .Z(o[4513]) );
  AND U12194 ( .A(p_input[24513]), .B(p_input[14513]), .Z(n6097) );
  AND U12195 ( .A(n6098), .B(p_input[4512]), .Z(o[4512]) );
  AND U12196 ( .A(p_input[24512]), .B(p_input[14512]), .Z(n6098) );
  AND U12197 ( .A(n6099), .B(p_input[4511]), .Z(o[4511]) );
  AND U12198 ( .A(p_input[24511]), .B(p_input[14511]), .Z(n6099) );
  AND U12199 ( .A(n6100), .B(p_input[4510]), .Z(o[4510]) );
  AND U12200 ( .A(p_input[24510]), .B(p_input[14510]), .Z(n6100) );
  AND U12201 ( .A(n6101), .B(p_input[450]), .Z(o[450]) );
  AND U12202 ( .A(p_input[20450]), .B(p_input[10450]), .Z(n6101) );
  AND U12203 ( .A(n6102), .B(p_input[4509]), .Z(o[4509]) );
  AND U12204 ( .A(p_input[24509]), .B(p_input[14509]), .Z(n6102) );
  AND U12205 ( .A(n6103), .B(p_input[4508]), .Z(o[4508]) );
  AND U12206 ( .A(p_input[24508]), .B(p_input[14508]), .Z(n6103) );
  AND U12207 ( .A(n6104), .B(p_input[4507]), .Z(o[4507]) );
  AND U12208 ( .A(p_input[24507]), .B(p_input[14507]), .Z(n6104) );
  AND U12209 ( .A(n6105), .B(p_input[4506]), .Z(o[4506]) );
  AND U12210 ( .A(p_input[24506]), .B(p_input[14506]), .Z(n6105) );
  AND U12211 ( .A(n6106), .B(p_input[4505]), .Z(o[4505]) );
  AND U12212 ( .A(p_input[24505]), .B(p_input[14505]), .Z(n6106) );
  AND U12213 ( .A(n6107), .B(p_input[4504]), .Z(o[4504]) );
  AND U12214 ( .A(p_input[24504]), .B(p_input[14504]), .Z(n6107) );
  AND U12215 ( .A(n6108), .B(p_input[4503]), .Z(o[4503]) );
  AND U12216 ( .A(p_input[24503]), .B(p_input[14503]), .Z(n6108) );
  AND U12217 ( .A(n6109), .B(p_input[4502]), .Z(o[4502]) );
  AND U12218 ( .A(p_input[24502]), .B(p_input[14502]), .Z(n6109) );
  AND U12219 ( .A(n6110), .B(p_input[4501]), .Z(o[4501]) );
  AND U12220 ( .A(p_input[24501]), .B(p_input[14501]), .Z(n6110) );
  AND U12221 ( .A(n6111), .B(p_input[4500]), .Z(o[4500]) );
  AND U12222 ( .A(p_input[24500]), .B(p_input[14500]), .Z(n6111) );
  AND U12223 ( .A(n6112), .B(p_input[44]), .Z(o[44]) );
  AND U12224 ( .A(p_input[20044]), .B(p_input[10044]), .Z(n6112) );
  AND U12225 ( .A(n6113), .B(p_input[449]), .Z(o[449]) );
  AND U12226 ( .A(p_input[20449]), .B(p_input[10449]), .Z(n6113) );
  AND U12227 ( .A(n6114), .B(p_input[4499]), .Z(o[4499]) );
  AND U12228 ( .A(p_input[24499]), .B(p_input[14499]), .Z(n6114) );
  AND U12229 ( .A(n6115), .B(p_input[4498]), .Z(o[4498]) );
  AND U12230 ( .A(p_input[24498]), .B(p_input[14498]), .Z(n6115) );
  AND U12231 ( .A(n6116), .B(p_input[4497]), .Z(o[4497]) );
  AND U12232 ( .A(p_input[24497]), .B(p_input[14497]), .Z(n6116) );
  AND U12233 ( .A(n6117), .B(p_input[4496]), .Z(o[4496]) );
  AND U12234 ( .A(p_input[24496]), .B(p_input[14496]), .Z(n6117) );
  AND U12235 ( .A(n6118), .B(p_input[4495]), .Z(o[4495]) );
  AND U12236 ( .A(p_input[24495]), .B(p_input[14495]), .Z(n6118) );
  AND U12237 ( .A(n6119), .B(p_input[4494]), .Z(o[4494]) );
  AND U12238 ( .A(p_input[24494]), .B(p_input[14494]), .Z(n6119) );
  AND U12239 ( .A(n6120), .B(p_input[4493]), .Z(o[4493]) );
  AND U12240 ( .A(p_input[24493]), .B(p_input[14493]), .Z(n6120) );
  AND U12241 ( .A(n6121), .B(p_input[4492]), .Z(o[4492]) );
  AND U12242 ( .A(p_input[24492]), .B(p_input[14492]), .Z(n6121) );
  AND U12243 ( .A(n6122), .B(p_input[4491]), .Z(o[4491]) );
  AND U12244 ( .A(p_input[24491]), .B(p_input[14491]), .Z(n6122) );
  AND U12245 ( .A(n6123), .B(p_input[4490]), .Z(o[4490]) );
  AND U12246 ( .A(p_input[24490]), .B(p_input[14490]), .Z(n6123) );
  AND U12247 ( .A(n6124), .B(p_input[448]), .Z(o[448]) );
  AND U12248 ( .A(p_input[20448]), .B(p_input[10448]), .Z(n6124) );
  AND U12249 ( .A(n6125), .B(p_input[4489]), .Z(o[4489]) );
  AND U12250 ( .A(p_input[24489]), .B(p_input[14489]), .Z(n6125) );
  AND U12251 ( .A(n6126), .B(p_input[4488]), .Z(o[4488]) );
  AND U12252 ( .A(p_input[24488]), .B(p_input[14488]), .Z(n6126) );
  AND U12253 ( .A(n6127), .B(p_input[4487]), .Z(o[4487]) );
  AND U12254 ( .A(p_input[24487]), .B(p_input[14487]), .Z(n6127) );
  AND U12255 ( .A(n6128), .B(p_input[4486]), .Z(o[4486]) );
  AND U12256 ( .A(p_input[24486]), .B(p_input[14486]), .Z(n6128) );
  AND U12257 ( .A(n6129), .B(p_input[4485]), .Z(o[4485]) );
  AND U12258 ( .A(p_input[24485]), .B(p_input[14485]), .Z(n6129) );
  AND U12259 ( .A(n6130), .B(p_input[4484]), .Z(o[4484]) );
  AND U12260 ( .A(p_input[24484]), .B(p_input[14484]), .Z(n6130) );
  AND U12261 ( .A(n6131), .B(p_input[4483]), .Z(o[4483]) );
  AND U12262 ( .A(p_input[24483]), .B(p_input[14483]), .Z(n6131) );
  AND U12263 ( .A(n6132), .B(p_input[4482]), .Z(o[4482]) );
  AND U12264 ( .A(p_input[24482]), .B(p_input[14482]), .Z(n6132) );
  AND U12265 ( .A(n6133), .B(p_input[4481]), .Z(o[4481]) );
  AND U12266 ( .A(p_input[24481]), .B(p_input[14481]), .Z(n6133) );
  AND U12267 ( .A(n6134), .B(p_input[4480]), .Z(o[4480]) );
  AND U12268 ( .A(p_input[24480]), .B(p_input[14480]), .Z(n6134) );
  AND U12269 ( .A(n6135), .B(p_input[447]), .Z(o[447]) );
  AND U12270 ( .A(p_input[20447]), .B(p_input[10447]), .Z(n6135) );
  AND U12271 ( .A(n6136), .B(p_input[4479]), .Z(o[4479]) );
  AND U12272 ( .A(p_input[24479]), .B(p_input[14479]), .Z(n6136) );
  AND U12273 ( .A(n6137), .B(p_input[4478]), .Z(o[4478]) );
  AND U12274 ( .A(p_input[24478]), .B(p_input[14478]), .Z(n6137) );
  AND U12275 ( .A(n6138), .B(p_input[4477]), .Z(o[4477]) );
  AND U12276 ( .A(p_input[24477]), .B(p_input[14477]), .Z(n6138) );
  AND U12277 ( .A(n6139), .B(p_input[4476]), .Z(o[4476]) );
  AND U12278 ( .A(p_input[24476]), .B(p_input[14476]), .Z(n6139) );
  AND U12279 ( .A(n6140), .B(p_input[4475]), .Z(o[4475]) );
  AND U12280 ( .A(p_input[24475]), .B(p_input[14475]), .Z(n6140) );
  AND U12281 ( .A(n6141), .B(p_input[4474]), .Z(o[4474]) );
  AND U12282 ( .A(p_input[24474]), .B(p_input[14474]), .Z(n6141) );
  AND U12283 ( .A(n6142), .B(p_input[4473]), .Z(o[4473]) );
  AND U12284 ( .A(p_input[24473]), .B(p_input[14473]), .Z(n6142) );
  AND U12285 ( .A(n6143), .B(p_input[4472]), .Z(o[4472]) );
  AND U12286 ( .A(p_input[24472]), .B(p_input[14472]), .Z(n6143) );
  AND U12287 ( .A(n6144), .B(p_input[4471]), .Z(o[4471]) );
  AND U12288 ( .A(p_input[24471]), .B(p_input[14471]), .Z(n6144) );
  AND U12289 ( .A(n6145), .B(p_input[4470]), .Z(o[4470]) );
  AND U12290 ( .A(p_input[24470]), .B(p_input[14470]), .Z(n6145) );
  AND U12291 ( .A(n6146), .B(p_input[446]), .Z(o[446]) );
  AND U12292 ( .A(p_input[20446]), .B(p_input[10446]), .Z(n6146) );
  AND U12293 ( .A(n6147), .B(p_input[4469]), .Z(o[4469]) );
  AND U12294 ( .A(p_input[24469]), .B(p_input[14469]), .Z(n6147) );
  AND U12295 ( .A(n6148), .B(p_input[4468]), .Z(o[4468]) );
  AND U12296 ( .A(p_input[24468]), .B(p_input[14468]), .Z(n6148) );
  AND U12297 ( .A(n6149), .B(p_input[4467]), .Z(o[4467]) );
  AND U12298 ( .A(p_input[24467]), .B(p_input[14467]), .Z(n6149) );
  AND U12299 ( .A(n6150), .B(p_input[4466]), .Z(o[4466]) );
  AND U12300 ( .A(p_input[24466]), .B(p_input[14466]), .Z(n6150) );
  AND U12301 ( .A(n6151), .B(p_input[4465]), .Z(o[4465]) );
  AND U12302 ( .A(p_input[24465]), .B(p_input[14465]), .Z(n6151) );
  AND U12303 ( .A(n6152), .B(p_input[4464]), .Z(o[4464]) );
  AND U12304 ( .A(p_input[24464]), .B(p_input[14464]), .Z(n6152) );
  AND U12305 ( .A(n6153), .B(p_input[4463]), .Z(o[4463]) );
  AND U12306 ( .A(p_input[24463]), .B(p_input[14463]), .Z(n6153) );
  AND U12307 ( .A(n6154), .B(p_input[4462]), .Z(o[4462]) );
  AND U12308 ( .A(p_input[24462]), .B(p_input[14462]), .Z(n6154) );
  AND U12309 ( .A(n6155), .B(p_input[4461]), .Z(o[4461]) );
  AND U12310 ( .A(p_input[24461]), .B(p_input[14461]), .Z(n6155) );
  AND U12311 ( .A(n6156), .B(p_input[4460]), .Z(o[4460]) );
  AND U12312 ( .A(p_input[24460]), .B(p_input[14460]), .Z(n6156) );
  AND U12313 ( .A(n6157), .B(p_input[445]), .Z(o[445]) );
  AND U12314 ( .A(p_input[20445]), .B(p_input[10445]), .Z(n6157) );
  AND U12315 ( .A(n6158), .B(p_input[4459]), .Z(o[4459]) );
  AND U12316 ( .A(p_input[24459]), .B(p_input[14459]), .Z(n6158) );
  AND U12317 ( .A(n6159), .B(p_input[4458]), .Z(o[4458]) );
  AND U12318 ( .A(p_input[24458]), .B(p_input[14458]), .Z(n6159) );
  AND U12319 ( .A(n6160), .B(p_input[4457]), .Z(o[4457]) );
  AND U12320 ( .A(p_input[24457]), .B(p_input[14457]), .Z(n6160) );
  AND U12321 ( .A(n6161), .B(p_input[4456]), .Z(o[4456]) );
  AND U12322 ( .A(p_input[24456]), .B(p_input[14456]), .Z(n6161) );
  AND U12323 ( .A(n6162), .B(p_input[4455]), .Z(o[4455]) );
  AND U12324 ( .A(p_input[24455]), .B(p_input[14455]), .Z(n6162) );
  AND U12325 ( .A(n6163), .B(p_input[4454]), .Z(o[4454]) );
  AND U12326 ( .A(p_input[24454]), .B(p_input[14454]), .Z(n6163) );
  AND U12327 ( .A(n6164), .B(p_input[4453]), .Z(o[4453]) );
  AND U12328 ( .A(p_input[24453]), .B(p_input[14453]), .Z(n6164) );
  AND U12329 ( .A(n6165), .B(p_input[4452]), .Z(o[4452]) );
  AND U12330 ( .A(p_input[24452]), .B(p_input[14452]), .Z(n6165) );
  AND U12331 ( .A(n6166), .B(p_input[4451]), .Z(o[4451]) );
  AND U12332 ( .A(p_input[24451]), .B(p_input[14451]), .Z(n6166) );
  AND U12333 ( .A(n6167), .B(p_input[4450]), .Z(o[4450]) );
  AND U12334 ( .A(p_input[24450]), .B(p_input[14450]), .Z(n6167) );
  AND U12335 ( .A(n6168), .B(p_input[444]), .Z(o[444]) );
  AND U12336 ( .A(p_input[20444]), .B(p_input[10444]), .Z(n6168) );
  AND U12337 ( .A(n6169), .B(p_input[4449]), .Z(o[4449]) );
  AND U12338 ( .A(p_input[24449]), .B(p_input[14449]), .Z(n6169) );
  AND U12339 ( .A(n6170), .B(p_input[4448]), .Z(o[4448]) );
  AND U12340 ( .A(p_input[24448]), .B(p_input[14448]), .Z(n6170) );
  AND U12341 ( .A(n6171), .B(p_input[4447]), .Z(o[4447]) );
  AND U12342 ( .A(p_input[24447]), .B(p_input[14447]), .Z(n6171) );
  AND U12343 ( .A(n6172), .B(p_input[4446]), .Z(o[4446]) );
  AND U12344 ( .A(p_input[24446]), .B(p_input[14446]), .Z(n6172) );
  AND U12345 ( .A(n6173), .B(p_input[4445]), .Z(o[4445]) );
  AND U12346 ( .A(p_input[24445]), .B(p_input[14445]), .Z(n6173) );
  AND U12347 ( .A(n6174), .B(p_input[4444]), .Z(o[4444]) );
  AND U12348 ( .A(p_input[24444]), .B(p_input[14444]), .Z(n6174) );
  AND U12349 ( .A(n6175), .B(p_input[4443]), .Z(o[4443]) );
  AND U12350 ( .A(p_input[24443]), .B(p_input[14443]), .Z(n6175) );
  AND U12351 ( .A(n6176), .B(p_input[4442]), .Z(o[4442]) );
  AND U12352 ( .A(p_input[24442]), .B(p_input[14442]), .Z(n6176) );
  AND U12353 ( .A(n6177), .B(p_input[4441]), .Z(o[4441]) );
  AND U12354 ( .A(p_input[24441]), .B(p_input[14441]), .Z(n6177) );
  AND U12355 ( .A(n6178), .B(p_input[4440]), .Z(o[4440]) );
  AND U12356 ( .A(p_input[24440]), .B(p_input[14440]), .Z(n6178) );
  AND U12357 ( .A(n6179), .B(p_input[443]), .Z(o[443]) );
  AND U12358 ( .A(p_input[20443]), .B(p_input[10443]), .Z(n6179) );
  AND U12359 ( .A(n6180), .B(p_input[4439]), .Z(o[4439]) );
  AND U12360 ( .A(p_input[24439]), .B(p_input[14439]), .Z(n6180) );
  AND U12361 ( .A(n6181), .B(p_input[4438]), .Z(o[4438]) );
  AND U12362 ( .A(p_input[24438]), .B(p_input[14438]), .Z(n6181) );
  AND U12363 ( .A(n6182), .B(p_input[4437]), .Z(o[4437]) );
  AND U12364 ( .A(p_input[24437]), .B(p_input[14437]), .Z(n6182) );
  AND U12365 ( .A(n6183), .B(p_input[4436]), .Z(o[4436]) );
  AND U12366 ( .A(p_input[24436]), .B(p_input[14436]), .Z(n6183) );
  AND U12367 ( .A(n6184), .B(p_input[4435]), .Z(o[4435]) );
  AND U12368 ( .A(p_input[24435]), .B(p_input[14435]), .Z(n6184) );
  AND U12369 ( .A(n6185), .B(p_input[4434]), .Z(o[4434]) );
  AND U12370 ( .A(p_input[24434]), .B(p_input[14434]), .Z(n6185) );
  AND U12371 ( .A(n6186), .B(p_input[4433]), .Z(o[4433]) );
  AND U12372 ( .A(p_input[24433]), .B(p_input[14433]), .Z(n6186) );
  AND U12373 ( .A(n6187), .B(p_input[4432]), .Z(o[4432]) );
  AND U12374 ( .A(p_input[24432]), .B(p_input[14432]), .Z(n6187) );
  AND U12375 ( .A(n6188), .B(p_input[4431]), .Z(o[4431]) );
  AND U12376 ( .A(p_input[24431]), .B(p_input[14431]), .Z(n6188) );
  AND U12377 ( .A(n6189), .B(p_input[4430]), .Z(o[4430]) );
  AND U12378 ( .A(p_input[24430]), .B(p_input[14430]), .Z(n6189) );
  AND U12379 ( .A(n6190), .B(p_input[442]), .Z(o[442]) );
  AND U12380 ( .A(p_input[20442]), .B(p_input[10442]), .Z(n6190) );
  AND U12381 ( .A(n6191), .B(p_input[4429]), .Z(o[4429]) );
  AND U12382 ( .A(p_input[24429]), .B(p_input[14429]), .Z(n6191) );
  AND U12383 ( .A(n6192), .B(p_input[4428]), .Z(o[4428]) );
  AND U12384 ( .A(p_input[24428]), .B(p_input[14428]), .Z(n6192) );
  AND U12385 ( .A(n6193), .B(p_input[4427]), .Z(o[4427]) );
  AND U12386 ( .A(p_input[24427]), .B(p_input[14427]), .Z(n6193) );
  AND U12387 ( .A(n6194), .B(p_input[4426]), .Z(o[4426]) );
  AND U12388 ( .A(p_input[24426]), .B(p_input[14426]), .Z(n6194) );
  AND U12389 ( .A(n6195), .B(p_input[4425]), .Z(o[4425]) );
  AND U12390 ( .A(p_input[24425]), .B(p_input[14425]), .Z(n6195) );
  AND U12391 ( .A(n6196), .B(p_input[4424]), .Z(o[4424]) );
  AND U12392 ( .A(p_input[24424]), .B(p_input[14424]), .Z(n6196) );
  AND U12393 ( .A(n6197), .B(p_input[4423]), .Z(o[4423]) );
  AND U12394 ( .A(p_input[24423]), .B(p_input[14423]), .Z(n6197) );
  AND U12395 ( .A(n6198), .B(p_input[4422]), .Z(o[4422]) );
  AND U12396 ( .A(p_input[24422]), .B(p_input[14422]), .Z(n6198) );
  AND U12397 ( .A(n6199), .B(p_input[4421]), .Z(o[4421]) );
  AND U12398 ( .A(p_input[24421]), .B(p_input[14421]), .Z(n6199) );
  AND U12399 ( .A(n6200), .B(p_input[4420]), .Z(o[4420]) );
  AND U12400 ( .A(p_input[24420]), .B(p_input[14420]), .Z(n6200) );
  AND U12401 ( .A(n6201), .B(p_input[441]), .Z(o[441]) );
  AND U12402 ( .A(p_input[20441]), .B(p_input[10441]), .Z(n6201) );
  AND U12403 ( .A(n6202), .B(p_input[4419]), .Z(o[4419]) );
  AND U12404 ( .A(p_input[24419]), .B(p_input[14419]), .Z(n6202) );
  AND U12405 ( .A(n6203), .B(p_input[4418]), .Z(o[4418]) );
  AND U12406 ( .A(p_input[24418]), .B(p_input[14418]), .Z(n6203) );
  AND U12407 ( .A(n6204), .B(p_input[4417]), .Z(o[4417]) );
  AND U12408 ( .A(p_input[24417]), .B(p_input[14417]), .Z(n6204) );
  AND U12409 ( .A(n6205), .B(p_input[4416]), .Z(o[4416]) );
  AND U12410 ( .A(p_input[24416]), .B(p_input[14416]), .Z(n6205) );
  AND U12411 ( .A(n6206), .B(p_input[4415]), .Z(o[4415]) );
  AND U12412 ( .A(p_input[24415]), .B(p_input[14415]), .Z(n6206) );
  AND U12413 ( .A(n6207), .B(p_input[4414]), .Z(o[4414]) );
  AND U12414 ( .A(p_input[24414]), .B(p_input[14414]), .Z(n6207) );
  AND U12415 ( .A(n6208), .B(p_input[4413]), .Z(o[4413]) );
  AND U12416 ( .A(p_input[24413]), .B(p_input[14413]), .Z(n6208) );
  AND U12417 ( .A(n6209), .B(p_input[4412]), .Z(o[4412]) );
  AND U12418 ( .A(p_input[24412]), .B(p_input[14412]), .Z(n6209) );
  AND U12419 ( .A(n6210), .B(p_input[4411]), .Z(o[4411]) );
  AND U12420 ( .A(p_input[24411]), .B(p_input[14411]), .Z(n6210) );
  AND U12421 ( .A(n6211), .B(p_input[4410]), .Z(o[4410]) );
  AND U12422 ( .A(p_input[24410]), .B(p_input[14410]), .Z(n6211) );
  AND U12423 ( .A(n6212), .B(p_input[440]), .Z(o[440]) );
  AND U12424 ( .A(p_input[20440]), .B(p_input[10440]), .Z(n6212) );
  AND U12425 ( .A(n6213), .B(p_input[4409]), .Z(o[4409]) );
  AND U12426 ( .A(p_input[24409]), .B(p_input[14409]), .Z(n6213) );
  AND U12427 ( .A(n6214), .B(p_input[4408]), .Z(o[4408]) );
  AND U12428 ( .A(p_input[24408]), .B(p_input[14408]), .Z(n6214) );
  AND U12429 ( .A(n6215), .B(p_input[4407]), .Z(o[4407]) );
  AND U12430 ( .A(p_input[24407]), .B(p_input[14407]), .Z(n6215) );
  AND U12431 ( .A(n6216), .B(p_input[4406]), .Z(o[4406]) );
  AND U12432 ( .A(p_input[24406]), .B(p_input[14406]), .Z(n6216) );
  AND U12433 ( .A(n6217), .B(p_input[4405]), .Z(o[4405]) );
  AND U12434 ( .A(p_input[24405]), .B(p_input[14405]), .Z(n6217) );
  AND U12435 ( .A(n6218), .B(p_input[4404]), .Z(o[4404]) );
  AND U12436 ( .A(p_input[24404]), .B(p_input[14404]), .Z(n6218) );
  AND U12437 ( .A(n6219), .B(p_input[4403]), .Z(o[4403]) );
  AND U12438 ( .A(p_input[24403]), .B(p_input[14403]), .Z(n6219) );
  AND U12439 ( .A(n6220), .B(p_input[4402]), .Z(o[4402]) );
  AND U12440 ( .A(p_input[24402]), .B(p_input[14402]), .Z(n6220) );
  AND U12441 ( .A(n6221), .B(p_input[4401]), .Z(o[4401]) );
  AND U12442 ( .A(p_input[24401]), .B(p_input[14401]), .Z(n6221) );
  AND U12443 ( .A(n6222), .B(p_input[4400]), .Z(o[4400]) );
  AND U12444 ( .A(p_input[24400]), .B(p_input[14400]), .Z(n6222) );
  AND U12445 ( .A(n6223), .B(p_input[43]), .Z(o[43]) );
  AND U12446 ( .A(p_input[20043]), .B(p_input[10043]), .Z(n6223) );
  AND U12447 ( .A(n6224), .B(p_input[439]), .Z(o[439]) );
  AND U12448 ( .A(p_input[20439]), .B(p_input[10439]), .Z(n6224) );
  AND U12449 ( .A(n6225), .B(p_input[4399]), .Z(o[4399]) );
  AND U12450 ( .A(p_input[24399]), .B(p_input[14399]), .Z(n6225) );
  AND U12451 ( .A(n6226), .B(p_input[4398]), .Z(o[4398]) );
  AND U12452 ( .A(p_input[24398]), .B(p_input[14398]), .Z(n6226) );
  AND U12453 ( .A(n6227), .B(p_input[4397]), .Z(o[4397]) );
  AND U12454 ( .A(p_input[24397]), .B(p_input[14397]), .Z(n6227) );
  AND U12455 ( .A(n6228), .B(p_input[4396]), .Z(o[4396]) );
  AND U12456 ( .A(p_input[24396]), .B(p_input[14396]), .Z(n6228) );
  AND U12457 ( .A(n6229), .B(p_input[4395]), .Z(o[4395]) );
  AND U12458 ( .A(p_input[24395]), .B(p_input[14395]), .Z(n6229) );
  AND U12459 ( .A(n6230), .B(p_input[4394]), .Z(o[4394]) );
  AND U12460 ( .A(p_input[24394]), .B(p_input[14394]), .Z(n6230) );
  AND U12461 ( .A(n6231), .B(p_input[4393]), .Z(o[4393]) );
  AND U12462 ( .A(p_input[24393]), .B(p_input[14393]), .Z(n6231) );
  AND U12463 ( .A(n6232), .B(p_input[4392]), .Z(o[4392]) );
  AND U12464 ( .A(p_input[24392]), .B(p_input[14392]), .Z(n6232) );
  AND U12465 ( .A(n6233), .B(p_input[4391]), .Z(o[4391]) );
  AND U12466 ( .A(p_input[24391]), .B(p_input[14391]), .Z(n6233) );
  AND U12467 ( .A(n6234), .B(p_input[4390]), .Z(o[4390]) );
  AND U12468 ( .A(p_input[24390]), .B(p_input[14390]), .Z(n6234) );
  AND U12469 ( .A(n6235), .B(p_input[438]), .Z(o[438]) );
  AND U12470 ( .A(p_input[20438]), .B(p_input[10438]), .Z(n6235) );
  AND U12471 ( .A(n6236), .B(p_input[4389]), .Z(o[4389]) );
  AND U12472 ( .A(p_input[24389]), .B(p_input[14389]), .Z(n6236) );
  AND U12473 ( .A(n6237), .B(p_input[4388]), .Z(o[4388]) );
  AND U12474 ( .A(p_input[24388]), .B(p_input[14388]), .Z(n6237) );
  AND U12475 ( .A(n6238), .B(p_input[4387]), .Z(o[4387]) );
  AND U12476 ( .A(p_input[24387]), .B(p_input[14387]), .Z(n6238) );
  AND U12477 ( .A(n6239), .B(p_input[4386]), .Z(o[4386]) );
  AND U12478 ( .A(p_input[24386]), .B(p_input[14386]), .Z(n6239) );
  AND U12479 ( .A(n6240), .B(p_input[4385]), .Z(o[4385]) );
  AND U12480 ( .A(p_input[24385]), .B(p_input[14385]), .Z(n6240) );
  AND U12481 ( .A(n6241), .B(p_input[4384]), .Z(o[4384]) );
  AND U12482 ( .A(p_input[24384]), .B(p_input[14384]), .Z(n6241) );
  AND U12483 ( .A(n6242), .B(p_input[4383]), .Z(o[4383]) );
  AND U12484 ( .A(p_input[24383]), .B(p_input[14383]), .Z(n6242) );
  AND U12485 ( .A(n6243), .B(p_input[4382]), .Z(o[4382]) );
  AND U12486 ( .A(p_input[24382]), .B(p_input[14382]), .Z(n6243) );
  AND U12487 ( .A(n6244), .B(p_input[4381]), .Z(o[4381]) );
  AND U12488 ( .A(p_input[24381]), .B(p_input[14381]), .Z(n6244) );
  AND U12489 ( .A(n6245), .B(p_input[4380]), .Z(o[4380]) );
  AND U12490 ( .A(p_input[24380]), .B(p_input[14380]), .Z(n6245) );
  AND U12491 ( .A(n6246), .B(p_input[437]), .Z(o[437]) );
  AND U12492 ( .A(p_input[20437]), .B(p_input[10437]), .Z(n6246) );
  AND U12493 ( .A(n6247), .B(p_input[4379]), .Z(o[4379]) );
  AND U12494 ( .A(p_input[24379]), .B(p_input[14379]), .Z(n6247) );
  AND U12495 ( .A(n6248), .B(p_input[4378]), .Z(o[4378]) );
  AND U12496 ( .A(p_input[24378]), .B(p_input[14378]), .Z(n6248) );
  AND U12497 ( .A(n6249), .B(p_input[4377]), .Z(o[4377]) );
  AND U12498 ( .A(p_input[24377]), .B(p_input[14377]), .Z(n6249) );
  AND U12499 ( .A(n6250), .B(p_input[4376]), .Z(o[4376]) );
  AND U12500 ( .A(p_input[24376]), .B(p_input[14376]), .Z(n6250) );
  AND U12501 ( .A(n6251), .B(p_input[4375]), .Z(o[4375]) );
  AND U12502 ( .A(p_input[24375]), .B(p_input[14375]), .Z(n6251) );
  AND U12503 ( .A(n6252), .B(p_input[4374]), .Z(o[4374]) );
  AND U12504 ( .A(p_input[24374]), .B(p_input[14374]), .Z(n6252) );
  AND U12505 ( .A(n6253), .B(p_input[4373]), .Z(o[4373]) );
  AND U12506 ( .A(p_input[24373]), .B(p_input[14373]), .Z(n6253) );
  AND U12507 ( .A(n6254), .B(p_input[4372]), .Z(o[4372]) );
  AND U12508 ( .A(p_input[24372]), .B(p_input[14372]), .Z(n6254) );
  AND U12509 ( .A(n6255), .B(p_input[4371]), .Z(o[4371]) );
  AND U12510 ( .A(p_input[24371]), .B(p_input[14371]), .Z(n6255) );
  AND U12511 ( .A(n6256), .B(p_input[4370]), .Z(o[4370]) );
  AND U12512 ( .A(p_input[24370]), .B(p_input[14370]), .Z(n6256) );
  AND U12513 ( .A(n6257), .B(p_input[436]), .Z(o[436]) );
  AND U12514 ( .A(p_input[20436]), .B(p_input[10436]), .Z(n6257) );
  AND U12515 ( .A(n6258), .B(p_input[4369]), .Z(o[4369]) );
  AND U12516 ( .A(p_input[24369]), .B(p_input[14369]), .Z(n6258) );
  AND U12517 ( .A(n6259), .B(p_input[4368]), .Z(o[4368]) );
  AND U12518 ( .A(p_input[24368]), .B(p_input[14368]), .Z(n6259) );
  AND U12519 ( .A(n6260), .B(p_input[4367]), .Z(o[4367]) );
  AND U12520 ( .A(p_input[24367]), .B(p_input[14367]), .Z(n6260) );
  AND U12521 ( .A(n6261), .B(p_input[4366]), .Z(o[4366]) );
  AND U12522 ( .A(p_input[24366]), .B(p_input[14366]), .Z(n6261) );
  AND U12523 ( .A(n6262), .B(p_input[4365]), .Z(o[4365]) );
  AND U12524 ( .A(p_input[24365]), .B(p_input[14365]), .Z(n6262) );
  AND U12525 ( .A(n6263), .B(p_input[4364]), .Z(o[4364]) );
  AND U12526 ( .A(p_input[24364]), .B(p_input[14364]), .Z(n6263) );
  AND U12527 ( .A(n6264), .B(p_input[4363]), .Z(o[4363]) );
  AND U12528 ( .A(p_input[24363]), .B(p_input[14363]), .Z(n6264) );
  AND U12529 ( .A(n6265), .B(p_input[4362]), .Z(o[4362]) );
  AND U12530 ( .A(p_input[24362]), .B(p_input[14362]), .Z(n6265) );
  AND U12531 ( .A(n6266), .B(p_input[4361]), .Z(o[4361]) );
  AND U12532 ( .A(p_input[24361]), .B(p_input[14361]), .Z(n6266) );
  AND U12533 ( .A(n6267), .B(p_input[4360]), .Z(o[4360]) );
  AND U12534 ( .A(p_input[24360]), .B(p_input[14360]), .Z(n6267) );
  AND U12535 ( .A(n6268), .B(p_input[435]), .Z(o[435]) );
  AND U12536 ( .A(p_input[20435]), .B(p_input[10435]), .Z(n6268) );
  AND U12537 ( .A(n6269), .B(p_input[4359]), .Z(o[4359]) );
  AND U12538 ( .A(p_input[24359]), .B(p_input[14359]), .Z(n6269) );
  AND U12539 ( .A(n6270), .B(p_input[4358]), .Z(o[4358]) );
  AND U12540 ( .A(p_input[24358]), .B(p_input[14358]), .Z(n6270) );
  AND U12541 ( .A(n6271), .B(p_input[4357]), .Z(o[4357]) );
  AND U12542 ( .A(p_input[24357]), .B(p_input[14357]), .Z(n6271) );
  AND U12543 ( .A(n6272), .B(p_input[4356]), .Z(o[4356]) );
  AND U12544 ( .A(p_input[24356]), .B(p_input[14356]), .Z(n6272) );
  AND U12545 ( .A(n6273), .B(p_input[4355]), .Z(o[4355]) );
  AND U12546 ( .A(p_input[24355]), .B(p_input[14355]), .Z(n6273) );
  AND U12547 ( .A(n6274), .B(p_input[4354]), .Z(o[4354]) );
  AND U12548 ( .A(p_input[24354]), .B(p_input[14354]), .Z(n6274) );
  AND U12549 ( .A(n6275), .B(p_input[4353]), .Z(o[4353]) );
  AND U12550 ( .A(p_input[24353]), .B(p_input[14353]), .Z(n6275) );
  AND U12551 ( .A(n6276), .B(p_input[4352]), .Z(o[4352]) );
  AND U12552 ( .A(p_input[24352]), .B(p_input[14352]), .Z(n6276) );
  AND U12553 ( .A(n6277), .B(p_input[4351]), .Z(o[4351]) );
  AND U12554 ( .A(p_input[24351]), .B(p_input[14351]), .Z(n6277) );
  AND U12555 ( .A(n6278), .B(p_input[4350]), .Z(o[4350]) );
  AND U12556 ( .A(p_input[24350]), .B(p_input[14350]), .Z(n6278) );
  AND U12557 ( .A(n6279), .B(p_input[434]), .Z(o[434]) );
  AND U12558 ( .A(p_input[20434]), .B(p_input[10434]), .Z(n6279) );
  AND U12559 ( .A(n6280), .B(p_input[4349]), .Z(o[4349]) );
  AND U12560 ( .A(p_input[24349]), .B(p_input[14349]), .Z(n6280) );
  AND U12561 ( .A(n6281), .B(p_input[4348]), .Z(o[4348]) );
  AND U12562 ( .A(p_input[24348]), .B(p_input[14348]), .Z(n6281) );
  AND U12563 ( .A(n6282), .B(p_input[4347]), .Z(o[4347]) );
  AND U12564 ( .A(p_input[24347]), .B(p_input[14347]), .Z(n6282) );
  AND U12565 ( .A(n6283), .B(p_input[4346]), .Z(o[4346]) );
  AND U12566 ( .A(p_input[24346]), .B(p_input[14346]), .Z(n6283) );
  AND U12567 ( .A(n6284), .B(p_input[4345]), .Z(o[4345]) );
  AND U12568 ( .A(p_input[24345]), .B(p_input[14345]), .Z(n6284) );
  AND U12569 ( .A(n6285), .B(p_input[4344]), .Z(o[4344]) );
  AND U12570 ( .A(p_input[24344]), .B(p_input[14344]), .Z(n6285) );
  AND U12571 ( .A(n6286), .B(p_input[4343]), .Z(o[4343]) );
  AND U12572 ( .A(p_input[24343]), .B(p_input[14343]), .Z(n6286) );
  AND U12573 ( .A(n6287), .B(p_input[4342]), .Z(o[4342]) );
  AND U12574 ( .A(p_input[24342]), .B(p_input[14342]), .Z(n6287) );
  AND U12575 ( .A(n6288), .B(p_input[4341]), .Z(o[4341]) );
  AND U12576 ( .A(p_input[24341]), .B(p_input[14341]), .Z(n6288) );
  AND U12577 ( .A(n6289), .B(p_input[4340]), .Z(o[4340]) );
  AND U12578 ( .A(p_input[24340]), .B(p_input[14340]), .Z(n6289) );
  AND U12579 ( .A(n6290), .B(p_input[433]), .Z(o[433]) );
  AND U12580 ( .A(p_input[20433]), .B(p_input[10433]), .Z(n6290) );
  AND U12581 ( .A(n6291), .B(p_input[4339]), .Z(o[4339]) );
  AND U12582 ( .A(p_input[24339]), .B(p_input[14339]), .Z(n6291) );
  AND U12583 ( .A(n6292), .B(p_input[4338]), .Z(o[4338]) );
  AND U12584 ( .A(p_input[24338]), .B(p_input[14338]), .Z(n6292) );
  AND U12585 ( .A(n6293), .B(p_input[4337]), .Z(o[4337]) );
  AND U12586 ( .A(p_input[24337]), .B(p_input[14337]), .Z(n6293) );
  AND U12587 ( .A(n6294), .B(p_input[4336]), .Z(o[4336]) );
  AND U12588 ( .A(p_input[24336]), .B(p_input[14336]), .Z(n6294) );
  AND U12589 ( .A(n6295), .B(p_input[4335]), .Z(o[4335]) );
  AND U12590 ( .A(p_input[24335]), .B(p_input[14335]), .Z(n6295) );
  AND U12591 ( .A(n6296), .B(p_input[4334]), .Z(o[4334]) );
  AND U12592 ( .A(p_input[24334]), .B(p_input[14334]), .Z(n6296) );
  AND U12593 ( .A(n6297), .B(p_input[4333]), .Z(o[4333]) );
  AND U12594 ( .A(p_input[24333]), .B(p_input[14333]), .Z(n6297) );
  AND U12595 ( .A(n6298), .B(p_input[4332]), .Z(o[4332]) );
  AND U12596 ( .A(p_input[24332]), .B(p_input[14332]), .Z(n6298) );
  AND U12597 ( .A(n6299), .B(p_input[4331]), .Z(o[4331]) );
  AND U12598 ( .A(p_input[24331]), .B(p_input[14331]), .Z(n6299) );
  AND U12599 ( .A(n6300), .B(p_input[4330]), .Z(o[4330]) );
  AND U12600 ( .A(p_input[24330]), .B(p_input[14330]), .Z(n6300) );
  AND U12601 ( .A(n6301), .B(p_input[432]), .Z(o[432]) );
  AND U12602 ( .A(p_input[20432]), .B(p_input[10432]), .Z(n6301) );
  AND U12603 ( .A(n6302), .B(p_input[4329]), .Z(o[4329]) );
  AND U12604 ( .A(p_input[24329]), .B(p_input[14329]), .Z(n6302) );
  AND U12605 ( .A(n6303), .B(p_input[4328]), .Z(o[4328]) );
  AND U12606 ( .A(p_input[24328]), .B(p_input[14328]), .Z(n6303) );
  AND U12607 ( .A(n6304), .B(p_input[4327]), .Z(o[4327]) );
  AND U12608 ( .A(p_input[24327]), .B(p_input[14327]), .Z(n6304) );
  AND U12609 ( .A(n6305), .B(p_input[4326]), .Z(o[4326]) );
  AND U12610 ( .A(p_input[24326]), .B(p_input[14326]), .Z(n6305) );
  AND U12611 ( .A(n6306), .B(p_input[4325]), .Z(o[4325]) );
  AND U12612 ( .A(p_input[24325]), .B(p_input[14325]), .Z(n6306) );
  AND U12613 ( .A(n6307), .B(p_input[4324]), .Z(o[4324]) );
  AND U12614 ( .A(p_input[24324]), .B(p_input[14324]), .Z(n6307) );
  AND U12615 ( .A(n6308), .B(p_input[4323]), .Z(o[4323]) );
  AND U12616 ( .A(p_input[24323]), .B(p_input[14323]), .Z(n6308) );
  AND U12617 ( .A(n6309), .B(p_input[4322]), .Z(o[4322]) );
  AND U12618 ( .A(p_input[24322]), .B(p_input[14322]), .Z(n6309) );
  AND U12619 ( .A(n6310), .B(p_input[4321]), .Z(o[4321]) );
  AND U12620 ( .A(p_input[24321]), .B(p_input[14321]), .Z(n6310) );
  AND U12621 ( .A(n6311), .B(p_input[4320]), .Z(o[4320]) );
  AND U12622 ( .A(p_input[24320]), .B(p_input[14320]), .Z(n6311) );
  AND U12623 ( .A(n6312), .B(p_input[431]), .Z(o[431]) );
  AND U12624 ( .A(p_input[20431]), .B(p_input[10431]), .Z(n6312) );
  AND U12625 ( .A(n6313), .B(p_input[4319]), .Z(o[4319]) );
  AND U12626 ( .A(p_input[24319]), .B(p_input[14319]), .Z(n6313) );
  AND U12627 ( .A(n6314), .B(p_input[4318]), .Z(o[4318]) );
  AND U12628 ( .A(p_input[24318]), .B(p_input[14318]), .Z(n6314) );
  AND U12629 ( .A(n6315), .B(p_input[4317]), .Z(o[4317]) );
  AND U12630 ( .A(p_input[24317]), .B(p_input[14317]), .Z(n6315) );
  AND U12631 ( .A(n6316), .B(p_input[4316]), .Z(o[4316]) );
  AND U12632 ( .A(p_input[24316]), .B(p_input[14316]), .Z(n6316) );
  AND U12633 ( .A(n6317), .B(p_input[4315]), .Z(o[4315]) );
  AND U12634 ( .A(p_input[24315]), .B(p_input[14315]), .Z(n6317) );
  AND U12635 ( .A(n6318), .B(p_input[4314]), .Z(o[4314]) );
  AND U12636 ( .A(p_input[24314]), .B(p_input[14314]), .Z(n6318) );
  AND U12637 ( .A(n6319), .B(p_input[4313]), .Z(o[4313]) );
  AND U12638 ( .A(p_input[24313]), .B(p_input[14313]), .Z(n6319) );
  AND U12639 ( .A(n6320), .B(p_input[4312]), .Z(o[4312]) );
  AND U12640 ( .A(p_input[24312]), .B(p_input[14312]), .Z(n6320) );
  AND U12641 ( .A(n6321), .B(p_input[4311]), .Z(o[4311]) );
  AND U12642 ( .A(p_input[24311]), .B(p_input[14311]), .Z(n6321) );
  AND U12643 ( .A(n6322), .B(p_input[4310]), .Z(o[4310]) );
  AND U12644 ( .A(p_input[24310]), .B(p_input[14310]), .Z(n6322) );
  AND U12645 ( .A(n6323), .B(p_input[430]), .Z(o[430]) );
  AND U12646 ( .A(p_input[20430]), .B(p_input[10430]), .Z(n6323) );
  AND U12647 ( .A(n6324), .B(p_input[4309]), .Z(o[4309]) );
  AND U12648 ( .A(p_input[24309]), .B(p_input[14309]), .Z(n6324) );
  AND U12649 ( .A(n6325), .B(p_input[4308]), .Z(o[4308]) );
  AND U12650 ( .A(p_input[24308]), .B(p_input[14308]), .Z(n6325) );
  AND U12651 ( .A(n6326), .B(p_input[4307]), .Z(o[4307]) );
  AND U12652 ( .A(p_input[24307]), .B(p_input[14307]), .Z(n6326) );
  AND U12653 ( .A(n6327), .B(p_input[4306]), .Z(o[4306]) );
  AND U12654 ( .A(p_input[24306]), .B(p_input[14306]), .Z(n6327) );
  AND U12655 ( .A(n6328), .B(p_input[4305]), .Z(o[4305]) );
  AND U12656 ( .A(p_input[24305]), .B(p_input[14305]), .Z(n6328) );
  AND U12657 ( .A(n6329), .B(p_input[4304]), .Z(o[4304]) );
  AND U12658 ( .A(p_input[24304]), .B(p_input[14304]), .Z(n6329) );
  AND U12659 ( .A(n6330), .B(p_input[4303]), .Z(o[4303]) );
  AND U12660 ( .A(p_input[24303]), .B(p_input[14303]), .Z(n6330) );
  AND U12661 ( .A(n6331), .B(p_input[4302]), .Z(o[4302]) );
  AND U12662 ( .A(p_input[24302]), .B(p_input[14302]), .Z(n6331) );
  AND U12663 ( .A(n6332), .B(p_input[4301]), .Z(o[4301]) );
  AND U12664 ( .A(p_input[24301]), .B(p_input[14301]), .Z(n6332) );
  AND U12665 ( .A(n6333), .B(p_input[4300]), .Z(o[4300]) );
  AND U12666 ( .A(p_input[24300]), .B(p_input[14300]), .Z(n6333) );
  AND U12667 ( .A(n6334), .B(p_input[42]), .Z(o[42]) );
  AND U12668 ( .A(p_input[20042]), .B(p_input[10042]), .Z(n6334) );
  AND U12669 ( .A(n6335), .B(p_input[429]), .Z(o[429]) );
  AND U12670 ( .A(p_input[20429]), .B(p_input[10429]), .Z(n6335) );
  AND U12671 ( .A(n6336), .B(p_input[4299]), .Z(o[4299]) );
  AND U12672 ( .A(p_input[24299]), .B(p_input[14299]), .Z(n6336) );
  AND U12673 ( .A(n6337), .B(p_input[4298]), .Z(o[4298]) );
  AND U12674 ( .A(p_input[24298]), .B(p_input[14298]), .Z(n6337) );
  AND U12675 ( .A(n6338), .B(p_input[4297]), .Z(o[4297]) );
  AND U12676 ( .A(p_input[24297]), .B(p_input[14297]), .Z(n6338) );
  AND U12677 ( .A(n6339), .B(p_input[4296]), .Z(o[4296]) );
  AND U12678 ( .A(p_input[24296]), .B(p_input[14296]), .Z(n6339) );
  AND U12679 ( .A(n6340), .B(p_input[4295]), .Z(o[4295]) );
  AND U12680 ( .A(p_input[24295]), .B(p_input[14295]), .Z(n6340) );
  AND U12681 ( .A(n6341), .B(p_input[4294]), .Z(o[4294]) );
  AND U12682 ( .A(p_input[24294]), .B(p_input[14294]), .Z(n6341) );
  AND U12683 ( .A(n6342), .B(p_input[4293]), .Z(o[4293]) );
  AND U12684 ( .A(p_input[24293]), .B(p_input[14293]), .Z(n6342) );
  AND U12685 ( .A(n6343), .B(p_input[4292]), .Z(o[4292]) );
  AND U12686 ( .A(p_input[24292]), .B(p_input[14292]), .Z(n6343) );
  AND U12687 ( .A(n6344), .B(p_input[4291]), .Z(o[4291]) );
  AND U12688 ( .A(p_input[24291]), .B(p_input[14291]), .Z(n6344) );
  AND U12689 ( .A(n6345), .B(p_input[4290]), .Z(o[4290]) );
  AND U12690 ( .A(p_input[24290]), .B(p_input[14290]), .Z(n6345) );
  AND U12691 ( .A(n6346), .B(p_input[428]), .Z(o[428]) );
  AND U12692 ( .A(p_input[20428]), .B(p_input[10428]), .Z(n6346) );
  AND U12693 ( .A(n6347), .B(p_input[4289]), .Z(o[4289]) );
  AND U12694 ( .A(p_input[24289]), .B(p_input[14289]), .Z(n6347) );
  AND U12695 ( .A(n6348), .B(p_input[4288]), .Z(o[4288]) );
  AND U12696 ( .A(p_input[24288]), .B(p_input[14288]), .Z(n6348) );
  AND U12697 ( .A(n6349), .B(p_input[4287]), .Z(o[4287]) );
  AND U12698 ( .A(p_input[24287]), .B(p_input[14287]), .Z(n6349) );
  AND U12699 ( .A(n6350), .B(p_input[4286]), .Z(o[4286]) );
  AND U12700 ( .A(p_input[24286]), .B(p_input[14286]), .Z(n6350) );
  AND U12701 ( .A(n6351), .B(p_input[4285]), .Z(o[4285]) );
  AND U12702 ( .A(p_input[24285]), .B(p_input[14285]), .Z(n6351) );
  AND U12703 ( .A(n6352), .B(p_input[4284]), .Z(o[4284]) );
  AND U12704 ( .A(p_input[24284]), .B(p_input[14284]), .Z(n6352) );
  AND U12705 ( .A(n6353), .B(p_input[4283]), .Z(o[4283]) );
  AND U12706 ( .A(p_input[24283]), .B(p_input[14283]), .Z(n6353) );
  AND U12707 ( .A(n6354), .B(p_input[4282]), .Z(o[4282]) );
  AND U12708 ( .A(p_input[24282]), .B(p_input[14282]), .Z(n6354) );
  AND U12709 ( .A(n6355), .B(p_input[4281]), .Z(o[4281]) );
  AND U12710 ( .A(p_input[24281]), .B(p_input[14281]), .Z(n6355) );
  AND U12711 ( .A(n6356), .B(p_input[4280]), .Z(o[4280]) );
  AND U12712 ( .A(p_input[24280]), .B(p_input[14280]), .Z(n6356) );
  AND U12713 ( .A(n6357), .B(p_input[427]), .Z(o[427]) );
  AND U12714 ( .A(p_input[20427]), .B(p_input[10427]), .Z(n6357) );
  AND U12715 ( .A(n6358), .B(p_input[4279]), .Z(o[4279]) );
  AND U12716 ( .A(p_input[24279]), .B(p_input[14279]), .Z(n6358) );
  AND U12717 ( .A(n6359), .B(p_input[4278]), .Z(o[4278]) );
  AND U12718 ( .A(p_input[24278]), .B(p_input[14278]), .Z(n6359) );
  AND U12719 ( .A(n6360), .B(p_input[4277]), .Z(o[4277]) );
  AND U12720 ( .A(p_input[24277]), .B(p_input[14277]), .Z(n6360) );
  AND U12721 ( .A(n6361), .B(p_input[4276]), .Z(o[4276]) );
  AND U12722 ( .A(p_input[24276]), .B(p_input[14276]), .Z(n6361) );
  AND U12723 ( .A(n6362), .B(p_input[4275]), .Z(o[4275]) );
  AND U12724 ( .A(p_input[24275]), .B(p_input[14275]), .Z(n6362) );
  AND U12725 ( .A(n6363), .B(p_input[4274]), .Z(o[4274]) );
  AND U12726 ( .A(p_input[24274]), .B(p_input[14274]), .Z(n6363) );
  AND U12727 ( .A(n6364), .B(p_input[4273]), .Z(o[4273]) );
  AND U12728 ( .A(p_input[24273]), .B(p_input[14273]), .Z(n6364) );
  AND U12729 ( .A(n6365), .B(p_input[4272]), .Z(o[4272]) );
  AND U12730 ( .A(p_input[24272]), .B(p_input[14272]), .Z(n6365) );
  AND U12731 ( .A(n6366), .B(p_input[4271]), .Z(o[4271]) );
  AND U12732 ( .A(p_input[24271]), .B(p_input[14271]), .Z(n6366) );
  AND U12733 ( .A(n6367), .B(p_input[4270]), .Z(o[4270]) );
  AND U12734 ( .A(p_input[24270]), .B(p_input[14270]), .Z(n6367) );
  AND U12735 ( .A(n6368), .B(p_input[426]), .Z(o[426]) );
  AND U12736 ( .A(p_input[20426]), .B(p_input[10426]), .Z(n6368) );
  AND U12737 ( .A(n6369), .B(p_input[4269]), .Z(o[4269]) );
  AND U12738 ( .A(p_input[24269]), .B(p_input[14269]), .Z(n6369) );
  AND U12739 ( .A(n6370), .B(p_input[4268]), .Z(o[4268]) );
  AND U12740 ( .A(p_input[24268]), .B(p_input[14268]), .Z(n6370) );
  AND U12741 ( .A(n6371), .B(p_input[4267]), .Z(o[4267]) );
  AND U12742 ( .A(p_input[24267]), .B(p_input[14267]), .Z(n6371) );
  AND U12743 ( .A(n6372), .B(p_input[4266]), .Z(o[4266]) );
  AND U12744 ( .A(p_input[24266]), .B(p_input[14266]), .Z(n6372) );
  AND U12745 ( .A(n6373), .B(p_input[4265]), .Z(o[4265]) );
  AND U12746 ( .A(p_input[24265]), .B(p_input[14265]), .Z(n6373) );
  AND U12747 ( .A(n6374), .B(p_input[4264]), .Z(o[4264]) );
  AND U12748 ( .A(p_input[24264]), .B(p_input[14264]), .Z(n6374) );
  AND U12749 ( .A(n6375), .B(p_input[4263]), .Z(o[4263]) );
  AND U12750 ( .A(p_input[24263]), .B(p_input[14263]), .Z(n6375) );
  AND U12751 ( .A(n6376), .B(p_input[4262]), .Z(o[4262]) );
  AND U12752 ( .A(p_input[24262]), .B(p_input[14262]), .Z(n6376) );
  AND U12753 ( .A(n6377), .B(p_input[4261]), .Z(o[4261]) );
  AND U12754 ( .A(p_input[24261]), .B(p_input[14261]), .Z(n6377) );
  AND U12755 ( .A(n6378), .B(p_input[4260]), .Z(o[4260]) );
  AND U12756 ( .A(p_input[24260]), .B(p_input[14260]), .Z(n6378) );
  AND U12757 ( .A(n6379), .B(p_input[425]), .Z(o[425]) );
  AND U12758 ( .A(p_input[20425]), .B(p_input[10425]), .Z(n6379) );
  AND U12759 ( .A(n6380), .B(p_input[4259]), .Z(o[4259]) );
  AND U12760 ( .A(p_input[24259]), .B(p_input[14259]), .Z(n6380) );
  AND U12761 ( .A(n6381), .B(p_input[4258]), .Z(o[4258]) );
  AND U12762 ( .A(p_input[24258]), .B(p_input[14258]), .Z(n6381) );
  AND U12763 ( .A(n6382), .B(p_input[4257]), .Z(o[4257]) );
  AND U12764 ( .A(p_input[24257]), .B(p_input[14257]), .Z(n6382) );
  AND U12765 ( .A(n6383), .B(p_input[4256]), .Z(o[4256]) );
  AND U12766 ( .A(p_input[24256]), .B(p_input[14256]), .Z(n6383) );
  AND U12767 ( .A(n6384), .B(p_input[4255]), .Z(o[4255]) );
  AND U12768 ( .A(p_input[24255]), .B(p_input[14255]), .Z(n6384) );
  AND U12769 ( .A(n6385), .B(p_input[4254]), .Z(o[4254]) );
  AND U12770 ( .A(p_input[24254]), .B(p_input[14254]), .Z(n6385) );
  AND U12771 ( .A(n6386), .B(p_input[4253]), .Z(o[4253]) );
  AND U12772 ( .A(p_input[24253]), .B(p_input[14253]), .Z(n6386) );
  AND U12773 ( .A(n6387), .B(p_input[4252]), .Z(o[4252]) );
  AND U12774 ( .A(p_input[24252]), .B(p_input[14252]), .Z(n6387) );
  AND U12775 ( .A(n6388), .B(p_input[4251]), .Z(o[4251]) );
  AND U12776 ( .A(p_input[24251]), .B(p_input[14251]), .Z(n6388) );
  AND U12777 ( .A(n6389), .B(p_input[4250]), .Z(o[4250]) );
  AND U12778 ( .A(p_input[24250]), .B(p_input[14250]), .Z(n6389) );
  AND U12779 ( .A(n6390), .B(p_input[424]), .Z(o[424]) );
  AND U12780 ( .A(p_input[20424]), .B(p_input[10424]), .Z(n6390) );
  AND U12781 ( .A(n6391), .B(p_input[4249]), .Z(o[4249]) );
  AND U12782 ( .A(p_input[24249]), .B(p_input[14249]), .Z(n6391) );
  AND U12783 ( .A(n6392), .B(p_input[4248]), .Z(o[4248]) );
  AND U12784 ( .A(p_input[24248]), .B(p_input[14248]), .Z(n6392) );
  AND U12785 ( .A(n6393), .B(p_input[4247]), .Z(o[4247]) );
  AND U12786 ( .A(p_input[24247]), .B(p_input[14247]), .Z(n6393) );
  AND U12787 ( .A(n6394), .B(p_input[4246]), .Z(o[4246]) );
  AND U12788 ( .A(p_input[24246]), .B(p_input[14246]), .Z(n6394) );
  AND U12789 ( .A(n6395), .B(p_input[4245]), .Z(o[4245]) );
  AND U12790 ( .A(p_input[24245]), .B(p_input[14245]), .Z(n6395) );
  AND U12791 ( .A(n6396), .B(p_input[4244]), .Z(o[4244]) );
  AND U12792 ( .A(p_input[24244]), .B(p_input[14244]), .Z(n6396) );
  AND U12793 ( .A(n6397), .B(p_input[4243]), .Z(o[4243]) );
  AND U12794 ( .A(p_input[24243]), .B(p_input[14243]), .Z(n6397) );
  AND U12795 ( .A(n6398), .B(p_input[4242]), .Z(o[4242]) );
  AND U12796 ( .A(p_input[24242]), .B(p_input[14242]), .Z(n6398) );
  AND U12797 ( .A(n6399), .B(p_input[4241]), .Z(o[4241]) );
  AND U12798 ( .A(p_input[24241]), .B(p_input[14241]), .Z(n6399) );
  AND U12799 ( .A(n6400), .B(p_input[4240]), .Z(o[4240]) );
  AND U12800 ( .A(p_input[24240]), .B(p_input[14240]), .Z(n6400) );
  AND U12801 ( .A(n6401), .B(p_input[423]), .Z(o[423]) );
  AND U12802 ( .A(p_input[20423]), .B(p_input[10423]), .Z(n6401) );
  AND U12803 ( .A(n6402), .B(p_input[4239]), .Z(o[4239]) );
  AND U12804 ( .A(p_input[24239]), .B(p_input[14239]), .Z(n6402) );
  AND U12805 ( .A(n6403), .B(p_input[4238]), .Z(o[4238]) );
  AND U12806 ( .A(p_input[24238]), .B(p_input[14238]), .Z(n6403) );
  AND U12807 ( .A(n6404), .B(p_input[4237]), .Z(o[4237]) );
  AND U12808 ( .A(p_input[24237]), .B(p_input[14237]), .Z(n6404) );
  AND U12809 ( .A(n6405), .B(p_input[4236]), .Z(o[4236]) );
  AND U12810 ( .A(p_input[24236]), .B(p_input[14236]), .Z(n6405) );
  AND U12811 ( .A(n6406), .B(p_input[4235]), .Z(o[4235]) );
  AND U12812 ( .A(p_input[24235]), .B(p_input[14235]), .Z(n6406) );
  AND U12813 ( .A(n6407), .B(p_input[4234]), .Z(o[4234]) );
  AND U12814 ( .A(p_input[24234]), .B(p_input[14234]), .Z(n6407) );
  AND U12815 ( .A(n6408), .B(p_input[4233]), .Z(o[4233]) );
  AND U12816 ( .A(p_input[24233]), .B(p_input[14233]), .Z(n6408) );
  AND U12817 ( .A(n6409), .B(p_input[4232]), .Z(o[4232]) );
  AND U12818 ( .A(p_input[24232]), .B(p_input[14232]), .Z(n6409) );
  AND U12819 ( .A(n6410), .B(p_input[4231]), .Z(o[4231]) );
  AND U12820 ( .A(p_input[24231]), .B(p_input[14231]), .Z(n6410) );
  AND U12821 ( .A(n6411), .B(p_input[4230]), .Z(o[4230]) );
  AND U12822 ( .A(p_input[24230]), .B(p_input[14230]), .Z(n6411) );
  AND U12823 ( .A(n6412), .B(p_input[422]), .Z(o[422]) );
  AND U12824 ( .A(p_input[20422]), .B(p_input[10422]), .Z(n6412) );
  AND U12825 ( .A(n6413), .B(p_input[4229]), .Z(o[4229]) );
  AND U12826 ( .A(p_input[24229]), .B(p_input[14229]), .Z(n6413) );
  AND U12827 ( .A(n6414), .B(p_input[4228]), .Z(o[4228]) );
  AND U12828 ( .A(p_input[24228]), .B(p_input[14228]), .Z(n6414) );
  AND U12829 ( .A(n6415), .B(p_input[4227]), .Z(o[4227]) );
  AND U12830 ( .A(p_input[24227]), .B(p_input[14227]), .Z(n6415) );
  AND U12831 ( .A(n6416), .B(p_input[4226]), .Z(o[4226]) );
  AND U12832 ( .A(p_input[24226]), .B(p_input[14226]), .Z(n6416) );
  AND U12833 ( .A(n6417), .B(p_input[4225]), .Z(o[4225]) );
  AND U12834 ( .A(p_input[24225]), .B(p_input[14225]), .Z(n6417) );
  AND U12835 ( .A(n6418), .B(p_input[4224]), .Z(o[4224]) );
  AND U12836 ( .A(p_input[24224]), .B(p_input[14224]), .Z(n6418) );
  AND U12837 ( .A(n6419), .B(p_input[4223]), .Z(o[4223]) );
  AND U12838 ( .A(p_input[24223]), .B(p_input[14223]), .Z(n6419) );
  AND U12839 ( .A(n6420), .B(p_input[4222]), .Z(o[4222]) );
  AND U12840 ( .A(p_input[24222]), .B(p_input[14222]), .Z(n6420) );
  AND U12841 ( .A(n6421), .B(p_input[4221]), .Z(o[4221]) );
  AND U12842 ( .A(p_input[24221]), .B(p_input[14221]), .Z(n6421) );
  AND U12843 ( .A(n6422), .B(p_input[4220]), .Z(o[4220]) );
  AND U12844 ( .A(p_input[24220]), .B(p_input[14220]), .Z(n6422) );
  AND U12845 ( .A(n6423), .B(p_input[421]), .Z(o[421]) );
  AND U12846 ( .A(p_input[20421]), .B(p_input[10421]), .Z(n6423) );
  AND U12847 ( .A(n6424), .B(p_input[4219]), .Z(o[4219]) );
  AND U12848 ( .A(p_input[24219]), .B(p_input[14219]), .Z(n6424) );
  AND U12849 ( .A(n6425), .B(p_input[4218]), .Z(o[4218]) );
  AND U12850 ( .A(p_input[24218]), .B(p_input[14218]), .Z(n6425) );
  AND U12851 ( .A(n6426), .B(p_input[4217]), .Z(o[4217]) );
  AND U12852 ( .A(p_input[24217]), .B(p_input[14217]), .Z(n6426) );
  AND U12853 ( .A(n6427), .B(p_input[4216]), .Z(o[4216]) );
  AND U12854 ( .A(p_input[24216]), .B(p_input[14216]), .Z(n6427) );
  AND U12855 ( .A(n6428), .B(p_input[4215]), .Z(o[4215]) );
  AND U12856 ( .A(p_input[24215]), .B(p_input[14215]), .Z(n6428) );
  AND U12857 ( .A(n6429), .B(p_input[4214]), .Z(o[4214]) );
  AND U12858 ( .A(p_input[24214]), .B(p_input[14214]), .Z(n6429) );
  AND U12859 ( .A(n6430), .B(p_input[4213]), .Z(o[4213]) );
  AND U12860 ( .A(p_input[24213]), .B(p_input[14213]), .Z(n6430) );
  AND U12861 ( .A(n6431), .B(p_input[4212]), .Z(o[4212]) );
  AND U12862 ( .A(p_input[24212]), .B(p_input[14212]), .Z(n6431) );
  AND U12863 ( .A(n6432), .B(p_input[4211]), .Z(o[4211]) );
  AND U12864 ( .A(p_input[24211]), .B(p_input[14211]), .Z(n6432) );
  AND U12865 ( .A(n6433), .B(p_input[4210]), .Z(o[4210]) );
  AND U12866 ( .A(p_input[24210]), .B(p_input[14210]), .Z(n6433) );
  AND U12867 ( .A(n6434), .B(p_input[420]), .Z(o[420]) );
  AND U12868 ( .A(p_input[20420]), .B(p_input[10420]), .Z(n6434) );
  AND U12869 ( .A(n6435), .B(p_input[4209]), .Z(o[4209]) );
  AND U12870 ( .A(p_input[24209]), .B(p_input[14209]), .Z(n6435) );
  AND U12871 ( .A(n6436), .B(p_input[4208]), .Z(o[4208]) );
  AND U12872 ( .A(p_input[24208]), .B(p_input[14208]), .Z(n6436) );
  AND U12873 ( .A(n6437), .B(p_input[4207]), .Z(o[4207]) );
  AND U12874 ( .A(p_input[24207]), .B(p_input[14207]), .Z(n6437) );
  AND U12875 ( .A(n6438), .B(p_input[4206]), .Z(o[4206]) );
  AND U12876 ( .A(p_input[24206]), .B(p_input[14206]), .Z(n6438) );
  AND U12877 ( .A(n6439), .B(p_input[4205]), .Z(o[4205]) );
  AND U12878 ( .A(p_input[24205]), .B(p_input[14205]), .Z(n6439) );
  AND U12879 ( .A(n6440), .B(p_input[4204]), .Z(o[4204]) );
  AND U12880 ( .A(p_input[24204]), .B(p_input[14204]), .Z(n6440) );
  AND U12881 ( .A(n6441), .B(p_input[4203]), .Z(o[4203]) );
  AND U12882 ( .A(p_input[24203]), .B(p_input[14203]), .Z(n6441) );
  AND U12883 ( .A(n6442), .B(p_input[4202]), .Z(o[4202]) );
  AND U12884 ( .A(p_input[24202]), .B(p_input[14202]), .Z(n6442) );
  AND U12885 ( .A(n6443), .B(p_input[4201]), .Z(o[4201]) );
  AND U12886 ( .A(p_input[24201]), .B(p_input[14201]), .Z(n6443) );
  AND U12887 ( .A(n6444), .B(p_input[4200]), .Z(o[4200]) );
  AND U12888 ( .A(p_input[24200]), .B(p_input[14200]), .Z(n6444) );
  AND U12889 ( .A(n6445), .B(p_input[41]), .Z(o[41]) );
  AND U12890 ( .A(p_input[20041]), .B(p_input[10041]), .Z(n6445) );
  AND U12891 ( .A(n6446), .B(p_input[419]), .Z(o[419]) );
  AND U12892 ( .A(p_input[20419]), .B(p_input[10419]), .Z(n6446) );
  AND U12893 ( .A(n6447), .B(p_input[4199]), .Z(o[4199]) );
  AND U12894 ( .A(p_input[24199]), .B(p_input[14199]), .Z(n6447) );
  AND U12895 ( .A(n6448), .B(p_input[4198]), .Z(o[4198]) );
  AND U12896 ( .A(p_input[24198]), .B(p_input[14198]), .Z(n6448) );
  AND U12897 ( .A(n6449), .B(p_input[4197]), .Z(o[4197]) );
  AND U12898 ( .A(p_input[24197]), .B(p_input[14197]), .Z(n6449) );
  AND U12899 ( .A(n6450), .B(p_input[4196]), .Z(o[4196]) );
  AND U12900 ( .A(p_input[24196]), .B(p_input[14196]), .Z(n6450) );
  AND U12901 ( .A(n6451), .B(p_input[4195]), .Z(o[4195]) );
  AND U12902 ( .A(p_input[24195]), .B(p_input[14195]), .Z(n6451) );
  AND U12903 ( .A(n6452), .B(p_input[4194]), .Z(o[4194]) );
  AND U12904 ( .A(p_input[24194]), .B(p_input[14194]), .Z(n6452) );
  AND U12905 ( .A(n6453), .B(p_input[4193]), .Z(o[4193]) );
  AND U12906 ( .A(p_input[24193]), .B(p_input[14193]), .Z(n6453) );
  AND U12907 ( .A(n6454), .B(p_input[4192]), .Z(o[4192]) );
  AND U12908 ( .A(p_input[24192]), .B(p_input[14192]), .Z(n6454) );
  AND U12909 ( .A(n6455), .B(p_input[4191]), .Z(o[4191]) );
  AND U12910 ( .A(p_input[24191]), .B(p_input[14191]), .Z(n6455) );
  AND U12911 ( .A(n6456), .B(p_input[4190]), .Z(o[4190]) );
  AND U12912 ( .A(p_input[24190]), .B(p_input[14190]), .Z(n6456) );
  AND U12913 ( .A(n6457), .B(p_input[418]), .Z(o[418]) );
  AND U12914 ( .A(p_input[20418]), .B(p_input[10418]), .Z(n6457) );
  AND U12915 ( .A(n6458), .B(p_input[4189]), .Z(o[4189]) );
  AND U12916 ( .A(p_input[24189]), .B(p_input[14189]), .Z(n6458) );
  AND U12917 ( .A(n6459), .B(p_input[4188]), .Z(o[4188]) );
  AND U12918 ( .A(p_input[24188]), .B(p_input[14188]), .Z(n6459) );
  AND U12919 ( .A(n6460), .B(p_input[4187]), .Z(o[4187]) );
  AND U12920 ( .A(p_input[24187]), .B(p_input[14187]), .Z(n6460) );
  AND U12921 ( .A(n6461), .B(p_input[4186]), .Z(o[4186]) );
  AND U12922 ( .A(p_input[24186]), .B(p_input[14186]), .Z(n6461) );
  AND U12923 ( .A(n6462), .B(p_input[4185]), .Z(o[4185]) );
  AND U12924 ( .A(p_input[24185]), .B(p_input[14185]), .Z(n6462) );
  AND U12925 ( .A(n6463), .B(p_input[4184]), .Z(o[4184]) );
  AND U12926 ( .A(p_input[24184]), .B(p_input[14184]), .Z(n6463) );
  AND U12927 ( .A(n6464), .B(p_input[4183]), .Z(o[4183]) );
  AND U12928 ( .A(p_input[24183]), .B(p_input[14183]), .Z(n6464) );
  AND U12929 ( .A(n6465), .B(p_input[4182]), .Z(o[4182]) );
  AND U12930 ( .A(p_input[24182]), .B(p_input[14182]), .Z(n6465) );
  AND U12931 ( .A(n6466), .B(p_input[4181]), .Z(o[4181]) );
  AND U12932 ( .A(p_input[24181]), .B(p_input[14181]), .Z(n6466) );
  AND U12933 ( .A(n6467), .B(p_input[4180]), .Z(o[4180]) );
  AND U12934 ( .A(p_input[24180]), .B(p_input[14180]), .Z(n6467) );
  AND U12935 ( .A(n6468), .B(p_input[417]), .Z(o[417]) );
  AND U12936 ( .A(p_input[20417]), .B(p_input[10417]), .Z(n6468) );
  AND U12937 ( .A(n6469), .B(p_input[4179]), .Z(o[4179]) );
  AND U12938 ( .A(p_input[24179]), .B(p_input[14179]), .Z(n6469) );
  AND U12939 ( .A(n6470), .B(p_input[4178]), .Z(o[4178]) );
  AND U12940 ( .A(p_input[24178]), .B(p_input[14178]), .Z(n6470) );
  AND U12941 ( .A(n6471), .B(p_input[4177]), .Z(o[4177]) );
  AND U12942 ( .A(p_input[24177]), .B(p_input[14177]), .Z(n6471) );
  AND U12943 ( .A(n6472), .B(p_input[4176]), .Z(o[4176]) );
  AND U12944 ( .A(p_input[24176]), .B(p_input[14176]), .Z(n6472) );
  AND U12945 ( .A(n6473), .B(p_input[4175]), .Z(o[4175]) );
  AND U12946 ( .A(p_input[24175]), .B(p_input[14175]), .Z(n6473) );
  AND U12947 ( .A(n6474), .B(p_input[4174]), .Z(o[4174]) );
  AND U12948 ( .A(p_input[24174]), .B(p_input[14174]), .Z(n6474) );
  AND U12949 ( .A(n6475), .B(p_input[4173]), .Z(o[4173]) );
  AND U12950 ( .A(p_input[24173]), .B(p_input[14173]), .Z(n6475) );
  AND U12951 ( .A(n6476), .B(p_input[4172]), .Z(o[4172]) );
  AND U12952 ( .A(p_input[24172]), .B(p_input[14172]), .Z(n6476) );
  AND U12953 ( .A(n6477), .B(p_input[4171]), .Z(o[4171]) );
  AND U12954 ( .A(p_input[24171]), .B(p_input[14171]), .Z(n6477) );
  AND U12955 ( .A(n6478), .B(p_input[4170]), .Z(o[4170]) );
  AND U12956 ( .A(p_input[24170]), .B(p_input[14170]), .Z(n6478) );
  AND U12957 ( .A(n6479), .B(p_input[416]), .Z(o[416]) );
  AND U12958 ( .A(p_input[20416]), .B(p_input[10416]), .Z(n6479) );
  AND U12959 ( .A(n6480), .B(p_input[4169]), .Z(o[4169]) );
  AND U12960 ( .A(p_input[24169]), .B(p_input[14169]), .Z(n6480) );
  AND U12961 ( .A(n6481), .B(p_input[4168]), .Z(o[4168]) );
  AND U12962 ( .A(p_input[24168]), .B(p_input[14168]), .Z(n6481) );
  AND U12963 ( .A(n6482), .B(p_input[4167]), .Z(o[4167]) );
  AND U12964 ( .A(p_input[24167]), .B(p_input[14167]), .Z(n6482) );
  AND U12965 ( .A(n6483), .B(p_input[4166]), .Z(o[4166]) );
  AND U12966 ( .A(p_input[24166]), .B(p_input[14166]), .Z(n6483) );
  AND U12967 ( .A(n6484), .B(p_input[4165]), .Z(o[4165]) );
  AND U12968 ( .A(p_input[24165]), .B(p_input[14165]), .Z(n6484) );
  AND U12969 ( .A(n6485), .B(p_input[4164]), .Z(o[4164]) );
  AND U12970 ( .A(p_input[24164]), .B(p_input[14164]), .Z(n6485) );
  AND U12971 ( .A(n6486), .B(p_input[4163]), .Z(o[4163]) );
  AND U12972 ( .A(p_input[24163]), .B(p_input[14163]), .Z(n6486) );
  AND U12973 ( .A(n6487), .B(p_input[4162]), .Z(o[4162]) );
  AND U12974 ( .A(p_input[24162]), .B(p_input[14162]), .Z(n6487) );
  AND U12975 ( .A(n6488), .B(p_input[4161]), .Z(o[4161]) );
  AND U12976 ( .A(p_input[24161]), .B(p_input[14161]), .Z(n6488) );
  AND U12977 ( .A(n6489), .B(p_input[4160]), .Z(o[4160]) );
  AND U12978 ( .A(p_input[24160]), .B(p_input[14160]), .Z(n6489) );
  AND U12979 ( .A(n6490), .B(p_input[415]), .Z(o[415]) );
  AND U12980 ( .A(p_input[20415]), .B(p_input[10415]), .Z(n6490) );
  AND U12981 ( .A(n6491), .B(p_input[4159]), .Z(o[4159]) );
  AND U12982 ( .A(p_input[24159]), .B(p_input[14159]), .Z(n6491) );
  AND U12983 ( .A(n6492), .B(p_input[4158]), .Z(o[4158]) );
  AND U12984 ( .A(p_input[24158]), .B(p_input[14158]), .Z(n6492) );
  AND U12985 ( .A(n6493), .B(p_input[4157]), .Z(o[4157]) );
  AND U12986 ( .A(p_input[24157]), .B(p_input[14157]), .Z(n6493) );
  AND U12987 ( .A(n6494), .B(p_input[4156]), .Z(o[4156]) );
  AND U12988 ( .A(p_input[24156]), .B(p_input[14156]), .Z(n6494) );
  AND U12989 ( .A(n6495), .B(p_input[4155]), .Z(o[4155]) );
  AND U12990 ( .A(p_input[24155]), .B(p_input[14155]), .Z(n6495) );
  AND U12991 ( .A(n6496), .B(p_input[4154]), .Z(o[4154]) );
  AND U12992 ( .A(p_input[24154]), .B(p_input[14154]), .Z(n6496) );
  AND U12993 ( .A(n6497), .B(p_input[4153]), .Z(o[4153]) );
  AND U12994 ( .A(p_input[24153]), .B(p_input[14153]), .Z(n6497) );
  AND U12995 ( .A(n6498), .B(p_input[4152]), .Z(o[4152]) );
  AND U12996 ( .A(p_input[24152]), .B(p_input[14152]), .Z(n6498) );
  AND U12997 ( .A(n6499), .B(p_input[4151]), .Z(o[4151]) );
  AND U12998 ( .A(p_input[24151]), .B(p_input[14151]), .Z(n6499) );
  AND U12999 ( .A(n6500), .B(p_input[4150]), .Z(o[4150]) );
  AND U13000 ( .A(p_input[24150]), .B(p_input[14150]), .Z(n6500) );
  AND U13001 ( .A(n6501), .B(p_input[414]), .Z(o[414]) );
  AND U13002 ( .A(p_input[20414]), .B(p_input[10414]), .Z(n6501) );
  AND U13003 ( .A(n6502), .B(p_input[4149]), .Z(o[4149]) );
  AND U13004 ( .A(p_input[24149]), .B(p_input[14149]), .Z(n6502) );
  AND U13005 ( .A(n6503), .B(p_input[4148]), .Z(o[4148]) );
  AND U13006 ( .A(p_input[24148]), .B(p_input[14148]), .Z(n6503) );
  AND U13007 ( .A(n6504), .B(p_input[4147]), .Z(o[4147]) );
  AND U13008 ( .A(p_input[24147]), .B(p_input[14147]), .Z(n6504) );
  AND U13009 ( .A(n6505), .B(p_input[4146]), .Z(o[4146]) );
  AND U13010 ( .A(p_input[24146]), .B(p_input[14146]), .Z(n6505) );
  AND U13011 ( .A(n6506), .B(p_input[4145]), .Z(o[4145]) );
  AND U13012 ( .A(p_input[24145]), .B(p_input[14145]), .Z(n6506) );
  AND U13013 ( .A(n6507), .B(p_input[4144]), .Z(o[4144]) );
  AND U13014 ( .A(p_input[24144]), .B(p_input[14144]), .Z(n6507) );
  AND U13015 ( .A(n6508), .B(p_input[4143]), .Z(o[4143]) );
  AND U13016 ( .A(p_input[24143]), .B(p_input[14143]), .Z(n6508) );
  AND U13017 ( .A(n6509), .B(p_input[4142]), .Z(o[4142]) );
  AND U13018 ( .A(p_input[24142]), .B(p_input[14142]), .Z(n6509) );
  AND U13019 ( .A(n6510), .B(p_input[4141]), .Z(o[4141]) );
  AND U13020 ( .A(p_input[24141]), .B(p_input[14141]), .Z(n6510) );
  AND U13021 ( .A(n6511), .B(p_input[4140]), .Z(o[4140]) );
  AND U13022 ( .A(p_input[24140]), .B(p_input[14140]), .Z(n6511) );
  AND U13023 ( .A(n6512), .B(p_input[413]), .Z(o[413]) );
  AND U13024 ( .A(p_input[20413]), .B(p_input[10413]), .Z(n6512) );
  AND U13025 ( .A(n6513), .B(p_input[4139]), .Z(o[4139]) );
  AND U13026 ( .A(p_input[24139]), .B(p_input[14139]), .Z(n6513) );
  AND U13027 ( .A(n6514), .B(p_input[4138]), .Z(o[4138]) );
  AND U13028 ( .A(p_input[24138]), .B(p_input[14138]), .Z(n6514) );
  AND U13029 ( .A(n6515), .B(p_input[4137]), .Z(o[4137]) );
  AND U13030 ( .A(p_input[24137]), .B(p_input[14137]), .Z(n6515) );
  AND U13031 ( .A(n6516), .B(p_input[4136]), .Z(o[4136]) );
  AND U13032 ( .A(p_input[24136]), .B(p_input[14136]), .Z(n6516) );
  AND U13033 ( .A(n6517), .B(p_input[4135]), .Z(o[4135]) );
  AND U13034 ( .A(p_input[24135]), .B(p_input[14135]), .Z(n6517) );
  AND U13035 ( .A(n6518), .B(p_input[4134]), .Z(o[4134]) );
  AND U13036 ( .A(p_input[24134]), .B(p_input[14134]), .Z(n6518) );
  AND U13037 ( .A(n6519), .B(p_input[4133]), .Z(o[4133]) );
  AND U13038 ( .A(p_input[24133]), .B(p_input[14133]), .Z(n6519) );
  AND U13039 ( .A(n6520), .B(p_input[4132]), .Z(o[4132]) );
  AND U13040 ( .A(p_input[24132]), .B(p_input[14132]), .Z(n6520) );
  AND U13041 ( .A(n6521), .B(p_input[4131]), .Z(o[4131]) );
  AND U13042 ( .A(p_input[24131]), .B(p_input[14131]), .Z(n6521) );
  AND U13043 ( .A(n6522), .B(p_input[4130]), .Z(o[4130]) );
  AND U13044 ( .A(p_input[24130]), .B(p_input[14130]), .Z(n6522) );
  AND U13045 ( .A(n6523), .B(p_input[412]), .Z(o[412]) );
  AND U13046 ( .A(p_input[20412]), .B(p_input[10412]), .Z(n6523) );
  AND U13047 ( .A(n6524), .B(p_input[4129]), .Z(o[4129]) );
  AND U13048 ( .A(p_input[24129]), .B(p_input[14129]), .Z(n6524) );
  AND U13049 ( .A(n6525), .B(p_input[4128]), .Z(o[4128]) );
  AND U13050 ( .A(p_input[24128]), .B(p_input[14128]), .Z(n6525) );
  AND U13051 ( .A(n6526), .B(p_input[4127]), .Z(o[4127]) );
  AND U13052 ( .A(p_input[24127]), .B(p_input[14127]), .Z(n6526) );
  AND U13053 ( .A(n6527), .B(p_input[4126]), .Z(o[4126]) );
  AND U13054 ( .A(p_input[24126]), .B(p_input[14126]), .Z(n6527) );
  AND U13055 ( .A(n6528), .B(p_input[4125]), .Z(o[4125]) );
  AND U13056 ( .A(p_input[24125]), .B(p_input[14125]), .Z(n6528) );
  AND U13057 ( .A(n6529), .B(p_input[4124]), .Z(o[4124]) );
  AND U13058 ( .A(p_input[24124]), .B(p_input[14124]), .Z(n6529) );
  AND U13059 ( .A(n6530), .B(p_input[4123]), .Z(o[4123]) );
  AND U13060 ( .A(p_input[24123]), .B(p_input[14123]), .Z(n6530) );
  AND U13061 ( .A(n6531), .B(p_input[4122]), .Z(o[4122]) );
  AND U13062 ( .A(p_input[24122]), .B(p_input[14122]), .Z(n6531) );
  AND U13063 ( .A(n6532), .B(p_input[4121]), .Z(o[4121]) );
  AND U13064 ( .A(p_input[24121]), .B(p_input[14121]), .Z(n6532) );
  AND U13065 ( .A(n6533), .B(p_input[4120]), .Z(o[4120]) );
  AND U13066 ( .A(p_input[24120]), .B(p_input[14120]), .Z(n6533) );
  AND U13067 ( .A(n6534), .B(p_input[411]), .Z(o[411]) );
  AND U13068 ( .A(p_input[20411]), .B(p_input[10411]), .Z(n6534) );
  AND U13069 ( .A(n6535), .B(p_input[4119]), .Z(o[4119]) );
  AND U13070 ( .A(p_input[24119]), .B(p_input[14119]), .Z(n6535) );
  AND U13071 ( .A(n6536), .B(p_input[4118]), .Z(o[4118]) );
  AND U13072 ( .A(p_input[24118]), .B(p_input[14118]), .Z(n6536) );
  AND U13073 ( .A(n6537), .B(p_input[4117]), .Z(o[4117]) );
  AND U13074 ( .A(p_input[24117]), .B(p_input[14117]), .Z(n6537) );
  AND U13075 ( .A(n6538), .B(p_input[4116]), .Z(o[4116]) );
  AND U13076 ( .A(p_input[24116]), .B(p_input[14116]), .Z(n6538) );
  AND U13077 ( .A(n6539), .B(p_input[4115]), .Z(o[4115]) );
  AND U13078 ( .A(p_input[24115]), .B(p_input[14115]), .Z(n6539) );
  AND U13079 ( .A(n6540), .B(p_input[4114]), .Z(o[4114]) );
  AND U13080 ( .A(p_input[24114]), .B(p_input[14114]), .Z(n6540) );
  AND U13081 ( .A(n6541), .B(p_input[4113]), .Z(o[4113]) );
  AND U13082 ( .A(p_input[24113]), .B(p_input[14113]), .Z(n6541) );
  AND U13083 ( .A(n6542), .B(p_input[4112]), .Z(o[4112]) );
  AND U13084 ( .A(p_input[24112]), .B(p_input[14112]), .Z(n6542) );
  AND U13085 ( .A(n6543), .B(p_input[4111]), .Z(o[4111]) );
  AND U13086 ( .A(p_input[24111]), .B(p_input[14111]), .Z(n6543) );
  AND U13087 ( .A(n6544), .B(p_input[4110]), .Z(o[4110]) );
  AND U13088 ( .A(p_input[24110]), .B(p_input[14110]), .Z(n6544) );
  AND U13089 ( .A(n6545), .B(p_input[410]), .Z(o[410]) );
  AND U13090 ( .A(p_input[20410]), .B(p_input[10410]), .Z(n6545) );
  AND U13091 ( .A(n6546), .B(p_input[4109]), .Z(o[4109]) );
  AND U13092 ( .A(p_input[24109]), .B(p_input[14109]), .Z(n6546) );
  AND U13093 ( .A(n6547), .B(p_input[4108]), .Z(o[4108]) );
  AND U13094 ( .A(p_input[24108]), .B(p_input[14108]), .Z(n6547) );
  AND U13095 ( .A(n6548), .B(p_input[4107]), .Z(o[4107]) );
  AND U13096 ( .A(p_input[24107]), .B(p_input[14107]), .Z(n6548) );
  AND U13097 ( .A(n6549), .B(p_input[4106]), .Z(o[4106]) );
  AND U13098 ( .A(p_input[24106]), .B(p_input[14106]), .Z(n6549) );
  AND U13099 ( .A(n6550), .B(p_input[4105]), .Z(o[4105]) );
  AND U13100 ( .A(p_input[24105]), .B(p_input[14105]), .Z(n6550) );
  AND U13101 ( .A(n6551), .B(p_input[4104]), .Z(o[4104]) );
  AND U13102 ( .A(p_input[24104]), .B(p_input[14104]), .Z(n6551) );
  AND U13103 ( .A(n6552), .B(p_input[4103]), .Z(o[4103]) );
  AND U13104 ( .A(p_input[24103]), .B(p_input[14103]), .Z(n6552) );
  AND U13105 ( .A(n6553), .B(p_input[4102]), .Z(o[4102]) );
  AND U13106 ( .A(p_input[24102]), .B(p_input[14102]), .Z(n6553) );
  AND U13107 ( .A(n6554), .B(p_input[4101]), .Z(o[4101]) );
  AND U13108 ( .A(p_input[24101]), .B(p_input[14101]), .Z(n6554) );
  AND U13109 ( .A(n6555), .B(p_input[4100]), .Z(o[4100]) );
  AND U13110 ( .A(p_input[24100]), .B(p_input[14100]), .Z(n6555) );
  AND U13111 ( .A(n6556), .B(p_input[40]), .Z(o[40]) );
  AND U13112 ( .A(p_input[20040]), .B(p_input[10040]), .Z(n6556) );
  AND U13113 ( .A(n6557), .B(p_input[409]), .Z(o[409]) );
  AND U13114 ( .A(p_input[20409]), .B(p_input[10409]), .Z(n6557) );
  AND U13115 ( .A(n6558), .B(p_input[4099]), .Z(o[4099]) );
  AND U13116 ( .A(p_input[24099]), .B(p_input[14099]), .Z(n6558) );
  AND U13117 ( .A(n6559), .B(p_input[4098]), .Z(o[4098]) );
  AND U13118 ( .A(p_input[24098]), .B(p_input[14098]), .Z(n6559) );
  AND U13119 ( .A(n6560), .B(p_input[4097]), .Z(o[4097]) );
  AND U13120 ( .A(p_input[24097]), .B(p_input[14097]), .Z(n6560) );
  AND U13121 ( .A(n6561), .B(p_input[4096]), .Z(o[4096]) );
  AND U13122 ( .A(p_input[24096]), .B(p_input[14096]), .Z(n6561) );
  AND U13123 ( .A(n6562), .B(p_input[4095]), .Z(o[4095]) );
  AND U13124 ( .A(p_input[24095]), .B(p_input[14095]), .Z(n6562) );
  AND U13125 ( .A(n6563), .B(p_input[4094]), .Z(o[4094]) );
  AND U13126 ( .A(p_input[24094]), .B(p_input[14094]), .Z(n6563) );
  AND U13127 ( .A(n6564), .B(p_input[4093]), .Z(o[4093]) );
  AND U13128 ( .A(p_input[24093]), .B(p_input[14093]), .Z(n6564) );
  AND U13129 ( .A(n6565), .B(p_input[4092]), .Z(o[4092]) );
  AND U13130 ( .A(p_input[24092]), .B(p_input[14092]), .Z(n6565) );
  AND U13131 ( .A(n6566), .B(p_input[4091]), .Z(o[4091]) );
  AND U13132 ( .A(p_input[24091]), .B(p_input[14091]), .Z(n6566) );
  AND U13133 ( .A(n6567), .B(p_input[4090]), .Z(o[4090]) );
  AND U13134 ( .A(p_input[24090]), .B(p_input[14090]), .Z(n6567) );
  AND U13135 ( .A(n6568), .B(p_input[408]), .Z(o[408]) );
  AND U13136 ( .A(p_input[20408]), .B(p_input[10408]), .Z(n6568) );
  AND U13137 ( .A(n6569), .B(p_input[4089]), .Z(o[4089]) );
  AND U13138 ( .A(p_input[24089]), .B(p_input[14089]), .Z(n6569) );
  AND U13139 ( .A(n6570), .B(p_input[4088]), .Z(o[4088]) );
  AND U13140 ( .A(p_input[24088]), .B(p_input[14088]), .Z(n6570) );
  AND U13141 ( .A(n6571), .B(p_input[4087]), .Z(o[4087]) );
  AND U13142 ( .A(p_input[24087]), .B(p_input[14087]), .Z(n6571) );
  AND U13143 ( .A(n6572), .B(p_input[4086]), .Z(o[4086]) );
  AND U13144 ( .A(p_input[24086]), .B(p_input[14086]), .Z(n6572) );
  AND U13145 ( .A(n6573), .B(p_input[4085]), .Z(o[4085]) );
  AND U13146 ( .A(p_input[24085]), .B(p_input[14085]), .Z(n6573) );
  AND U13147 ( .A(n6574), .B(p_input[4084]), .Z(o[4084]) );
  AND U13148 ( .A(p_input[24084]), .B(p_input[14084]), .Z(n6574) );
  AND U13149 ( .A(n6575), .B(p_input[4083]), .Z(o[4083]) );
  AND U13150 ( .A(p_input[24083]), .B(p_input[14083]), .Z(n6575) );
  AND U13151 ( .A(n6576), .B(p_input[4082]), .Z(o[4082]) );
  AND U13152 ( .A(p_input[24082]), .B(p_input[14082]), .Z(n6576) );
  AND U13153 ( .A(n6577), .B(p_input[4081]), .Z(o[4081]) );
  AND U13154 ( .A(p_input[24081]), .B(p_input[14081]), .Z(n6577) );
  AND U13155 ( .A(n6578), .B(p_input[4080]), .Z(o[4080]) );
  AND U13156 ( .A(p_input[24080]), .B(p_input[14080]), .Z(n6578) );
  AND U13157 ( .A(n6579), .B(p_input[407]), .Z(o[407]) );
  AND U13158 ( .A(p_input[20407]), .B(p_input[10407]), .Z(n6579) );
  AND U13159 ( .A(n6580), .B(p_input[4079]), .Z(o[4079]) );
  AND U13160 ( .A(p_input[24079]), .B(p_input[14079]), .Z(n6580) );
  AND U13161 ( .A(n6581), .B(p_input[4078]), .Z(o[4078]) );
  AND U13162 ( .A(p_input[24078]), .B(p_input[14078]), .Z(n6581) );
  AND U13163 ( .A(n6582), .B(p_input[4077]), .Z(o[4077]) );
  AND U13164 ( .A(p_input[24077]), .B(p_input[14077]), .Z(n6582) );
  AND U13165 ( .A(n6583), .B(p_input[4076]), .Z(o[4076]) );
  AND U13166 ( .A(p_input[24076]), .B(p_input[14076]), .Z(n6583) );
  AND U13167 ( .A(n6584), .B(p_input[4075]), .Z(o[4075]) );
  AND U13168 ( .A(p_input[24075]), .B(p_input[14075]), .Z(n6584) );
  AND U13169 ( .A(n6585), .B(p_input[4074]), .Z(o[4074]) );
  AND U13170 ( .A(p_input[24074]), .B(p_input[14074]), .Z(n6585) );
  AND U13171 ( .A(n6586), .B(p_input[4073]), .Z(o[4073]) );
  AND U13172 ( .A(p_input[24073]), .B(p_input[14073]), .Z(n6586) );
  AND U13173 ( .A(n6587), .B(p_input[4072]), .Z(o[4072]) );
  AND U13174 ( .A(p_input[24072]), .B(p_input[14072]), .Z(n6587) );
  AND U13175 ( .A(n6588), .B(p_input[4071]), .Z(o[4071]) );
  AND U13176 ( .A(p_input[24071]), .B(p_input[14071]), .Z(n6588) );
  AND U13177 ( .A(n6589), .B(p_input[4070]), .Z(o[4070]) );
  AND U13178 ( .A(p_input[24070]), .B(p_input[14070]), .Z(n6589) );
  AND U13179 ( .A(n6590), .B(p_input[406]), .Z(o[406]) );
  AND U13180 ( .A(p_input[20406]), .B(p_input[10406]), .Z(n6590) );
  AND U13181 ( .A(n6591), .B(p_input[4069]), .Z(o[4069]) );
  AND U13182 ( .A(p_input[24069]), .B(p_input[14069]), .Z(n6591) );
  AND U13183 ( .A(n6592), .B(p_input[4068]), .Z(o[4068]) );
  AND U13184 ( .A(p_input[24068]), .B(p_input[14068]), .Z(n6592) );
  AND U13185 ( .A(n6593), .B(p_input[4067]), .Z(o[4067]) );
  AND U13186 ( .A(p_input[24067]), .B(p_input[14067]), .Z(n6593) );
  AND U13187 ( .A(n6594), .B(p_input[4066]), .Z(o[4066]) );
  AND U13188 ( .A(p_input[24066]), .B(p_input[14066]), .Z(n6594) );
  AND U13189 ( .A(n6595), .B(p_input[4065]), .Z(o[4065]) );
  AND U13190 ( .A(p_input[24065]), .B(p_input[14065]), .Z(n6595) );
  AND U13191 ( .A(n6596), .B(p_input[4064]), .Z(o[4064]) );
  AND U13192 ( .A(p_input[24064]), .B(p_input[14064]), .Z(n6596) );
  AND U13193 ( .A(n6597), .B(p_input[4063]), .Z(o[4063]) );
  AND U13194 ( .A(p_input[24063]), .B(p_input[14063]), .Z(n6597) );
  AND U13195 ( .A(n6598), .B(p_input[4062]), .Z(o[4062]) );
  AND U13196 ( .A(p_input[24062]), .B(p_input[14062]), .Z(n6598) );
  AND U13197 ( .A(n6599), .B(p_input[4061]), .Z(o[4061]) );
  AND U13198 ( .A(p_input[24061]), .B(p_input[14061]), .Z(n6599) );
  AND U13199 ( .A(n6600), .B(p_input[4060]), .Z(o[4060]) );
  AND U13200 ( .A(p_input[24060]), .B(p_input[14060]), .Z(n6600) );
  AND U13201 ( .A(n6601), .B(p_input[405]), .Z(o[405]) );
  AND U13202 ( .A(p_input[20405]), .B(p_input[10405]), .Z(n6601) );
  AND U13203 ( .A(n6602), .B(p_input[4059]), .Z(o[4059]) );
  AND U13204 ( .A(p_input[24059]), .B(p_input[14059]), .Z(n6602) );
  AND U13205 ( .A(n6603), .B(p_input[4058]), .Z(o[4058]) );
  AND U13206 ( .A(p_input[24058]), .B(p_input[14058]), .Z(n6603) );
  AND U13207 ( .A(n6604), .B(p_input[4057]), .Z(o[4057]) );
  AND U13208 ( .A(p_input[24057]), .B(p_input[14057]), .Z(n6604) );
  AND U13209 ( .A(n6605), .B(p_input[4056]), .Z(o[4056]) );
  AND U13210 ( .A(p_input[24056]), .B(p_input[14056]), .Z(n6605) );
  AND U13211 ( .A(n6606), .B(p_input[4055]), .Z(o[4055]) );
  AND U13212 ( .A(p_input[24055]), .B(p_input[14055]), .Z(n6606) );
  AND U13213 ( .A(n6607), .B(p_input[4054]), .Z(o[4054]) );
  AND U13214 ( .A(p_input[24054]), .B(p_input[14054]), .Z(n6607) );
  AND U13215 ( .A(n6608), .B(p_input[4053]), .Z(o[4053]) );
  AND U13216 ( .A(p_input[24053]), .B(p_input[14053]), .Z(n6608) );
  AND U13217 ( .A(n6609), .B(p_input[4052]), .Z(o[4052]) );
  AND U13218 ( .A(p_input[24052]), .B(p_input[14052]), .Z(n6609) );
  AND U13219 ( .A(n6610), .B(p_input[4051]), .Z(o[4051]) );
  AND U13220 ( .A(p_input[24051]), .B(p_input[14051]), .Z(n6610) );
  AND U13221 ( .A(n6611), .B(p_input[4050]), .Z(o[4050]) );
  AND U13222 ( .A(p_input[24050]), .B(p_input[14050]), .Z(n6611) );
  AND U13223 ( .A(n6612), .B(p_input[404]), .Z(o[404]) );
  AND U13224 ( .A(p_input[20404]), .B(p_input[10404]), .Z(n6612) );
  AND U13225 ( .A(n6613), .B(p_input[4049]), .Z(o[4049]) );
  AND U13226 ( .A(p_input[24049]), .B(p_input[14049]), .Z(n6613) );
  AND U13227 ( .A(n6614), .B(p_input[4048]), .Z(o[4048]) );
  AND U13228 ( .A(p_input[24048]), .B(p_input[14048]), .Z(n6614) );
  AND U13229 ( .A(n6615), .B(p_input[4047]), .Z(o[4047]) );
  AND U13230 ( .A(p_input[24047]), .B(p_input[14047]), .Z(n6615) );
  AND U13231 ( .A(n6616), .B(p_input[4046]), .Z(o[4046]) );
  AND U13232 ( .A(p_input[24046]), .B(p_input[14046]), .Z(n6616) );
  AND U13233 ( .A(n6617), .B(p_input[4045]), .Z(o[4045]) );
  AND U13234 ( .A(p_input[24045]), .B(p_input[14045]), .Z(n6617) );
  AND U13235 ( .A(n6618), .B(p_input[4044]), .Z(o[4044]) );
  AND U13236 ( .A(p_input[24044]), .B(p_input[14044]), .Z(n6618) );
  AND U13237 ( .A(n6619), .B(p_input[4043]), .Z(o[4043]) );
  AND U13238 ( .A(p_input[24043]), .B(p_input[14043]), .Z(n6619) );
  AND U13239 ( .A(n6620), .B(p_input[4042]), .Z(o[4042]) );
  AND U13240 ( .A(p_input[24042]), .B(p_input[14042]), .Z(n6620) );
  AND U13241 ( .A(n6621), .B(p_input[4041]), .Z(o[4041]) );
  AND U13242 ( .A(p_input[24041]), .B(p_input[14041]), .Z(n6621) );
  AND U13243 ( .A(n6622), .B(p_input[4040]), .Z(o[4040]) );
  AND U13244 ( .A(p_input[24040]), .B(p_input[14040]), .Z(n6622) );
  AND U13245 ( .A(n6623), .B(p_input[403]), .Z(o[403]) );
  AND U13246 ( .A(p_input[20403]), .B(p_input[10403]), .Z(n6623) );
  AND U13247 ( .A(n6624), .B(p_input[4039]), .Z(o[4039]) );
  AND U13248 ( .A(p_input[24039]), .B(p_input[14039]), .Z(n6624) );
  AND U13249 ( .A(n6625), .B(p_input[4038]), .Z(o[4038]) );
  AND U13250 ( .A(p_input[24038]), .B(p_input[14038]), .Z(n6625) );
  AND U13251 ( .A(n6626), .B(p_input[4037]), .Z(o[4037]) );
  AND U13252 ( .A(p_input[24037]), .B(p_input[14037]), .Z(n6626) );
  AND U13253 ( .A(n6627), .B(p_input[4036]), .Z(o[4036]) );
  AND U13254 ( .A(p_input[24036]), .B(p_input[14036]), .Z(n6627) );
  AND U13255 ( .A(n6628), .B(p_input[4035]), .Z(o[4035]) );
  AND U13256 ( .A(p_input[24035]), .B(p_input[14035]), .Z(n6628) );
  AND U13257 ( .A(n6629), .B(p_input[4034]), .Z(o[4034]) );
  AND U13258 ( .A(p_input[24034]), .B(p_input[14034]), .Z(n6629) );
  AND U13259 ( .A(n6630), .B(p_input[4033]), .Z(o[4033]) );
  AND U13260 ( .A(p_input[24033]), .B(p_input[14033]), .Z(n6630) );
  AND U13261 ( .A(n6631), .B(p_input[4032]), .Z(o[4032]) );
  AND U13262 ( .A(p_input[24032]), .B(p_input[14032]), .Z(n6631) );
  AND U13263 ( .A(n6632), .B(p_input[4031]), .Z(o[4031]) );
  AND U13264 ( .A(p_input[24031]), .B(p_input[14031]), .Z(n6632) );
  AND U13265 ( .A(n6633), .B(p_input[4030]), .Z(o[4030]) );
  AND U13266 ( .A(p_input[24030]), .B(p_input[14030]), .Z(n6633) );
  AND U13267 ( .A(n6634), .B(p_input[402]), .Z(o[402]) );
  AND U13268 ( .A(p_input[20402]), .B(p_input[10402]), .Z(n6634) );
  AND U13269 ( .A(n6635), .B(p_input[4029]), .Z(o[4029]) );
  AND U13270 ( .A(p_input[24029]), .B(p_input[14029]), .Z(n6635) );
  AND U13271 ( .A(n6636), .B(p_input[4028]), .Z(o[4028]) );
  AND U13272 ( .A(p_input[24028]), .B(p_input[14028]), .Z(n6636) );
  AND U13273 ( .A(n6637), .B(p_input[4027]), .Z(o[4027]) );
  AND U13274 ( .A(p_input[24027]), .B(p_input[14027]), .Z(n6637) );
  AND U13275 ( .A(n6638), .B(p_input[4026]), .Z(o[4026]) );
  AND U13276 ( .A(p_input[24026]), .B(p_input[14026]), .Z(n6638) );
  AND U13277 ( .A(n6639), .B(p_input[4025]), .Z(o[4025]) );
  AND U13278 ( .A(p_input[24025]), .B(p_input[14025]), .Z(n6639) );
  AND U13279 ( .A(n6640), .B(p_input[4024]), .Z(o[4024]) );
  AND U13280 ( .A(p_input[24024]), .B(p_input[14024]), .Z(n6640) );
  AND U13281 ( .A(n6641), .B(p_input[4023]), .Z(o[4023]) );
  AND U13282 ( .A(p_input[24023]), .B(p_input[14023]), .Z(n6641) );
  AND U13283 ( .A(n6642), .B(p_input[4022]), .Z(o[4022]) );
  AND U13284 ( .A(p_input[24022]), .B(p_input[14022]), .Z(n6642) );
  AND U13285 ( .A(n6643), .B(p_input[4021]), .Z(o[4021]) );
  AND U13286 ( .A(p_input[24021]), .B(p_input[14021]), .Z(n6643) );
  AND U13287 ( .A(n6644), .B(p_input[4020]), .Z(o[4020]) );
  AND U13288 ( .A(p_input[24020]), .B(p_input[14020]), .Z(n6644) );
  AND U13289 ( .A(n6645), .B(p_input[401]), .Z(o[401]) );
  AND U13290 ( .A(p_input[20401]), .B(p_input[10401]), .Z(n6645) );
  AND U13291 ( .A(n6646), .B(p_input[4019]), .Z(o[4019]) );
  AND U13292 ( .A(p_input[24019]), .B(p_input[14019]), .Z(n6646) );
  AND U13293 ( .A(n6647), .B(p_input[4018]), .Z(o[4018]) );
  AND U13294 ( .A(p_input[24018]), .B(p_input[14018]), .Z(n6647) );
  AND U13295 ( .A(n6648), .B(p_input[4017]), .Z(o[4017]) );
  AND U13296 ( .A(p_input[24017]), .B(p_input[14017]), .Z(n6648) );
  AND U13297 ( .A(n6649), .B(p_input[4016]), .Z(o[4016]) );
  AND U13298 ( .A(p_input[24016]), .B(p_input[14016]), .Z(n6649) );
  AND U13299 ( .A(n6650), .B(p_input[4015]), .Z(o[4015]) );
  AND U13300 ( .A(p_input[24015]), .B(p_input[14015]), .Z(n6650) );
  AND U13301 ( .A(n6651), .B(p_input[4014]), .Z(o[4014]) );
  AND U13302 ( .A(p_input[24014]), .B(p_input[14014]), .Z(n6651) );
  AND U13303 ( .A(n6652), .B(p_input[4013]), .Z(o[4013]) );
  AND U13304 ( .A(p_input[24013]), .B(p_input[14013]), .Z(n6652) );
  AND U13305 ( .A(n6653), .B(p_input[4012]), .Z(o[4012]) );
  AND U13306 ( .A(p_input[24012]), .B(p_input[14012]), .Z(n6653) );
  AND U13307 ( .A(n6654), .B(p_input[4011]), .Z(o[4011]) );
  AND U13308 ( .A(p_input[24011]), .B(p_input[14011]), .Z(n6654) );
  AND U13309 ( .A(n6655), .B(p_input[4010]), .Z(o[4010]) );
  AND U13310 ( .A(p_input[24010]), .B(p_input[14010]), .Z(n6655) );
  AND U13311 ( .A(n6656), .B(p_input[400]), .Z(o[400]) );
  AND U13312 ( .A(p_input[20400]), .B(p_input[10400]), .Z(n6656) );
  AND U13313 ( .A(n6657), .B(p_input[4009]), .Z(o[4009]) );
  AND U13314 ( .A(p_input[24009]), .B(p_input[14009]), .Z(n6657) );
  AND U13315 ( .A(n6658), .B(p_input[4008]), .Z(o[4008]) );
  AND U13316 ( .A(p_input[24008]), .B(p_input[14008]), .Z(n6658) );
  AND U13317 ( .A(n6659), .B(p_input[4007]), .Z(o[4007]) );
  AND U13318 ( .A(p_input[24007]), .B(p_input[14007]), .Z(n6659) );
  AND U13319 ( .A(n6660), .B(p_input[4006]), .Z(o[4006]) );
  AND U13320 ( .A(p_input[24006]), .B(p_input[14006]), .Z(n6660) );
  AND U13321 ( .A(n6661), .B(p_input[4005]), .Z(o[4005]) );
  AND U13322 ( .A(p_input[24005]), .B(p_input[14005]), .Z(n6661) );
  AND U13323 ( .A(n6662), .B(p_input[4004]), .Z(o[4004]) );
  AND U13324 ( .A(p_input[24004]), .B(p_input[14004]), .Z(n6662) );
  AND U13325 ( .A(n6663), .B(p_input[4003]), .Z(o[4003]) );
  AND U13326 ( .A(p_input[24003]), .B(p_input[14003]), .Z(n6663) );
  AND U13327 ( .A(n6664), .B(p_input[4002]), .Z(o[4002]) );
  AND U13328 ( .A(p_input[24002]), .B(p_input[14002]), .Z(n6664) );
  AND U13329 ( .A(n6665), .B(p_input[4001]), .Z(o[4001]) );
  AND U13330 ( .A(p_input[24001]), .B(p_input[14001]), .Z(n6665) );
  AND U13331 ( .A(n6666), .B(p_input[4000]), .Z(o[4000]) );
  AND U13332 ( .A(p_input[24000]), .B(p_input[14000]), .Z(n6666) );
  AND U13333 ( .A(n6667), .B(p_input[3]), .Z(o[3]) );
  AND U13334 ( .A(p_input[20003]), .B(p_input[10003]), .Z(n6667) );
  AND U13335 ( .A(n6668), .B(p_input[39]), .Z(o[39]) );
  AND U13336 ( .A(p_input[20039]), .B(p_input[10039]), .Z(n6668) );
  AND U13337 ( .A(n6669), .B(p_input[399]), .Z(o[399]) );
  AND U13338 ( .A(p_input[20399]), .B(p_input[10399]), .Z(n6669) );
  AND U13339 ( .A(n6670), .B(p_input[3999]), .Z(o[3999]) );
  AND U13340 ( .A(p_input[23999]), .B(p_input[13999]), .Z(n6670) );
  AND U13341 ( .A(n6671), .B(p_input[3998]), .Z(o[3998]) );
  AND U13342 ( .A(p_input[23998]), .B(p_input[13998]), .Z(n6671) );
  AND U13343 ( .A(n6672), .B(p_input[3997]), .Z(o[3997]) );
  AND U13344 ( .A(p_input[23997]), .B(p_input[13997]), .Z(n6672) );
  AND U13345 ( .A(n6673), .B(p_input[3996]), .Z(o[3996]) );
  AND U13346 ( .A(p_input[23996]), .B(p_input[13996]), .Z(n6673) );
  AND U13347 ( .A(n6674), .B(p_input[3995]), .Z(o[3995]) );
  AND U13348 ( .A(p_input[23995]), .B(p_input[13995]), .Z(n6674) );
  AND U13349 ( .A(n6675), .B(p_input[3994]), .Z(o[3994]) );
  AND U13350 ( .A(p_input[23994]), .B(p_input[13994]), .Z(n6675) );
  AND U13351 ( .A(n6676), .B(p_input[3993]), .Z(o[3993]) );
  AND U13352 ( .A(p_input[23993]), .B(p_input[13993]), .Z(n6676) );
  AND U13353 ( .A(n6677), .B(p_input[3992]), .Z(o[3992]) );
  AND U13354 ( .A(p_input[23992]), .B(p_input[13992]), .Z(n6677) );
  AND U13355 ( .A(n6678), .B(p_input[3991]), .Z(o[3991]) );
  AND U13356 ( .A(p_input[23991]), .B(p_input[13991]), .Z(n6678) );
  AND U13357 ( .A(n6679), .B(p_input[3990]), .Z(o[3990]) );
  AND U13358 ( .A(p_input[23990]), .B(p_input[13990]), .Z(n6679) );
  AND U13359 ( .A(n6680), .B(p_input[398]), .Z(o[398]) );
  AND U13360 ( .A(p_input[20398]), .B(p_input[10398]), .Z(n6680) );
  AND U13361 ( .A(n6681), .B(p_input[3989]), .Z(o[3989]) );
  AND U13362 ( .A(p_input[23989]), .B(p_input[13989]), .Z(n6681) );
  AND U13363 ( .A(n6682), .B(p_input[3988]), .Z(o[3988]) );
  AND U13364 ( .A(p_input[23988]), .B(p_input[13988]), .Z(n6682) );
  AND U13365 ( .A(n6683), .B(p_input[3987]), .Z(o[3987]) );
  AND U13366 ( .A(p_input[23987]), .B(p_input[13987]), .Z(n6683) );
  AND U13367 ( .A(n6684), .B(p_input[3986]), .Z(o[3986]) );
  AND U13368 ( .A(p_input[23986]), .B(p_input[13986]), .Z(n6684) );
  AND U13369 ( .A(n6685), .B(p_input[3985]), .Z(o[3985]) );
  AND U13370 ( .A(p_input[23985]), .B(p_input[13985]), .Z(n6685) );
  AND U13371 ( .A(n6686), .B(p_input[3984]), .Z(o[3984]) );
  AND U13372 ( .A(p_input[23984]), .B(p_input[13984]), .Z(n6686) );
  AND U13373 ( .A(n6687), .B(p_input[3983]), .Z(o[3983]) );
  AND U13374 ( .A(p_input[23983]), .B(p_input[13983]), .Z(n6687) );
  AND U13375 ( .A(n6688), .B(p_input[3982]), .Z(o[3982]) );
  AND U13376 ( .A(p_input[23982]), .B(p_input[13982]), .Z(n6688) );
  AND U13377 ( .A(n6689), .B(p_input[3981]), .Z(o[3981]) );
  AND U13378 ( .A(p_input[23981]), .B(p_input[13981]), .Z(n6689) );
  AND U13379 ( .A(n6690), .B(p_input[3980]), .Z(o[3980]) );
  AND U13380 ( .A(p_input[23980]), .B(p_input[13980]), .Z(n6690) );
  AND U13381 ( .A(n6691), .B(p_input[397]), .Z(o[397]) );
  AND U13382 ( .A(p_input[20397]), .B(p_input[10397]), .Z(n6691) );
  AND U13383 ( .A(n6692), .B(p_input[3979]), .Z(o[3979]) );
  AND U13384 ( .A(p_input[23979]), .B(p_input[13979]), .Z(n6692) );
  AND U13385 ( .A(n6693), .B(p_input[3978]), .Z(o[3978]) );
  AND U13386 ( .A(p_input[23978]), .B(p_input[13978]), .Z(n6693) );
  AND U13387 ( .A(n6694), .B(p_input[3977]), .Z(o[3977]) );
  AND U13388 ( .A(p_input[23977]), .B(p_input[13977]), .Z(n6694) );
  AND U13389 ( .A(n6695), .B(p_input[3976]), .Z(o[3976]) );
  AND U13390 ( .A(p_input[23976]), .B(p_input[13976]), .Z(n6695) );
  AND U13391 ( .A(n6696), .B(p_input[3975]), .Z(o[3975]) );
  AND U13392 ( .A(p_input[23975]), .B(p_input[13975]), .Z(n6696) );
  AND U13393 ( .A(n6697), .B(p_input[3974]), .Z(o[3974]) );
  AND U13394 ( .A(p_input[23974]), .B(p_input[13974]), .Z(n6697) );
  AND U13395 ( .A(n6698), .B(p_input[3973]), .Z(o[3973]) );
  AND U13396 ( .A(p_input[23973]), .B(p_input[13973]), .Z(n6698) );
  AND U13397 ( .A(n6699), .B(p_input[3972]), .Z(o[3972]) );
  AND U13398 ( .A(p_input[23972]), .B(p_input[13972]), .Z(n6699) );
  AND U13399 ( .A(n6700), .B(p_input[3971]), .Z(o[3971]) );
  AND U13400 ( .A(p_input[23971]), .B(p_input[13971]), .Z(n6700) );
  AND U13401 ( .A(n6701), .B(p_input[3970]), .Z(o[3970]) );
  AND U13402 ( .A(p_input[23970]), .B(p_input[13970]), .Z(n6701) );
  AND U13403 ( .A(n6702), .B(p_input[396]), .Z(o[396]) );
  AND U13404 ( .A(p_input[20396]), .B(p_input[10396]), .Z(n6702) );
  AND U13405 ( .A(n6703), .B(p_input[3969]), .Z(o[3969]) );
  AND U13406 ( .A(p_input[23969]), .B(p_input[13969]), .Z(n6703) );
  AND U13407 ( .A(n6704), .B(p_input[3968]), .Z(o[3968]) );
  AND U13408 ( .A(p_input[23968]), .B(p_input[13968]), .Z(n6704) );
  AND U13409 ( .A(n6705), .B(p_input[3967]), .Z(o[3967]) );
  AND U13410 ( .A(p_input[23967]), .B(p_input[13967]), .Z(n6705) );
  AND U13411 ( .A(n6706), .B(p_input[3966]), .Z(o[3966]) );
  AND U13412 ( .A(p_input[23966]), .B(p_input[13966]), .Z(n6706) );
  AND U13413 ( .A(n6707), .B(p_input[3965]), .Z(o[3965]) );
  AND U13414 ( .A(p_input[23965]), .B(p_input[13965]), .Z(n6707) );
  AND U13415 ( .A(n6708), .B(p_input[3964]), .Z(o[3964]) );
  AND U13416 ( .A(p_input[23964]), .B(p_input[13964]), .Z(n6708) );
  AND U13417 ( .A(n6709), .B(p_input[3963]), .Z(o[3963]) );
  AND U13418 ( .A(p_input[23963]), .B(p_input[13963]), .Z(n6709) );
  AND U13419 ( .A(n6710), .B(p_input[3962]), .Z(o[3962]) );
  AND U13420 ( .A(p_input[23962]), .B(p_input[13962]), .Z(n6710) );
  AND U13421 ( .A(n6711), .B(p_input[3961]), .Z(o[3961]) );
  AND U13422 ( .A(p_input[23961]), .B(p_input[13961]), .Z(n6711) );
  AND U13423 ( .A(n6712), .B(p_input[3960]), .Z(o[3960]) );
  AND U13424 ( .A(p_input[23960]), .B(p_input[13960]), .Z(n6712) );
  AND U13425 ( .A(n6713), .B(p_input[395]), .Z(o[395]) );
  AND U13426 ( .A(p_input[20395]), .B(p_input[10395]), .Z(n6713) );
  AND U13427 ( .A(n6714), .B(p_input[3959]), .Z(o[3959]) );
  AND U13428 ( .A(p_input[23959]), .B(p_input[13959]), .Z(n6714) );
  AND U13429 ( .A(n6715), .B(p_input[3958]), .Z(o[3958]) );
  AND U13430 ( .A(p_input[23958]), .B(p_input[13958]), .Z(n6715) );
  AND U13431 ( .A(n6716), .B(p_input[3957]), .Z(o[3957]) );
  AND U13432 ( .A(p_input[23957]), .B(p_input[13957]), .Z(n6716) );
  AND U13433 ( .A(n6717), .B(p_input[3956]), .Z(o[3956]) );
  AND U13434 ( .A(p_input[23956]), .B(p_input[13956]), .Z(n6717) );
  AND U13435 ( .A(n6718), .B(p_input[3955]), .Z(o[3955]) );
  AND U13436 ( .A(p_input[23955]), .B(p_input[13955]), .Z(n6718) );
  AND U13437 ( .A(n6719), .B(p_input[3954]), .Z(o[3954]) );
  AND U13438 ( .A(p_input[23954]), .B(p_input[13954]), .Z(n6719) );
  AND U13439 ( .A(n6720), .B(p_input[3953]), .Z(o[3953]) );
  AND U13440 ( .A(p_input[23953]), .B(p_input[13953]), .Z(n6720) );
  AND U13441 ( .A(n6721), .B(p_input[3952]), .Z(o[3952]) );
  AND U13442 ( .A(p_input[23952]), .B(p_input[13952]), .Z(n6721) );
  AND U13443 ( .A(n6722), .B(p_input[3951]), .Z(o[3951]) );
  AND U13444 ( .A(p_input[23951]), .B(p_input[13951]), .Z(n6722) );
  AND U13445 ( .A(n6723), .B(p_input[3950]), .Z(o[3950]) );
  AND U13446 ( .A(p_input[23950]), .B(p_input[13950]), .Z(n6723) );
  AND U13447 ( .A(n6724), .B(p_input[394]), .Z(o[394]) );
  AND U13448 ( .A(p_input[20394]), .B(p_input[10394]), .Z(n6724) );
  AND U13449 ( .A(n6725), .B(p_input[3949]), .Z(o[3949]) );
  AND U13450 ( .A(p_input[23949]), .B(p_input[13949]), .Z(n6725) );
  AND U13451 ( .A(n6726), .B(p_input[3948]), .Z(o[3948]) );
  AND U13452 ( .A(p_input[23948]), .B(p_input[13948]), .Z(n6726) );
  AND U13453 ( .A(n6727), .B(p_input[3947]), .Z(o[3947]) );
  AND U13454 ( .A(p_input[23947]), .B(p_input[13947]), .Z(n6727) );
  AND U13455 ( .A(n6728), .B(p_input[3946]), .Z(o[3946]) );
  AND U13456 ( .A(p_input[23946]), .B(p_input[13946]), .Z(n6728) );
  AND U13457 ( .A(n6729), .B(p_input[3945]), .Z(o[3945]) );
  AND U13458 ( .A(p_input[23945]), .B(p_input[13945]), .Z(n6729) );
  AND U13459 ( .A(n6730), .B(p_input[3944]), .Z(o[3944]) );
  AND U13460 ( .A(p_input[23944]), .B(p_input[13944]), .Z(n6730) );
  AND U13461 ( .A(n6731), .B(p_input[3943]), .Z(o[3943]) );
  AND U13462 ( .A(p_input[23943]), .B(p_input[13943]), .Z(n6731) );
  AND U13463 ( .A(n6732), .B(p_input[3942]), .Z(o[3942]) );
  AND U13464 ( .A(p_input[23942]), .B(p_input[13942]), .Z(n6732) );
  AND U13465 ( .A(n6733), .B(p_input[3941]), .Z(o[3941]) );
  AND U13466 ( .A(p_input[23941]), .B(p_input[13941]), .Z(n6733) );
  AND U13467 ( .A(n6734), .B(p_input[3940]), .Z(o[3940]) );
  AND U13468 ( .A(p_input[23940]), .B(p_input[13940]), .Z(n6734) );
  AND U13469 ( .A(n6735), .B(p_input[393]), .Z(o[393]) );
  AND U13470 ( .A(p_input[20393]), .B(p_input[10393]), .Z(n6735) );
  AND U13471 ( .A(n6736), .B(p_input[3939]), .Z(o[3939]) );
  AND U13472 ( .A(p_input[23939]), .B(p_input[13939]), .Z(n6736) );
  AND U13473 ( .A(n6737), .B(p_input[3938]), .Z(o[3938]) );
  AND U13474 ( .A(p_input[23938]), .B(p_input[13938]), .Z(n6737) );
  AND U13475 ( .A(n6738), .B(p_input[3937]), .Z(o[3937]) );
  AND U13476 ( .A(p_input[23937]), .B(p_input[13937]), .Z(n6738) );
  AND U13477 ( .A(n6739), .B(p_input[3936]), .Z(o[3936]) );
  AND U13478 ( .A(p_input[23936]), .B(p_input[13936]), .Z(n6739) );
  AND U13479 ( .A(n6740), .B(p_input[3935]), .Z(o[3935]) );
  AND U13480 ( .A(p_input[23935]), .B(p_input[13935]), .Z(n6740) );
  AND U13481 ( .A(n6741), .B(p_input[3934]), .Z(o[3934]) );
  AND U13482 ( .A(p_input[23934]), .B(p_input[13934]), .Z(n6741) );
  AND U13483 ( .A(n6742), .B(p_input[3933]), .Z(o[3933]) );
  AND U13484 ( .A(p_input[23933]), .B(p_input[13933]), .Z(n6742) );
  AND U13485 ( .A(n6743), .B(p_input[3932]), .Z(o[3932]) );
  AND U13486 ( .A(p_input[23932]), .B(p_input[13932]), .Z(n6743) );
  AND U13487 ( .A(n6744), .B(p_input[3931]), .Z(o[3931]) );
  AND U13488 ( .A(p_input[23931]), .B(p_input[13931]), .Z(n6744) );
  AND U13489 ( .A(n6745), .B(p_input[3930]), .Z(o[3930]) );
  AND U13490 ( .A(p_input[23930]), .B(p_input[13930]), .Z(n6745) );
  AND U13491 ( .A(n6746), .B(p_input[392]), .Z(o[392]) );
  AND U13492 ( .A(p_input[20392]), .B(p_input[10392]), .Z(n6746) );
  AND U13493 ( .A(n6747), .B(p_input[3929]), .Z(o[3929]) );
  AND U13494 ( .A(p_input[23929]), .B(p_input[13929]), .Z(n6747) );
  AND U13495 ( .A(n6748), .B(p_input[3928]), .Z(o[3928]) );
  AND U13496 ( .A(p_input[23928]), .B(p_input[13928]), .Z(n6748) );
  AND U13497 ( .A(n6749), .B(p_input[3927]), .Z(o[3927]) );
  AND U13498 ( .A(p_input[23927]), .B(p_input[13927]), .Z(n6749) );
  AND U13499 ( .A(n6750), .B(p_input[3926]), .Z(o[3926]) );
  AND U13500 ( .A(p_input[23926]), .B(p_input[13926]), .Z(n6750) );
  AND U13501 ( .A(n6751), .B(p_input[3925]), .Z(o[3925]) );
  AND U13502 ( .A(p_input[23925]), .B(p_input[13925]), .Z(n6751) );
  AND U13503 ( .A(n6752), .B(p_input[3924]), .Z(o[3924]) );
  AND U13504 ( .A(p_input[23924]), .B(p_input[13924]), .Z(n6752) );
  AND U13505 ( .A(n6753), .B(p_input[3923]), .Z(o[3923]) );
  AND U13506 ( .A(p_input[23923]), .B(p_input[13923]), .Z(n6753) );
  AND U13507 ( .A(n6754), .B(p_input[3922]), .Z(o[3922]) );
  AND U13508 ( .A(p_input[23922]), .B(p_input[13922]), .Z(n6754) );
  AND U13509 ( .A(n6755), .B(p_input[3921]), .Z(o[3921]) );
  AND U13510 ( .A(p_input[23921]), .B(p_input[13921]), .Z(n6755) );
  AND U13511 ( .A(n6756), .B(p_input[3920]), .Z(o[3920]) );
  AND U13512 ( .A(p_input[23920]), .B(p_input[13920]), .Z(n6756) );
  AND U13513 ( .A(n6757), .B(p_input[391]), .Z(o[391]) );
  AND U13514 ( .A(p_input[20391]), .B(p_input[10391]), .Z(n6757) );
  AND U13515 ( .A(n6758), .B(p_input[3919]), .Z(o[3919]) );
  AND U13516 ( .A(p_input[23919]), .B(p_input[13919]), .Z(n6758) );
  AND U13517 ( .A(n6759), .B(p_input[3918]), .Z(o[3918]) );
  AND U13518 ( .A(p_input[23918]), .B(p_input[13918]), .Z(n6759) );
  AND U13519 ( .A(n6760), .B(p_input[3917]), .Z(o[3917]) );
  AND U13520 ( .A(p_input[23917]), .B(p_input[13917]), .Z(n6760) );
  AND U13521 ( .A(n6761), .B(p_input[3916]), .Z(o[3916]) );
  AND U13522 ( .A(p_input[23916]), .B(p_input[13916]), .Z(n6761) );
  AND U13523 ( .A(n6762), .B(p_input[3915]), .Z(o[3915]) );
  AND U13524 ( .A(p_input[23915]), .B(p_input[13915]), .Z(n6762) );
  AND U13525 ( .A(n6763), .B(p_input[3914]), .Z(o[3914]) );
  AND U13526 ( .A(p_input[23914]), .B(p_input[13914]), .Z(n6763) );
  AND U13527 ( .A(n6764), .B(p_input[3913]), .Z(o[3913]) );
  AND U13528 ( .A(p_input[23913]), .B(p_input[13913]), .Z(n6764) );
  AND U13529 ( .A(n6765), .B(p_input[3912]), .Z(o[3912]) );
  AND U13530 ( .A(p_input[23912]), .B(p_input[13912]), .Z(n6765) );
  AND U13531 ( .A(n6766), .B(p_input[3911]), .Z(o[3911]) );
  AND U13532 ( .A(p_input[23911]), .B(p_input[13911]), .Z(n6766) );
  AND U13533 ( .A(n6767), .B(p_input[3910]), .Z(o[3910]) );
  AND U13534 ( .A(p_input[23910]), .B(p_input[13910]), .Z(n6767) );
  AND U13535 ( .A(n6768), .B(p_input[390]), .Z(o[390]) );
  AND U13536 ( .A(p_input[20390]), .B(p_input[10390]), .Z(n6768) );
  AND U13537 ( .A(n6769), .B(p_input[3909]), .Z(o[3909]) );
  AND U13538 ( .A(p_input[23909]), .B(p_input[13909]), .Z(n6769) );
  AND U13539 ( .A(n6770), .B(p_input[3908]), .Z(o[3908]) );
  AND U13540 ( .A(p_input[23908]), .B(p_input[13908]), .Z(n6770) );
  AND U13541 ( .A(n6771), .B(p_input[3907]), .Z(o[3907]) );
  AND U13542 ( .A(p_input[23907]), .B(p_input[13907]), .Z(n6771) );
  AND U13543 ( .A(n6772), .B(p_input[3906]), .Z(o[3906]) );
  AND U13544 ( .A(p_input[23906]), .B(p_input[13906]), .Z(n6772) );
  AND U13545 ( .A(n6773), .B(p_input[3905]), .Z(o[3905]) );
  AND U13546 ( .A(p_input[23905]), .B(p_input[13905]), .Z(n6773) );
  AND U13547 ( .A(n6774), .B(p_input[3904]), .Z(o[3904]) );
  AND U13548 ( .A(p_input[23904]), .B(p_input[13904]), .Z(n6774) );
  AND U13549 ( .A(n6775), .B(p_input[3903]), .Z(o[3903]) );
  AND U13550 ( .A(p_input[23903]), .B(p_input[13903]), .Z(n6775) );
  AND U13551 ( .A(n6776), .B(p_input[3902]), .Z(o[3902]) );
  AND U13552 ( .A(p_input[23902]), .B(p_input[13902]), .Z(n6776) );
  AND U13553 ( .A(n6777), .B(p_input[3901]), .Z(o[3901]) );
  AND U13554 ( .A(p_input[23901]), .B(p_input[13901]), .Z(n6777) );
  AND U13555 ( .A(n6778), .B(p_input[3900]), .Z(o[3900]) );
  AND U13556 ( .A(p_input[23900]), .B(p_input[13900]), .Z(n6778) );
  AND U13557 ( .A(n6779), .B(p_input[38]), .Z(o[38]) );
  AND U13558 ( .A(p_input[20038]), .B(p_input[10038]), .Z(n6779) );
  AND U13559 ( .A(n6780), .B(p_input[389]), .Z(o[389]) );
  AND U13560 ( .A(p_input[20389]), .B(p_input[10389]), .Z(n6780) );
  AND U13561 ( .A(n6781), .B(p_input[3899]), .Z(o[3899]) );
  AND U13562 ( .A(p_input[23899]), .B(p_input[13899]), .Z(n6781) );
  AND U13563 ( .A(n6782), .B(p_input[3898]), .Z(o[3898]) );
  AND U13564 ( .A(p_input[23898]), .B(p_input[13898]), .Z(n6782) );
  AND U13565 ( .A(n6783), .B(p_input[3897]), .Z(o[3897]) );
  AND U13566 ( .A(p_input[23897]), .B(p_input[13897]), .Z(n6783) );
  AND U13567 ( .A(n6784), .B(p_input[3896]), .Z(o[3896]) );
  AND U13568 ( .A(p_input[23896]), .B(p_input[13896]), .Z(n6784) );
  AND U13569 ( .A(n6785), .B(p_input[3895]), .Z(o[3895]) );
  AND U13570 ( .A(p_input[23895]), .B(p_input[13895]), .Z(n6785) );
  AND U13571 ( .A(n6786), .B(p_input[3894]), .Z(o[3894]) );
  AND U13572 ( .A(p_input[23894]), .B(p_input[13894]), .Z(n6786) );
  AND U13573 ( .A(n6787), .B(p_input[3893]), .Z(o[3893]) );
  AND U13574 ( .A(p_input[23893]), .B(p_input[13893]), .Z(n6787) );
  AND U13575 ( .A(n6788), .B(p_input[3892]), .Z(o[3892]) );
  AND U13576 ( .A(p_input[23892]), .B(p_input[13892]), .Z(n6788) );
  AND U13577 ( .A(n6789), .B(p_input[3891]), .Z(o[3891]) );
  AND U13578 ( .A(p_input[23891]), .B(p_input[13891]), .Z(n6789) );
  AND U13579 ( .A(n6790), .B(p_input[3890]), .Z(o[3890]) );
  AND U13580 ( .A(p_input[23890]), .B(p_input[13890]), .Z(n6790) );
  AND U13581 ( .A(n6791), .B(p_input[388]), .Z(o[388]) );
  AND U13582 ( .A(p_input[20388]), .B(p_input[10388]), .Z(n6791) );
  AND U13583 ( .A(n6792), .B(p_input[3889]), .Z(o[3889]) );
  AND U13584 ( .A(p_input[23889]), .B(p_input[13889]), .Z(n6792) );
  AND U13585 ( .A(n6793), .B(p_input[3888]), .Z(o[3888]) );
  AND U13586 ( .A(p_input[23888]), .B(p_input[13888]), .Z(n6793) );
  AND U13587 ( .A(n6794), .B(p_input[3887]), .Z(o[3887]) );
  AND U13588 ( .A(p_input[23887]), .B(p_input[13887]), .Z(n6794) );
  AND U13589 ( .A(n6795), .B(p_input[3886]), .Z(o[3886]) );
  AND U13590 ( .A(p_input[23886]), .B(p_input[13886]), .Z(n6795) );
  AND U13591 ( .A(n6796), .B(p_input[3885]), .Z(o[3885]) );
  AND U13592 ( .A(p_input[23885]), .B(p_input[13885]), .Z(n6796) );
  AND U13593 ( .A(n6797), .B(p_input[3884]), .Z(o[3884]) );
  AND U13594 ( .A(p_input[23884]), .B(p_input[13884]), .Z(n6797) );
  AND U13595 ( .A(n6798), .B(p_input[3883]), .Z(o[3883]) );
  AND U13596 ( .A(p_input[23883]), .B(p_input[13883]), .Z(n6798) );
  AND U13597 ( .A(n6799), .B(p_input[3882]), .Z(o[3882]) );
  AND U13598 ( .A(p_input[23882]), .B(p_input[13882]), .Z(n6799) );
  AND U13599 ( .A(n6800), .B(p_input[3881]), .Z(o[3881]) );
  AND U13600 ( .A(p_input[23881]), .B(p_input[13881]), .Z(n6800) );
  AND U13601 ( .A(n6801), .B(p_input[3880]), .Z(o[3880]) );
  AND U13602 ( .A(p_input[23880]), .B(p_input[13880]), .Z(n6801) );
  AND U13603 ( .A(n6802), .B(p_input[387]), .Z(o[387]) );
  AND U13604 ( .A(p_input[20387]), .B(p_input[10387]), .Z(n6802) );
  AND U13605 ( .A(n6803), .B(p_input[3879]), .Z(o[3879]) );
  AND U13606 ( .A(p_input[23879]), .B(p_input[13879]), .Z(n6803) );
  AND U13607 ( .A(n6804), .B(p_input[3878]), .Z(o[3878]) );
  AND U13608 ( .A(p_input[23878]), .B(p_input[13878]), .Z(n6804) );
  AND U13609 ( .A(n6805), .B(p_input[3877]), .Z(o[3877]) );
  AND U13610 ( .A(p_input[23877]), .B(p_input[13877]), .Z(n6805) );
  AND U13611 ( .A(n6806), .B(p_input[3876]), .Z(o[3876]) );
  AND U13612 ( .A(p_input[23876]), .B(p_input[13876]), .Z(n6806) );
  AND U13613 ( .A(n6807), .B(p_input[3875]), .Z(o[3875]) );
  AND U13614 ( .A(p_input[23875]), .B(p_input[13875]), .Z(n6807) );
  AND U13615 ( .A(n6808), .B(p_input[3874]), .Z(o[3874]) );
  AND U13616 ( .A(p_input[23874]), .B(p_input[13874]), .Z(n6808) );
  AND U13617 ( .A(n6809), .B(p_input[3873]), .Z(o[3873]) );
  AND U13618 ( .A(p_input[23873]), .B(p_input[13873]), .Z(n6809) );
  AND U13619 ( .A(n6810), .B(p_input[3872]), .Z(o[3872]) );
  AND U13620 ( .A(p_input[23872]), .B(p_input[13872]), .Z(n6810) );
  AND U13621 ( .A(n6811), .B(p_input[3871]), .Z(o[3871]) );
  AND U13622 ( .A(p_input[23871]), .B(p_input[13871]), .Z(n6811) );
  AND U13623 ( .A(n6812), .B(p_input[3870]), .Z(o[3870]) );
  AND U13624 ( .A(p_input[23870]), .B(p_input[13870]), .Z(n6812) );
  AND U13625 ( .A(n6813), .B(p_input[386]), .Z(o[386]) );
  AND U13626 ( .A(p_input[20386]), .B(p_input[10386]), .Z(n6813) );
  AND U13627 ( .A(n6814), .B(p_input[3869]), .Z(o[3869]) );
  AND U13628 ( .A(p_input[23869]), .B(p_input[13869]), .Z(n6814) );
  AND U13629 ( .A(n6815), .B(p_input[3868]), .Z(o[3868]) );
  AND U13630 ( .A(p_input[23868]), .B(p_input[13868]), .Z(n6815) );
  AND U13631 ( .A(n6816), .B(p_input[3867]), .Z(o[3867]) );
  AND U13632 ( .A(p_input[23867]), .B(p_input[13867]), .Z(n6816) );
  AND U13633 ( .A(n6817), .B(p_input[3866]), .Z(o[3866]) );
  AND U13634 ( .A(p_input[23866]), .B(p_input[13866]), .Z(n6817) );
  AND U13635 ( .A(n6818), .B(p_input[3865]), .Z(o[3865]) );
  AND U13636 ( .A(p_input[23865]), .B(p_input[13865]), .Z(n6818) );
  AND U13637 ( .A(n6819), .B(p_input[3864]), .Z(o[3864]) );
  AND U13638 ( .A(p_input[23864]), .B(p_input[13864]), .Z(n6819) );
  AND U13639 ( .A(n6820), .B(p_input[3863]), .Z(o[3863]) );
  AND U13640 ( .A(p_input[23863]), .B(p_input[13863]), .Z(n6820) );
  AND U13641 ( .A(n6821), .B(p_input[3862]), .Z(o[3862]) );
  AND U13642 ( .A(p_input[23862]), .B(p_input[13862]), .Z(n6821) );
  AND U13643 ( .A(n6822), .B(p_input[3861]), .Z(o[3861]) );
  AND U13644 ( .A(p_input[23861]), .B(p_input[13861]), .Z(n6822) );
  AND U13645 ( .A(n6823), .B(p_input[3860]), .Z(o[3860]) );
  AND U13646 ( .A(p_input[23860]), .B(p_input[13860]), .Z(n6823) );
  AND U13647 ( .A(n6824), .B(p_input[385]), .Z(o[385]) );
  AND U13648 ( .A(p_input[20385]), .B(p_input[10385]), .Z(n6824) );
  AND U13649 ( .A(n6825), .B(p_input[3859]), .Z(o[3859]) );
  AND U13650 ( .A(p_input[23859]), .B(p_input[13859]), .Z(n6825) );
  AND U13651 ( .A(n6826), .B(p_input[3858]), .Z(o[3858]) );
  AND U13652 ( .A(p_input[23858]), .B(p_input[13858]), .Z(n6826) );
  AND U13653 ( .A(n6827), .B(p_input[3857]), .Z(o[3857]) );
  AND U13654 ( .A(p_input[23857]), .B(p_input[13857]), .Z(n6827) );
  AND U13655 ( .A(n6828), .B(p_input[3856]), .Z(o[3856]) );
  AND U13656 ( .A(p_input[23856]), .B(p_input[13856]), .Z(n6828) );
  AND U13657 ( .A(n6829), .B(p_input[3855]), .Z(o[3855]) );
  AND U13658 ( .A(p_input[23855]), .B(p_input[13855]), .Z(n6829) );
  AND U13659 ( .A(n6830), .B(p_input[3854]), .Z(o[3854]) );
  AND U13660 ( .A(p_input[23854]), .B(p_input[13854]), .Z(n6830) );
  AND U13661 ( .A(n6831), .B(p_input[3853]), .Z(o[3853]) );
  AND U13662 ( .A(p_input[23853]), .B(p_input[13853]), .Z(n6831) );
  AND U13663 ( .A(n6832), .B(p_input[3852]), .Z(o[3852]) );
  AND U13664 ( .A(p_input[23852]), .B(p_input[13852]), .Z(n6832) );
  AND U13665 ( .A(n6833), .B(p_input[3851]), .Z(o[3851]) );
  AND U13666 ( .A(p_input[23851]), .B(p_input[13851]), .Z(n6833) );
  AND U13667 ( .A(n6834), .B(p_input[3850]), .Z(o[3850]) );
  AND U13668 ( .A(p_input[23850]), .B(p_input[13850]), .Z(n6834) );
  AND U13669 ( .A(n6835), .B(p_input[384]), .Z(o[384]) );
  AND U13670 ( .A(p_input[20384]), .B(p_input[10384]), .Z(n6835) );
  AND U13671 ( .A(n6836), .B(p_input[3849]), .Z(o[3849]) );
  AND U13672 ( .A(p_input[23849]), .B(p_input[13849]), .Z(n6836) );
  AND U13673 ( .A(n6837), .B(p_input[3848]), .Z(o[3848]) );
  AND U13674 ( .A(p_input[23848]), .B(p_input[13848]), .Z(n6837) );
  AND U13675 ( .A(n6838), .B(p_input[3847]), .Z(o[3847]) );
  AND U13676 ( .A(p_input[23847]), .B(p_input[13847]), .Z(n6838) );
  AND U13677 ( .A(n6839), .B(p_input[3846]), .Z(o[3846]) );
  AND U13678 ( .A(p_input[23846]), .B(p_input[13846]), .Z(n6839) );
  AND U13679 ( .A(n6840), .B(p_input[3845]), .Z(o[3845]) );
  AND U13680 ( .A(p_input[23845]), .B(p_input[13845]), .Z(n6840) );
  AND U13681 ( .A(n6841), .B(p_input[3844]), .Z(o[3844]) );
  AND U13682 ( .A(p_input[23844]), .B(p_input[13844]), .Z(n6841) );
  AND U13683 ( .A(n6842), .B(p_input[3843]), .Z(o[3843]) );
  AND U13684 ( .A(p_input[23843]), .B(p_input[13843]), .Z(n6842) );
  AND U13685 ( .A(n6843), .B(p_input[3842]), .Z(o[3842]) );
  AND U13686 ( .A(p_input[23842]), .B(p_input[13842]), .Z(n6843) );
  AND U13687 ( .A(n6844), .B(p_input[3841]), .Z(o[3841]) );
  AND U13688 ( .A(p_input[23841]), .B(p_input[13841]), .Z(n6844) );
  AND U13689 ( .A(n6845), .B(p_input[3840]), .Z(o[3840]) );
  AND U13690 ( .A(p_input[23840]), .B(p_input[13840]), .Z(n6845) );
  AND U13691 ( .A(n6846), .B(p_input[383]), .Z(o[383]) );
  AND U13692 ( .A(p_input[20383]), .B(p_input[10383]), .Z(n6846) );
  AND U13693 ( .A(n6847), .B(p_input[3839]), .Z(o[3839]) );
  AND U13694 ( .A(p_input[23839]), .B(p_input[13839]), .Z(n6847) );
  AND U13695 ( .A(n6848), .B(p_input[3838]), .Z(o[3838]) );
  AND U13696 ( .A(p_input[23838]), .B(p_input[13838]), .Z(n6848) );
  AND U13697 ( .A(n6849), .B(p_input[3837]), .Z(o[3837]) );
  AND U13698 ( .A(p_input[23837]), .B(p_input[13837]), .Z(n6849) );
  AND U13699 ( .A(n6850), .B(p_input[3836]), .Z(o[3836]) );
  AND U13700 ( .A(p_input[23836]), .B(p_input[13836]), .Z(n6850) );
  AND U13701 ( .A(n6851), .B(p_input[3835]), .Z(o[3835]) );
  AND U13702 ( .A(p_input[23835]), .B(p_input[13835]), .Z(n6851) );
  AND U13703 ( .A(n6852), .B(p_input[3834]), .Z(o[3834]) );
  AND U13704 ( .A(p_input[23834]), .B(p_input[13834]), .Z(n6852) );
  AND U13705 ( .A(n6853), .B(p_input[3833]), .Z(o[3833]) );
  AND U13706 ( .A(p_input[23833]), .B(p_input[13833]), .Z(n6853) );
  AND U13707 ( .A(n6854), .B(p_input[3832]), .Z(o[3832]) );
  AND U13708 ( .A(p_input[23832]), .B(p_input[13832]), .Z(n6854) );
  AND U13709 ( .A(n6855), .B(p_input[3831]), .Z(o[3831]) );
  AND U13710 ( .A(p_input[23831]), .B(p_input[13831]), .Z(n6855) );
  AND U13711 ( .A(n6856), .B(p_input[3830]), .Z(o[3830]) );
  AND U13712 ( .A(p_input[23830]), .B(p_input[13830]), .Z(n6856) );
  AND U13713 ( .A(n6857), .B(p_input[382]), .Z(o[382]) );
  AND U13714 ( .A(p_input[20382]), .B(p_input[10382]), .Z(n6857) );
  AND U13715 ( .A(n6858), .B(p_input[3829]), .Z(o[3829]) );
  AND U13716 ( .A(p_input[23829]), .B(p_input[13829]), .Z(n6858) );
  AND U13717 ( .A(n6859), .B(p_input[3828]), .Z(o[3828]) );
  AND U13718 ( .A(p_input[23828]), .B(p_input[13828]), .Z(n6859) );
  AND U13719 ( .A(n6860), .B(p_input[3827]), .Z(o[3827]) );
  AND U13720 ( .A(p_input[23827]), .B(p_input[13827]), .Z(n6860) );
  AND U13721 ( .A(n6861), .B(p_input[3826]), .Z(o[3826]) );
  AND U13722 ( .A(p_input[23826]), .B(p_input[13826]), .Z(n6861) );
  AND U13723 ( .A(n6862), .B(p_input[3825]), .Z(o[3825]) );
  AND U13724 ( .A(p_input[23825]), .B(p_input[13825]), .Z(n6862) );
  AND U13725 ( .A(n6863), .B(p_input[3824]), .Z(o[3824]) );
  AND U13726 ( .A(p_input[23824]), .B(p_input[13824]), .Z(n6863) );
  AND U13727 ( .A(n6864), .B(p_input[3823]), .Z(o[3823]) );
  AND U13728 ( .A(p_input[23823]), .B(p_input[13823]), .Z(n6864) );
  AND U13729 ( .A(n6865), .B(p_input[3822]), .Z(o[3822]) );
  AND U13730 ( .A(p_input[23822]), .B(p_input[13822]), .Z(n6865) );
  AND U13731 ( .A(n6866), .B(p_input[3821]), .Z(o[3821]) );
  AND U13732 ( .A(p_input[23821]), .B(p_input[13821]), .Z(n6866) );
  AND U13733 ( .A(n6867), .B(p_input[3820]), .Z(o[3820]) );
  AND U13734 ( .A(p_input[23820]), .B(p_input[13820]), .Z(n6867) );
  AND U13735 ( .A(n6868), .B(p_input[381]), .Z(o[381]) );
  AND U13736 ( .A(p_input[20381]), .B(p_input[10381]), .Z(n6868) );
  AND U13737 ( .A(n6869), .B(p_input[3819]), .Z(o[3819]) );
  AND U13738 ( .A(p_input[23819]), .B(p_input[13819]), .Z(n6869) );
  AND U13739 ( .A(n6870), .B(p_input[3818]), .Z(o[3818]) );
  AND U13740 ( .A(p_input[23818]), .B(p_input[13818]), .Z(n6870) );
  AND U13741 ( .A(n6871), .B(p_input[3817]), .Z(o[3817]) );
  AND U13742 ( .A(p_input[23817]), .B(p_input[13817]), .Z(n6871) );
  AND U13743 ( .A(n6872), .B(p_input[3816]), .Z(o[3816]) );
  AND U13744 ( .A(p_input[23816]), .B(p_input[13816]), .Z(n6872) );
  AND U13745 ( .A(n6873), .B(p_input[3815]), .Z(o[3815]) );
  AND U13746 ( .A(p_input[23815]), .B(p_input[13815]), .Z(n6873) );
  AND U13747 ( .A(n6874), .B(p_input[3814]), .Z(o[3814]) );
  AND U13748 ( .A(p_input[23814]), .B(p_input[13814]), .Z(n6874) );
  AND U13749 ( .A(n6875), .B(p_input[3813]), .Z(o[3813]) );
  AND U13750 ( .A(p_input[23813]), .B(p_input[13813]), .Z(n6875) );
  AND U13751 ( .A(n6876), .B(p_input[3812]), .Z(o[3812]) );
  AND U13752 ( .A(p_input[23812]), .B(p_input[13812]), .Z(n6876) );
  AND U13753 ( .A(n6877), .B(p_input[3811]), .Z(o[3811]) );
  AND U13754 ( .A(p_input[23811]), .B(p_input[13811]), .Z(n6877) );
  AND U13755 ( .A(n6878), .B(p_input[3810]), .Z(o[3810]) );
  AND U13756 ( .A(p_input[23810]), .B(p_input[13810]), .Z(n6878) );
  AND U13757 ( .A(n6879), .B(p_input[380]), .Z(o[380]) );
  AND U13758 ( .A(p_input[20380]), .B(p_input[10380]), .Z(n6879) );
  AND U13759 ( .A(n6880), .B(p_input[3809]), .Z(o[3809]) );
  AND U13760 ( .A(p_input[23809]), .B(p_input[13809]), .Z(n6880) );
  AND U13761 ( .A(n6881), .B(p_input[3808]), .Z(o[3808]) );
  AND U13762 ( .A(p_input[23808]), .B(p_input[13808]), .Z(n6881) );
  AND U13763 ( .A(n6882), .B(p_input[3807]), .Z(o[3807]) );
  AND U13764 ( .A(p_input[23807]), .B(p_input[13807]), .Z(n6882) );
  AND U13765 ( .A(n6883), .B(p_input[3806]), .Z(o[3806]) );
  AND U13766 ( .A(p_input[23806]), .B(p_input[13806]), .Z(n6883) );
  AND U13767 ( .A(n6884), .B(p_input[3805]), .Z(o[3805]) );
  AND U13768 ( .A(p_input[23805]), .B(p_input[13805]), .Z(n6884) );
  AND U13769 ( .A(n6885), .B(p_input[3804]), .Z(o[3804]) );
  AND U13770 ( .A(p_input[23804]), .B(p_input[13804]), .Z(n6885) );
  AND U13771 ( .A(n6886), .B(p_input[3803]), .Z(o[3803]) );
  AND U13772 ( .A(p_input[23803]), .B(p_input[13803]), .Z(n6886) );
  AND U13773 ( .A(n6887), .B(p_input[3802]), .Z(o[3802]) );
  AND U13774 ( .A(p_input[23802]), .B(p_input[13802]), .Z(n6887) );
  AND U13775 ( .A(n6888), .B(p_input[3801]), .Z(o[3801]) );
  AND U13776 ( .A(p_input[23801]), .B(p_input[13801]), .Z(n6888) );
  AND U13777 ( .A(n6889), .B(p_input[3800]), .Z(o[3800]) );
  AND U13778 ( .A(p_input[23800]), .B(p_input[13800]), .Z(n6889) );
  AND U13779 ( .A(n6890), .B(p_input[37]), .Z(o[37]) );
  AND U13780 ( .A(p_input[20037]), .B(p_input[10037]), .Z(n6890) );
  AND U13781 ( .A(n6891), .B(p_input[379]), .Z(o[379]) );
  AND U13782 ( .A(p_input[20379]), .B(p_input[10379]), .Z(n6891) );
  AND U13783 ( .A(n6892), .B(p_input[3799]), .Z(o[3799]) );
  AND U13784 ( .A(p_input[23799]), .B(p_input[13799]), .Z(n6892) );
  AND U13785 ( .A(n6893), .B(p_input[3798]), .Z(o[3798]) );
  AND U13786 ( .A(p_input[23798]), .B(p_input[13798]), .Z(n6893) );
  AND U13787 ( .A(n6894), .B(p_input[3797]), .Z(o[3797]) );
  AND U13788 ( .A(p_input[23797]), .B(p_input[13797]), .Z(n6894) );
  AND U13789 ( .A(n6895), .B(p_input[3796]), .Z(o[3796]) );
  AND U13790 ( .A(p_input[23796]), .B(p_input[13796]), .Z(n6895) );
  AND U13791 ( .A(n6896), .B(p_input[3795]), .Z(o[3795]) );
  AND U13792 ( .A(p_input[23795]), .B(p_input[13795]), .Z(n6896) );
  AND U13793 ( .A(n6897), .B(p_input[3794]), .Z(o[3794]) );
  AND U13794 ( .A(p_input[23794]), .B(p_input[13794]), .Z(n6897) );
  AND U13795 ( .A(n6898), .B(p_input[3793]), .Z(o[3793]) );
  AND U13796 ( .A(p_input[23793]), .B(p_input[13793]), .Z(n6898) );
  AND U13797 ( .A(n6899), .B(p_input[3792]), .Z(o[3792]) );
  AND U13798 ( .A(p_input[23792]), .B(p_input[13792]), .Z(n6899) );
  AND U13799 ( .A(n6900), .B(p_input[3791]), .Z(o[3791]) );
  AND U13800 ( .A(p_input[23791]), .B(p_input[13791]), .Z(n6900) );
  AND U13801 ( .A(n6901), .B(p_input[3790]), .Z(o[3790]) );
  AND U13802 ( .A(p_input[23790]), .B(p_input[13790]), .Z(n6901) );
  AND U13803 ( .A(n6902), .B(p_input[378]), .Z(o[378]) );
  AND U13804 ( .A(p_input[20378]), .B(p_input[10378]), .Z(n6902) );
  AND U13805 ( .A(n6903), .B(p_input[3789]), .Z(o[3789]) );
  AND U13806 ( .A(p_input[23789]), .B(p_input[13789]), .Z(n6903) );
  AND U13807 ( .A(n6904), .B(p_input[3788]), .Z(o[3788]) );
  AND U13808 ( .A(p_input[23788]), .B(p_input[13788]), .Z(n6904) );
  AND U13809 ( .A(n6905), .B(p_input[3787]), .Z(o[3787]) );
  AND U13810 ( .A(p_input[23787]), .B(p_input[13787]), .Z(n6905) );
  AND U13811 ( .A(n6906), .B(p_input[3786]), .Z(o[3786]) );
  AND U13812 ( .A(p_input[23786]), .B(p_input[13786]), .Z(n6906) );
  AND U13813 ( .A(n6907), .B(p_input[3785]), .Z(o[3785]) );
  AND U13814 ( .A(p_input[23785]), .B(p_input[13785]), .Z(n6907) );
  AND U13815 ( .A(n6908), .B(p_input[3784]), .Z(o[3784]) );
  AND U13816 ( .A(p_input[23784]), .B(p_input[13784]), .Z(n6908) );
  AND U13817 ( .A(n6909), .B(p_input[3783]), .Z(o[3783]) );
  AND U13818 ( .A(p_input[23783]), .B(p_input[13783]), .Z(n6909) );
  AND U13819 ( .A(n6910), .B(p_input[3782]), .Z(o[3782]) );
  AND U13820 ( .A(p_input[23782]), .B(p_input[13782]), .Z(n6910) );
  AND U13821 ( .A(n6911), .B(p_input[3781]), .Z(o[3781]) );
  AND U13822 ( .A(p_input[23781]), .B(p_input[13781]), .Z(n6911) );
  AND U13823 ( .A(n6912), .B(p_input[3780]), .Z(o[3780]) );
  AND U13824 ( .A(p_input[23780]), .B(p_input[13780]), .Z(n6912) );
  AND U13825 ( .A(n6913), .B(p_input[377]), .Z(o[377]) );
  AND U13826 ( .A(p_input[20377]), .B(p_input[10377]), .Z(n6913) );
  AND U13827 ( .A(n6914), .B(p_input[3779]), .Z(o[3779]) );
  AND U13828 ( .A(p_input[23779]), .B(p_input[13779]), .Z(n6914) );
  AND U13829 ( .A(n6915), .B(p_input[3778]), .Z(o[3778]) );
  AND U13830 ( .A(p_input[23778]), .B(p_input[13778]), .Z(n6915) );
  AND U13831 ( .A(n6916), .B(p_input[3777]), .Z(o[3777]) );
  AND U13832 ( .A(p_input[23777]), .B(p_input[13777]), .Z(n6916) );
  AND U13833 ( .A(n6917), .B(p_input[3776]), .Z(o[3776]) );
  AND U13834 ( .A(p_input[23776]), .B(p_input[13776]), .Z(n6917) );
  AND U13835 ( .A(n6918), .B(p_input[3775]), .Z(o[3775]) );
  AND U13836 ( .A(p_input[23775]), .B(p_input[13775]), .Z(n6918) );
  AND U13837 ( .A(n6919), .B(p_input[3774]), .Z(o[3774]) );
  AND U13838 ( .A(p_input[23774]), .B(p_input[13774]), .Z(n6919) );
  AND U13839 ( .A(n6920), .B(p_input[3773]), .Z(o[3773]) );
  AND U13840 ( .A(p_input[23773]), .B(p_input[13773]), .Z(n6920) );
  AND U13841 ( .A(n6921), .B(p_input[3772]), .Z(o[3772]) );
  AND U13842 ( .A(p_input[23772]), .B(p_input[13772]), .Z(n6921) );
  AND U13843 ( .A(n6922), .B(p_input[3771]), .Z(o[3771]) );
  AND U13844 ( .A(p_input[23771]), .B(p_input[13771]), .Z(n6922) );
  AND U13845 ( .A(n6923), .B(p_input[3770]), .Z(o[3770]) );
  AND U13846 ( .A(p_input[23770]), .B(p_input[13770]), .Z(n6923) );
  AND U13847 ( .A(n6924), .B(p_input[376]), .Z(o[376]) );
  AND U13848 ( .A(p_input[20376]), .B(p_input[10376]), .Z(n6924) );
  AND U13849 ( .A(n6925), .B(p_input[3769]), .Z(o[3769]) );
  AND U13850 ( .A(p_input[23769]), .B(p_input[13769]), .Z(n6925) );
  AND U13851 ( .A(n6926), .B(p_input[3768]), .Z(o[3768]) );
  AND U13852 ( .A(p_input[23768]), .B(p_input[13768]), .Z(n6926) );
  AND U13853 ( .A(n6927), .B(p_input[3767]), .Z(o[3767]) );
  AND U13854 ( .A(p_input[23767]), .B(p_input[13767]), .Z(n6927) );
  AND U13855 ( .A(n6928), .B(p_input[3766]), .Z(o[3766]) );
  AND U13856 ( .A(p_input[23766]), .B(p_input[13766]), .Z(n6928) );
  AND U13857 ( .A(n6929), .B(p_input[3765]), .Z(o[3765]) );
  AND U13858 ( .A(p_input[23765]), .B(p_input[13765]), .Z(n6929) );
  AND U13859 ( .A(n6930), .B(p_input[3764]), .Z(o[3764]) );
  AND U13860 ( .A(p_input[23764]), .B(p_input[13764]), .Z(n6930) );
  AND U13861 ( .A(n6931), .B(p_input[3763]), .Z(o[3763]) );
  AND U13862 ( .A(p_input[23763]), .B(p_input[13763]), .Z(n6931) );
  AND U13863 ( .A(n6932), .B(p_input[3762]), .Z(o[3762]) );
  AND U13864 ( .A(p_input[23762]), .B(p_input[13762]), .Z(n6932) );
  AND U13865 ( .A(n6933), .B(p_input[3761]), .Z(o[3761]) );
  AND U13866 ( .A(p_input[23761]), .B(p_input[13761]), .Z(n6933) );
  AND U13867 ( .A(n6934), .B(p_input[3760]), .Z(o[3760]) );
  AND U13868 ( .A(p_input[23760]), .B(p_input[13760]), .Z(n6934) );
  AND U13869 ( .A(n6935), .B(p_input[375]), .Z(o[375]) );
  AND U13870 ( .A(p_input[20375]), .B(p_input[10375]), .Z(n6935) );
  AND U13871 ( .A(n6936), .B(p_input[3759]), .Z(o[3759]) );
  AND U13872 ( .A(p_input[23759]), .B(p_input[13759]), .Z(n6936) );
  AND U13873 ( .A(n6937), .B(p_input[3758]), .Z(o[3758]) );
  AND U13874 ( .A(p_input[23758]), .B(p_input[13758]), .Z(n6937) );
  AND U13875 ( .A(n6938), .B(p_input[3757]), .Z(o[3757]) );
  AND U13876 ( .A(p_input[23757]), .B(p_input[13757]), .Z(n6938) );
  AND U13877 ( .A(n6939), .B(p_input[3756]), .Z(o[3756]) );
  AND U13878 ( .A(p_input[23756]), .B(p_input[13756]), .Z(n6939) );
  AND U13879 ( .A(n6940), .B(p_input[3755]), .Z(o[3755]) );
  AND U13880 ( .A(p_input[23755]), .B(p_input[13755]), .Z(n6940) );
  AND U13881 ( .A(n6941), .B(p_input[3754]), .Z(o[3754]) );
  AND U13882 ( .A(p_input[23754]), .B(p_input[13754]), .Z(n6941) );
  AND U13883 ( .A(n6942), .B(p_input[3753]), .Z(o[3753]) );
  AND U13884 ( .A(p_input[23753]), .B(p_input[13753]), .Z(n6942) );
  AND U13885 ( .A(n6943), .B(p_input[3752]), .Z(o[3752]) );
  AND U13886 ( .A(p_input[23752]), .B(p_input[13752]), .Z(n6943) );
  AND U13887 ( .A(n6944), .B(p_input[3751]), .Z(o[3751]) );
  AND U13888 ( .A(p_input[23751]), .B(p_input[13751]), .Z(n6944) );
  AND U13889 ( .A(n6945), .B(p_input[3750]), .Z(o[3750]) );
  AND U13890 ( .A(p_input[23750]), .B(p_input[13750]), .Z(n6945) );
  AND U13891 ( .A(n6946), .B(p_input[374]), .Z(o[374]) );
  AND U13892 ( .A(p_input[20374]), .B(p_input[10374]), .Z(n6946) );
  AND U13893 ( .A(n6947), .B(p_input[3749]), .Z(o[3749]) );
  AND U13894 ( .A(p_input[23749]), .B(p_input[13749]), .Z(n6947) );
  AND U13895 ( .A(n6948), .B(p_input[3748]), .Z(o[3748]) );
  AND U13896 ( .A(p_input[23748]), .B(p_input[13748]), .Z(n6948) );
  AND U13897 ( .A(n6949), .B(p_input[3747]), .Z(o[3747]) );
  AND U13898 ( .A(p_input[23747]), .B(p_input[13747]), .Z(n6949) );
  AND U13899 ( .A(n6950), .B(p_input[3746]), .Z(o[3746]) );
  AND U13900 ( .A(p_input[23746]), .B(p_input[13746]), .Z(n6950) );
  AND U13901 ( .A(n6951), .B(p_input[3745]), .Z(o[3745]) );
  AND U13902 ( .A(p_input[23745]), .B(p_input[13745]), .Z(n6951) );
  AND U13903 ( .A(n6952), .B(p_input[3744]), .Z(o[3744]) );
  AND U13904 ( .A(p_input[23744]), .B(p_input[13744]), .Z(n6952) );
  AND U13905 ( .A(n6953), .B(p_input[3743]), .Z(o[3743]) );
  AND U13906 ( .A(p_input[23743]), .B(p_input[13743]), .Z(n6953) );
  AND U13907 ( .A(n6954), .B(p_input[3742]), .Z(o[3742]) );
  AND U13908 ( .A(p_input[23742]), .B(p_input[13742]), .Z(n6954) );
  AND U13909 ( .A(n6955), .B(p_input[3741]), .Z(o[3741]) );
  AND U13910 ( .A(p_input[23741]), .B(p_input[13741]), .Z(n6955) );
  AND U13911 ( .A(n6956), .B(p_input[3740]), .Z(o[3740]) );
  AND U13912 ( .A(p_input[23740]), .B(p_input[13740]), .Z(n6956) );
  AND U13913 ( .A(n6957), .B(p_input[373]), .Z(o[373]) );
  AND U13914 ( .A(p_input[20373]), .B(p_input[10373]), .Z(n6957) );
  AND U13915 ( .A(n6958), .B(p_input[3739]), .Z(o[3739]) );
  AND U13916 ( .A(p_input[23739]), .B(p_input[13739]), .Z(n6958) );
  AND U13917 ( .A(n6959), .B(p_input[3738]), .Z(o[3738]) );
  AND U13918 ( .A(p_input[23738]), .B(p_input[13738]), .Z(n6959) );
  AND U13919 ( .A(n6960), .B(p_input[3737]), .Z(o[3737]) );
  AND U13920 ( .A(p_input[23737]), .B(p_input[13737]), .Z(n6960) );
  AND U13921 ( .A(n6961), .B(p_input[3736]), .Z(o[3736]) );
  AND U13922 ( .A(p_input[23736]), .B(p_input[13736]), .Z(n6961) );
  AND U13923 ( .A(n6962), .B(p_input[3735]), .Z(o[3735]) );
  AND U13924 ( .A(p_input[23735]), .B(p_input[13735]), .Z(n6962) );
  AND U13925 ( .A(n6963), .B(p_input[3734]), .Z(o[3734]) );
  AND U13926 ( .A(p_input[23734]), .B(p_input[13734]), .Z(n6963) );
  AND U13927 ( .A(n6964), .B(p_input[3733]), .Z(o[3733]) );
  AND U13928 ( .A(p_input[23733]), .B(p_input[13733]), .Z(n6964) );
  AND U13929 ( .A(n6965), .B(p_input[3732]), .Z(o[3732]) );
  AND U13930 ( .A(p_input[23732]), .B(p_input[13732]), .Z(n6965) );
  AND U13931 ( .A(n6966), .B(p_input[3731]), .Z(o[3731]) );
  AND U13932 ( .A(p_input[23731]), .B(p_input[13731]), .Z(n6966) );
  AND U13933 ( .A(n6967), .B(p_input[3730]), .Z(o[3730]) );
  AND U13934 ( .A(p_input[23730]), .B(p_input[13730]), .Z(n6967) );
  AND U13935 ( .A(n6968), .B(p_input[372]), .Z(o[372]) );
  AND U13936 ( .A(p_input[20372]), .B(p_input[10372]), .Z(n6968) );
  AND U13937 ( .A(n6969), .B(p_input[3729]), .Z(o[3729]) );
  AND U13938 ( .A(p_input[23729]), .B(p_input[13729]), .Z(n6969) );
  AND U13939 ( .A(n6970), .B(p_input[3728]), .Z(o[3728]) );
  AND U13940 ( .A(p_input[23728]), .B(p_input[13728]), .Z(n6970) );
  AND U13941 ( .A(n6971), .B(p_input[3727]), .Z(o[3727]) );
  AND U13942 ( .A(p_input[23727]), .B(p_input[13727]), .Z(n6971) );
  AND U13943 ( .A(n6972), .B(p_input[3726]), .Z(o[3726]) );
  AND U13944 ( .A(p_input[23726]), .B(p_input[13726]), .Z(n6972) );
  AND U13945 ( .A(n6973), .B(p_input[3725]), .Z(o[3725]) );
  AND U13946 ( .A(p_input[23725]), .B(p_input[13725]), .Z(n6973) );
  AND U13947 ( .A(n6974), .B(p_input[3724]), .Z(o[3724]) );
  AND U13948 ( .A(p_input[23724]), .B(p_input[13724]), .Z(n6974) );
  AND U13949 ( .A(n6975), .B(p_input[3723]), .Z(o[3723]) );
  AND U13950 ( .A(p_input[23723]), .B(p_input[13723]), .Z(n6975) );
  AND U13951 ( .A(n6976), .B(p_input[3722]), .Z(o[3722]) );
  AND U13952 ( .A(p_input[23722]), .B(p_input[13722]), .Z(n6976) );
  AND U13953 ( .A(n6977), .B(p_input[3721]), .Z(o[3721]) );
  AND U13954 ( .A(p_input[23721]), .B(p_input[13721]), .Z(n6977) );
  AND U13955 ( .A(n6978), .B(p_input[3720]), .Z(o[3720]) );
  AND U13956 ( .A(p_input[23720]), .B(p_input[13720]), .Z(n6978) );
  AND U13957 ( .A(n6979), .B(p_input[371]), .Z(o[371]) );
  AND U13958 ( .A(p_input[20371]), .B(p_input[10371]), .Z(n6979) );
  AND U13959 ( .A(n6980), .B(p_input[3719]), .Z(o[3719]) );
  AND U13960 ( .A(p_input[23719]), .B(p_input[13719]), .Z(n6980) );
  AND U13961 ( .A(n6981), .B(p_input[3718]), .Z(o[3718]) );
  AND U13962 ( .A(p_input[23718]), .B(p_input[13718]), .Z(n6981) );
  AND U13963 ( .A(n6982), .B(p_input[3717]), .Z(o[3717]) );
  AND U13964 ( .A(p_input[23717]), .B(p_input[13717]), .Z(n6982) );
  AND U13965 ( .A(n6983), .B(p_input[3716]), .Z(o[3716]) );
  AND U13966 ( .A(p_input[23716]), .B(p_input[13716]), .Z(n6983) );
  AND U13967 ( .A(n6984), .B(p_input[3715]), .Z(o[3715]) );
  AND U13968 ( .A(p_input[23715]), .B(p_input[13715]), .Z(n6984) );
  AND U13969 ( .A(n6985), .B(p_input[3714]), .Z(o[3714]) );
  AND U13970 ( .A(p_input[23714]), .B(p_input[13714]), .Z(n6985) );
  AND U13971 ( .A(n6986), .B(p_input[3713]), .Z(o[3713]) );
  AND U13972 ( .A(p_input[23713]), .B(p_input[13713]), .Z(n6986) );
  AND U13973 ( .A(n6987), .B(p_input[3712]), .Z(o[3712]) );
  AND U13974 ( .A(p_input[23712]), .B(p_input[13712]), .Z(n6987) );
  AND U13975 ( .A(n6988), .B(p_input[3711]), .Z(o[3711]) );
  AND U13976 ( .A(p_input[23711]), .B(p_input[13711]), .Z(n6988) );
  AND U13977 ( .A(n6989), .B(p_input[3710]), .Z(o[3710]) );
  AND U13978 ( .A(p_input[23710]), .B(p_input[13710]), .Z(n6989) );
  AND U13979 ( .A(n6990), .B(p_input[370]), .Z(o[370]) );
  AND U13980 ( .A(p_input[20370]), .B(p_input[10370]), .Z(n6990) );
  AND U13981 ( .A(n6991), .B(p_input[3709]), .Z(o[3709]) );
  AND U13982 ( .A(p_input[23709]), .B(p_input[13709]), .Z(n6991) );
  AND U13983 ( .A(n6992), .B(p_input[3708]), .Z(o[3708]) );
  AND U13984 ( .A(p_input[23708]), .B(p_input[13708]), .Z(n6992) );
  AND U13985 ( .A(n6993), .B(p_input[3707]), .Z(o[3707]) );
  AND U13986 ( .A(p_input[23707]), .B(p_input[13707]), .Z(n6993) );
  AND U13987 ( .A(n6994), .B(p_input[3706]), .Z(o[3706]) );
  AND U13988 ( .A(p_input[23706]), .B(p_input[13706]), .Z(n6994) );
  AND U13989 ( .A(n6995), .B(p_input[3705]), .Z(o[3705]) );
  AND U13990 ( .A(p_input[23705]), .B(p_input[13705]), .Z(n6995) );
  AND U13991 ( .A(n6996), .B(p_input[3704]), .Z(o[3704]) );
  AND U13992 ( .A(p_input[23704]), .B(p_input[13704]), .Z(n6996) );
  AND U13993 ( .A(n6997), .B(p_input[3703]), .Z(o[3703]) );
  AND U13994 ( .A(p_input[23703]), .B(p_input[13703]), .Z(n6997) );
  AND U13995 ( .A(n6998), .B(p_input[3702]), .Z(o[3702]) );
  AND U13996 ( .A(p_input[23702]), .B(p_input[13702]), .Z(n6998) );
  AND U13997 ( .A(n6999), .B(p_input[3701]), .Z(o[3701]) );
  AND U13998 ( .A(p_input[23701]), .B(p_input[13701]), .Z(n6999) );
  AND U13999 ( .A(n7000), .B(p_input[3700]), .Z(o[3700]) );
  AND U14000 ( .A(p_input[23700]), .B(p_input[13700]), .Z(n7000) );
  AND U14001 ( .A(n7001), .B(p_input[36]), .Z(o[36]) );
  AND U14002 ( .A(p_input[20036]), .B(p_input[10036]), .Z(n7001) );
  AND U14003 ( .A(n7002), .B(p_input[369]), .Z(o[369]) );
  AND U14004 ( .A(p_input[20369]), .B(p_input[10369]), .Z(n7002) );
  AND U14005 ( .A(n7003), .B(p_input[3699]), .Z(o[3699]) );
  AND U14006 ( .A(p_input[23699]), .B(p_input[13699]), .Z(n7003) );
  AND U14007 ( .A(n7004), .B(p_input[3698]), .Z(o[3698]) );
  AND U14008 ( .A(p_input[23698]), .B(p_input[13698]), .Z(n7004) );
  AND U14009 ( .A(n7005), .B(p_input[3697]), .Z(o[3697]) );
  AND U14010 ( .A(p_input[23697]), .B(p_input[13697]), .Z(n7005) );
  AND U14011 ( .A(n7006), .B(p_input[3696]), .Z(o[3696]) );
  AND U14012 ( .A(p_input[23696]), .B(p_input[13696]), .Z(n7006) );
  AND U14013 ( .A(n7007), .B(p_input[3695]), .Z(o[3695]) );
  AND U14014 ( .A(p_input[23695]), .B(p_input[13695]), .Z(n7007) );
  AND U14015 ( .A(n7008), .B(p_input[3694]), .Z(o[3694]) );
  AND U14016 ( .A(p_input[23694]), .B(p_input[13694]), .Z(n7008) );
  AND U14017 ( .A(n7009), .B(p_input[3693]), .Z(o[3693]) );
  AND U14018 ( .A(p_input[23693]), .B(p_input[13693]), .Z(n7009) );
  AND U14019 ( .A(n7010), .B(p_input[3692]), .Z(o[3692]) );
  AND U14020 ( .A(p_input[23692]), .B(p_input[13692]), .Z(n7010) );
  AND U14021 ( .A(n7011), .B(p_input[3691]), .Z(o[3691]) );
  AND U14022 ( .A(p_input[23691]), .B(p_input[13691]), .Z(n7011) );
  AND U14023 ( .A(n7012), .B(p_input[3690]), .Z(o[3690]) );
  AND U14024 ( .A(p_input[23690]), .B(p_input[13690]), .Z(n7012) );
  AND U14025 ( .A(n7013), .B(p_input[368]), .Z(o[368]) );
  AND U14026 ( .A(p_input[20368]), .B(p_input[10368]), .Z(n7013) );
  AND U14027 ( .A(n7014), .B(p_input[3689]), .Z(o[3689]) );
  AND U14028 ( .A(p_input[23689]), .B(p_input[13689]), .Z(n7014) );
  AND U14029 ( .A(n7015), .B(p_input[3688]), .Z(o[3688]) );
  AND U14030 ( .A(p_input[23688]), .B(p_input[13688]), .Z(n7015) );
  AND U14031 ( .A(n7016), .B(p_input[3687]), .Z(o[3687]) );
  AND U14032 ( .A(p_input[23687]), .B(p_input[13687]), .Z(n7016) );
  AND U14033 ( .A(n7017), .B(p_input[3686]), .Z(o[3686]) );
  AND U14034 ( .A(p_input[23686]), .B(p_input[13686]), .Z(n7017) );
  AND U14035 ( .A(n7018), .B(p_input[3685]), .Z(o[3685]) );
  AND U14036 ( .A(p_input[23685]), .B(p_input[13685]), .Z(n7018) );
  AND U14037 ( .A(n7019), .B(p_input[3684]), .Z(o[3684]) );
  AND U14038 ( .A(p_input[23684]), .B(p_input[13684]), .Z(n7019) );
  AND U14039 ( .A(n7020), .B(p_input[3683]), .Z(o[3683]) );
  AND U14040 ( .A(p_input[23683]), .B(p_input[13683]), .Z(n7020) );
  AND U14041 ( .A(n7021), .B(p_input[3682]), .Z(o[3682]) );
  AND U14042 ( .A(p_input[23682]), .B(p_input[13682]), .Z(n7021) );
  AND U14043 ( .A(n7022), .B(p_input[3681]), .Z(o[3681]) );
  AND U14044 ( .A(p_input[23681]), .B(p_input[13681]), .Z(n7022) );
  AND U14045 ( .A(n7023), .B(p_input[3680]), .Z(o[3680]) );
  AND U14046 ( .A(p_input[23680]), .B(p_input[13680]), .Z(n7023) );
  AND U14047 ( .A(n7024), .B(p_input[367]), .Z(o[367]) );
  AND U14048 ( .A(p_input[20367]), .B(p_input[10367]), .Z(n7024) );
  AND U14049 ( .A(n7025), .B(p_input[3679]), .Z(o[3679]) );
  AND U14050 ( .A(p_input[23679]), .B(p_input[13679]), .Z(n7025) );
  AND U14051 ( .A(n7026), .B(p_input[3678]), .Z(o[3678]) );
  AND U14052 ( .A(p_input[23678]), .B(p_input[13678]), .Z(n7026) );
  AND U14053 ( .A(n7027), .B(p_input[3677]), .Z(o[3677]) );
  AND U14054 ( .A(p_input[23677]), .B(p_input[13677]), .Z(n7027) );
  AND U14055 ( .A(n7028), .B(p_input[3676]), .Z(o[3676]) );
  AND U14056 ( .A(p_input[23676]), .B(p_input[13676]), .Z(n7028) );
  AND U14057 ( .A(n7029), .B(p_input[3675]), .Z(o[3675]) );
  AND U14058 ( .A(p_input[23675]), .B(p_input[13675]), .Z(n7029) );
  AND U14059 ( .A(n7030), .B(p_input[3674]), .Z(o[3674]) );
  AND U14060 ( .A(p_input[23674]), .B(p_input[13674]), .Z(n7030) );
  AND U14061 ( .A(n7031), .B(p_input[3673]), .Z(o[3673]) );
  AND U14062 ( .A(p_input[23673]), .B(p_input[13673]), .Z(n7031) );
  AND U14063 ( .A(n7032), .B(p_input[3672]), .Z(o[3672]) );
  AND U14064 ( .A(p_input[23672]), .B(p_input[13672]), .Z(n7032) );
  AND U14065 ( .A(n7033), .B(p_input[3671]), .Z(o[3671]) );
  AND U14066 ( .A(p_input[23671]), .B(p_input[13671]), .Z(n7033) );
  AND U14067 ( .A(n7034), .B(p_input[3670]), .Z(o[3670]) );
  AND U14068 ( .A(p_input[23670]), .B(p_input[13670]), .Z(n7034) );
  AND U14069 ( .A(n7035), .B(p_input[366]), .Z(o[366]) );
  AND U14070 ( .A(p_input[20366]), .B(p_input[10366]), .Z(n7035) );
  AND U14071 ( .A(n7036), .B(p_input[3669]), .Z(o[3669]) );
  AND U14072 ( .A(p_input[23669]), .B(p_input[13669]), .Z(n7036) );
  AND U14073 ( .A(n7037), .B(p_input[3668]), .Z(o[3668]) );
  AND U14074 ( .A(p_input[23668]), .B(p_input[13668]), .Z(n7037) );
  AND U14075 ( .A(n7038), .B(p_input[3667]), .Z(o[3667]) );
  AND U14076 ( .A(p_input[23667]), .B(p_input[13667]), .Z(n7038) );
  AND U14077 ( .A(n7039), .B(p_input[3666]), .Z(o[3666]) );
  AND U14078 ( .A(p_input[23666]), .B(p_input[13666]), .Z(n7039) );
  AND U14079 ( .A(n7040), .B(p_input[3665]), .Z(o[3665]) );
  AND U14080 ( .A(p_input[23665]), .B(p_input[13665]), .Z(n7040) );
  AND U14081 ( .A(n7041), .B(p_input[3664]), .Z(o[3664]) );
  AND U14082 ( .A(p_input[23664]), .B(p_input[13664]), .Z(n7041) );
  AND U14083 ( .A(n7042), .B(p_input[3663]), .Z(o[3663]) );
  AND U14084 ( .A(p_input[23663]), .B(p_input[13663]), .Z(n7042) );
  AND U14085 ( .A(n7043), .B(p_input[3662]), .Z(o[3662]) );
  AND U14086 ( .A(p_input[23662]), .B(p_input[13662]), .Z(n7043) );
  AND U14087 ( .A(n7044), .B(p_input[3661]), .Z(o[3661]) );
  AND U14088 ( .A(p_input[23661]), .B(p_input[13661]), .Z(n7044) );
  AND U14089 ( .A(n7045), .B(p_input[3660]), .Z(o[3660]) );
  AND U14090 ( .A(p_input[23660]), .B(p_input[13660]), .Z(n7045) );
  AND U14091 ( .A(n7046), .B(p_input[365]), .Z(o[365]) );
  AND U14092 ( .A(p_input[20365]), .B(p_input[10365]), .Z(n7046) );
  AND U14093 ( .A(n7047), .B(p_input[3659]), .Z(o[3659]) );
  AND U14094 ( .A(p_input[23659]), .B(p_input[13659]), .Z(n7047) );
  AND U14095 ( .A(n7048), .B(p_input[3658]), .Z(o[3658]) );
  AND U14096 ( .A(p_input[23658]), .B(p_input[13658]), .Z(n7048) );
  AND U14097 ( .A(n7049), .B(p_input[3657]), .Z(o[3657]) );
  AND U14098 ( .A(p_input[23657]), .B(p_input[13657]), .Z(n7049) );
  AND U14099 ( .A(n7050), .B(p_input[3656]), .Z(o[3656]) );
  AND U14100 ( .A(p_input[23656]), .B(p_input[13656]), .Z(n7050) );
  AND U14101 ( .A(n7051), .B(p_input[3655]), .Z(o[3655]) );
  AND U14102 ( .A(p_input[23655]), .B(p_input[13655]), .Z(n7051) );
  AND U14103 ( .A(n7052), .B(p_input[3654]), .Z(o[3654]) );
  AND U14104 ( .A(p_input[23654]), .B(p_input[13654]), .Z(n7052) );
  AND U14105 ( .A(n7053), .B(p_input[3653]), .Z(o[3653]) );
  AND U14106 ( .A(p_input[23653]), .B(p_input[13653]), .Z(n7053) );
  AND U14107 ( .A(n7054), .B(p_input[3652]), .Z(o[3652]) );
  AND U14108 ( .A(p_input[23652]), .B(p_input[13652]), .Z(n7054) );
  AND U14109 ( .A(n7055), .B(p_input[3651]), .Z(o[3651]) );
  AND U14110 ( .A(p_input[23651]), .B(p_input[13651]), .Z(n7055) );
  AND U14111 ( .A(n7056), .B(p_input[3650]), .Z(o[3650]) );
  AND U14112 ( .A(p_input[23650]), .B(p_input[13650]), .Z(n7056) );
  AND U14113 ( .A(n7057), .B(p_input[364]), .Z(o[364]) );
  AND U14114 ( .A(p_input[20364]), .B(p_input[10364]), .Z(n7057) );
  AND U14115 ( .A(n7058), .B(p_input[3649]), .Z(o[3649]) );
  AND U14116 ( .A(p_input[23649]), .B(p_input[13649]), .Z(n7058) );
  AND U14117 ( .A(n7059), .B(p_input[3648]), .Z(o[3648]) );
  AND U14118 ( .A(p_input[23648]), .B(p_input[13648]), .Z(n7059) );
  AND U14119 ( .A(n7060), .B(p_input[3647]), .Z(o[3647]) );
  AND U14120 ( .A(p_input[23647]), .B(p_input[13647]), .Z(n7060) );
  AND U14121 ( .A(n7061), .B(p_input[3646]), .Z(o[3646]) );
  AND U14122 ( .A(p_input[23646]), .B(p_input[13646]), .Z(n7061) );
  AND U14123 ( .A(n7062), .B(p_input[3645]), .Z(o[3645]) );
  AND U14124 ( .A(p_input[23645]), .B(p_input[13645]), .Z(n7062) );
  AND U14125 ( .A(n7063), .B(p_input[3644]), .Z(o[3644]) );
  AND U14126 ( .A(p_input[23644]), .B(p_input[13644]), .Z(n7063) );
  AND U14127 ( .A(n7064), .B(p_input[3643]), .Z(o[3643]) );
  AND U14128 ( .A(p_input[23643]), .B(p_input[13643]), .Z(n7064) );
  AND U14129 ( .A(n7065), .B(p_input[3642]), .Z(o[3642]) );
  AND U14130 ( .A(p_input[23642]), .B(p_input[13642]), .Z(n7065) );
  AND U14131 ( .A(n7066), .B(p_input[3641]), .Z(o[3641]) );
  AND U14132 ( .A(p_input[23641]), .B(p_input[13641]), .Z(n7066) );
  AND U14133 ( .A(n7067), .B(p_input[3640]), .Z(o[3640]) );
  AND U14134 ( .A(p_input[23640]), .B(p_input[13640]), .Z(n7067) );
  AND U14135 ( .A(n7068), .B(p_input[363]), .Z(o[363]) );
  AND U14136 ( .A(p_input[20363]), .B(p_input[10363]), .Z(n7068) );
  AND U14137 ( .A(n7069), .B(p_input[3639]), .Z(o[3639]) );
  AND U14138 ( .A(p_input[23639]), .B(p_input[13639]), .Z(n7069) );
  AND U14139 ( .A(n7070), .B(p_input[3638]), .Z(o[3638]) );
  AND U14140 ( .A(p_input[23638]), .B(p_input[13638]), .Z(n7070) );
  AND U14141 ( .A(n7071), .B(p_input[3637]), .Z(o[3637]) );
  AND U14142 ( .A(p_input[23637]), .B(p_input[13637]), .Z(n7071) );
  AND U14143 ( .A(n7072), .B(p_input[3636]), .Z(o[3636]) );
  AND U14144 ( .A(p_input[23636]), .B(p_input[13636]), .Z(n7072) );
  AND U14145 ( .A(n7073), .B(p_input[3635]), .Z(o[3635]) );
  AND U14146 ( .A(p_input[23635]), .B(p_input[13635]), .Z(n7073) );
  AND U14147 ( .A(n7074), .B(p_input[3634]), .Z(o[3634]) );
  AND U14148 ( .A(p_input[23634]), .B(p_input[13634]), .Z(n7074) );
  AND U14149 ( .A(n7075), .B(p_input[3633]), .Z(o[3633]) );
  AND U14150 ( .A(p_input[23633]), .B(p_input[13633]), .Z(n7075) );
  AND U14151 ( .A(n7076), .B(p_input[3632]), .Z(o[3632]) );
  AND U14152 ( .A(p_input[23632]), .B(p_input[13632]), .Z(n7076) );
  AND U14153 ( .A(n7077), .B(p_input[3631]), .Z(o[3631]) );
  AND U14154 ( .A(p_input[23631]), .B(p_input[13631]), .Z(n7077) );
  AND U14155 ( .A(n7078), .B(p_input[3630]), .Z(o[3630]) );
  AND U14156 ( .A(p_input[23630]), .B(p_input[13630]), .Z(n7078) );
  AND U14157 ( .A(n7079), .B(p_input[362]), .Z(o[362]) );
  AND U14158 ( .A(p_input[20362]), .B(p_input[10362]), .Z(n7079) );
  AND U14159 ( .A(n7080), .B(p_input[3629]), .Z(o[3629]) );
  AND U14160 ( .A(p_input[23629]), .B(p_input[13629]), .Z(n7080) );
  AND U14161 ( .A(n7081), .B(p_input[3628]), .Z(o[3628]) );
  AND U14162 ( .A(p_input[23628]), .B(p_input[13628]), .Z(n7081) );
  AND U14163 ( .A(n7082), .B(p_input[3627]), .Z(o[3627]) );
  AND U14164 ( .A(p_input[23627]), .B(p_input[13627]), .Z(n7082) );
  AND U14165 ( .A(n7083), .B(p_input[3626]), .Z(o[3626]) );
  AND U14166 ( .A(p_input[23626]), .B(p_input[13626]), .Z(n7083) );
  AND U14167 ( .A(n7084), .B(p_input[3625]), .Z(o[3625]) );
  AND U14168 ( .A(p_input[23625]), .B(p_input[13625]), .Z(n7084) );
  AND U14169 ( .A(n7085), .B(p_input[3624]), .Z(o[3624]) );
  AND U14170 ( .A(p_input[23624]), .B(p_input[13624]), .Z(n7085) );
  AND U14171 ( .A(n7086), .B(p_input[3623]), .Z(o[3623]) );
  AND U14172 ( .A(p_input[23623]), .B(p_input[13623]), .Z(n7086) );
  AND U14173 ( .A(n7087), .B(p_input[3622]), .Z(o[3622]) );
  AND U14174 ( .A(p_input[23622]), .B(p_input[13622]), .Z(n7087) );
  AND U14175 ( .A(n7088), .B(p_input[3621]), .Z(o[3621]) );
  AND U14176 ( .A(p_input[23621]), .B(p_input[13621]), .Z(n7088) );
  AND U14177 ( .A(n7089), .B(p_input[3620]), .Z(o[3620]) );
  AND U14178 ( .A(p_input[23620]), .B(p_input[13620]), .Z(n7089) );
  AND U14179 ( .A(n7090), .B(p_input[361]), .Z(o[361]) );
  AND U14180 ( .A(p_input[20361]), .B(p_input[10361]), .Z(n7090) );
  AND U14181 ( .A(n7091), .B(p_input[3619]), .Z(o[3619]) );
  AND U14182 ( .A(p_input[23619]), .B(p_input[13619]), .Z(n7091) );
  AND U14183 ( .A(n7092), .B(p_input[3618]), .Z(o[3618]) );
  AND U14184 ( .A(p_input[23618]), .B(p_input[13618]), .Z(n7092) );
  AND U14185 ( .A(n7093), .B(p_input[3617]), .Z(o[3617]) );
  AND U14186 ( .A(p_input[23617]), .B(p_input[13617]), .Z(n7093) );
  AND U14187 ( .A(n7094), .B(p_input[3616]), .Z(o[3616]) );
  AND U14188 ( .A(p_input[23616]), .B(p_input[13616]), .Z(n7094) );
  AND U14189 ( .A(n7095), .B(p_input[3615]), .Z(o[3615]) );
  AND U14190 ( .A(p_input[23615]), .B(p_input[13615]), .Z(n7095) );
  AND U14191 ( .A(n7096), .B(p_input[3614]), .Z(o[3614]) );
  AND U14192 ( .A(p_input[23614]), .B(p_input[13614]), .Z(n7096) );
  AND U14193 ( .A(n7097), .B(p_input[3613]), .Z(o[3613]) );
  AND U14194 ( .A(p_input[23613]), .B(p_input[13613]), .Z(n7097) );
  AND U14195 ( .A(n7098), .B(p_input[3612]), .Z(o[3612]) );
  AND U14196 ( .A(p_input[23612]), .B(p_input[13612]), .Z(n7098) );
  AND U14197 ( .A(n7099), .B(p_input[3611]), .Z(o[3611]) );
  AND U14198 ( .A(p_input[23611]), .B(p_input[13611]), .Z(n7099) );
  AND U14199 ( .A(n7100), .B(p_input[3610]), .Z(o[3610]) );
  AND U14200 ( .A(p_input[23610]), .B(p_input[13610]), .Z(n7100) );
  AND U14201 ( .A(n7101), .B(p_input[360]), .Z(o[360]) );
  AND U14202 ( .A(p_input[20360]), .B(p_input[10360]), .Z(n7101) );
  AND U14203 ( .A(n7102), .B(p_input[3609]), .Z(o[3609]) );
  AND U14204 ( .A(p_input[23609]), .B(p_input[13609]), .Z(n7102) );
  AND U14205 ( .A(n7103), .B(p_input[3608]), .Z(o[3608]) );
  AND U14206 ( .A(p_input[23608]), .B(p_input[13608]), .Z(n7103) );
  AND U14207 ( .A(n7104), .B(p_input[3607]), .Z(o[3607]) );
  AND U14208 ( .A(p_input[23607]), .B(p_input[13607]), .Z(n7104) );
  AND U14209 ( .A(n7105), .B(p_input[3606]), .Z(o[3606]) );
  AND U14210 ( .A(p_input[23606]), .B(p_input[13606]), .Z(n7105) );
  AND U14211 ( .A(n7106), .B(p_input[3605]), .Z(o[3605]) );
  AND U14212 ( .A(p_input[23605]), .B(p_input[13605]), .Z(n7106) );
  AND U14213 ( .A(n7107), .B(p_input[3604]), .Z(o[3604]) );
  AND U14214 ( .A(p_input[23604]), .B(p_input[13604]), .Z(n7107) );
  AND U14215 ( .A(n7108), .B(p_input[3603]), .Z(o[3603]) );
  AND U14216 ( .A(p_input[23603]), .B(p_input[13603]), .Z(n7108) );
  AND U14217 ( .A(n7109), .B(p_input[3602]), .Z(o[3602]) );
  AND U14218 ( .A(p_input[23602]), .B(p_input[13602]), .Z(n7109) );
  AND U14219 ( .A(n7110), .B(p_input[3601]), .Z(o[3601]) );
  AND U14220 ( .A(p_input[23601]), .B(p_input[13601]), .Z(n7110) );
  AND U14221 ( .A(n7111), .B(p_input[3600]), .Z(o[3600]) );
  AND U14222 ( .A(p_input[23600]), .B(p_input[13600]), .Z(n7111) );
  AND U14223 ( .A(n7112), .B(p_input[35]), .Z(o[35]) );
  AND U14224 ( .A(p_input[20035]), .B(p_input[10035]), .Z(n7112) );
  AND U14225 ( .A(n7113), .B(p_input[359]), .Z(o[359]) );
  AND U14226 ( .A(p_input[20359]), .B(p_input[10359]), .Z(n7113) );
  AND U14227 ( .A(n7114), .B(p_input[3599]), .Z(o[3599]) );
  AND U14228 ( .A(p_input[23599]), .B(p_input[13599]), .Z(n7114) );
  AND U14229 ( .A(n7115), .B(p_input[3598]), .Z(o[3598]) );
  AND U14230 ( .A(p_input[23598]), .B(p_input[13598]), .Z(n7115) );
  AND U14231 ( .A(n7116), .B(p_input[3597]), .Z(o[3597]) );
  AND U14232 ( .A(p_input[23597]), .B(p_input[13597]), .Z(n7116) );
  AND U14233 ( .A(n7117), .B(p_input[3596]), .Z(o[3596]) );
  AND U14234 ( .A(p_input[23596]), .B(p_input[13596]), .Z(n7117) );
  AND U14235 ( .A(n7118), .B(p_input[3595]), .Z(o[3595]) );
  AND U14236 ( .A(p_input[23595]), .B(p_input[13595]), .Z(n7118) );
  AND U14237 ( .A(n7119), .B(p_input[3594]), .Z(o[3594]) );
  AND U14238 ( .A(p_input[23594]), .B(p_input[13594]), .Z(n7119) );
  AND U14239 ( .A(n7120), .B(p_input[3593]), .Z(o[3593]) );
  AND U14240 ( .A(p_input[23593]), .B(p_input[13593]), .Z(n7120) );
  AND U14241 ( .A(n7121), .B(p_input[3592]), .Z(o[3592]) );
  AND U14242 ( .A(p_input[23592]), .B(p_input[13592]), .Z(n7121) );
  AND U14243 ( .A(n7122), .B(p_input[3591]), .Z(o[3591]) );
  AND U14244 ( .A(p_input[23591]), .B(p_input[13591]), .Z(n7122) );
  AND U14245 ( .A(n7123), .B(p_input[3590]), .Z(o[3590]) );
  AND U14246 ( .A(p_input[23590]), .B(p_input[13590]), .Z(n7123) );
  AND U14247 ( .A(n7124), .B(p_input[358]), .Z(o[358]) );
  AND U14248 ( .A(p_input[20358]), .B(p_input[10358]), .Z(n7124) );
  AND U14249 ( .A(n7125), .B(p_input[3589]), .Z(o[3589]) );
  AND U14250 ( .A(p_input[23589]), .B(p_input[13589]), .Z(n7125) );
  AND U14251 ( .A(n7126), .B(p_input[3588]), .Z(o[3588]) );
  AND U14252 ( .A(p_input[23588]), .B(p_input[13588]), .Z(n7126) );
  AND U14253 ( .A(n7127), .B(p_input[3587]), .Z(o[3587]) );
  AND U14254 ( .A(p_input[23587]), .B(p_input[13587]), .Z(n7127) );
  AND U14255 ( .A(n7128), .B(p_input[3586]), .Z(o[3586]) );
  AND U14256 ( .A(p_input[23586]), .B(p_input[13586]), .Z(n7128) );
  AND U14257 ( .A(n7129), .B(p_input[3585]), .Z(o[3585]) );
  AND U14258 ( .A(p_input[23585]), .B(p_input[13585]), .Z(n7129) );
  AND U14259 ( .A(n7130), .B(p_input[3584]), .Z(o[3584]) );
  AND U14260 ( .A(p_input[23584]), .B(p_input[13584]), .Z(n7130) );
  AND U14261 ( .A(n7131), .B(p_input[3583]), .Z(o[3583]) );
  AND U14262 ( .A(p_input[23583]), .B(p_input[13583]), .Z(n7131) );
  AND U14263 ( .A(n7132), .B(p_input[3582]), .Z(o[3582]) );
  AND U14264 ( .A(p_input[23582]), .B(p_input[13582]), .Z(n7132) );
  AND U14265 ( .A(n7133), .B(p_input[3581]), .Z(o[3581]) );
  AND U14266 ( .A(p_input[23581]), .B(p_input[13581]), .Z(n7133) );
  AND U14267 ( .A(n7134), .B(p_input[3580]), .Z(o[3580]) );
  AND U14268 ( .A(p_input[23580]), .B(p_input[13580]), .Z(n7134) );
  AND U14269 ( .A(n7135), .B(p_input[357]), .Z(o[357]) );
  AND U14270 ( .A(p_input[20357]), .B(p_input[10357]), .Z(n7135) );
  AND U14271 ( .A(n7136), .B(p_input[3579]), .Z(o[3579]) );
  AND U14272 ( .A(p_input[23579]), .B(p_input[13579]), .Z(n7136) );
  AND U14273 ( .A(n7137), .B(p_input[3578]), .Z(o[3578]) );
  AND U14274 ( .A(p_input[23578]), .B(p_input[13578]), .Z(n7137) );
  AND U14275 ( .A(n7138), .B(p_input[3577]), .Z(o[3577]) );
  AND U14276 ( .A(p_input[23577]), .B(p_input[13577]), .Z(n7138) );
  AND U14277 ( .A(n7139), .B(p_input[3576]), .Z(o[3576]) );
  AND U14278 ( .A(p_input[23576]), .B(p_input[13576]), .Z(n7139) );
  AND U14279 ( .A(n7140), .B(p_input[3575]), .Z(o[3575]) );
  AND U14280 ( .A(p_input[23575]), .B(p_input[13575]), .Z(n7140) );
  AND U14281 ( .A(n7141), .B(p_input[3574]), .Z(o[3574]) );
  AND U14282 ( .A(p_input[23574]), .B(p_input[13574]), .Z(n7141) );
  AND U14283 ( .A(n7142), .B(p_input[3573]), .Z(o[3573]) );
  AND U14284 ( .A(p_input[23573]), .B(p_input[13573]), .Z(n7142) );
  AND U14285 ( .A(n7143), .B(p_input[3572]), .Z(o[3572]) );
  AND U14286 ( .A(p_input[23572]), .B(p_input[13572]), .Z(n7143) );
  AND U14287 ( .A(n7144), .B(p_input[3571]), .Z(o[3571]) );
  AND U14288 ( .A(p_input[23571]), .B(p_input[13571]), .Z(n7144) );
  AND U14289 ( .A(n7145), .B(p_input[3570]), .Z(o[3570]) );
  AND U14290 ( .A(p_input[23570]), .B(p_input[13570]), .Z(n7145) );
  AND U14291 ( .A(n7146), .B(p_input[356]), .Z(o[356]) );
  AND U14292 ( .A(p_input[20356]), .B(p_input[10356]), .Z(n7146) );
  AND U14293 ( .A(n7147), .B(p_input[3569]), .Z(o[3569]) );
  AND U14294 ( .A(p_input[23569]), .B(p_input[13569]), .Z(n7147) );
  AND U14295 ( .A(n7148), .B(p_input[3568]), .Z(o[3568]) );
  AND U14296 ( .A(p_input[23568]), .B(p_input[13568]), .Z(n7148) );
  AND U14297 ( .A(n7149), .B(p_input[3567]), .Z(o[3567]) );
  AND U14298 ( .A(p_input[23567]), .B(p_input[13567]), .Z(n7149) );
  AND U14299 ( .A(n7150), .B(p_input[3566]), .Z(o[3566]) );
  AND U14300 ( .A(p_input[23566]), .B(p_input[13566]), .Z(n7150) );
  AND U14301 ( .A(n7151), .B(p_input[3565]), .Z(o[3565]) );
  AND U14302 ( .A(p_input[23565]), .B(p_input[13565]), .Z(n7151) );
  AND U14303 ( .A(n7152), .B(p_input[3564]), .Z(o[3564]) );
  AND U14304 ( .A(p_input[23564]), .B(p_input[13564]), .Z(n7152) );
  AND U14305 ( .A(n7153), .B(p_input[3563]), .Z(o[3563]) );
  AND U14306 ( .A(p_input[23563]), .B(p_input[13563]), .Z(n7153) );
  AND U14307 ( .A(n7154), .B(p_input[3562]), .Z(o[3562]) );
  AND U14308 ( .A(p_input[23562]), .B(p_input[13562]), .Z(n7154) );
  AND U14309 ( .A(n7155), .B(p_input[3561]), .Z(o[3561]) );
  AND U14310 ( .A(p_input[23561]), .B(p_input[13561]), .Z(n7155) );
  AND U14311 ( .A(n7156), .B(p_input[3560]), .Z(o[3560]) );
  AND U14312 ( .A(p_input[23560]), .B(p_input[13560]), .Z(n7156) );
  AND U14313 ( .A(n7157), .B(p_input[355]), .Z(o[355]) );
  AND U14314 ( .A(p_input[20355]), .B(p_input[10355]), .Z(n7157) );
  AND U14315 ( .A(n7158), .B(p_input[3559]), .Z(o[3559]) );
  AND U14316 ( .A(p_input[23559]), .B(p_input[13559]), .Z(n7158) );
  AND U14317 ( .A(n7159), .B(p_input[3558]), .Z(o[3558]) );
  AND U14318 ( .A(p_input[23558]), .B(p_input[13558]), .Z(n7159) );
  AND U14319 ( .A(n7160), .B(p_input[3557]), .Z(o[3557]) );
  AND U14320 ( .A(p_input[23557]), .B(p_input[13557]), .Z(n7160) );
  AND U14321 ( .A(n7161), .B(p_input[3556]), .Z(o[3556]) );
  AND U14322 ( .A(p_input[23556]), .B(p_input[13556]), .Z(n7161) );
  AND U14323 ( .A(n7162), .B(p_input[3555]), .Z(o[3555]) );
  AND U14324 ( .A(p_input[23555]), .B(p_input[13555]), .Z(n7162) );
  AND U14325 ( .A(n7163), .B(p_input[3554]), .Z(o[3554]) );
  AND U14326 ( .A(p_input[23554]), .B(p_input[13554]), .Z(n7163) );
  AND U14327 ( .A(n7164), .B(p_input[3553]), .Z(o[3553]) );
  AND U14328 ( .A(p_input[23553]), .B(p_input[13553]), .Z(n7164) );
  AND U14329 ( .A(n7165), .B(p_input[3552]), .Z(o[3552]) );
  AND U14330 ( .A(p_input[23552]), .B(p_input[13552]), .Z(n7165) );
  AND U14331 ( .A(n7166), .B(p_input[3551]), .Z(o[3551]) );
  AND U14332 ( .A(p_input[23551]), .B(p_input[13551]), .Z(n7166) );
  AND U14333 ( .A(n7167), .B(p_input[3550]), .Z(o[3550]) );
  AND U14334 ( .A(p_input[23550]), .B(p_input[13550]), .Z(n7167) );
  AND U14335 ( .A(n7168), .B(p_input[354]), .Z(o[354]) );
  AND U14336 ( .A(p_input[20354]), .B(p_input[10354]), .Z(n7168) );
  AND U14337 ( .A(n7169), .B(p_input[3549]), .Z(o[3549]) );
  AND U14338 ( .A(p_input[23549]), .B(p_input[13549]), .Z(n7169) );
  AND U14339 ( .A(n7170), .B(p_input[3548]), .Z(o[3548]) );
  AND U14340 ( .A(p_input[23548]), .B(p_input[13548]), .Z(n7170) );
  AND U14341 ( .A(n7171), .B(p_input[3547]), .Z(o[3547]) );
  AND U14342 ( .A(p_input[23547]), .B(p_input[13547]), .Z(n7171) );
  AND U14343 ( .A(n7172), .B(p_input[3546]), .Z(o[3546]) );
  AND U14344 ( .A(p_input[23546]), .B(p_input[13546]), .Z(n7172) );
  AND U14345 ( .A(n7173), .B(p_input[3545]), .Z(o[3545]) );
  AND U14346 ( .A(p_input[23545]), .B(p_input[13545]), .Z(n7173) );
  AND U14347 ( .A(n7174), .B(p_input[3544]), .Z(o[3544]) );
  AND U14348 ( .A(p_input[23544]), .B(p_input[13544]), .Z(n7174) );
  AND U14349 ( .A(n7175), .B(p_input[3543]), .Z(o[3543]) );
  AND U14350 ( .A(p_input[23543]), .B(p_input[13543]), .Z(n7175) );
  AND U14351 ( .A(n7176), .B(p_input[3542]), .Z(o[3542]) );
  AND U14352 ( .A(p_input[23542]), .B(p_input[13542]), .Z(n7176) );
  AND U14353 ( .A(n7177), .B(p_input[3541]), .Z(o[3541]) );
  AND U14354 ( .A(p_input[23541]), .B(p_input[13541]), .Z(n7177) );
  AND U14355 ( .A(n7178), .B(p_input[3540]), .Z(o[3540]) );
  AND U14356 ( .A(p_input[23540]), .B(p_input[13540]), .Z(n7178) );
  AND U14357 ( .A(n7179), .B(p_input[353]), .Z(o[353]) );
  AND U14358 ( .A(p_input[20353]), .B(p_input[10353]), .Z(n7179) );
  AND U14359 ( .A(n7180), .B(p_input[3539]), .Z(o[3539]) );
  AND U14360 ( .A(p_input[23539]), .B(p_input[13539]), .Z(n7180) );
  AND U14361 ( .A(n7181), .B(p_input[3538]), .Z(o[3538]) );
  AND U14362 ( .A(p_input[23538]), .B(p_input[13538]), .Z(n7181) );
  AND U14363 ( .A(n7182), .B(p_input[3537]), .Z(o[3537]) );
  AND U14364 ( .A(p_input[23537]), .B(p_input[13537]), .Z(n7182) );
  AND U14365 ( .A(n7183), .B(p_input[3536]), .Z(o[3536]) );
  AND U14366 ( .A(p_input[23536]), .B(p_input[13536]), .Z(n7183) );
  AND U14367 ( .A(n7184), .B(p_input[3535]), .Z(o[3535]) );
  AND U14368 ( .A(p_input[23535]), .B(p_input[13535]), .Z(n7184) );
  AND U14369 ( .A(n7185), .B(p_input[3534]), .Z(o[3534]) );
  AND U14370 ( .A(p_input[23534]), .B(p_input[13534]), .Z(n7185) );
  AND U14371 ( .A(n7186), .B(p_input[3533]), .Z(o[3533]) );
  AND U14372 ( .A(p_input[23533]), .B(p_input[13533]), .Z(n7186) );
  AND U14373 ( .A(n7187), .B(p_input[3532]), .Z(o[3532]) );
  AND U14374 ( .A(p_input[23532]), .B(p_input[13532]), .Z(n7187) );
  AND U14375 ( .A(n7188), .B(p_input[3531]), .Z(o[3531]) );
  AND U14376 ( .A(p_input[23531]), .B(p_input[13531]), .Z(n7188) );
  AND U14377 ( .A(n7189), .B(p_input[3530]), .Z(o[3530]) );
  AND U14378 ( .A(p_input[23530]), .B(p_input[13530]), .Z(n7189) );
  AND U14379 ( .A(n7190), .B(p_input[352]), .Z(o[352]) );
  AND U14380 ( .A(p_input[20352]), .B(p_input[10352]), .Z(n7190) );
  AND U14381 ( .A(n7191), .B(p_input[3529]), .Z(o[3529]) );
  AND U14382 ( .A(p_input[23529]), .B(p_input[13529]), .Z(n7191) );
  AND U14383 ( .A(n7192), .B(p_input[3528]), .Z(o[3528]) );
  AND U14384 ( .A(p_input[23528]), .B(p_input[13528]), .Z(n7192) );
  AND U14385 ( .A(n7193), .B(p_input[3527]), .Z(o[3527]) );
  AND U14386 ( .A(p_input[23527]), .B(p_input[13527]), .Z(n7193) );
  AND U14387 ( .A(n7194), .B(p_input[3526]), .Z(o[3526]) );
  AND U14388 ( .A(p_input[23526]), .B(p_input[13526]), .Z(n7194) );
  AND U14389 ( .A(n7195), .B(p_input[3525]), .Z(o[3525]) );
  AND U14390 ( .A(p_input[23525]), .B(p_input[13525]), .Z(n7195) );
  AND U14391 ( .A(n7196), .B(p_input[3524]), .Z(o[3524]) );
  AND U14392 ( .A(p_input[23524]), .B(p_input[13524]), .Z(n7196) );
  AND U14393 ( .A(n7197), .B(p_input[3523]), .Z(o[3523]) );
  AND U14394 ( .A(p_input[23523]), .B(p_input[13523]), .Z(n7197) );
  AND U14395 ( .A(n7198), .B(p_input[3522]), .Z(o[3522]) );
  AND U14396 ( .A(p_input[23522]), .B(p_input[13522]), .Z(n7198) );
  AND U14397 ( .A(n7199), .B(p_input[3521]), .Z(o[3521]) );
  AND U14398 ( .A(p_input[23521]), .B(p_input[13521]), .Z(n7199) );
  AND U14399 ( .A(n7200), .B(p_input[3520]), .Z(o[3520]) );
  AND U14400 ( .A(p_input[23520]), .B(p_input[13520]), .Z(n7200) );
  AND U14401 ( .A(n7201), .B(p_input[351]), .Z(o[351]) );
  AND U14402 ( .A(p_input[20351]), .B(p_input[10351]), .Z(n7201) );
  AND U14403 ( .A(n7202), .B(p_input[3519]), .Z(o[3519]) );
  AND U14404 ( .A(p_input[23519]), .B(p_input[13519]), .Z(n7202) );
  AND U14405 ( .A(n7203), .B(p_input[3518]), .Z(o[3518]) );
  AND U14406 ( .A(p_input[23518]), .B(p_input[13518]), .Z(n7203) );
  AND U14407 ( .A(n7204), .B(p_input[3517]), .Z(o[3517]) );
  AND U14408 ( .A(p_input[23517]), .B(p_input[13517]), .Z(n7204) );
  AND U14409 ( .A(n7205), .B(p_input[3516]), .Z(o[3516]) );
  AND U14410 ( .A(p_input[23516]), .B(p_input[13516]), .Z(n7205) );
  AND U14411 ( .A(n7206), .B(p_input[3515]), .Z(o[3515]) );
  AND U14412 ( .A(p_input[23515]), .B(p_input[13515]), .Z(n7206) );
  AND U14413 ( .A(n7207), .B(p_input[3514]), .Z(o[3514]) );
  AND U14414 ( .A(p_input[23514]), .B(p_input[13514]), .Z(n7207) );
  AND U14415 ( .A(n7208), .B(p_input[3513]), .Z(o[3513]) );
  AND U14416 ( .A(p_input[23513]), .B(p_input[13513]), .Z(n7208) );
  AND U14417 ( .A(n7209), .B(p_input[3512]), .Z(o[3512]) );
  AND U14418 ( .A(p_input[23512]), .B(p_input[13512]), .Z(n7209) );
  AND U14419 ( .A(n7210), .B(p_input[3511]), .Z(o[3511]) );
  AND U14420 ( .A(p_input[23511]), .B(p_input[13511]), .Z(n7210) );
  AND U14421 ( .A(n7211), .B(p_input[3510]), .Z(o[3510]) );
  AND U14422 ( .A(p_input[23510]), .B(p_input[13510]), .Z(n7211) );
  AND U14423 ( .A(n7212), .B(p_input[350]), .Z(o[350]) );
  AND U14424 ( .A(p_input[20350]), .B(p_input[10350]), .Z(n7212) );
  AND U14425 ( .A(n7213), .B(p_input[3509]), .Z(o[3509]) );
  AND U14426 ( .A(p_input[23509]), .B(p_input[13509]), .Z(n7213) );
  AND U14427 ( .A(n7214), .B(p_input[3508]), .Z(o[3508]) );
  AND U14428 ( .A(p_input[23508]), .B(p_input[13508]), .Z(n7214) );
  AND U14429 ( .A(n7215), .B(p_input[3507]), .Z(o[3507]) );
  AND U14430 ( .A(p_input[23507]), .B(p_input[13507]), .Z(n7215) );
  AND U14431 ( .A(n7216), .B(p_input[3506]), .Z(o[3506]) );
  AND U14432 ( .A(p_input[23506]), .B(p_input[13506]), .Z(n7216) );
  AND U14433 ( .A(n7217), .B(p_input[3505]), .Z(o[3505]) );
  AND U14434 ( .A(p_input[23505]), .B(p_input[13505]), .Z(n7217) );
  AND U14435 ( .A(n7218), .B(p_input[3504]), .Z(o[3504]) );
  AND U14436 ( .A(p_input[23504]), .B(p_input[13504]), .Z(n7218) );
  AND U14437 ( .A(n7219), .B(p_input[3503]), .Z(o[3503]) );
  AND U14438 ( .A(p_input[23503]), .B(p_input[13503]), .Z(n7219) );
  AND U14439 ( .A(n7220), .B(p_input[3502]), .Z(o[3502]) );
  AND U14440 ( .A(p_input[23502]), .B(p_input[13502]), .Z(n7220) );
  AND U14441 ( .A(n7221), .B(p_input[3501]), .Z(o[3501]) );
  AND U14442 ( .A(p_input[23501]), .B(p_input[13501]), .Z(n7221) );
  AND U14443 ( .A(n7222), .B(p_input[3500]), .Z(o[3500]) );
  AND U14444 ( .A(p_input[23500]), .B(p_input[13500]), .Z(n7222) );
  AND U14445 ( .A(n7223), .B(p_input[34]), .Z(o[34]) );
  AND U14446 ( .A(p_input[20034]), .B(p_input[10034]), .Z(n7223) );
  AND U14447 ( .A(n7224), .B(p_input[349]), .Z(o[349]) );
  AND U14448 ( .A(p_input[20349]), .B(p_input[10349]), .Z(n7224) );
  AND U14449 ( .A(n7225), .B(p_input[3499]), .Z(o[3499]) );
  AND U14450 ( .A(p_input[23499]), .B(p_input[13499]), .Z(n7225) );
  AND U14451 ( .A(n7226), .B(p_input[3498]), .Z(o[3498]) );
  AND U14452 ( .A(p_input[23498]), .B(p_input[13498]), .Z(n7226) );
  AND U14453 ( .A(n7227), .B(p_input[3497]), .Z(o[3497]) );
  AND U14454 ( .A(p_input[23497]), .B(p_input[13497]), .Z(n7227) );
  AND U14455 ( .A(n7228), .B(p_input[3496]), .Z(o[3496]) );
  AND U14456 ( .A(p_input[23496]), .B(p_input[13496]), .Z(n7228) );
  AND U14457 ( .A(n7229), .B(p_input[3495]), .Z(o[3495]) );
  AND U14458 ( .A(p_input[23495]), .B(p_input[13495]), .Z(n7229) );
  AND U14459 ( .A(n7230), .B(p_input[3494]), .Z(o[3494]) );
  AND U14460 ( .A(p_input[23494]), .B(p_input[13494]), .Z(n7230) );
  AND U14461 ( .A(n7231), .B(p_input[3493]), .Z(o[3493]) );
  AND U14462 ( .A(p_input[23493]), .B(p_input[13493]), .Z(n7231) );
  AND U14463 ( .A(n7232), .B(p_input[3492]), .Z(o[3492]) );
  AND U14464 ( .A(p_input[23492]), .B(p_input[13492]), .Z(n7232) );
  AND U14465 ( .A(n7233), .B(p_input[3491]), .Z(o[3491]) );
  AND U14466 ( .A(p_input[23491]), .B(p_input[13491]), .Z(n7233) );
  AND U14467 ( .A(n7234), .B(p_input[3490]), .Z(o[3490]) );
  AND U14468 ( .A(p_input[23490]), .B(p_input[13490]), .Z(n7234) );
  AND U14469 ( .A(n7235), .B(p_input[348]), .Z(o[348]) );
  AND U14470 ( .A(p_input[20348]), .B(p_input[10348]), .Z(n7235) );
  AND U14471 ( .A(n7236), .B(p_input[3489]), .Z(o[3489]) );
  AND U14472 ( .A(p_input[23489]), .B(p_input[13489]), .Z(n7236) );
  AND U14473 ( .A(n7237), .B(p_input[3488]), .Z(o[3488]) );
  AND U14474 ( .A(p_input[23488]), .B(p_input[13488]), .Z(n7237) );
  AND U14475 ( .A(n7238), .B(p_input[3487]), .Z(o[3487]) );
  AND U14476 ( .A(p_input[23487]), .B(p_input[13487]), .Z(n7238) );
  AND U14477 ( .A(n7239), .B(p_input[3486]), .Z(o[3486]) );
  AND U14478 ( .A(p_input[23486]), .B(p_input[13486]), .Z(n7239) );
  AND U14479 ( .A(n7240), .B(p_input[3485]), .Z(o[3485]) );
  AND U14480 ( .A(p_input[23485]), .B(p_input[13485]), .Z(n7240) );
  AND U14481 ( .A(n7241), .B(p_input[3484]), .Z(o[3484]) );
  AND U14482 ( .A(p_input[23484]), .B(p_input[13484]), .Z(n7241) );
  AND U14483 ( .A(n7242), .B(p_input[3483]), .Z(o[3483]) );
  AND U14484 ( .A(p_input[23483]), .B(p_input[13483]), .Z(n7242) );
  AND U14485 ( .A(n7243), .B(p_input[3482]), .Z(o[3482]) );
  AND U14486 ( .A(p_input[23482]), .B(p_input[13482]), .Z(n7243) );
  AND U14487 ( .A(n7244), .B(p_input[3481]), .Z(o[3481]) );
  AND U14488 ( .A(p_input[23481]), .B(p_input[13481]), .Z(n7244) );
  AND U14489 ( .A(n7245), .B(p_input[3480]), .Z(o[3480]) );
  AND U14490 ( .A(p_input[23480]), .B(p_input[13480]), .Z(n7245) );
  AND U14491 ( .A(n7246), .B(p_input[347]), .Z(o[347]) );
  AND U14492 ( .A(p_input[20347]), .B(p_input[10347]), .Z(n7246) );
  AND U14493 ( .A(n7247), .B(p_input[3479]), .Z(o[3479]) );
  AND U14494 ( .A(p_input[23479]), .B(p_input[13479]), .Z(n7247) );
  AND U14495 ( .A(n7248), .B(p_input[3478]), .Z(o[3478]) );
  AND U14496 ( .A(p_input[23478]), .B(p_input[13478]), .Z(n7248) );
  AND U14497 ( .A(n7249), .B(p_input[3477]), .Z(o[3477]) );
  AND U14498 ( .A(p_input[23477]), .B(p_input[13477]), .Z(n7249) );
  AND U14499 ( .A(n7250), .B(p_input[3476]), .Z(o[3476]) );
  AND U14500 ( .A(p_input[23476]), .B(p_input[13476]), .Z(n7250) );
  AND U14501 ( .A(n7251), .B(p_input[3475]), .Z(o[3475]) );
  AND U14502 ( .A(p_input[23475]), .B(p_input[13475]), .Z(n7251) );
  AND U14503 ( .A(n7252), .B(p_input[3474]), .Z(o[3474]) );
  AND U14504 ( .A(p_input[23474]), .B(p_input[13474]), .Z(n7252) );
  AND U14505 ( .A(n7253), .B(p_input[3473]), .Z(o[3473]) );
  AND U14506 ( .A(p_input[23473]), .B(p_input[13473]), .Z(n7253) );
  AND U14507 ( .A(n7254), .B(p_input[3472]), .Z(o[3472]) );
  AND U14508 ( .A(p_input[23472]), .B(p_input[13472]), .Z(n7254) );
  AND U14509 ( .A(n7255), .B(p_input[3471]), .Z(o[3471]) );
  AND U14510 ( .A(p_input[23471]), .B(p_input[13471]), .Z(n7255) );
  AND U14511 ( .A(n7256), .B(p_input[3470]), .Z(o[3470]) );
  AND U14512 ( .A(p_input[23470]), .B(p_input[13470]), .Z(n7256) );
  AND U14513 ( .A(n7257), .B(p_input[346]), .Z(o[346]) );
  AND U14514 ( .A(p_input[20346]), .B(p_input[10346]), .Z(n7257) );
  AND U14515 ( .A(n7258), .B(p_input[3469]), .Z(o[3469]) );
  AND U14516 ( .A(p_input[23469]), .B(p_input[13469]), .Z(n7258) );
  AND U14517 ( .A(n7259), .B(p_input[3468]), .Z(o[3468]) );
  AND U14518 ( .A(p_input[23468]), .B(p_input[13468]), .Z(n7259) );
  AND U14519 ( .A(n7260), .B(p_input[3467]), .Z(o[3467]) );
  AND U14520 ( .A(p_input[23467]), .B(p_input[13467]), .Z(n7260) );
  AND U14521 ( .A(n7261), .B(p_input[3466]), .Z(o[3466]) );
  AND U14522 ( .A(p_input[23466]), .B(p_input[13466]), .Z(n7261) );
  AND U14523 ( .A(n7262), .B(p_input[3465]), .Z(o[3465]) );
  AND U14524 ( .A(p_input[23465]), .B(p_input[13465]), .Z(n7262) );
  AND U14525 ( .A(n7263), .B(p_input[3464]), .Z(o[3464]) );
  AND U14526 ( .A(p_input[23464]), .B(p_input[13464]), .Z(n7263) );
  AND U14527 ( .A(n7264), .B(p_input[3463]), .Z(o[3463]) );
  AND U14528 ( .A(p_input[23463]), .B(p_input[13463]), .Z(n7264) );
  AND U14529 ( .A(n7265), .B(p_input[3462]), .Z(o[3462]) );
  AND U14530 ( .A(p_input[23462]), .B(p_input[13462]), .Z(n7265) );
  AND U14531 ( .A(n7266), .B(p_input[3461]), .Z(o[3461]) );
  AND U14532 ( .A(p_input[23461]), .B(p_input[13461]), .Z(n7266) );
  AND U14533 ( .A(n7267), .B(p_input[3460]), .Z(o[3460]) );
  AND U14534 ( .A(p_input[23460]), .B(p_input[13460]), .Z(n7267) );
  AND U14535 ( .A(n7268), .B(p_input[345]), .Z(o[345]) );
  AND U14536 ( .A(p_input[20345]), .B(p_input[10345]), .Z(n7268) );
  AND U14537 ( .A(n7269), .B(p_input[3459]), .Z(o[3459]) );
  AND U14538 ( .A(p_input[23459]), .B(p_input[13459]), .Z(n7269) );
  AND U14539 ( .A(n7270), .B(p_input[3458]), .Z(o[3458]) );
  AND U14540 ( .A(p_input[23458]), .B(p_input[13458]), .Z(n7270) );
  AND U14541 ( .A(n7271), .B(p_input[3457]), .Z(o[3457]) );
  AND U14542 ( .A(p_input[23457]), .B(p_input[13457]), .Z(n7271) );
  AND U14543 ( .A(n7272), .B(p_input[3456]), .Z(o[3456]) );
  AND U14544 ( .A(p_input[23456]), .B(p_input[13456]), .Z(n7272) );
  AND U14545 ( .A(n7273), .B(p_input[3455]), .Z(o[3455]) );
  AND U14546 ( .A(p_input[23455]), .B(p_input[13455]), .Z(n7273) );
  AND U14547 ( .A(n7274), .B(p_input[3454]), .Z(o[3454]) );
  AND U14548 ( .A(p_input[23454]), .B(p_input[13454]), .Z(n7274) );
  AND U14549 ( .A(n7275), .B(p_input[3453]), .Z(o[3453]) );
  AND U14550 ( .A(p_input[23453]), .B(p_input[13453]), .Z(n7275) );
  AND U14551 ( .A(n7276), .B(p_input[3452]), .Z(o[3452]) );
  AND U14552 ( .A(p_input[23452]), .B(p_input[13452]), .Z(n7276) );
  AND U14553 ( .A(n7277), .B(p_input[3451]), .Z(o[3451]) );
  AND U14554 ( .A(p_input[23451]), .B(p_input[13451]), .Z(n7277) );
  AND U14555 ( .A(n7278), .B(p_input[3450]), .Z(o[3450]) );
  AND U14556 ( .A(p_input[23450]), .B(p_input[13450]), .Z(n7278) );
  AND U14557 ( .A(n7279), .B(p_input[344]), .Z(o[344]) );
  AND U14558 ( .A(p_input[20344]), .B(p_input[10344]), .Z(n7279) );
  AND U14559 ( .A(n7280), .B(p_input[3449]), .Z(o[3449]) );
  AND U14560 ( .A(p_input[23449]), .B(p_input[13449]), .Z(n7280) );
  AND U14561 ( .A(n7281), .B(p_input[3448]), .Z(o[3448]) );
  AND U14562 ( .A(p_input[23448]), .B(p_input[13448]), .Z(n7281) );
  AND U14563 ( .A(n7282), .B(p_input[3447]), .Z(o[3447]) );
  AND U14564 ( .A(p_input[23447]), .B(p_input[13447]), .Z(n7282) );
  AND U14565 ( .A(n7283), .B(p_input[3446]), .Z(o[3446]) );
  AND U14566 ( .A(p_input[23446]), .B(p_input[13446]), .Z(n7283) );
  AND U14567 ( .A(n7284), .B(p_input[3445]), .Z(o[3445]) );
  AND U14568 ( .A(p_input[23445]), .B(p_input[13445]), .Z(n7284) );
  AND U14569 ( .A(n7285), .B(p_input[3444]), .Z(o[3444]) );
  AND U14570 ( .A(p_input[23444]), .B(p_input[13444]), .Z(n7285) );
  AND U14571 ( .A(n7286), .B(p_input[3443]), .Z(o[3443]) );
  AND U14572 ( .A(p_input[23443]), .B(p_input[13443]), .Z(n7286) );
  AND U14573 ( .A(n7287), .B(p_input[3442]), .Z(o[3442]) );
  AND U14574 ( .A(p_input[23442]), .B(p_input[13442]), .Z(n7287) );
  AND U14575 ( .A(n7288), .B(p_input[3441]), .Z(o[3441]) );
  AND U14576 ( .A(p_input[23441]), .B(p_input[13441]), .Z(n7288) );
  AND U14577 ( .A(n7289), .B(p_input[3440]), .Z(o[3440]) );
  AND U14578 ( .A(p_input[23440]), .B(p_input[13440]), .Z(n7289) );
  AND U14579 ( .A(n7290), .B(p_input[343]), .Z(o[343]) );
  AND U14580 ( .A(p_input[20343]), .B(p_input[10343]), .Z(n7290) );
  AND U14581 ( .A(n7291), .B(p_input[3439]), .Z(o[3439]) );
  AND U14582 ( .A(p_input[23439]), .B(p_input[13439]), .Z(n7291) );
  AND U14583 ( .A(n7292), .B(p_input[3438]), .Z(o[3438]) );
  AND U14584 ( .A(p_input[23438]), .B(p_input[13438]), .Z(n7292) );
  AND U14585 ( .A(n7293), .B(p_input[3437]), .Z(o[3437]) );
  AND U14586 ( .A(p_input[23437]), .B(p_input[13437]), .Z(n7293) );
  AND U14587 ( .A(n7294), .B(p_input[3436]), .Z(o[3436]) );
  AND U14588 ( .A(p_input[23436]), .B(p_input[13436]), .Z(n7294) );
  AND U14589 ( .A(n7295), .B(p_input[3435]), .Z(o[3435]) );
  AND U14590 ( .A(p_input[23435]), .B(p_input[13435]), .Z(n7295) );
  AND U14591 ( .A(n7296), .B(p_input[3434]), .Z(o[3434]) );
  AND U14592 ( .A(p_input[23434]), .B(p_input[13434]), .Z(n7296) );
  AND U14593 ( .A(n7297), .B(p_input[3433]), .Z(o[3433]) );
  AND U14594 ( .A(p_input[23433]), .B(p_input[13433]), .Z(n7297) );
  AND U14595 ( .A(n7298), .B(p_input[3432]), .Z(o[3432]) );
  AND U14596 ( .A(p_input[23432]), .B(p_input[13432]), .Z(n7298) );
  AND U14597 ( .A(n7299), .B(p_input[3431]), .Z(o[3431]) );
  AND U14598 ( .A(p_input[23431]), .B(p_input[13431]), .Z(n7299) );
  AND U14599 ( .A(n7300), .B(p_input[3430]), .Z(o[3430]) );
  AND U14600 ( .A(p_input[23430]), .B(p_input[13430]), .Z(n7300) );
  AND U14601 ( .A(n7301), .B(p_input[342]), .Z(o[342]) );
  AND U14602 ( .A(p_input[20342]), .B(p_input[10342]), .Z(n7301) );
  AND U14603 ( .A(n7302), .B(p_input[3429]), .Z(o[3429]) );
  AND U14604 ( .A(p_input[23429]), .B(p_input[13429]), .Z(n7302) );
  AND U14605 ( .A(n7303), .B(p_input[3428]), .Z(o[3428]) );
  AND U14606 ( .A(p_input[23428]), .B(p_input[13428]), .Z(n7303) );
  AND U14607 ( .A(n7304), .B(p_input[3427]), .Z(o[3427]) );
  AND U14608 ( .A(p_input[23427]), .B(p_input[13427]), .Z(n7304) );
  AND U14609 ( .A(n7305), .B(p_input[3426]), .Z(o[3426]) );
  AND U14610 ( .A(p_input[23426]), .B(p_input[13426]), .Z(n7305) );
  AND U14611 ( .A(n7306), .B(p_input[3425]), .Z(o[3425]) );
  AND U14612 ( .A(p_input[23425]), .B(p_input[13425]), .Z(n7306) );
  AND U14613 ( .A(n7307), .B(p_input[3424]), .Z(o[3424]) );
  AND U14614 ( .A(p_input[23424]), .B(p_input[13424]), .Z(n7307) );
  AND U14615 ( .A(n7308), .B(p_input[3423]), .Z(o[3423]) );
  AND U14616 ( .A(p_input[23423]), .B(p_input[13423]), .Z(n7308) );
  AND U14617 ( .A(n7309), .B(p_input[3422]), .Z(o[3422]) );
  AND U14618 ( .A(p_input[23422]), .B(p_input[13422]), .Z(n7309) );
  AND U14619 ( .A(n7310), .B(p_input[3421]), .Z(o[3421]) );
  AND U14620 ( .A(p_input[23421]), .B(p_input[13421]), .Z(n7310) );
  AND U14621 ( .A(n7311), .B(p_input[3420]), .Z(o[3420]) );
  AND U14622 ( .A(p_input[23420]), .B(p_input[13420]), .Z(n7311) );
  AND U14623 ( .A(n7312), .B(p_input[341]), .Z(o[341]) );
  AND U14624 ( .A(p_input[20341]), .B(p_input[10341]), .Z(n7312) );
  AND U14625 ( .A(n7313), .B(p_input[3419]), .Z(o[3419]) );
  AND U14626 ( .A(p_input[23419]), .B(p_input[13419]), .Z(n7313) );
  AND U14627 ( .A(n7314), .B(p_input[3418]), .Z(o[3418]) );
  AND U14628 ( .A(p_input[23418]), .B(p_input[13418]), .Z(n7314) );
  AND U14629 ( .A(n7315), .B(p_input[3417]), .Z(o[3417]) );
  AND U14630 ( .A(p_input[23417]), .B(p_input[13417]), .Z(n7315) );
  AND U14631 ( .A(n7316), .B(p_input[3416]), .Z(o[3416]) );
  AND U14632 ( .A(p_input[23416]), .B(p_input[13416]), .Z(n7316) );
  AND U14633 ( .A(n7317), .B(p_input[3415]), .Z(o[3415]) );
  AND U14634 ( .A(p_input[23415]), .B(p_input[13415]), .Z(n7317) );
  AND U14635 ( .A(n7318), .B(p_input[3414]), .Z(o[3414]) );
  AND U14636 ( .A(p_input[23414]), .B(p_input[13414]), .Z(n7318) );
  AND U14637 ( .A(n7319), .B(p_input[3413]), .Z(o[3413]) );
  AND U14638 ( .A(p_input[23413]), .B(p_input[13413]), .Z(n7319) );
  AND U14639 ( .A(n7320), .B(p_input[3412]), .Z(o[3412]) );
  AND U14640 ( .A(p_input[23412]), .B(p_input[13412]), .Z(n7320) );
  AND U14641 ( .A(n7321), .B(p_input[3411]), .Z(o[3411]) );
  AND U14642 ( .A(p_input[23411]), .B(p_input[13411]), .Z(n7321) );
  AND U14643 ( .A(n7322), .B(p_input[3410]), .Z(o[3410]) );
  AND U14644 ( .A(p_input[23410]), .B(p_input[13410]), .Z(n7322) );
  AND U14645 ( .A(n7323), .B(p_input[340]), .Z(o[340]) );
  AND U14646 ( .A(p_input[20340]), .B(p_input[10340]), .Z(n7323) );
  AND U14647 ( .A(n7324), .B(p_input[3409]), .Z(o[3409]) );
  AND U14648 ( .A(p_input[23409]), .B(p_input[13409]), .Z(n7324) );
  AND U14649 ( .A(n7325), .B(p_input[3408]), .Z(o[3408]) );
  AND U14650 ( .A(p_input[23408]), .B(p_input[13408]), .Z(n7325) );
  AND U14651 ( .A(n7326), .B(p_input[3407]), .Z(o[3407]) );
  AND U14652 ( .A(p_input[23407]), .B(p_input[13407]), .Z(n7326) );
  AND U14653 ( .A(n7327), .B(p_input[3406]), .Z(o[3406]) );
  AND U14654 ( .A(p_input[23406]), .B(p_input[13406]), .Z(n7327) );
  AND U14655 ( .A(n7328), .B(p_input[3405]), .Z(o[3405]) );
  AND U14656 ( .A(p_input[23405]), .B(p_input[13405]), .Z(n7328) );
  AND U14657 ( .A(n7329), .B(p_input[3404]), .Z(o[3404]) );
  AND U14658 ( .A(p_input[23404]), .B(p_input[13404]), .Z(n7329) );
  AND U14659 ( .A(n7330), .B(p_input[3403]), .Z(o[3403]) );
  AND U14660 ( .A(p_input[23403]), .B(p_input[13403]), .Z(n7330) );
  AND U14661 ( .A(n7331), .B(p_input[3402]), .Z(o[3402]) );
  AND U14662 ( .A(p_input[23402]), .B(p_input[13402]), .Z(n7331) );
  AND U14663 ( .A(n7332), .B(p_input[3401]), .Z(o[3401]) );
  AND U14664 ( .A(p_input[23401]), .B(p_input[13401]), .Z(n7332) );
  AND U14665 ( .A(n7333), .B(p_input[3400]), .Z(o[3400]) );
  AND U14666 ( .A(p_input[23400]), .B(p_input[13400]), .Z(n7333) );
  AND U14667 ( .A(n7334), .B(p_input[33]), .Z(o[33]) );
  AND U14668 ( .A(p_input[20033]), .B(p_input[10033]), .Z(n7334) );
  AND U14669 ( .A(n7335), .B(p_input[339]), .Z(o[339]) );
  AND U14670 ( .A(p_input[20339]), .B(p_input[10339]), .Z(n7335) );
  AND U14671 ( .A(n7336), .B(p_input[3399]), .Z(o[3399]) );
  AND U14672 ( .A(p_input[23399]), .B(p_input[13399]), .Z(n7336) );
  AND U14673 ( .A(n7337), .B(p_input[3398]), .Z(o[3398]) );
  AND U14674 ( .A(p_input[23398]), .B(p_input[13398]), .Z(n7337) );
  AND U14675 ( .A(n7338), .B(p_input[3397]), .Z(o[3397]) );
  AND U14676 ( .A(p_input[23397]), .B(p_input[13397]), .Z(n7338) );
  AND U14677 ( .A(n7339), .B(p_input[3396]), .Z(o[3396]) );
  AND U14678 ( .A(p_input[23396]), .B(p_input[13396]), .Z(n7339) );
  AND U14679 ( .A(n7340), .B(p_input[3395]), .Z(o[3395]) );
  AND U14680 ( .A(p_input[23395]), .B(p_input[13395]), .Z(n7340) );
  AND U14681 ( .A(n7341), .B(p_input[3394]), .Z(o[3394]) );
  AND U14682 ( .A(p_input[23394]), .B(p_input[13394]), .Z(n7341) );
  AND U14683 ( .A(n7342), .B(p_input[3393]), .Z(o[3393]) );
  AND U14684 ( .A(p_input[23393]), .B(p_input[13393]), .Z(n7342) );
  AND U14685 ( .A(n7343), .B(p_input[3392]), .Z(o[3392]) );
  AND U14686 ( .A(p_input[23392]), .B(p_input[13392]), .Z(n7343) );
  AND U14687 ( .A(n7344), .B(p_input[3391]), .Z(o[3391]) );
  AND U14688 ( .A(p_input[23391]), .B(p_input[13391]), .Z(n7344) );
  AND U14689 ( .A(n7345), .B(p_input[3390]), .Z(o[3390]) );
  AND U14690 ( .A(p_input[23390]), .B(p_input[13390]), .Z(n7345) );
  AND U14691 ( .A(n7346), .B(p_input[338]), .Z(o[338]) );
  AND U14692 ( .A(p_input[20338]), .B(p_input[10338]), .Z(n7346) );
  AND U14693 ( .A(n7347), .B(p_input[3389]), .Z(o[3389]) );
  AND U14694 ( .A(p_input[23389]), .B(p_input[13389]), .Z(n7347) );
  AND U14695 ( .A(n7348), .B(p_input[3388]), .Z(o[3388]) );
  AND U14696 ( .A(p_input[23388]), .B(p_input[13388]), .Z(n7348) );
  AND U14697 ( .A(n7349), .B(p_input[3387]), .Z(o[3387]) );
  AND U14698 ( .A(p_input[23387]), .B(p_input[13387]), .Z(n7349) );
  AND U14699 ( .A(n7350), .B(p_input[3386]), .Z(o[3386]) );
  AND U14700 ( .A(p_input[23386]), .B(p_input[13386]), .Z(n7350) );
  AND U14701 ( .A(n7351), .B(p_input[3385]), .Z(o[3385]) );
  AND U14702 ( .A(p_input[23385]), .B(p_input[13385]), .Z(n7351) );
  AND U14703 ( .A(n7352), .B(p_input[3384]), .Z(o[3384]) );
  AND U14704 ( .A(p_input[23384]), .B(p_input[13384]), .Z(n7352) );
  AND U14705 ( .A(n7353), .B(p_input[3383]), .Z(o[3383]) );
  AND U14706 ( .A(p_input[23383]), .B(p_input[13383]), .Z(n7353) );
  AND U14707 ( .A(n7354), .B(p_input[3382]), .Z(o[3382]) );
  AND U14708 ( .A(p_input[23382]), .B(p_input[13382]), .Z(n7354) );
  AND U14709 ( .A(n7355), .B(p_input[3381]), .Z(o[3381]) );
  AND U14710 ( .A(p_input[23381]), .B(p_input[13381]), .Z(n7355) );
  AND U14711 ( .A(n7356), .B(p_input[3380]), .Z(o[3380]) );
  AND U14712 ( .A(p_input[23380]), .B(p_input[13380]), .Z(n7356) );
  AND U14713 ( .A(n7357), .B(p_input[337]), .Z(o[337]) );
  AND U14714 ( .A(p_input[20337]), .B(p_input[10337]), .Z(n7357) );
  AND U14715 ( .A(n7358), .B(p_input[3379]), .Z(o[3379]) );
  AND U14716 ( .A(p_input[23379]), .B(p_input[13379]), .Z(n7358) );
  AND U14717 ( .A(n7359), .B(p_input[3378]), .Z(o[3378]) );
  AND U14718 ( .A(p_input[23378]), .B(p_input[13378]), .Z(n7359) );
  AND U14719 ( .A(n7360), .B(p_input[3377]), .Z(o[3377]) );
  AND U14720 ( .A(p_input[23377]), .B(p_input[13377]), .Z(n7360) );
  AND U14721 ( .A(n7361), .B(p_input[3376]), .Z(o[3376]) );
  AND U14722 ( .A(p_input[23376]), .B(p_input[13376]), .Z(n7361) );
  AND U14723 ( .A(n7362), .B(p_input[3375]), .Z(o[3375]) );
  AND U14724 ( .A(p_input[23375]), .B(p_input[13375]), .Z(n7362) );
  AND U14725 ( .A(n7363), .B(p_input[3374]), .Z(o[3374]) );
  AND U14726 ( .A(p_input[23374]), .B(p_input[13374]), .Z(n7363) );
  AND U14727 ( .A(n7364), .B(p_input[3373]), .Z(o[3373]) );
  AND U14728 ( .A(p_input[23373]), .B(p_input[13373]), .Z(n7364) );
  AND U14729 ( .A(n7365), .B(p_input[3372]), .Z(o[3372]) );
  AND U14730 ( .A(p_input[23372]), .B(p_input[13372]), .Z(n7365) );
  AND U14731 ( .A(n7366), .B(p_input[3371]), .Z(o[3371]) );
  AND U14732 ( .A(p_input[23371]), .B(p_input[13371]), .Z(n7366) );
  AND U14733 ( .A(n7367), .B(p_input[3370]), .Z(o[3370]) );
  AND U14734 ( .A(p_input[23370]), .B(p_input[13370]), .Z(n7367) );
  AND U14735 ( .A(n7368), .B(p_input[336]), .Z(o[336]) );
  AND U14736 ( .A(p_input[20336]), .B(p_input[10336]), .Z(n7368) );
  AND U14737 ( .A(n7369), .B(p_input[3369]), .Z(o[3369]) );
  AND U14738 ( .A(p_input[23369]), .B(p_input[13369]), .Z(n7369) );
  AND U14739 ( .A(n7370), .B(p_input[3368]), .Z(o[3368]) );
  AND U14740 ( .A(p_input[23368]), .B(p_input[13368]), .Z(n7370) );
  AND U14741 ( .A(n7371), .B(p_input[3367]), .Z(o[3367]) );
  AND U14742 ( .A(p_input[23367]), .B(p_input[13367]), .Z(n7371) );
  AND U14743 ( .A(n7372), .B(p_input[3366]), .Z(o[3366]) );
  AND U14744 ( .A(p_input[23366]), .B(p_input[13366]), .Z(n7372) );
  AND U14745 ( .A(n7373), .B(p_input[3365]), .Z(o[3365]) );
  AND U14746 ( .A(p_input[23365]), .B(p_input[13365]), .Z(n7373) );
  AND U14747 ( .A(n7374), .B(p_input[3364]), .Z(o[3364]) );
  AND U14748 ( .A(p_input[23364]), .B(p_input[13364]), .Z(n7374) );
  AND U14749 ( .A(n7375), .B(p_input[3363]), .Z(o[3363]) );
  AND U14750 ( .A(p_input[23363]), .B(p_input[13363]), .Z(n7375) );
  AND U14751 ( .A(n7376), .B(p_input[3362]), .Z(o[3362]) );
  AND U14752 ( .A(p_input[23362]), .B(p_input[13362]), .Z(n7376) );
  AND U14753 ( .A(n7377), .B(p_input[3361]), .Z(o[3361]) );
  AND U14754 ( .A(p_input[23361]), .B(p_input[13361]), .Z(n7377) );
  AND U14755 ( .A(n7378), .B(p_input[3360]), .Z(o[3360]) );
  AND U14756 ( .A(p_input[23360]), .B(p_input[13360]), .Z(n7378) );
  AND U14757 ( .A(n7379), .B(p_input[335]), .Z(o[335]) );
  AND U14758 ( .A(p_input[20335]), .B(p_input[10335]), .Z(n7379) );
  AND U14759 ( .A(n7380), .B(p_input[3359]), .Z(o[3359]) );
  AND U14760 ( .A(p_input[23359]), .B(p_input[13359]), .Z(n7380) );
  AND U14761 ( .A(n7381), .B(p_input[3358]), .Z(o[3358]) );
  AND U14762 ( .A(p_input[23358]), .B(p_input[13358]), .Z(n7381) );
  AND U14763 ( .A(n7382), .B(p_input[3357]), .Z(o[3357]) );
  AND U14764 ( .A(p_input[23357]), .B(p_input[13357]), .Z(n7382) );
  AND U14765 ( .A(n7383), .B(p_input[3356]), .Z(o[3356]) );
  AND U14766 ( .A(p_input[23356]), .B(p_input[13356]), .Z(n7383) );
  AND U14767 ( .A(n7384), .B(p_input[3355]), .Z(o[3355]) );
  AND U14768 ( .A(p_input[23355]), .B(p_input[13355]), .Z(n7384) );
  AND U14769 ( .A(n7385), .B(p_input[3354]), .Z(o[3354]) );
  AND U14770 ( .A(p_input[23354]), .B(p_input[13354]), .Z(n7385) );
  AND U14771 ( .A(n7386), .B(p_input[3353]), .Z(o[3353]) );
  AND U14772 ( .A(p_input[23353]), .B(p_input[13353]), .Z(n7386) );
  AND U14773 ( .A(n7387), .B(p_input[3352]), .Z(o[3352]) );
  AND U14774 ( .A(p_input[23352]), .B(p_input[13352]), .Z(n7387) );
  AND U14775 ( .A(n7388), .B(p_input[3351]), .Z(o[3351]) );
  AND U14776 ( .A(p_input[23351]), .B(p_input[13351]), .Z(n7388) );
  AND U14777 ( .A(n7389), .B(p_input[3350]), .Z(o[3350]) );
  AND U14778 ( .A(p_input[23350]), .B(p_input[13350]), .Z(n7389) );
  AND U14779 ( .A(n7390), .B(p_input[334]), .Z(o[334]) );
  AND U14780 ( .A(p_input[20334]), .B(p_input[10334]), .Z(n7390) );
  AND U14781 ( .A(n7391), .B(p_input[3349]), .Z(o[3349]) );
  AND U14782 ( .A(p_input[23349]), .B(p_input[13349]), .Z(n7391) );
  AND U14783 ( .A(n7392), .B(p_input[3348]), .Z(o[3348]) );
  AND U14784 ( .A(p_input[23348]), .B(p_input[13348]), .Z(n7392) );
  AND U14785 ( .A(n7393), .B(p_input[3347]), .Z(o[3347]) );
  AND U14786 ( .A(p_input[23347]), .B(p_input[13347]), .Z(n7393) );
  AND U14787 ( .A(n7394), .B(p_input[3346]), .Z(o[3346]) );
  AND U14788 ( .A(p_input[23346]), .B(p_input[13346]), .Z(n7394) );
  AND U14789 ( .A(n7395), .B(p_input[3345]), .Z(o[3345]) );
  AND U14790 ( .A(p_input[23345]), .B(p_input[13345]), .Z(n7395) );
  AND U14791 ( .A(n7396), .B(p_input[3344]), .Z(o[3344]) );
  AND U14792 ( .A(p_input[23344]), .B(p_input[13344]), .Z(n7396) );
  AND U14793 ( .A(n7397), .B(p_input[3343]), .Z(o[3343]) );
  AND U14794 ( .A(p_input[23343]), .B(p_input[13343]), .Z(n7397) );
  AND U14795 ( .A(n7398), .B(p_input[3342]), .Z(o[3342]) );
  AND U14796 ( .A(p_input[23342]), .B(p_input[13342]), .Z(n7398) );
  AND U14797 ( .A(n7399), .B(p_input[3341]), .Z(o[3341]) );
  AND U14798 ( .A(p_input[23341]), .B(p_input[13341]), .Z(n7399) );
  AND U14799 ( .A(n7400), .B(p_input[3340]), .Z(o[3340]) );
  AND U14800 ( .A(p_input[23340]), .B(p_input[13340]), .Z(n7400) );
  AND U14801 ( .A(n7401), .B(p_input[333]), .Z(o[333]) );
  AND U14802 ( .A(p_input[20333]), .B(p_input[10333]), .Z(n7401) );
  AND U14803 ( .A(n7402), .B(p_input[3339]), .Z(o[3339]) );
  AND U14804 ( .A(p_input[23339]), .B(p_input[13339]), .Z(n7402) );
  AND U14805 ( .A(n7403), .B(p_input[3338]), .Z(o[3338]) );
  AND U14806 ( .A(p_input[23338]), .B(p_input[13338]), .Z(n7403) );
  AND U14807 ( .A(n7404), .B(p_input[3337]), .Z(o[3337]) );
  AND U14808 ( .A(p_input[23337]), .B(p_input[13337]), .Z(n7404) );
  AND U14809 ( .A(n7405), .B(p_input[3336]), .Z(o[3336]) );
  AND U14810 ( .A(p_input[23336]), .B(p_input[13336]), .Z(n7405) );
  AND U14811 ( .A(n7406), .B(p_input[3335]), .Z(o[3335]) );
  AND U14812 ( .A(p_input[23335]), .B(p_input[13335]), .Z(n7406) );
  AND U14813 ( .A(n7407), .B(p_input[3334]), .Z(o[3334]) );
  AND U14814 ( .A(p_input[23334]), .B(p_input[13334]), .Z(n7407) );
  AND U14815 ( .A(n7408), .B(p_input[3333]), .Z(o[3333]) );
  AND U14816 ( .A(p_input[23333]), .B(p_input[13333]), .Z(n7408) );
  AND U14817 ( .A(n7409), .B(p_input[3332]), .Z(o[3332]) );
  AND U14818 ( .A(p_input[23332]), .B(p_input[13332]), .Z(n7409) );
  AND U14819 ( .A(n7410), .B(p_input[3331]), .Z(o[3331]) );
  AND U14820 ( .A(p_input[23331]), .B(p_input[13331]), .Z(n7410) );
  AND U14821 ( .A(n7411), .B(p_input[3330]), .Z(o[3330]) );
  AND U14822 ( .A(p_input[23330]), .B(p_input[13330]), .Z(n7411) );
  AND U14823 ( .A(n7412), .B(p_input[332]), .Z(o[332]) );
  AND U14824 ( .A(p_input[20332]), .B(p_input[10332]), .Z(n7412) );
  AND U14825 ( .A(n7413), .B(p_input[3329]), .Z(o[3329]) );
  AND U14826 ( .A(p_input[23329]), .B(p_input[13329]), .Z(n7413) );
  AND U14827 ( .A(n7414), .B(p_input[3328]), .Z(o[3328]) );
  AND U14828 ( .A(p_input[23328]), .B(p_input[13328]), .Z(n7414) );
  AND U14829 ( .A(n7415), .B(p_input[3327]), .Z(o[3327]) );
  AND U14830 ( .A(p_input[23327]), .B(p_input[13327]), .Z(n7415) );
  AND U14831 ( .A(n7416), .B(p_input[3326]), .Z(o[3326]) );
  AND U14832 ( .A(p_input[23326]), .B(p_input[13326]), .Z(n7416) );
  AND U14833 ( .A(n7417), .B(p_input[3325]), .Z(o[3325]) );
  AND U14834 ( .A(p_input[23325]), .B(p_input[13325]), .Z(n7417) );
  AND U14835 ( .A(n7418), .B(p_input[3324]), .Z(o[3324]) );
  AND U14836 ( .A(p_input[23324]), .B(p_input[13324]), .Z(n7418) );
  AND U14837 ( .A(n7419), .B(p_input[3323]), .Z(o[3323]) );
  AND U14838 ( .A(p_input[23323]), .B(p_input[13323]), .Z(n7419) );
  AND U14839 ( .A(n7420), .B(p_input[3322]), .Z(o[3322]) );
  AND U14840 ( .A(p_input[23322]), .B(p_input[13322]), .Z(n7420) );
  AND U14841 ( .A(n7421), .B(p_input[3321]), .Z(o[3321]) );
  AND U14842 ( .A(p_input[23321]), .B(p_input[13321]), .Z(n7421) );
  AND U14843 ( .A(n7422), .B(p_input[3320]), .Z(o[3320]) );
  AND U14844 ( .A(p_input[23320]), .B(p_input[13320]), .Z(n7422) );
  AND U14845 ( .A(n7423), .B(p_input[331]), .Z(o[331]) );
  AND U14846 ( .A(p_input[20331]), .B(p_input[10331]), .Z(n7423) );
  AND U14847 ( .A(n7424), .B(p_input[3319]), .Z(o[3319]) );
  AND U14848 ( .A(p_input[23319]), .B(p_input[13319]), .Z(n7424) );
  AND U14849 ( .A(n7425), .B(p_input[3318]), .Z(o[3318]) );
  AND U14850 ( .A(p_input[23318]), .B(p_input[13318]), .Z(n7425) );
  AND U14851 ( .A(n7426), .B(p_input[3317]), .Z(o[3317]) );
  AND U14852 ( .A(p_input[23317]), .B(p_input[13317]), .Z(n7426) );
  AND U14853 ( .A(n7427), .B(p_input[3316]), .Z(o[3316]) );
  AND U14854 ( .A(p_input[23316]), .B(p_input[13316]), .Z(n7427) );
  AND U14855 ( .A(n7428), .B(p_input[3315]), .Z(o[3315]) );
  AND U14856 ( .A(p_input[23315]), .B(p_input[13315]), .Z(n7428) );
  AND U14857 ( .A(n7429), .B(p_input[3314]), .Z(o[3314]) );
  AND U14858 ( .A(p_input[23314]), .B(p_input[13314]), .Z(n7429) );
  AND U14859 ( .A(n7430), .B(p_input[3313]), .Z(o[3313]) );
  AND U14860 ( .A(p_input[23313]), .B(p_input[13313]), .Z(n7430) );
  AND U14861 ( .A(n7431), .B(p_input[3312]), .Z(o[3312]) );
  AND U14862 ( .A(p_input[23312]), .B(p_input[13312]), .Z(n7431) );
  AND U14863 ( .A(n7432), .B(p_input[3311]), .Z(o[3311]) );
  AND U14864 ( .A(p_input[23311]), .B(p_input[13311]), .Z(n7432) );
  AND U14865 ( .A(n7433), .B(p_input[3310]), .Z(o[3310]) );
  AND U14866 ( .A(p_input[23310]), .B(p_input[13310]), .Z(n7433) );
  AND U14867 ( .A(n7434), .B(p_input[330]), .Z(o[330]) );
  AND U14868 ( .A(p_input[20330]), .B(p_input[10330]), .Z(n7434) );
  AND U14869 ( .A(n7435), .B(p_input[3309]), .Z(o[3309]) );
  AND U14870 ( .A(p_input[23309]), .B(p_input[13309]), .Z(n7435) );
  AND U14871 ( .A(n7436), .B(p_input[3308]), .Z(o[3308]) );
  AND U14872 ( .A(p_input[23308]), .B(p_input[13308]), .Z(n7436) );
  AND U14873 ( .A(n7437), .B(p_input[3307]), .Z(o[3307]) );
  AND U14874 ( .A(p_input[23307]), .B(p_input[13307]), .Z(n7437) );
  AND U14875 ( .A(n7438), .B(p_input[3306]), .Z(o[3306]) );
  AND U14876 ( .A(p_input[23306]), .B(p_input[13306]), .Z(n7438) );
  AND U14877 ( .A(n7439), .B(p_input[3305]), .Z(o[3305]) );
  AND U14878 ( .A(p_input[23305]), .B(p_input[13305]), .Z(n7439) );
  AND U14879 ( .A(n7440), .B(p_input[3304]), .Z(o[3304]) );
  AND U14880 ( .A(p_input[23304]), .B(p_input[13304]), .Z(n7440) );
  AND U14881 ( .A(n7441), .B(p_input[3303]), .Z(o[3303]) );
  AND U14882 ( .A(p_input[23303]), .B(p_input[13303]), .Z(n7441) );
  AND U14883 ( .A(n7442), .B(p_input[3302]), .Z(o[3302]) );
  AND U14884 ( .A(p_input[23302]), .B(p_input[13302]), .Z(n7442) );
  AND U14885 ( .A(n7443), .B(p_input[3301]), .Z(o[3301]) );
  AND U14886 ( .A(p_input[23301]), .B(p_input[13301]), .Z(n7443) );
  AND U14887 ( .A(n7444), .B(p_input[3300]), .Z(o[3300]) );
  AND U14888 ( .A(p_input[23300]), .B(p_input[13300]), .Z(n7444) );
  AND U14889 ( .A(n7445), .B(p_input[32]), .Z(o[32]) );
  AND U14890 ( .A(p_input[20032]), .B(p_input[10032]), .Z(n7445) );
  AND U14891 ( .A(n7446), .B(p_input[329]), .Z(o[329]) );
  AND U14892 ( .A(p_input[20329]), .B(p_input[10329]), .Z(n7446) );
  AND U14893 ( .A(n7447), .B(p_input[3299]), .Z(o[3299]) );
  AND U14894 ( .A(p_input[23299]), .B(p_input[13299]), .Z(n7447) );
  AND U14895 ( .A(n7448), .B(p_input[3298]), .Z(o[3298]) );
  AND U14896 ( .A(p_input[23298]), .B(p_input[13298]), .Z(n7448) );
  AND U14897 ( .A(n7449), .B(p_input[3297]), .Z(o[3297]) );
  AND U14898 ( .A(p_input[23297]), .B(p_input[13297]), .Z(n7449) );
  AND U14899 ( .A(n7450), .B(p_input[3296]), .Z(o[3296]) );
  AND U14900 ( .A(p_input[23296]), .B(p_input[13296]), .Z(n7450) );
  AND U14901 ( .A(n7451), .B(p_input[3295]), .Z(o[3295]) );
  AND U14902 ( .A(p_input[23295]), .B(p_input[13295]), .Z(n7451) );
  AND U14903 ( .A(n7452), .B(p_input[3294]), .Z(o[3294]) );
  AND U14904 ( .A(p_input[23294]), .B(p_input[13294]), .Z(n7452) );
  AND U14905 ( .A(n7453), .B(p_input[3293]), .Z(o[3293]) );
  AND U14906 ( .A(p_input[23293]), .B(p_input[13293]), .Z(n7453) );
  AND U14907 ( .A(n7454), .B(p_input[3292]), .Z(o[3292]) );
  AND U14908 ( .A(p_input[23292]), .B(p_input[13292]), .Z(n7454) );
  AND U14909 ( .A(n7455), .B(p_input[3291]), .Z(o[3291]) );
  AND U14910 ( .A(p_input[23291]), .B(p_input[13291]), .Z(n7455) );
  AND U14911 ( .A(n7456), .B(p_input[3290]), .Z(o[3290]) );
  AND U14912 ( .A(p_input[23290]), .B(p_input[13290]), .Z(n7456) );
  AND U14913 ( .A(n7457), .B(p_input[328]), .Z(o[328]) );
  AND U14914 ( .A(p_input[20328]), .B(p_input[10328]), .Z(n7457) );
  AND U14915 ( .A(n7458), .B(p_input[3289]), .Z(o[3289]) );
  AND U14916 ( .A(p_input[23289]), .B(p_input[13289]), .Z(n7458) );
  AND U14917 ( .A(n7459), .B(p_input[3288]), .Z(o[3288]) );
  AND U14918 ( .A(p_input[23288]), .B(p_input[13288]), .Z(n7459) );
  AND U14919 ( .A(n7460), .B(p_input[3287]), .Z(o[3287]) );
  AND U14920 ( .A(p_input[23287]), .B(p_input[13287]), .Z(n7460) );
  AND U14921 ( .A(n7461), .B(p_input[3286]), .Z(o[3286]) );
  AND U14922 ( .A(p_input[23286]), .B(p_input[13286]), .Z(n7461) );
  AND U14923 ( .A(n7462), .B(p_input[3285]), .Z(o[3285]) );
  AND U14924 ( .A(p_input[23285]), .B(p_input[13285]), .Z(n7462) );
  AND U14925 ( .A(n7463), .B(p_input[3284]), .Z(o[3284]) );
  AND U14926 ( .A(p_input[23284]), .B(p_input[13284]), .Z(n7463) );
  AND U14927 ( .A(n7464), .B(p_input[3283]), .Z(o[3283]) );
  AND U14928 ( .A(p_input[23283]), .B(p_input[13283]), .Z(n7464) );
  AND U14929 ( .A(n7465), .B(p_input[3282]), .Z(o[3282]) );
  AND U14930 ( .A(p_input[23282]), .B(p_input[13282]), .Z(n7465) );
  AND U14931 ( .A(n7466), .B(p_input[3281]), .Z(o[3281]) );
  AND U14932 ( .A(p_input[23281]), .B(p_input[13281]), .Z(n7466) );
  AND U14933 ( .A(n7467), .B(p_input[3280]), .Z(o[3280]) );
  AND U14934 ( .A(p_input[23280]), .B(p_input[13280]), .Z(n7467) );
  AND U14935 ( .A(n7468), .B(p_input[327]), .Z(o[327]) );
  AND U14936 ( .A(p_input[20327]), .B(p_input[10327]), .Z(n7468) );
  AND U14937 ( .A(n7469), .B(p_input[3279]), .Z(o[3279]) );
  AND U14938 ( .A(p_input[23279]), .B(p_input[13279]), .Z(n7469) );
  AND U14939 ( .A(n7470), .B(p_input[3278]), .Z(o[3278]) );
  AND U14940 ( .A(p_input[23278]), .B(p_input[13278]), .Z(n7470) );
  AND U14941 ( .A(n7471), .B(p_input[3277]), .Z(o[3277]) );
  AND U14942 ( .A(p_input[23277]), .B(p_input[13277]), .Z(n7471) );
  AND U14943 ( .A(n7472), .B(p_input[3276]), .Z(o[3276]) );
  AND U14944 ( .A(p_input[23276]), .B(p_input[13276]), .Z(n7472) );
  AND U14945 ( .A(n7473), .B(p_input[3275]), .Z(o[3275]) );
  AND U14946 ( .A(p_input[23275]), .B(p_input[13275]), .Z(n7473) );
  AND U14947 ( .A(n7474), .B(p_input[3274]), .Z(o[3274]) );
  AND U14948 ( .A(p_input[23274]), .B(p_input[13274]), .Z(n7474) );
  AND U14949 ( .A(n7475), .B(p_input[3273]), .Z(o[3273]) );
  AND U14950 ( .A(p_input[23273]), .B(p_input[13273]), .Z(n7475) );
  AND U14951 ( .A(n7476), .B(p_input[3272]), .Z(o[3272]) );
  AND U14952 ( .A(p_input[23272]), .B(p_input[13272]), .Z(n7476) );
  AND U14953 ( .A(n7477), .B(p_input[3271]), .Z(o[3271]) );
  AND U14954 ( .A(p_input[23271]), .B(p_input[13271]), .Z(n7477) );
  AND U14955 ( .A(n7478), .B(p_input[3270]), .Z(o[3270]) );
  AND U14956 ( .A(p_input[23270]), .B(p_input[13270]), .Z(n7478) );
  AND U14957 ( .A(n7479), .B(p_input[326]), .Z(o[326]) );
  AND U14958 ( .A(p_input[20326]), .B(p_input[10326]), .Z(n7479) );
  AND U14959 ( .A(n7480), .B(p_input[3269]), .Z(o[3269]) );
  AND U14960 ( .A(p_input[23269]), .B(p_input[13269]), .Z(n7480) );
  AND U14961 ( .A(n7481), .B(p_input[3268]), .Z(o[3268]) );
  AND U14962 ( .A(p_input[23268]), .B(p_input[13268]), .Z(n7481) );
  AND U14963 ( .A(n7482), .B(p_input[3267]), .Z(o[3267]) );
  AND U14964 ( .A(p_input[23267]), .B(p_input[13267]), .Z(n7482) );
  AND U14965 ( .A(n7483), .B(p_input[3266]), .Z(o[3266]) );
  AND U14966 ( .A(p_input[23266]), .B(p_input[13266]), .Z(n7483) );
  AND U14967 ( .A(n7484), .B(p_input[3265]), .Z(o[3265]) );
  AND U14968 ( .A(p_input[23265]), .B(p_input[13265]), .Z(n7484) );
  AND U14969 ( .A(n7485), .B(p_input[3264]), .Z(o[3264]) );
  AND U14970 ( .A(p_input[23264]), .B(p_input[13264]), .Z(n7485) );
  AND U14971 ( .A(n7486), .B(p_input[3263]), .Z(o[3263]) );
  AND U14972 ( .A(p_input[23263]), .B(p_input[13263]), .Z(n7486) );
  AND U14973 ( .A(n7487), .B(p_input[3262]), .Z(o[3262]) );
  AND U14974 ( .A(p_input[23262]), .B(p_input[13262]), .Z(n7487) );
  AND U14975 ( .A(n7488), .B(p_input[3261]), .Z(o[3261]) );
  AND U14976 ( .A(p_input[23261]), .B(p_input[13261]), .Z(n7488) );
  AND U14977 ( .A(n7489), .B(p_input[3260]), .Z(o[3260]) );
  AND U14978 ( .A(p_input[23260]), .B(p_input[13260]), .Z(n7489) );
  AND U14979 ( .A(n7490), .B(p_input[325]), .Z(o[325]) );
  AND U14980 ( .A(p_input[20325]), .B(p_input[10325]), .Z(n7490) );
  AND U14981 ( .A(n7491), .B(p_input[3259]), .Z(o[3259]) );
  AND U14982 ( .A(p_input[23259]), .B(p_input[13259]), .Z(n7491) );
  AND U14983 ( .A(n7492), .B(p_input[3258]), .Z(o[3258]) );
  AND U14984 ( .A(p_input[23258]), .B(p_input[13258]), .Z(n7492) );
  AND U14985 ( .A(n7493), .B(p_input[3257]), .Z(o[3257]) );
  AND U14986 ( .A(p_input[23257]), .B(p_input[13257]), .Z(n7493) );
  AND U14987 ( .A(n7494), .B(p_input[3256]), .Z(o[3256]) );
  AND U14988 ( .A(p_input[23256]), .B(p_input[13256]), .Z(n7494) );
  AND U14989 ( .A(n7495), .B(p_input[3255]), .Z(o[3255]) );
  AND U14990 ( .A(p_input[23255]), .B(p_input[13255]), .Z(n7495) );
  AND U14991 ( .A(n7496), .B(p_input[3254]), .Z(o[3254]) );
  AND U14992 ( .A(p_input[23254]), .B(p_input[13254]), .Z(n7496) );
  AND U14993 ( .A(n7497), .B(p_input[3253]), .Z(o[3253]) );
  AND U14994 ( .A(p_input[23253]), .B(p_input[13253]), .Z(n7497) );
  AND U14995 ( .A(n7498), .B(p_input[3252]), .Z(o[3252]) );
  AND U14996 ( .A(p_input[23252]), .B(p_input[13252]), .Z(n7498) );
  AND U14997 ( .A(n7499), .B(p_input[3251]), .Z(o[3251]) );
  AND U14998 ( .A(p_input[23251]), .B(p_input[13251]), .Z(n7499) );
  AND U14999 ( .A(n7500), .B(p_input[3250]), .Z(o[3250]) );
  AND U15000 ( .A(p_input[23250]), .B(p_input[13250]), .Z(n7500) );
  AND U15001 ( .A(n7501), .B(p_input[324]), .Z(o[324]) );
  AND U15002 ( .A(p_input[20324]), .B(p_input[10324]), .Z(n7501) );
  AND U15003 ( .A(n7502), .B(p_input[3249]), .Z(o[3249]) );
  AND U15004 ( .A(p_input[23249]), .B(p_input[13249]), .Z(n7502) );
  AND U15005 ( .A(n7503), .B(p_input[3248]), .Z(o[3248]) );
  AND U15006 ( .A(p_input[23248]), .B(p_input[13248]), .Z(n7503) );
  AND U15007 ( .A(n7504), .B(p_input[3247]), .Z(o[3247]) );
  AND U15008 ( .A(p_input[23247]), .B(p_input[13247]), .Z(n7504) );
  AND U15009 ( .A(n7505), .B(p_input[3246]), .Z(o[3246]) );
  AND U15010 ( .A(p_input[23246]), .B(p_input[13246]), .Z(n7505) );
  AND U15011 ( .A(n7506), .B(p_input[3245]), .Z(o[3245]) );
  AND U15012 ( .A(p_input[23245]), .B(p_input[13245]), .Z(n7506) );
  AND U15013 ( .A(n7507), .B(p_input[3244]), .Z(o[3244]) );
  AND U15014 ( .A(p_input[23244]), .B(p_input[13244]), .Z(n7507) );
  AND U15015 ( .A(n7508), .B(p_input[3243]), .Z(o[3243]) );
  AND U15016 ( .A(p_input[23243]), .B(p_input[13243]), .Z(n7508) );
  AND U15017 ( .A(n7509), .B(p_input[3242]), .Z(o[3242]) );
  AND U15018 ( .A(p_input[23242]), .B(p_input[13242]), .Z(n7509) );
  AND U15019 ( .A(n7510), .B(p_input[3241]), .Z(o[3241]) );
  AND U15020 ( .A(p_input[23241]), .B(p_input[13241]), .Z(n7510) );
  AND U15021 ( .A(n7511), .B(p_input[3240]), .Z(o[3240]) );
  AND U15022 ( .A(p_input[23240]), .B(p_input[13240]), .Z(n7511) );
  AND U15023 ( .A(n7512), .B(p_input[323]), .Z(o[323]) );
  AND U15024 ( .A(p_input[20323]), .B(p_input[10323]), .Z(n7512) );
  AND U15025 ( .A(n7513), .B(p_input[3239]), .Z(o[3239]) );
  AND U15026 ( .A(p_input[23239]), .B(p_input[13239]), .Z(n7513) );
  AND U15027 ( .A(n7514), .B(p_input[3238]), .Z(o[3238]) );
  AND U15028 ( .A(p_input[23238]), .B(p_input[13238]), .Z(n7514) );
  AND U15029 ( .A(n7515), .B(p_input[3237]), .Z(o[3237]) );
  AND U15030 ( .A(p_input[23237]), .B(p_input[13237]), .Z(n7515) );
  AND U15031 ( .A(n7516), .B(p_input[3236]), .Z(o[3236]) );
  AND U15032 ( .A(p_input[23236]), .B(p_input[13236]), .Z(n7516) );
  AND U15033 ( .A(n7517), .B(p_input[3235]), .Z(o[3235]) );
  AND U15034 ( .A(p_input[23235]), .B(p_input[13235]), .Z(n7517) );
  AND U15035 ( .A(n7518), .B(p_input[3234]), .Z(o[3234]) );
  AND U15036 ( .A(p_input[23234]), .B(p_input[13234]), .Z(n7518) );
  AND U15037 ( .A(n7519), .B(p_input[3233]), .Z(o[3233]) );
  AND U15038 ( .A(p_input[23233]), .B(p_input[13233]), .Z(n7519) );
  AND U15039 ( .A(n7520), .B(p_input[3232]), .Z(o[3232]) );
  AND U15040 ( .A(p_input[23232]), .B(p_input[13232]), .Z(n7520) );
  AND U15041 ( .A(n7521), .B(p_input[3231]), .Z(o[3231]) );
  AND U15042 ( .A(p_input[23231]), .B(p_input[13231]), .Z(n7521) );
  AND U15043 ( .A(n7522), .B(p_input[3230]), .Z(o[3230]) );
  AND U15044 ( .A(p_input[23230]), .B(p_input[13230]), .Z(n7522) );
  AND U15045 ( .A(n7523), .B(p_input[322]), .Z(o[322]) );
  AND U15046 ( .A(p_input[20322]), .B(p_input[10322]), .Z(n7523) );
  AND U15047 ( .A(n7524), .B(p_input[3229]), .Z(o[3229]) );
  AND U15048 ( .A(p_input[23229]), .B(p_input[13229]), .Z(n7524) );
  AND U15049 ( .A(n7525), .B(p_input[3228]), .Z(o[3228]) );
  AND U15050 ( .A(p_input[23228]), .B(p_input[13228]), .Z(n7525) );
  AND U15051 ( .A(n7526), .B(p_input[3227]), .Z(o[3227]) );
  AND U15052 ( .A(p_input[23227]), .B(p_input[13227]), .Z(n7526) );
  AND U15053 ( .A(n7527), .B(p_input[3226]), .Z(o[3226]) );
  AND U15054 ( .A(p_input[23226]), .B(p_input[13226]), .Z(n7527) );
  AND U15055 ( .A(n7528), .B(p_input[3225]), .Z(o[3225]) );
  AND U15056 ( .A(p_input[23225]), .B(p_input[13225]), .Z(n7528) );
  AND U15057 ( .A(n7529), .B(p_input[3224]), .Z(o[3224]) );
  AND U15058 ( .A(p_input[23224]), .B(p_input[13224]), .Z(n7529) );
  AND U15059 ( .A(n7530), .B(p_input[3223]), .Z(o[3223]) );
  AND U15060 ( .A(p_input[23223]), .B(p_input[13223]), .Z(n7530) );
  AND U15061 ( .A(n7531), .B(p_input[3222]), .Z(o[3222]) );
  AND U15062 ( .A(p_input[23222]), .B(p_input[13222]), .Z(n7531) );
  AND U15063 ( .A(n7532), .B(p_input[3221]), .Z(o[3221]) );
  AND U15064 ( .A(p_input[23221]), .B(p_input[13221]), .Z(n7532) );
  AND U15065 ( .A(n7533), .B(p_input[3220]), .Z(o[3220]) );
  AND U15066 ( .A(p_input[23220]), .B(p_input[13220]), .Z(n7533) );
  AND U15067 ( .A(n7534), .B(p_input[321]), .Z(o[321]) );
  AND U15068 ( .A(p_input[20321]), .B(p_input[10321]), .Z(n7534) );
  AND U15069 ( .A(n7535), .B(p_input[3219]), .Z(o[3219]) );
  AND U15070 ( .A(p_input[23219]), .B(p_input[13219]), .Z(n7535) );
  AND U15071 ( .A(n7536), .B(p_input[3218]), .Z(o[3218]) );
  AND U15072 ( .A(p_input[23218]), .B(p_input[13218]), .Z(n7536) );
  AND U15073 ( .A(n7537), .B(p_input[3217]), .Z(o[3217]) );
  AND U15074 ( .A(p_input[23217]), .B(p_input[13217]), .Z(n7537) );
  AND U15075 ( .A(n7538), .B(p_input[3216]), .Z(o[3216]) );
  AND U15076 ( .A(p_input[23216]), .B(p_input[13216]), .Z(n7538) );
  AND U15077 ( .A(n7539), .B(p_input[3215]), .Z(o[3215]) );
  AND U15078 ( .A(p_input[23215]), .B(p_input[13215]), .Z(n7539) );
  AND U15079 ( .A(n7540), .B(p_input[3214]), .Z(o[3214]) );
  AND U15080 ( .A(p_input[23214]), .B(p_input[13214]), .Z(n7540) );
  AND U15081 ( .A(n7541), .B(p_input[3213]), .Z(o[3213]) );
  AND U15082 ( .A(p_input[23213]), .B(p_input[13213]), .Z(n7541) );
  AND U15083 ( .A(n7542), .B(p_input[3212]), .Z(o[3212]) );
  AND U15084 ( .A(p_input[23212]), .B(p_input[13212]), .Z(n7542) );
  AND U15085 ( .A(n7543), .B(p_input[3211]), .Z(o[3211]) );
  AND U15086 ( .A(p_input[23211]), .B(p_input[13211]), .Z(n7543) );
  AND U15087 ( .A(n7544), .B(p_input[3210]), .Z(o[3210]) );
  AND U15088 ( .A(p_input[23210]), .B(p_input[13210]), .Z(n7544) );
  AND U15089 ( .A(n7545), .B(p_input[320]), .Z(o[320]) );
  AND U15090 ( .A(p_input[20320]), .B(p_input[10320]), .Z(n7545) );
  AND U15091 ( .A(n7546), .B(p_input[3209]), .Z(o[3209]) );
  AND U15092 ( .A(p_input[23209]), .B(p_input[13209]), .Z(n7546) );
  AND U15093 ( .A(n7547), .B(p_input[3208]), .Z(o[3208]) );
  AND U15094 ( .A(p_input[23208]), .B(p_input[13208]), .Z(n7547) );
  AND U15095 ( .A(n7548), .B(p_input[3207]), .Z(o[3207]) );
  AND U15096 ( .A(p_input[23207]), .B(p_input[13207]), .Z(n7548) );
  AND U15097 ( .A(n7549), .B(p_input[3206]), .Z(o[3206]) );
  AND U15098 ( .A(p_input[23206]), .B(p_input[13206]), .Z(n7549) );
  AND U15099 ( .A(n7550), .B(p_input[3205]), .Z(o[3205]) );
  AND U15100 ( .A(p_input[23205]), .B(p_input[13205]), .Z(n7550) );
  AND U15101 ( .A(n7551), .B(p_input[3204]), .Z(o[3204]) );
  AND U15102 ( .A(p_input[23204]), .B(p_input[13204]), .Z(n7551) );
  AND U15103 ( .A(n7552), .B(p_input[3203]), .Z(o[3203]) );
  AND U15104 ( .A(p_input[23203]), .B(p_input[13203]), .Z(n7552) );
  AND U15105 ( .A(n7553), .B(p_input[3202]), .Z(o[3202]) );
  AND U15106 ( .A(p_input[23202]), .B(p_input[13202]), .Z(n7553) );
  AND U15107 ( .A(n7554), .B(p_input[3201]), .Z(o[3201]) );
  AND U15108 ( .A(p_input[23201]), .B(p_input[13201]), .Z(n7554) );
  AND U15109 ( .A(n7555), .B(p_input[3200]), .Z(o[3200]) );
  AND U15110 ( .A(p_input[23200]), .B(p_input[13200]), .Z(n7555) );
  AND U15111 ( .A(n7556), .B(p_input[31]), .Z(o[31]) );
  AND U15112 ( .A(p_input[20031]), .B(p_input[10031]), .Z(n7556) );
  AND U15113 ( .A(n7557), .B(p_input[319]), .Z(o[319]) );
  AND U15114 ( .A(p_input[20319]), .B(p_input[10319]), .Z(n7557) );
  AND U15115 ( .A(n7558), .B(p_input[3199]), .Z(o[3199]) );
  AND U15116 ( .A(p_input[23199]), .B(p_input[13199]), .Z(n7558) );
  AND U15117 ( .A(n7559), .B(p_input[3198]), .Z(o[3198]) );
  AND U15118 ( .A(p_input[23198]), .B(p_input[13198]), .Z(n7559) );
  AND U15119 ( .A(n7560), .B(p_input[3197]), .Z(o[3197]) );
  AND U15120 ( .A(p_input[23197]), .B(p_input[13197]), .Z(n7560) );
  AND U15121 ( .A(n7561), .B(p_input[3196]), .Z(o[3196]) );
  AND U15122 ( .A(p_input[23196]), .B(p_input[13196]), .Z(n7561) );
  AND U15123 ( .A(n7562), .B(p_input[3195]), .Z(o[3195]) );
  AND U15124 ( .A(p_input[23195]), .B(p_input[13195]), .Z(n7562) );
  AND U15125 ( .A(n7563), .B(p_input[3194]), .Z(o[3194]) );
  AND U15126 ( .A(p_input[23194]), .B(p_input[13194]), .Z(n7563) );
  AND U15127 ( .A(n7564), .B(p_input[3193]), .Z(o[3193]) );
  AND U15128 ( .A(p_input[23193]), .B(p_input[13193]), .Z(n7564) );
  AND U15129 ( .A(n7565), .B(p_input[3192]), .Z(o[3192]) );
  AND U15130 ( .A(p_input[23192]), .B(p_input[13192]), .Z(n7565) );
  AND U15131 ( .A(n7566), .B(p_input[3191]), .Z(o[3191]) );
  AND U15132 ( .A(p_input[23191]), .B(p_input[13191]), .Z(n7566) );
  AND U15133 ( .A(n7567), .B(p_input[3190]), .Z(o[3190]) );
  AND U15134 ( .A(p_input[23190]), .B(p_input[13190]), .Z(n7567) );
  AND U15135 ( .A(n7568), .B(p_input[318]), .Z(o[318]) );
  AND U15136 ( .A(p_input[20318]), .B(p_input[10318]), .Z(n7568) );
  AND U15137 ( .A(n7569), .B(p_input[3189]), .Z(o[3189]) );
  AND U15138 ( .A(p_input[23189]), .B(p_input[13189]), .Z(n7569) );
  AND U15139 ( .A(n7570), .B(p_input[3188]), .Z(o[3188]) );
  AND U15140 ( .A(p_input[23188]), .B(p_input[13188]), .Z(n7570) );
  AND U15141 ( .A(n7571), .B(p_input[3187]), .Z(o[3187]) );
  AND U15142 ( .A(p_input[23187]), .B(p_input[13187]), .Z(n7571) );
  AND U15143 ( .A(n7572), .B(p_input[3186]), .Z(o[3186]) );
  AND U15144 ( .A(p_input[23186]), .B(p_input[13186]), .Z(n7572) );
  AND U15145 ( .A(n7573), .B(p_input[3185]), .Z(o[3185]) );
  AND U15146 ( .A(p_input[23185]), .B(p_input[13185]), .Z(n7573) );
  AND U15147 ( .A(n7574), .B(p_input[3184]), .Z(o[3184]) );
  AND U15148 ( .A(p_input[23184]), .B(p_input[13184]), .Z(n7574) );
  AND U15149 ( .A(n7575), .B(p_input[3183]), .Z(o[3183]) );
  AND U15150 ( .A(p_input[23183]), .B(p_input[13183]), .Z(n7575) );
  AND U15151 ( .A(n7576), .B(p_input[3182]), .Z(o[3182]) );
  AND U15152 ( .A(p_input[23182]), .B(p_input[13182]), .Z(n7576) );
  AND U15153 ( .A(n7577), .B(p_input[3181]), .Z(o[3181]) );
  AND U15154 ( .A(p_input[23181]), .B(p_input[13181]), .Z(n7577) );
  AND U15155 ( .A(n7578), .B(p_input[3180]), .Z(o[3180]) );
  AND U15156 ( .A(p_input[23180]), .B(p_input[13180]), .Z(n7578) );
  AND U15157 ( .A(n7579), .B(p_input[317]), .Z(o[317]) );
  AND U15158 ( .A(p_input[20317]), .B(p_input[10317]), .Z(n7579) );
  AND U15159 ( .A(n7580), .B(p_input[3179]), .Z(o[3179]) );
  AND U15160 ( .A(p_input[23179]), .B(p_input[13179]), .Z(n7580) );
  AND U15161 ( .A(n7581), .B(p_input[3178]), .Z(o[3178]) );
  AND U15162 ( .A(p_input[23178]), .B(p_input[13178]), .Z(n7581) );
  AND U15163 ( .A(n7582), .B(p_input[3177]), .Z(o[3177]) );
  AND U15164 ( .A(p_input[23177]), .B(p_input[13177]), .Z(n7582) );
  AND U15165 ( .A(n7583), .B(p_input[3176]), .Z(o[3176]) );
  AND U15166 ( .A(p_input[23176]), .B(p_input[13176]), .Z(n7583) );
  AND U15167 ( .A(n7584), .B(p_input[3175]), .Z(o[3175]) );
  AND U15168 ( .A(p_input[23175]), .B(p_input[13175]), .Z(n7584) );
  AND U15169 ( .A(n7585), .B(p_input[3174]), .Z(o[3174]) );
  AND U15170 ( .A(p_input[23174]), .B(p_input[13174]), .Z(n7585) );
  AND U15171 ( .A(n7586), .B(p_input[3173]), .Z(o[3173]) );
  AND U15172 ( .A(p_input[23173]), .B(p_input[13173]), .Z(n7586) );
  AND U15173 ( .A(n7587), .B(p_input[3172]), .Z(o[3172]) );
  AND U15174 ( .A(p_input[23172]), .B(p_input[13172]), .Z(n7587) );
  AND U15175 ( .A(n7588), .B(p_input[3171]), .Z(o[3171]) );
  AND U15176 ( .A(p_input[23171]), .B(p_input[13171]), .Z(n7588) );
  AND U15177 ( .A(n7589), .B(p_input[3170]), .Z(o[3170]) );
  AND U15178 ( .A(p_input[23170]), .B(p_input[13170]), .Z(n7589) );
  AND U15179 ( .A(n7590), .B(p_input[316]), .Z(o[316]) );
  AND U15180 ( .A(p_input[20316]), .B(p_input[10316]), .Z(n7590) );
  AND U15181 ( .A(n7591), .B(p_input[3169]), .Z(o[3169]) );
  AND U15182 ( .A(p_input[23169]), .B(p_input[13169]), .Z(n7591) );
  AND U15183 ( .A(n7592), .B(p_input[3168]), .Z(o[3168]) );
  AND U15184 ( .A(p_input[23168]), .B(p_input[13168]), .Z(n7592) );
  AND U15185 ( .A(n7593), .B(p_input[3167]), .Z(o[3167]) );
  AND U15186 ( .A(p_input[23167]), .B(p_input[13167]), .Z(n7593) );
  AND U15187 ( .A(n7594), .B(p_input[3166]), .Z(o[3166]) );
  AND U15188 ( .A(p_input[23166]), .B(p_input[13166]), .Z(n7594) );
  AND U15189 ( .A(n7595), .B(p_input[3165]), .Z(o[3165]) );
  AND U15190 ( .A(p_input[23165]), .B(p_input[13165]), .Z(n7595) );
  AND U15191 ( .A(n7596), .B(p_input[3164]), .Z(o[3164]) );
  AND U15192 ( .A(p_input[23164]), .B(p_input[13164]), .Z(n7596) );
  AND U15193 ( .A(n7597), .B(p_input[3163]), .Z(o[3163]) );
  AND U15194 ( .A(p_input[23163]), .B(p_input[13163]), .Z(n7597) );
  AND U15195 ( .A(n7598), .B(p_input[3162]), .Z(o[3162]) );
  AND U15196 ( .A(p_input[23162]), .B(p_input[13162]), .Z(n7598) );
  AND U15197 ( .A(n7599), .B(p_input[3161]), .Z(o[3161]) );
  AND U15198 ( .A(p_input[23161]), .B(p_input[13161]), .Z(n7599) );
  AND U15199 ( .A(n7600), .B(p_input[3160]), .Z(o[3160]) );
  AND U15200 ( .A(p_input[23160]), .B(p_input[13160]), .Z(n7600) );
  AND U15201 ( .A(n7601), .B(p_input[315]), .Z(o[315]) );
  AND U15202 ( .A(p_input[20315]), .B(p_input[10315]), .Z(n7601) );
  AND U15203 ( .A(n7602), .B(p_input[3159]), .Z(o[3159]) );
  AND U15204 ( .A(p_input[23159]), .B(p_input[13159]), .Z(n7602) );
  AND U15205 ( .A(n7603), .B(p_input[3158]), .Z(o[3158]) );
  AND U15206 ( .A(p_input[23158]), .B(p_input[13158]), .Z(n7603) );
  AND U15207 ( .A(n7604), .B(p_input[3157]), .Z(o[3157]) );
  AND U15208 ( .A(p_input[23157]), .B(p_input[13157]), .Z(n7604) );
  AND U15209 ( .A(n7605), .B(p_input[3156]), .Z(o[3156]) );
  AND U15210 ( .A(p_input[23156]), .B(p_input[13156]), .Z(n7605) );
  AND U15211 ( .A(n7606), .B(p_input[3155]), .Z(o[3155]) );
  AND U15212 ( .A(p_input[23155]), .B(p_input[13155]), .Z(n7606) );
  AND U15213 ( .A(n7607), .B(p_input[3154]), .Z(o[3154]) );
  AND U15214 ( .A(p_input[23154]), .B(p_input[13154]), .Z(n7607) );
  AND U15215 ( .A(n7608), .B(p_input[3153]), .Z(o[3153]) );
  AND U15216 ( .A(p_input[23153]), .B(p_input[13153]), .Z(n7608) );
  AND U15217 ( .A(n7609), .B(p_input[3152]), .Z(o[3152]) );
  AND U15218 ( .A(p_input[23152]), .B(p_input[13152]), .Z(n7609) );
  AND U15219 ( .A(n7610), .B(p_input[3151]), .Z(o[3151]) );
  AND U15220 ( .A(p_input[23151]), .B(p_input[13151]), .Z(n7610) );
  AND U15221 ( .A(n7611), .B(p_input[3150]), .Z(o[3150]) );
  AND U15222 ( .A(p_input[23150]), .B(p_input[13150]), .Z(n7611) );
  AND U15223 ( .A(n7612), .B(p_input[314]), .Z(o[314]) );
  AND U15224 ( .A(p_input[20314]), .B(p_input[10314]), .Z(n7612) );
  AND U15225 ( .A(n7613), .B(p_input[3149]), .Z(o[3149]) );
  AND U15226 ( .A(p_input[23149]), .B(p_input[13149]), .Z(n7613) );
  AND U15227 ( .A(n7614), .B(p_input[3148]), .Z(o[3148]) );
  AND U15228 ( .A(p_input[23148]), .B(p_input[13148]), .Z(n7614) );
  AND U15229 ( .A(n7615), .B(p_input[3147]), .Z(o[3147]) );
  AND U15230 ( .A(p_input[23147]), .B(p_input[13147]), .Z(n7615) );
  AND U15231 ( .A(n7616), .B(p_input[3146]), .Z(o[3146]) );
  AND U15232 ( .A(p_input[23146]), .B(p_input[13146]), .Z(n7616) );
  AND U15233 ( .A(n7617), .B(p_input[3145]), .Z(o[3145]) );
  AND U15234 ( .A(p_input[23145]), .B(p_input[13145]), .Z(n7617) );
  AND U15235 ( .A(n7618), .B(p_input[3144]), .Z(o[3144]) );
  AND U15236 ( .A(p_input[23144]), .B(p_input[13144]), .Z(n7618) );
  AND U15237 ( .A(n7619), .B(p_input[3143]), .Z(o[3143]) );
  AND U15238 ( .A(p_input[23143]), .B(p_input[13143]), .Z(n7619) );
  AND U15239 ( .A(n7620), .B(p_input[3142]), .Z(o[3142]) );
  AND U15240 ( .A(p_input[23142]), .B(p_input[13142]), .Z(n7620) );
  AND U15241 ( .A(n7621), .B(p_input[3141]), .Z(o[3141]) );
  AND U15242 ( .A(p_input[23141]), .B(p_input[13141]), .Z(n7621) );
  AND U15243 ( .A(n7622), .B(p_input[3140]), .Z(o[3140]) );
  AND U15244 ( .A(p_input[23140]), .B(p_input[13140]), .Z(n7622) );
  AND U15245 ( .A(n7623), .B(p_input[313]), .Z(o[313]) );
  AND U15246 ( .A(p_input[20313]), .B(p_input[10313]), .Z(n7623) );
  AND U15247 ( .A(n7624), .B(p_input[3139]), .Z(o[3139]) );
  AND U15248 ( .A(p_input[23139]), .B(p_input[13139]), .Z(n7624) );
  AND U15249 ( .A(n7625), .B(p_input[3138]), .Z(o[3138]) );
  AND U15250 ( .A(p_input[23138]), .B(p_input[13138]), .Z(n7625) );
  AND U15251 ( .A(n7626), .B(p_input[3137]), .Z(o[3137]) );
  AND U15252 ( .A(p_input[23137]), .B(p_input[13137]), .Z(n7626) );
  AND U15253 ( .A(n7627), .B(p_input[3136]), .Z(o[3136]) );
  AND U15254 ( .A(p_input[23136]), .B(p_input[13136]), .Z(n7627) );
  AND U15255 ( .A(n7628), .B(p_input[3135]), .Z(o[3135]) );
  AND U15256 ( .A(p_input[23135]), .B(p_input[13135]), .Z(n7628) );
  AND U15257 ( .A(n7629), .B(p_input[3134]), .Z(o[3134]) );
  AND U15258 ( .A(p_input[23134]), .B(p_input[13134]), .Z(n7629) );
  AND U15259 ( .A(n7630), .B(p_input[3133]), .Z(o[3133]) );
  AND U15260 ( .A(p_input[23133]), .B(p_input[13133]), .Z(n7630) );
  AND U15261 ( .A(n7631), .B(p_input[3132]), .Z(o[3132]) );
  AND U15262 ( .A(p_input[23132]), .B(p_input[13132]), .Z(n7631) );
  AND U15263 ( .A(n7632), .B(p_input[3131]), .Z(o[3131]) );
  AND U15264 ( .A(p_input[23131]), .B(p_input[13131]), .Z(n7632) );
  AND U15265 ( .A(n7633), .B(p_input[3130]), .Z(o[3130]) );
  AND U15266 ( .A(p_input[23130]), .B(p_input[13130]), .Z(n7633) );
  AND U15267 ( .A(n7634), .B(p_input[312]), .Z(o[312]) );
  AND U15268 ( .A(p_input[20312]), .B(p_input[10312]), .Z(n7634) );
  AND U15269 ( .A(n7635), .B(p_input[3129]), .Z(o[3129]) );
  AND U15270 ( .A(p_input[23129]), .B(p_input[13129]), .Z(n7635) );
  AND U15271 ( .A(n7636), .B(p_input[3128]), .Z(o[3128]) );
  AND U15272 ( .A(p_input[23128]), .B(p_input[13128]), .Z(n7636) );
  AND U15273 ( .A(n7637), .B(p_input[3127]), .Z(o[3127]) );
  AND U15274 ( .A(p_input[23127]), .B(p_input[13127]), .Z(n7637) );
  AND U15275 ( .A(n7638), .B(p_input[3126]), .Z(o[3126]) );
  AND U15276 ( .A(p_input[23126]), .B(p_input[13126]), .Z(n7638) );
  AND U15277 ( .A(n7639), .B(p_input[3125]), .Z(o[3125]) );
  AND U15278 ( .A(p_input[23125]), .B(p_input[13125]), .Z(n7639) );
  AND U15279 ( .A(n7640), .B(p_input[3124]), .Z(o[3124]) );
  AND U15280 ( .A(p_input[23124]), .B(p_input[13124]), .Z(n7640) );
  AND U15281 ( .A(n7641), .B(p_input[3123]), .Z(o[3123]) );
  AND U15282 ( .A(p_input[23123]), .B(p_input[13123]), .Z(n7641) );
  AND U15283 ( .A(n7642), .B(p_input[3122]), .Z(o[3122]) );
  AND U15284 ( .A(p_input[23122]), .B(p_input[13122]), .Z(n7642) );
  AND U15285 ( .A(n7643), .B(p_input[3121]), .Z(o[3121]) );
  AND U15286 ( .A(p_input[23121]), .B(p_input[13121]), .Z(n7643) );
  AND U15287 ( .A(n7644), .B(p_input[3120]), .Z(o[3120]) );
  AND U15288 ( .A(p_input[23120]), .B(p_input[13120]), .Z(n7644) );
  AND U15289 ( .A(n7645), .B(p_input[311]), .Z(o[311]) );
  AND U15290 ( .A(p_input[20311]), .B(p_input[10311]), .Z(n7645) );
  AND U15291 ( .A(n7646), .B(p_input[3119]), .Z(o[3119]) );
  AND U15292 ( .A(p_input[23119]), .B(p_input[13119]), .Z(n7646) );
  AND U15293 ( .A(n7647), .B(p_input[3118]), .Z(o[3118]) );
  AND U15294 ( .A(p_input[23118]), .B(p_input[13118]), .Z(n7647) );
  AND U15295 ( .A(n7648), .B(p_input[3117]), .Z(o[3117]) );
  AND U15296 ( .A(p_input[23117]), .B(p_input[13117]), .Z(n7648) );
  AND U15297 ( .A(n7649), .B(p_input[3116]), .Z(o[3116]) );
  AND U15298 ( .A(p_input[23116]), .B(p_input[13116]), .Z(n7649) );
  AND U15299 ( .A(n7650), .B(p_input[3115]), .Z(o[3115]) );
  AND U15300 ( .A(p_input[23115]), .B(p_input[13115]), .Z(n7650) );
  AND U15301 ( .A(n7651), .B(p_input[3114]), .Z(o[3114]) );
  AND U15302 ( .A(p_input[23114]), .B(p_input[13114]), .Z(n7651) );
  AND U15303 ( .A(n7652), .B(p_input[3113]), .Z(o[3113]) );
  AND U15304 ( .A(p_input[23113]), .B(p_input[13113]), .Z(n7652) );
  AND U15305 ( .A(n7653), .B(p_input[3112]), .Z(o[3112]) );
  AND U15306 ( .A(p_input[23112]), .B(p_input[13112]), .Z(n7653) );
  AND U15307 ( .A(n7654), .B(p_input[3111]), .Z(o[3111]) );
  AND U15308 ( .A(p_input[23111]), .B(p_input[13111]), .Z(n7654) );
  AND U15309 ( .A(n7655), .B(p_input[3110]), .Z(o[3110]) );
  AND U15310 ( .A(p_input[23110]), .B(p_input[13110]), .Z(n7655) );
  AND U15311 ( .A(n7656), .B(p_input[310]), .Z(o[310]) );
  AND U15312 ( .A(p_input[20310]), .B(p_input[10310]), .Z(n7656) );
  AND U15313 ( .A(n7657), .B(p_input[3109]), .Z(o[3109]) );
  AND U15314 ( .A(p_input[23109]), .B(p_input[13109]), .Z(n7657) );
  AND U15315 ( .A(n7658), .B(p_input[3108]), .Z(o[3108]) );
  AND U15316 ( .A(p_input[23108]), .B(p_input[13108]), .Z(n7658) );
  AND U15317 ( .A(n7659), .B(p_input[3107]), .Z(o[3107]) );
  AND U15318 ( .A(p_input[23107]), .B(p_input[13107]), .Z(n7659) );
  AND U15319 ( .A(n7660), .B(p_input[3106]), .Z(o[3106]) );
  AND U15320 ( .A(p_input[23106]), .B(p_input[13106]), .Z(n7660) );
  AND U15321 ( .A(n7661), .B(p_input[3105]), .Z(o[3105]) );
  AND U15322 ( .A(p_input[23105]), .B(p_input[13105]), .Z(n7661) );
  AND U15323 ( .A(n7662), .B(p_input[3104]), .Z(o[3104]) );
  AND U15324 ( .A(p_input[23104]), .B(p_input[13104]), .Z(n7662) );
  AND U15325 ( .A(n7663), .B(p_input[3103]), .Z(o[3103]) );
  AND U15326 ( .A(p_input[23103]), .B(p_input[13103]), .Z(n7663) );
  AND U15327 ( .A(n7664), .B(p_input[3102]), .Z(o[3102]) );
  AND U15328 ( .A(p_input[23102]), .B(p_input[13102]), .Z(n7664) );
  AND U15329 ( .A(n7665), .B(p_input[3101]), .Z(o[3101]) );
  AND U15330 ( .A(p_input[23101]), .B(p_input[13101]), .Z(n7665) );
  AND U15331 ( .A(n7666), .B(p_input[3100]), .Z(o[3100]) );
  AND U15332 ( .A(p_input[23100]), .B(p_input[13100]), .Z(n7666) );
  AND U15333 ( .A(n7667), .B(p_input[30]), .Z(o[30]) );
  AND U15334 ( .A(p_input[20030]), .B(p_input[10030]), .Z(n7667) );
  AND U15335 ( .A(n7668), .B(p_input[309]), .Z(o[309]) );
  AND U15336 ( .A(p_input[20309]), .B(p_input[10309]), .Z(n7668) );
  AND U15337 ( .A(n7669), .B(p_input[3099]), .Z(o[3099]) );
  AND U15338 ( .A(p_input[23099]), .B(p_input[13099]), .Z(n7669) );
  AND U15339 ( .A(n7670), .B(p_input[3098]), .Z(o[3098]) );
  AND U15340 ( .A(p_input[23098]), .B(p_input[13098]), .Z(n7670) );
  AND U15341 ( .A(n7671), .B(p_input[3097]), .Z(o[3097]) );
  AND U15342 ( .A(p_input[23097]), .B(p_input[13097]), .Z(n7671) );
  AND U15343 ( .A(n7672), .B(p_input[3096]), .Z(o[3096]) );
  AND U15344 ( .A(p_input[23096]), .B(p_input[13096]), .Z(n7672) );
  AND U15345 ( .A(n7673), .B(p_input[3095]), .Z(o[3095]) );
  AND U15346 ( .A(p_input[23095]), .B(p_input[13095]), .Z(n7673) );
  AND U15347 ( .A(n7674), .B(p_input[3094]), .Z(o[3094]) );
  AND U15348 ( .A(p_input[23094]), .B(p_input[13094]), .Z(n7674) );
  AND U15349 ( .A(n7675), .B(p_input[3093]), .Z(o[3093]) );
  AND U15350 ( .A(p_input[23093]), .B(p_input[13093]), .Z(n7675) );
  AND U15351 ( .A(n7676), .B(p_input[3092]), .Z(o[3092]) );
  AND U15352 ( .A(p_input[23092]), .B(p_input[13092]), .Z(n7676) );
  AND U15353 ( .A(n7677), .B(p_input[3091]), .Z(o[3091]) );
  AND U15354 ( .A(p_input[23091]), .B(p_input[13091]), .Z(n7677) );
  AND U15355 ( .A(n7678), .B(p_input[3090]), .Z(o[3090]) );
  AND U15356 ( .A(p_input[23090]), .B(p_input[13090]), .Z(n7678) );
  AND U15357 ( .A(n7679), .B(p_input[308]), .Z(o[308]) );
  AND U15358 ( .A(p_input[20308]), .B(p_input[10308]), .Z(n7679) );
  AND U15359 ( .A(n7680), .B(p_input[3089]), .Z(o[3089]) );
  AND U15360 ( .A(p_input[23089]), .B(p_input[13089]), .Z(n7680) );
  AND U15361 ( .A(n7681), .B(p_input[3088]), .Z(o[3088]) );
  AND U15362 ( .A(p_input[23088]), .B(p_input[13088]), .Z(n7681) );
  AND U15363 ( .A(n7682), .B(p_input[3087]), .Z(o[3087]) );
  AND U15364 ( .A(p_input[23087]), .B(p_input[13087]), .Z(n7682) );
  AND U15365 ( .A(n7683), .B(p_input[3086]), .Z(o[3086]) );
  AND U15366 ( .A(p_input[23086]), .B(p_input[13086]), .Z(n7683) );
  AND U15367 ( .A(n7684), .B(p_input[3085]), .Z(o[3085]) );
  AND U15368 ( .A(p_input[23085]), .B(p_input[13085]), .Z(n7684) );
  AND U15369 ( .A(n7685), .B(p_input[3084]), .Z(o[3084]) );
  AND U15370 ( .A(p_input[23084]), .B(p_input[13084]), .Z(n7685) );
  AND U15371 ( .A(n7686), .B(p_input[3083]), .Z(o[3083]) );
  AND U15372 ( .A(p_input[23083]), .B(p_input[13083]), .Z(n7686) );
  AND U15373 ( .A(n7687), .B(p_input[3082]), .Z(o[3082]) );
  AND U15374 ( .A(p_input[23082]), .B(p_input[13082]), .Z(n7687) );
  AND U15375 ( .A(n7688), .B(p_input[3081]), .Z(o[3081]) );
  AND U15376 ( .A(p_input[23081]), .B(p_input[13081]), .Z(n7688) );
  AND U15377 ( .A(n7689), .B(p_input[3080]), .Z(o[3080]) );
  AND U15378 ( .A(p_input[23080]), .B(p_input[13080]), .Z(n7689) );
  AND U15379 ( .A(n7690), .B(p_input[307]), .Z(o[307]) );
  AND U15380 ( .A(p_input[20307]), .B(p_input[10307]), .Z(n7690) );
  AND U15381 ( .A(n7691), .B(p_input[3079]), .Z(o[3079]) );
  AND U15382 ( .A(p_input[23079]), .B(p_input[13079]), .Z(n7691) );
  AND U15383 ( .A(n7692), .B(p_input[3078]), .Z(o[3078]) );
  AND U15384 ( .A(p_input[23078]), .B(p_input[13078]), .Z(n7692) );
  AND U15385 ( .A(n7693), .B(p_input[3077]), .Z(o[3077]) );
  AND U15386 ( .A(p_input[23077]), .B(p_input[13077]), .Z(n7693) );
  AND U15387 ( .A(n7694), .B(p_input[3076]), .Z(o[3076]) );
  AND U15388 ( .A(p_input[23076]), .B(p_input[13076]), .Z(n7694) );
  AND U15389 ( .A(n7695), .B(p_input[3075]), .Z(o[3075]) );
  AND U15390 ( .A(p_input[23075]), .B(p_input[13075]), .Z(n7695) );
  AND U15391 ( .A(n7696), .B(p_input[3074]), .Z(o[3074]) );
  AND U15392 ( .A(p_input[23074]), .B(p_input[13074]), .Z(n7696) );
  AND U15393 ( .A(n7697), .B(p_input[3073]), .Z(o[3073]) );
  AND U15394 ( .A(p_input[23073]), .B(p_input[13073]), .Z(n7697) );
  AND U15395 ( .A(n7698), .B(p_input[3072]), .Z(o[3072]) );
  AND U15396 ( .A(p_input[23072]), .B(p_input[13072]), .Z(n7698) );
  AND U15397 ( .A(n7699), .B(p_input[3071]), .Z(o[3071]) );
  AND U15398 ( .A(p_input[23071]), .B(p_input[13071]), .Z(n7699) );
  AND U15399 ( .A(n7700), .B(p_input[3070]), .Z(o[3070]) );
  AND U15400 ( .A(p_input[23070]), .B(p_input[13070]), .Z(n7700) );
  AND U15401 ( .A(n7701), .B(p_input[306]), .Z(o[306]) );
  AND U15402 ( .A(p_input[20306]), .B(p_input[10306]), .Z(n7701) );
  AND U15403 ( .A(n7702), .B(p_input[3069]), .Z(o[3069]) );
  AND U15404 ( .A(p_input[23069]), .B(p_input[13069]), .Z(n7702) );
  AND U15405 ( .A(n7703), .B(p_input[3068]), .Z(o[3068]) );
  AND U15406 ( .A(p_input[23068]), .B(p_input[13068]), .Z(n7703) );
  AND U15407 ( .A(n7704), .B(p_input[3067]), .Z(o[3067]) );
  AND U15408 ( .A(p_input[23067]), .B(p_input[13067]), .Z(n7704) );
  AND U15409 ( .A(n7705), .B(p_input[3066]), .Z(o[3066]) );
  AND U15410 ( .A(p_input[23066]), .B(p_input[13066]), .Z(n7705) );
  AND U15411 ( .A(n7706), .B(p_input[3065]), .Z(o[3065]) );
  AND U15412 ( .A(p_input[23065]), .B(p_input[13065]), .Z(n7706) );
  AND U15413 ( .A(n7707), .B(p_input[3064]), .Z(o[3064]) );
  AND U15414 ( .A(p_input[23064]), .B(p_input[13064]), .Z(n7707) );
  AND U15415 ( .A(n7708), .B(p_input[3063]), .Z(o[3063]) );
  AND U15416 ( .A(p_input[23063]), .B(p_input[13063]), .Z(n7708) );
  AND U15417 ( .A(n7709), .B(p_input[3062]), .Z(o[3062]) );
  AND U15418 ( .A(p_input[23062]), .B(p_input[13062]), .Z(n7709) );
  AND U15419 ( .A(n7710), .B(p_input[3061]), .Z(o[3061]) );
  AND U15420 ( .A(p_input[23061]), .B(p_input[13061]), .Z(n7710) );
  AND U15421 ( .A(n7711), .B(p_input[3060]), .Z(o[3060]) );
  AND U15422 ( .A(p_input[23060]), .B(p_input[13060]), .Z(n7711) );
  AND U15423 ( .A(n7712), .B(p_input[305]), .Z(o[305]) );
  AND U15424 ( .A(p_input[20305]), .B(p_input[10305]), .Z(n7712) );
  AND U15425 ( .A(n7713), .B(p_input[3059]), .Z(o[3059]) );
  AND U15426 ( .A(p_input[23059]), .B(p_input[13059]), .Z(n7713) );
  AND U15427 ( .A(n7714), .B(p_input[3058]), .Z(o[3058]) );
  AND U15428 ( .A(p_input[23058]), .B(p_input[13058]), .Z(n7714) );
  AND U15429 ( .A(n7715), .B(p_input[3057]), .Z(o[3057]) );
  AND U15430 ( .A(p_input[23057]), .B(p_input[13057]), .Z(n7715) );
  AND U15431 ( .A(n7716), .B(p_input[3056]), .Z(o[3056]) );
  AND U15432 ( .A(p_input[23056]), .B(p_input[13056]), .Z(n7716) );
  AND U15433 ( .A(n7717), .B(p_input[3055]), .Z(o[3055]) );
  AND U15434 ( .A(p_input[23055]), .B(p_input[13055]), .Z(n7717) );
  AND U15435 ( .A(n7718), .B(p_input[3054]), .Z(o[3054]) );
  AND U15436 ( .A(p_input[23054]), .B(p_input[13054]), .Z(n7718) );
  AND U15437 ( .A(n7719), .B(p_input[3053]), .Z(o[3053]) );
  AND U15438 ( .A(p_input[23053]), .B(p_input[13053]), .Z(n7719) );
  AND U15439 ( .A(n7720), .B(p_input[3052]), .Z(o[3052]) );
  AND U15440 ( .A(p_input[23052]), .B(p_input[13052]), .Z(n7720) );
  AND U15441 ( .A(n7721), .B(p_input[3051]), .Z(o[3051]) );
  AND U15442 ( .A(p_input[23051]), .B(p_input[13051]), .Z(n7721) );
  AND U15443 ( .A(n7722), .B(p_input[3050]), .Z(o[3050]) );
  AND U15444 ( .A(p_input[23050]), .B(p_input[13050]), .Z(n7722) );
  AND U15445 ( .A(n7723), .B(p_input[304]), .Z(o[304]) );
  AND U15446 ( .A(p_input[20304]), .B(p_input[10304]), .Z(n7723) );
  AND U15447 ( .A(n7724), .B(p_input[3049]), .Z(o[3049]) );
  AND U15448 ( .A(p_input[23049]), .B(p_input[13049]), .Z(n7724) );
  AND U15449 ( .A(n7725), .B(p_input[3048]), .Z(o[3048]) );
  AND U15450 ( .A(p_input[23048]), .B(p_input[13048]), .Z(n7725) );
  AND U15451 ( .A(n7726), .B(p_input[3047]), .Z(o[3047]) );
  AND U15452 ( .A(p_input[23047]), .B(p_input[13047]), .Z(n7726) );
  AND U15453 ( .A(n7727), .B(p_input[3046]), .Z(o[3046]) );
  AND U15454 ( .A(p_input[23046]), .B(p_input[13046]), .Z(n7727) );
  AND U15455 ( .A(n7728), .B(p_input[3045]), .Z(o[3045]) );
  AND U15456 ( .A(p_input[23045]), .B(p_input[13045]), .Z(n7728) );
  AND U15457 ( .A(n7729), .B(p_input[3044]), .Z(o[3044]) );
  AND U15458 ( .A(p_input[23044]), .B(p_input[13044]), .Z(n7729) );
  AND U15459 ( .A(n7730), .B(p_input[3043]), .Z(o[3043]) );
  AND U15460 ( .A(p_input[23043]), .B(p_input[13043]), .Z(n7730) );
  AND U15461 ( .A(n7731), .B(p_input[3042]), .Z(o[3042]) );
  AND U15462 ( .A(p_input[23042]), .B(p_input[13042]), .Z(n7731) );
  AND U15463 ( .A(n7732), .B(p_input[3041]), .Z(o[3041]) );
  AND U15464 ( .A(p_input[23041]), .B(p_input[13041]), .Z(n7732) );
  AND U15465 ( .A(n7733), .B(p_input[3040]), .Z(o[3040]) );
  AND U15466 ( .A(p_input[23040]), .B(p_input[13040]), .Z(n7733) );
  AND U15467 ( .A(n7734), .B(p_input[303]), .Z(o[303]) );
  AND U15468 ( .A(p_input[20303]), .B(p_input[10303]), .Z(n7734) );
  AND U15469 ( .A(n7735), .B(p_input[3039]), .Z(o[3039]) );
  AND U15470 ( .A(p_input[23039]), .B(p_input[13039]), .Z(n7735) );
  AND U15471 ( .A(n7736), .B(p_input[3038]), .Z(o[3038]) );
  AND U15472 ( .A(p_input[23038]), .B(p_input[13038]), .Z(n7736) );
  AND U15473 ( .A(n7737), .B(p_input[3037]), .Z(o[3037]) );
  AND U15474 ( .A(p_input[23037]), .B(p_input[13037]), .Z(n7737) );
  AND U15475 ( .A(n7738), .B(p_input[3036]), .Z(o[3036]) );
  AND U15476 ( .A(p_input[23036]), .B(p_input[13036]), .Z(n7738) );
  AND U15477 ( .A(n7739), .B(p_input[3035]), .Z(o[3035]) );
  AND U15478 ( .A(p_input[23035]), .B(p_input[13035]), .Z(n7739) );
  AND U15479 ( .A(n7740), .B(p_input[3034]), .Z(o[3034]) );
  AND U15480 ( .A(p_input[23034]), .B(p_input[13034]), .Z(n7740) );
  AND U15481 ( .A(n7741), .B(p_input[3033]), .Z(o[3033]) );
  AND U15482 ( .A(p_input[23033]), .B(p_input[13033]), .Z(n7741) );
  AND U15483 ( .A(n7742), .B(p_input[3032]), .Z(o[3032]) );
  AND U15484 ( .A(p_input[23032]), .B(p_input[13032]), .Z(n7742) );
  AND U15485 ( .A(n7743), .B(p_input[3031]), .Z(o[3031]) );
  AND U15486 ( .A(p_input[23031]), .B(p_input[13031]), .Z(n7743) );
  AND U15487 ( .A(n7744), .B(p_input[3030]), .Z(o[3030]) );
  AND U15488 ( .A(p_input[23030]), .B(p_input[13030]), .Z(n7744) );
  AND U15489 ( .A(n7745), .B(p_input[302]), .Z(o[302]) );
  AND U15490 ( .A(p_input[20302]), .B(p_input[10302]), .Z(n7745) );
  AND U15491 ( .A(n7746), .B(p_input[3029]), .Z(o[3029]) );
  AND U15492 ( .A(p_input[23029]), .B(p_input[13029]), .Z(n7746) );
  AND U15493 ( .A(n7747), .B(p_input[3028]), .Z(o[3028]) );
  AND U15494 ( .A(p_input[23028]), .B(p_input[13028]), .Z(n7747) );
  AND U15495 ( .A(n7748), .B(p_input[3027]), .Z(o[3027]) );
  AND U15496 ( .A(p_input[23027]), .B(p_input[13027]), .Z(n7748) );
  AND U15497 ( .A(n7749), .B(p_input[3026]), .Z(o[3026]) );
  AND U15498 ( .A(p_input[23026]), .B(p_input[13026]), .Z(n7749) );
  AND U15499 ( .A(n7750), .B(p_input[3025]), .Z(o[3025]) );
  AND U15500 ( .A(p_input[23025]), .B(p_input[13025]), .Z(n7750) );
  AND U15501 ( .A(n7751), .B(p_input[3024]), .Z(o[3024]) );
  AND U15502 ( .A(p_input[23024]), .B(p_input[13024]), .Z(n7751) );
  AND U15503 ( .A(n7752), .B(p_input[3023]), .Z(o[3023]) );
  AND U15504 ( .A(p_input[23023]), .B(p_input[13023]), .Z(n7752) );
  AND U15505 ( .A(n7753), .B(p_input[3022]), .Z(o[3022]) );
  AND U15506 ( .A(p_input[23022]), .B(p_input[13022]), .Z(n7753) );
  AND U15507 ( .A(n7754), .B(p_input[3021]), .Z(o[3021]) );
  AND U15508 ( .A(p_input[23021]), .B(p_input[13021]), .Z(n7754) );
  AND U15509 ( .A(n7755), .B(p_input[3020]), .Z(o[3020]) );
  AND U15510 ( .A(p_input[23020]), .B(p_input[13020]), .Z(n7755) );
  AND U15511 ( .A(n7756), .B(p_input[301]), .Z(o[301]) );
  AND U15512 ( .A(p_input[20301]), .B(p_input[10301]), .Z(n7756) );
  AND U15513 ( .A(n7757), .B(p_input[3019]), .Z(o[3019]) );
  AND U15514 ( .A(p_input[23019]), .B(p_input[13019]), .Z(n7757) );
  AND U15515 ( .A(n7758), .B(p_input[3018]), .Z(o[3018]) );
  AND U15516 ( .A(p_input[23018]), .B(p_input[13018]), .Z(n7758) );
  AND U15517 ( .A(n7759), .B(p_input[3017]), .Z(o[3017]) );
  AND U15518 ( .A(p_input[23017]), .B(p_input[13017]), .Z(n7759) );
  AND U15519 ( .A(n7760), .B(p_input[3016]), .Z(o[3016]) );
  AND U15520 ( .A(p_input[23016]), .B(p_input[13016]), .Z(n7760) );
  AND U15521 ( .A(n7761), .B(p_input[3015]), .Z(o[3015]) );
  AND U15522 ( .A(p_input[23015]), .B(p_input[13015]), .Z(n7761) );
  AND U15523 ( .A(n7762), .B(p_input[3014]), .Z(o[3014]) );
  AND U15524 ( .A(p_input[23014]), .B(p_input[13014]), .Z(n7762) );
  AND U15525 ( .A(n7763), .B(p_input[3013]), .Z(o[3013]) );
  AND U15526 ( .A(p_input[23013]), .B(p_input[13013]), .Z(n7763) );
  AND U15527 ( .A(n7764), .B(p_input[3012]), .Z(o[3012]) );
  AND U15528 ( .A(p_input[23012]), .B(p_input[13012]), .Z(n7764) );
  AND U15529 ( .A(n7765), .B(p_input[3011]), .Z(o[3011]) );
  AND U15530 ( .A(p_input[23011]), .B(p_input[13011]), .Z(n7765) );
  AND U15531 ( .A(n7766), .B(p_input[3010]), .Z(o[3010]) );
  AND U15532 ( .A(p_input[23010]), .B(p_input[13010]), .Z(n7766) );
  AND U15533 ( .A(n7767), .B(p_input[300]), .Z(o[300]) );
  AND U15534 ( .A(p_input[20300]), .B(p_input[10300]), .Z(n7767) );
  AND U15535 ( .A(n7768), .B(p_input[3009]), .Z(o[3009]) );
  AND U15536 ( .A(p_input[23009]), .B(p_input[13009]), .Z(n7768) );
  AND U15537 ( .A(n7769), .B(p_input[3008]), .Z(o[3008]) );
  AND U15538 ( .A(p_input[23008]), .B(p_input[13008]), .Z(n7769) );
  AND U15539 ( .A(n7770), .B(p_input[3007]), .Z(o[3007]) );
  AND U15540 ( .A(p_input[23007]), .B(p_input[13007]), .Z(n7770) );
  AND U15541 ( .A(n7771), .B(p_input[3006]), .Z(o[3006]) );
  AND U15542 ( .A(p_input[23006]), .B(p_input[13006]), .Z(n7771) );
  AND U15543 ( .A(n7772), .B(p_input[3005]), .Z(o[3005]) );
  AND U15544 ( .A(p_input[23005]), .B(p_input[13005]), .Z(n7772) );
  AND U15545 ( .A(n7773), .B(p_input[3004]), .Z(o[3004]) );
  AND U15546 ( .A(p_input[23004]), .B(p_input[13004]), .Z(n7773) );
  AND U15547 ( .A(n7774), .B(p_input[3003]), .Z(o[3003]) );
  AND U15548 ( .A(p_input[23003]), .B(p_input[13003]), .Z(n7774) );
  AND U15549 ( .A(n7775), .B(p_input[3002]), .Z(o[3002]) );
  AND U15550 ( .A(p_input[23002]), .B(p_input[13002]), .Z(n7775) );
  AND U15551 ( .A(n7776), .B(p_input[3001]), .Z(o[3001]) );
  AND U15552 ( .A(p_input[23001]), .B(p_input[13001]), .Z(n7776) );
  AND U15553 ( .A(n7777), .B(p_input[3000]), .Z(o[3000]) );
  AND U15554 ( .A(p_input[23000]), .B(p_input[13000]), .Z(n7777) );
  AND U15555 ( .A(n7778), .B(p_input[2]), .Z(o[2]) );
  AND U15556 ( .A(p_input[20002]), .B(p_input[10002]), .Z(n7778) );
  AND U15557 ( .A(n7779), .B(p_input[29]), .Z(o[29]) );
  AND U15558 ( .A(p_input[20029]), .B(p_input[10029]), .Z(n7779) );
  AND U15559 ( .A(n7780), .B(p_input[299]), .Z(o[299]) );
  AND U15560 ( .A(p_input[20299]), .B(p_input[10299]), .Z(n7780) );
  AND U15561 ( .A(n7781), .B(p_input[2999]), .Z(o[2999]) );
  AND U15562 ( .A(p_input[22999]), .B(p_input[12999]), .Z(n7781) );
  AND U15563 ( .A(n7782), .B(p_input[2998]), .Z(o[2998]) );
  AND U15564 ( .A(p_input[22998]), .B(p_input[12998]), .Z(n7782) );
  AND U15565 ( .A(n7783), .B(p_input[2997]), .Z(o[2997]) );
  AND U15566 ( .A(p_input[22997]), .B(p_input[12997]), .Z(n7783) );
  AND U15567 ( .A(n7784), .B(p_input[2996]), .Z(o[2996]) );
  AND U15568 ( .A(p_input[22996]), .B(p_input[12996]), .Z(n7784) );
  AND U15569 ( .A(n7785), .B(p_input[2995]), .Z(o[2995]) );
  AND U15570 ( .A(p_input[22995]), .B(p_input[12995]), .Z(n7785) );
  AND U15571 ( .A(n7786), .B(p_input[2994]), .Z(o[2994]) );
  AND U15572 ( .A(p_input[22994]), .B(p_input[12994]), .Z(n7786) );
  AND U15573 ( .A(n7787), .B(p_input[2993]), .Z(o[2993]) );
  AND U15574 ( .A(p_input[22993]), .B(p_input[12993]), .Z(n7787) );
  AND U15575 ( .A(n7788), .B(p_input[2992]), .Z(o[2992]) );
  AND U15576 ( .A(p_input[22992]), .B(p_input[12992]), .Z(n7788) );
  AND U15577 ( .A(n7789), .B(p_input[2991]), .Z(o[2991]) );
  AND U15578 ( .A(p_input[22991]), .B(p_input[12991]), .Z(n7789) );
  AND U15579 ( .A(n7790), .B(p_input[2990]), .Z(o[2990]) );
  AND U15580 ( .A(p_input[22990]), .B(p_input[12990]), .Z(n7790) );
  AND U15581 ( .A(n7791), .B(p_input[298]), .Z(o[298]) );
  AND U15582 ( .A(p_input[20298]), .B(p_input[10298]), .Z(n7791) );
  AND U15583 ( .A(n7792), .B(p_input[2989]), .Z(o[2989]) );
  AND U15584 ( .A(p_input[22989]), .B(p_input[12989]), .Z(n7792) );
  AND U15585 ( .A(n7793), .B(p_input[2988]), .Z(o[2988]) );
  AND U15586 ( .A(p_input[22988]), .B(p_input[12988]), .Z(n7793) );
  AND U15587 ( .A(n7794), .B(p_input[2987]), .Z(o[2987]) );
  AND U15588 ( .A(p_input[22987]), .B(p_input[12987]), .Z(n7794) );
  AND U15589 ( .A(n7795), .B(p_input[2986]), .Z(o[2986]) );
  AND U15590 ( .A(p_input[22986]), .B(p_input[12986]), .Z(n7795) );
  AND U15591 ( .A(n7796), .B(p_input[2985]), .Z(o[2985]) );
  AND U15592 ( .A(p_input[22985]), .B(p_input[12985]), .Z(n7796) );
  AND U15593 ( .A(n7797), .B(p_input[2984]), .Z(o[2984]) );
  AND U15594 ( .A(p_input[22984]), .B(p_input[12984]), .Z(n7797) );
  AND U15595 ( .A(n7798), .B(p_input[2983]), .Z(o[2983]) );
  AND U15596 ( .A(p_input[22983]), .B(p_input[12983]), .Z(n7798) );
  AND U15597 ( .A(n7799), .B(p_input[2982]), .Z(o[2982]) );
  AND U15598 ( .A(p_input[22982]), .B(p_input[12982]), .Z(n7799) );
  AND U15599 ( .A(n7800), .B(p_input[2981]), .Z(o[2981]) );
  AND U15600 ( .A(p_input[22981]), .B(p_input[12981]), .Z(n7800) );
  AND U15601 ( .A(n7801), .B(p_input[2980]), .Z(o[2980]) );
  AND U15602 ( .A(p_input[22980]), .B(p_input[12980]), .Z(n7801) );
  AND U15603 ( .A(n7802), .B(p_input[297]), .Z(o[297]) );
  AND U15604 ( .A(p_input[20297]), .B(p_input[10297]), .Z(n7802) );
  AND U15605 ( .A(n7803), .B(p_input[2979]), .Z(o[2979]) );
  AND U15606 ( .A(p_input[22979]), .B(p_input[12979]), .Z(n7803) );
  AND U15607 ( .A(n7804), .B(p_input[2978]), .Z(o[2978]) );
  AND U15608 ( .A(p_input[22978]), .B(p_input[12978]), .Z(n7804) );
  AND U15609 ( .A(n7805), .B(p_input[2977]), .Z(o[2977]) );
  AND U15610 ( .A(p_input[22977]), .B(p_input[12977]), .Z(n7805) );
  AND U15611 ( .A(n7806), .B(p_input[2976]), .Z(o[2976]) );
  AND U15612 ( .A(p_input[22976]), .B(p_input[12976]), .Z(n7806) );
  AND U15613 ( .A(n7807), .B(p_input[2975]), .Z(o[2975]) );
  AND U15614 ( .A(p_input[22975]), .B(p_input[12975]), .Z(n7807) );
  AND U15615 ( .A(n7808), .B(p_input[2974]), .Z(o[2974]) );
  AND U15616 ( .A(p_input[22974]), .B(p_input[12974]), .Z(n7808) );
  AND U15617 ( .A(n7809), .B(p_input[2973]), .Z(o[2973]) );
  AND U15618 ( .A(p_input[22973]), .B(p_input[12973]), .Z(n7809) );
  AND U15619 ( .A(n7810), .B(p_input[2972]), .Z(o[2972]) );
  AND U15620 ( .A(p_input[22972]), .B(p_input[12972]), .Z(n7810) );
  AND U15621 ( .A(n7811), .B(p_input[2971]), .Z(o[2971]) );
  AND U15622 ( .A(p_input[22971]), .B(p_input[12971]), .Z(n7811) );
  AND U15623 ( .A(n7812), .B(p_input[2970]), .Z(o[2970]) );
  AND U15624 ( .A(p_input[22970]), .B(p_input[12970]), .Z(n7812) );
  AND U15625 ( .A(n7813), .B(p_input[296]), .Z(o[296]) );
  AND U15626 ( .A(p_input[20296]), .B(p_input[10296]), .Z(n7813) );
  AND U15627 ( .A(n7814), .B(p_input[2969]), .Z(o[2969]) );
  AND U15628 ( .A(p_input[22969]), .B(p_input[12969]), .Z(n7814) );
  AND U15629 ( .A(n7815), .B(p_input[2968]), .Z(o[2968]) );
  AND U15630 ( .A(p_input[22968]), .B(p_input[12968]), .Z(n7815) );
  AND U15631 ( .A(n7816), .B(p_input[2967]), .Z(o[2967]) );
  AND U15632 ( .A(p_input[22967]), .B(p_input[12967]), .Z(n7816) );
  AND U15633 ( .A(n7817), .B(p_input[2966]), .Z(o[2966]) );
  AND U15634 ( .A(p_input[22966]), .B(p_input[12966]), .Z(n7817) );
  AND U15635 ( .A(n7818), .B(p_input[2965]), .Z(o[2965]) );
  AND U15636 ( .A(p_input[22965]), .B(p_input[12965]), .Z(n7818) );
  AND U15637 ( .A(n7819), .B(p_input[2964]), .Z(o[2964]) );
  AND U15638 ( .A(p_input[22964]), .B(p_input[12964]), .Z(n7819) );
  AND U15639 ( .A(n7820), .B(p_input[2963]), .Z(o[2963]) );
  AND U15640 ( .A(p_input[22963]), .B(p_input[12963]), .Z(n7820) );
  AND U15641 ( .A(n7821), .B(p_input[2962]), .Z(o[2962]) );
  AND U15642 ( .A(p_input[22962]), .B(p_input[12962]), .Z(n7821) );
  AND U15643 ( .A(n7822), .B(p_input[2961]), .Z(o[2961]) );
  AND U15644 ( .A(p_input[22961]), .B(p_input[12961]), .Z(n7822) );
  AND U15645 ( .A(n7823), .B(p_input[2960]), .Z(o[2960]) );
  AND U15646 ( .A(p_input[22960]), .B(p_input[12960]), .Z(n7823) );
  AND U15647 ( .A(n7824), .B(p_input[295]), .Z(o[295]) );
  AND U15648 ( .A(p_input[20295]), .B(p_input[10295]), .Z(n7824) );
  AND U15649 ( .A(n7825), .B(p_input[2959]), .Z(o[2959]) );
  AND U15650 ( .A(p_input[22959]), .B(p_input[12959]), .Z(n7825) );
  AND U15651 ( .A(n7826), .B(p_input[2958]), .Z(o[2958]) );
  AND U15652 ( .A(p_input[22958]), .B(p_input[12958]), .Z(n7826) );
  AND U15653 ( .A(n7827), .B(p_input[2957]), .Z(o[2957]) );
  AND U15654 ( .A(p_input[22957]), .B(p_input[12957]), .Z(n7827) );
  AND U15655 ( .A(n7828), .B(p_input[2956]), .Z(o[2956]) );
  AND U15656 ( .A(p_input[22956]), .B(p_input[12956]), .Z(n7828) );
  AND U15657 ( .A(n7829), .B(p_input[2955]), .Z(o[2955]) );
  AND U15658 ( .A(p_input[22955]), .B(p_input[12955]), .Z(n7829) );
  AND U15659 ( .A(n7830), .B(p_input[2954]), .Z(o[2954]) );
  AND U15660 ( .A(p_input[22954]), .B(p_input[12954]), .Z(n7830) );
  AND U15661 ( .A(n7831), .B(p_input[2953]), .Z(o[2953]) );
  AND U15662 ( .A(p_input[22953]), .B(p_input[12953]), .Z(n7831) );
  AND U15663 ( .A(n7832), .B(p_input[2952]), .Z(o[2952]) );
  AND U15664 ( .A(p_input[22952]), .B(p_input[12952]), .Z(n7832) );
  AND U15665 ( .A(n7833), .B(p_input[2951]), .Z(o[2951]) );
  AND U15666 ( .A(p_input[22951]), .B(p_input[12951]), .Z(n7833) );
  AND U15667 ( .A(n7834), .B(p_input[2950]), .Z(o[2950]) );
  AND U15668 ( .A(p_input[22950]), .B(p_input[12950]), .Z(n7834) );
  AND U15669 ( .A(n7835), .B(p_input[294]), .Z(o[294]) );
  AND U15670 ( .A(p_input[20294]), .B(p_input[10294]), .Z(n7835) );
  AND U15671 ( .A(n7836), .B(p_input[2949]), .Z(o[2949]) );
  AND U15672 ( .A(p_input[22949]), .B(p_input[12949]), .Z(n7836) );
  AND U15673 ( .A(n7837), .B(p_input[2948]), .Z(o[2948]) );
  AND U15674 ( .A(p_input[22948]), .B(p_input[12948]), .Z(n7837) );
  AND U15675 ( .A(n7838), .B(p_input[2947]), .Z(o[2947]) );
  AND U15676 ( .A(p_input[22947]), .B(p_input[12947]), .Z(n7838) );
  AND U15677 ( .A(n7839), .B(p_input[2946]), .Z(o[2946]) );
  AND U15678 ( .A(p_input[22946]), .B(p_input[12946]), .Z(n7839) );
  AND U15679 ( .A(n7840), .B(p_input[2945]), .Z(o[2945]) );
  AND U15680 ( .A(p_input[22945]), .B(p_input[12945]), .Z(n7840) );
  AND U15681 ( .A(n7841), .B(p_input[2944]), .Z(o[2944]) );
  AND U15682 ( .A(p_input[22944]), .B(p_input[12944]), .Z(n7841) );
  AND U15683 ( .A(n7842), .B(p_input[2943]), .Z(o[2943]) );
  AND U15684 ( .A(p_input[22943]), .B(p_input[12943]), .Z(n7842) );
  AND U15685 ( .A(n7843), .B(p_input[2942]), .Z(o[2942]) );
  AND U15686 ( .A(p_input[22942]), .B(p_input[12942]), .Z(n7843) );
  AND U15687 ( .A(n7844), .B(p_input[2941]), .Z(o[2941]) );
  AND U15688 ( .A(p_input[22941]), .B(p_input[12941]), .Z(n7844) );
  AND U15689 ( .A(n7845), .B(p_input[2940]), .Z(o[2940]) );
  AND U15690 ( .A(p_input[22940]), .B(p_input[12940]), .Z(n7845) );
  AND U15691 ( .A(n7846), .B(p_input[293]), .Z(o[293]) );
  AND U15692 ( .A(p_input[20293]), .B(p_input[10293]), .Z(n7846) );
  AND U15693 ( .A(n7847), .B(p_input[2939]), .Z(o[2939]) );
  AND U15694 ( .A(p_input[22939]), .B(p_input[12939]), .Z(n7847) );
  AND U15695 ( .A(n7848), .B(p_input[2938]), .Z(o[2938]) );
  AND U15696 ( .A(p_input[22938]), .B(p_input[12938]), .Z(n7848) );
  AND U15697 ( .A(n7849), .B(p_input[2937]), .Z(o[2937]) );
  AND U15698 ( .A(p_input[22937]), .B(p_input[12937]), .Z(n7849) );
  AND U15699 ( .A(n7850), .B(p_input[2936]), .Z(o[2936]) );
  AND U15700 ( .A(p_input[22936]), .B(p_input[12936]), .Z(n7850) );
  AND U15701 ( .A(n7851), .B(p_input[2935]), .Z(o[2935]) );
  AND U15702 ( .A(p_input[22935]), .B(p_input[12935]), .Z(n7851) );
  AND U15703 ( .A(n7852), .B(p_input[2934]), .Z(o[2934]) );
  AND U15704 ( .A(p_input[22934]), .B(p_input[12934]), .Z(n7852) );
  AND U15705 ( .A(n7853), .B(p_input[2933]), .Z(o[2933]) );
  AND U15706 ( .A(p_input[22933]), .B(p_input[12933]), .Z(n7853) );
  AND U15707 ( .A(n7854), .B(p_input[2932]), .Z(o[2932]) );
  AND U15708 ( .A(p_input[22932]), .B(p_input[12932]), .Z(n7854) );
  AND U15709 ( .A(n7855), .B(p_input[2931]), .Z(o[2931]) );
  AND U15710 ( .A(p_input[22931]), .B(p_input[12931]), .Z(n7855) );
  AND U15711 ( .A(n7856), .B(p_input[2930]), .Z(o[2930]) );
  AND U15712 ( .A(p_input[22930]), .B(p_input[12930]), .Z(n7856) );
  AND U15713 ( .A(n7857), .B(p_input[292]), .Z(o[292]) );
  AND U15714 ( .A(p_input[20292]), .B(p_input[10292]), .Z(n7857) );
  AND U15715 ( .A(n7858), .B(p_input[2929]), .Z(o[2929]) );
  AND U15716 ( .A(p_input[22929]), .B(p_input[12929]), .Z(n7858) );
  AND U15717 ( .A(n7859), .B(p_input[2928]), .Z(o[2928]) );
  AND U15718 ( .A(p_input[22928]), .B(p_input[12928]), .Z(n7859) );
  AND U15719 ( .A(n7860), .B(p_input[2927]), .Z(o[2927]) );
  AND U15720 ( .A(p_input[22927]), .B(p_input[12927]), .Z(n7860) );
  AND U15721 ( .A(n7861), .B(p_input[2926]), .Z(o[2926]) );
  AND U15722 ( .A(p_input[22926]), .B(p_input[12926]), .Z(n7861) );
  AND U15723 ( .A(n7862), .B(p_input[2925]), .Z(o[2925]) );
  AND U15724 ( .A(p_input[22925]), .B(p_input[12925]), .Z(n7862) );
  AND U15725 ( .A(n7863), .B(p_input[2924]), .Z(o[2924]) );
  AND U15726 ( .A(p_input[22924]), .B(p_input[12924]), .Z(n7863) );
  AND U15727 ( .A(n7864), .B(p_input[2923]), .Z(o[2923]) );
  AND U15728 ( .A(p_input[22923]), .B(p_input[12923]), .Z(n7864) );
  AND U15729 ( .A(n7865), .B(p_input[2922]), .Z(o[2922]) );
  AND U15730 ( .A(p_input[22922]), .B(p_input[12922]), .Z(n7865) );
  AND U15731 ( .A(n7866), .B(p_input[2921]), .Z(o[2921]) );
  AND U15732 ( .A(p_input[22921]), .B(p_input[12921]), .Z(n7866) );
  AND U15733 ( .A(n7867), .B(p_input[2920]), .Z(o[2920]) );
  AND U15734 ( .A(p_input[22920]), .B(p_input[12920]), .Z(n7867) );
  AND U15735 ( .A(n7868), .B(p_input[291]), .Z(o[291]) );
  AND U15736 ( .A(p_input[20291]), .B(p_input[10291]), .Z(n7868) );
  AND U15737 ( .A(n7869), .B(p_input[2919]), .Z(o[2919]) );
  AND U15738 ( .A(p_input[22919]), .B(p_input[12919]), .Z(n7869) );
  AND U15739 ( .A(n7870), .B(p_input[2918]), .Z(o[2918]) );
  AND U15740 ( .A(p_input[22918]), .B(p_input[12918]), .Z(n7870) );
  AND U15741 ( .A(n7871), .B(p_input[2917]), .Z(o[2917]) );
  AND U15742 ( .A(p_input[22917]), .B(p_input[12917]), .Z(n7871) );
  AND U15743 ( .A(n7872), .B(p_input[2916]), .Z(o[2916]) );
  AND U15744 ( .A(p_input[22916]), .B(p_input[12916]), .Z(n7872) );
  AND U15745 ( .A(n7873), .B(p_input[2915]), .Z(o[2915]) );
  AND U15746 ( .A(p_input[22915]), .B(p_input[12915]), .Z(n7873) );
  AND U15747 ( .A(n7874), .B(p_input[2914]), .Z(o[2914]) );
  AND U15748 ( .A(p_input[22914]), .B(p_input[12914]), .Z(n7874) );
  AND U15749 ( .A(n7875), .B(p_input[2913]), .Z(o[2913]) );
  AND U15750 ( .A(p_input[22913]), .B(p_input[12913]), .Z(n7875) );
  AND U15751 ( .A(n7876), .B(p_input[2912]), .Z(o[2912]) );
  AND U15752 ( .A(p_input[22912]), .B(p_input[12912]), .Z(n7876) );
  AND U15753 ( .A(n7877), .B(p_input[2911]), .Z(o[2911]) );
  AND U15754 ( .A(p_input[22911]), .B(p_input[12911]), .Z(n7877) );
  AND U15755 ( .A(n7878), .B(p_input[2910]), .Z(o[2910]) );
  AND U15756 ( .A(p_input[22910]), .B(p_input[12910]), .Z(n7878) );
  AND U15757 ( .A(n7879), .B(p_input[290]), .Z(o[290]) );
  AND U15758 ( .A(p_input[20290]), .B(p_input[10290]), .Z(n7879) );
  AND U15759 ( .A(n7880), .B(p_input[2909]), .Z(o[2909]) );
  AND U15760 ( .A(p_input[22909]), .B(p_input[12909]), .Z(n7880) );
  AND U15761 ( .A(n7881), .B(p_input[2908]), .Z(o[2908]) );
  AND U15762 ( .A(p_input[22908]), .B(p_input[12908]), .Z(n7881) );
  AND U15763 ( .A(n7882), .B(p_input[2907]), .Z(o[2907]) );
  AND U15764 ( .A(p_input[22907]), .B(p_input[12907]), .Z(n7882) );
  AND U15765 ( .A(n7883), .B(p_input[2906]), .Z(o[2906]) );
  AND U15766 ( .A(p_input[22906]), .B(p_input[12906]), .Z(n7883) );
  AND U15767 ( .A(n7884), .B(p_input[2905]), .Z(o[2905]) );
  AND U15768 ( .A(p_input[22905]), .B(p_input[12905]), .Z(n7884) );
  AND U15769 ( .A(n7885), .B(p_input[2904]), .Z(o[2904]) );
  AND U15770 ( .A(p_input[22904]), .B(p_input[12904]), .Z(n7885) );
  AND U15771 ( .A(n7886), .B(p_input[2903]), .Z(o[2903]) );
  AND U15772 ( .A(p_input[22903]), .B(p_input[12903]), .Z(n7886) );
  AND U15773 ( .A(n7887), .B(p_input[2902]), .Z(o[2902]) );
  AND U15774 ( .A(p_input[22902]), .B(p_input[12902]), .Z(n7887) );
  AND U15775 ( .A(n7888), .B(p_input[2901]), .Z(o[2901]) );
  AND U15776 ( .A(p_input[22901]), .B(p_input[12901]), .Z(n7888) );
  AND U15777 ( .A(n7889), .B(p_input[2900]), .Z(o[2900]) );
  AND U15778 ( .A(p_input[22900]), .B(p_input[12900]), .Z(n7889) );
  AND U15779 ( .A(n7890), .B(p_input[28]), .Z(o[28]) );
  AND U15780 ( .A(p_input[20028]), .B(p_input[10028]), .Z(n7890) );
  AND U15781 ( .A(n7891), .B(p_input[289]), .Z(o[289]) );
  AND U15782 ( .A(p_input[20289]), .B(p_input[10289]), .Z(n7891) );
  AND U15783 ( .A(n7892), .B(p_input[2899]), .Z(o[2899]) );
  AND U15784 ( .A(p_input[22899]), .B(p_input[12899]), .Z(n7892) );
  AND U15785 ( .A(n7893), .B(p_input[2898]), .Z(o[2898]) );
  AND U15786 ( .A(p_input[22898]), .B(p_input[12898]), .Z(n7893) );
  AND U15787 ( .A(n7894), .B(p_input[2897]), .Z(o[2897]) );
  AND U15788 ( .A(p_input[22897]), .B(p_input[12897]), .Z(n7894) );
  AND U15789 ( .A(n7895), .B(p_input[2896]), .Z(o[2896]) );
  AND U15790 ( .A(p_input[22896]), .B(p_input[12896]), .Z(n7895) );
  AND U15791 ( .A(n7896), .B(p_input[2895]), .Z(o[2895]) );
  AND U15792 ( .A(p_input[22895]), .B(p_input[12895]), .Z(n7896) );
  AND U15793 ( .A(n7897), .B(p_input[2894]), .Z(o[2894]) );
  AND U15794 ( .A(p_input[22894]), .B(p_input[12894]), .Z(n7897) );
  AND U15795 ( .A(n7898), .B(p_input[2893]), .Z(o[2893]) );
  AND U15796 ( .A(p_input[22893]), .B(p_input[12893]), .Z(n7898) );
  AND U15797 ( .A(n7899), .B(p_input[2892]), .Z(o[2892]) );
  AND U15798 ( .A(p_input[22892]), .B(p_input[12892]), .Z(n7899) );
  AND U15799 ( .A(n7900), .B(p_input[2891]), .Z(o[2891]) );
  AND U15800 ( .A(p_input[22891]), .B(p_input[12891]), .Z(n7900) );
  AND U15801 ( .A(n7901), .B(p_input[2890]), .Z(o[2890]) );
  AND U15802 ( .A(p_input[22890]), .B(p_input[12890]), .Z(n7901) );
  AND U15803 ( .A(n7902), .B(p_input[288]), .Z(o[288]) );
  AND U15804 ( .A(p_input[20288]), .B(p_input[10288]), .Z(n7902) );
  AND U15805 ( .A(n7903), .B(p_input[2889]), .Z(o[2889]) );
  AND U15806 ( .A(p_input[22889]), .B(p_input[12889]), .Z(n7903) );
  AND U15807 ( .A(n7904), .B(p_input[2888]), .Z(o[2888]) );
  AND U15808 ( .A(p_input[22888]), .B(p_input[12888]), .Z(n7904) );
  AND U15809 ( .A(n7905), .B(p_input[2887]), .Z(o[2887]) );
  AND U15810 ( .A(p_input[22887]), .B(p_input[12887]), .Z(n7905) );
  AND U15811 ( .A(n7906), .B(p_input[2886]), .Z(o[2886]) );
  AND U15812 ( .A(p_input[22886]), .B(p_input[12886]), .Z(n7906) );
  AND U15813 ( .A(n7907), .B(p_input[2885]), .Z(o[2885]) );
  AND U15814 ( .A(p_input[22885]), .B(p_input[12885]), .Z(n7907) );
  AND U15815 ( .A(n7908), .B(p_input[2884]), .Z(o[2884]) );
  AND U15816 ( .A(p_input[22884]), .B(p_input[12884]), .Z(n7908) );
  AND U15817 ( .A(n7909), .B(p_input[2883]), .Z(o[2883]) );
  AND U15818 ( .A(p_input[22883]), .B(p_input[12883]), .Z(n7909) );
  AND U15819 ( .A(n7910), .B(p_input[2882]), .Z(o[2882]) );
  AND U15820 ( .A(p_input[22882]), .B(p_input[12882]), .Z(n7910) );
  AND U15821 ( .A(n7911), .B(p_input[2881]), .Z(o[2881]) );
  AND U15822 ( .A(p_input[22881]), .B(p_input[12881]), .Z(n7911) );
  AND U15823 ( .A(n7912), .B(p_input[2880]), .Z(o[2880]) );
  AND U15824 ( .A(p_input[22880]), .B(p_input[12880]), .Z(n7912) );
  AND U15825 ( .A(n7913), .B(p_input[287]), .Z(o[287]) );
  AND U15826 ( .A(p_input[20287]), .B(p_input[10287]), .Z(n7913) );
  AND U15827 ( .A(n7914), .B(p_input[2879]), .Z(o[2879]) );
  AND U15828 ( .A(p_input[22879]), .B(p_input[12879]), .Z(n7914) );
  AND U15829 ( .A(n7915), .B(p_input[2878]), .Z(o[2878]) );
  AND U15830 ( .A(p_input[22878]), .B(p_input[12878]), .Z(n7915) );
  AND U15831 ( .A(n7916), .B(p_input[2877]), .Z(o[2877]) );
  AND U15832 ( .A(p_input[22877]), .B(p_input[12877]), .Z(n7916) );
  AND U15833 ( .A(n7917), .B(p_input[2876]), .Z(o[2876]) );
  AND U15834 ( .A(p_input[22876]), .B(p_input[12876]), .Z(n7917) );
  AND U15835 ( .A(n7918), .B(p_input[2875]), .Z(o[2875]) );
  AND U15836 ( .A(p_input[22875]), .B(p_input[12875]), .Z(n7918) );
  AND U15837 ( .A(n7919), .B(p_input[2874]), .Z(o[2874]) );
  AND U15838 ( .A(p_input[22874]), .B(p_input[12874]), .Z(n7919) );
  AND U15839 ( .A(n7920), .B(p_input[2873]), .Z(o[2873]) );
  AND U15840 ( .A(p_input[22873]), .B(p_input[12873]), .Z(n7920) );
  AND U15841 ( .A(n7921), .B(p_input[2872]), .Z(o[2872]) );
  AND U15842 ( .A(p_input[22872]), .B(p_input[12872]), .Z(n7921) );
  AND U15843 ( .A(n7922), .B(p_input[2871]), .Z(o[2871]) );
  AND U15844 ( .A(p_input[22871]), .B(p_input[12871]), .Z(n7922) );
  AND U15845 ( .A(n7923), .B(p_input[2870]), .Z(o[2870]) );
  AND U15846 ( .A(p_input[22870]), .B(p_input[12870]), .Z(n7923) );
  AND U15847 ( .A(n7924), .B(p_input[286]), .Z(o[286]) );
  AND U15848 ( .A(p_input[20286]), .B(p_input[10286]), .Z(n7924) );
  AND U15849 ( .A(n7925), .B(p_input[2869]), .Z(o[2869]) );
  AND U15850 ( .A(p_input[22869]), .B(p_input[12869]), .Z(n7925) );
  AND U15851 ( .A(n7926), .B(p_input[2868]), .Z(o[2868]) );
  AND U15852 ( .A(p_input[22868]), .B(p_input[12868]), .Z(n7926) );
  AND U15853 ( .A(n7927), .B(p_input[2867]), .Z(o[2867]) );
  AND U15854 ( .A(p_input[22867]), .B(p_input[12867]), .Z(n7927) );
  AND U15855 ( .A(n7928), .B(p_input[2866]), .Z(o[2866]) );
  AND U15856 ( .A(p_input[22866]), .B(p_input[12866]), .Z(n7928) );
  AND U15857 ( .A(n7929), .B(p_input[2865]), .Z(o[2865]) );
  AND U15858 ( .A(p_input[22865]), .B(p_input[12865]), .Z(n7929) );
  AND U15859 ( .A(n7930), .B(p_input[2864]), .Z(o[2864]) );
  AND U15860 ( .A(p_input[22864]), .B(p_input[12864]), .Z(n7930) );
  AND U15861 ( .A(n7931), .B(p_input[2863]), .Z(o[2863]) );
  AND U15862 ( .A(p_input[22863]), .B(p_input[12863]), .Z(n7931) );
  AND U15863 ( .A(n7932), .B(p_input[2862]), .Z(o[2862]) );
  AND U15864 ( .A(p_input[22862]), .B(p_input[12862]), .Z(n7932) );
  AND U15865 ( .A(n7933), .B(p_input[2861]), .Z(o[2861]) );
  AND U15866 ( .A(p_input[22861]), .B(p_input[12861]), .Z(n7933) );
  AND U15867 ( .A(n7934), .B(p_input[2860]), .Z(o[2860]) );
  AND U15868 ( .A(p_input[22860]), .B(p_input[12860]), .Z(n7934) );
  AND U15869 ( .A(n7935), .B(p_input[285]), .Z(o[285]) );
  AND U15870 ( .A(p_input[20285]), .B(p_input[10285]), .Z(n7935) );
  AND U15871 ( .A(n7936), .B(p_input[2859]), .Z(o[2859]) );
  AND U15872 ( .A(p_input[22859]), .B(p_input[12859]), .Z(n7936) );
  AND U15873 ( .A(n7937), .B(p_input[2858]), .Z(o[2858]) );
  AND U15874 ( .A(p_input[22858]), .B(p_input[12858]), .Z(n7937) );
  AND U15875 ( .A(n7938), .B(p_input[2857]), .Z(o[2857]) );
  AND U15876 ( .A(p_input[22857]), .B(p_input[12857]), .Z(n7938) );
  AND U15877 ( .A(n7939), .B(p_input[2856]), .Z(o[2856]) );
  AND U15878 ( .A(p_input[22856]), .B(p_input[12856]), .Z(n7939) );
  AND U15879 ( .A(n7940), .B(p_input[2855]), .Z(o[2855]) );
  AND U15880 ( .A(p_input[22855]), .B(p_input[12855]), .Z(n7940) );
  AND U15881 ( .A(n7941), .B(p_input[2854]), .Z(o[2854]) );
  AND U15882 ( .A(p_input[22854]), .B(p_input[12854]), .Z(n7941) );
  AND U15883 ( .A(n7942), .B(p_input[2853]), .Z(o[2853]) );
  AND U15884 ( .A(p_input[22853]), .B(p_input[12853]), .Z(n7942) );
  AND U15885 ( .A(n7943), .B(p_input[2852]), .Z(o[2852]) );
  AND U15886 ( .A(p_input[22852]), .B(p_input[12852]), .Z(n7943) );
  AND U15887 ( .A(n7944), .B(p_input[2851]), .Z(o[2851]) );
  AND U15888 ( .A(p_input[22851]), .B(p_input[12851]), .Z(n7944) );
  AND U15889 ( .A(n7945), .B(p_input[2850]), .Z(o[2850]) );
  AND U15890 ( .A(p_input[22850]), .B(p_input[12850]), .Z(n7945) );
  AND U15891 ( .A(n7946), .B(p_input[284]), .Z(o[284]) );
  AND U15892 ( .A(p_input[20284]), .B(p_input[10284]), .Z(n7946) );
  AND U15893 ( .A(n7947), .B(p_input[2849]), .Z(o[2849]) );
  AND U15894 ( .A(p_input[22849]), .B(p_input[12849]), .Z(n7947) );
  AND U15895 ( .A(n7948), .B(p_input[2848]), .Z(o[2848]) );
  AND U15896 ( .A(p_input[22848]), .B(p_input[12848]), .Z(n7948) );
  AND U15897 ( .A(n7949), .B(p_input[2847]), .Z(o[2847]) );
  AND U15898 ( .A(p_input[22847]), .B(p_input[12847]), .Z(n7949) );
  AND U15899 ( .A(n7950), .B(p_input[2846]), .Z(o[2846]) );
  AND U15900 ( .A(p_input[22846]), .B(p_input[12846]), .Z(n7950) );
  AND U15901 ( .A(n7951), .B(p_input[2845]), .Z(o[2845]) );
  AND U15902 ( .A(p_input[22845]), .B(p_input[12845]), .Z(n7951) );
  AND U15903 ( .A(n7952), .B(p_input[2844]), .Z(o[2844]) );
  AND U15904 ( .A(p_input[22844]), .B(p_input[12844]), .Z(n7952) );
  AND U15905 ( .A(n7953), .B(p_input[2843]), .Z(o[2843]) );
  AND U15906 ( .A(p_input[22843]), .B(p_input[12843]), .Z(n7953) );
  AND U15907 ( .A(n7954), .B(p_input[2842]), .Z(o[2842]) );
  AND U15908 ( .A(p_input[22842]), .B(p_input[12842]), .Z(n7954) );
  AND U15909 ( .A(n7955), .B(p_input[2841]), .Z(o[2841]) );
  AND U15910 ( .A(p_input[22841]), .B(p_input[12841]), .Z(n7955) );
  AND U15911 ( .A(n7956), .B(p_input[2840]), .Z(o[2840]) );
  AND U15912 ( .A(p_input[22840]), .B(p_input[12840]), .Z(n7956) );
  AND U15913 ( .A(n7957), .B(p_input[283]), .Z(o[283]) );
  AND U15914 ( .A(p_input[20283]), .B(p_input[10283]), .Z(n7957) );
  AND U15915 ( .A(n7958), .B(p_input[2839]), .Z(o[2839]) );
  AND U15916 ( .A(p_input[22839]), .B(p_input[12839]), .Z(n7958) );
  AND U15917 ( .A(n7959), .B(p_input[2838]), .Z(o[2838]) );
  AND U15918 ( .A(p_input[22838]), .B(p_input[12838]), .Z(n7959) );
  AND U15919 ( .A(n7960), .B(p_input[2837]), .Z(o[2837]) );
  AND U15920 ( .A(p_input[22837]), .B(p_input[12837]), .Z(n7960) );
  AND U15921 ( .A(n7961), .B(p_input[2836]), .Z(o[2836]) );
  AND U15922 ( .A(p_input[22836]), .B(p_input[12836]), .Z(n7961) );
  AND U15923 ( .A(n7962), .B(p_input[2835]), .Z(o[2835]) );
  AND U15924 ( .A(p_input[22835]), .B(p_input[12835]), .Z(n7962) );
  AND U15925 ( .A(n7963), .B(p_input[2834]), .Z(o[2834]) );
  AND U15926 ( .A(p_input[22834]), .B(p_input[12834]), .Z(n7963) );
  AND U15927 ( .A(n7964), .B(p_input[2833]), .Z(o[2833]) );
  AND U15928 ( .A(p_input[22833]), .B(p_input[12833]), .Z(n7964) );
  AND U15929 ( .A(n7965), .B(p_input[2832]), .Z(o[2832]) );
  AND U15930 ( .A(p_input[22832]), .B(p_input[12832]), .Z(n7965) );
  AND U15931 ( .A(n7966), .B(p_input[2831]), .Z(o[2831]) );
  AND U15932 ( .A(p_input[22831]), .B(p_input[12831]), .Z(n7966) );
  AND U15933 ( .A(n7967), .B(p_input[2830]), .Z(o[2830]) );
  AND U15934 ( .A(p_input[22830]), .B(p_input[12830]), .Z(n7967) );
  AND U15935 ( .A(n7968), .B(p_input[282]), .Z(o[282]) );
  AND U15936 ( .A(p_input[20282]), .B(p_input[10282]), .Z(n7968) );
  AND U15937 ( .A(n7969), .B(p_input[2829]), .Z(o[2829]) );
  AND U15938 ( .A(p_input[22829]), .B(p_input[12829]), .Z(n7969) );
  AND U15939 ( .A(n7970), .B(p_input[2828]), .Z(o[2828]) );
  AND U15940 ( .A(p_input[22828]), .B(p_input[12828]), .Z(n7970) );
  AND U15941 ( .A(n7971), .B(p_input[2827]), .Z(o[2827]) );
  AND U15942 ( .A(p_input[22827]), .B(p_input[12827]), .Z(n7971) );
  AND U15943 ( .A(n7972), .B(p_input[2826]), .Z(o[2826]) );
  AND U15944 ( .A(p_input[22826]), .B(p_input[12826]), .Z(n7972) );
  AND U15945 ( .A(n7973), .B(p_input[2825]), .Z(o[2825]) );
  AND U15946 ( .A(p_input[22825]), .B(p_input[12825]), .Z(n7973) );
  AND U15947 ( .A(n7974), .B(p_input[2824]), .Z(o[2824]) );
  AND U15948 ( .A(p_input[22824]), .B(p_input[12824]), .Z(n7974) );
  AND U15949 ( .A(n7975), .B(p_input[2823]), .Z(o[2823]) );
  AND U15950 ( .A(p_input[22823]), .B(p_input[12823]), .Z(n7975) );
  AND U15951 ( .A(n7976), .B(p_input[2822]), .Z(o[2822]) );
  AND U15952 ( .A(p_input[22822]), .B(p_input[12822]), .Z(n7976) );
  AND U15953 ( .A(n7977), .B(p_input[2821]), .Z(o[2821]) );
  AND U15954 ( .A(p_input[22821]), .B(p_input[12821]), .Z(n7977) );
  AND U15955 ( .A(n7978), .B(p_input[2820]), .Z(o[2820]) );
  AND U15956 ( .A(p_input[22820]), .B(p_input[12820]), .Z(n7978) );
  AND U15957 ( .A(n7979), .B(p_input[281]), .Z(o[281]) );
  AND U15958 ( .A(p_input[20281]), .B(p_input[10281]), .Z(n7979) );
  AND U15959 ( .A(n7980), .B(p_input[2819]), .Z(o[2819]) );
  AND U15960 ( .A(p_input[22819]), .B(p_input[12819]), .Z(n7980) );
  AND U15961 ( .A(n7981), .B(p_input[2818]), .Z(o[2818]) );
  AND U15962 ( .A(p_input[22818]), .B(p_input[12818]), .Z(n7981) );
  AND U15963 ( .A(n7982), .B(p_input[2817]), .Z(o[2817]) );
  AND U15964 ( .A(p_input[22817]), .B(p_input[12817]), .Z(n7982) );
  AND U15965 ( .A(n7983), .B(p_input[2816]), .Z(o[2816]) );
  AND U15966 ( .A(p_input[22816]), .B(p_input[12816]), .Z(n7983) );
  AND U15967 ( .A(n7984), .B(p_input[2815]), .Z(o[2815]) );
  AND U15968 ( .A(p_input[22815]), .B(p_input[12815]), .Z(n7984) );
  AND U15969 ( .A(n7985), .B(p_input[2814]), .Z(o[2814]) );
  AND U15970 ( .A(p_input[22814]), .B(p_input[12814]), .Z(n7985) );
  AND U15971 ( .A(n7986), .B(p_input[2813]), .Z(o[2813]) );
  AND U15972 ( .A(p_input[22813]), .B(p_input[12813]), .Z(n7986) );
  AND U15973 ( .A(n7987), .B(p_input[2812]), .Z(o[2812]) );
  AND U15974 ( .A(p_input[22812]), .B(p_input[12812]), .Z(n7987) );
  AND U15975 ( .A(n7988), .B(p_input[2811]), .Z(o[2811]) );
  AND U15976 ( .A(p_input[22811]), .B(p_input[12811]), .Z(n7988) );
  AND U15977 ( .A(n7989), .B(p_input[2810]), .Z(o[2810]) );
  AND U15978 ( .A(p_input[22810]), .B(p_input[12810]), .Z(n7989) );
  AND U15979 ( .A(n7990), .B(p_input[280]), .Z(o[280]) );
  AND U15980 ( .A(p_input[20280]), .B(p_input[10280]), .Z(n7990) );
  AND U15981 ( .A(n7991), .B(p_input[2809]), .Z(o[2809]) );
  AND U15982 ( .A(p_input[22809]), .B(p_input[12809]), .Z(n7991) );
  AND U15983 ( .A(n7992), .B(p_input[2808]), .Z(o[2808]) );
  AND U15984 ( .A(p_input[22808]), .B(p_input[12808]), .Z(n7992) );
  AND U15985 ( .A(n7993), .B(p_input[2807]), .Z(o[2807]) );
  AND U15986 ( .A(p_input[22807]), .B(p_input[12807]), .Z(n7993) );
  AND U15987 ( .A(n7994), .B(p_input[2806]), .Z(o[2806]) );
  AND U15988 ( .A(p_input[22806]), .B(p_input[12806]), .Z(n7994) );
  AND U15989 ( .A(n7995), .B(p_input[2805]), .Z(o[2805]) );
  AND U15990 ( .A(p_input[22805]), .B(p_input[12805]), .Z(n7995) );
  AND U15991 ( .A(n7996), .B(p_input[2804]), .Z(o[2804]) );
  AND U15992 ( .A(p_input[22804]), .B(p_input[12804]), .Z(n7996) );
  AND U15993 ( .A(n7997), .B(p_input[2803]), .Z(o[2803]) );
  AND U15994 ( .A(p_input[22803]), .B(p_input[12803]), .Z(n7997) );
  AND U15995 ( .A(n7998), .B(p_input[2802]), .Z(o[2802]) );
  AND U15996 ( .A(p_input[22802]), .B(p_input[12802]), .Z(n7998) );
  AND U15997 ( .A(n7999), .B(p_input[2801]), .Z(o[2801]) );
  AND U15998 ( .A(p_input[22801]), .B(p_input[12801]), .Z(n7999) );
  AND U15999 ( .A(n8000), .B(p_input[2800]), .Z(o[2800]) );
  AND U16000 ( .A(p_input[22800]), .B(p_input[12800]), .Z(n8000) );
  AND U16001 ( .A(n8001), .B(p_input[27]), .Z(o[27]) );
  AND U16002 ( .A(p_input[20027]), .B(p_input[10027]), .Z(n8001) );
  AND U16003 ( .A(n8002), .B(p_input[279]), .Z(o[279]) );
  AND U16004 ( .A(p_input[20279]), .B(p_input[10279]), .Z(n8002) );
  AND U16005 ( .A(n8003), .B(p_input[2799]), .Z(o[2799]) );
  AND U16006 ( .A(p_input[22799]), .B(p_input[12799]), .Z(n8003) );
  AND U16007 ( .A(n8004), .B(p_input[2798]), .Z(o[2798]) );
  AND U16008 ( .A(p_input[22798]), .B(p_input[12798]), .Z(n8004) );
  AND U16009 ( .A(n8005), .B(p_input[2797]), .Z(o[2797]) );
  AND U16010 ( .A(p_input[22797]), .B(p_input[12797]), .Z(n8005) );
  AND U16011 ( .A(n8006), .B(p_input[2796]), .Z(o[2796]) );
  AND U16012 ( .A(p_input[22796]), .B(p_input[12796]), .Z(n8006) );
  AND U16013 ( .A(n8007), .B(p_input[2795]), .Z(o[2795]) );
  AND U16014 ( .A(p_input[22795]), .B(p_input[12795]), .Z(n8007) );
  AND U16015 ( .A(n8008), .B(p_input[2794]), .Z(o[2794]) );
  AND U16016 ( .A(p_input[22794]), .B(p_input[12794]), .Z(n8008) );
  AND U16017 ( .A(n8009), .B(p_input[2793]), .Z(o[2793]) );
  AND U16018 ( .A(p_input[22793]), .B(p_input[12793]), .Z(n8009) );
  AND U16019 ( .A(n8010), .B(p_input[2792]), .Z(o[2792]) );
  AND U16020 ( .A(p_input[22792]), .B(p_input[12792]), .Z(n8010) );
  AND U16021 ( .A(n8011), .B(p_input[2791]), .Z(o[2791]) );
  AND U16022 ( .A(p_input[22791]), .B(p_input[12791]), .Z(n8011) );
  AND U16023 ( .A(n8012), .B(p_input[2790]), .Z(o[2790]) );
  AND U16024 ( .A(p_input[22790]), .B(p_input[12790]), .Z(n8012) );
  AND U16025 ( .A(n8013), .B(p_input[278]), .Z(o[278]) );
  AND U16026 ( .A(p_input[20278]), .B(p_input[10278]), .Z(n8013) );
  AND U16027 ( .A(n8014), .B(p_input[2789]), .Z(o[2789]) );
  AND U16028 ( .A(p_input[22789]), .B(p_input[12789]), .Z(n8014) );
  AND U16029 ( .A(n8015), .B(p_input[2788]), .Z(o[2788]) );
  AND U16030 ( .A(p_input[22788]), .B(p_input[12788]), .Z(n8015) );
  AND U16031 ( .A(n8016), .B(p_input[2787]), .Z(o[2787]) );
  AND U16032 ( .A(p_input[22787]), .B(p_input[12787]), .Z(n8016) );
  AND U16033 ( .A(n8017), .B(p_input[2786]), .Z(o[2786]) );
  AND U16034 ( .A(p_input[22786]), .B(p_input[12786]), .Z(n8017) );
  AND U16035 ( .A(n8018), .B(p_input[2785]), .Z(o[2785]) );
  AND U16036 ( .A(p_input[22785]), .B(p_input[12785]), .Z(n8018) );
  AND U16037 ( .A(n8019), .B(p_input[2784]), .Z(o[2784]) );
  AND U16038 ( .A(p_input[22784]), .B(p_input[12784]), .Z(n8019) );
  AND U16039 ( .A(n8020), .B(p_input[2783]), .Z(o[2783]) );
  AND U16040 ( .A(p_input[22783]), .B(p_input[12783]), .Z(n8020) );
  AND U16041 ( .A(n8021), .B(p_input[2782]), .Z(o[2782]) );
  AND U16042 ( .A(p_input[22782]), .B(p_input[12782]), .Z(n8021) );
  AND U16043 ( .A(n8022), .B(p_input[2781]), .Z(o[2781]) );
  AND U16044 ( .A(p_input[22781]), .B(p_input[12781]), .Z(n8022) );
  AND U16045 ( .A(n8023), .B(p_input[2780]), .Z(o[2780]) );
  AND U16046 ( .A(p_input[22780]), .B(p_input[12780]), .Z(n8023) );
  AND U16047 ( .A(n8024), .B(p_input[277]), .Z(o[277]) );
  AND U16048 ( .A(p_input[20277]), .B(p_input[10277]), .Z(n8024) );
  AND U16049 ( .A(n8025), .B(p_input[2779]), .Z(o[2779]) );
  AND U16050 ( .A(p_input[22779]), .B(p_input[12779]), .Z(n8025) );
  AND U16051 ( .A(n8026), .B(p_input[2778]), .Z(o[2778]) );
  AND U16052 ( .A(p_input[22778]), .B(p_input[12778]), .Z(n8026) );
  AND U16053 ( .A(n8027), .B(p_input[2777]), .Z(o[2777]) );
  AND U16054 ( .A(p_input[22777]), .B(p_input[12777]), .Z(n8027) );
  AND U16055 ( .A(n8028), .B(p_input[2776]), .Z(o[2776]) );
  AND U16056 ( .A(p_input[22776]), .B(p_input[12776]), .Z(n8028) );
  AND U16057 ( .A(n8029), .B(p_input[2775]), .Z(o[2775]) );
  AND U16058 ( .A(p_input[22775]), .B(p_input[12775]), .Z(n8029) );
  AND U16059 ( .A(n8030), .B(p_input[2774]), .Z(o[2774]) );
  AND U16060 ( .A(p_input[22774]), .B(p_input[12774]), .Z(n8030) );
  AND U16061 ( .A(n8031), .B(p_input[2773]), .Z(o[2773]) );
  AND U16062 ( .A(p_input[22773]), .B(p_input[12773]), .Z(n8031) );
  AND U16063 ( .A(n8032), .B(p_input[2772]), .Z(o[2772]) );
  AND U16064 ( .A(p_input[22772]), .B(p_input[12772]), .Z(n8032) );
  AND U16065 ( .A(n8033), .B(p_input[2771]), .Z(o[2771]) );
  AND U16066 ( .A(p_input[22771]), .B(p_input[12771]), .Z(n8033) );
  AND U16067 ( .A(n8034), .B(p_input[2770]), .Z(o[2770]) );
  AND U16068 ( .A(p_input[22770]), .B(p_input[12770]), .Z(n8034) );
  AND U16069 ( .A(n8035), .B(p_input[276]), .Z(o[276]) );
  AND U16070 ( .A(p_input[20276]), .B(p_input[10276]), .Z(n8035) );
  AND U16071 ( .A(n8036), .B(p_input[2769]), .Z(o[2769]) );
  AND U16072 ( .A(p_input[22769]), .B(p_input[12769]), .Z(n8036) );
  AND U16073 ( .A(n8037), .B(p_input[2768]), .Z(o[2768]) );
  AND U16074 ( .A(p_input[22768]), .B(p_input[12768]), .Z(n8037) );
  AND U16075 ( .A(n8038), .B(p_input[2767]), .Z(o[2767]) );
  AND U16076 ( .A(p_input[22767]), .B(p_input[12767]), .Z(n8038) );
  AND U16077 ( .A(n8039), .B(p_input[2766]), .Z(o[2766]) );
  AND U16078 ( .A(p_input[22766]), .B(p_input[12766]), .Z(n8039) );
  AND U16079 ( .A(n8040), .B(p_input[2765]), .Z(o[2765]) );
  AND U16080 ( .A(p_input[22765]), .B(p_input[12765]), .Z(n8040) );
  AND U16081 ( .A(n8041), .B(p_input[2764]), .Z(o[2764]) );
  AND U16082 ( .A(p_input[22764]), .B(p_input[12764]), .Z(n8041) );
  AND U16083 ( .A(n8042), .B(p_input[2763]), .Z(o[2763]) );
  AND U16084 ( .A(p_input[22763]), .B(p_input[12763]), .Z(n8042) );
  AND U16085 ( .A(n8043), .B(p_input[2762]), .Z(o[2762]) );
  AND U16086 ( .A(p_input[22762]), .B(p_input[12762]), .Z(n8043) );
  AND U16087 ( .A(n8044), .B(p_input[2761]), .Z(o[2761]) );
  AND U16088 ( .A(p_input[22761]), .B(p_input[12761]), .Z(n8044) );
  AND U16089 ( .A(n8045), .B(p_input[2760]), .Z(o[2760]) );
  AND U16090 ( .A(p_input[22760]), .B(p_input[12760]), .Z(n8045) );
  AND U16091 ( .A(n8046), .B(p_input[275]), .Z(o[275]) );
  AND U16092 ( .A(p_input[20275]), .B(p_input[10275]), .Z(n8046) );
  AND U16093 ( .A(n8047), .B(p_input[2759]), .Z(o[2759]) );
  AND U16094 ( .A(p_input[22759]), .B(p_input[12759]), .Z(n8047) );
  AND U16095 ( .A(n8048), .B(p_input[2758]), .Z(o[2758]) );
  AND U16096 ( .A(p_input[22758]), .B(p_input[12758]), .Z(n8048) );
  AND U16097 ( .A(n8049), .B(p_input[2757]), .Z(o[2757]) );
  AND U16098 ( .A(p_input[22757]), .B(p_input[12757]), .Z(n8049) );
  AND U16099 ( .A(n8050), .B(p_input[2756]), .Z(o[2756]) );
  AND U16100 ( .A(p_input[22756]), .B(p_input[12756]), .Z(n8050) );
  AND U16101 ( .A(n8051), .B(p_input[2755]), .Z(o[2755]) );
  AND U16102 ( .A(p_input[22755]), .B(p_input[12755]), .Z(n8051) );
  AND U16103 ( .A(n8052), .B(p_input[2754]), .Z(o[2754]) );
  AND U16104 ( .A(p_input[22754]), .B(p_input[12754]), .Z(n8052) );
  AND U16105 ( .A(n8053), .B(p_input[2753]), .Z(o[2753]) );
  AND U16106 ( .A(p_input[22753]), .B(p_input[12753]), .Z(n8053) );
  AND U16107 ( .A(n8054), .B(p_input[2752]), .Z(o[2752]) );
  AND U16108 ( .A(p_input[22752]), .B(p_input[12752]), .Z(n8054) );
  AND U16109 ( .A(n8055), .B(p_input[2751]), .Z(o[2751]) );
  AND U16110 ( .A(p_input[22751]), .B(p_input[12751]), .Z(n8055) );
  AND U16111 ( .A(n8056), .B(p_input[2750]), .Z(o[2750]) );
  AND U16112 ( .A(p_input[22750]), .B(p_input[12750]), .Z(n8056) );
  AND U16113 ( .A(n8057), .B(p_input[274]), .Z(o[274]) );
  AND U16114 ( .A(p_input[20274]), .B(p_input[10274]), .Z(n8057) );
  AND U16115 ( .A(n8058), .B(p_input[2749]), .Z(o[2749]) );
  AND U16116 ( .A(p_input[22749]), .B(p_input[12749]), .Z(n8058) );
  AND U16117 ( .A(n8059), .B(p_input[2748]), .Z(o[2748]) );
  AND U16118 ( .A(p_input[22748]), .B(p_input[12748]), .Z(n8059) );
  AND U16119 ( .A(n8060), .B(p_input[2747]), .Z(o[2747]) );
  AND U16120 ( .A(p_input[22747]), .B(p_input[12747]), .Z(n8060) );
  AND U16121 ( .A(n8061), .B(p_input[2746]), .Z(o[2746]) );
  AND U16122 ( .A(p_input[22746]), .B(p_input[12746]), .Z(n8061) );
  AND U16123 ( .A(n8062), .B(p_input[2745]), .Z(o[2745]) );
  AND U16124 ( .A(p_input[22745]), .B(p_input[12745]), .Z(n8062) );
  AND U16125 ( .A(n8063), .B(p_input[2744]), .Z(o[2744]) );
  AND U16126 ( .A(p_input[22744]), .B(p_input[12744]), .Z(n8063) );
  AND U16127 ( .A(n8064), .B(p_input[2743]), .Z(o[2743]) );
  AND U16128 ( .A(p_input[22743]), .B(p_input[12743]), .Z(n8064) );
  AND U16129 ( .A(n8065), .B(p_input[2742]), .Z(o[2742]) );
  AND U16130 ( .A(p_input[22742]), .B(p_input[12742]), .Z(n8065) );
  AND U16131 ( .A(n8066), .B(p_input[2741]), .Z(o[2741]) );
  AND U16132 ( .A(p_input[22741]), .B(p_input[12741]), .Z(n8066) );
  AND U16133 ( .A(n8067), .B(p_input[2740]), .Z(o[2740]) );
  AND U16134 ( .A(p_input[22740]), .B(p_input[12740]), .Z(n8067) );
  AND U16135 ( .A(n8068), .B(p_input[273]), .Z(o[273]) );
  AND U16136 ( .A(p_input[20273]), .B(p_input[10273]), .Z(n8068) );
  AND U16137 ( .A(n8069), .B(p_input[2739]), .Z(o[2739]) );
  AND U16138 ( .A(p_input[22739]), .B(p_input[12739]), .Z(n8069) );
  AND U16139 ( .A(n8070), .B(p_input[2738]), .Z(o[2738]) );
  AND U16140 ( .A(p_input[22738]), .B(p_input[12738]), .Z(n8070) );
  AND U16141 ( .A(n8071), .B(p_input[2737]), .Z(o[2737]) );
  AND U16142 ( .A(p_input[22737]), .B(p_input[12737]), .Z(n8071) );
  AND U16143 ( .A(n8072), .B(p_input[2736]), .Z(o[2736]) );
  AND U16144 ( .A(p_input[22736]), .B(p_input[12736]), .Z(n8072) );
  AND U16145 ( .A(n8073), .B(p_input[2735]), .Z(o[2735]) );
  AND U16146 ( .A(p_input[22735]), .B(p_input[12735]), .Z(n8073) );
  AND U16147 ( .A(n8074), .B(p_input[2734]), .Z(o[2734]) );
  AND U16148 ( .A(p_input[22734]), .B(p_input[12734]), .Z(n8074) );
  AND U16149 ( .A(n8075), .B(p_input[2733]), .Z(o[2733]) );
  AND U16150 ( .A(p_input[22733]), .B(p_input[12733]), .Z(n8075) );
  AND U16151 ( .A(n8076), .B(p_input[2732]), .Z(o[2732]) );
  AND U16152 ( .A(p_input[22732]), .B(p_input[12732]), .Z(n8076) );
  AND U16153 ( .A(n8077), .B(p_input[2731]), .Z(o[2731]) );
  AND U16154 ( .A(p_input[22731]), .B(p_input[12731]), .Z(n8077) );
  AND U16155 ( .A(n8078), .B(p_input[2730]), .Z(o[2730]) );
  AND U16156 ( .A(p_input[22730]), .B(p_input[12730]), .Z(n8078) );
  AND U16157 ( .A(n8079), .B(p_input[272]), .Z(o[272]) );
  AND U16158 ( .A(p_input[20272]), .B(p_input[10272]), .Z(n8079) );
  AND U16159 ( .A(n8080), .B(p_input[2729]), .Z(o[2729]) );
  AND U16160 ( .A(p_input[22729]), .B(p_input[12729]), .Z(n8080) );
  AND U16161 ( .A(n8081), .B(p_input[2728]), .Z(o[2728]) );
  AND U16162 ( .A(p_input[22728]), .B(p_input[12728]), .Z(n8081) );
  AND U16163 ( .A(n8082), .B(p_input[2727]), .Z(o[2727]) );
  AND U16164 ( .A(p_input[22727]), .B(p_input[12727]), .Z(n8082) );
  AND U16165 ( .A(n8083), .B(p_input[2726]), .Z(o[2726]) );
  AND U16166 ( .A(p_input[22726]), .B(p_input[12726]), .Z(n8083) );
  AND U16167 ( .A(n8084), .B(p_input[2725]), .Z(o[2725]) );
  AND U16168 ( .A(p_input[22725]), .B(p_input[12725]), .Z(n8084) );
  AND U16169 ( .A(n8085), .B(p_input[2724]), .Z(o[2724]) );
  AND U16170 ( .A(p_input[22724]), .B(p_input[12724]), .Z(n8085) );
  AND U16171 ( .A(n8086), .B(p_input[2723]), .Z(o[2723]) );
  AND U16172 ( .A(p_input[22723]), .B(p_input[12723]), .Z(n8086) );
  AND U16173 ( .A(n8087), .B(p_input[2722]), .Z(o[2722]) );
  AND U16174 ( .A(p_input[22722]), .B(p_input[12722]), .Z(n8087) );
  AND U16175 ( .A(n8088), .B(p_input[2721]), .Z(o[2721]) );
  AND U16176 ( .A(p_input[22721]), .B(p_input[12721]), .Z(n8088) );
  AND U16177 ( .A(n8089), .B(p_input[2720]), .Z(o[2720]) );
  AND U16178 ( .A(p_input[22720]), .B(p_input[12720]), .Z(n8089) );
  AND U16179 ( .A(n8090), .B(p_input[271]), .Z(o[271]) );
  AND U16180 ( .A(p_input[20271]), .B(p_input[10271]), .Z(n8090) );
  AND U16181 ( .A(n8091), .B(p_input[2719]), .Z(o[2719]) );
  AND U16182 ( .A(p_input[22719]), .B(p_input[12719]), .Z(n8091) );
  AND U16183 ( .A(n8092), .B(p_input[2718]), .Z(o[2718]) );
  AND U16184 ( .A(p_input[22718]), .B(p_input[12718]), .Z(n8092) );
  AND U16185 ( .A(n8093), .B(p_input[2717]), .Z(o[2717]) );
  AND U16186 ( .A(p_input[22717]), .B(p_input[12717]), .Z(n8093) );
  AND U16187 ( .A(n8094), .B(p_input[2716]), .Z(o[2716]) );
  AND U16188 ( .A(p_input[22716]), .B(p_input[12716]), .Z(n8094) );
  AND U16189 ( .A(n8095), .B(p_input[2715]), .Z(o[2715]) );
  AND U16190 ( .A(p_input[22715]), .B(p_input[12715]), .Z(n8095) );
  AND U16191 ( .A(n8096), .B(p_input[2714]), .Z(o[2714]) );
  AND U16192 ( .A(p_input[22714]), .B(p_input[12714]), .Z(n8096) );
  AND U16193 ( .A(n8097), .B(p_input[2713]), .Z(o[2713]) );
  AND U16194 ( .A(p_input[22713]), .B(p_input[12713]), .Z(n8097) );
  AND U16195 ( .A(n8098), .B(p_input[2712]), .Z(o[2712]) );
  AND U16196 ( .A(p_input[22712]), .B(p_input[12712]), .Z(n8098) );
  AND U16197 ( .A(n8099), .B(p_input[2711]), .Z(o[2711]) );
  AND U16198 ( .A(p_input[22711]), .B(p_input[12711]), .Z(n8099) );
  AND U16199 ( .A(n8100), .B(p_input[2710]), .Z(o[2710]) );
  AND U16200 ( .A(p_input[22710]), .B(p_input[12710]), .Z(n8100) );
  AND U16201 ( .A(n8101), .B(p_input[270]), .Z(o[270]) );
  AND U16202 ( .A(p_input[20270]), .B(p_input[10270]), .Z(n8101) );
  AND U16203 ( .A(n8102), .B(p_input[2709]), .Z(o[2709]) );
  AND U16204 ( .A(p_input[22709]), .B(p_input[12709]), .Z(n8102) );
  AND U16205 ( .A(n8103), .B(p_input[2708]), .Z(o[2708]) );
  AND U16206 ( .A(p_input[22708]), .B(p_input[12708]), .Z(n8103) );
  AND U16207 ( .A(n8104), .B(p_input[2707]), .Z(o[2707]) );
  AND U16208 ( .A(p_input[22707]), .B(p_input[12707]), .Z(n8104) );
  AND U16209 ( .A(n8105), .B(p_input[2706]), .Z(o[2706]) );
  AND U16210 ( .A(p_input[22706]), .B(p_input[12706]), .Z(n8105) );
  AND U16211 ( .A(n8106), .B(p_input[2705]), .Z(o[2705]) );
  AND U16212 ( .A(p_input[22705]), .B(p_input[12705]), .Z(n8106) );
  AND U16213 ( .A(n8107), .B(p_input[2704]), .Z(o[2704]) );
  AND U16214 ( .A(p_input[22704]), .B(p_input[12704]), .Z(n8107) );
  AND U16215 ( .A(n8108), .B(p_input[2703]), .Z(o[2703]) );
  AND U16216 ( .A(p_input[22703]), .B(p_input[12703]), .Z(n8108) );
  AND U16217 ( .A(n8109), .B(p_input[2702]), .Z(o[2702]) );
  AND U16218 ( .A(p_input[22702]), .B(p_input[12702]), .Z(n8109) );
  AND U16219 ( .A(n8110), .B(p_input[2701]), .Z(o[2701]) );
  AND U16220 ( .A(p_input[22701]), .B(p_input[12701]), .Z(n8110) );
  AND U16221 ( .A(n8111), .B(p_input[2700]), .Z(o[2700]) );
  AND U16222 ( .A(p_input[22700]), .B(p_input[12700]), .Z(n8111) );
  AND U16223 ( .A(n8112), .B(p_input[26]), .Z(o[26]) );
  AND U16224 ( .A(p_input[20026]), .B(p_input[10026]), .Z(n8112) );
  AND U16225 ( .A(n8113), .B(p_input[269]), .Z(o[269]) );
  AND U16226 ( .A(p_input[20269]), .B(p_input[10269]), .Z(n8113) );
  AND U16227 ( .A(n8114), .B(p_input[2699]), .Z(o[2699]) );
  AND U16228 ( .A(p_input[22699]), .B(p_input[12699]), .Z(n8114) );
  AND U16229 ( .A(n8115), .B(p_input[2698]), .Z(o[2698]) );
  AND U16230 ( .A(p_input[22698]), .B(p_input[12698]), .Z(n8115) );
  AND U16231 ( .A(n8116), .B(p_input[2697]), .Z(o[2697]) );
  AND U16232 ( .A(p_input[22697]), .B(p_input[12697]), .Z(n8116) );
  AND U16233 ( .A(n8117), .B(p_input[2696]), .Z(o[2696]) );
  AND U16234 ( .A(p_input[22696]), .B(p_input[12696]), .Z(n8117) );
  AND U16235 ( .A(n8118), .B(p_input[2695]), .Z(o[2695]) );
  AND U16236 ( .A(p_input[22695]), .B(p_input[12695]), .Z(n8118) );
  AND U16237 ( .A(n8119), .B(p_input[2694]), .Z(o[2694]) );
  AND U16238 ( .A(p_input[22694]), .B(p_input[12694]), .Z(n8119) );
  AND U16239 ( .A(n8120), .B(p_input[2693]), .Z(o[2693]) );
  AND U16240 ( .A(p_input[22693]), .B(p_input[12693]), .Z(n8120) );
  AND U16241 ( .A(n8121), .B(p_input[2692]), .Z(o[2692]) );
  AND U16242 ( .A(p_input[22692]), .B(p_input[12692]), .Z(n8121) );
  AND U16243 ( .A(n8122), .B(p_input[2691]), .Z(o[2691]) );
  AND U16244 ( .A(p_input[22691]), .B(p_input[12691]), .Z(n8122) );
  AND U16245 ( .A(n8123), .B(p_input[2690]), .Z(o[2690]) );
  AND U16246 ( .A(p_input[22690]), .B(p_input[12690]), .Z(n8123) );
  AND U16247 ( .A(n8124), .B(p_input[268]), .Z(o[268]) );
  AND U16248 ( .A(p_input[20268]), .B(p_input[10268]), .Z(n8124) );
  AND U16249 ( .A(n8125), .B(p_input[2689]), .Z(o[2689]) );
  AND U16250 ( .A(p_input[22689]), .B(p_input[12689]), .Z(n8125) );
  AND U16251 ( .A(n8126), .B(p_input[2688]), .Z(o[2688]) );
  AND U16252 ( .A(p_input[22688]), .B(p_input[12688]), .Z(n8126) );
  AND U16253 ( .A(n8127), .B(p_input[2687]), .Z(o[2687]) );
  AND U16254 ( .A(p_input[22687]), .B(p_input[12687]), .Z(n8127) );
  AND U16255 ( .A(n8128), .B(p_input[2686]), .Z(o[2686]) );
  AND U16256 ( .A(p_input[22686]), .B(p_input[12686]), .Z(n8128) );
  AND U16257 ( .A(n8129), .B(p_input[2685]), .Z(o[2685]) );
  AND U16258 ( .A(p_input[22685]), .B(p_input[12685]), .Z(n8129) );
  AND U16259 ( .A(n8130), .B(p_input[2684]), .Z(o[2684]) );
  AND U16260 ( .A(p_input[22684]), .B(p_input[12684]), .Z(n8130) );
  AND U16261 ( .A(n8131), .B(p_input[2683]), .Z(o[2683]) );
  AND U16262 ( .A(p_input[22683]), .B(p_input[12683]), .Z(n8131) );
  AND U16263 ( .A(n8132), .B(p_input[2682]), .Z(o[2682]) );
  AND U16264 ( .A(p_input[22682]), .B(p_input[12682]), .Z(n8132) );
  AND U16265 ( .A(n8133), .B(p_input[2681]), .Z(o[2681]) );
  AND U16266 ( .A(p_input[22681]), .B(p_input[12681]), .Z(n8133) );
  AND U16267 ( .A(n8134), .B(p_input[2680]), .Z(o[2680]) );
  AND U16268 ( .A(p_input[22680]), .B(p_input[12680]), .Z(n8134) );
  AND U16269 ( .A(n8135), .B(p_input[267]), .Z(o[267]) );
  AND U16270 ( .A(p_input[20267]), .B(p_input[10267]), .Z(n8135) );
  AND U16271 ( .A(n8136), .B(p_input[2679]), .Z(o[2679]) );
  AND U16272 ( .A(p_input[22679]), .B(p_input[12679]), .Z(n8136) );
  AND U16273 ( .A(n8137), .B(p_input[2678]), .Z(o[2678]) );
  AND U16274 ( .A(p_input[22678]), .B(p_input[12678]), .Z(n8137) );
  AND U16275 ( .A(n8138), .B(p_input[2677]), .Z(o[2677]) );
  AND U16276 ( .A(p_input[22677]), .B(p_input[12677]), .Z(n8138) );
  AND U16277 ( .A(n8139), .B(p_input[2676]), .Z(o[2676]) );
  AND U16278 ( .A(p_input[22676]), .B(p_input[12676]), .Z(n8139) );
  AND U16279 ( .A(n8140), .B(p_input[2675]), .Z(o[2675]) );
  AND U16280 ( .A(p_input[22675]), .B(p_input[12675]), .Z(n8140) );
  AND U16281 ( .A(n8141), .B(p_input[2674]), .Z(o[2674]) );
  AND U16282 ( .A(p_input[22674]), .B(p_input[12674]), .Z(n8141) );
  AND U16283 ( .A(n8142), .B(p_input[2673]), .Z(o[2673]) );
  AND U16284 ( .A(p_input[22673]), .B(p_input[12673]), .Z(n8142) );
  AND U16285 ( .A(n8143), .B(p_input[2672]), .Z(o[2672]) );
  AND U16286 ( .A(p_input[22672]), .B(p_input[12672]), .Z(n8143) );
  AND U16287 ( .A(n8144), .B(p_input[2671]), .Z(o[2671]) );
  AND U16288 ( .A(p_input[22671]), .B(p_input[12671]), .Z(n8144) );
  AND U16289 ( .A(n8145), .B(p_input[2670]), .Z(o[2670]) );
  AND U16290 ( .A(p_input[22670]), .B(p_input[12670]), .Z(n8145) );
  AND U16291 ( .A(n8146), .B(p_input[266]), .Z(o[266]) );
  AND U16292 ( .A(p_input[20266]), .B(p_input[10266]), .Z(n8146) );
  AND U16293 ( .A(n8147), .B(p_input[2669]), .Z(o[2669]) );
  AND U16294 ( .A(p_input[22669]), .B(p_input[12669]), .Z(n8147) );
  AND U16295 ( .A(n8148), .B(p_input[2668]), .Z(o[2668]) );
  AND U16296 ( .A(p_input[22668]), .B(p_input[12668]), .Z(n8148) );
  AND U16297 ( .A(n8149), .B(p_input[2667]), .Z(o[2667]) );
  AND U16298 ( .A(p_input[22667]), .B(p_input[12667]), .Z(n8149) );
  AND U16299 ( .A(n8150), .B(p_input[2666]), .Z(o[2666]) );
  AND U16300 ( .A(p_input[22666]), .B(p_input[12666]), .Z(n8150) );
  AND U16301 ( .A(n8151), .B(p_input[2665]), .Z(o[2665]) );
  AND U16302 ( .A(p_input[22665]), .B(p_input[12665]), .Z(n8151) );
  AND U16303 ( .A(n8152), .B(p_input[2664]), .Z(o[2664]) );
  AND U16304 ( .A(p_input[22664]), .B(p_input[12664]), .Z(n8152) );
  AND U16305 ( .A(n8153), .B(p_input[2663]), .Z(o[2663]) );
  AND U16306 ( .A(p_input[22663]), .B(p_input[12663]), .Z(n8153) );
  AND U16307 ( .A(n8154), .B(p_input[2662]), .Z(o[2662]) );
  AND U16308 ( .A(p_input[22662]), .B(p_input[12662]), .Z(n8154) );
  AND U16309 ( .A(n8155), .B(p_input[2661]), .Z(o[2661]) );
  AND U16310 ( .A(p_input[22661]), .B(p_input[12661]), .Z(n8155) );
  AND U16311 ( .A(n8156), .B(p_input[2660]), .Z(o[2660]) );
  AND U16312 ( .A(p_input[22660]), .B(p_input[12660]), .Z(n8156) );
  AND U16313 ( .A(n8157), .B(p_input[265]), .Z(o[265]) );
  AND U16314 ( .A(p_input[20265]), .B(p_input[10265]), .Z(n8157) );
  AND U16315 ( .A(n8158), .B(p_input[2659]), .Z(o[2659]) );
  AND U16316 ( .A(p_input[22659]), .B(p_input[12659]), .Z(n8158) );
  AND U16317 ( .A(n8159), .B(p_input[2658]), .Z(o[2658]) );
  AND U16318 ( .A(p_input[22658]), .B(p_input[12658]), .Z(n8159) );
  AND U16319 ( .A(n8160), .B(p_input[2657]), .Z(o[2657]) );
  AND U16320 ( .A(p_input[22657]), .B(p_input[12657]), .Z(n8160) );
  AND U16321 ( .A(n8161), .B(p_input[2656]), .Z(o[2656]) );
  AND U16322 ( .A(p_input[22656]), .B(p_input[12656]), .Z(n8161) );
  AND U16323 ( .A(n8162), .B(p_input[2655]), .Z(o[2655]) );
  AND U16324 ( .A(p_input[22655]), .B(p_input[12655]), .Z(n8162) );
  AND U16325 ( .A(n8163), .B(p_input[2654]), .Z(o[2654]) );
  AND U16326 ( .A(p_input[22654]), .B(p_input[12654]), .Z(n8163) );
  AND U16327 ( .A(n8164), .B(p_input[2653]), .Z(o[2653]) );
  AND U16328 ( .A(p_input[22653]), .B(p_input[12653]), .Z(n8164) );
  AND U16329 ( .A(n8165), .B(p_input[2652]), .Z(o[2652]) );
  AND U16330 ( .A(p_input[22652]), .B(p_input[12652]), .Z(n8165) );
  AND U16331 ( .A(n8166), .B(p_input[2651]), .Z(o[2651]) );
  AND U16332 ( .A(p_input[22651]), .B(p_input[12651]), .Z(n8166) );
  AND U16333 ( .A(n8167), .B(p_input[2650]), .Z(o[2650]) );
  AND U16334 ( .A(p_input[22650]), .B(p_input[12650]), .Z(n8167) );
  AND U16335 ( .A(n8168), .B(p_input[264]), .Z(o[264]) );
  AND U16336 ( .A(p_input[20264]), .B(p_input[10264]), .Z(n8168) );
  AND U16337 ( .A(n8169), .B(p_input[2649]), .Z(o[2649]) );
  AND U16338 ( .A(p_input[22649]), .B(p_input[12649]), .Z(n8169) );
  AND U16339 ( .A(n8170), .B(p_input[2648]), .Z(o[2648]) );
  AND U16340 ( .A(p_input[22648]), .B(p_input[12648]), .Z(n8170) );
  AND U16341 ( .A(n8171), .B(p_input[2647]), .Z(o[2647]) );
  AND U16342 ( .A(p_input[22647]), .B(p_input[12647]), .Z(n8171) );
  AND U16343 ( .A(n8172), .B(p_input[2646]), .Z(o[2646]) );
  AND U16344 ( .A(p_input[22646]), .B(p_input[12646]), .Z(n8172) );
  AND U16345 ( .A(n8173), .B(p_input[2645]), .Z(o[2645]) );
  AND U16346 ( .A(p_input[22645]), .B(p_input[12645]), .Z(n8173) );
  AND U16347 ( .A(n8174), .B(p_input[2644]), .Z(o[2644]) );
  AND U16348 ( .A(p_input[22644]), .B(p_input[12644]), .Z(n8174) );
  AND U16349 ( .A(n8175), .B(p_input[2643]), .Z(o[2643]) );
  AND U16350 ( .A(p_input[22643]), .B(p_input[12643]), .Z(n8175) );
  AND U16351 ( .A(n8176), .B(p_input[2642]), .Z(o[2642]) );
  AND U16352 ( .A(p_input[22642]), .B(p_input[12642]), .Z(n8176) );
  AND U16353 ( .A(n8177), .B(p_input[2641]), .Z(o[2641]) );
  AND U16354 ( .A(p_input[22641]), .B(p_input[12641]), .Z(n8177) );
  AND U16355 ( .A(n8178), .B(p_input[2640]), .Z(o[2640]) );
  AND U16356 ( .A(p_input[22640]), .B(p_input[12640]), .Z(n8178) );
  AND U16357 ( .A(n8179), .B(p_input[263]), .Z(o[263]) );
  AND U16358 ( .A(p_input[20263]), .B(p_input[10263]), .Z(n8179) );
  AND U16359 ( .A(n8180), .B(p_input[2639]), .Z(o[2639]) );
  AND U16360 ( .A(p_input[22639]), .B(p_input[12639]), .Z(n8180) );
  AND U16361 ( .A(n8181), .B(p_input[2638]), .Z(o[2638]) );
  AND U16362 ( .A(p_input[22638]), .B(p_input[12638]), .Z(n8181) );
  AND U16363 ( .A(n8182), .B(p_input[2637]), .Z(o[2637]) );
  AND U16364 ( .A(p_input[22637]), .B(p_input[12637]), .Z(n8182) );
  AND U16365 ( .A(n8183), .B(p_input[2636]), .Z(o[2636]) );
  AND U16366 ( .A(p_input[22636]), .B(p_input[12636]), .Z(n8183) );
  AND U16367 ( .A(n8184), .B(p_input[2635]), .Z(o[2635]) );
  AND U16368 ( .A(p_input[22635]), .B(p_input[12635]), .Z(n8184) );
  AND U16369 ( .A(n8185), .B(p_input[2634]), .Z(o[2634]) );
  AND U16370 ( .A(p_input[22634]), .B(p_input[12634]), .Z(n8185) );
  AND U16371 ( .A(n8186), .B(p_input[2633]), .Z(o[2633]) );
  AND U16372 ( .A(p_input[22633]), .B(p_input[12633]), .Z(n8186) );
  AND U16373 ( .A(n8187), .B(p_input[2632]), .Z(o[2632]) );
  AND U16374 ( .A(p_input[22632]), .B(p_input[12632]), .Z(n8187) );
  AND U16375 ( .A(n8188), .B(p_input[2631]), .Z(o[2631]) );
  AND U16376 ( .A(p_input[22631]), .B(p_input[12631]), .Z(n8188) );
  AND U16377 ( .A(n8189), .B(p_input[2630]), .Z(o[2630]) );
  AND U16378 ( .A(p_input[22630]), .B(p_input[12630]), .Z(n8189) );
  AND U16379 ( .A(n8190), .B(p_input[262]), .Z(o[262]) );
  AND U16380 ( .A(p_input[20262]), .B(p_input[10262]), .Z(n8190) );
  AND U16381 ( .A(n8191), .B(p_input[2629]), .Z(o[2629]) );
  AND U16382 ( .A(p_input[22629]), .B(p_input[12629]), .Z(n8191) );
  AND U16383 ( .A(n8192), .B(p_input[2628]), .Z(o[2628]) );
  AND U16384 ( .A(p_input[22628]), .B(p_input[12628]), .Z(n8192) );
  AND U16385 ( .A(n8193), .B(p_input[2627]), .Z(o[2627]) );
  AND U16386 ( .A(p_input[22627]), .B(p_input[12627]), .Z(n8193) );
  AND U16387 ( .A(n8194), .B(p_input[2626]), .Z(o[2626]) );
  AND U16388 ( .A(p_input[22626]), .B(p_input[12626]), .Z(n8194) );
  AND U16389 ( .A(n8195), .B(p_input[2625]), .Z(o[2625]) );
  AND U16390 ( .A(p_input[22625]), .B(p_input[12625]), .Z(n8195) );
  AND U16391 ( .A(n8196), .B(p_input[2624]), .Z(o[2624]) );
  AND U16392 ( .A(p_input[22624]), .B(p_input[12624]), .Z(n8196) );
  AND U16393 ( .A(n8197), .B(p_input[2623]), .Z(o[2623]) );
  AND U16394 ( .A(p_input[22623]), .B(p_input[12623]), .Z(n8197) );
  AND U16395 ( .A(n8198), .B(p_input[2622]), .Z(o[2622]) );
  AND U16396 ( .A(p_input[22622]), .B(p_input[12622]), .Z(n8198) );
  AND U16397 ( .A(n8199), .B(p_input[2621]), .Z(o[2621]) );
  AND U16398 ( .A(p_input[22621]), .B(p_input[12621]), .Z(n8199) );
  AND U16399 ( .A(n8200), .B(p_input[2620]), .Z(o[2620]) );
  AND U16400 ( .A(p_input[22620]), .B(p_input[12620]), .Z(n8200) );
  AND U16401 ( .A(n8201), .B(p_input[261]), .Z(o[261]) );
  AND U16402 ( .A(p_input[20261]), .B(p_input[10261]), .Z(n8201) );
  AND U16403 ( .A(n8202), .B(p_input[2619]), .Z(o[2619]) );
  AND U16404 ( .A(p_input[22619]), .B(p_input[12619]), .Z(n8202) );
  AND U16405 ( .A(n8203), .B(p_input[2618]), .Z(o[2618]) );
  AND U16406 ( .A(p_input[22618]), .B(p_input[12618]), .Z(n8203) );
  AND U16407 ( .A(n8204), .B(p_input[2617]), .Z(o[2617]) );
  AND U16408 ( .A(p_input[22617]), .B(p_input[12617]), .Z(n8204) );
  AND U16409 ( .A(n8205), .B(p_input[2616]), .Z(o[2616]) );
  AND U16410 ( .A(p_input[22616]), .B(p_input[12616]), .Z(n8205) );
  AND U16411 ( .A(n8206), .B(p_input[2615]), .Z(o[2615]) );
  AND U16412 ( .A(p_input[22615]), .B(p_input[12615]), .Z(n8206) );
  AND U16413 ( .A(n8207), .B(p_input[2614]), .Z(o[2614]) );
  AND U16414 ( .A(p_input[22614]), .B(p_input[12614]), .Z(n8207) );
  AND U16415 ( .A(n8208), .B(p_input[2613]), .Z(o[2613]) );
  AND U16416 ( .A(p_input[22613]), .B(p_input[12613]), .Z(n8208) );
  AND U16417 ( .A(n8209), .B(p_input[2612]), .Z(o[2612]) );
  AND U16418 ( .A(p_input[22612]), .B(p_input[12612]), .Z(n8209) );
  AND U16419 ( .A(n8210), .B(p_input[2611]), .Z(o[2611]) );
  AND U16420 ( .A(p_input[22611]), .B(p_input[12611]), .Z(n8210) );
  AND U16421 ( .A(n8211), .B(p_input[2610]), .Z(o[2610]) );
  AND U16422 ( .A(p_input[22610]), .B(p_input[12610]), .Z(n8211) );
  AND U16423 ( .A(n8212), .B(p_input[260]), .Z(o[260]) );
  AND U16424 ( .A(p_input[20260]), .B(p_input[10260]), .Z(n8212) );
  AND U16425 ( .A(n8213), .B(p_input[2609]), .Z(o[2609]) );
  AND U16426 ( .A(p_input[22609]), .B(p_input[12609]), .Z(n8213) );
  AND U16427 ( .A(n8214), .B(p_input[2608]), .Z(o[2608]) );
  AND U16428 ( .A(p_input[22608]), .B(p_input[12608]), .Z(n8214) );
  AND U16429 ( .A(n8215), .B(p_input[2607]), .Z(o[2607]) );
  AND U16430 ( .A(p_input[22607]), .B(p_input[12607]), .Z(n8215) );
  AND U16431 ( .A(n8216), .B(p_input[2606]), .Z(o[2606]) );
  AND U16432 ( .A(p_input[22606]), .B(p_input[12606]), .Z(n8216) );
  AND U16433 ( .A(n8217), .B(p_input[2605]), .Z(o[2605]) );
  AND U16434 ( .A(p_input[22605]), .B(p_input[12605]), .Z(n8217) );
  AND U16435 ( .A(n8218), .B(p_input[2604]), .Z(o[2604]) );
  AND U16436 ( .A(p_input[22604]), .B(p_input[12604]), .Z(n8218) );
  AND U16437 ( .A(n8219), .B(p_input[2603]), .Z(o[2603]) );
  AND U16438 ( .A(p_input[22603]), .B(p_input[12603]), .Z(n8219) );
  AND U16439 ( .A(n8220), .B(p_input[2602]), .Z(o[2602]) );
  AND U16440 ( .A(p_input[22602]), .B(p_input[12602]), .Z(n8220) );
  AND U16441 ( .A(n8221), .B(p_input[2601]), .Z(o[2601]) );
  AND U16442 ( .A(p_input[22601]), .B(p_input[12601]), .Z(n8221) );
  AND U16443 ( .A(n8222), .B(p_input[2600]), .Z(o[2600]) );
  AND U16444 ( .A(p_input[22600]), .B(p_input[12600]), .Z(n8222) );
  AND U16445 ( .A(n8223), .B(p_input[25]), .Z(o[25]) );
  AND U16446 ( .A(p_input[20025]), .B(p_input[10025]), .Z(n8223) );
  AND U16447 ( .A(n8224), .B(p_input[259]), .Z(o[259]) );
  AND U16448 ( .A(p_input[20259]), .B(p_input[10259]), .Z(n8224) );
  AND U16449 ( .A(n8225), .B(p_input[2599]), .Z(o[2599]) );
  AND U16450 ( .A(p_input[22599]), .B(p_input[12599]), .Z(n8225) );
  AND U16451 ( .A(n8226), .B(p_input[2598]), .Z(o[2598]) );
  AND U16452 ( .A(p_input[22598]), .B(p_input[12598]), .Z(n8226) );
  AND U16453 ( .A(n8227), .B(p_input[2597]), .Z(o[2597]) );
  AND U16454 ( .A(p_input[22597]), .B(p_input[12597]), .Z(n8227) );
  AND U16455 ( .A(n8228), .B(p_input[2596]), .Z(o[2596]) );
  AND U16456 ( .A(p_input[22596]), .B(p_input[12596]), .Z(n8228) );
  AND U16457 ( .A(n8229), .B(p_input[2595]), .Z(o[2595]) );
  AND U16458 ( .A(p_input[22595]), .B(p_input[12595]), .Z(n8229) );
  AND U16459 ( .A(n8230), .B(p_input[2594]), .Z(o[2594]) );
  AND U16460 ( .A(p_input[22594]), .B(p_input[12594]), .Z(n8230) );
  AND U16461 ( .A(n8231), .B(p_input[2593]), .Z(o[2593]) );
  AND U16462 ( .A(p_input[22593]), .B(p_input[12593]), .Z(n8231) );
  AND U16463 ( .A(n8232), .B(p_input[2592]), .Z(o[2592]) );
  AND U16464 ( .A(p_input[22592]), .B(p_input[12592]), .Z(n8232) );
  AND U16465 ( .A(n8233), .B(p_input[2591]), .Z(o[2591]) );
  AND U16466 ( .A(p_input[22591]), .B(p_input[12591]), .Z(n8233) );
  AND U16467 ( .A(n8234), .B(p_input[2590]), .Z(o[2590]) );
  AND U16468 ( .A(p_input[22590]), .B(p_input[12590]), .Z(n8234) );
  AND U16469 ( .A(n8235), .B(p_input[258]), .Z(o[258]) );
  AND U16470 ( .A(p_input[20258]), .B(p_input[10258]), .Z(n8235) );
  AND U16471 ( .A(n8236), .B(p_input[2589]), .Z(o[2589]) );
  AND U16472 ( .A(p_input[22589]), .B(p_input[12589]), .Z(n8236) );
  AND U16473 ( .A(n8237), .B(p_input[2588]), .Z(o[2588]) );
  AND U16474 ( .A(p_input[22588]), .B(p_input[12588]), .Z(n8237) );
  AND U16475 ( .A(n8238), .B(p_input[2587]), .Z(o[2587]) );
  AND U16476 ( .A(p_input[22587]), .B(p_input[12587]), .Z(n8238) );
  AND U16477 ( .A(n8239), .B(p_input[2586]), .Z(o[2586]) );
  AND U16478 ( .A(p_input[22586]), .B(p_input[12586]), .Z(n8239) );
  AND U16479 ( .A(n8240), .B(p_input[2585]), .Z(o[2585]) );
  AND U16480 ( .A(p_input[22585]), .B(p_input[12585]), .Z(n8240) );
  AND U16481 ( .A(n8241), .B(p_input[2584]), .Z(o[2584]) );
  AND U16482 ( .A(p_input[22584]), .B(p_input[12584]), .Z(n8241) );
  AND U16483 ( .A(n8242), .B(p_input[2583]), .Z(o[2583]) );
  AND U16484 ( .A(p_input[22583]), .B(p_input[12583]), .Z(n8242) );
  AND U16485 ( .A(n8243), .B(p_input[2582]), .Z(o[2582]) );
  AND U16486 ( .A(p_input[22582]), .B(p_input[12582]), .Z(n8243) );
  AND U16487 ( .A(n8244), .B(p_input[2581]), .Z(o[2581]) );
  AND U16488 ( .A(p_input[22581]), .B(p_input[12581]), .Z(n8244) );
  AND U16489 ( .A(n8245), .B(p_input[2580]), .Z(o[2580]) );
  AND U16490 ( .A(p_input[22580]), .B(p_input[12580]), .Z(n8245) );
  AND U16491 ( .A(n8246), .B(p_input[257]), .Z(o[257]) );
  AND U16492 ( .A(p_input[20257]), .B(p_input[10257]), .Z(n8246) );
  AND U16493 ( .A(n8247), .B(p_input[2579]), .Z(o[2579]) );
  AND U16494 ( .A(p_input[22579]), .B(p_input[12579]), .Z(n8247) );
  AND U16495 ( .A(n8248), .B(p_input[2578]), .Z(o[2578]) );
  AND U16496 ( .A(p_input[22578]), .B(p_input[12578]), .Z(n8248) );
  AND U16497 ( .A(n8249), .B(p_input[2577]), .Z(o[2577]) );
  AND U16498 ( .A(p_input[22577]), .B(p_input[12577]), .Z(n8249) );
  AND U16499 ( .A(n8250), .B(p_input[2576]), .Z(o[2576]) );
  AND U16500 ( .A(p_input[22576]), .B(p_input[12576]), .Z(n8250) );
  AND U16501 ( .A(n8251), .B(p_input[2575]), .Z(o[2575]) );
  AND U16502 ( .A(p_input[22575]), .B(p_input[12575]), .Z(n8251) );
  AND U16503 ( .A(n8252), .B(p_input[2574]), .Z(o[2574]) );
  AND U16504 ( .A(p_input[22574]), .B(p_input[12574]), .Z(n8252) );
  AND U16505 ( .A(n8253), .B(p_input[2573]), .Z(o[2573]) );
  AND U16506 ( .A(p_input[22573]), .B(p_input[12573]), .Z(n8253) );
  AND U16507 ( .A(n8254), .B(p_input[2572]), .Z(o[2572]) );
  AND U16508 ( .A(p_input[22572]), .B(p_input[12572]), .Z(n8254) );
  AND U16509 ( .A(n8255), .B(p_input[2571]), .Z(o[2571]) );
  AND U16510 ( .A(p_input[22571]), .B(p_input[12571]), .Z(n8255) );
  AND U16511 ( .A(n8256), .B(p_input[2570]), .Z(o[2570]) );
  AND U16512 ( .A(p_input[22570]), .B(p_input[12570]), .Z(n8256) );
  AND U16513 ( .A(n8257), .B(p_input[256]), .Z(o[256]) );
  AND U16514 ( .A(p_input[20256]), .B(p_input[10256]), .Z(n8257) );
  AND U16515 ( .A(n8258), .B(p_input[2569]), .Z(o[2569]) );
  AND U16516 ( .A(p_input[22569]), .B(p_input[12569]), .Z(n8258) );
  AND U16517 ( .A(n8259), .B(p_input[2568]), .Z(o[2568]) );
  AND U16518 ( .A(p_input[22568]), .B(p_input[12568]), .Z(n8259) );
  AND U16519 ( .A(n8260), .B(p_input[2567]), .Z(o[2567]) );
  AND U16520 ( .A(p_input[22567]), .B(p_input[12567]), .Z(n8260) );
  AND U16521 ( .A(n8261), .B(p_input[2566]), .Z(o[2566]) );
  AND U16522 ( .A(p_input[22566]), .B(p_input[12566]), .Z(n8261) );
  AND U16523 ( .A(n8262), .B(p_input[2565]), .Z(o[2565]) );
  AND U16524 ( .A(p_input[22565]), .B(p_input[12565]), .Z(n8262) );
  AND U16525 ( .A(n8263), .B(p_input[2564]), .Z(o[2564]) );
  AND U16526 ( .A(p_input[22564]), .B(p_input[12564]), .Z(n8263) );
  AND U16527 ( .A(n8264), .B(p_input[2563]), .Z(o[2563]) );
  AND U16528 ( .A(p_input[22563]), .B(p_input[12563]), .Z(n8264) );
  AND U16529 ( .A(n8265), .B(p_input[2562]), .Z(o[2562]) );
  AND U16530 ( .A(p_input[22562]), .B(p_input[12562]), .Z(n8265) );
  AND U16531 ( .A(n8266), .B(p_input[2561]), .Z(o[2561]) );
  AND U16532 ( .A(p_input[22561]), .B(p_input[12561]), .Z(n8266) );
  AND U16533 ( .A(n8267), .B(p_input[2560]), .Z(o[2560]) );
  AND U16534 ( .A(p_input[22560]), .B(p_input[12560]), .Z(n8267) );
  AND U16535 ( .A(n8268), .B(p_input[255]), .Z(o[255]) );
  AND U16536 ( .A(p_input[20255]), .B(p_input[10255]), .Z(n8268) );
  AND U16537 ( .A(n8269), .B(p_input[2559]), .Z(o[2559]) );
  AND U16538 ( .A(p_input[22559]), .B(p_input[12559]), .Z(n8269) );
  AND U16539 ( .A(n8270), .B(p_input[2558]), .Z(o[2558]) );
  AND U16540 ( .A(p_input[22558]), .B(p_input[12558]), .Z(n8270) );
  AND U16541 ( .A(n8271), .B(p_input[2557]), .Z(o[2557]) );
  AND U16542 ( .A(p_input[22557]), .B(p_input[12557]), .Z(n8271) );
  AND U16543 ( .A(n8272), .B(p_input[2556]), .Z(o[2556]) );
  AND U16544 ( .A(p_input[22556]), .B(p_input[12556]), .Z(n8272) );
  AND U16545 ( .A(n8273), .B(p_input[2555]), .Z(o[2555]) );
  AND U16546 ( .A(p_input[22555]), .B(p_input[12555]), .Z(n8273) );
  AND U16547 ( .A(n8274), .B(p_input[2554]), .Z(o[2554]) );
  AND U16548 ( .A(p_input[22554]), .B(p_input[12554]), .Z(n8274) );
  AND U16549 ( .A(n8275), .B(p_input[2553]), .Z(o[2553]) );
  AND U16550 ( .A(p_input[22553]), .B(p_input[12553]), .Z(n8275) );
  AND U16551 ( .A(n8276), .B(p_input[2552]), .Z(o[2552]) );
  AND U16552 ( .A(p_input[22552]), .B(p_input[12552]), .Z(n8276) );
  AND U16553 ( .A(n8277), .B(p_input[2551]), .Z(o[2551]) );
  AND U16554 ( .A(p_input[22551]), .B(p_input[12551]), .Z(n8277) );
  AND U16555 ( .A(n8278), .B(p_input[2550]), .Z(o[2550]) );
  AND U16556 ( .A(p_input[22550]), .B(p_input[12550]), .Z(n8278) );
  AND U16557 ( .A(n8279), .B(p_input[254]), .Z(o[254]) );
  AND U16558 ( .A(p_input[20254]), .B(p_input[10254]), .Z(n8279) );
  AND U16559 ( .A(n8280), .B(p_input[2549]), .Z(o[2549]) );
  AND U16560 ( .A(p_input[22549]), .B(p_input[12549]), .Z(n8280) );
  AND U16561 ( .A(n8281), .B(p_input[2548]), .Z(o[2548]) );
  AND U16562 ( .A(p_input[22548]), .B(p_input[12548]), .Z(n8281) );
  AND U16563 ( .A(n8282), .B(p_input[2547]), .Z(o[2547]) );
  AND U16564 ( .A(p_input[22547]), .B(p_input[12547]), .Z(n8282) );
  AND U16565 ( .A(n8283), .B(p_input[2546]), .Z(o[2546]) );
  AND U16566 ( .A(p_input[22546]), .B(p_input[12546]), .Z(n8283) );
  AND U16567 ( .A(n8284), .B(p_input[2545]), .Z(o[2545]) );
  AND U16568 ( .A(p_input[22545]), .B(p_input[12545]), .Z(n8284) );
  AND U16569 ( .A(n8285), .B(p_input[2544]), .Z(o[2544]) );
  AND U16570 ( .A(p_input[22544]), .B(p_input[12544]), .Z(n8285) );
  AND U16571 ( .A(n8286), .B(p_input[2543]), .Z(o[2543]) );
  AND U16572 ( .A(p_input[22543]), .B(p_input[12543]), .Z(n8286) );
  AND U16573 ( .A(n8287), .B(p_input[2542]), .Z(o[2542]) );
  AND U16574 ( .A(p_input[22542]), .B(p_input[12542]), .Z(n8287) );
  AND U16575 ( .A(n8288), .B(p_input[2541]), .Z(o[2541]) );
  AND U16576 ( .A(p_input[22541]), .B(p_input[12541]), .Z(n8288) );
  AND U16577 ( .A(n8289), .B(p_input[2540]), .Z(o[2540]) );
  AND U16578 ( .A(p_input[22540]), .B(p_input[12540]), .Z(n8289) );
  AND U16579 ( .A(n8290), .B(p_input[253]), .Z(o[253]) );
  AND U16580 ( .A(p_input[20253]), .B(p_input[10253]), .Z(n8290) );
  AND U16581 ( .A(n8291), .B(p_input[2539]), .Z(o[2539]) );
  AND U16582 ( .A(p_input[22539]), .B(p_input[12539]), .Z(n8291) );
  AND U16583 ( .A(n8292), .B(p_input[2538]), .Z(o[2538]) );
  AND U16584 ( .A(p_input[22538]), .B(p_input[12538]), .Z(n8292) );
  AND U16585 ( .A(n8293), .B(p_input[2537]), .Z(o[2537]) );
  AND U16586 ( .A(p_input[22537]), .B(p_input[12537]), .Z(n8293) );
  AND U16587 ( .A(n8294), .B(p_input[2536]), .Z(o[2536]) );
  AND U16588 ( .A(p_input[22536]), .B(p_input[12536]), .Z(n8294) );
  AND U16589 ( .A(n8295), .B(p_input[2535]), .Z(o[2535]) );
  AND U16590 ( .A(p_input[22535]), .B(p_input[12535]), .Z(n8295) );
  AND U16591 ( .A(n8296), .B(p_input[2534]), .Z(o[2534]) );
  AND U16592 ( .A(p_input[22534]), .B(p_input[12534]), .Z(n8296) );
  AND U16593 ( .A(n8297), .B(p_input[2533]), .Z(o[2533]) );
  AND U16594 ( .A(p_input[22533]), .B(p_input[12533]), .Z(n8297) );
  AND U16595 ( .A(n8298), .B(p_input[2532]), .Z(o[2532]) );
  AND U16596 ( .A(p_input[22532]), .B(p_input[12532]), .Z(n8298) );
  AND U16597 ( .A(n8299), .B(p_input[2531]), .Z(o[2531]) );
  AND U16598 ( .A(p_input[22531]), .B(p_input[12531]), .Z(n8299) );
  AND U16599 ( .A(n8300), .B(p_input[2530]), .Z(o[2530]) );
  AND U16600 ( .A(p_input[22530]), .B(p_input[12530]), .Z(n8300) );
  AND U16601 ( .A(n8301), .B(p_input[252]), .Z(o[252]) );
  AND U16602 ( .A(p_input[20252]), .B(p_input[10252]), .Z(n8301) );
  AND U16603 ( .A(n8302), .B(p_input[2529]), .Z(o[2529]) );
  AND U16604 ( .A(p_input[22529]), .B(p_input[12529]), .Z(n8302) );
  AND U16605 ( .A(n8303), .B(p_input[2528]), .Z(o[2528]) );
  AND U16606 ( .A(p_input[22528]), .B(p_input[12528]), .Z(n8303) );
  AND U16607 ( .A(n8304), .B(p_input[2527]), .Z(o[2527]) );
  AND U16608 ( .A(p_input[22527]), .B(p_input[12527]), .Z(n8304) );
  AND U16609 ( .A(n8305), .B(p_input[2526]), .Z(o[2526]) );
  AND U16610 ( .A(p_input[22526]), .B(p_input[12526]), .Z(n8305) );
  AND U16611 ( .A(n8306), .B(p_input[2525]), .Z(o[2525]) );
  AND U16612 ( .A(p_input[22525]), .B(p_input[12525]), .Z(n8306) );
  AND U16613 ( .A(n8307), .B(p_input[2524]), .Z(o[2524]) );
  AND U16614 ( .A(p_input[22524]), .B(p_input[12524]), .Z(n8307) );
  AND U16615 ( .A(n8308), .B(p_input[2523]), .Z(o[2523]) );
  AND U16616 ( .A(p_input[22523]), .B(p_input[12523]), .Z(n8308) );
  AND U16617 ( .A(n8309), .B(p_input[2522]), .Z(o[2522]) );
  AND U16618 ( .A(p_input[22522]), .B(p_input[12522]), .Z(n8309) );
  AND U16619 ( .A(n8310), .B(p_input[2521]), .Z(o[2521]) );
  AND U16620 ( .A(p_input[22521]), .B(p_input[12521]), .Z(n8310) );
  AND U16621 ( .A(n8311), .B(p_input[2520]), .Z(o[2520]) );
  AND U16622 ( .A(p_input[22520]), .B(p_input[12520]), .Z(n8311) );
  AND U16623 ( .A(n8312), .B(p_input[251]), .Z(o[251]) );
  AND U16624 ( .A(p_input[20251]), .B(p_input[10251]), .Z(n8312) );
  AND U16625 ( .A(n8313), .B(p_input[2519]), .Z(o[2519]) );
  AND U16626 ( .A(p_input[22519]), .B(p_input[12519]), .Z(n8313) );
  AND U16627 ( .A(n8314), .B(p_input[2518]), .Z(o[2518]) );
  AND U16628 ( .A(p_input[22518]), .B(p_input[12518]), .Z(n8314) );
  AND U16629 ( .A(n8315), .B(p_input[2517]), .Z(o[2517]) );
  AND U16630 ( .A(p_input[22517]), .B(p_input[12517]), .Z(n8315) );
  AND U16631 ( .A(n8316), .B(p_input[2516]), .Z(o[2516]) );
  AND U16632 ( .A(p_input[22516]), .B(p_input[12516]), .Z(n8316) );
  AND U16633 ( .A(n8317), .B(p_input[2515]), .Z(o[2515]) );
  AND U16634 ( .A(p_input[22515]), .B(p_input[12515]), .Z(n8317) );
  AND U16635 ( .A(n8318), .B(p_input[2514]), .Z(o[2514]) );
  AND U16636 ( .A(p_input[22514]), .B(p_input[12514]), .Z(n8318) );
  AND U16637 ( .A(n8319), .B(p_input[2513]), .Z(o[2513]) );
  AND U16638 ( .A(p_input[22513]), .B(p_input[12513]), .Z(n8319) );
  AND U16639 ( .A(n8320), .B(p_input[2512]), .Z(o[2512]) );
  AND U16640 ( .A(p_input[22512]), .B(p_input[12512]), .Z(n8320) );
  AND U16641 ( .A(n8321), .B(p_input[2511]), .Z(o[2511]) );
  AND U16642 ( .A(p_input[22511]), .B(p_input[12511]), .Z(n8321) );
  AND U16643 ( .A(n8322), .B(p_input[2510]), .Z(o[2510]) );
  AND U16644 ( .A(p_input[22510]), .B(p_input[12510]), .Z(n8322) );
  AND U16645 ( .A(n8323), .B(p_input[250]), .Z(o[250]) );
  AND U16646 ( .A(p_input[20250]), .B(p_input[10250]), .Z(n8323) );
  AND U16647 ( .A(n8324), .B(p_input[2509]), .Z(o[2509]) );
  AND U16648 ( .A(p_input[22509]), .B(p_input[12509]), .Z(n8324) );
  AND U16649 ( .A(n8325), .B(p_input[2508]), .Z(o[2508]) );
  AND U16650 ( .A(p_input[22508]), .B(p_input[12508]), .Z(n8325) );
  AND U16651 ( .A(n8326), .B(p_input[2507]), .Z(o[2507]) );
  AND U16652 ( .A(p_input[22507]), .B(p_input[12507]), .Z(n8326) );
  AND U16653 ( .A(n8327), .B(p_input[2506]), .Z(o[2506]) );
  AND U16654 ( .A(p_input[22506]), .B(p_input[12506]), .Z(n8327) );
  AND U16655 ( .A(n8328), .B(p_input[2505]), .Z(o[2505]) );
  AND U16656 ( .A(p_input[22505]), .B(p_input[12505]), .Z(n8328) );
  AND U16657 ( .A(n8329), .B(p_input[2504]), .Z(o[2504]) );
  AND U16658 ( .A(p_input[22504]), .B(p_input[12504]), .Z(n8329) );
  AND U16659 ( .A(n8330), .B(p_input[2503]), .Z(o[2503]) );
  AND U16660 ( .A(p_input[22503]), .B(p_input[12503]), .Z(n8330) );
  AND U16661 ( .A(n8331), .B(p_input[2502]), .Z(o[2502]) );
  AND U16662 ( .A(p_input[22502]), .B(p_input[12502]), .Z(n8331) );
  AND U16663 ( .A(n8332), .B(p_input[2501]), .Z(o[2501]) );
  AND U16664 ( .A(p_input[22501]), .B(p_input[12501]), .Z(n8332) );
  AND U16665 ( .A(n8333), .B(p_input[2500]), .Z(o[2500]) );
  AND U16666 ( .A(p_input[22500]), .B(p_input[12500]), .Z(n8333) );
  AND U16667 ( .A(n8334), .B(p_input[24]), .Z(o[24]) );
  AND U16668 ( .A(p_input[20024]), .B(p_input[10024]), .Z(n8334) );
  AND U16669 ( .A(n8335), .B(p_input[249]), .Z(o[249]) );
  AND U16670 ( .A(p_input[20249]), .B(p_input[10249]), .Z(n8335) );
  AND U16671 ( .A(n8336), .B(p_input[2499]), .Z(o[2499]) );
  AND U16672 ( .A(p_input[22499]), .B(p_input[12499]), .Z(n8336) );
  AND U16673 ( .A(n8337), .B(p_input[2498]), .Z(o[2498]) );
  AND U16674 ( .A(p_input[22498]), .B(p_input[12498]), .Z(n8337) );
  AND U16675 ( .A(n8338), .B(p_input[2497]), .Z(o[2497]) );
  AND U16676 ( .A(p_input[22497]), .B(p_input[12497]), .Z(n8338) );
  AND U16677 ( .A(n8339), .B(p_input[2496]), .Z(o[2496]) );
  AND U16678 ( .A(p_input[22496]), .B(p_input[12496]), .Z(n8339) );
  AND U16679 ( .A(n8340), .B(p_input[2495]), .Z(o[2495]) );
  AND U16680 ( .A(p_input[22495]), .B(p_input[12495]), .Z(n8340) );
  AND U16681 ( .A(n8341), .B(p_input[2494]), .Z(o[2494]) );
  AND U16682 ( .A(p_input[22494]), .B(p_input[12494]), .Z(n8341) );
  AND U16683 ( .A(n8342), .B(p_input[2493]), .Z(o[2493]) );
  AND U16684 ( .A(p_input[22493]), .B(p_input[12493]), .Z(n8342) );
  AND U16685 ( .A(n8343), .B(p_input[2492]), .Z(o[2492]) );
  AND U16686 ( .A(p_input[22492]), .B(p_input[12492]), .Z(n8343) );
  AND U16687 ( .A(n8344), .B(p_input[2491]), .Z(o[2491]) );
  AND U16688 ( .A(p_input[22491]), .B(p_input[12491]), .Z(n8344) );
  AND U16689 ( .A(n8345), .B(p_input[2490]), .Z(o[2490]) );
  AND U16690 ( .A(p_input[22490]), .B(p_input[12490]), .Z(n8345) );
  AND U16691 ( .A(n8346), .B(p_input[248]), .Z(o[248]) );
  AND U16692 ( .A(p_input[20248]), .B(p_input[10248]), .Z(n8346) );
  AND U16693 ( .A(n8347), .B(p_input[2489]), .Z(o[2489]) );
  AND U16694 ( .A(p_input[22489]), .B(p_input[12489]), .Z(n8347) );
  AND U16695 ( .A(n8348), .B(p_input[2488]), .Z(o[2488]) );
  AND U16696 ( .A(p_input[22488]), .B(p_input[12488]), .Z(n8348) );
  AND U16697 ( .A(n8349), .B(p_input[2487]), .Z(o[2487]) );
  AND U16698 ( .A(p_input[22487]), .B(p_input[12487]), .Z(n8349) );
  AND U16699 ( .A(n8350), .B(p_input[2486]), .Z(o[2486]) );
  AND U16700 ( .A(p_input[22486]), .B(p_input[12486]), .Z(n8350) );
  AND U16701 ( .A(n8351), .B(p_input[2485]), .Z(o[2485]) );
  AND U16702 ( .A(p_input[22485]), .B(p_input[12485]), .Z(n8351) );
  AND U16703 ( .A(n8352), .B(p_input[2484]), .Z(o[2484]) );
  AND U16704 ( .A(p_input[22484]), .B(p_input[12484]), .Z(n8352) );
  AND U16705 ( .A(n8353), .B(p_input[2483]), .Z(o[2483]) );
  AND U16706 ( .A(p_input[22483]), .B(p_input[12483]), .Z(n8353) );
  AND U16707 ( .A(n8354), .B(p_input[2482]), .Z(o[2482]) );
  AND U16708 ( .A(p_input[22482]), .B(p_input[12482]), .Z(n8354) );
  AND U16709 ( .A(n8355), .B(p_input[2481]), .Z(o[2481]) );
  AND U16710 ( .A(p_input[22481]), .B(p_input[12481]), .Z(n8355) );
  AND U16711 ( .A(n8356), .B(p_input[2480]), .Z(o[2480]) );
  AND U16712 ( .A(p_input[22480]), .B(p_input[12480]), .Z(n8356) );
  AND U16713 ( .A(n8357), .B(p_input[247]), .Z(o[247]) );
  AND U16714 ( .A(p_input[20247]), .B(p_input[10247]), .Z(n8357) );
  AND U16715 ( .A(n8358), .B(p_input[2479]), .Z(o[2479]) );
  AND U16716 ( .A(p_input[22479]), .B(p_input[12479]), .Z(n8358) );
  AND U16717 ( .A(n8359), .B(p_input[2478]), .Z(o[2478]) );
  AND U16718 ( .A(p_input[22478]), .B(p_input[12478]), .Z(n8359) );
  AND U16719 ( .A(n8360), .B(p_input[2477]), .Z(o[2477]) );
  AND U16720 ( .A(p_input[22477]), .B(p_input[12477]), .Z(n8360) );
  AND U16721 ( .A(n8361), .B(p_input[2476]), .Z(o[2476]) );
  AND U16722 ( .A(p_input[22476]), .B(p_input[12476]), .Z(n8361) );
  AND U16723 ( .A(n8362), .B(p_input[2475]), .Z(o[2475]) );
  AND U16724 ( .A(p_input[22475]), .B(p_input[12475]), .Z(n8362) );
  AND U16725 ( .A(n8363), .B(p_input[2474]), .Z(o[2474]) );
  AND U16726 ( .A(p_input[22474]), .B(p_input[12474]), .Z(n8363) );
  AND U16727 ( .A(n8364), .B(p_input[2473]), .Z(o[2473]) );
  AND U16728 ( .A(p_input[22473]), .B(p_input[12473]), .Z(n8364) );
  AND U16729 ( .A(n8365), .B(p_input[2472]), .Z(o[2472]) );
  AND U16730 ( .A(p_input[22472]), .B(p_input[12472]), .Z(n8365) );
  AND U16731 ( .A(n8366), .B(p_input[2471]), .Z(o[2471]) );
  AND U16732 ( .A(p_input[22471]), .B(p_input[12471]), .Z(n8366) );
  AND U16733 ( .A(n8367), .B(p_input[2470]), .Z(o[2470]) );
  AND U16734 ( .A(p_input[22470]), .B(p_input[12470]), .Z(n8367) );
  AND U16735 ( .A(n8368), .B(p_input[246]), .Z(o[246]) );
  AND U16736 ( .A(p_input[20246]), .B(p_input[10246]), .Z(n8368) );
  AND U16737 ( .A(n8369), .B(p_input[2469]), .Z(o[2469]) );
  AND U16738 ( .A(p_input[22469]), .B(p_input[12469]), .Z(n8369) );
  AND U16739 ( .A(n8370), .B(p_input[2468]), .Z(o[2468]) );
  AND U16740 ( .A(p_input[22468]), .B(p_input[12468]), .Z(n8370) );
  AND U16741 ( .A(n8371), .B(p_input[2467]), .Z(o[2467]) );
  AND U16742 ( .A(p_input[22467]), .B(p_input[12467]), .Z(n8371) );
  AND U16743 ( .A(n8372), .B(p_input[2466]), .Z(o[2466]) );
  AND U16744 ( .A(p_input[22466]), .B(p_input[12466]), .Z(n8372) );
  AND U16745 ( .A(n8373), .B(p_input[2465]), .Z(o[2465]) );
  AND U16746 ( .A(p_input[22465]), .B(p_input[12465]), .Z(n8373) );
  AND U16747 ( .A(n8374), .B(p_input[2464]), .Z(o[2464]) );
  AND U16748 ( .A(p_input[22464]), .B(p_input[12464]), .Z(n8374) );
  AND U16749 ( .A(n8375), .B(p_input[2463]), .Z(o[2463]) );
  AND U16750 ( .A(p_input[22463]), .B(p_input[12463]), .Z(n8375) );
  AND U16751 ( .A(n8376), .B(p_input[2462]), .Z(o[2462]) );
  AND U16752 ( .A(p_input[22462]), .B(p_input[12462]), .Z(n8376) );
  AND U16753 ( .A(n8377), .B(p_input[2461]), .Z(o[2461]) );
  AND U16754 ( .A(p_input[22461]), .B(p_input[12461]), .Z(n8377) );
  AND U16755 ( .A(n8378), .B(p_input[2460]), .Z(o[2460]) );
  AND U16756 ( .A(p_input[22460]), .B(p_input[12460]), .Z(n8378) );
  AND U16757 ( .A(n8379), .B(p_input[245]), .Z(o[245]) );
  AND U16758 ( .A(p_input[20245]), .B(p_input[10245]), .Z(n8379) );
  AND U16759 ( .A(n8380), .B(p_input[2459]), .Z(o[2459]) );
  AND U16760 ( .A(p_input[22459]), .B(p_input[12459]), .Z(n8380) );
  AND U16761 ( .A(n8381), .B(p_input[2458]), .Z(o[2458]) );
  AND U16762 ( .A(p_input[22458]), .B(p_input[12458]), .Z(n8381) );
  AND U16763 ( .A(n8382), .B(p_input[2457]), .Z(o[2457]) );
  AND U16764 ( .A(p_input[22457]), .B(p_input[12457]), .Z(n8382) );
  AND U16765 ( .A(n8383), .B(p_input[2456]), .Z(o[2456]) );
  AND U16766 ( .A(p_input[22456]), .B(p_input[12456]), .Z(n8383) );
  AND U16767 ( .A(n8384), .B(p_input[2455]), .Z(o[2455]) );
  AND U16768 ( .A(p_input[22455]), .B(p_input[12455]), .Z(n8384) );
  AND U16769 ( .A(n8385), .B(p_input[2454]), .Z(o[2454]) );
  AND U16770 ( .A(p_input[22454]), .B(p_input[12454]), .Z(n8385) );
  AND U16771 ( .A(n8386), .B(p_input[2453]), .Z(o[2453]) );
  AND U16772 ( .A(p_input[22453]), .B(p_input[12453]), .Z(n8386) );
  AND U16773 ( .A(n8387), .B(p_input[2452]), .Z(o[2452]) );
  AND U16774 ( .A(p_input[22452]), .B(p_input[12452]), .Z(n8387) );
  AND U16775 ( .A(n8388), .B(p_input[2451]), .Z(o[2451]) );
  AND U16776 ( .A(p_input[22451]), .B(p_input[12451]), .Z(n8388) );
  AND U16777 ( .A(n8389), .B(p_input[2450]), .Z(o[2450]) );
  AND U16778 ( .A(p_input[22450]), .B(p_input[12450]), .Z(n8389) );
  AND U16779 ( .A(n8390), .B(p_input[244]), .Z(o[244]) );
  AND U16780 ( .A(p_input[20244]), .B(p_input[10244]), .Z(n8390) );
  AND U16781 ( .A(n8391), .B(p_input[2449]), .Z(o[2449]) );
  AND U16782 ( .A(p_input[22449]), .B(p_input[12449]), .Z(n8391) );
  AND U16783 ( .A(n8392), .B(p_input[2448]), .Z(o[2448]) );
  AND U16784 ( .A(p_input[22448]), .B(p_input[12448]), .Z(n8392) );
  AND U16785 ( .A(n8393), .B(p_input[2447]), .Z(o[2447]) );
  AND U16786 ( .A(p_input[22447]), .B(p_input[12447]), .Z(n8393) );
  AND U16787 ( .A(n8394), .B(p_input[2446]), .Z(o[2446]) );
  AND U16788 ( .A(p_input[22446]), .B(p_input[12446]), .Z(n8394) );
  AND U16789 ( .A(n8395), .B(p_input[2445]), .Z(o[2445]) );
  AND U16790 ( .A(p_input[22445]), .B(p_input[12445]), .Z(n8395) );
  AND U16791 ( .A(n8396), .B(p_input[2444]), .Z(o[2444]) );
  AND U16792 ( .A(p_input[22444]), .B(p_input[12444]), .Z(n8396) );
  AND U16793 ( .A(n8397), .B(p_input[2443]), .Z(o[2443]) );
  AND U16794 ( .A(p_input[22443]), .B(p_input[12443]), .Z(n8397) );
  AND U16795 ( .A(n8398), .B(p_input[2442]), .Z(o[2442]) );
  AND U16796 ( .A(p_input[22442]), .B(p_input[12442]), .Z(n8398) );
  AND U16797 ( .A(n8399), .B(p_input[2441]), .Z(o[2441]) );
  AND U16798 ( .A(p_input[22441]), .B(p_input[12441]), .Z(n8399) );
  AND U16799 ( .A(n8400), .B(p_input[2440]), .Z(o[2440]) );
  AND U16800 ( .A(p_input[22440]), .B(p_input[12440]), .Z(n8400) );
  AND U16801 ( .A(n8401), .B(p_input[243]), .Z(o[243]) );
  AND U16802 ( .A(p_input[20243]), .B(p_input[10243]), .Z(n8401) );
  AND U16803 ( .A(n8402), .B(p_input[2439]), .Z(o[2439]) );
  AND U16804 ( .A(p_input[22439]), .B(p_input[12439]), .Z(n8402) );
  AND U16805 ( .A(n8403), .B(p_input[2438]), .Z(o[2438]) );
  AND U16806 ( .A(p_input[22438]), .B(p_input[12438]), .Z(n8403) );
  AND U16807 ( .A(n8404), .B(p_input[2437]), .Z(o[2437]) );
  AND U16808 ( .A(p_input[22437]), .B(p_input[12437]), .Z(n8404) );
  AND U16809 ( .A(n8405), .B(p_input[2436]), .Z(o[2436]) );
  AND U16810 ( .A(p_input[22436]), .B(p_input[12436]), .Z(n8405) );
  AND U16811 ( .A(n8406), .B(p_input[2435]), .Z(o[2435]) );
  AND U16812 ( .A(p_input[22435]), .B(p_input[12435]), .Z(n8406) );
  AND U16813 ( .A(n8407), .B(p_input[2434]), .Z(o[2434]) );
  AND U16814 ( .A(p_input[22434]), .B(p_input[12434]), .Z(n8407) );
  AND U16815 ( .A(n8408), .B(p_input[2433]), .Z(o[2433]) );
  AND U16816 ( .A(p_input[22433]), .B(p_input[12433]), .Z(n8408) );
  AND U16817 ( .A(n8409), .B(p_input[2432]), .Z(o[2432]) );
  AND U16818 ( .A(p_input[22432]), .B(p_input[12432]), .Z(n8409) );
  AND U16819 ( .A(n8410), .B(p_input[2431]), .Z(o[2431]) );
  AND U16820 ( .A(p_input[22431]), .B(p_input[12431]), .Z(n8410) );
  AND U16821 ( .A(n8411), .B(p_input[2430]), .Z(o[2430]) );
  AND U16822 ( .A(p_input[22430]), .B(p_input[12430]), .Z(n8411) );
  AND U16823 ( .A(n8412), .B(p_input[242]), .Z(o[242]) );
  AND U16824 ( .A(p_input[20242]), .B(p_input[10242]), .Z(n8412) );
  AND U16825 ( .A(n8413), .B(p_input[2429]), .Z(o[2429]) );
  AND U16826 ( .A(p_input[22429]), .B(p_input[12429]), .Z(n8413) );
  AND U16827 ( .A(n8414), .B(p_input[2428]), .Z(o[2428]) );
  AND U16828 ( .A(p_input[22428]), .B(p_input[12428]), .Z(n8414) );
  AND U16829 ( .A(n8415), .B(p_input[2427]), .Z(o[2427]) );
  AND U16830 ( .A(p_input[22427]), .B(p_input[12427]), .Z(n8415) );
  AND U16831 ( .A(n8416), .B(p_input[2426]), .Z(o[2426]) );
  AND U16832 ( .A(p_input[22426]), .B(p_input[12426]), .Z(n8416) );
  AND U16833 ( .A(n8417), .B(p_input[2425]), .Z(o[2425]) );
  AND U16834 ( .A(p_input[22425]), .B(p_input[12425]), .Z(n8417) );
  AND U16835 ( .A(n8418), .B(p_input[2424]), .Z(o[2424]) );
  AND U16836 ( .A(p_input[22424]), .B(p_input[12424]), .Z(n8418) );
  AND U16837 ( .A(n8419), .B(p_input[2423]), .Z(o[2423]) );
  AND U16838 ( .A(p_input[22423]), .B(p_input[12423]), .Z(n8419) );
  AND U16839 ( .A(n8420), .B(p_input[2422]), .Z(o[2422]) );
  AND U16840 ( .A(p_input[22422]), .B(p_input[12422]), .Z(n8420) );
  AND U16841 ( .A(n8421), .B(p_input[2421]), .Z(o[2421]) );
  AND U16842 ( .A(p_input[22421]), .B(p_input[12421]), .Z(n8421) );
  AND U16843 ( .A(n8422), .B(p_input[2420]), .Z(o[2420]) );
  AND U16844 ( .A(p_input[22420]), .B(p_input[12420]), .Z(n8422) );
  AND U16845 ( .A(n8423), .B(p_input[241]), .Z(o[241]) );
  AND U16846 ( .A(p_input[20241]), .B(p_input[10241]), .Z(n8423) );
  AND U16847 ( .A(n8424), .B(p_input[2419]), .Z(o[2419]) );
  AND U16848 ( .A(p_input[22419]), .B(p_input[12419]), .Z(n8424) );
  AND U16849 ( .A(n8425), .B(p_input[2418]), .Z(o[2418]) );
  AND U16850 ( .A(p_input[22418]), .B(p_input[12418]), .Z(n8425) );
  AND U16851 ( .A(n8426), .B(p_input[2417]), .Z(o[2417]) );
  AND U16852 ( .A(p_input[22417]), .B(p_input[12417]), .Z(n8426) );
  AND U16853 ( .A(n8427), .B(p_input[2416]), .Z(o[2416]) );
  AND U16854 ( .A(p_input[22416]), .B(p_input[12416]), .Z(n8427) );
  AND U16855 ( .A(n8428), .B(p_input[2415]), .Z(o[2415]) );
  AND U16856 ( .A(p_input[22415]), .B(p_input[12415]), .Z(n8428) );
  AND U16857 ( .A(n8429), .B(p_input[2414]), .Z(o[2414]) );
  AND U16858 ( .A(p_input[22414]), .B(p_input[12414]), .Z(n8429) );
  AND U16859 ( .A(n8430), .B(p_input[2413]), .Z(o[2413]) );
  AND U16860 ( .A(p_input[22413]), .B(p_input[12413]), .Z(n8430) );
  AND U16861 ( .A(n8431), .B(p_input[2412]), .Z(o[2412]) );
  AND U16862 ( .A(p_input[22412]), .B(p_input[12412]), .Z(n8431) );
  AND U16863 ( .A(n8432), .B(p_input[2411]), .Z(o[2411]) );
  AND U16864 ( .A(p_input[22411]), .B(p_input[12411]), .Z(n8432) );
  AND U16865 ( .A(n8433), .B(p_input[2410]), .Z(o[2410]) );
  AND U16866 ( .A(p_input[22410]), .B(p_input[12410]), .Z(n8433) );
  AND U16867 ( .A(n8434), .B(p_input[240]), .Z(o[240]) );
  AND U16868 ( .A(p_input[20240]), .B(p_input[10240]), .Z(n8434) );
  AND U16869 ( .A(n8435), .B(p_input[2409]), .Z(o[2409]) );
  AND U16870 ( .A(p_input[22409]), .B(p_input[12409]), .Z(n8435) );
  AND U16871 ( .A(n8436), .B(p_input[2408]), .Z(o[2408]) );
  AND U16872 ( .A(p_input[22408]), .B(p_input[12408]), .Z(n8436) );
  AND U16873 ( .A(n8437), .B(p_input[2407]), .Z(o[2407]) );
  AND U16874 ( .A(p_input[22407]), .B(p_input[12407]), .Z(n8437) );
  AND U16875 ( .A(n8438), .B(p_input[2406]), .Z(o[2406]) );
  AND U16876 ( .A(p_input[22406]), .B(p_input[12406]), .Z(n8438) );
  AND U16877 ( .A(n8439), .B(p_input[2405]), .Z(o[2405]) );
  AND U16878 ( .A(p_input[22405]), .B(p_input[12405]), .Z(n8439) );
  AND U16879 ( .A(n8440), .B(p_input[2404]), .Z(o[2404]) );
  AND U16880 ( .A(p_input[22404]), .B(p_input[12404]), .Z(n8440) );
  AND U16881 ( .A(n8441), .B(p_input[2403]), .Z(o[2403]) );
  AND U16882 ( .A(p_input[22403]), .B(p_input[12403]), .Z(n8441) );
  AND U16883 ( .A(n8442), .B(p_input[2402]), .Z(o[2402]) );
  AND U16884 ( .A(p_input[22402]), .B(p_input[12402]), .Z(n8442) );
  AND U16885 ( .A(n8443), .B(p_input[2401]), .Z(o[2401]) );
  AND U16886 ( .A(p_input[22401]), .B(p_input[12401]), .Z(n8443) );
  AND U16887 ( .A(n8444), .B(p_input[2400]), .Z(o[2400]) );
  AND U16888 ( .A(p_input[22400]), .B(p_input[12400]), .Z(n8444) );
  AND U16889 ( .A(n8445), .B(p_input[23]), .Z(o[23]) );
  AND U16890 ( .A(p_input[20023]), .B(p_input[10023]), .Z(n8445) );
  AND U16891 ( .A(n8446), .B(p_input[239]), .Z(o[239]) );
  AND U16892 ( .A(p_input[20239]), .B(p_input[10239]), .Z(n8446) );
  AND U16893 ( .A(n8447), .B(p_input[2399]), .Z(o[2399]) );
  AND U16894 ( .A(p_input[22399]), .B(p_input[12399]), .Z(n8447) );
  AND U16895 ( .A(n8448), .B(p_input[2398]), .Z(o[2398]) );
  AND U16896 ( .A(p_input[22398]), .B(p_input[12398]), .Z(n8448) );
  AND U16897 ( .A(n8449), .B(p_input[2397]), .Z(o[2397]) );
  AND U16898 ( .A(p_input[22397]), .B(p_input[12397]), .Z(n8449) );
  AND U16899 ( .A(n8450), .B(p_input[2396]), .Z(o[2396]) );
  AND U16900 ( .A(p_input[22396]), .B(p_input[12396]), .Z(n8450) );
  AND U16901 ( .A(n8451), .B(p_input[2395]), .Z(o[2395]) );
  AND U16902 ( .A(p_input[22395]), .B(p_input[12395]), .Z(n8451) );
  AND U16903 ( .A(n8452), .B(p_input[2394]), .Z(o[2394]) );
  AND U16904 ( .A(p_input[22394]), .B(p_input[12394]), .Z(n8452) );
  AND U16905 ( .A(n8453), .B(p_input[2393]), .Z(o[2393]) );
  AND U16906 ( .A(p_input[22393]), .B(p_input[12393]), .Z(n8453) );
  AND U16907 ( .A(n8454), .B(p_input[2392]), .Z(o[2392]) );
  AND U16908 ( .A(p_input[22392]), .B(p_input[12392]), .Z(n8454) );
  AND U16909 ( .A(n8455), .B(p_input[2391]), .Z(o[2391]) );
  AND U16910 ( .A(p_input[22391]), .B(p_input[12391]), .Z(n8455) );
  AND U16911 ( .A(n8456), .B(p_input[2390]), .Z(o[2390]) );
  AND U16912 ( .A(p_input[22390]), .B(p_input[12390]), .Z(n8456) );
  AND U16913 ( .A(n8457), .B(p_input[238]), .Z(o[238]) );
  AND U16914 ( .A(p_input[20238]), .B(p_input[10238]), .Z(n8457) );
  AND U16915 ( .A(n8458), .B(p_input[2389]), .Z(o[2389]) );
  AND U16916 ( .A(p_input[22389]), .B(p_input[12389]), .Z(n8458) );
  AND U16917 ( .A(n8459), .B(p_input[2388]), .Z(o[2388]) );
  AND U16918 ( .A(p_input[22388]), .B(p_input[12388]), .Z(n8459) );
  AND U16919 ( .A(n8460), .B(p_input[2387]), .Z(o[2387]) );
  AND U16920 ( .A(p_input[22387]), .B(p_input[12387]), .Z(n8460) );
  AND U16921 ( .A(n8461), .B(p_input[2386]), .Z(o[2386]) );
  AND U16922 ( .A(p_input[22386]), .B(p_input[12386]), .Z(n8461) );
  AND U16923 ( .A(n8462), .B(p_input[2385]), .Z(o[2385]) );
  AND U16924 ( .A(p_input[22385]), .B(p_input[12385]), .Z(n8462) );
  AND U16925 ( .A(n8463), .B(p_input[2384]), .Z(o[2384]) );
  AND U16926 ( .A(p_input[22384]), .B(p_input[12384]), .Z(n8463) );
  AND U16927 ( .A(n8464), .B(p_input[2383]), .Z(o[2383]) );
  AND U16928 ( .A(p_input[22383]), .B(p_input[12383]), .Z(n8464) );
  AND U16929 ( .A(n8465), .B(p_input[2382]), .Z(o[2382]) );
  AND U16930 ( .A(p_input[22382]), .B(p_input[12382]), .Z(n8465) );
  AND U16931 ( .A(n8466), .B(p_input[2381]), .Z(o[2381]) );
  AND U16932 ( .A(p_input[22381]), .B(p_input[12381]), .Z(n8466) );
  AND U16933 ( .A(n8467), .B(p_input[2380]), .Z(o[2380]) );
  AND U16934 ( .A(p_input[22380]), .B(p_input[12380]), .Z(n8467) );
  AND U16935 ( .A(n8468), .B(p_input[237]), .Z(o[237]) );
  AND U16936 ( .A(p_input[20237]), .B(p_input[10237]), .Z(n8468) );
  AND U16937 ( .A(n8469), .B(p_input[2379]), .Z(o[2379]) );
  AND U16938 ( .A(p_input[22379]), .B(p_input[12379]), .Z(n8469) );
  AND U16939 ( .A(n8470), .B(p_input[2378]), .Z(o[2378]) );
  AND U16940 ( .A(p_input[22378]), .B(p_input[12378]), .Z(n8470) );
  AND U16941 ( .A(n8471), .B(p_input[2377]), .Z(o[2377]) );
  AND U16942 ( .A(p_input[22377]), .B(p_input[12377]), .Z(n8471) );
  AND U16943 ( .A(n8472), .B(p_input[2376]), .Z(o[2376]) );
  AND U16944 ( .A(p_input[22376]), .B(p_input[12376]), .Z(n8472) );
  AND U16945 ( .A(n8473), .B(p_input[2375]), .Z(o[2375]) );
  AND U16946 ( .A(p_input[22375]), .B(p_input[12375]), .Z(n8473) );
  AND U16947 ( .A(n8474), .B(p_input[2374]), .Z(o[2374]) );
  AND U16948 ( .A(p_input[22374]), .B(p_input[12374]), .Z(n8474) );
  AND U16949 ( .A(n8475), .B(p_input[2373]), .Z(o[2373]) );
  AND U16950 ( .A(p_input[22373]), .B(p_input[12373]), .Z(n8475) );
  AND U16951 ( .A(n8476), .B(p_input[2372]), .Z(o[2372]) );
  AND U16952 ( .A(p_input[22372]), .B(p_input[12372]), .Z(n8476) );
  AND U16953 ( .A(n8477), .B(p_input[2371]), .Z(o[2371]) );
  AND U16954 ( .A(p_input[22371]), .B(p_input[12371]), .Z(n8477) );
  AND U16955 ( .A(n8478), .B(p_input[2370]), .Z(o[2370]) );
  AND U16956 ( .A(p_input[22370]), .B(p_input[12370]), .Z(n8478) );
  AND U16957 ( .A(n8479), .B(p_input[236]), .Z(o[236]) );
  AND U16958 ( .A(p_input[20236]), .B(p_input[10236]), .Z(n8479) );
  AND U16959 ( .A(n8480), .B(p_input[2369]), .Z(o[2369]) );
  AND U16960 ( .A(p_input[22369]), .B(p_input[12369]), .Z(n8480) );
  AND U16961 ( .A(n8481), .B(p_input[2368]), .Z(o[2368]) );
  AND U16962 ( .A(p_input[22368]), .B(p_input[12368]), .Z(n8481) );
  AND U16963 ( .A(n8482), .B(p_input[2367]), .Z(o[2367]) );
  AND U16964 ( .A(p_input[22367]), .B(p_input[12367]), .Z(n8482) );
  AND U16965 ( .A(n8483), .B(p_input[2366]), .Z(o[2366]) );
  AND U16966 ( .A(p_input[22366]), .B(p_input[12366]), .Z(n8483) );
  AND U16967 ( .A(n8484), .B(p_input[2365]), .Z(o[2365]) );
  AND U16968 ( .A(p_input[22365]), .B(p_input[12365]), .Z(n8484) );
  AND U16969 ( .A(n8485), .B(p_input[2364]), .Z(o[2364]) );
  AND U16970 ( .A(p_input[22364]), .B(p_input[12364]), .Z(n8485) );
  AND U16971 ( .A(n8486), .B(p_input[2363]), .Z(o[2363]) );
  AND U16972 ( .A(p_input[22363]), .B(p_input[12363]), .Z(n8486) );
  AND U16973 ( .A(n8487), .B(p_input[2362]), .Z(o[2362]) );
  AND U16974 ( .A(p_input[22362]), .B(p_input[12362]), .Z(n8487) );
  AND U16975 ( .A(n8488), .B(p_input[2361]), .Z(o[2361]) );
  AND U16976 ( .A(p_input[22361]), .B(p_input[12361]), .Z(n8488) );
  AND U16977 ( .A(n8489), .B(p_input[2360]), .Z(o[2360]) );
  AND U16978 ( .A(p_input[22360]), .B(p_input[12360]), .Z(n8489) );
  AND U16979 ( .A(n8490), .B(p_input[235]), .Z(o[235]) );
  AND U16980 ( .A(p_input[20235]), .B(p_input[10235]), .Z(n8490) );
  AND U16981 ( .A(n8491), .B(p_input[2359]), .Z(o[2359]) );
  AND U16982 ( .A(p_input[22359]), .B(p_input[12359]), .Z(n8491) );
  AND U16983 ( .A(n8492), .B(p_input[2358]), .Z(o[2358]) );
  AND U16984 ( .A(p_input[22358]), .B(p_input[12358]), .Z(n8492) );
  AND U16985 ( .A(n8493), .B(p_input[2357]), .Z(o[2357]) );
  AND U16986 ( .A(p_input[22357]), .B(p_input[12357]), .Z(n8493) );
  AND U16987 ( .A(n8494), .B(p_input[2356]), .Z(o[2356]) );
  AND U16988 ( .A(p_input[22356]), .B(p_input[12356]), .Z(n8494) );
  AND U16989 ( .A(n8495), .B(p_input[2355]), .Z(o[2355]) );
  AND U16990 ( .A(p_input[22355]), .B(p_input[12355]), .Z(n8495) );
  AND U16991 ( .A(n8496), .B(p_input[2354]), .Z(o[2354]) );
  AND U16992 ( .A(p_input[22354]), .B(p_input[12354]), .Z(n8496) );
  AND U16993 ( .A(n8497), .B(p_input[2353]), .Z(o[2353]) );
  AND U16994 ( .A(p_input[22353]), .B(p_input[12353]), .Z(n8497) );
  AND U16995 ( .A(n8498), .B(p_input[2352]), .Z(o[2352]) );
  AND U16996 ( .A(p_input[22352]), .B(p_input[12352]), .Z(n8498) );
  AND U16997 ( .A(n8499), .B(p_input[2351]), .Z(o[2351]) );
  AND U16998 ( .A(p_input[22351]), .B(p_input[12351]), .Z(n8499) );
  AND U16999 ( .A(n8500), .B(p_input[2350]), .Z(o[2350]) );
  AND U17000 ( .A(p_input[22350]), .B(p_input[12350]), .Z(n8500) );
  AND U17001 ( .A(n8501), .B(p_input[234]), .Z(o[234]) );
  AND U17002 ( .A(p_input[20234]), .B(p_input[10234]), .Z(n8501) );
  AND U17003 ( .A(n8502), .B(p_input[2349]), .Z(o[2349]) );
  AND U17004 ( .A(p_input[22349]), .B(p_input[12349]), .Z(n8502) );
  AND U17005 ( .A(n8503), .B(p_input[2348]), .Z(o[2348]) );
  AND U17006 ( .A(p_input[22348]), .B(p_input[12348]), .Z(n8503) );
  AND U17007 ( .A(n8504), .B(p_input[2347]), .Z(o[2347]) );
  AND U17008 ( .A(p_input[22347]), .B(p_input[12347]), .Z(n8504) );
  AND U17009 ( .A(n8505), .B(p_input[2346]), .Z(o[2346]) );
  AND U17010 ( .A(p_input[22346]), .B(p_input[12346]), .Z(n8505) );
  AND U17011 ( .A(n8506), .B(p_input[2345]), .Z(o[2345]) );
  AND U17012 ( .A(p_input[22345]), .B(p_input[12345]), .Z(n8506) );
  AND U17013 ( .A(n8507), .B(p_input[2344]), .Z(o[2344]) );
  AND U17014 ( .A(p_input[22344]), .B(p_input[12344]), .Z(n8507) );
  AND U17015 ( .A(n8508), .B(p_input[2343]), .Z(o[2343]) );
  AND U17016 ( .A(p_input[22343]), .B(p_input[12343]), .Z(n8508) );
  AND U17017 ( .A(n8509), .B(p_input[2342]), .Z(o[2342]) );
  AND U17018 ( .A(p_input[22342]), .B(p_input[12342]), .Z(n8509) );
  AND U17019 ( .A(n8510), .B(p_input[2341]), .Z(o[2341]) );
  AND U17020 ( .A(p_input[22341]), .B(p_input[12341]), .Z(n8510) );
  AND U17021 ( .A(n8511), .B(p_input[2340]), .Z(o[2340]) );
  AND U17022 ( .A(p_input[22340]), .B(p_input[12340]), .Z(n8511) );
  AND U17023 ( .A(n8512), .B(p_input[233]), .Z(o[233]) );
  AND U17024 ( .A(p_input[20233]), .B(p_input[10233]), .Z(n8512) );
  AND U17025 ( .A(n8513), .B(p_input[2339]), .Z(o[2339]) );
  AND U17026 ( .A(p_input[22339]), .B(p_input[12339]), .Z(n8513) );
  AND U17027 ( .A(n8514), .B(p_input[2338]), .Z(o[2338]) );
  AND U17028 ( .A(p_input[22338]), .B(p_input[12338]), .Z(n8514) );
  AND U17029 ( .A(n8515), .B(p_input[2337]), .Z(o[2337]) );
  AND U17030 ( .A(p_input[22337]), .B(p_input[12337]), .Z(n8515) );
  AND U17031 ( .A(n8516), .B(p_input[2336]), .Z(o[2336]) );
  AND U17032 ( .A(p_input[22336]), .B(p_input[12336]), .Z(n8516) );
  AND U17033 ( .A(n8517), .B(p_input[2335]), .Z(o[2335]) );
  AND U17034 ( .A(p_input[22335]), .B(p_input[12335]), .Z(n8517) );
  AND U17035 ( .A(n8518), .B(p_input[2334]), .Z(o[2334]) );
  AND U17036 ( .A(p_input[22334]), .B(p_input[12334]), .Z(n8518) );
  AND U17037 ( .A(n8519), .B(p_input[2333]), .Z(o[2333]) );
  AND U17038 ( .A(p_input[22333]), .B(p_input[12333]), .Z(n8519) );
  AND U17039 ( .A(n8520), .B(p_input[2332]), .Z(o[2332]) );
  AND U17040 ( .A(p_input[22332]), .B(p_input[12332]), .Z(n8520) );
  AND U17041 ( .A(n8521), .B(p_input[2331]), .Z(o[2331]) );
  AND U17042 ( .A(p_input[22331]), .B(p_input[12331]), .Z(n8521) );
  AND U17043 ( .A(n8522), .B(p_input[2330]), .Z(o[2330]) );
  AND U17044 ( .A(p_input[22330]), .B(p_input[12330]), .Z(n8522) );
  AND U17045 ( .A(n8523), .B(p_input[232]), .Z(o[232]) );
  AND U17046 ( .A(p_input[20232]), .B(p_input[10232]), .Z(n8523) );
  AND U17047 ( .A(n8524), .B(p_input[2329]), .Z(o[2329]) );
  AND U17048 ( .A(p_input[22329]), .B(p_input[12329]), .Z(n8524) );
  AND U17049 ( .A(n8525), .B(p_input[2328]), .Z(o[2328]) );
  AND U17050 ( .A(p_input[22328]), .B(p_input[12328]), .Z(n8525) );
  AND U17051 ( .A(n8526), .B(p_input[2327]), .Z(o[2327]) );
  AND U17052 ( .A(p_input[22327]), .B(p_input[12327]), .Z(n8526) );
  AND U17053 ( .A(n8527), .B(p_input[2326]), .Z(o[2326]) );
  AND U17054 ( .A(p_input[22326]), .B(p_input[12326]), .Z(n8527) );
  AND U17055 ( .A(n8528), .B(p_input[2325]), .Z(o[2325]) );
  AND U17056 ( .A(p_input[22325]), .B(p_input[12325]), .Z(n8528) );
  AND U17057 ( .A(n8529), .B(p_input[2324]), .Z(o[2324]) );
  AND U17058 ( .A(p_input[22324]), .B(p_input[12324]), .Z(n8529) );
  AND U17059 ( .A(n8530), .B(p_input[2323]), .Z(o[2323]) );
  AND U17060 ( .A(p_input[22323]), .B(p_input[12323]), .Z(n8530) );
  AND U17061 ( .A(n8531), .B(p_input[2322]), .Z(o[2322]) );
  AND U17062 ( .A(p_input[22322]), .B(p_input[12322]), .Z(n8531) );
  AND U17063 ( .A(n8532), .B(p_input[2321]), .Z(o[2321]) );
  AND U17064 ( .A(p_input[22321]), .B(p_input[12321]), .Z(n8532) );
  AND U17065 ( .A(n8533), .B(p_input[2320]), .Z(o[2320]) );
  AND U17066 ( .A(p_input[22320]), .B(p_input[12320]), .Z(n8533) );
  AND U17067 ( .A(n8534), .B(p_input[231]), .Z(o[231]) );
  AND U17068 ( .A(p_input[20231]), .B(p_input[10231]), .Z(n8534) );
  AND U17069 ( .A(n8535), .B(p_input[2319]), .Z(o[2319]) );
  AND U17070 ( .A(p_input[22319]), .B(p_input[12319]), .Z(n8535) );
  AND U17071 ( .A(n8536), .B(p_input[2318]), .Z(o[2318]) );
  AND U17072 ( .A(p_input[22318]), .B(p_input[12318]), .Z(n8536) );
  AND U17073 ( .A(n8537), .B(p_input[2317]), .Z(o[2317]) );
  AND U17074 ( .A(p_input[22317]), .B(p_input[12317]), .Z(n8537) );
  AND U17075 ( .A(n8538), .B(p_input[2316]), .Z(o[2316]) );
  AND U17076 ( .A(p_input[22316]), .B(p_input[12316]), .Z(n8538) );
  AND U17077 ( .A(n8539), .B(p_input[2315]), .Z(o[2315]) );
  AND U17078 ( .A(p_input[22315]), .B(p_input[12315]), .Z(n8539) );
  AND U17079 ( .A(n8540), .B(p_input[2314]), .Z(o[2314]) );
  AND U17080 ( .A(p_input[22314]), .B(p_input[12314]), .Z(n8540) );
  AND U17081 ( .A(n8541), .B(p_input[2313]), .Z(o[2313]) );
  AND U17082 ( .A(p_input[22313]), .B(p_input[12313]), .Z(n8541) );
  AND U17083 ( .A(n8542), .B(p_input[2312]), .Z(o[2312]) );
  AND U17084 ( .A(p_input[22312]), .B(p_input[12312]), .Z(n8542) );
  AND U17085 ( .A(n8543), .B(p_input[2311]), .Z(o[2311]) );
  AND U17086 ( .A(p_input[22311]), .B(p_input[12311]), .Z(n8543) );
  AND U17087 ( .A(n8544), .B(p_input[2310]), .Z(o[2310]) );
  AND U17088 ( .A(p_input[22310]), .B(p_input[12310]), .Z(n8544) );
  AND U17089 ( .A(n8545), .B(p_input[230]), .Z(o[230]) );
  AND U17090 ( .A(p_input[20230]), .B(p_input[10230]), .Z(n8545) );
  AND U17091 ( .A(n8546), .B(p_input[2309]), .Z(o[2309]) );
  AND U17092 ( .A(p_input[22309]), .B(p_input[12309]), .Z(n8546) );
  AND U17093 ( .A(n8547), .B(p_input[2308]), .Z(o[2308]) );
  AND U17094 ( .A(p_input[22308]), .B(p_input[12308]), .Z(n8547) );
  AND U17095 ( .A(n8548), .B(p_input[2307]), .Z(o[2307]) );
  AND U17096 ( .A(p_input[22307]), .B(p_input[12307]), .Z(n8548) );
  AND U17097 ( .A(n8549), .B(p_input[2306]), .Z(o[2306]) );
  AND U17098 ( .A(p_input[22306]), .B(p_input[12306]), .Z(n8549) );
  AND U17099 ( .A(n8550), .B(p_input[2305]), .Z(o[2305]) );
  AND U17100 ( .A(p_input[22305]), .B(p_input[12305]), .Z(n8550) );
  AND U17101 ( .A(n8551), .B(p_input[2304]), .Z(o[2304]) );
  AND U17102 ( .A(p_input[22304]), .B(p_input[12304]), .Z(n8551) );
  AND U17103 ( .A(n8552), .B(p_input[2303]), .Z(o[2303]) );
  AND U17104 ( .A(p_input[22303]), .B(p_input[12303]), .Z(n8552) );
  AND U17105 ( .A(n8553), .B(p_input[2302]), .Z(o[2302]) );
  AND U17106 ( .A(p_input[22302]), .B(p_input[12302]), .Z(n8553) );
  AND U17107 ( .A(n8554), .B(p_input[2301]), .Z(o[2301]) );
  AND U17108 ( .A(p_input[22301]), .B(p_input[12301]), .Z(n8554) );
  AND U17109 ( .A(n8555), .B(p_input[2300]), .Z(o[2300]) );
  AND U17110 ( .A(p_input[22300]), .B(p_input[12300]), .Z(n8555) );
  AND U17111 ( .A(n8556), .B(p_input[22]), .Z(o[22]) );
  AND U17112 ( .A(p_input[20022]), .B(p_input[10022]), .Z(n8556) );
  AND U17113 ( .A(n8557), .B(p_input[229]), .Z(o[229]) );
  AND U17114 ( .A(p_input[20229]), .B(p_input[10229]), .Z(n8557) );
  AND U17115 ( .A(n8558), .B(p_input[2299]), .Z(o[2299]) );
  AND U17116 ( .A(p_input[22299]), .B(p_input[12299]), .Z(n8558) );
  AND U17117 ( .A(n8559), .B(p_input[2298]), .Z(o[2298]) );
  AND U17118 ( .A(p_input[22298]), .B(p_input[12298]), .Z(n8559) );
  AND U17119 ( .A(n8560), .B(p_input[2297]), .Z(o[2297]) );
  AND U17120 ( .A(p_input[22297]), .B(p_input[12297]), .Z(n8560) );
  AND U17121 ( .A(n8561), .B(p_input[2296]), .Z(o[2296]) );
  AND U17122 ( .A(p_input[22296]), .B(p_input[12296]), .Z(n8561) );
  AND U17123 ( .A(n8562), .B(p_input[2295]), .Z(o[2295]) );
  AND U17124 ( .A(p_input[22295]), .B(p_input[12295]), .Z(n8562) );
  AND U17125 ( .A(n8563), .B(p_input[2294]), .Z(o[2294]) );
  AND U17126 ( .A(p_input[22294]), .B(p_input[12294]), .Z(n8563) );
  AND U17127 ( .A(n8564), .B(p_input[2293]), .Z(o[2293]) );
  AND U17128 ( .A(p_input[22293]), .B(p_input[12293]), .Z(n8564) );
  AND U17129 ( .A(n8565), .B(p_input[2292]), .Z(o[2292]) );
  AND U17130 ( .A(p_input[22292]), .B(p_input[12292]), .Z(n8565) );
  AND U17131 ( .A(n8566), .B(p_input[2291]), .Z(o[2291]) );
  AND U17132 ( .A(p_input[22291]), .B(p_input[12291]), .Z(n8566) );
  AND U17133 ( .A(n8567), .B(p_input[2290]), .Z(o[2290]) );
  AND U17134 ( .A(p_input[22290]), .B(p_input[12290]), .Z(n8567) );
  AND U17135 ( .A(n8568), .B(p_input[228]), .Z(o[228]) );
  AND U17136 ( .A(p_input[20228]), .B(p_input[10228]), .Z(n8568) );
  AND U17137 ( .A(n8569), .B(p_input[2289]), .Z(o[2289]) );
  AND U17138 ( .A(p_input[22289]), .B(p_input[12289]), .Z(n8569) );
  AND U17139 ( .A(n8570), .B(p_input[2288]), .Z(o[2288]) );
  AND U17140 ( .A(p_input[22288]), .B(p_input[12288]), .Z(n8570) );
  AND U17141 ( .A(n8571), .B(p_input[2287]), .Z(o[2287]) );
  AND U17142 ( .A(p_input[22287]), .B(p_input[12287]), .Z(n8571) );
  AND U17143 ( .A(n8572), .B(p_input[2286]), .Z(o[2286]) );
  AND U17144 ( .A(p_input[22286]), .B(p_input[12286]), .Z(n8572) );
  AND U17145 ( .A(n8573), .B(p_input[2285]), .Z(o[2285]) );
  AND U17146 ( .A(p_input[22285]), .B(p_input[12285]), .Z(n8573) );
  AND U17147 ( .A(n8574), .B(p_input[2284]), .Z(o[2284]) );
  AND U17148 ( .A(p_input[22284]), .B(p_input[12284]), .Z(n8574) );
  AND U17149 ( .A(n8575), .B(p_input[2283]), .Z(o[2283]) );
  AND U17150 ( .A(p_input[22283]), .B(p_input[12283]), .Z(n8575) );
  AND U17151 ( .A(n8576), .B(p_input[2282]), .Z(o[2282]) );
  AND U17152 ( .A(p_input[22282]), .B(p_input[12282]), .Z(n8576) );
  AND U17153 ( .A(n8577), .B(p_input[2281]), .Z(o[2281]) );
  AND U17154 ( .A(p_input[22281]), .B(p_input[12281]), .Z(n8577) );
  AND U17155 ( .A(n8578), .B(p_input[2280]), .Z(o[2280]) );
  AND U17156 ( .A(p_input[22280]), .B(p_input[12280]), .Z(n8578) );
  AND U17157 ( .A(n8579), .B(p_input[227]), .Z(o[227]) );
  AND U17158 ( .A(p_input[20227]), .B(p_input[10227]), .Z(n8579) );
  AND U17159 ( .A(n8580), .B(p_input[2279]), .Z(o[2279]) );
  AND U17160 ( .A(p_input[22279]), .B(p_input[12279]), .Z(n8580) );
  AND U17161 ( .A(n8581), .B(p_input[2278]), .Z(o[2278]) );
  AND U17162 ( .A(p_input[22278]), .B(p_input[12278]), .Z(n8581) );
  AND U17163 ( .A(n8582), .B(p_input[2277]), .Z(o[2277]) );
  AND U17164 ( .A(p_input[22277]), .B(p_input[12277]), .Z(n8582) );
  AND U17165 ( .A(n8583), .B(p_input[2276]), .Z(o[2276]) );
  AND U17166 ( .A(p_input[22276]), .B(p_input[12276]), .Z(n8583) );
  AND U17167 ( .A(n8584), .B(p_input[2275]), .Z(o[2275]) );
  AND U17168 ( .A(p_input[22275]), .B(p_input[12275]), .Z(n8584) );
  AND U17169 ( .A(n8585), .B(p_input[2274]), .Z(o[2274]) );
  AND U17170 ( .A(p_input[22274]), .B(p_input[12274]), .Z(n8585) );
  AND U17171 ( .A(n8586), .B(p_input[2273]), .Z(o[2273]) );
  AND U17172 ( .A(p_input[22273]), .B(p_input[12273]), .Z(n8586) );
  AND U17173 ( .A(n8587), .B(p_input[2272]), .Z(o[2272]) );
  AND U17174 ( .A(p_input[22272]), .B(p_input[12272]), .Z(n8587) );
  AND U17175 ( .A(n8588), .B(p_input[2271]), .Z(o[2271]) );
  AND U17176 ( .A(p_input[22271]), .B(p_input[12271]), .Z(n8588) );
  AND U17177 ( .A(n8589), .B(p_input[2270]), .Z(o[2270]) );
  AND U17178 ( .A(p_input[22270]), .B(p_input[12270]), .Z(n8589) );
  AND U17179 ( .A(n8590), .B(p_input[226]), .Z(o[226]) );
  AND U17180 ( .A(p_input[20226]), .B(p_input[10226]), .Z(n8590) );
  AND U17181 ( .A(n8591), .B(p_input[2269]), .Z(o[2269]) );
  AND U17182 ( .A(p_input[22269]), .B(p_input[12269]), .Z(n8591) );
  AND U17183 ( .A(n8592), .B(p_input[2268]), .Z(o[2268]) );
  AND U17184 ( .A(p_input[22268]), .B(p_input[12268]), .Z(n8592) );
  AND U17185 ( .A(n8593), .B(p_input[2267]), .Z(o[2267]) );
  AND U17186 ( .A(p_input[22267]), .B(p_input[12267]), .Z(n8593) );
  AND U17187 ( .A(n8594), .B(p_input[2266]), .Z(o[2266]) );
  AND U17188 ( .A(p_input[22266]), .B(p_input[12266]), .Z(n8594) );
  AND U17189 ( .A(n8595), .B(p_input[2265]), .Z(o[2265]) );
  AND U17190 ( .A(p_input[22265]), .B(p_input[12265]), .Z(n8595) );
  AND U17191 ( .A(n8596), .B(p_input[2264]), .Z(o[2264]) );
  AND U17192 ( .A(p_input[22264]), .B(p_input[12264]), .Z(n8596) );
  AND U17193 ( .A(n8597), .B(p_input[2263]), .Z(o[2263]) );
  AND U17194 ( .A(p_input[22263]), .B(p_input[12263]), .Z(n8597) );
  AND U17195 ( .A(n8598), .B(p_input[2262]), .Z(o[2262]) );
  AND U17196 ( .A(p_input[22262]), .B(p_input[12262]), .Z(n8598) );
  AND U17197 ( .A(n8599), .B(p_input[2261]), .Z(o[2261]) );
  AND U17198 ( .A(p_input[22261]), .B(p_input[12261]), .Z(n8599) );
  AND U17199 ( .A(n8600), .B(p_input[2260]), .Z(o[2260]) );
  AND U17200 ( .A(p_input[22260]), .B(p_input[12260]), .Z(n8600) );
  AND U17201 ( .A(n8601), .B(p_input[225]), .Z(o[225]) );
  AND U17202 ( .A(p_input[20225]), .B(p_input[10225]), .Z(n8601) );
  AND U17203 ( .A(n8602), .B(p_input[2259]), .Z(o[2259]) );
  AND U17204 ( .A(p_input[22259]), .B(p_input[12259]), .Z(n8602) );
  AND U17205 ( .A(n8603), .B(p_input[2258]), .Z(o[2258]) );
  AND U17206 ( .A(p_input[22258]), .B(p_input[12258]), .Z(n8603) );
  AND U17207 ( .A(n8604), .B(p_input[2257]), .Z(o[2257]) );
  AND U17208 ( .A(p_input[22257]), .B(p_input[12257]), .Z(n8604) );
  AND U17209 ( .A(n8605), .B(p_input[2256]), .Z(o[2256]) );
  AND U17210 ( .A(p_input[22256]), .B(p_input[12256]), .Z(n8605) );
  AND U17211 ( .A(n8606), .B(p_input[2255]), .Z(o[2255]) );
  AND U17212 ( .A(p_input[22255]), .B(p_input[12255]), .Z(n8606) );
  AND U17213 ( .A(n8607), .B(p_input[2254]), .Z(o[2254]) );
  AND U17214 ( .A(p_input[22254]), .B(p_input[12254]), .Z(n8607) );
  AND U17215 ( .A(n8608), .B(p_input[2253]), .Z(o[2253]) );
  AND U17216 ( .A(p_input[22253]), .B(p_input[12253]), .Z(n8608) );
  AND U17217 ( .A(n8609), .B(p_input[2252]), .Z(o[2252]) );
  AND U17218 ( .A(p_input[22252]), .B(p_input[12252]), .Z(n8609) );
  AND U17219 ( .A(n8610), .B(p_input[2251]), .Z(o[2251]) );
  AND U17220 ( .A(p_input[22251]), .B(p_input[12251]), .Z(n8610) );
  AND U17221 ( .A(n8611), .B(p_input[2250]), .Z(o[2250]) );
  AND U17222 ( .A(p_input[22250]), .B(p_input[12250]), .Z(n8611) );
  AND U17223 ( .A(n8612), .B(p_input[224]), .Z(o[224]) );
  AND U17224 ( .A(p_input[20224]), .B(p_input[10224]), .Z(n8612) );
  AND U17225 ( .A(n8613), .B(p_input[2249]), .Z(o[2249]) );
  AND U17226 ( .A(p_input[22249]), .B(p_input[12249]), .Z(n8613) );
  AND U17227 ( .A(n8614), .B(p_input[2248]), .Z(o[2248]) );
  AND U17228 ( .A(p_input[22248]), .B(p_input[12248]), .Z(n8614) );
  AND U17229 ( .A(n8615), .B(p_input[2247]), .Z(o[2247]) );
  AND U17230 ( .A(p_input[22247]), .B(p_input[12247]), .Z(n8615) );
  AND U17231 ( .A(n8616), .B(p_input[2246]), .Z(o[2246]) );
  AND U17232 ( .A(p_input[22246]), .B(p_input[12246]), .Z(n8616) );
  AND U17233 ( .A(n8617), .B(p_input[2245]), .Z(o[2245]) );
  AND U17234 ( .A(p_input[22245]), .B(p_input[12245]), .Z(n8617) );
  AND U17235 ( .A(n8618), .B(p_input[2244]), .Z(o[2244]) );
  AND U17236 ( .A(p_input[22244]), .B(p_input[12244]), .Z(n8618) );
  AND U17237 ( .A(n8619), .B(p_input[2243]), .Z(o[2243]) );
  AND U17238 ( .A(p_input[22243]), .B(p_input[12243]), .Z(n8619) );
  AND U17239 ( .A(n8620), .B(p_input[2242]), .Z(o[2242]) );
  AND U17240 ( .A(p_input[22242]), .B(p_input[12242]), .Z(n8620) );
  AND U17241 ( .A(n8621), .B(p_input[2241]), .Z(o[2241]) );
  AND U17242 ( .A(p_input[22241]), .B(p_input[12241]), .Z(n8621) );
  AND U17243 ( .A(n8622), .B(p_input[2240]), .Z(o[2240]) );
  AND U17244 ( .A(p_input[22240]), .B(p_input[12240]), .Z(n8622) );
  AND U17245 ( .A(n8623), .B(p_input[223]), .Z(o[223]) );
  AND U17246 ( .A(p_input[20223]), .B(p_input[10223]), .Z(n8623) );
  AND U17247 ( .A(n8624), .B(p_input[2239]), .Z(o[2239]) );
  AND U17248 ( .A(p_input[22239]), .B(p_input[12239]), .Z(n8624) );
  AND U17249 ( .A(n8625), .B(p_input[2238]), .Z(o[2238]) );
  AND U17250 ( .A(p_input[22238]), .B(p_input[12238]), .Z(n8625) );
  AND U17251 ( .A(n8626), .B(p_input[2237]), .Z(o[2237]) );
  AND U17252 ( .A(p_input[22237]), .B(p_input[12237]), .Z(n8626) );
  AND U17253 ( .A(n8627), .B(p_input[2236]), .Z(o[2236]) );
  AND U17254 ( .A(p_input[22236]), .B(p_input[12236]), .Z(n8627) );
  AND U17255 ( .A(n8628), .B(p_input[2235]), .Z(o[2235]) );
  AND U17256 ( .A(p_input[22235]), .B(p_input[12235]), .Z(n8628) );
  AND U17257 ( .A(n8629), .B(p_input[2234]), .Z(o[2234]) );
  AND U17258 ( .A(p_input[22234]), .B(p_input[12234]), .Z(n8629) );
  AND U17259 ( .A(n8630), .B(p_input[2233]), .Z(o[2233]) );
  AND U17260 ( .A(p_input[22233]), .B(p_input[12233]), .Z(n8630) );
  AND U17261 ( .A(n8631), .B(p_input[2232]), .Z(o[2232]) );
  AND U17262 ( .A(p_input[22232]), .B(p_input[12232]), .Z(n8631) );
  AND U17263 ( .A(n8632), .B(p_input[2231]), .Z(o[2231]) );
  AND U17264 ( .A(p_input[22231]), .B(p_input[12231]), .Z(n8632) );
  AND U17265 ( .A(n8633), .B(p_input[2230]), .Z(o[2230]) );
  AND U17266 ( .A(p_input[22230]), .B(p_input[12230]), .Z(n8633) );
  AND U17267 ( .A(n8634), .B(p_input[222]), .Z(o[222]) );
  AND U17268 ( .A(p_input[20222]), .B(p_input[10222]), .Z(n8634) );
  AND U17269 ( .A(n8635), .B(p_input[2229]), .Z(o[2229]) );
  AND U17270 ( .A(p_input[22229]), .B(p_input[12229]), .Z(n8635) );
  AND U17271 ( .A(n8636), .B(p_input[2228]), .Z(o[2228]) );
  AND U17272 ( .A(p_input[22228]), .B(p_input[12228]), .Z(n8636) );
  AND U17273 ( .A(n8637), .B(p_input[2227]), .Z(o[2227]) );
  AND U17274 ( .A(p_input[22227]), .B(p_input[12227]), .Z(n8637) );
  AND U17275 ( .A(n8638), .B(p_input[2226]), .Z(o[2226]) );
  AND U17276 ( .A(p_input[22226]), .B(p_input[12226]), .Z(n8638) );
  AND U17277 ( .A(n8639), .B(p_input[2225]), .Z(o[2225]) );
  AND U17278 ( .A(p_input[22225]), .B(p_input[12225]), .Z(n8639) );
  AND U17279 ( .A(n8640), .B(p_input[2224]), .Z(o[2224]) );
  AND U17280 ( .A(p_input[22224]), .B(p_input[12224]), .Z(n8640) );
  AND U17281 ( .A(n8641), .B(p_input[2223]), .Z(o[2223]) );
  AND U17282 ( .A(p_input[22223]), .B(p_input[12223]), .Z(n8641) );
  AND U17283 ( .A(n8642), .B(p_input[2222]), .Z(o[2222]) );
  AND U17284 ( .A(p_input[22222]), .B(p_input[12222]), .Z(n8642) );
  AND U17285 ( .A(n8643), .B(p_input[22221]), .Z(o[2221]) );
  AND U17286 ( .A(p_input[2221]), .B(p_input[12221]), .Z(n8643) );
  AND U17287 ( .A(n8644), .B(p_input[22220]), .Z(o[2220]) );
  AND U17288 ( .A(p_input[2220]), .B(p_input[12220]), .Z(n8644) );
  AND U17289 ( .A(n8645), .B(p_input[221]), .Z(o[221]) );
  AND U17290 ( .A(p_input[20221]), .B(p_input[10221]), .Z(n8645) );
  AND U17291 ( .A(n8646), .B(p_input[22219]), .Z(o[2219]) );
  AND U17292 ( .A(p_input[2219]), .B(p_input[12219]), .Z(n8646) );
  AND U17293 ( .A(n8647), .B(p_input[22218]), .Z(o[2218]) );
  AND U17294 ( .A(p_input[2218]), .B(p_input[12218]), .Z(n8647) );
  AND U17295 ( .A(n8648), .B(p_input[22217]), .Z(o[2217]) );
  AND U17296 ( .A(p_input[2217]), .B(p_input[12217]), .Z(n8648) );
  AND U17297 ( .A(n8649), .B(p_input[22216]), .Z(o[2216]) );
  AND U17298 ( .A(p_input[2216]), .B(p_input[12216]), .Z(n8649) );
  AND U17299 ( .A(n8650), .B(p_input[22215]), .Z(o[2215]) );
  AND U17300 ( .A(p_input[2215]), .B(p_input[12215]), .Z(n8650) );
  AND U17301 ( .A(n8651), .B(p_input[22214]), .Z(o[2214]) );
  AND U17302 ( .A(p_input[2214]), .B(p_input[12214]), .Z(n8651) );
  AND U17303 ( .A(n8652), .B(p_input[22213]), .Z(o[2213]) );
  AND U17304 ( .A(p_input[2213]), .B(p_input[12213]), .Z(n8652) );
  AND U17305 ( .A(n8653), .B(p_input[22212]), .Z(o[2212]) );
  AND U17306 ( .A(p_input[2212]), .B(p_input[12212]), .Z(n8653) );
  AND U17307 ( .A(n8654), .B(p_input[22211]), .Z(o[2211]) );
  AND U17308 ( .A(p_input[2211]), .B(p_input[12211]), .Z(n8654) );
  AND U17309 ( .A(n8655), .B(p_input[22210]), .Z(o[2210]) );
  AND U17310 ( .A(p_input[2210]), .B(p_input[12210]), .Z(n8655) );
  AND U17311 ( .A(n8656), .B(p_input[220]), .Z(o[220]) );
  AND U17312 ( .A(p_input[20220]), .B(p_input[10220]), .Z(n8656) );
  AND U17313 ( .A(n8657), .B(p_input[22209]), .Z(o[2209]) );
  AND U17314 ( .A(p_input[2209]), .B(p_input[12209]), .Z(n8657) );
  AND U17315 ( .A(n8658), .B(p_input[22208]), .Z(o[2208]) );
  AND U17316 ( .A(p_input[2208]), .B(p_input[12208]), .Z(n8658) );
  AND U17317 ( .A(n8659), .B(p_input[22207]), .Z(o[2207]) );
  AND U17318 ( .A(p_input[2207]), .B(p_input[12207]), .Z(n8659) );
  AND U17319 ( .A(n8660), .B(p_input[22206]), .Z(o[2206]) );
  AND U17320 ( .A(p_input[2206]), .B(p_input[12206]), .Z(n8660) );
  AND U17321 ( .A(n8661), .B(p_input[22205]), .Z(o[2205]) );
  AND U17322 ( .A(p_input[2205]), .B(p_input[12205]), .Z(n8661) );
  AND U17323 ( .A(n8662), .B(p_input[22204]), .Z(o[2204]) );
  AND U17324 ( .A(p_input[2204]), .B(p_input[12204]), .Z(n8662) );
  AND U17325 ( .A(n8663), .B(p_input[22203]), .Z(o[2203]) );
  AND U17326 ( .A(p_input[2203]), .B(p_input[12203]), .Z(n8663) );
  AND U17327 ( .A(n8664), .B(p_input[22202]), .Z(o[2202]) );
  AND U17328 ( .A(p_input[2202]), .B(p_input[12202]), .Z(n8664) );
  AND U17329 ( .A(n8665), .B(p_input[22201]), .Z(o[2201]) );
  AND U17330 ( .A(p_input[2201]), .B(p_input[12201]), .Z(n8665) );
  AND U17331 ( .A(n8666), .B(p_input[22200]), .Z(o[2200]) );
  AND U17332 ( .A(p_input[2200]), .B(p_input[12200]), .Z(n8666) );
  AND U17333 ( .A(n8667), .B(p_input[21]), .Z(o[21]) );
  AND U17334 ( .A(p_input[20021]), .B(p_input[10021]), .Z(n8667) );
  AND U17335 ( .A(n8668), .B(p_input[219]), .Z(o[219]) );
  AND U17336 ( .A(p_input[20219]), .B(p_input[10219]), .Z(n8668) );
  AND U17337 ( .A(n8669), .B(p_input[22199]), .Z(o[2199]) );
  AND U17338 ( .A(p_input[2199]), .B(p_input[12199]), .Z(n8669) );
  AND U17339 ( .A(n8670), .B(p_input[22198]), .Z(o[2198]) );
  AND U17340 ( .A(p_input[2198]), .B(p_input[12198]), .Z(n8670) );
  AND U17341 ( .A(n8671), .B(p_input[22197]), .Z(o[2197]) );
  AND U17342 ( .A(p_input[2197]), .B(p_input[12197]), .Z(n8671) );
  AND U17343 ( .A(n8672), .B(p_input[22196]), .Z(o[2196]) );
  AND U17344 ( .A(p_input[2196]), .B(p_input[12196]), .Z(n8672) );
  AND U17345 ( .A(n8673), .B(p_input[22195]), .Z(o[2195]) );
  AND U17346 ( .A(p_input[2195]), .B(p_input[12195]), .Z(n8673) );
  AND U17347 ( .A(n8674), .B(p_input[22194]), .Z(o[2194]) );
  AND U17348 ( .A(p_input[2194]), .B(p_input[12194]), .Z(n8674) );
  AND U17349 ( .A(n8675), .B(p_input[22193]), .Z(o[2193]) );
  AND U17350 ( .A(p_input[2193]), .B(p_input[12193]), .Z(n8675) );
  AND U17351 ( .A(n8676), .B(p_input[22192]), .Z(o[2192]) );
  AND U17352 ( .A(p_input[2192]), .B(p_input[12192]), .Z(n8676) );
  AND U17353 ( .A(n8677), .B(p_input[22191]), .Z(o[2191]) );
  AND U17354 ( .A(p_input[2191]), .B(p_input[12191]), .Z(n8677) );
  AND U17355 ( .A(n8678), .B(p_input[22190]), .Z(o[2190]) );
  AND U17356 ( .A(p_input[2190]), .B(p_input[12190]), .Z(n8678) );
  AND U17357 ( .A(n8679), .B(p_input[218]), .Z(o[218]) );
  AND U17358 ( .A(p_input[20218]), .B(p_input[10218]), .Z(n8679) );
  AND U17359 ( .A(n8680), .B(p_input[22189]), .Z(o[2189]) );
  AND U17360 ( .A(p_input[2189]), .B(p_input[12189]), .Z(n8680) );
  AND U17361 ( .A(n8681), .B(p_input[22188]), .Z(o[2188]) );
  AND U17362 ( .A(p_input[2188]), .B(p_input[12188]), .Z(n8681) );
  AND U17363 ( .A(n8682), .B(p_input[22187]), .Z(o[2187]) );
  AND U17364 ( .A(p_input[2187]), .B(p_input[12187]), .Z(n8682) );
  AND U17365 ( .A(n8683), .B(p_input[22186]), .Z(o[2186]) );
  AND U17366 ( .A(p_input[2186]), .B(p_input[12186]), .Z(n8683) );
  AND U17367 ( .A(n8684), .B(p_input[22185]), .Z(o[2185]) );
  AND U17368 ( .A(p_input[2185]), .B(p_input[12185]), .Z(n8684) );
  AND U17369 ( .A(n8685), .B(p_input[22184]), .Z(o[2184]) );
  AND U17370 ( .A(p_input[2184]), .B(p_input[12184]), .Z(n8685) );
  AND U17371 ( .A(n8686), .B(p_input[22183]), .Z(o[2183]) );
  AND U17372 ( .A(p_input[2183]), .B(p_input[12183]), .Z(n8686) );
  AND U17373 ( .A(n8687), .B(p_input[22182]), .Z(o[2182]) );
  AND U17374 ( .A(p_input[2182]), .B(p_input[12182]), .Z(n8687) );
  AND U17375 ( .A(n8688), .B(p_input[22181]), .Z(o[2181]) );
  AND U17376 ( .A(p_input[2181]), .B(p_input[12181]), .Z(n8688) );
  AND U17377 ( .A(n8689), .B(p_input[22180]), .Z(o[2180]) );
  AND U17378 ( .A(p_input[2180]), .B(p_input[12180]), .Z(n8689) );
  AND U17379 ( .A(n8690), .B(p_input[217]), .Z(o[217]) );
  AND U17380 ( .A(p_input[20217]), .B(p_input[10217]), .Z(n8690) );
  AND U17381 ( .A(n8691), .B(p_input[22179]), .Z(o[2179]) );
  AND U17382 ( .A(p_input[2179]), .B(p_input[12179]), .Z(n8691) );
  AND U17383 ( .A(n8692), .B(p_input[22178]), .Z(o[2178]) );
  AND U17384 ( .A(p_input[2178]), .B(p_input[12178]), .Z(n8692) );
  AND U17385 ( .A(n8693), .B(p_input[22177]), .Z(o[2177]) );
  AND U17386 ( .A(p_input[2177]), .B(p_input[12177]), .Z(n8693) );
  AND U17387 ( .A(n8694), .B(p_input[22176]), .Z(o[2176]) );
  AND U17388 ( .A(p_input[2176]), .B(p_input[12176]), .Z(n8694) );
  AND U17389 ( .A(n8695), .B(p_input[22175]), .Z(o[2175]) );
  AND U17390 ( .A(p_input[2175]), .B(p_input[12175]), .Z(n8695) );
  AND U17391 ( .A(n8696), .B(p_input[22174]), .Z(o[2174]) );
  AND U17392 ( .A(p_input[2174]), .B(p_input[12174]), .Z(n8696) );
  AND U17393 ( .A(n8697), .B(p_input[22173]), .Z(o[2173]) );
  AND U17394 ( .A(p_input[2173]), .B(p_input[12173]), .Z(n8697) );
  AND U17395 ( .A(n8698), .B(p_input[22172]), .Z(o[2172]) );
  AND U17396 ( .A(p_input[2172]), .B(p_input[12172]), .Z(n8698) );
  AND U17397 ( .A(n8699), .B(p_input[22171]), .Z(o[2171]) );
  AND U17398 ( .A(p_input[2171]), .B(p_input[12171]), .Z(n8699) );
  AND U17399 ( .A(n8700), .B(p_input[22170]), .Z(o[2170]) );
  AND U17400 ( .A(p_input[2170]), .B(p_input[12170]), .Z(n8700) );
  AND U17401 ( .A(n8701), .B(p_input[216]), .Z(o[216]) );
  AND U17402 ( .A(p_input[20216]), .B(p_input[10216]), .Z(n8701) );
  AND U17403 ( .A(n8702), .B(p_input[22169]), .Z(o[2169]) );
  AND U17404 ( .A(p_input[2169]), .B(p_input[12169]), .Z(n8702) );
  AND U17405 ( .A(n8703), .B(p_input[22168]), .Z(o[2168]) );
  AND U17406 ( .A(p_input[2168]), .B(p_input[12168]), .Z(n8703) );
  AND U17407 ( .A(n8704), .B(p_input[22167]), .Z(o[2167]) );
  AND U17408 ( .A(p_input[2167]), .B(p_input[12167]), .Z(n8704) );
  AND U17409 ( .A(n8705), .B(p_input[22166]), .Z(o[2166]) );
  AND U17410 ( .A(p_input[2166]), .B(p_input[12166]), .Z(n8705) );
  AND U17411 ( .A(n8706), .B(p_input[22165]), .Z(o[2165]) );
  AND U17412 ( .A(p_input[2165]), .B(p_input[12165]), .Z(n8706) );
  AND U17413 ( .A(n8707), .B(p_input[22164]), .Z(o[2164]) );
  AND U17414 ( .A(p_input[2164]), .B(p_input[12164]), .Z(n8707) );
  AND U17415 ( .A(n8708), .B(p_input[22163]), .Z(o[2163]) );
  AND U17416 ( .A(p_input[2163]), .B(p_input[12163]), .Z(n8708) );
  AND U17417 ( .A(n8709), .B(p_input[22162]), .Z(o[2162]) );
  AND U17418 ( .A(p_input[2162]), .B(p_input[12162]), .Z(n8709) );
  AND U17419 ( .A(n8710), .B(p_input[22161]), .Z(o[2161]) );
  AND U17420 ( .A(p_input[2161]), .B(p_input[12161]), .Z(n8710) );
  AND U17421 ( .A(n8711), .B(p_input[22160]), .Z(o[2160]) );
  AND U17422 ( .A(p_input[2160]), .B(p_input[12160]), .Z(n8711) );
  AND U17423 ( .A(n8712), .B(p_input[215]), .Z(o[215]) );
  AND U17424 ( .A(p_input[20215]), .B(p_input[10215]), .Z(n8712) );
  AND U17425 ( .A(n8713), .B(p_input[22159]), .Z(o[2159]) );
  AND U17426 ( .A(p_input[2159]), .B(p_input[12159]), .Z(n8713) );
  AND U17427 ( .A(n8714), .B(p_input[22158]), .Z(o[2158]) );
  AND U17428 ( .A(p_input[2158]), .B(p_input[12158]), .Z(n8714) );
  AND U17429 ( .A(n8715), .B(p_input[22157]), .Z(o[2157]) );
  AND U17430 ( .A(p_input[2157]), .B(p_input[12157]), .Z(n8715) );
  AND U17431 ( .A(n8716), .B(p_input[22156]), .Z(o[2156]) );
  AND U17432 ( .A(p_input[2156]), .B(p_input[12156]), .Z(n8716) );
  AND U17433 ( .A(n8717), .B(p_input[22155]), .Z(o[2155]) );
  AND U17434 ( .A(p_input[2155]), .B(p_input[12155]), .Z(n8717) );
  AND U17435 ( .A(n8718), .B(p_input[22154]), .Z(o[2154]) );
  AND U17436 ( .A(p_input[2154]), .B(p_input[12154]), .Z(n8718) );
  AND U17437 ( .A(n8719), .B(p_input[22153]), .Z(o[2153]) );
  AND U17438 ( .A(p_input[2153]), .B(p_input[12153]), .Z(n8719) );
  AND U17439 ( .A(n8720), .B(p_input[22152]), .Z(o[2152]) );
  AND U17440 ( .A(p_input[2152]), .B(p_input[12152]), .Z(n8720) );
  AND U17441 ( .A(n8721), .B(p_input[22151]), .Z(o[2151]) );
  AND U17442 ( .A(p_input[2151]), .B(p_input[12151]), .Z(n8721) );
  AND U17443 ( .A(n8722), .B(p_input[22150]), .Z(o[2150]) );
  AND U17444 ( .A(p_input[2150]), .B(p_input[12150]), .Z(n8722) );
  AND U17445 ( .A(n8723), .B(p_input[214]), .Z(o[214]) );
  AND U17446 ( .A(p_input[20214]), .B(p_input[10214]), .Z(n8723) );
  AND U17447 ( .A(n8724), .B(p_input[22149]), .Z(o[2149]) );
  AND U17448 ( .A(p_input[2149]), .B(p_input[12149]), .Z(n8724) );
  AND U17449 ( .A(n8725), .B(p_input[22148]), .Z(o[2148]) );
  AND U17450 ( .A(p_input[2148]), .B(p_input[12148]), .Z(n8725) );
  AND U17451 ( .A(n8726), .B(p_input[22147]), .Z(o[2147]) );
  AND U17452 ( .A(p_input[2147]), .B(p_input[12147]), .Z(n8726) );
  AND U17453 ( .A(n8727), .B(p_input[22146]), .Z(o[2146]) );
  AND U17454 ( .A(p_input[2146]), .B(p_input[12146]), .Z(n8727) );
  AND U17455 ( .A(n8728), .B(p_input[22145]), .Z(o[2145]) );
  AND U17456 ( .A(p_input[2145]), .B(p_input[12145]), .Z(n8728) );
  AND U17457 ( .A(n8729), .B(p_input[22144]), .Z(o[2144]) );
  AND U17458 ( .A(p_input[2144]), .B(p_input[12144]), .Z(n8729) );
  AND U17459 ( .A(n8730), .B(p_input[22143]), .Z(o[2143]) );
  AND U17460 ( .A(p_input[2143]), .B(p_input[12143]), .Z(n8730) );
  AND U17461 ( .A(n8731), .B(p_input[22142]), .Z(o[2142]) );
  AND U17462 ( .A(p_input[2142]), .B(p_input[12142]), .Z(n8731) );
  AND U17463 ( .A(n8732), .B(p_input[22141]), .Z(o[2141]) );
  AND U17464 ( .A(p_input[2141]), .B(p_input[12141]), .Z(n8732) );
  AND U17465 ( .A(n8733), .B(p_input[22140]), .Z(o[2140]) );
  AND U17466 ( .A(p_input[2140]), .B(p_input[12140]), .Z(n8733) );
  AND U17467 ( .A(n8734), .B(p_input[213]), .Z(o[213]) );
  AND U17468 ( .A(p_input[20213]), .B(p_input[10213]), .Z(n8734) );
  AND U17469 ( .A(n8735), .B(p_input[22139]), .Z(o[2139]) );
  AND U17470 ( .A(p_input[2139]), .B(p_input[12139]), .Z(n8735) );
  AND U17471 ( .A(n8736), .B(p_input[22138]), .Z(o[2138]) );
  AND U17472 ( .A(p_input[2138]), .B(p_input[12138]), .Z(n8736) );
  AND U17473 ( .A(n8737), .B(p_input[22137]), .Z(o[2137]) );
  AND U17474 ( .A(p_input[2137]), .B(p_input[12137]), .Z(n8737) );
  AND U17475 ( .A(n8738), .B(p_input[22136]), .Z(o[2136]) );
  AND U17476 ( .A(p_input[2136]), .B(p_input[12136]), .Z(n8738) );
  AND U17477 ( .A(n8739), .B(p_input[22135]), .Z(o[2135]) );
  AND U17478 ( .A(p_input[2135]), .B(p_input[12135]), .Z(n8739) );
  AND U17479 ( .A(n8740), .B(p_input[22134]), .Z(o[2134]) );
  AND U17480 ( .A(p_input[2134]), .B(p_input[12134]), .Z(n8740) );
  AND U17481 ( .A(n8741), .B(p_input[22133]), .Z(o[2133]) );
  AND U17482 ( .A(p_input[2133]), .B(p_input[12133]), .Z(n8741) );
  AND U17483 ( .A(n8742), .B(p_input[22132]), .Z(o[2132]) );
  AND U17484 ( .A(p_input[2132]), .B(p_input[12132]), .Z(n8742) );
  AND U17485 ( .A(n8743), .B(p_input[22131]), .Z(o[2131]) );
  AND U17486 ( .A(p_input[2131]), .B(p_input[12131]), .Z(n8743) );
  AND U17487 ( .A(n8744), .B(p_input[22130]), .Z(o[2130]) );
  AND U17488 ( .A(p_input[2130]), .B(p_input[12130]), .Z(n8744) );
  AND U17489 ( .A(n8745), .B(p_input[212]), .Z(o[212]) );
  AND U17490 ( .A(p_input[20212]), .B(p_input[10212]), .Z(n8745) );
  AND U17491 ( .A(n8746), .B(p_input[22129]), .Z(o[2129]) );
  AND U17492 ( .A(p_input[2129]), .B(p_input[12129]), .Z(n8746) );
  AND U17493 ( .A(n8747), .B(p_input[22128]), .Z(o[2128]) );
  AND U17494 ( .A(p_input[2128]), .B(p_input[12128]), .Z(n8747) );
  AND U17495 ( .A(n8748), .B(p_input[22127]), .Z(o[2127]) );
  AND U17496 ( .A(p_input[2127]), .B(p_input[12127]), .Z(n8748) );
  AND U17497 ( .A(n8749), .B(p_input[22126]), .Z(o[2126]) );
  AND U17498 ( .A(p_input[2126]), .B(p_input[12126]), .Z(n8749) );
  AND U17499 ( .A(n8750), .B(p_input[22125]), .Z(o[2125]) );
  AND U17500 ( .A(p_input[2125]), .B(p_input[12125]), .Z(n8750) );
  AND U17501 ( .A(n8751), .B(p_input[22124]), .Z(o[2124]) );
  AND U17502 ( .A(p_input[2124]), .B(p_input[12124]), .Z(n8751) );
  AND U17503 ( .A(n8752), .B(p_input[22123]), .Z(o[2123]) );
  AND U17504 ( .A(p_input[2123]), .B(p_input[12123]), .Z(n8752) );
  AND U17505 ( .A(n8753), .B(p_input[22122]), .Z(o[2122]) );
  AND U17506 ( .A(p_input[2122]), .B(p_input[12122]), .Z(n8753) );
  AND U17507 ( .A(n8754), .B(p_input[22121]), .Z(o[2121]) );
  AND U17508 ( .A(p_input[2121]), .B(p_input[12121]), .Z(n8754) );
  AND U17509 ( .A(n8755), .B(p_input[22120]), .Z(o[2120]) );
  AND U17510 ( .A(p_input[2120]), .B(p_input[12120]), .Z(n8755) );
  AND U17511 ( .A(n8756), .B(p_input[211]), .Z(o[211]) );
  AND U17512 ( .A(p_input[20211]), .B(p_input[10211]), .Z(n8756) );
  AND U17513 ( .A(n8757), .B(p_input[22119]), .Z(o[2119]) );
  AND U17514 ( .A(p_input[2119]), .B(p_input[12119]), .Z(n8757) );
  AND U17515 ( .A(n8758), .B(p_input[22118]), .Z(o[2118]) );
  AND U17516 ( .A(p_input[2118]), .B(p_input[12118]), .Z(n8758) );
  AND U17517 ( .A(n8759), .B(p_input[22117]), .Z(o[2117]) );
  AND U17518 ( .A(p_input[2117]), .B(p_input[12117]), .Z(n8759) );
  AND U17519 ( .A(n8760), .B(p_input[22116]), .Z(o[2116]) );
  AND U17520 ( .A(p_input[2116]), .B(p_input[12116]), .Z(n8760) );
  AND U17521 ( .A(n8761), .B(p_input[22115]), .Z(o[2115]) );
  AND U17522 ( .A(p_input[2115]), .B(p_input[12115]), .Z(n8761) );
  AND U17523 ( .A(n8762), .B(p_input[22114]), .Z(o[2114]) );
  AND U17524 ( .A(p_input[2114]), .B(p_input[12114]), .Z(n8762) );
  AND U17525 ( .A(n8763), .B(p_input[22113]), .Z(o[2113]) );
  AND U17526 ( .A(p_input[2113]), .B(p_input[12113]), .Z(n8763) );
  AND U17527 ( .A(n8764), .B(p_input[22112]), .Z(o[2112]) );
  AND U17528 ( .A(p_input[2112]), .B(p_input[12112]), .Z(n8764) );
  AND U17529 ( .A(n8765), .B(p_input[22111]), .Z(o[2111]) );
  AND U17530 ( .A(p_input[2111]), .B(p_input[12111]), .Z(n8765) );
  AND U17531 ( .A(n8766), .B(p_input[22110]), .Z(o[2110]) );
  AND U17532 ( .A(p_input[2110]), .B(p_input[12110]), .Z(n8766) );
  AND U17533 ( .A(n8767), .B(p_input[210]), .Z(o[210]) );
  AND U17534 ( .A(p_input[20210]), .B(p_input[10210]), .Z(n8767) );
  AND U17535 ( .A(n8768), .B(p_input[22109]), .Z(o[2109]) );
  AND U17536 ( .A(p_input[2109]), .B(p_input[12109]), .Z(n8768) );
  AND U17537 ( .A(n8769), .B(p_input[22108]), .Z(o[2108]) );
  AND U17538 ( .A(p_input[2108]), .B(p_input[12108]), .Z(n8769) );
  AND U17539 ( .A(n8770), .B(p_input[22107]), .Z(o[2107]) );
  AND U17540 ( .A(p_input[2107]), .B(p_input[12107]), .Z(n8770) );
  AND U17541 ( .A(n8771), .B(p_input[22106]), .Z(o[2106]) );
  AND U17542 ( .A(p_input[2106]), .B(p_input[12106]), .Z(n8771) );
  AND U17543 ( .A(n8772), .B(p_input[22105]), .Z(o[2105]) );
  AND U17544 ( .A(p_input[2105]), .B(p_input[12105]), .Z(n8772) );
  AND U17545 ( .A(n8773), .B(p_input[22104]), .Z(o[2104]) );
  AND U17546 ( .A(p_input[2104]), .B(p_input[12104]), .Z(n8773) );
  AND U17547 ( .A(n8774), .B(p_input[22103]), .Z(o[2103]) );
  AND U17548 ( .A(p_input[2103]), .B(p_input[12103]), .Z(n8774) );
  AND U17549 ( .A(n8775), .B(p_input[22102]), .Z(o[2102]) );
  AND U17550 ( .A(p_input[2102]), .B(p_input[12102]), .Z(n8775) );
  AND U17551 ( .A(n8776), .B(p_input[22101]), .Z(o[2101]) );
  AND U17552 ( .A(p_input[2101]), .B(p_input[12101]), .Z(n8776) );
  AND U17553 ( .A(n8777), .B(p_input[22100]), .Z(o[2100]) );
  AND U17554 ( .A(p_input[2100]), .B(p_input[12100]), .Z(n8777) );
  AND U17555 ( .A(n8778), .B(p_input[20]), .Z(o[20]) );
  AND U17556 ( .A(p_input[20020]), .B(p_input[10020]), .Z(n8778) );
  AND U17557 ( .A(n8779), .B(p_input[209]), .Z(o[209]) );
  AND U17558 ( .A(p_input[20209]), .B(p_input[10209]), .Z(n8779) );
  AND U17559 ( .A(n8780), .B(p_input[22099]), .Z(o[2099]) );
  AND U17560 ( .A(p_input[2099]), .B(p_input[12099]), .Z(n8780) );
  AND U17561 ( .A(n8781), .B(p_input[22098]), .Z(o[2098]) );
  AND U17562 ( .A(p_input[2098]), .B(p_input[12098]), .Z(n8781) );
  AND U17563 ( .A(n8782), .B(p_input[22097]), .Z(o[2097]) );
  AND U17564 ( .A(p_input[2097]), .B(p_input[12097]), .Z(n8782) );
  AND U17565 ( .A(n8783), .B(p_input[22096]), .Z(o[2096]) );
  AND U17566 ( .A(p_input[2096]), .B(p_input[12096]), .Z(n8783) );
  AND U17567 ( .A(n8784), .B(p_input[22095]), .Z(o[2095]) );
  AND U17568 ( .A(p_input[2095]), .B(p_input[12095]), .Z(n8784) );
  AND U17569 ( .A(n8785), .B(p_input[22094]), .Z(o[2094]) );
  AND U17570 ( .A(p_input[2094]), .B(p_input[12094]), .Z(n8785) );
  AND U17571 ( .A(n8786), .B(p_input[22093]), .Z(o[2093]) );
  AND U17572 ( .A(p_input[2093]), .B(p_input[12093]), .Z(n8786) );
  AND U17573 ( .A(n8787), .B(p_input[22092]), .Z(o[2092]) );
  AND U17574 ( .A(p_input[2092]), .B(p_input[12092]), .Z(n8787) );
  AND U17575 ( .A(n8788), .B(p_input[22091]), .Z(o[2091]) );
  AND U17576 ( .A(p_input[2091]), .B(p_input[12091]), .Z(n8788) );
  AND U17577 ( .A(n8789), .B(p_input[22090]), .Z(o[2090]) );
  AND U17578 ( .A(p_input[2090]), .B(p_input[12090]), .Z(n8789) );
  AND U17579 ( .A(n8790), .B(p_input[208]), .Z(o[208]) );
  AND U17580 ( .A(p_input[20208]), .B(p_input[10208]), .Z(n8790) );
  AND U17581 ( .A(n8791), .B(p_input[22089]), .Z(o[2089]) );
  AND U17582 ( .A(p_input[2089]), .B(p_input[12089]), .Z(n8791) );
  AND U17583 ( .A(n8792), .B(p_input[22088]), .Z(o[2088]) );
  AND U17584 ( .A(p_input[2088]), .B(p_input[12088]), .Z(n8792) );
  AND U17585 ( .A(n8793), .B(p_input[22087]), .Z(o[2087]) );
  AND U17586 ( .A(p_input[2087]), .B(p_input[12087]), .Z(n8793) );
  AND U17587 ( .A(n8794), .B(p_input[22086]), .Z(o[2086]) );
  AND U17588 ( .A(p_input[2086]), .B(p_input[12086]), .Z(n8794) );
  AND U17589 ( .A(n8795), .B(p_input[22085]), .Z(o[2085]) );
  AND U17590 ( .A(p_input[2085]), .B(p_input[12085]), .Z(n8795) );
  AND U17591 ( .A(n8796), .B(p_input[22084]), .Z(o[2084]) );
  AND U17592 ( .A(p_input[2084]), .B(p_input[12084]), .Z(n8796) );
  AND U17593 ( .A(n8797), .B(p_input[22083]), .Z(o[2083]) );
  AND U17594 ( .A(p_input[2083]), .B(p_input[12083]), .Z(n8797) );
  AND U17595 ( .A(n8798), .B(p_input[22082]), .Z(o[2082]) );
  AND U17596 ( .A(p_input[2082]), .B(p_input[12082]), .Z(n8798) );
  AND U17597 ( .A(n8799), .B(p_input[22081]), .Z(o[2081]) );
  AND U17598 ( .A(p_input[2081]), .B(p_input[12081]), .Z(n8799) );
  AND U17599 ( .A(n8800), .B(p_input[22080]), .Z(o[2080]) );
  AND U17600 ( .A(p_input[2080]), .B(p_input[12080]), .Z(n8800) );
  AND U17601 ( .A(n8801), .B(p_input[207]), .Z(o[207]) );
  AND U17602 ( .A(p_input[20207]), .B(p_input[10207]), .Z(n8801) );
  AND U17603 ( .A(n8802), .B(p_input[22079]), .Z(o[2079]) );
  AND U17604 ( .A(p_input[2079]), .B(p_input[12079]), .Z(n8802) );
  AND U17605 ( .A(n8803), .B(p_input[22078]), .Z(o[2078]) );
  AND U17606 ( .A(p_input[2078]), .B(p_input[12078]), .Z(n8803) );
  AND U17607 ( .A(n8804), .B(p_input[22077]), .Z(o[2077]) );
  AND U17608 ( .A(p_input[2077]), .B(p_input[12077]), .Z(n8804) );
  AND U17609 ( .A(n8805), .B(p_input[22076]), .Z(o[2076]) );
  AND U17610 ( .A(p_input[2076]), .B(p_input[12076]), .Z(n8805) );
  AND U17611 ( .A(n8806), .B(p_input[22075]), .Z(o[2075]) );
  AND U17612 ( .A(p_input[2075]), .B(p_input[12075]), .Z(n8806) );
  AND U17613 ( .A(n8807), .B(p_input[22074]), .Z(o[2074]) );
  AND U17614 ( .A(p_input[2074]), .B(p_input[12074]), .Z(n8807) );
  AND U17615 ( .A(n8808), .B(p_input[22073]), .Z(o[2073]) );
  AND U17616 ( .A(p_input[2073]), .B(p_input[12073]), .Z(n8808) );
  AND U17617 ( .A(n8809), .B(p_input[22072]), .Z(o[2072]) );
  AND U17618 ( .A(p_input[2072]), .B(p_input[12072]), .Z(n8809) );
  AND U17619 ( .A(n8810), .B(p_input[22071]), .Z(o[2071]) );
  AND U17620 ( .A(p_input[2071]), .B(p_input[12071]), .Z(n8810) );
  AND U17621 ( .A(n8811), .B(p_input[22070]), .Z(o[2070]) );
  AND U17622 ( .A(p_input[2070]), .B(p_input[12070]), .Z(n8811) );
  AND U17623 ( .A(n8812), .B(p_input[206]), .Z(o[206]) );
  AND U17624 ( .A(p_input[20206]), .B(p_input[10206]), .Z(n8812) );
  AND U17625 ( .A(n8813), .B(p_input[22069]), .Z(o[2069]) );
  AND U17626 ( .A(p_input[2069]), .B(p_input[12069]), .Z(n8813) );
  AND U17627 ( .A(n8814), .B(p_input[22068]), .Z(o[2068]) );
  AND U17628 ( .A(p_input[2068]), .B(p_input[12068]), .Z(n8814) );
  AND U17629 ( .A(n8815), .B(p_input[22067]), .Z(o[2067]) );
  AND U17630 ( .A(p_input[2067]), .B(p_input[12067]), .Z(n8815) );
  AND U17631 ( .A(n8816), .B(p_input[22066]), .Z(o[2066]) );
  AND U17632 ( .A(p_input[2066]), .B(p_input[12066]), .Z(n8816) );
  AND U17633 ( .A(n8817), .B(p_input[22065]), .Z(o[2065]) );
  AND U17634 ( .A(p_input[2065]), .B(p_input[12065]), .Z(n8817) );
  AND U17635 ( .A(n8818), .B(p_input[22064]), .Z(o[2064]) );
  AND U17636 ( .A(p_input[2064]), .B(p_input[12064]), .Z(n8818) );
  AND U17637 ( .A(n8819), .B(p_input[22063]), .Z(o[2063]) );
  AND U17638 ( .A(p_input[2063]), .B(p_input[12063]), .Z(n8819) );
  AND U17639 ( .A(n8820), .B(p_input[22062]), .Z(o[2062]) );
  AND U17640 ( .A(p_input[2062]), .B(p_input[12062]), .Z(n8820) );
  AND U17641 ( .A(n8821), .B(p_input[22061]), .Z(o[2061]) );
  AND U17642 ( .A(p_input[2061]), .B(p_input[12061]), .Z(n8821) );
  AND U17643 ( .A(n8822), .B(p_input[22060]), .Z(o[2060]) );
  AND U17644 ( .A(p_input[2060]), .B(p_input[12060]), .Z(n8822) );
  AND U17645 ( .A(n8823), .B(p_input[205]), .Z(o[205]) );
  AND U17646 ( .A(p_input[20205]), .B(p_input[10205]), .Z(n8823) );
  AND U17647 ( .A(n8824), .B(p_input[22059]), .Z(o[2059]) );
  AND U17648 ( .A(p_input[2059]), .B(p_input[12059]), .Z(n8824) );
  AND U17649 ( .A(n8825), .B(p_input[22058]), .Z(o[2058]) );
  AND U17650 ( .A(p_input[2058]), .B(p_input[12058]), .Z(n8825) );
  AND U17651 ( .A(n8826), .B(p_input[22057]), .Z(o[2057]) );
  AND U17652 ( .A(p_input[2057]), .B(p_input[12057]), .Z(n8826) );
  AND U17653 ( .A(n8827), .B(p_input[22056]), .Z(o[2056]) );
  AND U17654 ( .A(p_input[2056]), .B(p_input[12056]), .Z(n8827) );
  AND U17655 ( .A(n8828), .B(p_input[22055]), .Z(o[2055]) );
  AND U17656 ( .A(p_input[2055]), .B(p_input[12055]), .Z(n8828) );
  AND U17657 ( .A(n8829), .B(p_input[22054]), .Z(o[2054]) );
  AND U17658 ( .A(p_input[2054]), .B(p_input[12054]), .Z(n8829) );
  AND U17659 ( .A(n8830), .B(p_input[22053]), .Z(o[2053]) );
  AND U17660 ( .A(p_input[2053]), .B(p_input[12053]), .Z(n8830) );
  AND U17661 ( .A(n8831), .B(p_input[22052]), .Z(o[2052]) );
  AND U17662 ( .A(p_input[2052]), .B(p_input[12052]), .Z(n8831) );
  AND U17663 ( .A(n8832), .B(p_input[22051]), .Z(o[2051]) );
  AND U17664 ( .A(p_input[2051]), .B(p_input[12051]), .Z(n8832) );
  AND U17665 ( .A(n8833), .B(p_input[22050]), .Z(o[2050]) );
  AND U17666 ( .A(p_input[2050]), .B(p_input[12050]), .Z(n8833) );
  AND U17667 ( .A(n8834), .B(p_input[204]), .Z(o[204]) );
  AND U17668 ( .A(p_input[20204]), .B(p_input[10204]), .Z(n8834) );
  AND U17669 ( .A(n8835), .B(p_input[22049]), .Z(o[2049]) );
  AND U17670 ( .A(p_input[2049]), .B(p_input[12049]), .Z(n8835) );
  AND U17671 ( .A(n8836), .B(p_input[22048]), .Z(o[2048]) );
  AND U17672 ( .A(p_input[2048]), .B(p_input[12048]), .Z(n8836) );
  AND U17673 ( .A(n8837), .B(p_input[22047]), .Z(o[2047]) );
  AND U17674 ( .A(p_input[2047]), .B(p_input[12047]), .Z(n8837) );
  AND U17675 ( .A(n8838), .B(p_input[22046]), .Z(o[2046]) );
  AND U17676 ( .A(p_input[2046]), .B(p_input[12046]), .Z(n8838) );
  AND U17677 ( .A(n8839), .B(p_input[22045]), .Z(o[2045]) );
  AND U17678 ( .A(p_input[2045]), .B(p_input[12045]), .Z(n8839) );
  AND U17679 ( .A(n8840), .B(p_input[22044]), .Z(o[2044]) );
  AND U17680 ( .A(p_input[2044]), .B(p_input[12044]), .Z(n8840) );
  AND U17681 ( .A(n8841), .B(p_input[22043]), .Z(o[2043]) );
  AND U17682 ( .A(p_input[2043]), .B(p_input[12043]), .Z(n8841) );
  AND U17683 ( .A(n8842), .B(p_input[22042]), .Z(o[2042]) );
  AND U17684 ( .A(p_input[2042]), .B(p_input[12042]), .Z(n8842) );
  AND U17685 ( .A(n8843), .B(p_input[22041]), .Z(o[2041]) );
  AND U17686 ( .A(p_input[2041]), .B(p_input[12041]), .Z(n8843) );
  AND U17687 ( .A(n8844), .B(p_input[22040]), .Z(o[2040]) );
  AND U17688 ( .A(p_input[2040]), .B(p_input[12040]), .Z(n8844) );
  AND U17689 ( .A(n8845), .B(p_input[203]), .Z(o[203]) );
  AND U17690 ( .A(p_input[20203]), .B(p_input[10203]), .Z(n8845) );
  AND U17691 ( .A(n8846), .B(p_input[22039]), .Z(o[2039]) );
  AND U17692 ( .A(p_input[2039]), .B(p_input[12039]), .Z(n8846) );
  AND U17693 ( .A(n8847), .B(p_input[22038]), .Z(o[2038]) );
  AND U17694 ( .A(p_input[2038]), .B(p_input[12038]), .Z(n8847) );
  AND U17695 ( .A(n8848), .B(p_input[22037]), .Z(o[2037]) );
  AND U17696 ( .A(p_input[2037]), .B(p_input[12037]), .Z(n8848) );
  AND U17697 ( .A(n8849), .B(p_input[22036]), .Z(o[2036]) );
  AND U17698 ( .A(p_input[2036]), .B(p_input[12036]), .Z(n8849) );
  AND U17699 ( .A(n8850), .B(p_input[22035]), .Z(o[2035]) );
  AND U17700 ( .A(p_input[2035]), .B(p_input[12035]), .Z(n8850) );
  AND U17701 ( .A(n8851), .B(p_input[22034]), .Z(o[2034]) );
  AND U17702 ( .A(p_input[2034]), .B(p_input[12034]), .Z(n8851) );
  AND U17703 ( .A(n8852), .B(p_input[22033]), .Z(o[2033]) );
  AND U17704 ( .A(p_input[2033]), .B(p_input[12033]), .Z(n8852) );
  AND U17705 ( .A(n8853), .B(p_input[22032]), .Z(o[2032]) );
  AND U17706 ( .A(p_input[2032]), .B(p_input[12032]), .Z(n8853) );
  AND U17707 ( .A(n8854), .B(p_input[22031]), .Z(o[2031]) );
  AND U17708 ( .A(p_input[2031]), .B(p_input[12031]), .Z(n8854) );
  AND U17709 ( .A(n8855), .B(p_input[22030]), .Z(o[2030]) );
  AND U17710 ( .A(p_input[2030]), .B(p_input[12030]), .Z(n8855) );
  AND U17711 ( .A(n8856), .B(p_input[202]), .Z(o[202]) );
  AND U17712 ( .A(p_input[20202]), .B(p_input[10202]), .Z(n8856) );
  AND U17713 ( .A(n8857), .B(p_input[22029]), .Z(o[2029]) );
  AND U17714 ( .A(p_input[2029]), .B(p_input[12029]), .Z(n8857) );
  AND U17715 ( .A(n8858), .B(p_input[22028]), .Z(o[2028]) );
  AND U17716 ( .A(p_input[2028]), .B(p_input[12028]), .Z(n8858) );
  AND U17717 ( .A(n8859), .B(p_input[22027]), .Z(o[2027]) );
  AND U17718 ( .A(p_input[2027]), .B(p_input[12027]), .Z(n8859) );
  AND U17719 ( .A(n8860), .B(p_input[22026]), .Z(o[2026]) );
  AND U17720 ( .A(p_input[2026]), .B(p_input[12026]), .Z(n8860) );
  AND U17721 ( .A(n8861), .B(p_input[22025]), .Z(o[2025]) );
  AND U17722 ( .A(p_input[2025]), .B(p_input[12025]), .Z(n8861) );
  AND U17723 ( .A(n8862), .B(p_input[22024]), .Z(o[2024]) );
  AND U17724 ( .A(p_input[2024]), .B(p_input[12024]), .Z(n8862) );
  AND U17725 ( .A(n8863), .B(p_input[22023]), .Z(o[2023]) );
  AND U17726 ( .A(p_input[2023]), .B(p_input[12023]), .Z(n8863) );
  AND U17727 ( .A(n8864), .B(p_input[22022]), .Z(o[2022]) );
  AND U17728 ( .A(p_input[2022]), .B(p_input[12022]), .Z(n8864) );
  AND U17729 ( .A(n8865), .B(p_input[22021]), .Z(o[2021]) );
  AND U17730 ( .A(p_input[2021]), .B(p_input[12021]), .Z(n8865) );
  AND U17731 ( .A(n8866), .B(p_input[22020]), .Z(o[2020]) );
  AND U17732 ( .A(p_input[2020]), .B(p_input[12020]), .Z(n8866) );
  AND U17733 ( .A(n8867), .B(p_input[20201]), .Z(o[201]) );
  AND U17734 ( .A(p_input[201]), .B(p_input[10201]), .Z(n8867) );
  AND U17735 ( .A(n8868), .B(p_input[22019]), .Z(o[2019]) );
  AND U17736 ( .A(p_input[2019]), .B(p_input[12019]), .Z(n8868) );
  AND U17737 ( .A(n8869), .B(p_input[22018]), .Z(o[2018]) );
  AND U17738 ( .A(p_input[2018]), .B(p_input[12018]), .Z(n8869) );
  AND U17739 ( .A(n8870), .B(p_input[22017]), .Z(o[2017]) );
  AND U17740 ( .A(p_input[2017]), .B(p_input[12017]), .Z(n8870) );
  AND U17741 ( .A(n8871), .B(p_input[22016]), .Z(o[2016]) );
  AND U17742 ( .A(p_input[2016]), .B(p_input[12016]), .Z(n8871) );
  AND U17743 ( .A(n8872), .B(p_input[22015]), .Z(o[2015]) );
  AND U17744 ( .A(p_input[2015]), .B(p_input[12015]), .Z(n8872) );
  AND U17745 ( .A(n8873), .B(p_input[22014]), .Z(o[2014]) );
  AND U17746 ( .A(p_input[2014]), .B(p_input[12014]), .Z(n8873) );
  AND U17747 ( .A(n8874), .B(p_input[22013]), .Z(o[2013]) );
  AND U17748 ( .A(p_input[2013]), .B(p_input[12013]), .Z(n8874) );
  AND U17749 ( .A(n8875), .B(p_input[22012]), .Z(o[2012]) );
  AND U17750 ( .A(p_input[2012]), .B(p_input[12012]), .Z(n8875) );
  AND U17751 ( .A(n8876), .B(p_input[22011]), .Z(o[2011]) );
  AND U17752 ( .A(p_input[2011]), .B(p_input[12011]), .Z(n8876) );
  AND U17753 ( .A(n8877), .B(p_input[22010]), .Z(o[2010]) );
  AND U17754 ( .A(p_input[2010]), .B(p_input[12010]), .Z(n8877) );
  AND U17755 ( .A(n8878), .B(p_input[20200]), .Z(o[200]) );
  AND U17756 ( .A(p_input[200]), .B(p_input[10200]), .Z(n8878) );
  AND U17757 ( .A(n8879), .B(p_input[22009]), .Z(o[2009]) );
  AND U17758 ( .A(p_input[2009]), .B(p_input[12009]), .Z(n8879) );
  AND U17759 ( .A(n8880), .B(p_input[22008]), .Z(o[2008]) );
  AND U17760 ( .A(p_input[2008]), .B(p_input[12008]), .Z(n8880) );
  AND U17761 ( .A(n8881), .B(p_input[22007]), .Z(o[2007]) );
  AND U17762 ( .A(p_input[2007]), .B(p_input[12007]), .Z(n8881) );
  AND U17763 ( .A(n8882), .B(p_input[22006]), .Z(o[2006]) );
  AND U17764 ( .A(p_input[2006]), .B(p_input[12006]), .Z(n8882) );
  AND U17765 ( .A(n8883), .B(p_input[22005]), .Z(o[2005]) );
  AND U17766 ( .A(p_input[2005]), .B(p_input[12005]), .Z(n8883) );
  AND U17767 ( .A(n8884), .B(p_input[22004]), .Z(o[2004]) );
  AND U17768 ( .A(p_input[2004]), .B(p_input[12004]), .Z(n8884) );
  AND U17769 ( .A(n8885), .B(p_input[22003]), .Z(o[2003]) );
  AND U17770 ( .A(p_input[2003]), .B(p_input[12003]), .Z(n8885) );
  AND U17771 ( .A(n8886), .B(p_input[22002]), .Z(o[2002]) );
  AND U17772 ( .A(p_input[2002]), .B(p_input[12002]), .Z(n8886) );
  AND U17773 ( .A(n8887), .B(p_input[22001]), .Z(o[2001]) );
  AND U17774 ( .A(p_input[2001]), .B(p_input[12001]), .Z(n8887) );
  AND U17775 ( .A(n8888), .B(p_input[22000]), .Z(o[2000]) );
  AND U17776 ( .A(p_input[2000]), .B(p_input[12000]), .Z(n8888) );
  AND U17777 ( .A(n8889), .B(p_input[20001]), .Z(o[1]) );
  AND U17778 ( .A(p_input[1]), .B(p_input[10001]), .Z(n8889) );
  AND U17779 ( .A(n8890), .B(p_input[20019]), .Z(o[19]) );
  AND U17780 ( .A(p_input[19]), .B(p_input[10019]), .Z(n8890) );
  AND U17781 ( .A(n8891), .B(p_input[20199]), .Z(o[199]) );
  AND U17782 ( .A(p_input[199]), .B(p_input[10199]), .Z(n8891) );
  AND U17783 ( .A(n8892), .B(p_input[21999]), .Z(o[1999]) );
  AND U17784 ( .A(p_input[1999]), .B(p_input[11999]), .Z(n8892) );
  AND U17785 ( .A(n8893), .B(p_input[21998]), .Z(o[1998]) );
  AND U17786 ( .A(p_input[1998]), .B(p_input[11998]), .Z(n8893) );
  AND U17787 ( .A(n8894), .B(p_input[21997]), .Z(o[1997]) );
  AND U17788 ( .A(p_input[1997]), .B(p_input[11997]), .Z(n8894) );
  AND U17789 ( .A(n8895), .B(p_input[21996]), .Z(o[1996]) );
  AND U17790 ( .A(p_input[1996]), .B(p_input[11996]), .Z(n8895) );
  AND U17791 ( .A(n8896), .B(p_input[21995]), .Z(o[1995]) );
  AND U17792 ( .A(p_input[1995]), .B(p_input[11995]), .Z(n8896) );
  AND U17793 ( .A(n8897), .B(p_input[21994]), .Z(o[1994]) );
  AND U17794 ( .A(p_input[1994]), .B(p_input[11994]), .Z(n8897) );
  AND U17795 ( .A(n8898), .B(p_input[21993]), .Z(o[1993]) );
  AND U17796 ( .A(p_input[1993]), .B(p_input[11993]), .Z(n8898) );
  AND U17797 ( .A(n8899), .B(p_input[21992]), .Z(o[1992]) );
  AND U17798 ( .A(p_input[1992]), .B(p_input[11992]), .Z(n8899) );
  AND U17799 ( .A(n8900), .B(p_input[21991]), .Z(o[1991]) );
  AND U17800 ( .A(p_input[1991]), .B(p_input[11991]), .Z(n8900) );
  AND U17801 ( .A(n8901), .B(p_input[21990]), .Z(o[1990]) );
  AND U17802 ( .A(p_input[1990]), .B(p_input[11990]), .Z(n8901) );
  AND U17803 ( .A(n8902), .B(p_input[20198]), .Z(o[198]) );
  AND U17804 ( .A(p_input[198]), .B(p_input[10198]), .Z(n8902) );
  AND U17805 ( .A(n8903), .B(p_input[21989]), .Z(o[1989]) );
  AND U17806 ( .A(p_input[1989]), .B(p_input[11989]), .Z(n8903) );
  AND U17807 ( .A(n8904), .B(p_input[21988]), .Z(o[1988]) );
  AND U17808 ( .A(p_input[1988]), .B(p_input[11988]), .Z(n8904) );
  AND U17809 ( .A(n8905), .B(p_input[21987]), .Z(o[1987]) );
  AND U17810 ( .A(p_input[1987]), .B(p_input[11987]), .Z(n8905) );
  AND U17811 ( .A(n8906), .B(p_input[21986]), .Z(o[1986]) );
  AND U17812 ( .A(p_input[1986]), .B(p_input[11986]), .Z(n8906) );
  AND U17813 ( .A(n8907), .B(p_input[21985]), .Z(o[1985]) );
  AND U17814 ( .A(p_input[1985]), .B(p_input[11985]), .Z(n8907) );
  AND U17815 ( .A(n8908), .B(p_input[21984]), .Z(o[1984]) );
  AND U17816 ( .A(p_input[1984]), .B(p_input[11984]), .Z(n8908) );
  AND U17817 ( .A(n8909), .B(p_input[21983]), .Z(o[1983]) );
  AND U17818 ( .A(p_input[1983]), .B(p_input[11983]), .Z(n8909) );
  AND U17819 ( .A(n8910), .B(p_input[21982]), .Z(o[1982]) );
  AND U17820 ( .A(p_input[1982]), .B(p_input[11982]), .Z(n8910) );
  AND U17821 ( .A(n8911), .B(p_input[21981]), .Z(o[1981]) );
  AND U17822 ( .A(p_input[1981]), .B(p_input[11981]), .Z(n8911) );
  AND U17823 ( .A(n8912), .B(p_input[21980]), .Z(o[1980]) );
  AND U17824 ( .A(p_input[1980]), .B(p_input[11980]), .Z(n8912) );
  AND U17825 ( .A(n8913), .B(p_input[20197]), .Z(o[197]) );
  AND U17826 ( .A(p_input[197]), .B(p_input[10197]), .Z(n8913) );
  AND U17827 ( .A(n8914), .B(p_input[21979]), .Z(o[1979]) );
  AND U17828 ( .A(p_input[1979]), .B(p_input[11979]), .Z(n8914) );
  AND U17829 ( .A(n8915), .B(p_input[21978]), .Z(o[1978]) );
  AND U17830 ( .A(p_input[1978]), .B(p_input[11978]), .Z(n8915) );
  AND U17831 ( .A(n8916), .B(p_input[21977]), .Z(o[1977]) );
  AND U17832 ( .A(p_input[1977]), .B(p_input[11977]), .Z(n8916) );
  AND U17833 ( .A(n8917), .B(p_input[21976]), .Z(o[1976]) );
  AND U17834 ( .A(p_input[1976]), .B(p_input[11976]), .Z(n8917) );
  AND U17835 ( .A(n8918), .B(p_input[21975]), .Z(o[1975]) );
  AND U17836 ( .A(p_input[1975]), .B(p_input[11975]), .Z(n8918) );
  AND U17837 ( .A(n8919), .B(p_input[21974]), .Z(o[1974]) );
  AND U17838 ( .A(p_input[1974]), .B(p_input[11974]), .Z(n8919) );
  AND U17839 ( .A(n8920), .B(p_input[21973]), .Z(o[1973]) );
  AND U17840 ( .A(p_input[1973]), .B(p_input[11973]), .Z(n8920) );
  AND U17841 ( .A(n8921), .B(p_input[21972]), .Z(o[1972]) );
  AND U17842 ( .A(p_input[1972]), .B(p_input[11972]), .Z(n8921) );
  AND U17843 ( .A(n8922), .B(p_input[21971]), .Z(o[1971]) );
  AND U17844 ( .A(p_input[1971]), .B(p_input[11971]), .Z(n8922) );
  AND U17845 ( .A(n8923), .B(p_input[21970]), .Z(o[1970]) );
  AND U17846 ( .A(p_input[1970]), .B(p_input[11970]), .Z(n8923) );
  AND U17847 ( .A(n8924), .B(p_input[20196]), .Z(o[196]) );
  AND U17848 ( .A(p_input[196]), .B(p_input[10196]), .Z(n8924) );
  AND U17849 ( .A(n8925), .B(p_input[21969]), .Z(o[1969]) );
  AND U17850 ( .A(p_input[1969]), .B(p_input[11969]), .Z(n8925) );
  AND U17851 ( .A(n8926), .B(p_input[21968]), .Z(o[1968]) );
  AND U17852 ( .A(p_input[1968]), .B(p_input[11968]), .Z(n8926) );
  AND U17853 ( .A(n8927), .B(p_input[21967]), .Z(o[1967]) );
  AND U17854 ( .A(p_input[1967]), .B(p_input[11967]), .Z(n8927) );
  AND U17855 ( .A(n8928), .B(p_input[21966]), .Z(o[1966]) );
  AND U17856 ( .A(p_input[1966]), .B(p_input[11966]), .Z(n8928) );
  AND U17857 ( .A(n8929), .B(p_input[21965]), .Z(o[1965]) );
  AND U17858 ( .A(p_input[1965]), .B(p_input[11965]), .Z(n8929) );
  AND U17859 ( .A(n8930), .B(p_input[21964]), .Z(o[1964]) );
  AND U17860 ( .A(p_input[1964]), .B(p_input[11964]), .Z(n8930) );
  AND U17861 ( .A(n8931), .B(p_input[21963]), .Z(o[1963]) );
  AND U17862 ( .A(p_input[1963]), .B(p_input[11963]), .Z(n8931) );
  AND U17863 ( .A(n8932), .B(p_input[21962]), .Z(o[1962]) );
  AND U17864 ( .A(p_input[1962]), .B(p_input[11962]), .Z(n8932) );
  AND U17865 ( .A(n8933), .B(p_input[21961]), .Z(o[1961]) );
  AND U17866 ( .A(p_input[1961]), .B(p_input[11961]), .Z(n8933) );
  AND U17867 ( .A(n8934), .B(p_input[21960]), .Z(o[1960]) );
  AND U17868 ( .A(p_input[1960]), .B(p_input[11960]), .Z(n8934) );
  AND U17869 ( .A(n8935), .B(p_input[20195]), .Z(o[195]) );
  AND U17870 ( .A(p_input[195]), .B(p_input[10195]), .Z(n8935) );
  AND U17871 ( .A(n8936), .B(p_input[21959]), .Z(o[1959]) );
  AND U17872 ( .A(p_input[1959]), .B(p_input[11959]), .Z(n8936) );
  AND U17873 ( .A(n8937), .B(p_input[21958]), .Z(o[1958]) );
  AND U17874 ( .A(p_input[1958]), .B(p_input[11958]), .Z(n8937) );
  AND U17875 ( .A(n8938), .B(p_input[21957]), .Z(o[1957]) );
  AND U17876 ( .A(p_input[1957]), .B(p_input[11957]), .Z(n8938) );
  AND U17877 ( .A(n8939), .B(p_input[21956]), .Z(o[1956]) );
  AND U17878 ( .A(p_input[1956]), .B(p_input[11956]), .Z(n8939) );
  AND U17879 ( .A(n8940), .B(p_input[21955]), .Z(o[1955]) );
  AND U17880 ( .A(p_input[1955]), .B(p_input[11955]), .Z(n8940) );
  AND U17881 ( .A(n8941), .B(p_input[21954]), .Z(o[1954]) );
  AND U17882 ( .A(p_input[1954]), .B(p_input[11954]), .Z(n8941) );
  AND U17883 ( .A(n8942), .B(p_input[21953]), .Z(o[1953]) );
  AND U17884 ( .A(p_input[1953]), .B(p_input[11953]), .Z(n8942) );
  AND U17885 ( .A(n8943), .B(p_input[21952]), .Z(o[1952]) );
  AND U17886 ( .A(p_input[1952]), .B(p_input[11952]), .Z(n8943) );
  AND U17887 ( .A(n8944), .B(p_input[21951]), .Z(o[1951]) );
  AND U17888 ( .A(p_input[1951]), .B(p_input[11951]), .Z(n8944) );
  AND U17889 ( .A(n8945), .B(p_input[21950]), .Z(o[1950]) );
  AND U17890 ( .A(p_input[1950]), .B(p_input[11950]), .Z(n8945) );
  AND U17891 ( .A(n8946), .B(p_input[20194]), .Z(o[194]) );
  AND U17892 ( .A(p_input[194]), .B(p_input[10194]), .Z(n8946) );
  AND U17893 ( .A(n8947), .B(p_input[21949]), .Z(o[1949]) );
  AND U17894 ( .A(p_input[1949]), .B(p_input[11949]), .Z(n8947) );
  AND U17895 ( .A(n8948), .B(p_input[21948]), .Z(o[1948]) );
  AND U17896 ( .A(p_input[1948]), .B(p_input[11948]), .Z(n8948) );
  AND U17897 ( .A(n8949), .B(p_input[21947]), .Z(o[1947]) );
  AND U17898 ( .A(p_input[1947]), .B(p_input[11947]), .Z(n8949) );
  AND U17899 ( .A(n8950), .B(p_input[21946]), .Z(o[1946]) );
  AND U17900 ( .A(p_input[1946]), .B(p_input[11946]), .Z(n8950) );
  AND U17901 ( .A(n8951), .B(p_input[21945]), .Z(o[1945]) );
  AND U17902 ( .A(p_input[1945]), .B(p_input[11945]), .Z(n8951) );
  AND U17903 ( .A(n8952), .B(p_input[21944]), .Z(o[1944]) );
  AND U17904 ( .A(p_input[1944]), .B(p_input[11944]), .Z(n8952) );
  AND U17905 ( .A(n8953), .B(p_input[21943]), .Z(o[1943]) );
  AND U17906 ( .A(p_input[1943]), .B(p_input[11943]), .Z(n8953) );
  AND U17907 ( .A(n8954), .B(p_input[21942]), .Z(o[1942]) );
  AND U17908 ( .A(p_input[1942]), .B(p_input[11942]), .Z(n8954) );
  AND U17909 ( .A(n8955), .B(p_input[21941]), .Z(o[1941]) );
  AND U17910 ( .A(p_input[1941]), .B(p_input[11941]), .Z(n8955) );
  AND U17911 ( .A(n8956), .B(p_input[21940]), .Z(o[1940]) );
  AND U17912 ( .A(p_input[1940]), .B(p_input[11940]), .Z(n8956) );
  AND U17913 ( .A(n8957), .B(p_input[20193]), .Z(o[193]) );
  AND U17914 ( .A(p_input[193]), .B(p_input[10193]), .Z(n8957) );
  AND U17915 ( .A(n8958), .B(p_input[21939]), .Z(o[1939]) );
  AND U17916 ( .A(p_input[1939]), .B(p_input[11939]), .Z(n8958) );
  AND U17917 ( .A(n8959), .B(p_input[21938]), .Z(o[1938]) );
  AND U17918 ( .A(p_input[1938]), .B(p_input[11938]), .Z(n8959) );
  AND U17919 ( .A(n8960), .B(p_input[21937]), .Z(o[1937]) );
  AND U17920 ( .A(p_input[1937]), .B(p_input[11937]), .Z(n8960) );
  AND U17921 ( .A(n8961), .B(p_input[21936]), .Z(o[1936]) );
  AND U17922 ( .A(p_input[1936]), .B(p_input[11936]), .Z(n8961) );
  AND U17923 ( .A(n8962), .B(p_input[21935]), .Z(o[1935]) );
  AND U17924 ( .A(p_input[1935]), .B(p_input[11935]), .Z(n8962) );
  AND U17925 ( .A(n8963), .B(p_input[21934]), .Z(o[1934]) );
  AND U17926 ( .A(p_input[1934]), .B(p_input[11934]), .Z(n8963) );
  AND U17927 ( .A(n8964), .B(p_input[21933]), .Z(o[1933]) );
  AND U17928 ( .A(p_input[1933]), .B(p_input[11933]), .Z(n8964) );
  AND U17929 ( .A(n8965), .B(p_input[21932]), .Z(o[1932]) );
  AND U17930 ( .A(p_input[1932]), .B(p_input[11932]), .Z(n8965) );
  AND U17931 ( .A(n8966), .B(p_input[21931]), .Z(o[1931]) );
  AND U17932 ( .A(p_input[1931]), .B(p_input[11931]), .Z(n8966) );
  AND U17933 ( .A(n8967), .B(p_input[21930]), .Z(o[1930]) );
  AND U17934 ( .A(p_input[1930]), .B(p_input[11930]), .Z(n8967) );
  AND U17935 ( .A(n8968), .B(p_input[20192]), .Z(o[192]) );
  AND U17936 ( .A(p_input[192]), .B(p_input[10192]), .Z(n8968) );
  AND U17937 ( .A(n8969), .B(p_input[21929]), .Z(o[1929]) );
  AND U17938 ( .A(p_input[1929]), .B(p_input[11929]), .Z(n8969) );
  AND U17939 ( .A(n8970), .B(p_input[21928]), .Z(o[1928]) );
  AND U17940 ( .A(p_input[1928]), .B(p_input[11928]), .Z(n8970) );
  AND U17941 ( .A(n8971), .B(p_input[21927]), .Z(o[1927]) );
  AND U17942 ( .A(p_input[1927]), .B(p_input[11927]), .Z(n8971) );
  AND U17943 ( .A(n8972), .B(p_input[21926]), .Z(o[1926]) );
  AND U17944 ( .A(p_input[1926]), .B(p_input[11926]), .Z(n8972) );
  AND U17945 ( .A(n8973), .B(p_input[21925]), .Z(o[1925]) );
  AND U17946 ( .A(p_input[1925]), .B(p_input[11925]), .Z(n8973) );
  AND U17947 ( .A(n8974), .B(p_input[21924]), .Z(o[1924]) );
  AND U17948 ( .A(p_input[1924]), .B(p_input[11924]), .Z(n8974) );
  AND U17949 ( .A(n8975), .B(p_input[21923]), .Z(o[1923]) );
  AND U17950 ( .A(p_input[1923]), .B(p_input[11923]), .Z(n8975) );
  AND U17951 ( .A(n8976), .B(p_input[21922]), .Z(o[1922]) );
  AND U17952 ( .A(p_input[1922]), .B(p_input[11922]), .Z(n8976) );
  AND U17953 ( .A(n8977), .B(p_input[21921]), .Z(o[1921]) );
  AND U17954 ( .A(p_input[1921]), .B(p_input[11921]), .Z(n8977) );
  AND U17955 ( .A(n8978), .B(p_input[21920]), .Z(o[1920]) );
  AND U17956 ( .A(p_input[1920]), .B(p_input[11920]), .Z(n8978) );
  AND U17957 ( .A(n8979), .B(p_input[20191]), .Z(o[191]) );
  AND U17958 ( .A(p_input[191]), .B(p_input[10191]), .Z(n8979) );
  AND U17959 ( .A(n8980), .B(p_input[21919]), .Z(o[1919]) );
  AND U17960 ( .A(p_input[1919]), .B(p_input[11919]), .Z(n8980) );
  AND U17961 ( .A(n8981), .B(p_input[21918]), .Z(o[1918]) );
  AND U17962 ( .A(p_input[1918]), .B(p_input[11918]), .Z(n8981) );
  AND U17963 ( .A(n8982), .B(p_input[21917]), .Z(o[1917]) );
  AND U17964 ( .A(p_input[1917]), .B(p_input[11917]), .Z(n8982) );
  AND U17965 ( .A(n8983), .B(p_input[21916]), .Z(o[1916]) );
  AND U17966 ( .A(p_input[1916]), .B(p_input[11916]), .Z(n8983) );
  AND U17967 ( .A(n8984), .B(p_input[21915]), .Z(o[1915]) );
  AND U17968 ( .A(p_input[1915]), .B(p_input[11915]), .Z(n8984) );
  AND U17969 ( .A(n8985), .B(p_input[21914]), .Z(o[1914]) );
  AND U17970 ( .A(p_input[1914]), .B(p_input[11914]), .Z(n8985) );
  AND U17971 ( .A(n8986), .B(p_input[21913]), .Z(o[1913]) );
  AND U17972 ( .A(p_input[1913]), .B(p_input[11913]), .Z(n8986) );
  AND U17973 ( .A(n8987), .B(p_input[21912]), .Z(o[1912]) );
  AND U17974 ( .A(p_input[1912]), .B(p_input[11912]), .Z(n8987) );
  AND U17975 ( .A(n8988), .B(p_input[21911]), .Z(o[1911]) );
  AND U17976 ( .A(p_input[1911]), .B(p_input[11911]), .Z(n8988) );
  AND U17977 ( .A(n8989), .B(p_input[21910]), .Z(o[1910]) );
  AND U17978 ( .A(p_input[1910]), .B(p_input[11910]), .Z(n8989) );
  AND U17979 ( .A(n8990), .B(p_input[20190]), .Z(o[190]) );
  AND U17980 ( .A(p_input[190]), .B(p_input[10190]), .Z(n8990) );
  AND U17981 ( .A(n8991), .B(p_input[21909]), .Z(o[1909]) );
  AND U17982 ( .A(p_input[1909]), .B(p_input[11909]), .Z(n8991) );
  AND U17983 ( .A(n8992), .B(p_input[21908]), .Z(o[1908]) );
  AND U17984 ( .A(p_input[1908]), .B(p_input[11908]), .Z(n8992) );
  AND U17985 ( .A(n8993), .B(p_input[21907]), .Z(o[1907]) );
  AND U17986 ( .A(p_input[1907]), .B(p_input[11907]), .Z(n8993) );
  AND U17987 ( .A(n8994), .B(p_input[21906]), .Z(o[1906]) );
  AND U17988 ( .A(p_input[1906]), .B(p_input[11906]), .Z(n8994) );
  AND U17989 ( .A(n8995), .B(p_input[21905]), .Z(o[1905]) );
  AND U17990 ( .A(p_input[1905]), .B(p_input[11905]), .Z(n8995) );
  AND U17991 ( .A(n8996), .B(p_input[21904]), .Z(o[1904]) );
  AND U17992 ( .A(p_input[1904]), .B(p_input[11904]), .Z(n8996) );
  AND U17993 ( .A(n8997), .B(p_input[21903]), .Z(o[1903]) );
  AND U17994 ( .A(p_input[1903]), .B(p_input[11903]), .Z(n8997) );
  AND U17995 ( .A(n8998), .B(p_input[21902]), .Z(o[1902]) );
  AND U17996 ( .A(p_input[1902]), .B(p_input[11902]), .Z(n8998) );
  AND U17997 ( .A(n8999), .B(p_input[21901]), .Z(o[1901]) );
  AND U17998 ( .A(p_input[1901]), .B(p_input[11901]), .Z(n8999) );
  AND U17999 ( .A(n9000), .B(p_input[21900]), .Z(o[1900]) );
  AND U18000 ( .A(p_input[1900]), .B(p_input[11900]), .Z(n9000) );
  AND U18001 ( .A(n9001), .B(p_input[20018]), .Z(o[18]) );
  AND U18002 ( .A(p_input[18]), .B(p_input[10018]), .Z(n9001) );
  AND U18003 ( .A(n9002), .B(p_input[20189]), .Z(o[189]) );
  AND U18004 ( .A(p_input[189]), .B(p_input[10189]), .Z(n9002) );
  AND U18005 ( .A(n9003), .B(p_input[21899]), .Z(o[1899]) );
  AND U18006 ( .A(p_input[1899]), .B(p_input[11899]), .Z(n9003) );
  AND U18007 ( .A(n9004), .B(p_input[21898]), .Z(o[1898]) );
  AND U18008 ( .A(p_input[1898]), .B(p_input[11898]), .Z(n9004) );
  AND U18009 ( .A(n9005), .B(p_input[21897]), .Z(o[1897]) );
  AND U18010 ( .A(p_input[1897]), .B(p_input[11897]), .Z(n9005) );
  AND U18011 ( .A(n9006), .B(p_input[21896]), .Z(o[1896]) );
  AND U18012 ( .A(p_input[1896]), .B(p_input[11896]), .Z(n9006) );
  AND U18013 ( .A(n9007), .B(p_input[21895]), .Z(o[1895]) );
  AND U18014 ( .A(p_input[1895]), .B(p_input[11895]), .Z(n9007) );
  AND U18015 ( .A(n9008), .B(p_input[21894]), .Z(o[1894]) );
  AND U18016 ( .A(p_input[1894]), .B(p_input[11894]), .Z(n9008) );
  AND U18017 ( .A(n9009), .B(p_input[21893]), .Z(o[1893]) );
  AND U18018 ( .A(p_input[1893]), .B(p_input[11893]), .Z(n9009) );
  AND U18019 ( .A(n9010), .B(p_input[21892]), .Z(o[1892]) );
  AND U18020 ( .A(p_input[1892]), .B(p_input[11892]), .Z(n9010) );
  AND U18021 ( .A(n9011), .B(p_input[21891]), .Z(o[1891]) );
  AND U18022 ( .A(p_input[1891]), .B(p_input[11891]), .Z(n9011) );
  AND U18023 ( .A(n9012), .B(p_input[21890]), .Z(o[1890]) );
  AND U18024 ( .A(p_input[1890]), .B(p_input[11890]), .Z(n9012) );
  AND U18025 ( .A(n9013), .B(p_input[20188]), .Z(o[188]) );
  AND U18026 ( .A(p_input[188]), .B(p_input[10188]), .Z(n9013) );
  AND U18027 ( .A(n9014), .B(p_input[21889]), .Z(o[1889]) );
  AND U18028 ( .A(p_input[1889]), .B(p_input[11889]), .Z(n9014) );
  AND U18029 ( .A(n9015), .B(p_input[21888]), .Z(o[1888]) );
  AND U18030 ( .A(p_input[1888]), .B(p_input[11888]), .Z(n9015) );
  AND U18031 ( .A(n9016), .B(p_input[21887]), .Z(o[1887]) );
  AND U18032 ( .A(p_input[1887]), .B(p_input[11887]), .Z(n9016) );
  AND U18033 ( .A(n9017), .B(p_input[21886]), .Z(o[1886]) );
  AND U18034 ( .A(p_input[1886]), .B(p_input[11886]), .Z(n9017) );
  AND U18035 ( .A(n9018), .B(p_input[21885]), .Z(o[1885]) );
  AND U18036 ( .A(p_input[1885]), .B(p_input[11885]), .Z(n9018) );
  AND U18037 ( .A(n9019), .B(p_input[21884]), .Z(o[1884]) );
  AND U18038 ( .A(p_input[1884]), .B(p_input[11884]), .Z(n9019) );
  AND U18039 ( .A(n9020), .B(p_input[21883]), .Z(o[1883]) );
  AND U18040 ( .A(p_input[1883]), .B(p_input[11883]), .Z(n9020) );
  AND U18041 ( .A(n9021), .B(p_input[21882]), .Z(o[1882]) );
  AND U18042 ( .A(p_input[1882]), .B(p_input[11882]), .Z(n9021) );
  AND U18043 ( .A(n9022), .B(p_input[21881]), .Z(o[1881]) );
  AND U18044 ( .A(p_input[1881]), .B(p_input[11881]), .Z(n9022) );
  AND U18045 ( .A(n9023), .B(p_input[21880]), .Z(o[1880]) );
  AND U18046 ( .A(p_input[1880]), .B(p_input[11880]), .Z(n9023) );
  AND U18047 ( .A(n9024), .B(p_input[20187]), .Z(o[187]) );
  AND U18048 ( .A(p_input[187]), .B(p_input[10187]), .Z(n9024) );
  AND U18049 ( .A(n9025), .B(p_input[21879]), .Z(o[1879]) );
  AND U18050 ( .A(p_input[1879]), .B(p_input[11879]), .Z(n9025) );
  AND U18051 ( .A(n9026), .B(p_input[21878]), .Z(o[1878]) );
  AND U18052 ( .A(p_input[1878]), .B(p_input[11878]), .Z(n9026) );
  AND U18053 ( .A(n9027), .B(p_input[21877]), .Z(o[1877]) );
  AND U18054 ( .A(p_input[1877]), .B(p_input[11877]), .Z(n9027) );
  AND U18055 ( .A(n9028), .B(p_input[21876]), .Z(o[1876]) );
  AND U18056 ( .A(p_input[1876]), .B(p_input[11876]), .Z(n9028) );
  AND U18057 ( .A(n9029), .B(p_input[21875]), .Z(o[1875]) );
  AND U18058 ( .A(p_input[1875]), .B(p_input[11875]), .Z(n9029) );
  AND U18059 ( .A(n9030), .B(p_input[21874]), .Z(o[1874]) );
  AND U18060 ( .A(p_input[1874]), .B(p_input[11874]), .Z(n9030) );
  AND U18061 ( .A(n9031), .B(p_input[21873]), .Z(o[1873]) );
  AND U18062 ( .A(p_input[1873]), .B(p_input[11873]), .Z(n9031) );
  AND U18063 ( .A(n9032), .B(p_input[21872]), .Z(o[1872]) );
  AND U18064 ( .A(p_input[1872]), .B(p_input[11872]), .Z(n9032) );
  AND U18065 ( .A(n9033), .B(p_input[21871]), .Z(o[1871]) );
  AND U18066 ( .A(p_input[1871]), .B(p_input[11871]), .Z(n9033) );
  AND U18067 ( .A(n9034), .B(p_input[21870]), .Z(o[1870]) );
  AND U18068 ( .A(p_input[1870]), .B(p_input[11870]), .Z(n9034) );
  AND U18069 ( .A(n9035), .B(p_input[20186]), .Z(o[186]) );
  AND U18070 ( .A(p_input[186]), .B(p_input[10186]), .Z(n9035) );
  AND U18071 ( .A(n9036), .B(p_input[21869]), .Z(o[1869]) );
  AND U18072 ( .A(p_input[1869]), .B(p_input[11869]), .Z(n9036) );
  AND U18073 ( .A(n9037), .B(p_input[21868]), .Z(o[1868]) );
  AND U18074 ( .A(p_input[1868]), .B(p_input[11868]), .Z(n9037) );
  AND U18075 ( .A(n9038), .B(p_input[21867]), .Z(o[1867]) );
  AND U18076 ( .A(p_input[1867]), .B(p_input[11867]), .Z(n9038) );
  AND U18077 ( .A(n9039), .B(p_input[21866]), .Z(o[1866]) );
  AND U18078 ( .A(p_input[1866]), .B(p_input[11866]), .Z(n9039) );
  AND U18079 ( .A(n9040), .B(p_input[21865]), .Z(o[1865]) );
  AND U18080 ( .A(p_input[1865]), .B(p_input[11865]), .Z(n9040) );
  AND U18081 ( .A(n9041), .B(p_input[21864]), .Z(o[1864]) );
  AND U18082 ( .A(p_input[1864]), .B(p_input[11864]), .Z(n9041) );
  AND U18083 ( .A(n9042), .B(p_input[21863]), .Z(o[1863]) );
  AND U18084 ( .A(p_input[1863]), .B(p_input[11863]), .Z(n9042) );
  AND U18085 ( .A(n9043), .B(p_input[21862]), .Z(o[1862]) );
  AND U18086 ( .A(p_input[1862]), .B(p_input[11862]), .Z(n9043) );
  AND U18087 ( .A(n9044), .B(p_input[21861]), .Z(o[1861]) );
  AND U18088 ( .A(p_input[1861]), .B(p_input[11861]), .Z(n9044) );
  AND U18089 ( .A(n9045), .B(p_input[21860]), .Z(o[1860]) );
  AND U18090 ( .A(p_input[1860]), .B(p_input[11860]), .Z(n9045) );
  AND U18091 ( .A(n9046), .B(p_input[20185]), .Z(o[185]) );
  AND U18092 ( .A(p_input[185]), .B(p_input[10185]), .Z(n9046) );
  AND U18093 ( .A(n9047), .B(p_input[21859]), .Z(o[1859]) );
  AND U18094 ( .A(p_input[1859]), .B(p_input[11859]), .Z(n9047) );
  AND U18095 ( .A(n9048), .B(p_input[21858]), .Z(o[1858]) );
  AND U18096 ( .A(p_input[1858]), .B(p_input[11858]), .Z(n9048) );
  AND U18097 ( .A(n9049), .B(p_input[21857]), .Z(o[1857]) );
  AND U18098 ( .A(p_input[1857]), .B(p_input[11857]), .Z(n9049) );
  AND U18099 ( .A(n9050), .B(p_input[21856]), .Z(o[1856]) );
  AND U18100 ( .A(p_input[1856]), .B(p_input[11856]), .Z(n9050) );
  AND U18101 ( .A(n9051), .B(p_input[21855]), .Z(o[1855]) );
  AND U18102 ( .A(p_input[1855]), .B(p_input[11855]), .Z(n9051) );
  AND U18103 ( .A(n9052), .B(p_input[21854]), .Z(o[1854]) );
  AND U18104 ( .A(p_input[1854]), .B(p_input[11854]), .Z(n9052) );
  AND U18105 ( .A(n9053), .B(p_input[21853]), .Z(o[1853]) );
  AND U18106 ( .A(p_input[1853]), .B(p_input[11853]), .Z(n9053) );
  AND U18107 ( .A(n9054), .B(p_input[21852]), .Z(o[1852]) );
  AND U18108 ( .A(p_input[1852]), .B(p_input[11852]), .Z(n9054) );
  AND U18109 ( .A(n9055), .B(p_input[21851]), .Z(o[1851]) );
  AND U18110 ( .A(p_input[1851]), .B(p_input[11851]), .Z(n9055) );
  AND U18111 ( .A(n9056), .B(p_input[21850]), .Z(o[1850]) );
  AND U18112 ( .A(p_input[1850]), .B(p_input[11850]), .Z(n9056) );
  AND U18113 ( .A(n9057), .B(p_input[20184]), .Z(o[184]) );
  AND U18114 ( .A(p_input[184]), .B(p_input[10184]), .Z(n9057) );
  AND U18115 ( .A(n9058), .B(p_input[21849]), .Z(o[1849]) );
  AND U18116 ( .A(p_input[1849]), .B(p_input[11849]), .Z(n9058) );
  AND U18117 ( .A(n9059), .B(p_input[21848]), .Z(o[1848]) );
  AND U18118 ( .A(p_input[1848]), .B(p_input[11848]), .Z(n9059) );
  AND U18119 ( .A(n9060), .B(p_input[21847]), .Z(o[1847]) );
  AND U18120 ( .A(p_input[1847]), .B(p_input[11847]), .Z(n9060) );
  AND U18121 ( .A(n9061), .B(p_input[21846]), .Z(o[1846]) );
  AND U18122 ( .A(p_input[1846]), .B(p_input[11846]), .Z(n9061) );
  AND U18123 ( .A(n9062), .B(p_input[21845]), .Z(o[1845]) );
  AND U18124 ( .A(p_input[1845]), .B(p_input[11845]), .Z(n9062) );
  AND U18125 ( .A(n9063), .B(p_input[21844]), .Z(o[1844]) );
  AND U18126 ( .A(p_input[1844]), .B(p_input[11844]), .Z(n9063) );
  AND U18127 ( .A(n9064), .B(p_input[21843]), .Z(o[1843]) );
  AND U18128 ( .A(p_input[1843]), .B(p_input[11843]), .Z(n9064) );
  AND U18129 ( .A(n9065), .B(p_input[21842]), .Z(o[1842]) );
  AND U18130 ( .A(p_input[1842]), .B(p_input[11842]), .Z(n9065) );
  AND U18131 ( .A(n9066), .B(p_input[21841]), .Z(o[1841]) );
  AND U18132 ( .A(p_input[1841]), .B(p_input[11841]), .Z(n9066) );
  AND U18133 ( .A(n9067), .B(p_input[21840]), .Z(o[1840]) );
  AND U18134 ( .A(p_input[1840]), .B(p_input[11840]), .Z(n9067) );
  AND U18135 ( .A(n9068), .B(p_input[20183]), .Z(o[183]) );
  AND U18136 ( .A(p_input[183]), .B(p_input[10183]), .Z(n9068) );
  AND U18137 ( .A(n9069), .B(p_input[21839]), .Z(o[1839]) );
  AND U18138 ( .A(p_input[1839]), .B(p_input[11839]), .Z(n9069) );
  AND U18139 ( .A(n9070), .B(p_input[21838]), .Z(o[1838]) );
  AND U18140 ( .A(p_input[1838]), .B(p_input[11838]), .Z(n9070) );
  AND U18141 ( .A(n9071), .B(p_input[21837]), .Z(o[1837]) );
  AND U18142 ( .A(p_input[1837]), .B(p_input[11837]), .Z(n9071) );
  AND U18143 ( .A(n9072), .B(p_input[21836]), .Z(o[1836]) );
  AND U18144 ( .A(p_input[1836]), .B(p_input[11836]), .Z(n9072) );
  AND U18145 ( .A(n9073), .B(p_input[21835]), .Z(o[1835]) );
  AND U18146 ( .A(p_input[1835]), .B(p_input[11835]), .Z(n9073) );
  AND U18147 ( .A(n9074), .B(p_input[21834]), .Z(o[1834]) );
  AND U18148 ( .A(p_input[1834]), .B(p_input[11834]), .Z(n9074) );
  AND U18149 ( .A(n9075), .B(p_input[21833]), .Z(o[1833]) );
  AND U18150 ( .A(p_input[1833]), .B(p_input[11833]), .Z(n9075) );
  AND U18151 ( .A(n9076), .B(p_input[21832]), .Z(o[1832]) );
  AND U18152 ( .A(p_input[1832]), .B(p_input[11832]), .Z(n9076) );
  AND U18153 ( .A(n9077), .B(p_input[21831]), .Z(o[1831]) );
  AND U18154 ( .A(p_input[1831]), .B(p_input[11831]), .Z(n9077) );
  AND U18155 ( .A(n9078), .B(p_input[21830]), .Z(o[1830]) );
  AND U18156 ( .A(p_input[1830]), .B(p_input[11830]), .Z(n9078) );
  AND U18157 ( .A(n9079), .B(p_input[20182]), .Z(o[182]) );
  AND U18158 ( .A(p_input[182]), .B(p_input[10182]), .Z(n9079) );
  AND U18159 ( .A(n9080), .B(p_input[21829]), .Z(o[1829]) );
  AND U18160 ( .A(p_input[1829]), .B(p_input[11829]), .Z(n9080) );
  AND U18161 ( .A(n9081), .B(p_input[21828]), .Z(o[1828]) );
  AND U18162 ( .A(p_input[1828]), .B(p_input[11828]), .Z(n9081) );
  AND U18163 ( .A(n9082), .B(p_input[21827]), .Z(o[1827]) );
  AND U18164 ( .A(p_input[1827]), .B(p_input[11827]), .Z(n9082) );
  AND U18165 ( .A(n9083), .B(p_input[21826]), .Z(o[1826]) );
  AND U18166 ( .A(p_input[1826]), .B(p_input[11826]), .Z(n9083) );
  AND U18167 ( .A(n9084), .B(p_input[21825]), .Z(o[1825]) );
  AND U18168 ( .A(p_input[1825]), .B(p_input[11825]), .Z(n9084) );
  AND U18169 ( .A(n9085), .B(p_input[21824]), .Z(o[1824]) );
  AND U18170 ( .A(p_input[1824]), .B(p_input[11824]), .Z(n9085) );
  AND U18171 ( .A(n9086), .B(p_input[21823]), .Z(o[1823]) );
  AND U18172 ( .A(p_input[1823]), .B(p_input[11823]), .Z(n9086) );
  AND U18173 ( .A(n9087), .B(p_input[21822]), .Z(o[1822]) );
  AND U18174 ( .A(p_input[1822]), .B(p_input[11822]), .Z(n9087) );
  AND U18175 ( .A(n9088), .B(p_input[21821]), .Z(o[1821]) );
  AND U18176 ( .A(p_input[1821]), .B(p_input[11821]), .Z(n9088) );
  AND U18177 ( .A(n9089), .B(p_input[21820]), .Z(o[1820]) );
  AND U18178 ( .A(p_input[1820]), .B(p_input[11820]), .Z(n9089) );
  AND U18179 ( .A(n9090), .B(p_input[20181]), .Z(o[181]) );
  AND U18180 ( .A(p_input[181]), .B(p_input[10181]), .Z(n9090) );
  AND U18181 ( .A(n9091), .B(p_input[21819]), .Z(o[1819]) );
  AND U18182 ( .A(p_input[1819]), .B(p_input[11819]), .Z(n9091) );
  AND U18183 ( .A(n9092), .B(p_input[21818]), .Z(o[1818]) );
  AND U18184 ( .A(p_input[1818]), .B(p_input[11818]), .Z(n9092) );
  AND U18185 ( .A(n9093), .B(p_input[21817]), .Z(o[1817]) );
  AND U18186 ( .A(p_input[1817]), .B(p_input[11817]), .Z(n9093) );
  AND U18187 ( .A(n9094), .B(p_input[21816]), .Z(o[1816]) );
  AND U18188 ( .A(p_input[1816]), .B(p_input[11816]), .Z(n9094) );
  AND U18189 ( .A(n9095), .B(p_input[21815]), .Z(o[1815]) );
  AND U18190 ( .A(p_input[1815]), .B(p_input[11815]), .Z(n9095) );
  AND U18191 ( .A(n9096), .B(p_input[21814]), .Z(o[1814]) );
  AND U18192 ( .A(p_input[1814]), .B(p_input[11814]), .Z(n9096) );
  AND U18193 ( .A(n9097), .B(p_input[21813]), .Z(o[1813]) );
  AND U18194 ( .A(p_input[1813]), .B(p_input[11813]), .Z(n9097) );
  AND U18195 ( .A(n9098), .B(p_input[21812]), .Z(o[1812]) );
  AND U18196 ( .A(p_input[1812]), .B(p_input[11812]), .Z(n9098) );
  AND U18197 ( .A(n9099), .B(p_input[21811]), .Z(o[1811]) );
  AND U18198 ( .A(p_input[1811]), .B(p_input[11811]), .Z(n9099) );
  AND U18199 ( .A(n9100), .B(p_input[21810]), .Z(o[1810]) );
  AND U18200 ( .A(p_input[1810]), .B(p_input[11810]), .Z(n9100) );
  AND U18201 ( .A(n9101), .B(p_input[20180]), .Z(o[180]) );
  AND U18202 ( .A(p_input[180]), .B(p_input[10180]), .Z(n9101) );
  AND U18203 ( .A(n9102), .B(p_input[21809]), .Z(o[1809]) );
  AND U18204 ( .A(p_input[1809]), .B(p_input[11809]), .Z(n9102) );
  AND U18205 ( .A(n9103), .B(p_input[21808]), .Z(o[1808]) );
  AND U18206 ( .A(p_input[1808]), .B(p_input[11808]), .Z(n9103) );
  AND U18207 ( .A(n9104), .B(p_input[21807]), .Z(o[1807]) );
  AND U18208 ( .A(p_input[1807]), .B(p_input[11807]), .Z(n9104) );
  AND U18209 ( .A(n9105), .B(p_input[21806]), .Z(o[1806]) );
  AND U18210 ( .A(p_input[1806]), .B(p_input[11806]), .Z(n9105) );
  AND U18211 ( .A(n9106), .B(p_input[21805]), .Z(o[1805]) );
  AND U18212 ( .A(p_input[1805]), .B(p_input[11805]), .Z(n9106) );
  AND U18213 ( .A(n9107), .B(p_input[21804]), .Z(o[1804]) );
  AND U18214 ( .A(p_input[1804]), .B(p_input[11804]), .Z(n9107) );
  AND U18215 ( .A(n9108), .B(p_input[21803]), .Z(o[1803]) );
  AND U18216 ( .A(p_input[1803]), .B(p_input[11803]), .Z(n9108) );
  AND U18217 ( .A(n9109), .B(p_input[21802]), .Z(o[1802]) );
  AND U18218 ( .A(p_input[1802]), .B(p_input[11802]), .Z(n9109) );
  AND U18219 ( .A(n9110), .B(p_input[21801]), .Z(o[1801]) );
  AND U18220 ( .A(p_input[1801]), .B(p_input[11801]), .Z(n9110) );
  AND U18221 ( .A(n9111), .B(p_input[21800]), .Z(o[1800]) );
  AND U18222 ( .A(p_input[1800]), .B(p_input[11800]), .Z(n9111) );
  AND U18223 ( .A(n9112), .B(p_input[20017]), .Z(o[17]) );
  AND U18224 ( .A(p_input[17]), .B(p_input[10017]), .Z(n9112) );
  AND U18225 ( .A(n9113), .B(p_input[20179]), .Z(o[179]) );
  AND U18226 ( .A(p_input[179]), .B(p_input[10179]), .Z(n9113) );
  AND U18227 ( .A(n9114), .B(p_input[21799]), .Z(o[1799]) );
  AND U18228 ( .A(p_input[1799]), .B(p_input[11799]), .Z(n9114) );
  AND U18229 ( .A(n9115), .B(p_input[21798]), .Z(o[1798]) );
  AND U18230 ( .A(p_input[1798]), .B(p_input[11798]), .Z(n9115) );
  AND U18231 ( .A(n9116), .B(p_input[21797]), .Z(o[1797]) );
  AND U18232 ( .A(p_input[1797]), .B(p_input[11797]), .Z(n9116) );
  AND U18233 ( .A(n9117), .B(p_input[21796]), .Z(o[1796]) );
  AND U18234 ( .A(p_input[1796]), .B(p_input[11796]), .Z(n9117) );
  AND U18235 ( .A(n9118), .B(p_input[21795]), .Z(o[1795]) );
  AND U18236 ( .A(p_input[1795]), .B(p_input[11795]), .Z(n9118) );
  AND U18237 ( .A(n9119), .B(p_input[21794]), .Z(o[1794]) );
  AND U18238 ( .A(p_input[1794]), .B(p_input[11794]), .Z(n9119) );
  AND U18239 ( .A(n9120), .B(p_input[21793]), .Z(o[1793]) );
  AND U18240 ( .A(p_input[1793]), .B(p_input[11793]), .Z(n9120) );
  AND U18241 ( .A(n9121), .B(p_input[21792]), .Z(o[1792]) );
  AND U18242 ( .A(p_input[1792]), .B(p_input[11792]), .Z(n9121) );
  AND U18243 ( .A(n9122), .B(p_input[21791]), .Z(o[1791]) );
  AND U18244 ( .A(p_input[1791]), .B(p_input[11791]), .Z(n9122) );
  AND U18245 ( .A(n9123), .B(p_input[21790]), .Z(o[1790]) );
  AND U18246 ( .A(p_input[1790]), .B(p_input[11790]), .Z(n9123) );
  AND U18247 ( .A(n9124), .B(p_input[20178]), .Z(o[178]) );
  AND U18248 ( .A(p_input[178]), .B(p_input[10178]), .Z(n9124) );
  AND U18249 ( .A(n9125), .B(p_input[21789]), .Z(o[1789]) );
  AND U18250 ( .A(p_input[1789]), .B(p_input[11789]), .Z(n9125) );
  AND U18251 ( .A(n9126), .B(p_input[21788]), .Z(o[1788]) );
  AND U18252 ( .A(p_input[1788]), .B(p_input[11788]), .Z(n9126) );
  AND U18253 ( .A(n9127), .B(p_input[21787]), .Z(o[1787]) );
  AND U18254 ( .A(p_input[1787]), .B(p_input[11787]), .Z(n9127) );
  AND U18255 ( .A(n9128), .B(p_input[21786]), .Z(o[1786]) );
  AND U18256 ( .A(p_input[1786]), .B(p_input[11786]), .Z(n9128) );
  AND U18257 ( .A(n9129), .B(p_input[21785]), .Z(o[1785]) );
  AND U18258 ( .A(p_input[1785]), .B(p_input[11785]), .Z(n9129) );
  AND U18259 ( .A(n9130), .B(p_input[21784]), .Z(o[1784]) );
  AND U18260 ( .A(p_input[1784]), .B(p_input[11784]), .Z(n9130) );
  AND U18261 ( .A(n9131), .B(p_input[21783]), .Z(o[1783]) );
  AND U18262 ( .A(p_input[1783]), .B(p_input[11783]), .Z(n9131) );
  AND U18263 ( .A(n9132), .B(p_input[21782]), .Z(o[1782]) );
  AND U18264 ( .A(p_input[1782]), .B(p_input[11782]), .Z(n9132) );
  AND U18265 ( .A(n9133), .B(p_input[21781]), .Z(o[1781]) );
  AND U18266 ( .A(p_input[1781]), .B(p_input[11781]), .Z(n9133) );
  AND U18267 ( .A(n9134), .B(p_input[21780]), .Z(o[1780]) );
  AND U18268 ( .A(p_input[1780]), .B(p_input[11780]), .Z(n9134) );
  AND U18269 ( .A(n9135), .B(p_input[20177]), .Z(o[177]) );
  AND U18270 ( .A(p_input[177]), .B(p_input[10177]), .Z(n9135) );
  AND U18271 ( .A(n9136), .B(p_input[21779]), .Z(o[1779]) );
  AND U18272 ( .A(p_input[1779]), .B(p_input[11779]), .Z(n9136) );
  AND U18273 ( .A(n9137), .B(p_input[21778]), .Z(o[1778]) );
  AND U18274 ( .A(p_input[1778]), .B(p_input[11778]), .Z(n9137) );
  AND U18275 ( .A(n9138), .B(p_input[21777]), .Z(o[1777]) );
  AND U18276 ( .A(p_input[1777]), .B(p_input[11777]), .Z(n9138) );
  AND U18277 ( .A(n9139), .B(p_input[21776]), .Z(o[1776]) );
  AND U18278 ( .A(p_input[1776]), .B(p_input[11776]), .Z(n9139) );
  AND U18279 ( .A(n9140), .B(p_input[21775]), .Z(o[1775]) );
  AND U18280 ( .A(p_input[1775]), .B(p_input[11775]), .Z(n9140) );
  AND U18281 ( .A(n9141), .B(p_input[21774]), .Z(o[1774]) );
  AND U18282 ( .A(p_input[1774]), .B(p_input[11774]), .Z(n9141) );
  AND U18283 ( .A(n9142), .B(p_input[21773]), .Z(o[1773]) );
  AND U18284 ( .A(p_input[1773]), .B(p_input[11773]), .Z(n9142) );
  AND U18285 ( .A(n9143), .B(p_input[21772]), .Z(o[1772]) );
  AND U18286 ( .A(p_input[1772]), .B(p_input[11772]), .Z(n9143) );
  AND U18287 ( .A(n9144), .B(p_input[21771]), .Z(o[1771]) );
  AND U18288 ( .A(p_input[1771]), .B(p_input[11771]), .Z(n9144) );
  AND U18289 ( .A(n9145), .B(p_input[21770]), .Z(o[1770]) );
  AND U18290 ( .A(p_input[1770]), .B(p_input[11770]), .Z(n9145) );
  AND U18291 ( .A(n9146), .B(p_input[20176]), .Z(o[176]) );
  AND U18292 ( .A(p_input[176]), .B(p_input[10176]), .Z(n9146) );
  AND U18293 ( .A(n9147), .B(p_input[21769]), .Z(o[1769]) );
  AND U18294 ( .A(p_input[1769]), .B(p_input[11769]), .Z(n9147) );
  AND U18295 ( .A(n9148), .B(p_input[21768]), .Z(o[1768]) );
  AND U18296 ( .A(p_input[1768]), .B(p_input[11768]), .Z(n9148) );
  AND U18297 ( .A(n9149), .B(p_input[21767]), .Z(o[1767]) );
  AND U18298 ( .A(p_input[1767]), .B(p_input[11767]), .Z(n9149) );
  AND U18299 ( .A(n9150), .B(p_input[21766]), .Z(o[1766]) );
  AND U18300 ( .A(p_input[1766]), .B(p_input[11766]), .Z(n9150) );
  AND U18301 ( .A(n9151), .B(p_input[21765]), .Z(o[1765]) );
  AND U18302 ( .A(p_input[1765]), .B(p_input[11765]), .Z(n9151) );
  AND U18303 ( .A(n9152), .B(p_input[21764]), .Z(o[1764]) );
  AND U18304 ( .A(p_input[1764]), .B(p_input[11764]), .Z(n9152) );
  AND U18305 ( .A(n9153), .B(p_input[21763]), .Z(o[1763]) );
  AND U18306 ( .A(p_input[1763]), .B(p_input[11763]), .Z(n9153) );
  AND U18307 ( .A(n9154), .B(p_input[21762]), .Z(o[1762]) );
  AND U18308 ( .A(p_input[1762]), .B(p_input[11762]), .Z(n9154) );
  AND U18309 ( .A(n9155), .B(p_input[21761]), .Z(o[1761]) );
  AND U18310 ( .A(p_input[1761]), .B(p_input[11761]), .Z(n9155) );
  AND U18311 ( .A(n9156), .B(p_input[21760]), .Z(o[1760]) );
  AND U18312 ( .A(p_input[1760]), .B(p_input[11760]), .Z(n9156) );
  AND U18313 ( .A(n9157), .B(p_input[20175]), .Z(o[175]) );
  AND U18314 ( .A(p_input[175]), .B(p_input[10175]), .Z(n9157) );
  AND U18315 ( .A(n9158), .B(p_input[21759]), .Z(o[1759]) );
  AND U18316 ( .A(p_input[1759]), .B(p_input[11759]), .Z(n9158) );
  AND U18317 ( .A(n9159), .B(p_input[21758]), .Z(o[1758]) );
  AND U18318 ( .A(p_input[1758]), .B(p_input[11758]), .Z(n9159) );
  AND U18319 ( .A(n9160), .B(p_input[21757]), .Z(o[1757]) );
  AND U18320 ( .A(p_input[1757]), .B(p_input[11757]), .Z(n9160) );
  AND U18321 ( .A(n9161), .B(p_input[21756]), .Z(o[1756]) );
  AND U18322 ( .A(p_input[1756]), .B(p_input[11756]), .Z(n9161) );
  AND U18323 ( .A(n9162), .B(p_input[21755]), .Z(o[1755]) );
  AND U18324 ( .A(p_input[1755]), .B(p_input[11755]), .Z(n9162) );
  AND U18325 ( .A(n9163), .B(p_input[21754]), .Z(o[1754]) );
  AND U18326 ( .A(p_input[1754]), .B(p_input[11754]), .Z(n9163) );
  AND U18327 ( .A(n9164), .B(p_input[21753]), .Z(o[1753]) );
  AND U18328 ( .A(p_input[1753]), .B(p_input[11753]), .Z(n9164) );
  AND U18329 ( .A(n9165), .B(p_input[21752]), .Z(o[1752]) );
  AND U18330 ( .A(p_input[1752]), .B(p_input[11752]), .Z(n9165) );
  AND U18331 ( .A(n9166), .B(p_input[21751]), .Z(o[1751]) );
  AND U18332 ( .A(p_input[1751]), .B(p_input[11751]), .Z(n9166) );
  AND U18333 ( .A(n9167), .B(p_input[21750]), .Z(o[1750]) );
  AND U18334 ( .A(p_input[1750]), .B(p_input[11750]), .Z(n9167) );
  AND U18335 ( .A(n9168), .B(p_input[20174]), .Z(o[174]) );
  AND U18336 ( .A(p_input[174]), .B(p_input[10174]), .Z(n9168) );
  AND U18337 ( .A(n9169), .B(p_input[21749]), .Z(o[1749]) );
  AND U18338 ( .A(p_input[1749]), .B(p_input[11749]), .Z(n9169) );
  AND U18339 ( .A(n9170), .B(p_input[21748]), .Z(o[1748]) );
  AND U18340 ( .A(p_input[1748]), .B(p_input[11748]), .Z(n9170) );
  AND U18341 ( .A(n9171), .B(p_input[21747]), .Z(o[1747]) );
  AND U18342 ( .A(p_input[1747]), .B(p_input[11747]), .Z(n9171) );
  AND U18343 ( .A(n9172), .B(p_input[21746]), .Z(o[1746]) );
  AND U18344 ( .A(p_input[1746]), .B(p_input[11746]), .Z(n9172) );
  AND U18345 ( .A(n9173), .B(p_input[21745]), .Z(o[1745]) );
  AND U18346 ( .A(p_input[1745]), .B(p_input[11745]), .Z(n9173) );
  AND U18347 ( .A(n9174), .B(p_input[21744]), .Z(o[1744]) );
  AND U18348 ( .A(p_input[1744]), .B(p_input[11744]), .Z(n9174) );
  AND U18349 ( .A(n9175), .B(p_input[21743]), .Z(o[1743]) );
  AND U18350 ( .A(p_input[1743]), .B(p_input[11743]), .Z(n9175) );
  AND U18351 ( .A(n9176), .B(p_input[21742]), .Z(o[1742]) );
  AND U18352 ( .A(p_input[1742]), .B(p_input[11742]), .Z(n9176) );
  AND U18353 ( .A(n9177), .B(p_input[21741]), .Z(o[1741]) );
  AND U18354 ( .A(p_input[1741]), .B(p_input[11741]), .Z(n9177) );
  AND U18355 ( .A(n9178), .B(p_input[21740]), .Z(o[1740]) );
  AND U18356 ( .A(p_input[1740]), .B(p_input[11740]), .Z(n9178) );
  AND U18357 ( .A(n9179), .B(p_input[20173]), .Z(o[173]) );
  AND U18358 ( .A(p_input[173]), .B(p_input[10173]), .Z(n9179) );
  AND U18359 ( .A(n9180), .B(p_input[21739]), .Z(o[1739]) );
  AND U18360 ( .A(p_input[1739]), .B(p_input[11739]), .Z(n9180) );
  AND U18361 ( .A(n9181), .B(p_input[21738]), .Z(o[1738]) );
  AND U18362 ( .A(p_input[1738]), .B(p_input[11738]), .Z(n9181) );
  AND U18363 ( .A(n9182), .B(p_input[21737]), .Z(o[1737]) );
  AND U18364 ( .A(p_input[1737]), .B(p_input[11737]), .Z(n9182) );
  AND U18365 ( .A(n9183), .B(p_input[21736]), .Z(o[1736]) );
  AND U18366 ( .A(p_input[1736]), .B(p_input[11736]), .Z(n9183) );
  AND U18367 ( .A(n9184), .B(p_input[21735]), .Z(o[1735]) );
  AND U18368 ( .A(p_input[1735]), .B(p_input[11735]), .Z(n9184) );
  AND U18369 ( .A(n9185), .B(p_input[21734]), .Z(o[1734]) );
  AND U18370 ( .A(p_input[1734]), .B(p_input[11734]), .Z(n9185) );
  AND U18371 ( .A(n9186), .B(p_input[21733]), .Z(o[1733]) );
  AND U18372 ( .A(p_input[1733]), .B(p_input[11733]), .Z(n9186) );
  AND U18373 ( .A(n9187), .B(p_input[21732]), .Z(o[1732]) );
  AND U18374 ( .A(p_input[1732]), .B(p_input[11732]), .Z(n9187) );
  AND U18375 ( .A(n9188), .B(p_input[21731]), .Z(o[1731]) );
  AND U18376 ( .A(p_input[1731]), .B(p_input[11731]), .Z(n9188) );
  AND U18377 ( .A(n9189), .B(p_input[21730]), .Z(o[1730]) );
  AND U18378 ( .A(p_input[1730]), .B(p_input[11730]), .Z(n9189) );
  AND U18379 ( .A(n9190), .B(p_input[20172]), .Z(o[172]) );
  AND U18380 ( .A(p_input[172]), .B(p_input[10172]), .Z(n9190) );
  AND U18381 ( .A(n9191), .B(p_input[21729]), .Z(o[1729]) );
  AND U18382 ( .A(p_input[1729]), .B(p_input[11729]), .Z(n9191) );
  AND U18383 ( .A(n9192), .B(p_input[21728]), .Z(o[1728]) );
  AND U18384 ( .A(p_input[1728]), .B(p_input[11728]), .Z(n9192) );
  AND U18385 ( .A(n9193), .B(p_input[21727]), .Z(o[1727]) );
  AND U18386 ( .A(p_input[1727]), .B(p_input[11727]), .Z(n9193) );
  AND U18387 ( .A(n9194), .B(p_input[21726]), .Z(o[1726]) );
  AND U18388 ( .A(p_input[1726]), .B(p_input[11726]), .Z(n9194) );
  AND U18389 ( .A(n9195), .B(p_input[21725]), .Z(o[1725]) );
  AND U18390 ( .A(p_input[1725]), .B(p_input[11725]), .Z(n9195) );
  AND U18391 ( .A(n9196), .B(p_input[21724]), .Z(o[1724]) );
  AND U18392 ( .A(p_input[1724]), .B(p_input[11724]), .Z(n9196) );
  AND U18393 ( .A(n9197), .B(p_input[21723]), .Z(o[1723]) );
  AND U18394 ( .A(p_input[1723]), .B(p_input[11723]), .Z(n9197) );
  AND U18395 ( .A(n9198), .B(p_input[21722]), .Z(o[1722]) );
  AND U18396 ( .A(p_input[1722]), .B(p_input[11722]), .Z(n9198) );
  AND U18397 ( .A(n9199), .B(p_input[21721]), .Z(o[1721]) );
  AND U18398 ( .A(p_input[1721]), .B(p_input[11721]), .Z(n9199) );
  AND U18399 ( .A(n9200), .B(p_input[21720]), .Z(o[1720]) );
  AND U18400 ( .A(p_input[1720]), .B(p_input[11720]), .Z(n9200) );
  AND U18401 ( .A(n9201), .B(p_input[20171]), .Z(o[171]) );
  AND U18402 ( .A(p_input[171]), .B(p_input[10171]), .Z(n9201) );
  AND U18403 ( .A(n9202), .B(p_input[21719]), .Z(o[1719]) );
  AND U18404 ( .A(p_input[1719]), .B(p_input[11719]), .Z(n9202) );
  AND U18405 ( .A(n9203), .B(p_input[21718]), .Z(o[1718]) );
  AND U18406 ( .A(p_input[1718]), .B(p_input[11718]), .Z(n9203) );
  AND U18407 ( .A(n9204), .B(p_input[21717]), .Z(o[1717]) );
  AND U18408 ( .A(p_input[1717]), .B(p_input[11717]), .Z(n9204) );
  AND U18409 ( .A(n9205), .B(p_input[21716]), .Z(o[1716]) );
  AND U18410 ( .A(p_input[1716]), .B(p_input[11716]), .Z(n9205) );
  AND U18411 ( .A(n9206), .B(p_input[21715]), .Z(o[1715]) );
  AND U18412 ( .A(p_input[1715]), .B(p_input[11715]), .Z(n9206) );
  AND U18413 ( .A(n9207), .B(p_input[21714]), .Z(o[1714]) );
  AND U18414 ( .A(p_input[1714]), .B(p_input[11714]), .Z(n9207) );
  AND U18415 ( .A(n9208), .B(p_input[21713]), .Z(o[1713]) );
  AND U18416 ( .A(p_input[1713]), .B(p_input[11713]), .Z(n9208) );
  AND U18417 ( .A(n9209), .B(p_input[21712]), .Z(o[1712]) );
  AND U18418 ( .A(p_input[1712]), .B(p_input[11712]), .Z(n9209) );
  AND U18419 ( .A(n9210), .B(p_input[21711]), .Z(o[1711]) );
  AND U18420 ( .A(p_input[1711]), .B(p_input[11711]), .Z(n9210) );
  AND U18421 ( .A(n9211), .B(p_input[21710]), .Z(o[1710]) );
  AND U18422 ( .A(p_input[1710]), .B(p_input[11710]), .Z(n9211) );
  AND U18423 ( .A(n9212), .B(p_input[20170]), .Z(o[170]) );
  AND U18424 ( .A(p_input[170]), .B(p_input[10170]), .Z(n9212) );
  AND U18425 ( .A(n9213), .B(p_input[21709]), .Z(o[1709]) );
  AND U18426 ( .A(p_input[1709]), .B(p_input[11709]), .Z(n9213) );
  AND U18427 ( .A(n9214), .B(p_input[21708]), .Z(o[1708]) );
  AND U18428 ( .A(p_input[1708]), .B(p_input[11708]), .Z(n9214) );
  AND U18429 ( .A(n9215), .B(p_input[21707]), .Z(o[1707]) );
  AND U18430 ( .A(p_input[1707]), .B(p_input[11707]), .Z(n9215) );
  AND U18431 ( .A(n9216), .B(p_input[21706]), .Z(o[1706]) );
  AND U18432 ( .A(p_input[1706]), .B(p_input[11706]), .Z(n9216) );
  AND U18433 ( .A(n9217), .B(p_input[21705]), .Z(o[1705]) );
  AND U18434 ( .A(p_input[1705]), .B(p_input[11705]), .Z(n9217) );
  AND U18435 ( .A(n9218), .B(p_input[21704]), .Z(o[1704]) );
  AND U18436 ( .A(p_input[1704]), .B(p_input[11704]), .Z(n9218) );
  AND U18437 ( .A(n9219), .B(p_input[21703]), .Z(o[1703]) );
  AND U18438 ( .A(p_input[1703]), .B(p_input[11703]), .Z(n9219) );
  AND U18439 ( .A(n9220), .B(p_input[21702]), .Z(o[1702]) );
  AND U18440 ( .A(p_input[1702]), .B(p_input[11702]), .Z(n9220) );
  AND U18441 ( .A(n9221), .B(p_input[21701]), .Z(o[1701]) );
  AND U18442 ( .A(p_input[1701]), .B(p_input[11701]), .Z(n9221) );
  AND U18443 ( .A(n9222), .B(p_input[21700]), .Z(o[1700]) );
  AND U18444 ( .A(p_input[1700]), .B(p_input[11700]), .Z(n9222) );
  AND U18445 ( .A(n9223), .B(p_input[20016]), .Z(o[16]) );
  AND U18446 ( .A(p_input[16]), .B(p_input[10016]), .Z(n9223) );
  AND U18447 ( .A(n9224), .B(p_input[20169]), .Z(o[169]) );
  AND U18448 ( .A(p_input[169]), .B(p_input[10169]), .Z(n9224) );
  AND U18449 ( .A(n9225), .B(p_input[21699]), .Z(o[1699]) );
  AND U18450 ( .A(p_input[1699]), .B(p_input[11699]), .Z(n9225) );
  AND U18451 ( .A(n9226), .B(p_input[21698]), .Z(o[1698]) );
  AND U18452 ( .A(p_input[1698]), .B(p_input[11698]), .Z(n9226) );
  AND U18453 ( .A(n9227), .B(p_input[21697]), .Z(o[1697]) );
  AND U18454 ( .A(p_input[1697]), .B(p_input[11697]), .Z(n9227) );
  AND U18455 ( .A(n9228), .B(p_input[21696]), .Z(o[1696]) );
  AND U18456 ( .A(p_input[1696]), .B(p_input[11696]), .Z(n9228) );
  AND U18457 ( .A(n9229), .B(p_input[21695]), .Z(o[1695]) );
  AND U18458 ( .A(p_input[1695]), .B(p_input[11695]), .Z(n9229) );
  AND U18459 ( .A(n9230), .B(p_input[21694]), .Z(o[1694]) );
  AND U18460 ( .A(p_input[1694]), .B(p_input[11694]), .Z(n9230) );
  AND U18461 ( .A(n9231), .B(p_input[21693]), .Z(o[1693]) );
  AND U18462 ( .A(p_input[1693]), .B(p_input[11693]), .Z(n9231) );
  AND U18463 ( .A(n9232), .B(p_input[21692]), .Z(o[1692]) );
  AND U18464 ( .A(p_input[1692]), .B(p_input[11692]), .Z(n9232) );
  AND U18465 ( .A(n9233), .B(p_input[21691]), .Z(o[1691]) );
  AND U18466 ( .A(p_input[1691]), .B(p_input[11691]), .Z(n9233) );
  AND U18467 ( .A(n9234), .B(p_input[21690]), .Z(o[1690]) );
  AND U18468 ( .A(p_input[1690]), .B(p_input[11690]), .Z(n9234) );
  AND U18469 ( .A(n9235), .B(p_input[20168]), .Z(o[168]) );
  AND U18470 ( .A(p_input[168]), .B(p_input[10168]), .Z(n9235) );
  AND U18471 ( .A(n9236), .B(p_input[21689]), .Z(o[1689]) );
  AND U18472 ( .A(p_input[1689]), .B(p_input[11689]), .Z(n9236) );
  AND U18473 ( .A(n9237), .B(p_input[21688]), .Z(o[1688]) );
  AND U18474 ( .A(p_input[1688]), .B(p_input[11688]), .Z(n9237) );
  AND U18475 ( .A(n9238), .B(p_input[21687]), .Z(o[1687]) );
  AND U18476 ( .A(p_input[1687]), .B(p_input[11687]), .Z(n9238) );
  AND U18477 ( .A(n9239), .B(p_input[21686]), .Z(o[1686]) );
  AND U18478 ( .A(p_input[1686]), .B(p_input[11686]), .Z(n9239) );
  AND U18479 ( .A(n9240), .B(p_input[21685]), .Z(o[1685]) );
  AND U18480 ( .A(p_input[1685]), .B(p_input[11685]), .Z(n9240) );
  AND U18481 ( .A(n9241), .B(p_input[21684]), .Z(o[1684]) );
  AND U18482 ( .A(p_input[1684]), .B(p_input[11684]), .Z(n9241) );
  AND U18483 ( .A(n9242), .B(p_input[21683]), .Z(o[1683]) );
  AND U18484 ( .A(p_input[1683]), .B(p_input[11683]), .Z(n9242) );
  AND U18485 ( .A(n9243), .B(p_input[21682]), .Z(o[1682]) );
  AND U18486 ( .A(p_input[1682]), .B(p_input[11682]), .Z(n9243) );
  AND U18487 ( .A(n9244), .B(p_input[21681]), .Z(o[1681]) );
  AND U18488 ( .A(p_input[1681]), .B(p_input[11681]), .Z(n9244) );
  AND U18489 ( .A(n9245), .B(p_input[21680]), .Z(o[1680]) );
  AND U18490 ( .A(p_input[1680]), .B(p_input[11680]), .Z(n9245) );
  AND U18491 ( .A(n9246), .B(p_input[20167]), .Z(o[167]) );
  AND U18492 ( .A(p_input[167]), .B(p_input[10167]), .Z(n9246) );
  AND U18493 ( .A(n9247), .B(p_input[21679]), .Z(o[1679]) );
  AND U18494 ( .A(p_input[1679]), .B(p_input[11679]), .Z(n9247) );
  AND U18495 ( .A(n9248), .B(p_input[21678]), .Z(o[1678]) );
  AND U18496 ( .A(p_input[1678]), .B(p_input[11678]), .Z(n9248) );
  AND U18497 ( .A(n9249), .B(p_input[21677]), .Z(o[1677]) );
  AND U18498 ( .A(p_input[1677]), .B(p_input[11677]), .Z(n9249) );
  AND U18499 ( .A(n9250), .B(p_input[21676]), .Z(o[1676]) );
  AND U18500 ( .A(p_input[1676]), .B(p_input[11676]), .Z(n9250) );
  AND U18501 ( .A(n9251), .B(p_input[21675]), .Z(o[1675]) );
  AND U18502 ( .A(p_input[1675]), .B(p_input[11675]), .Z(n9251) );
  AND U18503 ( .A(n9252), .B(p_input[21674]), .Z(o[1674]) );
  AND U18504 ( .A(p_input[1674]), .B(p_input[11674]), .Z(n9252) );
  AND U18505 ( .A(n9253), .B(p_input[21673]), .Z(o[1673]) );
  AND U18506 ( .A(p_input[1673]), .B(p_input[11673]), .Z(n9253) );
  AND U18507 ( .A(n9254), .B(p_input[21672]), .Z(o[1672]) );
  AND U18508 ( .A(p_input[1672]), .B(p_input[11672]), .Z(n9254) );
  AND U18509 ( .A(n9255), .B(p_input[21671]), .Z(o[1671]) );
  AND U18510 ( .A(p_input[1671]), .B(p_input[11671]), .Z(n9255) );
  AND U18511 ( .A(n9256), .B(p_input[21670]), .Z(o[1670]) );
  AND U18512 ( .A(p_input[1670]), .B(p_input[11670]), .Z(n9256) );
  AND U18513 ( .A(n9257), .B(p_input[20166]), .Z(o[166]) );
  AND U18514 ( .A(p_input[166]), .B(p_input[10166]), .Z(n9257) );
  AND U18515 ( .A(n9258), .B(p_input[21669]), .Z(o[1669]) );
  AND U18516 ( .A(p_input[1669]), .B(p_input[11669]), .Z(n9258) );
  AND U18517 ( .A(n9259), .B(p_input[21668]), .Z(o[1668]) );
  AND U18518 ( .A(p_input[1668]), .B(p_input[11668]), .Z(n9259) );
  AND U18519 ( .A(n9260), .B(p_input[21667]), .Z(o[1667]) );
  AND U18520 ( .A(p_input[1667]), .B(p_input[11667]), .Z(n9260) );
  AND U18521 ( .A(n9261), .B(p_input[21666]), .Z(o[1666]) );
  AND U18522 ( .A(p_input[1666]), .B(p_input[11666]), .Z(n9261) );
  AND U18523 ( .A(n9262), .B(p_input[21665]), .Z(o[1665]) );
  AND U18524 ( .A(p_input[1665]), .B(p_input[11665]), .Z(n9262) );
  AND U18525 ( .A(n9263), .B(p_input[21664]), .Z(o[1664]) );
  AND U18526 ( .A(p_input[1664]), .B(p_input[11664]), .Z(n9263) );
  AND U18527 ( .A(n9264), .B(p_input[21663]), .Z(o[1663]) );
  AND U18528 ( .A(p_input[1663]), .B(p_input[11663]), .Z(n9264) );
  AND U18529 ( .A(n9265), .B(p_input[21662]), .Z(o[1662]) );
  AND U18530 ( .A(p_input[1662]), .B(p_input[11662]), .Z(n9265) );
  AND U18531 ( .A(n9266), .B(p_input[21661]), .Z(o[1661]) );
  AND U18532 ( .A(p_input[1661]), .B(p_input[11661]), .Z(n9266) );
  AND U18533 ( .A(n9267), .B(p_input[21660]), .Z(o[1660]) );
  AND U18534 ( .A(p_input[1660]), .B(p_input[11660]), .Z(n9267) );
  AND U18535 ( .A(n9268), .B(p_input[20165]), .Z(o[165]) );
  AND U18536 ( .A(p_input[165]), .B(p_input[10165]), .Z(n9268) );
  AND U18537 ( .A(n9269), .B(p_input[21659]), .Z(o[1659]) );
  AND U18538 ( .A(p_input[1659]), .B(p_input[11659]), .Z(n9269) );
  AND U18539 ( .A(n9270), .B(p_input[21658]), .Z(o[1658]) );
  AND U18540 ( .A(p_input[1658]), .B(p_input[11658]), .Z(n9270) );
  AND U18541 ( .A(n9271), .B(p_input[21657]), .Z(o[1657]) );
  AND U18542 ( .A(p_input[1657]), .B(p_input[11657]), .Z(n9271) );
  AND U18543 ( .A(n9272), .B(p_input[21656]), .Z(o[1656]) );
  AND U18544 ( .A(p_input[1656]), .B(p_input[11656]), .Z(n9272) );
  AND U18545 ( .A(n9273), .B(p_input[21655]), .Z(o[1655]) );
  AND U18546 ( .A(p_input[1655]), .B(p_input[11655]), .Z(n9273) );
  AND U18547 ( .A(n9274), .B(p_input[21654]), .Z(o[1654]) );
  AND U18548 ( .A(p_input[1654]), .B(p_input[11654]), .Z(n9274) );
  AND U18549 ( .A(n9275), .B(p_input[21653]), .Z(o[1653]) );
  AND U18550 ( .A(p_input[1653]), .B(p_input[11653]), .Z(n9275) );
  AND U18551 ( .A(n9276), .B(p_input[21652]), .Z(o[1652]) );
  AND U18552 ( .A(p_input[1652]), .B(p_input[11652]), .Z(n9276) );
  AND U18553 ( .A(n9277), .B(p_input[21651]), .Z(o[1651]) );
  AND U18554 ( .A(p_input[1651]), .B(p_input[11651]), .Z(n9277) );
  AND U18555 ( .A(n9278), .B(p_input[21650]), .Z(o[1650]) );
  AND U18556 ( .A(p_input[1650]), .B(p_input[11650]), .Z(n9278) );
  AND U18557 ( .A(n9279), .B(p_input[20164]), .Z(o[164]) );
  AND U18558 ( .A(p_input[164]), .B(p_input[10164]), .Z(n9279) );
  AND U18559 ( .A(n9280), .B(p_input[21649]), .Z(o[1649]) );
  AND U18560 ( .A(p_input[1649]), .B(p_input[11649]), .Z(n9280) );
  AND U18561 ( .A(n9281), .B(p_input[21648]), .Z(o[1648]) );
  AND U18562 ( .A(p_input[1648]), .B(p_input[11648]), .Z(n9281) );
  AND U18563 ( .A(n9282), .B(p_input[21647]), .Z(o[1647]) );
  AND U18564 ( .A(p_input[1647]), .B(p_input[11647]), .Z(n9282) );
  AND U18565 ( .A(n9283), .B(p_input[21646]), .Z(o[1646]) );
  AND U18566 ( .A(p_input[1646]), .B(p_input[11646]), .Z(n9283) );
  AND U18567 ( .A(n9284), .B(p_input[21645]), .Z(o[1645]) );
  AND U18568 ( .A(p_input[1645]), .B(p_input[11645]), .Z(n9284) );
  AND U18569 ( .A(n9285), .B(p_input[21644]), .Z(o[1644]) );
  AND U18570 ( .A(p_input[1644]), .B(p_input[11644]), .Z(n9285) );
  AND U18571 ( .A(n9286), .B(p_input[21643]), .Z(o[1643]) );
  AND U18572 ( .A(p_input[1643]), .B(p_input[11643]), .Z(n9286) );
  AND U18573 ( .A(n9287), .B(p_input[21642]), .Z(o[1642]) );
  AND U18574 ( .A(p_input[1642]), .B(p_input[11642]), .Z(n9287) );
  AND U18575 ( .A(n9288), .B(p_input[21641]), .Z(o[1641]) );
  AND U18576 ( .A(p_input[1641]), .B(p_input[11641]), .Z(n9288) );
  AND U18577 ( .A(n9289), .B(p_input[21640]), .Z(o[1640]) );
  AND U18578 ( .A(p_input[1640]), .B(p_input[11640]), .Z(n9289) );
  AND U18579 ( .A(n9290), .B(p_input[20163]), .Z(o[163]) );
  AND U18580 ( .A(p_input[163]), .B(p_input[10163]), .Z(n9290) );
  AND U18581 ( .A(n9291), .B(p_input[21639]), .Z(o[1639]) );
  AND U18582 ( .A(p_input[1639]), .B(p_input[11639]), .Z(n9291) );
  AND U18583 ( .A(n9292), .B(p_input[21638]), .Z(o[1638]) );
  AND U18584 ( .A(p_input[1638]), .B(p_input[11638]), .Z(n9292) );
  AND U18585 ( .A(n9293), .B(p_input[21637]), .Z(o[1637]) );
  AND U18586 ( .A(p_input[1637]), .B(p_input[11637]), .Z(n9293) );
  AND U18587 ( .A(n9294), .B(p_input[21636]), .Z(o[1636]) );
  AND U18588 ( .A(p_input[1636]), .B(p_input[11636]), .Z(n9294) );
  AND U18589 ( .A(n9295), .B(p_input[21635]), .Z(o[1635]) );
  AND U18590 ( .A(p_input[1635]), .B(p_input[11635]), .Z(n9295) );
  AND U18591 ( .A(n9296), .B(p_input[21634]), .Z(o[1634]) );
  AND U18592 ( .A(p_input[1634]), .B(p_input[11634]), .Z(n9296) );
  AND U18593 ( .A(n9297), .B(p_input[21633]), .Z(o[1633]) );
  AND U18594 ( .A(p_input[1633]), .B(p_input[11633]), .Z(n9297) );
  AND U18595 ( .A(n9298), .B(p_input[21632]), .Z(o[1632]) );
  AND U18596 ( .A(p_input[1632]), .B(p_input[11632]), .Z(n9298) );
  AND U18597 ( .A(n9299), .B(p_input[21631]), .Z(o[1631]) );
  AND U18598 ( .A(p_input[1631]), .B(p_input[11631]), .Z(n9299) );
  AND U18599 ( .A(n9300), .B(p_input[21630]), .Z(o[1630]) );
  AND U18600 ( .A(p_input[1630]), .B(p_input[11630]), .Z(n9300) );
  AND U18601 ( .A(n9301), .B(p_input[20162]), .Z(o[162]) );
  AND U18602 ( .A(p_input[162]), .B(p_input[10162]), .Z(n9301) );
  AND U18603 ( .A(n9302), .B(p_input[21629]), .Z(o[1629]) );
  AND U18604 ( .A(p_input[1629]), .B(p_input[11629]), .Z(n9302) );
  AND U18605 ( .A(n9303), .B(p_input[21628]), .Z(o[1628]) );
  AND U18606 ( .A(p_input[1628]), .B(p_input[11628]), .Z(n9303) );
  AND U18607 ( .A(n9304), .B(p_input[21627]), .Z(o[1627]) );
  AND U18608 ( .A(p_input[1627]), .B(p_input[11627]), .Z(n9304) );
  AND U18609 ( .A(n9305), .B(p_input[21626]), .Z(o[1626]) );
  AND U18610 ( .A(p_input[1626]), .B(p_input[11626]), .Z(n9305) );
  AND U18611 ( .A(n9306), .B(p_input[21625]), .Z(o[1625]) );
  AND U18612 ( .A(p_input[1625]), .B(p_input[11625]), .Z(n9306) );
  AND U18613 ( .A(n9307), .B(p_input[21624]), .Z(o[1624]) );
  AND U18614 ( .A(p_input[1624]), .B(p_input[11624]), .Z(n9307) );
  AND U18615 ( .A(n9308), .B(p_input[21623]), .Z(o[1623]) );
  AND U18616 ( .A(p_input[1623]), .B(p_input[11623]), .Z(n9308) );
  AND U18617 ( .A(n9309), .B(p_input[21622]), .Z(o[1622]) );
  AND U18618 ( .A(p_input[1622]), .B(p_input[11622]), .Z(n9309) );
  AND U18619 ( .A(n9310), .B(p_input[21621]), .Z(o[1621]) );
  AND U18620 ( .A(p_input[1621]), .B(p_input[11621]), .Z(n9310) );
  AND U18621 ( .A(n9311), .B(p_input[21620]), .Z(o[1620]) );
  AND U18622 ( .A(p_input[1620]), .B(p_input[11620]), .Z(n9311) );
  AND U18623 ( .A(n9312), .B(p_input[20161]), .Z(o[161]) );
  AND U18624 ( .A(p_input[161]), .B(p_input[10161]), .Z(n9312) );
  AND U18625 ( .A(n9313), .B(p_input[21619]), .Z(o[1619]) );
  AND U18626 ( .A(p_input[1619]), .B(p_input[11619]), .Z(n9313) );
  AND U18627 ( .A(n9314), .B(p_input[21618]), .Z(o[1618]) );
  AND U18628 ( .A(p_input[1618]), .B(p_input[11618]), .Z(n9314) );
  AND U18629 ( .A(n9315), .B(p_input[21617]), .Z(o[1617]) );
  AND U18630 ( .A(p_input[1617]), .B(p_input[11617]), .Z(n9315) );
  AND U18631 ( .A(n9316), .B(p_input[21616]), .Z(o[1616]) );
  AND U18632 ( .A(p_input[1616]), .B(p_input[11616]), .Z(n9316) );
  AND U18633 ( .A(n9317), .B(p_input[21615]), .Z(o[1615]) );
  AND U18634 ( .A(p_input[1615]), .B(p_input[11615]), .Z(n9317) );
  AND U18635 ( .A(n9318), .B(p_input[21614]), .Z(o[1614]) );
  AND U18636 ( .A(p_input[1614]), .B(p_input[11614]), .Z(n9318) );
  AND U18637 ( .A(n9319), .B(p_input[21613]), .Z(o[1613]) );
  AND U18638 ( .A(p_input[1613]), .B(p_input[11613]), .Z(n9319) );
  AND U18639 ( .A(n9320), .B(p_input[21612]), .Z(o[1612]) );
  AND U18640 ( .A(p_input[1612]), .B(p_input[11612]), .Z(n9320) );
  AND U18641 ( .A(n9321), .B(p_input[21611]), .Z(o[1611]) );
  AND U18642 ( .A(p_input[1611]), .B(p_input[11611]), .Z(n9321) );
  AND U18643 ( .A(n9322), .B(p_input[21610]), .Z(o[1610]) );
  AND U18644 ( .A(p_input[1610]), .B(p_input[11610]), .Z(n9322) );
  AND U18645 ( .A(n9323), .B(p_input[20160]), .Z(o[160]) );
  AND U18646 ( .A(p_input[160]), .B(p_input[10160]), .Z(n9323) );
  AND U18647 ( .A(n9324), .B(p_input[21609]), .Z(o[1609]) );
  AND U18648 ( .A(p_input[1609]), .B(p_input[11609]), .Z(n9324) );
  AND U18649 ( .A(n9325), .B(p_input[21608]), .Z(o[1608]) );
  AND U18650 ( .A(p_input[1608]), .B(p_input[11608]), .Z(n9325) );
  AND U18651 ( .A(n9326), .B(p_input[21607]), .Z(o[1607]) );
  AND U18652 ( .A(p_input[1607]), .B(p_input[11607]), .Z(n9326) );
  AND U18653 ( .A(n9327), .B(p_input[21606]), .Z(o[1606]) );
  AND U18654 ( .A(p_input[1606]), .B(p_input[11606]), .Z(n9327) );
  AND U18655 ( .A(n9328), .B(p_input[21605]), .Z(o[1605]) );
  AND U18656 ( .A(p_input[1605]), .B(p_input[11605]), .Z(n9328) );
  AND U18657 ( .A(n9329), .B(p_input[21604]), .Z(o[1604]) );
  AND U18658 ( .A(p_input[1604]), .B(p_input[11604]), .Z(n9329) );
  AND U18659 ( .A(n9330), .B(p_input[21603]), .Z(o[1603]) );
  AND U18660 ( .A(p_input[1603]), .B(p_input[11603]), .Z(n9330) );
  AND U18661 ( .A(n9331), .B(p_input[21602]), .Z(o[1602]) );
  AND U18662 ( .A(p_input[1602]), .B(p_input[11602]), .Z(n9331) );
  AND U18663 ( .A(n9332), .B(p_input[21601]), .Z(o[1601]) );
  AND U18664 ( .A(p_input[1601]), .B(p_input[11601]), .Z(n9332) );
  AND U18665 ( .A(n9333), .B(p_input[21600]), .Z(o[1600]) );
  AND U18666 ( .A(p_input[1600]), .B(p_input[11600]), .Z(n9333) );
  AND U18667 ( .A(n9334), .B(p_input[20015]), .Z(o[15]) );
  AND U18668 ( .A(p_input[15]), .B(p_input[10015]), .Z(n9334) );
  AND U18669 ( .A(n9335), .B(p_input[20159]), .Z(o[159]) );
  AND U18670 ( .A(p_input[159]), .B(p_input[10159]), .Z(n9335) );
  AND U18671 ( .A(n9336), .B(p_input[21599]), .Z(o[1599]) );
  AND U18672 ( .A(p_input[1599]), .B(p_input[11599]), .Z(n9336) );
  AND U18673 ( .A(n9337), .B(p_input[21598]), .Z(o[1598]) );
  AND U18674 ( .A(p_input[1598]), .B(p_input[11598]), .Z(n9337) );
  AND U18675 ( .A(n9338), .B(p_input[21597]), .Z(o[1597]) );
  AND U18676 ( .A(p_input[1597]), .B(p_input[11597]), .Z(n9338) );
  AND U18677 ( .A(n9339), .B(p_input[21596]), .Z(o[1596]) );
  AND U18678 ( .A(p_input[1596]), .B(p_input[11596]), .Z(n9339) );
  AND U18679 ( .A(n9340), .B(p_input[21595]), .Z(o[1595]) );
  AND U18680 ( .A(p_input[1595]), .B(p_input[11595]), .Z(n9340) );
  AND U18681 ( .A(n9341), .B(p_input[21594]), .Z(o[1594]) );
  AND U18682 ( .A(p_input[1594]), .B(p_input[11594]), .Z(n9341) );
  AND U18683 ( .A(n9342), .B(p_input[21593]), .Z(o[1593]) );
  AND U18684 ( .A(p_input[1593]), .B(p_input[11593]), .Z(n9342) );
  AND U18685 ( .A(n9343), .B(p_input[21592]), .Z(o[1592]) );
  AND U18686 ( .A(p_input[1592]), .B(p_input[11592]), .Z(n9343) );
  AND U18687 ( .A(n9344), .B(p_input[21591]), .Z(o[1591]) );
  AND U18688 ( .A(p_input[1591]), .B(p_input[11591]), .Z(n9344) );
  AND U18689 ( .A(n9345), .B(p_input[21590]), .Z(o[1590]) );
  AND U18690 ( .A(p_input[1590]), .B(p_input[11590]), .Z(n9345) );
  AND U18691 ( .A(n9346), .B(p_input[20158]), .Z(o[158]) );
  AND U18692 ( .A(p_input[158]), .B(p_input[10158]), .Z(n9346) );
  AND U18693 ( .A(n9347), .B(p_input[21589]), .Z(o[1589]) );
  AND U18694 ( .A(p_input[1589]), .B(p_input[11589]), .Z(n9347) );
  AND U18695 ( .A(n9348), .B(p_input[21588]), .Z(o[1588]) );
  AND U18696 ( .A(p_input[1588]), .B(p_input[11588]), .Z(n9348) );
  AND U18697 ( .A(n9349), .B(p_input[21587]), .Z(o[1587]) );
  AND U18698 ( .A(p_input[1587]), .B(p_input[11587]), .Z(n9349) );
  AND U18699 ( .A(n9350), .B(p_input[21586]), .Z(o[1586]) );
  AND U18700 ( .A(p_input[1586]), .B(p_input[11586]), .Z(n9350) );
  AND U18701 ( .A(n9351), .B(p_input[21585]), .Z(o[1585]) );
  AND U18702 ( .A(p_input[1585]), .B(p_input[11585]), .Z(n9351) );
  AND U18703 ( .A(n9352), .B(p_input[21584]), .Z(o[1584]) );
  AND U18704 ( .A(p_input[1584]), .B(p_input[11584]), .Z(n9352) );
  AND U18705 ( .A(n9353), .B(p_input[21583]), .Z(o[1583]) );
  AND U18706 ( .A(p_input[1583]), .B(p_input[11583]), .Z(n9353) );
  AND U18707 ( .A(n9354), .B(p_input[21582]), .Z(o[1582]) );
  AND U18708 ( .A(p_input[1582]), .B(p_input[11582]), .Z(n9354) );
  AND U18709 ( .A(n9355), .B(p_input[21581]), .Z(o[1581]) );
  AND U18710 ( .A(p_input[1581]), .B(p_input[11581]), .Z(n9355) );
  AND U18711 ( .A(n9356), .B(p_input[21580]), .Z(o[1580]) );
  AND U18712 ( .A(p_input[1580]), .B(p_input[11580]), .Z(n9356) );
  AND U18713 ( .A(n9357), .B(p_input[20157]), .Z(o[157]) );
  AND U18714 ( .A(p_input[157]), .B(p_input[10157]), .Z(n9357) );
  AND U18715 ( .A(n9358), .B(p_input[21579]), .Z(o[1579]) );
  AND U18716 ( .A(p_input[1579]), .B(p_input[11579]), .Z(n9358) );
  AND U18717 ( .A(n9359), .B(p_input[21578]), .Z(o[1578]) );
  AND U18718 ( .A(p_input[1578]), .B(p_input[11578]), .Z(n9359) );
  AND U18719 ( .A(n9360), .B(p_input[21577]), .Z(o[1577]) );
  AND U18720 ( .A(p_input[1577]), .B(p_input[11577]), .Z(n9360) );
  AND U18721 ( .A(n9361), .B(p_input[21576]), .Z(o[1576]) );
  AND U18722 ( .A(p_input[1576]), .B(p_input[11576]), .Z(n9361) );
  AND U18723 ( .A(n9362), .B(p_input[21575]), .Z(o[1575]) );
  AND U18724 ( .A(p_input[1575]), .B(p_input[11575]), .Z(n9362) );
  AND U18725 ( .A(n9363), .B(p_input[21574]), .Z(o[1574]) );
  AND U18726 ( .A(p_input[1574]), .B(p_input[11574]), .Z(n9363) );
  AND U18727 ( .A(n9364), .B(p_input[21573]), .Z(o[1573]) );
  AND U18728 ( .A(p_input[1573]), .B(p_input[11573]), .Z(n9364) );
  AND U18729 ( .A(n9365), .B(p_input[21572]), .Z(o[1572]) );
  AND U18730 ( .A(p_input[1572]), .B(p_input[11572]), .Z(n9365) );
  AND U18731 ( .A(n9366), .B(p_input[21571]), .Z(o[1571]) );
  AND U18732 ( .A(p_input[1571]), .B(p_input[11571]), .Z(n9366) );
  AND U18733 ( .A(n9367), .B(p_input[21570]), .Z(o[1570]) );
  AND U18734 ( .A(p_input[1570]), .B(p_input[11570]), .Z(n9367) );
  AND U18735 ( .A(n9368), .B(p_input[20156]), .Z(o[156]) );
  AND U18736 ( .A(p_input[156]), .B(p_input[10156]), .Z(n9368) );
  AND U18737 ( .A(n9369), .B(p_input[21569]), .Z(o[1569]) );
  AND U18738 ( .A(p_input[1569]), .B(p_input[11569]), .Z(n9369) );
  AND U18739 ( .A(n9370), .B(p_input[21568]), .Z(o[1568]) );
  AND U18740 ( .A(p_input[1568]), .B(p_input[11568]), .Z(n9370) );
  AND U18741 ( .A(n9371), .B(p_input[21567]), .Z(o[1567]) );
  AND U18742 ( .A(p_input[1567]), .B(p_input[11567]), .Z(n9371) );
  AND U18743 ( .A(n9372), .B(p_input[21566]), .Z(o[1566]) );
  AND U18744 ( .A(p_input[1566]), .B(p_input[11566]), .Z(n9372) );
  AND U18745 ( .A(n9373), .B(p_input[21565]), .Z(o[1565]) );
  AND U18746 ( .A(p_input[1565]), .B(p_input[11565]), .Z(n9373) );
  AND U18747 ( .A(n9374), .B(p_input[21564]), .Z(o[1564]) );
  AND U18748 ( .A(p_input[1564]), .B(p_input[11564]), .Z(n9374) );
  AND U18749 ( .A(n9375), .B(p_input[21563]), .Z(o[1563]) );
  AND U18750 ( .A(p_input[1563]), .B(p_input[11563]), .Z(n9375) );
  AND U18751 ( .A(n9376), .B(p_input[21562]), .Z(o[1562]) );
  AND U18752 ( .A(p_input[1562]), .B(p_input[11562]), .Z(n9376) );
  AND U18753 ( .A(n9377), .B(p_input[21561]), .Z(o[1561]) );
  AND U18754 ( .A(p_input[1561]), .B(p_input[11561]), .Z(n9377) );
  AND U18755 ( .A(n9378), .B(p_input[21560]), .Z(o[1560]) );
  AND U18756 ( .A(p_input[1560]), .B(p_input[11560]), .Z(n9378) );
  AND U18757 ( .A(n9379), .B(p_input[20155]), .Z(o[155]) );
  AND U18758 ( .A(p_input[155]), .B(p_input[10155]), .Z(n9379) );
  AND U18759 ( .A(n9380), .B(p_input[21559]), .Z(o[1559]) );
  AND U18760 ( .A(p_input[1559]), .B(p_input[11559]), .Z(n9380) );
  AND U18761 ( .A(n9381), .B(p_input[21558]), .Z(o[1558]) );
  AND U18762 ( .A(p_input[1558]), .B(p_input[11558]), .Z(n9381) );
  AND U18763 ( .A(n9382), .B(p_input[21557]), .Z(o[1557]) );
  AND U18764 ( .A(p_input[1557]), .B(p_input[11557]), .Z(n9382) );
  AND U18765 ( .A(n9383), .B(p_input[21556]), .Z(o[1556]) );
  AND U18766 ( .A(p_input[1556]), .B(p_input[11556]), .Z(n9383) );
  AND U18767 ( .A(n9384), .B(p_input[21555]), .Z(o[1555]) );
  AND U18768 ( .A(p_input[1555]), .B(p_input[11555]), .Z(n9384) );
  AND U18769 ( .A(n9385), .B(p_input[21554]), .Z(o[1554]) );
  AND U18770 ( .A(p_input[1554]), .B(p_input[11554]), .Z(n9385) );
  AND U18771 ( .A(n9386), .B(p_input[21553]), .Z(o[1553]) );
  AND U18772 ( .A(p_input[1553]), .B(p_input[11553]), .Z(n9386) );
  AND U18773 ( .A(n9387), .B(p_input[21552]), .Z(o[1552]) );
  AND U18774 ( .A(p_input[1552]), .B(p_input[11552]), .Z(n9387) );
  AND U18775 ( .A(n9388), .B(p_input[21551]), .Z(o[1551]) );
  AND U18776 ( .A(p_input[1551]), .B(p_input[11551]), .Z(n9388) );
  AND U18777 ( .A(n9389), .B(p_input[21550]), .Z(o[1550]) );
  AND U18778 ( .A(p_input[1550]), .B(p_input[11550]), .Z(n9389) );
  AND U18779 ( .A(n9390), .B(p_input[20154]), .Z(o[154]) );
  AND U18780 ( .A(p_input[154]), .B(p_input[10154]), .Z(n9390) );
  AND U18781 ( .A(n9391), .B(p_input[21549]), .Z(o[1549]) );
  AND U18782 ( .A(p_input[1549]), .B(p_input[11549]), .Z(n9391) );
  AND U18783 ( .A(n9392), .B(p_input[21548]), .Z(o[1548]) );
  AND U18784 ( .A(p_input[1548]), .B(p_input[11548]), .Z(n9392) );
  AND U18785 ( .A(n9393), .B(p_input[21547]), .Z(o[1547]) );
  AND U18786 ( .A(p_input[1547]), .B(p_input[11547]), .Z(n9393) );
  AND U18787 ( .A(n9394), .B(p_input[21546]), .Z(o[1546]) );
  AND U18788 ( .A(p_input[1546]), .B(p_input[11546]), .Z(n9394) );
  AND U18789 ( .A(n9395), .B(p_input[21545]), .Z(o[1545]) );
  AND U18790 ( .A(p_input[1545]), .B(p_input[11545]), .Z(n9395) );
  AND U18791 ( .A(n9396), .B(p_input[21544]), .Z(o[1544]) );
  AND U18792 ( .A(p_input[1544]), .B(p_input[11544]), .Z(n9396) );
  AND U18793 ( .A(n9397), .B(p_input[21543]), .Z(o[1543]) );
  AND U18794 ( .A(p_input[1543]), .B(p_input[11543]), .Z(n9397) );
  AND U18795 ( .A(n9398), .B(p_input[21542]), .Z(o[1542]) );
  AND U18796 ( .A(p_input[1542]), .B(p_input[11542]), .Z(n9398) );
  AND U18797 ( .A(n9399), .B(p_input[21541]), .Z(o[1541]) );
  AND U18798 ( .A(p_input[1541]), .B(p_input[11541]), .Z(n9399) );
  AND U18799 ( .A(n9400), .B(p_input[21540]), .Z(o[1540]) );
  AND U18800 ( .A(p_input[1540]), .B(p_input[11540]), .Z(n9400) );
  AND U18801 ( .A(n9401), .B(p_input[20153]), .Z(o[153]) );
  AND U18802 ( .A(p_input[153]), .B(p_input[10153]), .Z(n9401) );
  AND U18803 ( .A(n9402), .B(p_input[21539]), .Z(o[1539]) );
  AND U18804 ( .A(p_input[1539]), .B(p_input[11539]), .Z(n9402) );
  AND U18805 ( .A(n9403), .B(p_input[21538]), .Z(o[1538]) );
  AND U18806 ( .A(p_input[1538]), .B(p_input[11538]), .Z(n9403) );
  AND U18807 ( .A(n9404), .B(p_input[21537]), .Z(o[1537]) );
  AND U18808 ( .A(p_input[1537]), .B(p_input[11537]), .Z(n9404) );
  AND U18809 ( .A(n9405), .B(p_input[21536]), .Z(o[1536]) );
  AND U18810 ( .A(p_input[1536]), .B(p_input[11536]), .Z(n9405) );
  AND U18811 ( .A(n9406), .B(p_input[21535]), .Z(o[1535]) );
  AND U18812 ( .A(p_input[1535]), .B(p_input[11535]), .Z(n9406) );
  AND U18813 ( .A(n9407), .B(p_input[21534]), .Z(o[1534]) );
  AND U18814 ( .A(p_input[1534]), .B(p_input[11534]), .Z(n9407) );
  AND U18815 ( .A(n9408), .B(p_input[21533]), .Z(o[1533]) );
  AND U18816 ( .A(p_input[1533]), .B(p_input[11533]), .Z(n9408) );
  AND U18817 ( .A(n9409), .B(p_input[21532]), .Z(o[1532]) );
  AND U18818 ( .A(p_input[1532]), .B(p_input[11532]), .Z(n9409) );
  AND U18819 ( .A(n9410), .B(p_input[21531]), .Z(o[1531]) );
  AND U18820 ( .A(p_input[1531]), .B(p_input[11531]), .Z(n9410) );
  AND U18821 ( .A(n9411), .B(p_input[21530]), .Z(o[1530]) );
  AND U18822 ( .A(p_input[1530]), .B(p_input[11530]), .Z(n9411) );
  AND U18823 ( .A(n9412), .B(p_input[20152]), .Z(o[152]) );
  AND U18824 ( .A(p_input[152]), .B(p_input[10152]), .Z(n9412) );
  AND U18825 ( .A(n9413), .B(p_input[21529]), .Z(o[1529]) );
  AND U18826 ( .A(p_input[1529]), .B(p_input[11529]), .Z(n9413) );
  AND U18827 ( .A(n9414), .B(p_input[21528]), .Z(o[1528]) );
  AND U18828 ( .A(p_input[1528]), .B(p_input[11528]), .Z(n9414) );
  AND U18829 ( .A(n9415), .B(p_input[21527]), .Z(o[1527]) );
  AND U18830 ( .A(p_input[1527]), .B(p_input[11527]), .Z(n9415) );
  AND U18831 ( .A(n9416), .B(p_input[21526]), .Z(o[1526]) );
  AND U18832 ( .A(p_input[1526]), .B(p_input[11526]), .Z(n9416) );
  AND U18833 ( .A(n9417), .B(p_input[21525]), .Z(o[1525]) );
  AND U18834 ( .A(p_input[1525]), .B(p_input[11525]), .Z(n9417) );
  AND U18835 ( .A(n9418), .B(p_input[21524]), .Z(o[1524]) );
  AND U18836 ( .A(p_input[1524]), .B(p_input[11524]), .Z(n9418) );
  AND U18837 ( .A(n9419), .B(p_input[21523]), .Z(o[1523]) );
  AND U18838 ( .A(p_input[1523]), .B(p_input[11523]), .Z(n9419) );
  AND U18839 ( .A(n9420), .B(p_input[21522]), .Z(o[1522]) );
  AND U18840 ( .A(p_input[1522]), .B(p_input[11522]), .Z(n9420) );
  AND U18841 ( .A(n9421), .B(p_input[21521]), .Z(o[1521]) );
  AND U18842 ( .A(p_input[1521]), .B(p_input[11521]), .Z(n9421) );
  AND U18843 ( .A(n9422), .B(p_input[21520]), .Z(o[1520]) );
  AND U18844 ( .A(p_input[1520]), .B(p_input[11520]), .Z(n9422) );
  AND U18845 ( .A(n9423), .B(p_input[20151]), .Z(o[151]) );
  AND U18846 ( .A(p_input[151]), .B(p_input[10151]), .Z(n9423) );
  AND U18847 ( .A(n9424), .B(p_input[21519]), .Z(o[1519]) );
  AND U18848 ( .A(p_input[1519]), .B(p_input[11519]), .Z(n9424) );
  AND U18849 ( .A(n9425), .B(p_input[21518]), .Z(o[1518]) );
  AND U18850 ( .A(p_input[1518]), .B(p_input[11518]), .Z(n9425) );
  AND U18851 ( .A(n9426), .B(p_input[21517]), .Z(o[1517]) );
  AND U18852 ( .A(p_input[1517]), .B(p_input[11517]), .Z(n9426) );
  AND U18853 ( .A(n9427), .B(p_input[21516]), .Z(o[1516]) );
  AND U18854 ( .A(p_input[1516]), .B(p_input[11516]), .Z(n9427) );
  AND U18855 ( .A(n9428), .B(p_input[21515]), .Z(o[1515]) );
  AND U18856 ( .A(p_input[1515]), .B(p_input[11515]), .Z(n9428) );
  AND U18857 ( .A(n9429), .B(p_input[21514]), .Z(o[1514]) );
  AND U18858 ( .A(p_input[1514]), .B(p_input[11514]), .Z(n9429) );
  AND U18859 ( .A(n9430), .B(p_input[21513]), .Z(o[1513]) );
  AND U18860 ( .A(p_input[1513]), .B(p_input[11513]), .Z(n9430) );
  AND U18861 ( .A(n9431), .B(p_input[21512]), .Z(o[1512]) );
  AND U18862 ( .A(p_input[1512]), .B(p_input[11512]), .Z(n9431) );
  AND U18863 ( .A(n9432), .B(p_input[21511]), .Z(o[1511]) );
  AND U18864 ( .A(p_input[1511]), .B(p_input[11511]), .Z(n9432) );
  AND U18865 ( .A(n9433), .B(p_input[21510]), .Z(o[1510]) );
  AND U18866 ( .A(p_input[1510]), .B(p_input[11510]), .Z(n9433) );
  AND U18867 ( .A(n9434), .B(p_input[20150]), .Z(o[150]) );
  AND U18868 ( .A(p_input[150]), .B(p_input[10150]), .Z(n9434) );
  AND U18869 ( .A(n9435), .B(p_input[21509]), .Z(o[1509]) );
  AND U18870 ( .A(p_input[1509]), .B(p_input[11509]), .Z(n9435) );
  AND U18871 ( .A(n9436), .B(p_input[21508]), .Z(o[1508]) );
  AND U18872 ( .A(p_input[1508]), .B(p_input[11508]), .Z(n9436) );
  AND U18873 ( .A(n9437), .B(p_input[21507]), .Z(o[1507]) );
  AND U18874 ( .A(p_input[1507]), .B(p_input[11507]), .Z(n9437) );
  AND U18875 ( .A(n9438), .B(p_input[21506]), .Z(o[1506]) );
  AND U18876 ( .A(p_input[1506]), .B(p_input[11506]), .Z(n9438) );
  AND U18877 ( .A(n9439), .B(p_input[21505]), .Z(o[1505]) );
  AND U18878 ( .A(p_input[1505]), .B(p_input[11505]), .Z(n9439) );
  AND U18879 ( .A(n9440), .B(p_input[21504]), .Z(o[1504]) );
  AND U18880 ( .A(p_input[1504]), .B(p_input[11504]), .Z(n9440) );
  AND U18881 ( .A(n9441), .B(p_input[21503]), .Z(o[1503]) );
  AND U18882 ( .A(p_input[1503]), .B(p_input[11503]), .Z(n9441) );
  AND U18883 ( .A(n9442), .B(p_input[21502]), .Z(o[1502]) );
  AND U18884 ( .A(p_input[1502]), .B(p_input[11502]), .Z(n9442) );
  AND U18885 ( .A(n9443), .B(p_input[21501]), .Z(o[1501]) );
  AND U18886 ( .A(p_input[1501]), .B(p_input[11501]), .Z(n9443) );
  AND U18887 ( .A(n9444), .B(p_input[21500]), .Z(o[1500]) );
  AND U18888 ( .A(p_input[1500]), .B(p_input[11500]), .Z(n9444) );
  AND U18889 ( .A(n9445), .B(p_input[20014]), .Z(o[14]) );
  AND U18890 ( .A(p_input[14]), .B(p_input[10014]), .Z(n9445) );
  AND U18891 ( .A(n9446), .B(p_input[20149]), .Z(o[149]) );
  AND U18892 ( .A(p_input[149]), .B(p_input[10149]), .Z(n9446) );
  AND U18893 ( .A(n9447), .B(p_input[21499]), .Z(o[1499]) );
  AND U18894 ( .A(p_input[1499]), .B(p_input[11499]), .Z(n9447) );
  AND U18895 ( .A(n9448), .B(p_input[21498]), .Z(o[1498]) );
  AND U18896 ( .A(p_input[1498]), .B(p_input[11498]), .Z(n9448) );
  AND U18897 ( .A(n9449), .B(p_input[21497]), .Z(o[1497]) );
  AND U18898 ( .A(p_input[1497]), .B(p_input[11497]), .Z(n9449) );
  AND U18899 ( .A(n9450), .B(p_input[21496]), .Z(o[1496]) );
  AND U18900 ( .A(p_input[1496]), .B(p_input[11496]), .Z(n9450) );
  AND U18901 ( .A(n9451), .B(p_input[21495]), .Z(o[1495]) );
  AND U18902 ( .A(p_input[1495]), .B(p_input[11495]), .Z(n9451) );
  AND U18903 ( .A(n9452), .B(p_input[21494]), .Z(o[1494]) );
  AND U18904 ( .A(p_input[1494]), .B(p_input[11494]), .Z(n9452) );
  AND U18905 ( .A(n9453), .B(p_input[21493]), .Z(o[1493]) );
  AND U18906 ( .A(p_input[1493]), .B(p_input[11493]), .Z(n9453) );
  AND U18907 ( .A(n9454), .B(p_input[21492]), .Z(o[1492]) );
  AND U18908 ( .A(p_input[1492]), .B(p_input[11492]), .Z(n9454) );
  AND U18909 ( .A(n9455), .B(p_input[21491]), .Z(o[1491]) );
  AND U18910 ( .A(p_input[1491]), .B(p_input[11491]), .Z(n9455) );
  AND U18911 ( .A(n9456), .B(p_input[21490]), .Z(o[1490]) );
  AND U18912 ( .A(p_input[1490]), .B(p_input[11490]), .Z(n9456) );
  AND U18913 ( .A(n9457), .B(p_input[20148]), .Z(o[148]) );
  AND U18914 ( .A(p_input[148]), .B(p_input[10148]), .Z(n9457) );
  AND U18915 ( .A(n9458), .B(p_input[21489]), .Z(o[1489]) );
  AND U18916 ( .A(p_input[1489]), .B(p_input[11489]), .Z(n9458) );
  AND U18917 ( .A(n9459), .B(p_input[21488]), .Z(o[1488]) );
  AND U18918 ( .A(p_input[1488]), .B(p_input[11488]), .Z(n9459) );
  AND U18919 ( .A(n9460), .B(p_input[21487]), .Z(o[1487]) );
  AND U18920 ( .A(p_input[1487]), .B(p_input[11487]), .Z(n9460) );
  AND U18921 ( .A(n9461), .B(p_input[21486]), .Z(o[1486]) );
  AND U18922 ( .A(p_input[1486]), .B(p_input[11486]), .Z(n9461) );
  AND U18923 ( .A(n9462), .B(p_input[21485]), .Z(o[1485]) );
  AND U18924 ( .A(p_input[1485]), .B(p_input[11485]), .Z(n9462) );
  AND U18925 ( .A(n9463), .B(p_input[21484]), .Z(o[1484]) );
  AND U18926 ( .A(p_input[1484]), .B(p_input[11484]), .Z(n9463) );
  AND U18927 ( .A(n9464), .B(p_input[21483]), .Z(o[1483]) );
  AND U18928 ( .A(p_input[1483]), .B(p_input[11483]), .Z(n9464) );
  AND U18929 ( .A(n9465), .B(p_input[21482]), .Z(o[1482]) );
  AND U18930 ( .A(p_input[1482]), .B(p_input[11482]), .Z(n9465) );
  AND U18931 ( .A(n9466), .B(p_input[21481]), .Z(o[1481]) );
  AND U18932 ( .A(p_input[1481]), .B(p_input[11481]), .Z(n9466) );
  AND U18933 ( .A(n9467), .B(p_input[21480]), .Z(o[1480]) );
  AND U18934 ( .A(p_input[1480]), .B(p_input[11480]), .Z(n9467) );
  AND U18935 ( .A(n9468), .B(p_input[20147]), .Z(o[147]) );
  AND U18936 ( .A(p_input[147]), .B(p_input[10147]), .Z(n9468) );
  AND U18937 ( .A(n9469), .B(p_input[21479]), .Z(o[1479]) );
  AND U18938 ( .A(p_input[1479]), .B(p_input[11479]), .Z(n9469) );
  AND U18939 ( .A(n9470), .B(p_input[21478]), .Z(o[1478]) );
  AND U18940 ( .A(p_input[1478]), .B(p_input[11478]), .Z(n9470) );
  AND U18941 ( .A(n9471), .B(p_input[21477]), .Z(o[1477]) );
  AND U18942 ( .A(p_input[1477]), .B(p_input[11477]), .Z(n9471) );
  AND U18943 ( .A(n9472), .B(p_input[21476]), .Z(o[1476]) );
  AND U18944 ( .A(p_input[1476]), .B(p_input[11476]), .Z(n9472) );
  AND U18945 ( .A(n9473), .B(p_input[21475]), .Z(o[1475]) );
  AND U18946 ( .A(p_input[1475]), .B(p_input[11475]), .Z(n9473) );
  AND U18947 ( .A(n9474), .B(p_input[21474]), .Z(o[1474]) );
  AND U18948 ( .A(p_input[1474]), .B(p_input[11474]), .Z(n9474) );
  AND U18949 ( .A(n9475), .B(p_input[21473]), .Z(o[1473]) );
  AND U18950 ( .A(p_input[1473]), .B(p_input[11473]), .Z(n9475) );
  AND U18951 ( .A(n9476), .B(p_input[21472]), .Z(o[1472]) );
  AND U18952 ( .A(p_input[1472]), .B(p_input[11472]), .Z(n9476) );
  AND U18953 ( .A(n9477), .B(p_input[21471]), .Z(o[1471]) );
  AND U18954 ( .A(p_input[1471]), .B(p_input[11471]), .Z(n9477) );
  AND U18955 ( .A(n9478), .B(p_input[21470]), .Z(o[1470]) );
  AND U18956 ( .A(p_input[1470]), .B(p_input[11470]), .Z(n9478) );
  AND U18957 ( .A(n9479), .B(p_input[20146]), .Z(o[146]) );
  AND U18958 ( .A(p_input[146]), .B(p_input[10146]), .Z(n9479) );
  AND U18959 ( .A(n9480), .B(p_input[21469]), .Z(o[1469]) );
  AND U18960 ( .A(p_input[1469]), .B(p_input[11469]), .Z(n9480) );
  AND U18961 ( .A(n9481), .B(p_input[21468]), .Z(o[1468]) );
  AND U18962 ( .A(p_input[1468]), .B(p_input[11468]), .Z(n9481) );
  AND U18963 ( .A(n9482), .B(p_input[21467]), .Z(o[1467]) );
  AND U18964 ( .A(p_input[1467]), .B(p_input[11467]), .Z(n9482) );
  AND U18965 ( .A(n9483), .B(p_input[21466]), .Z(o[1466]) );
  AND U18966 ( .A(p_input[1466]), .B(p_input[11466]), .Z(n9483) );
  AND U18967 ( .A(n9484), .B(p_input[21465]), .Z(o[1465]) );
  AND U18968 ( .A(p_input[1465]), .B(p_input[11465]), .Z(n9484) );
  AND U18969 ( .A(n9485), .B(p_input[21464]), .Z(o[1464]) );
  AND U18970 ( .A(p_input[1464]), .B(p_input[11464]), .Z(n9485) );
  AND U18971 ( .A(n9486), .B(p_input[21463]), .Z(o[1463]) );
  AND U18972 ( .A(p_input[1463]), .B(p_input[11463]), .Z(n9486) );
  AND U18973 ( .A(n9487), .B(p_input[21462]), .Z(o[1462]) );
  AND U18974 ( .A(p_input[1462]), .B(p_input[11462]), .Z(n9487) );
  AND U18975 ( .A(n9488), .B(p_input[21461]), .Z(o[1461]) );
  AND U18976 ( .A(p_input[1461]), .B(p_input[11461]), .Z(n9488) );
  AND U18977 ( .A(n9489), .B(p_input[21460]), .Z(o[1460]) );
  AND U18978 ( .A(p_input[1460]), .B(p_input[11460]), .Z(n9489) );
  AND U18979 ( .A(n9490), .B(p_input[20145]), .Z(o[145]) );
  AND U18980 ( .A(p_input[145]), .B(p_input[10145]), .Z(n9490) );
  AND U18981 ( .A(n9491), .B(p_input[21459]), .Z(o[1459]) );
  AND U18982 ( .A(p_input[1459]), .B(p_input[11459]), .Z(n9491) );
  AND U18983 ( .A(n9492), .B(p_input[21458]), .Z(o[1458]) );
  AND U18984 ( .A(p_input[1458]), .B(p_input[11458]), .Z(n9492) );
  AND U18985 ( .A(n9493), .B(p_input[21457]), .Z(o[1457]) );
  AND U18986 ( .A(p_input[1457]), .B(p_input[11457]), .Z(n9493) );
  AND U18987 ( .A(n9494), .B(p_input[21456]), .Z(o[1456]) );
  AND U18988 ( .A(p_input[1456]), .B(p_input[11456]), .Z(n9494) );
  AND U18989 ( .A(n9495), .B(p_input[21455]), .Z(o[1455]) );
  AND U18990 ( .A(p_input[1455]), .B(p_input[11455]), .Z(n9495) );
  AND U18991 ( .A(n9496), .B(p_input[21454]), .Z(o[1454]) );
  AND U18992 ( .A(p_input[1454]), .B(p_input[11454]), .Z(n9496) );
  AND U18993 ( .A(n9497), .B(p_input[21453]), .Z(o[1453]) );
  AND U18994 ( .A(p_input[1453]), .B(p_input[11453]), .Z(n9497) );
  AND U18995 ( .A(n9498), .B(p_input[21452]), .Z(o[1452]) );
  AND U18996 ( .A(p_input[1452]), .B(p_input[11452]), .Z(n9498) );
  AND U18997 ( .A(n9499), .B(p_input[21451]), .Z(o[1451]) );
  AND U18998 ( .A(p_input[1451]), .B(p_input[11451]), .Z(n9499) );
  AND U18999 ( .A(n9500), .B(p_input[21450]), .Z(o[1450]) );
  AND U19000 ( .A(p_input[1450]), .B(p_input[11450]), .Z(n9500) );
  AND U19001 ( .A(n9501), .B(p_input[20144]), .Z(o[144]) );
  AND U19002 ( .A(p_input[144]), .B(p_input[10144]), .Z(n9501) );
  AND U19003 ( .A(n9502), .B(p_input[21449]), .Z(o[1449]) );
  AND U19004 ( .A(p_input[1449]), .B(p_input[11449]), .Z(n9502) );
  AND U19005 ( .A(n9503), .B(p_input[21448]), .Z(o[1448]) );
  AND U19006 ( .A(p_input[1448]), .B(p_input[11448]), .Z(n9503) );
  AND U19007 ( .A(n9504), .B(p_input[21447]), .Z(o[1447]) );
  AND U19008 ( .A(p_input[1447]), .B(p_input[11447]), .Z(n9504) );
  AND U19009 ( .A(n9505), .B(p_input[21446]), .Z(o[1446]) );
  AND U19010 ( .A(p_input[1446]), .B(p_input[11446]), .Z(n9505) );
  AND U19011 ( .A(n9506), .B(p_input[21445]), .Z(o[1445]) );
  AND U19012 ( .A(p_input[1445]), .B(p_input[11445]), .Z(n9506) );
  AND U19013 ( .A(n9507), .B(p_input[21444]), .Z(o[1444]) );
  AND U19014 ( .A(p_input[1444]), .B(p_input[11444]), .Z(n9507) );
  AND U19015 ( .A(n9508), .B(p_input[21443]), .Z(o[1443]) );
  AND U19016 ( .A(p_input[1443]), .B(p_input[11443]), .Z(n9508) );
  AND U19017 ( .A(n9509), .B(p_input[21442]), .Z(o[1442]) );
  AND U19018 ( .A(p_input[1442]), .B(p_input[11442]), .Z(n9509) );
  AND U19019 ( .A(n9510), .B(p_input[21441]), .Z(o[1441]) );
  AND U19020 ( .A(p_input[1441]), .B(p_input[11441]), .Z(n9510) );
  AND U19021 ( .A(n9511), .B(p_input[21440]), .Z(o[1440]) );
  AND U19022 ( .A(p_input[1440]), .B(p_input[11440]), .Z(n9511) );
  AND U19023 ( .A(n9512), .B(p_input[20143]), .Z(o[143]) );
  AND U19024 ( .A(p_input[143]), .B(p_input[10143]), .Z(n9512) );
  AND U19025 ( .A(n9513), .B(p_input[21439]), .Z(o[1439]) );
  AND U19026 ( .A(p_input[1439]), .B(p_input[11439]), .Z(n9513) );
  AND U19027 ( .A(n9514), .B(p_input[21438]), .Z(o[1438]) );
  AND U19028 ( .A(p_input[1438]), .B(p_input[11438]), .Z(n9514) );
  AND U19029 ( .A(n9515), .B(p_input[21437]), .Z(o[1437]) );
  AND U19030 ( .A(p_input[1437]), .B(p_input[11437]), .Z(n9515) );
  AND U19031 ( .A(n9516), .B(p_input[21436]), .Z(o[1436]) );
  AND U19032 ( .A(p_input[1436]), .B(p_input[11436]), .Z(n9516) );
  AND U19033 ( .A(n9517), .B(p_input[21435]), .Z(o[1435]) );
  AND U19034 ( .A(p_input[1435]), .B(p_input[11435]), .Z(n9517) );
  AND U19035 ( .A(n9518), .B(p_input[21434]), .Z(o[1434]) );
  AND U19036 ( .A(p_input[1434]), .B(p_input[11434]), .Z(n9518) );
  AND U19037 ( .A(n9519), .B(p_input[21433]), .Z(o[1433]) );
  AND U19038 ( .A(p_input[1433]), .B(p_input[11433]), .Z(n9519) );
  AND U19039 ( .A(n9520), .B(p_input[21432]), .Z(o[1432]) );
  AND U19040 ( .A(p_input[1432]), .B(p_input[11432]), .Z(n9520) );
  AND U19041 ( .A(n9521), .B(p_input[21431]), .Z(o[1431]) );
  AND U19042 ( .A(p_input[1431]), .B(p_input[11431]), .Z(n9521) );
  AND U19043 ( .A(n9522), .B(p_input[21430]), .Z(o[1430]) );
  AND U19044 ( .A(p_input[1430]), .B(p_input[11430]), .Z(n9522) );
  AND U19045 ( .A(n9523), .B(p_input[20142]), .Z(o[142]) );
  AND U19046 ( .A(p_input[142]), .B(p_input[10142]), .Z(n9523) );
  AND U19047 ( .A(n9524), .B(p_input[21429]), .Z(o[1429]) );
  AND U19048 ( .A(p_input[1429]), .B(p_input[11429]), .Z(n9524) );
  AND U19049 ( .A(n9525), .B(p_input[21428]), .Z(o[1428]) );
  AND U19050 ( .A(p_input[1428]), .B(p_input[11428]), .Z(n9525) );
  AND U19051 ( .A(n9526), .B(p_input[21427]), .Z(o[1427]) );
  AND U19052 ( .A(p_input[1427]), .B(p_input[11427]), .Z(n9526) );
  AND U19053 ( .A(n9527), .B(p_input[21426]), .Z(o[1426]) );
  AND U19054 ( .A(p_input[1426]), .B(p_input[11426]), .Z(n9527) );
  AND U19055 ( .A(n9528), .B(p_input[21425]), .Z(o[1425]) );
  AND U19056 ( .A(p_input[1425]), .B(p_input[11425]), .Z(n9528) );
  AND U19057 ( .A(n9529), .B(p_input[21424]), .Z(o[1424]) );
  AND U19058 ( .A(p_input[1424]), .B(p_input[11424]), .Z(n9529) );
  AND U19059 ( .A(n9530), .B(p_input[21423]), .Z(o[1423]) );
  AND U19060 ( .A(p_input[1423]), .B(p_input[11423]), .Z(n9530) );
  AND U19061 ( .A(n9531), .B(p_input[21422]), .Z(o[1422]) );
  AND U19062 ( .A(p_input[1422]), .B(p_input[11422]), .Z(n9531) );
  AND U19063 ( .A(n9532), .B(p_input[21421]), .Z(o[1421]) );
  AND U19064 ( .A(p_input[1421]), .B(p_input[11421]), .Z(n9532) );
  AND U19065 ( .A(n9533), .B(p_input[21420]), .Z(o[1420]) );
  AND U19066 ( .A(p_input[1420]), .B(p_input[11420]), .Z(n9533) );
  AND U19067 ( .A(n9534), .B(p_input[20141]), .Z(o[141]) );
  AND U19068 ( .A(p_input[141]), .B(p_input[10141]), .Z(n9534) );
  AND U19069 ( .A(n9535), .B(p_input[21419]), .Z(o[1419]) );
  AND U19070 ( .A(p_input[1419]), .B(p_input[11419]), .Z(n9535) );
  AND U19071 ( .A(n9536), .B(p_input[21418]), .Z(o[1418]) );
  AND U19072 ( .A(p_input[1418]), .B(p_input[11418]), .Z(n9536) );
  AND U19073 ( .A(n9537), .B(p_input[21417]), .Z(o[1417]) );
  AND U19074 ( .A(p_input[1417]), .B(p_input[11417]), .Z(n9537) );
  AND U19075 ( .A(n9538), .B(p_input[21416]), .Z(o[1416]) );
  AND U19076 ( .A(p_input[1416]), .B(p_input[11416]), .Z(n9538) );
  AND U19077 ( .A(n9539), .B(p_input[21415]), .Z(o[1415]) );
  AND U19078 ( .A(p_input[1415]), .B(p_input[11415]), .Z(n9539) );
  AND U19079 ( .A(n9540), .B(p_input[21414]), .Z(o[1414]) );
  AND U19080 ( .A(p_input[1414]), .B(p_input[11414]), .Z(n9540) );
  AND U19081 ( .A(n9541), .B(p_input[21413]), .Z(o[1413]) );
  AND U19082 ( .A(p_input[1413]), .B(p_input[11413]), .Z(n9541) );
  AND U19083 ( .A(n9542), .B(p_input[21412]), .Z(o[1412]) );
  AND U19084 ( .A(p_input[1412]), .B(p_input[11412]), .Z(n9542) );
  AND U19085 ( .A(n9543), .B(p_input[21411]), .Z(o[1411]) );
  AND U19086 ( .A(p_input[1411]), .B(p_input[11411]), .Z(n9543) );
  AND U19087 ( .A(n9544), .B(p_input[21410]), .Z(o[1410]) );
  AND U19088 ( .A(p_input[1410]), .B(p_input[11410]), .Z(n9544) );
  AND U19089 ( .A(n9545), .B(p_input[20140]), .Z(o[140]) );
  AND U19090 ( .A(p_input[140]), .B(p_input[10140]), .Z(n9545) );
  AND U19091 ( .A(n9546), .B(p_input[21409]), .Z(o[1409]) );
  AND U19092 ( .A(p_input[1409]), .B(p_input[11409]), .Z(n9546) );
  AND U19093 ( .A(n9547), .B(p_input[21408]), .Z(o[1408]) );
  AND U19094 ( .A(p_input[1408]), .B(p_input[11408]), .Z(n9547) );
  AND U19095 ( .A(n9548), .B(p_input[21407]), .Z(o[1407]) );
  AND U19096 ( .A(p_input[1407]), .B(p_input[11407]), .Z(n9548) );
  AND U19097 ( .A(n9549), .B(p_input[21406]), .Z(o[1406]) );
  AND U19098 ( .A(p_input[1406]), .B(p_input[11406]), .Z(n9549) );
  AND U19099 ( .A(n9550), .B(p_input[21405]), .Z(o[1405]) );
  AND U19100 ( .A(p_input[1405]), .B(p_input[11405]), .Z(n9550) );
  AND U19101 ( .A(n9551), .B(p_input[21404]), .Z(o[1404]) );
  AND U19102 ( .A(p_input[1404]), .B(p_input[11404]), .Z(n9551) );
  AND U19103 ( .A(n9552), .B(p_input[21403]), .Z(o[1403]) );
  AND U19104 ( .A(p_input[1403]), .B(p_input[11403]), .Z(n9552) );
  AND U19105 ( .A(n9553), .B(p_input[21402]), .Z(o[1402]) );
  AND U19106 ( .A(p_input[1402]), .B(p_input[11402]), .Z(n9553) );
  AND U19107 ( .A(n9554), .B(p_input[21401]), .Z(o[1401]) );
  AND U19108 ( .A(p_input[1401]), .B(p_input[11401]), .Z(n9554) );
  AND U19109 ( .A(n9555), .B(p_input[21400]), .Z(o[1400]) );
  AND U19110 ( .A(p_input[1400]), .B(p_input[11400]), .Z(n9555) );
  AND U19111 ( .A(n9556), .B(p_input[20013]), .Z(o[13]) );
  AND U19112 ( .A(p_input[13]), .B(p_input[10013]), .Z(n9556) );
  AND U19113 ( .A(n9557), .B(p_input[20139]), .Z(o[139]) );
  AND U19114 ( .A(p_input[139]), .B(p_input[10139]), .Z(n9557) );
  AND U19115 ( .A(n9558), .B(p_input[21399]), .Z(o[1399]) );
  AND U19116 ( .A(p_input[1399]), .B(p_input[11399]), .Z(n9558) );
  AND U19117 ( .A(n9559), .B(p_input[21398]), .Z(o[1398]) );
  AND U19118 ( .A(p_input[1398]), .B(p_input[11398]), .Z(n9559) );
  AND U19119 ( .A(n9560), .B(p_input[21397]), .Z(o[1397]) );
  AND U19120 ( .A(p_input[1397]), .B(p_input[11397]), .Z(n9560) );
  AND U19121 ( .A(n9561), .B(p_input[21396]), .Z(o[1396]) );
  AND U19122 ( .A(p_input[1396]), .B(p_input[11396]), .Z(n9561) );
  AND U19123 ( .A(n9562), .B(p_input[21395]), .Z(o[1395]) );
  AND U19124 ( .A(p_input[1395]), .B(p_input[11395]), .Z(n9562) );
  AND U19125 ( .A(n9563), .B(p_input[21394]), .Z(o[1394]) );
  AND U19126 ( .A(p_input[1394]), .B(p_input[11394]), .Z(n9563) );
  AND U19127 ( .A(n9564), .B(p_input[21393]), .Z(o[1393]) );
  AND U19128 ( .A(p_input[1393]), .B(p_input[11393]), .Z(n9564) );
  AND U19129 ( .A(n9565), .B(p_input[21392]), .Z(o[1392]) );
  AND U19130 ( .A(p_input[1392]), .B(p_input[11392]), .Z(n9565) );
  AND U19131 ( .A(n9566), .B(p_input[21391]), .Z(o[1391]) );
  AND U19132 ( .A(p_input[1391]), .B(p_input[11391]), .Z(n9566) );
  AND U19133 ( .A(n9567), .B(p_input[21390]), .Z(o[1390]) );
  AND U19134 ( .A(p_input[1390]), .B(p_input[11390]), .Z(n9567) );
  AND U19135 ( .A(n9568), .B(p_input[20138]), .Z(o[138]) );
  AND U19136 ( .A(p_input[138]), .B(p_input[10138]), .Z(n9568) );
  AND U19137 ( .A(n9569), .B(p_input[21389]), .Z(o[1389]) );
  AND U19138 ( .A(p_input[1389]), .B(p_input[11389]), .Z(n9569) );
  AND U19139 ( .A(n9570), .B(p_input[21388]), .Z(o[1388]) );
  AND U19140 ( .A(p_input[1388]), .B(p_input[11388]), .Z(n9570) );
  AND U19141 ( .A(n9571), .B(p_input[21387]), .Z(o[1387]) );
  AND U19142 ( .A(p_input[1387]), .B(p_input[11387]), .Z(n9571) );
  AND U19143 ( .A(n9572), .B(p_input[21386]), .Z(o[1386]) );
  AND U19144 ( .A(p_input[1386]), .B(p_input[11386]), .Z(n9572) );
  AND U19145 ( .A(n9573), .B(p_input[21385]), .Z(o[1385]) );
  AND U19146 ( .A(p_input[1385]), .B(p_input[11385]), .Z(n9573) );
  AND U19147 ( .A(n9574), .B(p_input[21384]), .Z(o[1384]) );
  AND U19148 ( .A(p_input[1384]), .B(p_input[11384]), .Z(n9574) );
  AND U19149 ( .A(n9575), .B(p_input[21383]), .Z(o[1383]) );
  AND U19150 ( .A(p_input[1383]), .B(p_input[11383]), .Z(n9575) );
  AND U19151 ( .A(n9576), .B(p_input[21382]), .Z(o[1382]) );
  AND U19152 ( .A(p_input[1382]), .B(p_input[11382]), .Z(n9576) );
  AND U19153 ( .A(n9577), .B(p_input[21381]), .Z(o[1381]) );
  AND U19154 ( .A(p_input[1381]), .B(p_input[11381]), .Z(n9577) );
  AND U19155 ( .A(n9578), .B(p_input[21380]), .Z(o[1380]) );
  AND U19156 ( .A(p_input[1380]), .B(p_input[11380]), .Z(n9578) );
  AND U19157 ( .A(n9579), .B(p_input[20137]), .Z(o[137]) );
  AND U19158 ( .A(p_input[137]), .B(p_input[10137]), .Z(n9579) );
  AND U19159 ( .A(n9580), .B(p_input[21379]), .Z(o[1379]) );
  AND U19160 ( .A(p_input[1379]), .B(p_input[11379]), .Z(n9580) );
  AND U19161 ( .A(n9581), .B(p_input[21378]), .Z(o[1378]) );
  AND U19162 ( .A(p_input[1378]), .B(p_input[11378]), .Z(n9581) );
  AND U19163 ( .A(n9582), .B(p_input[21377]), .Z(o[1377]) );
  AND U19164 ( .A(p_input[1377]), .B(p_input[11377]), .Z(n9582) );
  AND U19165 ( .A(n9583), .B(p_input[21376]), .Z(o[1376]) );
  AND U19166 ( .A(p_input[1376]), .B(p_input[11376]), .Z(n9583) );
  AND U19167 ( .A(n9584), .B(p_input[21375]), .Z(o[1375]) );
  AND U19168 ( .A(p_input[1375]), .B(p_input[11375]), .Z(n9584) );
  AND U19169 ( .A(n9585), .B(p_input[21374]), .Z(o[1374]) );
  AND U19170 ( .A(p_input[1374]), .B(p_input[11374]), .Z(n9585) );
  AND U19171 ( .A(n9586), .B(p_input[21373]), .Z(o[1373]) );
  AND U19172 ( .A(p_input[1373]), .B(p_input[11373]), .Z(n9586) );
  AND U19173 ( .A(n9587), .B(p_input[21372]), .Z(o[1372]) );
  AND U19174 ( .A(p_input[1372]), .B(p_input[11372]), .Z(n9587) );
  AND U19175 ( .A(n9588), .B(p_input[21371]), .Z(o[1371]) );
  AND U19176 ( .A(p_input[1371]), .B(p_input[11371]), .Z(n9588) );
  AND U19177 ( .A(n9589), .B(p_input[21370]), .Z(o[1370]) );
  AND U19178 ( .A(p_input[1370]), .B(p_input[11370]), .Z(n9589) );
  AND U19179 ( .A(n9590), .B(p_input[20136]), .Z(o[136]) );
  AND U19180 ( .A(p_input[136]), .B(p_input[10136]), .Z(n9590) );
  AND U19181 ( .A(n9591), .B(p_input[21369]), .Z(o[1369]) );
  AND U19182 ( .A(p_input[1369]), .B(p_input[11369]), .Z(n9591) );
  AND U19183 ( .A(n9592), .B(p_input[21368]), .Z(o[1368]) );
  AND U19184 ( .A(p_input[1368]), .B(p_input[11368]), .Z(n9592) );
  AND U19185 ( .A(n9593), .B(p_input[21367]), .Z(o[1367]) );
  AND U19186 ( .A(p_input[1367]), .B(p_input[11367]), .Z(n9593) );
  AND U19187 ( .A(n9594), .B(p_input[21366]), .Z(o[1366]) );
  AND U19188 ( .A(p_input[1366]), .B(p_input[11366]), .Z(n9594) );
  AND U19189 ( .A(n9595), .B(p_input[21365]), .Z(o[1365]) );
  AND U19190 ( .A(p_input[1365]), .B(p_input[11365]), .Z(n9595) );
  AND U19191 ( .A(n9596), .B(p_input[21364]), .Z(o[1364]) );
  AND U19192 ( .A(p_input[1364]), .B(p_input[11364]), .Z(n9596) );
  AND U19193 ( .A(n9597), .B(p_input[21363]), .Z(o[1363]) );
  AND U19194 ( .A(p_input[1363]), .B(p_input[11363]), .Z(n9597) );
  AND U19195 ( .A(n9598), .B(p_input[21362]), .Z(o[1362]) );
  AND U19196 ( .A(p_input[1362]), .B(p_input[11362]), .Z(n9598) );
  AND U19197 ( .A(n9599), .B(p_input[21361]), .Z(o[1361]) );
  AND U19198 ( .A(p_input[1361]), .B(p_input[11361]), .Z(n9599) );
  AND U19199 ( .A(n9600), .B(p_input[21360]), .Z(o[1360]) );
  AND U19200 ( .A(p_input[1360]), .B(p_input[11360]), .Z(n9600) );
  AND U19201 ( .A(n9601), .B(p_input[20135]), .Z(o[135]) );
  AND U19202 ( .A(p_input[135]), .B(p_input[10135]), .Z(n9601) );
  AND U19203 ( .A(n9602), .B(p_input[21359]), .Z(o[1359]) );
  AND U19204 ( .A(p_input[1359]), .B(p_input[11359]), .Z(n9602) );
  AND U19205 ( .A(n9603), .B(p_input[21358]), .Z(o[1358]) );
  AND U19206 ( .A(p_input[1358]), .B(p_input[11358]), .Z(n9603) );
  AND U19207 ( .A(n9604), .B(p_input[21357]), .Z(o[1357]) );
  AND U19208 ( .A(p_input[1357]), .B(p_input[11357]), .Z(n9604) );
  AND U19209 ( .A(n9605), .B(p_input[21356]), .Z(o[1356]) );
  AND U19210 ( .A(p_input[1356]), .B(p_input[11356]), .Z(n9605) );
  AND U19211 ( .A(n9606), .B(p_input[21355]), .Z(o[1355]) );
  AND U19212 ( .A(p_input[1355]), .B(p_input[11355]), .Z(n9606) );
  AND U19213 ( .A(n9607), .B(p_input[21354]), .Z(o[1354]) );
  AND U19214 ( .A(p_input[1354]), .B(p_input[11354]), .Z(n9607) );
  AND U19215 ( .A(n9608), .B(p_input[21353]), .Z(o[1353]) );
  AND U19216 ( .A(p_input[1353]), .B(p_input[11353]), .Z(n9608) );
  AND U19217 ( .A(n9609), .B(p_input[21352]), .Z(o[1352]) );
  AND U19218 ( .A(p_input[1352]), .B(p_input[11352]), .Z(n9609) );
  AND U19219 ( .A(n9610), .B(p_input[21351]), .Z(o[1351]) );
  AND U19220 ( .A(p_input[1351]), .B(p_input[11351]), .Z(n9610) );
  AND U19221 ( .A(n9611), .B(p_input[21350]), .Z(o[1350]) );
  AND U19222 ( .A(p_input[1350]), .B(p_input[11350]), .Z(n9611) );
  AND U19223 ( .A(n9612), .B(p_input[20134]), .Z(o[134]) );
  AND U19224 ( .A(p_input[134]), .B(p_input[10134]), .Z(n9612) );
  AND U19225 ( .A(n9613), .B(p_input[21349]), .Z(o[1349]) );
  AND U19226 ( .A(p_input[1349]), .B(p_input[11349]), .Z(n9613) );
  AND U19227 ( .A(n9614), .B(p_input[21348]), .Z(o[1348]) );
  AND U19228 ( .A(p_input[1348]), .B(p_input[11348]), .Z(n9614) );
  AND U19229 ( .A(n9615), .B(p_input[21347]), .Z(o[1347]) );
  AND U19230 ( .A(p_input[1347]), .B(p_input[11347]), .Z(n9615) );
  AND U19231 ( .A(n9616), .B(p_input[21346]), .Z(o[1346]) );
  AND U19232 ( .A(p_input[1346]), .B(p_input[11346]), .Z(n9616) );
  AND U19233 ( .A(n9617), .B(p_input[21345]), .Z(o[1345]) );
  AND U19234 ( .A(p_input[1345]), .B(p_input[11345]), .Z(n9617) );
  AND U19235 ( .A(n9618), .B(p_input[21344]), .Z(o[1344]) );
  AND U19236 ( .A(p_input[1344]), .B(p_input[11344]), .Z(n9618) );
  AND U19237 ( .A(n9619), .B(p_input[21343]), .Z(o[1343]) );
  AND U19238 ( .A(p_input[1343]), .B(p_input[11343]), .Z(n9619) );
  AND U19239 ( .A(n9620), .B(p_input[21342]), .Z(o[1342]) );
  AND U19240 ( .A(p_input[1342]), .B(p_input[11342]), .Z(n9620) );
  AND U19241 ( .A(n9621), .B(p_input[21341]), .Z(o[1341]) );
  AND U19242 ( .A(p_input[1341]), .B(p_input[11341]), .Z(n9621) );
  AND U19243 ( .A(n9622), .B(p_input[21340]), .Z(o[1340]) );
  AND U19244 ( .A(p_input[1340]), .B(p_input[11340]), .Z(n9622) );
  AND U19245 ( .A(n9623), .B(p_input[20133]), .Z(o[133]) );
  AND U19246 ( .A(p_input[133]), .B(p_input[10133]), .Z(n9623) );
  AND U19247 ( .A(n9624), .B(p_input[21339]), .Z(o[1339]) );
  AND U19248 ( .A(p_input[1339]), .B(p_input[11339]), .Z(n9624) );
  AND U19249 ( .A(n9625), .B(p_input[21338]), .Z(o[1338]) );
  AND U19250 ( .A(p_input[1338]), .B(p_input[11338]), .Z(n9625) );
  AND U19251 ( .A(n9626), .B(p_input[21337]), .Z(o[1337]) );
  AND U19252 ( .A(p_input[1337]), .B(p_input[11337]), .Z(n9626) );
  AND U19253 ( .A(n9627), .B(p_input[21336]), .Z(o[1336]) );
  AND U19254 ( .A(p_input[1336]), .B(p_input[11336]), .Z(n9627) );
  AND U19255 ( .A(n9628), .B(p_input[21335]), .Z(o[1335]) );
  AND U19256 ( .A(p_input[1335]), .B(p_input[11335]), .Z(n9628) );
  AND U19257 ( .A(n9629), .B(p_input[21334]), .Z(o[1334]) );
  AND U19258 ( .A(p_input[1334]), .B(p_input[11334]), .Z(n9629) );
  AND U19259 ( .A(n9630), .B(p_input[21333]), .Z(o[1333]) );
  AND U19260 ( .A(p_input[1333]), .B(p_input[11333]), .Z(n9630) );
  AND U19261 ( .A(n9631), .B(p_input[21332]), .Z(o[1332]) );
  AND U19262 ( .A(p_input[1332]), .B(p_input[11332]), .Z(n9631) );
  AND U19263 ( .A(n9632), .B(p_input[21331]), .Z(o[1331]) );
  AND U19264 ( .A(p_input[1331]), .B(p_input[11331]), .Z(n9632) );
  AND U19265 ( .A(n9633), .B(p_input[21330]), .Z(o[1330]) );
  AND U19266 ( .A(p_input[1330]), .B(p_input[11330]), .Z(n9633) );
  AND U19267 ( .A(n9634), .B(p_input[20132]), .Z(o[132]) );
  AND U19268 ( .A(p_input[132]), .B(p_input[10132]), .Z(n9634) );
  AND U19269 ( .A(n9635), .B(p_input[21329]), .Z(o[1329]) );
  AND U19270 ( .A(p_input[1329]), .B(p_input[11329]), .Z(n9635) );
  AND U19271 ( .A(n9636), .B(p_input[21328]), .Z(o[1328]) );
  AND U19272 ( .A(p_input[1328]), .B(p_input[11328]), .Z(n9636) );
  AND U19273 ( .A(n9637), .B(p_input[21327]), .Z(o[1327]) );
  AND U19274 ( .A(p_input[1327]), .B(p_input[11327]), .Z(n9637) );
  AND U19275 ( .A(n9638), .B(p_input[21326]), .Z(o[1326]) );
  AND U19276 ( .A(p_input[1326]), .B(p_input[11326]), .Z(n9638) );
  AND U19277 ( .A(n9639), .B(p_input[21325]), .Z(o[1325]) );
  AND U19278 ( .A(p_input[1325]), .B(p_input[11325]), .Z(n9639) );
  AND U19279 ( .A(n9640), .B(p_input[21324]), .Z(o[1324]) );
  AND U19280 ( .A(p_input[1324]), .B(p_input[11324]), .Z(n9640) );
  AND U19281 ( .A(n9641), .B(p_input[21323]), .Z(o[1323]) );
  AND U19282 ( .A(p_input[1323]), .B(p_input[11323]), .Z(n9641) );
  AND U19283 ( .A(n9642), .B(p_input[21322]), .Z(o[1322]) );
  AND U19284 ( .A(p_input[1322]), .B(p_input[11322]), .Z(n9642) );
  AND U19285 ( .A(n9643), .B(p_input[21321]), .Z(o[1321]) );
  AND U19286 ( .A(p_input[1321]), .B(p_input[11321]), .Z(n9643) );
  AND U19287 ( .A(n9644), .B(p_input[21320]), .Z(o[1320]) );
  AND U19288 ( .A(p_input[1320]), .B(p_input[11320]), .Z(n9644) );
  AND U19289 ( .A(n9645), .B(p_input[20131]), .Z(o[131]) );
  AND U19290 ( .A(p_input[131]), .B(p_input[10131]), .Z(n9645) );
  AND U19291 ( .A(n9646), .B(p_input[21319]), .Z(o[1319]) );
  AND U19292 ( .A(p_input[1319]), .B(p_input[11319]), .Z(n9646) );
  AND U19293 ( .A(n9647), .B(p_input[21318]), .Z(o[1318]) );
  AND U19294 ( .A(p_input[1318]), .B(p_input[11318]), .Z(n9647) );
  AND U19295 ( .A(n9648), .B(p_input[21317]), .Z(o[1317]) );
  AND U19296 ( .A(p_input[1317]), .B(p_input[11317]), .Z(n9648) );
  AND U19297 ( .A(n9649), .B(p_input[21316]), .Z(o[1316]) );
  AND U19298 ( .A(p_input[1316]), .B(p_input[11316]), .Z(n9649) );
  AND U19299 ( .A(n9650), .B(p_input[21315]), .Z(o[1315]) );
  AND U19300 ( .A(p_input[1315]), .B(p_input[11315]), .Z(n9650) );
  AND U19301 ( .A(n9651), .B(p_input[21314]), .Z(o[1314]) );
  AND U19302 ( .A(p_input[1314]), .B(p_input[11314]), .Z(n9651) );
  AND U19303 ( .A(n9652), .B(p_input[21313]), .Z(o[1313]) );
  AND U19304 ( .A(p_input[1313]), .B(p_input[11313]), .Z(n9652) );
  AND U19305 ( .A(n9653), .B(p_input[21312]), .Z(o[1312]) );
  AND U19306 ( .A(p_input[1312]), .B(p_input[11312]), .Z(n9653) );
  AND U19307 ( .A(n9654), .B(p_input[21311]), .Z(o[1311]) );
  AND U19308 ( .A(p_input[1311]), .B(p_input[11311]), .Z(n9654) );
  AND U19309 ( .A(n9655), .B(p_input[21310]), .Z(o[1310]) );
  AND U19310 ( .A(p_input[1310]), .B(p_input[11310]), .Z(n9655) );
  AND U19311 ( .A(n9656), .B(p_input[20130]), .Z(o[130]) );
  AND U19312 ( .A(p_input[130]), .B(p_input[10130]), .Z(n9656) );
  AND U19313 ( .A(n9657), .B(p_input[21309]), .Z(o[1309]) );
  AND U19314 ( .A(p_input[1309]), .B(p_input[11309]), .Z(n9657) );
  AND U19315 ( .A(n9658), .B(p_input[21308]), .Z(o[1308]) );
  AND U19316 ( .A(p_input[1308]), .B(p_input[11308]), .Z(n9658) );
  AND U19317 ( .A(n9659), .B(p_input[21307]), .Z(o[1307]) );
  AND U19318 ( .A(p_input[1307]), .B(p_input[11307]), .Z(n9659) );
  AND U19319 ( .A(n9660), .B(p_input[21306]), .Z(o[1306]) );
  AND U19320 ( .A(p_input[1306]), .B(p_input[11306]), .Z(n9660) );
  AND U19321 ( .A(n9661), .B(p_input[21305]), .Z(o[1305]) );
  AND U19322 ( .A(p_input[1305]), .B(p_input[11305]), .Z(n9661) );
  AND U19323 ( .A(n9662), .B(p_input[21304]), .Z(o[1304]) );
  AND U19324 ( .A(p_input[1304]), .B(p_input[11304]), .Z(n9662) );
  AND U19325 ( .A(n9663), .B(p_input[21303]), .Z(o[1303]) );
  AND U19326 ( .A(p_input[1303]), .B(p_input[11303]), .Z(n9663) );
  AND U19327 ( .A(n9664), .B(p_input[21302]), .Z(o[1302]) );
  AND U19328 ( .A(p_input[1302]), .B(p_input[11302]), .Z(n9664) );
  AND U19329 ( .A(n9665), .B(p_input[21301]), .Z(o[1301]) );
  AND U19330 ( .A(p_input[1301]), .B(p_input[11301]), .Z(n9665) );
  AND U19331 ( .A(n9666), .B(p_input[21300]), .Z(o[1300]) );
  AND U19332 ( .A(p_input[1300]), .B(p_input[11300]), .Z(n9666) );
  AND U19333 ( .A(n9667), .B(p_input[20012]), .Z(o[12]) );
  AND U19334 ( .A(p_input[12]), .B(p_input[10012]), .Z(n9667) );
  AND U19335 ( .A(n9668), .B(p_input[20129]), .Z(o[129]) );
  AND U19336 ( .A(p_input[129]), .B(p_input[10129]), .Z(n9668) );
  AND U19337 ( .A(n9669), .B(p_input[21299]), .Z(o[1299]) );
  AND U19338 ( .A(p_input[1299]), .B(p_input[11299]), .Z(n9669) );
  AND U19339 ( .A(n9670), .B(p_input[21298]), .Z(o[1298]) );
  AND U19340 ( .A(p_input[1298]), .B(p_input[11298]), .Z(n9670) );
  AND U19341 ( .A(n9671), .B(p_input[21297]), .Z(o[1297]) );
  AND U19342 ( .A(p_input[1297]), .B(p_input[11297]), .Z(n9671) );
  AND U19343 ( .A(n9672), .B(p_input[21296]), .Z(o[1296]) );
  AND U19344 ( .A(p_input[1296]), .B(p_input[11296]), .Z(n9672) );
  AND U19345 ( .A(n9673), .B(p_input[21295]), .Z(o[1295]) );
  AND U19346 ( .A(p_input[1295]), .B(p_input[11295]), .Z(n9673) );
  AND U19347 ( .A(n9674), .B(p_input[21294]), .Z(o[1294]) );
  AND U19348 ( .A(p_input[1294]), .B(p_input[11294]), .Z(n9674) );
  AND U19349 ( .A(n9675), .B(p_input[21293]), .Z(o[1293]) );
  AND U19350 ( .A(p_input[1293]), .B(p_input[11293]), .Z(n9675) );
  AND U19351 ( .A(n9676), .B(p_input[21292]), .Z(o[1292]) );
  AND U19352 ( .A(p_input[1292]), .B(p_input[11292]), .Z(n9676) );
  AND U19353 ( .A(n9677), .B(p_input[21291]), .Z(o[1291]) );
  AND U19354 ( .A(p_input[1291]), .B(p_input[11291]), .Z(n9677) );
  AND U19355 ( .A(n9678), .B(p_input[21290]), .Z(o[1290]) );
  AND U19356 ( .A(p_input[1290]), .B(p_input[11290]), .Z(n9678) );
  AND U19357 ( .A(n9679), .B(p_input[20128]), .Z(o[128]) );
  AND U19358 ( .A(p_input[128]), .B(p_input[10128]), .Z(n9679) );
  AND U19359 ( .A(n9680), .B(p_input[21289]), .Z(o[1289]) );
  AND U19360 ( .A(p_input[1289]), .B(p_input[11289]), .Z(n9680) );
  AND U19361 ( .A(n9681), .B(p_input[21288]), .Z(o[1288]) );
  AND U19362 ( .A(p_input[1288]), .B(p_input[11288]), .Z(n9681) );
  AND U19363 ( .A(n9682), .B(p_input[21287]), .Z(o[1287]) );
  AND U19364 ( .A(p_input[1287]), .B(p_input[11287]), .Z(n9682) );
  AND U19365 ( .A(n9683), .B(p_input[21286]), .Z(o[1286]) );
  AND U19366 ( .A(p_input[1286]), .B(p_input[11286]), .Z(n9683) );
  AND U19367 ( .A(n9684), .B(p_input[21285]), .Z(o[1285]) );
  AND U19368 ( .A(p_input[1285]), .B(p_input[11285]), .Z(n9684) );
  AND U19369 ( .A(n9685), .B(p_input[21284]), .Z(o[1284]) );
  AND U19370 ( .A(p_input[1284]), .B(p_input[11284]), .Z(n9685) );
  AND U19371 ( .A(n9686), .B(p_input[21283]), .Z(o[1283]) );
  AND U19372 ( .A(p_input[1283]), .B(p_input[11283]), .Z(n9686) );
  AND U19373 ( .A(n9687), .B(p_input[21282]), .Z(o[1282]) );
  AND U19374 ( .A(p_input[1282]), .B(p_input[11282]), .Z(n9687) );
  AND U19375 ( .A(n9688), .B(p_input[21281]), .Z(o[1281]) );
  AND U19376 ( .A(p_input[1281]), .B(p_input[11281]), .Z(n9688) );
  AND U19377 ( .A(n9689), .B(p_input[21280]), .Z(o[1280]) );
  AND U19378 ( .A(p_input[1280]), .B(p_input[11280]), .Z(n9689) );
  AND U19379 ( .A(n9690), .B(p_input[20127]), .Z(o[127]) );
  AND U19380 ( .A(p_input[127]), .B(p_input[10127]), .Z(n9690) );
  AND U19381 ( .A(n9691), .B(p_input[21279]), .Z(o[1279]) );
  AND U19382 ( .A(p_input[1279]), .B(p_input[11279]), .Z(n9691) );
  AND U19383 ( .A(n9692), .B(p_input[21278]), .Z(o[1278]) );
  AND U19384 ( .A(p_input[1278]), .B(p_input[11278]), .Z(n9692) );
  AND U19385 ( .A(n9693), .B(p_input[21277]), .Z(o[1277]) );
  AND U19386 ( .A(p_input[1277]), .B(p_input[11277]), .Z(n9693) );
  AND U19387 ( .A(n9694), .B(p_input[21276]), .Z(o[1276]) );
  AND U19388 ( .A(p_input[1276]), .B(p_input[11276]), .Z(n9694) );
  AND U19389 ( .A(n9695), .B(p_input[21275]), .Z(o[1275]) );
  AND U19390 ( .A(p_input[1275]), .B(p_input[11275]), .Z(n9695) );
  AND U19391 ( .A(n9696), .B(p_input[21274]), .Z(o[1274]) );
  AND U19392 ( .A(p_input[1274]), .B(p_input[11274]), .Z(n9696) );
  AND U19393 ( .A(n9697), .B(p_input[21273]), .Z(o[1273]) );
  AND U19394 ( .A(p_input[1273]), .B(p_input[11273]), .Z(n9697) );
  AND U19395 ( .A(n9698), .B(p_input[21272]), .Z(o[1272]) );
  AND U19396 ( .A(p_input[1272]), .B(p_input[11272]), .Z(n9698) );
  AND U19397 ( .A(n9699), .B(p_input[21271]), .Z(o[1271]) );
  AND U19398 ( .A(p_input[1271]), .B(p_input[11271]), .Z(n9699) );
  AND U19399 ( .A(n9700), .B(p_input[21270]), .Z(o[1270]) );
  AND U19400 ( .A(p_input[1270]), .B(p_input[11270]), .Z(n9700) );
  AND U19401 ( .A(n9701), .B(p_input[20126]), .Z(o[126]) );
  AND U19402 ( .A(p_input[126]), .B(p_input[10126]), .Z(n9701) );
  AND U19403 ( .A(n9702), .B(p_input[21269]), .Z(o[1269]) );
  AND U19404 ( .A(p_input[1269]), .B(p_input[11269]), .Z(n9702) );
  AND U19405 ( .A(n9703), .B(p_input[21268]), .Z(o[1268]) );
  AND U19406 ( .A(p_input[1268]), .B(p_input[11268]), .Z(n9703) );
  AND U19407 ( .A(n9704), .B(p_input[21267]), .Z(o[1267]) );
  AND U19408 ( .A(p_input[1267]), .B(p_input[11267]), .Z(n9704) );
  AND U19409 ( .A(n9705), .B(p_input[21266]), .Z(o[1266]) );
  AND U19410 ( .A(p_input[1266]), .B(p_input[11266]), .Z(n9705) );
  AND U19411 ( .A(n9706), .B(p_input[21265]), .Z(o[1265]) );
  AND U19412 ( .A(p_input[1265]), .B(p_input[11265]), .Z(n9706) );
  AND U19413 ( .A(n9707), .B(p_input[21264]), .Z(o[1264]) );
  AND U19414 ( .A(p_input[1264]), .B(p_input[11264]), .Z(n9707) );
  AND U19415 ( .A(n9708), .B(p_input[21263]), .Z(o[1263]) );
  AND U19416 ( .A(p_input[1263]), .B(p_input[11263]), .Z(n9708) );
  AND U19417 ( .A(n9709), .B(p_input[21262]), .Z(o[1262]) );
  AND U19418 ( .A(p_input[1262]), .B(p_input[11262]), .Z(n9709) );
  AND U19419 ( .A(n9710), .B(p_input[21261]), .Z(o[1261]) );
  AND U19420 ( .A(p_input[1261]), .B(p_input[11261]), .Z(n9710) );
  AND U19421 ( .A(n9711), .B(p_input[21260]), .Z(o[1260]) );
  AND U19422 ( .A(p_input[1260]), .B(p_input[11260]), .Z(n9711) );
  AND U19423 ( .A(n9712), .B(p_input[20125]), .Z(o[125]) );
  AND U19424 ( .A(p_input[125]), .B(p_input[10125]), .Z(n9712) );
  AND U19425 ( .A(n9713), .B(p_input[21259]), .Z(o[1259]) );
  AND U19426 ( .A(p_input[1259]), .B(p_input[11259]), .Z(n9713) );
  AND U19427 ( .A(n9714), .B(p_input[21258]), .Z(o[1258]) );
  AND U19428 ( .A(p_input[1258]), .B(p_input[11258]), .Z(n9714) );
  AND U19429 ( .A(n9715), .B(p_input[21257]), .Z(o[1257]) );
  AND U19430 ( .A(p_input[1257]), .B(p_input[11257]), .Z(n9715) );
  AND U19431 ( .A(n9716), .B(p_input[21256]), .Z(o[1256]) );
  AND U19432 ( .A(p_input[1256]), .B(p_input[11256]), .Z(n9716) );
  AND U19433 ( .A(n9717), .B(p_input[21255]), .Z(o[1255]) );
  AND U19434 ( .A(p_input[1255]), .B(p_input[11255]), .Z(n9717) );
  AND U19435 ( .A(n9718), .B(p_input[21254]), .Z(o[1254]) );
  AND U19436 ( .A(p_input[1254]), .B(p_input[11254]), .Z(n9718) );
  AND U19437 ( .A(n9719), .B(p_input[21253]), .Z(o[1253]) );
  AND U19438 ( .A(p_input[1253]), .B(p_input[11253]), .Z(n9719) );
  AND U19439 ( .A(n9720), .B(p_input[21252]), .Z(o[1252]) );
  AND U19440 ( .A(p_input[1252]), .B(p_input[11252]), .Z(n9720) );
  AND U19441 ( .A(n9721), .B(p_input[21251]), .Z(o[1251]) );
  AND U19442 ( .A(p_input[1251]), .B(p_input[11251]), .Z(n9721) );
  AND U19443 ( .A(n9722), .B(p_input[21250]), .Z(o[1250]) );
  AND U19444 ( .A(p_input[1250]), .B(p_input[11250]), .Z(n9722) );
  AND U19445 ( .A(n9723), .B(p_input[20124]), .Z(o[124]) );
  AND U19446 ( .A(p_input[124]), .B(p_input[10124]), .Z(n9723) );
  AND U19447 ( .A(n9724), .B(p_input[21249]), .Z(o[1249]) );
  AND U19448 ( .A(p_input[1249]), .B(p_input[11249]), .Z(n9724) );
  AND U19449 ( .A(n9725), .B(p_input[21248]), .Z(o[1248]) );
  AND U19450 ( .A(p_input[1248]), .B(p_input[11248]), .Z(n9725) );
  AND U19451 ( .A(n9726), .B(p_input[21247]), .Z(o[1247]) );
  AND U19452 ( .A(p_input[1247]), .B(p_input[11247]), .Z(n9726) );
  AND U19453 ( .A(n9727), .B(p_input[21246]), .Z(o[1246]) );
  AND U19454 ( .A(p_input[1246]), .B(p_input[11246]), .Z(n9727) );
  AND U19455 ( .A(n9728), .B(p_input[21245]), .Z(o[1245]) );
  AND U19456 ( .A(p_input[1245]), .B(p_input[11245]), .Z(n9728) );
  AND U19457 ( .A(n9729), .B(p_input[21244]), .Z(o[1244]) );
  AND U19458 ( .A(p_input[1244]), .B(p_input[11244]), .Z(n9729) );
  AND U19459 ( .A(n9730), .B(p_input[21243]), .Z(o[1243]) );
  AND U19460 ( .A(p_input[1243]), .B(p_input[11243]), .Z(n9730) );
  AND U19461 ( .A(n9731), .B(p_input[21242]), .Z(o[1242]) );
  AND U19462 ( .A(p_input[1242]), .B(p_input[11242]), .Z(n9731) );
  AND U19463 ( .A(n9732), .B(p_input[21241]), .Z(o[1241]) );
  AND U19464 ( .A(p_input[1241]), .B(p_input[11241]), .Z(n9732) );
  AND U19465 ( .A(n9733), .B(p_input[21240]), .Z(o[1240]) );
  AND U19466 ( .A(p_input[1240]), .B(p_input[11240]), .Z(n9733) );
  AND U19467 ( .A(n9734), .B(p_input[20123]), .Z(o[123]) );
  AND U19468 ( .A(p_input[123]), .B(p_input[10123]), .Z(n9734) );
  AND U19469 ( .A(n9735), .B(p_input[21239]), .Z(o[1239]) );
  AND U19470 ( .A(p_input[1239]), .B(p_input[11239]), .Z(n9735) );
  AND U19471 ( .A(n9736), .B(p_input[21238]), .Z(o[1238]) );
  AND U19472 ( .A(p_input[1238]), .B(p_input[11238]), .Z(n9736) );
  AND U19473 ( .A(n9737), .B(p_input[21237]), .Z(o[1237]) );
  AND U19474 ( .A(p_input[1237]), .B(p_input[11237]), .Z(n9737) );
  AND U19475 ( .A(n9738), .B(p_input[21236]), .Z(o[1236]) );
  AND U19476 ( .A(p_input[1236]), .B(p_input[11236]), .Z(n9738) );
  AND U19477 ( .A(n9739), .B(p_input[21235]), .Z(o[1235]) );
  AND U19478 ( .A(p_input[1235]), .B(p_input[11235]), .Z(n9739) );
  AND U19479 ( .A(n9740), .B(p_input[21234]), .Z(o[1234]) );
  AND U19480 ( .A(p_input[1234]), .B(p_input[11234]), .Z(n9740) );
  AND U19481 ( .A(n9741), .B(p_input[21233]), .Z(o[1233]) );
  AND U19482 ( .A(p_input[1233]), .B(p_input[11233]), .Z(n9741) );
  AND U19483 ( .A(n9742), .B(p_input[21232]), .Z(o[1232]) );
  AND U19484 ( .A(p_input[1232]), .B(p_input[11232]), .Z(n9742) );
  AND U19485 ( .A(n9743), .B(p_input[21231]), .Z(o[1231]) );
  AND U19486 ( .A(p_input[1231]), .B(p_input[11231]), .Z(n9743) );
  AND U19487 ( .A(n9744), .B(p_input[21230]), .Z(o[1230]) );
  AND U19488 ( .A(p_input[1230]), .B(p_input[11230]), .Z(n9744) );
  AND U19489 ( .A(n9745), .B(p_input[20122]), .Z(o[122]) );
  AND U19490 ( .A(p_input[122]), .B(p_input[10122]), .Z(n9745) );
  AND U19491 ( .A(n9746), .B(p_input[21229]), .Z(o[1229]) );
  AND U19492 ( .A(p_input[1229]), .B(p_input[11229]), .Z(n9746) );
  AND U19493 ( .A(n9747), .B(p_input[21228]), .Z(o[1228]) );
  AND U19494 ( .A(p_input[1228]), .B(p_input[11228]), .Z(n9747) );
  AND U19495 ( .A(n9748), .B(p_input[21227]), .Z(o[1227]) );
  AND U19496 ( .A(p_input[1227]), .B(p_input[11227]), .Z(n9748) );
  AND U19497 ( .A(n9749), .B(p_input[21226]), .Z(o[1226]) );
  AND U19498 ( .A(p_input[1226]), .B(p_input[11226]), .Z(n9749) );
  AND U19499 ( .A(n9750), .B(p_input[21225]), .Z(o[1225]) );
  AND U19500 ( .A(p_input[1225]), .B(p_input[11225]), .Z(n9750) );
  AND U19501 ( .A(n9751), .B(p_input[21224]), .Z(o[1224]) );
  AND U19502 ( .A(p_input[1224]), .B(p_input[11224]), .Z(n9751) );
  AND U19503 ( .A(n9752), .B(p_input[21223]), .Z(o[1223]) );
  AND U19504 ( .A(p_input[1223]), .B(p_input[11223]), .Z(n9752) );
  AND U19505 ( .A(n9753), .B(p_input[21222]), .Z(o[1222]) );
  AND U19506 ( .A(p_input[1222]), .B(p_input[11222]), .Z(n9753) );
  AND U19507 ( .A(n9754), .B(p_input[21221]), .Z(o[1221]) );
  AND U19508 ( .A(p_input[1221]), .B(p_input[11221]), .Z(n9754) );
  AND U19509 ( .A(n9755), .B(p_input[21220]), .Z(o[1220]) );
  AND U19510 ( .A(p_input[1220]), .B(p_input[11220]), .Z(n9755) );
  AND U19511 ( .A(n9756), .B(p_input[20121]), .Z(o[121]) );
  AND U19512 ( .A(p_input[121]), .B(p_input[10121]), .Z(n9756) );
  AND U19513 ( .A(n9757), .B(p_input[21219]), .Z(o[1219]) );
  AND U19514 ( .A(p_input[1219]), .B(p_input[11219]), .Z(n9757) );
  AND U19515 ( .A(n9758), .B(p_input[21218]), .Z(o[1218]) );
  AND U19516 ( .A(p_input[1218]), .B(p_input[11218]), .Z(n9758) );
  AND U19517 ( .A(n9759), .B(p_input[21217]), .Z(o[1217]) );
  AND U19518 ( .A(p_input[1217]), .B(p_input[11217]), .Z(n9759) );
  AND U19519 ( .A(n9760), .B(p_input[21216]), .Z(o[1216]) );
  AND U19520 ( .A(p_input[1216]), .B(p_input[11216]), .Z(n9760) );
  AND U19521 ( .A(n9761), .B(p_input[21215]), .Z(o[1215]) );
  AND U19522 ( .A(p_input[1215]), .B(p_input[11215]), .Z(n9761) );
  AND U19523 ( .A(n9762), .B(p_input[21214]), .Z(o[1214]) );
  AND U19524 ( .A(p_input[1214]), .B(p_input[11214]), .Z(n9762) );
  AND U19525 ( .A(n9763), .B(p_input[21213]), .Z(o[1213]) );
  AND U19526 ( .A(p_input[1213]), .B(p_input[11213]), .Z(n9763) );
  AND U19527 ( .A(n9764), .B(p_input[21212]), .Z(o[1212]) );
  AND U19528 ( .A(p_input[1212]), .B(p_input[11212]), .Z(n9764) );
  AND U19529 ( .A(n9765), .B(p_input[21211]), .Z(o[1211]) );
  AND U19530 ( .A(p_input[1211]), .B(p_input[11211]), .Z(n9765) );
  AND U19531 ( .A(n9766), .B(p_input[21210]), .Z(o[1210]) );
  AND U19532 ( .A(p_input[1210]), .B(p_input[11210]), .Z(n9766) );
  AND U19533 ( .A(n9767), .B(p_input[20120]), .Z(o[120]) );
  AND U19534 ( .A(p_input[120]), .B(p_input[10120]), .Z(n9767) );
  AND U19535 ( .A(n9768), .B(p_input[21209]), .Z(o[1209]) );
  AND U19536 ( .A(p_input[1209]), .B(p_input[11209]), .Z(n9768) );
  AND U19537 ( .A(n9769), .B(p_input[21208]), .Z(o[1208]) );
  AND U19538 ( .A(p_input[1208]), .B(p_input[11208]), .Z(n9769) );
  AND U19539 ( .A(n9770), .B(p_input[21207]), .Z(o[1207]) );
  AND U19540 ( .A(p_input[1207]), .B(p_input[11207]), .Z(n9770) );
  AND U19541 ( .A(n9771), .B(p_input[21206]), .Z(o[1206]) );
  AND U19542 ( .A(p_input[1206]), .B(p_input[11206]), .Z(n9771) );
  AND U19543 ( .A(n9772), .B(p_input[21205]), .Z(o[1205]) );
  AND U19544 ( .A(p_input[1205]), .B(p_input[11205]), .Z(n9772) );
  AND U19545 ( .A(n9773), .B(p_input[21204]), .Z(o[1204]) );
  AND U19546 ( .A(p_input[1204]), .B(p_input[11204]), .Z(n9773) );
  AND U19547 ( .A(n9774), .B(p_input[21203]), .Z(o[1203]) );
  AND U19548 ( .A(p_input[1203]), .B(p_input[11203]), .Z(n9774) );
  AND U19549 ( .A(n9775), .B(p_input[21202]), .Z(o[1202]) );
  AND U19550 ( .A(p_input[1202]), .B(p_input[11202]), .Z(n9775) );
  AND U19551 ( .A(n9776), .B(p_input[21201]), .Z(o[1201]) );
  AND U19552 ( .A(p_input[1201]), .B(p_input[11201]), .Z(n9776) );
  AND U19553 ( .A(n9777), .B(p_input[21200]), .Z(o[1200]) );
  AND U19554 ( .A(p_input[1200]), .B(p_input[11200]), .Z(n9777) );
  AND U19555 ( .A(n9778), .B(p_input[20011]), .Z(o[11]) );
  AND U19556 ( .A(p_input[11]), .B(p_input[10011]), .Z(n9778) );
  AND U19557 ( .A(n9779), .B(p_input[20119]), .Z(o[119]) );
  AND U19558 ( .A(p_input[119]), .B(p_input[10119]), .Z(n9779) );
  AND U19559 ( .A(n9780), .B(p_input[21199]), .Z(o[1199]) );
  AND U19560 ( .A(p_input[1199]), .B(p_input[11199]), .Z(n9780) );
  AND U19561 ( .A(n9781), .B(p_input[21198]), .Z(o[1198]) );
  AND U19562 ( .A(p_input[1198]), .B(p_input[11198]), .Z(n9781) );
  AND U19563 ( .A(n9782), .B(p_input[21197]), .Z(o[1197]) );
  AND U19564 ( .A(p_input[1197]), .B(p_input[11197]), .Z(n9782) );
  AND U19565 ( .A(n9783), .B(p_input[21196]), .Z(o[1196]) );
  AND U19566 ( .A(p_input[1196]), .B(p_input[11196]), .Z(n9783) );
  AND U19567 ( .A(n9784), .B(p_input[21195]), .Z(o[1195]) );
  AND U19568 ( .A(p_input[1195]), .B(p_input[11195]), .Z(n9784) );
  AND U19569 ( .A(n9785), .B(p_input[21194]), .Z(o[1194]) );
  AND U19570 ( .A(p_input[1194]), .B(p_input[11194]), .Z(n9785) );
  AND U19571 ( .A(n9786), .B(p_input[21193]), .Z(o[1193]) );
  AND U19572 ( .A(p_input[1193]), .B(p_input[11193]), .Z(n9786) );
  AND U19573 ( .A(n9787), .B(p_input[21192]), .Z(o[1192]) );
  AND U19574 ( .A(p_input[1192]), .B(p_input[11192]), .Z(n9787) );
  AND U19575 ( .A(n9788), .B(p_input[21191]), .Z(o[1191]) );
  AND U19576 ( .A(p_input[1191]), .B(p_input[11191]), .Z(n9788) );
  AND U19577 ( .A(n9789), .B(p_input[21190]), .Z(o[1190]) );
  AND U19578 ( .A(p_input[1190]), .B(p_input[11190]), .Z(n9789) );
  AND U19579 ( .A(n9790), .B(p_input[20118]), .Z(o[118]) );
  AND U19580 ( .A(p_input[118]), .B(p_input[10118]), .Z(n9790) );
  AND U19581 ( .A(n9791), .B(p_input[21189]), .Z(o[1189]) );
  AND U19582 ( .A(p_input[1189]), .B(p_input[11189]), .Z(n9791) );
  AND U19583 ( .A(n9792), .B(p_input[21188]), .Z(o[1188]) );
  AND U19584 ( .A(p_input[1188]), .B(p_input[11188]), .Z(n9792) );
  AND U19585 ( .A(n9793), .B(p_input[21187]), .Z(o[1187]) );
  AND U19586 ( .A(p_input[1187]), .B(p_input[11187]), .Z(n9793) );
  AND U19587 ( .A(n9794), .B(p_input[21186]), .Z(o[1186]) );
  AND U19588 ( .A(p_input[1186]), .B(p_input[11186]), .Z(n9794) );
  AND U19589 ( .A(n9795), .B(p_input[21185]), .Z(o[1185]) );
  AND U19590 ( .A(p_input[1185]), .B(p_input[11185]), .Z(n9795) );
  AND U19591 ( .A(n9796), .B(p_input[21184]), .Z(o[1184]) );
  AND U19592 ( .A(p_input[1184]), .B(p_input[11184]), .Z(n9796) );
  AND U19593 ( .A(n9797), .B(p_input[21183]), .Z(o[1183]) );
  AND U19594 ( .A(p_input[1183]), .B(p_input[11183]), .Z(n9797) );
  AND U19595 ( .A(n9798), .B(p_input[21182]), .Z(o[1182]) );
  AND U19596 ( .A(p_input[1182]), .B(p_input[11182]), .Z(n9798) );
  AND U19597 ( .A(n9799), .B(p_input[21181]), .Z(o[1181]) );
  AND U19598 ( .A(p_input[1181]), .B(p_input[11181]), .Z(n9799) );
  AND U19599 ( .A(n9800), .B(p_input[21180]), .Z(o[1180]) );
  AND U19600 ( .A(p_input[1180]), .B(p_input[11180]), .Z(n9800) );
  AND U19601 ( .A(n9801), .B(p_input[20117]), .Z(o[117]) );
  AND U19602 ( .A(p_input[117]), .B(p_input[10117]), .Z(n9801) );
  AND U19603 ( .A(n9802), .B(p_input[21179]), .Z(o[1179]) );
  AND U19604 ( .A(p_input[1179]), .B(p_input[11179]), .Z(n9802) );
  AND U19605 ( .A(n9803), .B(p_input[21178]), .Z(o[1178]) );
  AND U19606 ( .A(p_input[1178]), .B(p_input[11178]), .Z(n9803) );
  AND U19607 ( .A(n9804), .B(p_input[21177]), .Z(o[1177]) );
  AND U19608 ( .A(p_input[1177]), .B(p_input[11177]), .Z(n9804) );
  AND U19609 ( .A(n9805), .B(p_input[21176]), .Z(o[1176]) );
  AND U19610 ( .A(p_input[1176]), .B(p_input[11176]), .Z(n9805) );
  AND U19611 ( .A(n9806), .B(p_input[21175]), .Z(o[1175]) );
  AND U19612 ( .A(p_input[1175]), .B(p_input[11175]), .Z(n9806) );
  AND U19613 ( .A(n9807), .B(p_input[21174]), .Z(o[1174]) );
  AND U19614 ( .A(p_input[1174]), .B(p_input[11174]), .Z(n9807) );
  AND U19615 ( .A(n9808), .B(p_input[21173]), .Z(o[1173]) );
  AND U19616 ( .A(p_input[1173]), .B(p_input[11173]), .Z(n9808) );
  AND U19617 ( .A(n9809), .B(p_input[21172]), .Z(o[1172]) );
  AND U19618 ( .A(p_input[1172]), .B(p_input[11172]), .Z(n9809) );
  AND U19619 ( .A(n9810), .B(p_input[21171]), .Z(o[1171]) );
  AND U19620 ( .A(p_input[1171]), .B(p_input[11171]), .Z(n9810) );
  AND U19621 ( .A(n9811), .B(p_input[21170]), .Z(o[1170]) );
  AND U19622 ( .A(p_input[1170]), .B(p_input[11170]), .Z(n9811) );
  AND U19623 ( .A(n9812), .B(p_input[20116]), .Z(o[116]) );
  AND U19624 ( .A(p_input[116]), .B(p_input[10116]), .Z(n9812) );
  AND U19625 ( .A(n9813), .B(p_input[21169]), .Z(o[1169]) );
  AND U19626 ( .A(p_input[1169]), .B(p_input[11169]), .Z(n9813) );
  AND U19627 ( .A(n9814), .B(p_input[21168]), .Z(o[1168]) );
  AND U19628 ( .A(p_input[1168]), .B(p_input[11168]), .Z(n9814) );
  AND U19629 ( .A(n9815), .B(p_input[21167]), .Z(o[1167]) );
  AND U19630 ( .A(p_input[1167]), .B(p_input[11167]), .Z(n9815) );
  AND U19631 ( .A(n9816), .B(p_input[21166]), .Z(o[1166]) );
  AND U19632 ( .A(p_input[1166]), .B(p_input[11166]), .Z(n9816) );
  AND U19633 ( .A(n9817), .B(p_input[21165]), .Z(o[1165]) );
  AND U19634 ( .A(p_input[1165]), .B(p_input[11165]), .Z(n9817) );
  AND U19635 ( .A(n9818), .B(p_input[21164]), .Z(o[1164]) );
  AND U19636 ( .A(p_input[1164]), .B(p_input[11164]), .Z(n9818) );
  AND U19637 ( .A(n9819), .B(p_input[21163]), .Z(o[1163]) );
  AND U19638 ( .A(p_input[1163]), .B(p_input[11163]), .Z(n9819) );
  AND U19639 ( .A(n9820), .B(p_input[21162]), .Z(o[1162]) );
  AND U19640 ( .A(p_input[1162]), .B(p_input[11162]), .Z(n9820) );
  AND U19641 ( .A(n9821), .B(p_input[21161]), .Z(o[1161]) );
  AND U19642 ( .A(p_input[1161]), .B(p_input[11161]), .Z(n9821) );
  AND U19643 ( .A(n9822), .B(p_input[21160]), .Z(o[1160]) );
  AND U19644 ( .A(p_input[1160]), .B(p_input[11160]), .Z(n9822) );
  AND U19645 ( .A(n9823), .B(p_input[20115]), .Z(o[115]) );
  AND U19646 ( .A(p_input[115]), .B(p_input[10115]), .Z(n9823) );
  AND U19647 ( .A(n9824), .B(p_input[21159]), .Z(o[1159]) );
  AND U19648 ( .A(p_input[1159]), .B(p_input[11159]), .Z(n9824) );
  AND U19649 ( .A(n9825), .B(p_input[21158]), .Z(o[1158]) );
  AND U19650 ( .A(p_input[1158]), .B(p_input[11158]), .Z(n9825) );
  AND U19651 ( .A(n9826), .B(p_input[21157]), .Z(o[1157]) );
  AND U19652 ( .A(p_input[1157]), .B(p_input[11157]), .Z(n9826) );
  AND U19653 ( .A(n9827), .B(p_input[21156]), .Z(o[1156]) );
  AND U19654 ( .A(p_input[1156]), .B(p_input[11156]), .Z(n9827) );
  AND U19655 ( .A(n9828), .B(p_input[21155]), .Z(o[1155]) );
  AND U19656 ( .A(p_input[1155]), .B(p_input[11155]), .Z(n9828) );
  AND U19657 ( .A(n9829), .B(p_input[21154]), .Z(o[1154]) );
  AND U19658 ( .A(p_input[1154]), .B(p_input[11154]), .Z(n9829) );
  AND U19659 ( .A(n9830), .B(p_input[21153]), .Z(o[1153]) );
  AND U19660 ( .A(p_input[1153]), .B(p_input[11153]), .Z(n9830) );
  AND U19661 ( .A(n9831), .B(p_input[21152]), .Z(o[1152]) );
  AND U19662 ( .A(p_input[1152]), .B(p_input[11152]), .Z(n9831) );
  AND U19663 ( .A(n9832), .B(p_input[21151]), .Z(o[1151]) );
  AND U19664 ( .A(p_input[1151]), .B(p_input[11151]), .Z(n9832) );
  AND U19665 ( .A(n9833), .B(p_input[21150]), .Z(o[1150]) );
  AND U19666 ( .A(p_input[1150]), .B(p_input[11150]), .Z(n9833) );
  AND U19667 ( .A(n9834), .B(p_input[20114]), .Z(o[114]) );
  AND U19668 ( .A(p_input[114]), .B(p_input[10114]), .Z(n9834) );
  AND U19669 ( .A(n9835), .B(p_input[21149]), .Z(o[1149]) );
  AND U19670 ( .A(p_input[1149]), .B(p_input[11149]), .Z(n9835) );
  AND U19671 ( .A(n9836), .B(p_input[21148]), .Z(o[1148]) );
  AND U19672 ( .A(p_input[1148]), .B(p_input[11148]), .Z(n9836) );
  AND U19673 ( .A(n9837), .B(p_input[21147]), .Z(o[1147]) );
  AND U19674 ( .A(p_input[1147]), .B(p_input[11147]), .Z(n9837) );
  AND U19675 ( .A(n9838), .B(p_input[21146]), .Z(o[1146]) );
  AND U19676 ( .A(p_input[1146]), .B(p_input[11146]), .Z(n9838) );
  AND U19677 ( .A(n9839), .B(p_input[21145]), .Z(o[1145]) );
  AND U19678 ( .A(p_input[1145]), .B(p_input[11145]), .Z(n9839) );
  AND U19679 ( .A(n9840), .B(p_input[21144]), .Z(o[1144]) );
  AND U19680 ( .A(p_input[1144]), .B(p_input[11144]), .Z(n9840) );
  AND U19681 ( .A(n9841), .B(p_input[21143]), .Z(o[1143]) );
  AND U19682 ( .A(p_input[1143]), .B(p_input[11143]), .Z(n9841) );
  AND U19683 ( .A(n9842), .B(p_input[21142]), .Z(o[1142]) );
  AND U19684 ( .A(p_input[1142]), .B(p_input[11142]), .Z(n9842) );
  AND U19685 ( .A(n9843), .B(p_input[21141]), .Z(o[1141]) );
  AND U19686 ( .A(p_input[1141]), .B(p_input[11141]), .Z(n9843) );
  AND U19687 ( .A(n9844), .B(p_input[21140]), .Z(o[1140]) );
  AND U19688 ( .A(p_input[1140]), .B(p_input[11140]), .Z(n9844) );
  AND U19689 ( .A(n9845), .B(p_input[20113]), .Z(o[113]) );
  AND U19690 ( .A(p_input[113]), .B(p_input[10113]), .Z(n9845) );
  AND U19691 ( .A(n9846), .B(p_input[21139]), .Z(o[1139]) );
  AND U19692 ( .A(p_input[1139]), .B(p_input[11139]), .Z(n9846) );
  AND U19693 ( .A(n9847), .B(p_input[21138]), .Z(o[1138]) );
  AND U19694 ( .A(p_input[1138]), .B(p_input[11138]), .Z(n9847) );
  AND U19695 ( .A(n9848), .B(p_input[21137]), .Z(o[1137]) );
  AND U19696 ( .A(p_input[1137]), .B(p_input[11137]), .Z(n9848) );
  AND U19697 ( .A(n9849), .B(p_input[21136]), .Z(o[1136]) );
  AND U19698 ( .A(p_input[1136]), .B(p_input[11136]), .Z(n9849) );
  AND U19699 ( .A(n9850), .B(p_input[21135]), .Z(o[1135]) );
  AND U19700 ( .A(p_input[1135]), .B(p_input[11135]), .Z(n9850) );
  AND U19701 ( .A(n9851), .B(p_input[21134]), .Z(o[1134]) );
  AND U19702 ( .A(p_input[1134]), .B(p_input[11134]), .Z(n9851) );
  AND U19703 ( .A(n9852), .B(p_input[21133]), .Z(o[1133]) );
  AND U19704 ( .A(p_input[1133]), .B(p_input[11133]), .Z(n9852) );
  AND U19705 ( .A(n9853), .B(p_input[21132]), .Z(o[1132]) );
  AND U19706 ( .A(p_input[1132]), .B(p_input[11132]), .Z(n9853) );
  AND U19707 ( .A(n9854), .B(p_input[21131]), .Z(o[1131]) );
  AND U19708 ( .A(p_input[1131]), .B(p_input[11131]), .Z(n9854) );
  AND U19709 ( .A(n9855), .B(p_input[21130]), .Z(o[1130]) );
  AND U19710 ( .A(p_input[1130]), .B(p_input[11130]), .Z(n9855) );
  AND U19711 ( .A(n9856), .B(p_input[20112]), .Z(o[112]) );
  AND U19712 ( .A(p_input[112]), .B(p_input[10112]), .Z(n9856) );
  AND U19713 ( .A(n9857), .B(p_input[21129]), .Z(o[1129]) );
  AND U19714 ( .A(p_input[1129]), .B(p_input[11129]), .Z(n9857) );
  AND U19715 ( .A(n9858), .B(p_input[21128]), .Z(o[1128]) );
  AND U19716 ( .A(p_input[1128]), .B(p_input[11128]), .Z(n9858) );
  AND U19717 ( .A(n9859), .B(p_input[21127]), .Z(o[1127]) );
  AND U19718 ( .A(p_input[1127]), .B(p_input[11127]), .Z(n9859) );
  AND U19719 ( .A(n9860), .B(p_input[21126]), .Z(o[1126]) );
  AND U19720 ( .A(p_input[1126]), .B(p_input[11126]), .Z(n9860) );
  AND U19721 ( .A(n9861), .B(p_input[21125]), .Z(o[1125]) );
  AND U19722 ( .A(p_input[1125]), .B(p_input[11125]), .Z(n9861) );
  AND U19723 ( .A(n9862), .B(p_input[21124]), .Z(o[1124]) );
  AND U19724 ( .A(p_input[1124]), .B(p_input[11124]), .Z(n9862) );
  AND U19725 ( .A(n9863), .B(p_input[21123]), .Z(o[1123]) );
  AND U19726 ( .A(p_input[1123]), .B(p_input[11123]), .Z(n9863) );
  AND U19727 ( .A(n9864), .B(p_input[21122]), .Z(o[1122]) );
  AND U19728 ( .A(p_input[1122]), .B(p_input[11122]), .Z(n9864) );
  AND U19729 ( .A(n9865), .B(p_input[21121]), .Z(o[1121]) );
  AND U19730 ( .A(p_input[1121]), .B(p_input[11121]), .Z(n9865) );
  AND U19731 ( .A(n9866), .B(p_input[21120]), .Z(o[1120]) );
  AND U19732 ( .A(p_input[1120]), .B(p_input[11120]), .Z(n9866) );
  AND U19733 ( .A(n9867), .B(p_input[20111]), .Z(o[111]) );
  AND U19734 ( .A(p_input[111]), .B(p_input[10111]), .Z(n9867) );
  AND U19735 ( .A(n9868), .B(p_input[21119]), .Z(o[1119]) );
  AND U19736 ( .A(p_input[1119]), .B(p_input[11119]), .Z(n9868) );
  AND U19737 ( .A(n9869), .B(p_input[21118]), .Z(o[1118]) );
  AND U19738 ( .A(p_input[1118]), .B(p_input[11118]), .Z(n9869) );
  AND U19739 ( .A(n9870), .B(p_input[21117]), .Z(o[1117]) );
  AND U19740 ( .A(p_input[1117]), .B(p_input[11117]), .Z(n9870) );
  AND U19741 ( .A(n9871), .B(p_input[21116]), .Z(o[1116]) );
  AND U19742 ( .A(p_input[1116]), .B(p_input[11116]), .Z(n9871) );
  AND U19743 ( .A(n9872), .B(p_input[21115]), .Z(o[1115]) );
  AND U19744 ( .A(p_input[1115]), .B(p_input[11115]), .Z(n9872) );
  AND U19745 ( .A(n9873), .B(p_input[21114]), .Z(o[1114]) );
  AND U19746 ( .A(p_input[1114]), .B(p_input[11114]), .Z(n9873) );
  AND U19747 ( .A(n9874), .B(p_input[21113]), .Z(o[1113]) );
  AND U19748 ( .A(p_input[1113]), .B(p_input[11113]), .Z(n9874) );
  AND U19749 ( .A(n9875), .B(p_input[21112]), .Z(o[1112]) );
  AND U19750 ( .A(p_input[1112]), .B(p_input[11112]), .Z(n9875) );
  AND U19751 ( .A(n9876), .B(p_input[21111]), .Z(o[1111]) );
  AND U19752 ( .A(p_input[1111]), .B(p_input[11111]), .Z(n9876) );
  AND U19753 ( .A(n9877), .B(p_input[21110]), .Z(o[1110]) );
  AND U19754 ( .A(p_input[11110]), .B(p_input[1110]), .Z(n9877) );
  AND U19755 ( .A(n9878), .B(p_input[20110]), .Z(o[110]) );
  AND U19756 ( .A(p_input[110]), .B(p_input[10110]), .Z(n9878) );
  AND U19757 ( .A(n9879), .B(p_input[21109]), .Z(o[1109]) );
  AND U19758 ( .A(p_input[11109]), .B(p_input[1109]), .Z(n9879) );
  AND U19759 ( .A(n9880), .B(p_input[21108]), .Z(o[1108]) );
  AND U19760 ( .A(p_input[11108]), .B(p_input[1108]), .Z(n9880) );
  AND U19761 ( .A(n9881), .B(p_input[21107]), .Z(o[1107]) );
  AND U19762 ( .A(p_input[11107]), .B(p_input[1107]), .Z(n9881) );
  AND U19763 ( .A(n9882), .B(p_input[21106]), .Z(o[1106]) );
  AND U19764 ( .A(p_input[11106]), .B(p_input[1106]), .Z(n9882) );
  AND U19765 ( .A(n9883), .B(p_input[21105]), .Z(o[1105]) );
  AND U19766 ( .A(p_input[11105]), .B(p_input[1105]), .Z(n9883) );
  AND U19767 ( .A(n9884), .B(p_input[21104]), .Z(o[1104]) );
  AND U19768 ( .A(p_input[11104]), .B(p_input[1104]), .Z(n9884) );
  AND U19769 ( .A(n9885), .B(p_input[21103]), .Z(o[1103]) );
  AND U19770 ( .A(p_input[11103]), .B(p_input[1103]), .Z(n9885) );
  AND U19771 ( .A(n9886), .B(p_input[21102]), .Z(o[1102]) );
  AND U19772 ( .A(p_input[11102]), .B(p_input[1102]), .Z(n9886) );
  AND U19773 ( .A(n9887), .B(p_input[21101]), .Z(o[1101]) );
  AND U19774 ( .A(p_input[11101]), .B(p_input[1101]), .Z(n9887) );
  AND U19775 ( .A(n9888), .B(p_input[21100]), .Z(o[1100]) );
  AND U19776 ( .A(p_input[11100]), .B(p_input[1100]), .Z(n9888) );
  AND U19777 ( .A(n9889), .B(p_input[20010]), .Z(o[10]) );
  AND U19778 ( .A(p_input[10]), .B(p_input[10010]), .Z(n9889) );
  AND U19779 ( .A(n9890), .B(p_input[20109]), .Z(o[109]) );
  AND U19780 ( .A(p_input[109]), .B(p_input[10109]), .Z(n9890) );
  AND U19781 ( .A(n9891), .B(p_input[21099]), .Z(o[1099]) );
  AND U19782 ( .A(p_input[11099]), .B(p_input[1099]), .Z(n9891) );
  AND U19783 ( .A(n9892), .B(p_input[21098]), .Z(o[1098]) );
  AND U19784 ( .A(p_input[11098]), .B(p_input[1098]), .Z(n9892) );
  AND U19785 ( .A(n9893), .B(p_input[21097]), .Z(o[1097]) );
  AND U19786 ( .A(p_input[11097]), .B(p_input[1097]), .Z(n9893) );
  AND U19787 ( .A(n9894), .B(p_input[21096]), .Z(o[1096]) );
  AND U19788 ( .A(p_input[11096]), .B(p_input[1096]), .Z(n9894) );
  AND U19789 ( .A(n9895), .B(p_input[21095]), .Z(o[1095]) );
  AND U19790 ( .A(p_input[11095]), .B(p_input[1095]), .Z(n9895) );
  AND U19791 ( .A(n9896), .B(p_input[21094]), .Z(o[1094]) );
  AND U19792 ( .A(p_input[11094]), .B(p_input[1094]), .Z(n9896) );
  AND U19793 ( .A(n9897), .B(p_input[21093]), .Z(o[1093]) );
  AND U19794 ( .A(p_input[11093]), .B(p_input[1093]), .Z(n9897) );
  AND U19795 ( .A(n9898), .B(p_input[21092]), .Z(o[1092]) );
  AND U19796 ( .A(p_input[11092]), .B(p_input[1092]), .Z(n9898) );
  AND U19797 ( .A(n9899), .B(p_input[21091]), .Z(o[1091]) );
  AND U19798 ( .A(p_input[11091]), .B(p_input[1091]), .Z(n9899) );
  AND U19799 ( .A(n9900), .B(p_input[21090]), .Z(o[1090]) );
  AND U19800 ( .A(p_input[11090]), .B(p_input[1090]), .Z(n9900) );
  AND U19801 ( .A(n9901), .B(p_input[20108]), .Z(o[108]) );
  AND U19802 ( .A(p_input[108]), .B(p_input[10108]), .Z(n9901) );
  AND U19803 ( .A(n9902), .B(p_input[21089]), .Z(o[1089]) );
  AND U19804 ( .A(p_input[11089]), .B(p_input[1089]), .Z(n9902) );
  AND U19805 ( .A(n9903), .B(p_input[21088]), .Z(o[1088]) );
  AND U19806 ( .A(p_input[11088]), .B(p_input[1088]), .Z(n9903) );
  AND U19807 ( .A(n9904), .B(p_input[21087]), .Z(o[1087]) );
  AND U19808 ( .A(p_input[11087]), .B(p_input[1087]), .Z(n9904) );
  AND U19809 ( .A(n9905), .B(p_input[21086]), .Z(o[1086]) );
  AND U19810 ( .A(p_input[11086]), .B(p_input[1086]), .Z(n9905) );
  AND U19811 ( .A(n9906), .B(p_input[21085]), .Z(o[1085]) );
  AND U19812 ( .A(p_input[11085]), .B(p_input[1085]), .Z(n9906) );
  AND U19813 ( .A(n9907), .B(p_input[21084]), .Z(o[1084]) );
  AND U19814 ( .A(p_input[11084]), .B(p_input[1084]), .Z(n9907) );
  AND U19815 ( .A(n9908), .B(p_input[21083]), .Z(o[1083]) );
  AND U19816 ( .A(p_input[11083]), .B(p_input[1083]), .Z(n9908) );
  AND U19817 ( .A(n9909), .B(p_input[21082]), .Z(o[1082]) );
  AND U19818 ( .A(p_input[11082]), .B(p_input[1082]), .Z(n9909) );
  AND U19819 ( .A(n9910), .B(p_input[21081]), .Z(o[1081]) );
  AND U19820 ( .A(p_input[11081]), .B(p_input[1081]), .Z(n9910) );
  AND U19821 ( .A(n9911), .B(p_input[21080]), .Z(o[1080]) );
  AND U19822 ( .A(p_input[11080]), .B(p_input[1080]), .Z(n9911) );
  AND U19823 ( .A(n9912), .B(p_input[20107]), .Z(o[107]) );
  AND U19824 ( .A(p_input[107]), .B(p_input[10107]), .Z(n9912) );
  AND U19825 ( .A(n9913), .B(p_input[21079]), .Z(o[1079]) );
  AND U19826 ( .A(p_input[11079]), .B(p_input[1079]), .Z(n9913) );
  AND U19827 ( .A(n9914), .B(p_input[21078]), .Z(o[1078]) );
  AND U19828 ( .A(p_input[11078]), .B(p_input[1078]), .Z(n9914) );
  AND U19829 ( .A(n9915), .B(p_input[21077]), .Z(o[1077]) );
  AND U19830 ( .A(p_input[11077]), .B(p_input[1077]), .Z(n9915) );
  AND U19831 ( .A(n9916), .B(p_input[21076]), .Z(o[1076]) );
  AND U19832 ( .A(p_input[11076]), .B(p_input[1076]), .Z(n9916) );
  AND U19833 ( .A(n9917), .B(p_input[21075]), .Z(o[1075]) );
  AND U19834 ( .A(p_input[11075]), .B(p_input[1075]), .Z(n9917) );
  AND U19835 ( .A(n9918), .B(p_input[21074]), .Z(o[1074]) );
  AND U19836 ( .A(p_input[11074]), .B(p_input[1074]), .Z(n9918) );
  AND U19837 ( .A(n9919), .B(p_input[21073]), .Z(o[1073]) );
  AND U19838 ( .A(p_input[11073]), .B(p_input[1073]), .Z(n9919) );
  AND U19839 ( .A(n9920), .B(p_input[21072]), .Z(o[1072]) );
  AND U19840 ( .A(p_input[11072]), .B(p_input[1072]), .Z(n9920) );
  AND U19841 ( .A(n9921), .B(p_input[21071]), .Z(o[1071]) );
  AND U19842 ( .A(p_input[11071]), .B(p_input[1071]), .Z(n9921) );
  AND U19843 ( .A(n9922), .B(p_input[21070]), .Z(o[1070]) );
  AND U19844 ( .A(p_input[11070]), .B(p_input[1070]), .Z(n9922) );
  AND U19845 ( .A(n9923), .B(p_input[20106]), .Z(o[106]) );
  AND U19846 ( .A(p_input[106]), .B(p_input[10106]), .Z(n9923) );
  AND U19847 ( .A(n9924), .B(p_input[21069]), .Z(o[1069]) );
  AND U19848 ( .A(p_input[11069]), .B(p_input[1069]), .Z(n9924) );
  AND U19849 ( .A(n9925), .B(p_input[21068]), .Z(o[1068]) );
  AND U19850 ( .A(p_input[11068]), .B(p_input[1068]), .Z(n9925) );
  AND U19851 ( .A(n9926), .B(p_input[21067]), .Z(o[1067]) );
  AND U19852 ( .A(p_input[11067]), .B(p_input[1067]), .Z(n9926) );
  AND U19853 ( .A(n9927), .B(p_input[21066]), .Z(o[1066]) );
  AND U19854 ( .A(p_input[11066]), .B(p_input[1066]), .Z(n9927) );
  AND U19855 ( .A(n9928), .B(p_input[21065]), .Z(o[1065]) );
  AND U19856 ( .A(p_input[11065]), .B(p_input[1065]), .Z(n9928) );
  AND U19857 ( .A(n9929), .B(p_input[21064]), .Z(o[1064]) );
  AND U19858 ( .A(p_input[11064]), .B(p_input[1064]), .Z(n9929) );
  AND U19859 ( .A(n9930), .B(p_input[21063]), .Z(o[1063]) );
  AND U19860 ( .A(p_input[11063]), .B(p_input[1063]), .Z(n9930) );
  AND U19861 ( .A(n9931), .B(p_input[21062]), .Z(o[1062]) );
  AND U19862 ( .A(p_input[11062]), .B(p_input[1062]), .Z(n9931) );
  AND U19863 ( .A(n9932), .B(p_input[21061]), .Z(o[1061]) );
  AND U19864 ( .A(p_input[11061]), .B(p_input[1061]), .Z(n9932) );
  AND U19865 ( .A(n9933), .B(p_input[21060]), .Z(o[1060]) );
  AND U19866 ( .A(p_input[11060]), .B(p_input[1060]), .Z(n9933) );
  AND U19867 ( .A(n9934), .B(p_input[20105]), .Z(o[105]) );
  AND U19868 ( .A(p_input[105]), .B(p_input[10105]), .Z(n9934) );
  AND U19869 ( .A(n9935), .B(p_input[21059]), .Z(o[1059]) );
  AND U19870 ( .A(p_input[11059]), .B(p_input[1059]), .Z(n9935) );
  AND U19871 ( .A(n9936), .B(p_input[21058]), .Z(o[1058]) );
  AND U19872 ( .A(p_input[11058]), .B(p_input[1058]), .Z(n9936) );
  AND U19873 ( .A(n9937), .B(p_input[21057]), .Z(o[1057]) );
  AND U19874 ( .A(p_input[11057]), .B(p_input[1057]), .Z(n9937) );
  AND U19875 ( .A(n9938), .B(p_input[21056]), .Z(o[1056]) );
  AND U19876 ( .A(p_input[11056]), .B(p_input[1056]), .Z(n9938) );
  AND U19877 ( .A(n9939), .B(p_input[21055]), .Z(o[1055]) );
  AND U19878 ( .A(p_input[11055]), .B(p_input[1055]), .Z(n9939) );
  AND U19879 ( .A(n9940), .B(p_input[21054]), .Z(o[1054]) );
  AND U19880 ( .A(p_input[11054]), .B(p_input[1054]), .Z(n9940) );
  AND U19881 ( .A(n9941), .B(p_input[21053]), .Z(o[1053]) );
  AND U19882 ( .A(p_input[11053]), .B(p_input[1053]), .Z(n9941) );
  AND U19883 ( .A(n9942), .B(p_input[21052]), .Z(o[1052]) );
  AND U19884 ( .A(p_input[11052]), .B(p_input[1052]), .Z(n9942) );
  AND U19885 ( .A(n9943), .B(p_input[21051]), .Z(o[1051]) );
  AND U19886 ( .A(p_input[11051]), .B(p_input[1051]), .Z(n9943) );
  AND U19887 ( .A(n9944), .B(p_input[21050]), .Z(o[1050]) );
  AND U19888 ( .A(p_input[11050]), .B(p_input[1050]), .Z(n9944) );
  AND U19889 ( .A(n9945), .B(p_input[20104]), .Z(o[104]) );
  AND U19890 ( .A(p_input[104]), .B(p_input[10104]), .Z(n9945) );
  AND U19891 ( .A(n9946), .B(p_input[21049]), .Z(o[1049]) );
  AND U19892 ( .A(p_input[11049]), .B(p_input[1049]), .Z(n9946) );
  AND U19893 ( .A(n9947), .B(p_input[21048]), .Z(o[1048]) );
  AND U19894 ( .A(p_input[11048]), .B(p_input[1048]), .Z(n9947) );
  AND U19895 ( .A(n9948), .B(p_input[21047]), .Z(o[1047]) );
  AND U19896 ( .A(p_input[11047]), .B(p_input[1047]), .Z(n9948) );
  AND U19897 ( .A(n9949), .B(p_input[21046]), .Z(o[1046]) );
  AND U19898 ( .A(p_input[11046]), .B(p_input[1046]), .Z(n9949) );
  AND U19899 ( .A(n9950), .B(p_input[21045]), .Z(o[1045]) );
  AND U19900 ( .A(p_input[11045]), .B(p_input[1045]), .Z(n9950) );
  AND U19901 ( .A(n9951), .B(p_input[21044]), .Z(o[1044]) );
  AND U19902 ( .A(p_input[11044]), .B(p_input[1044]), .Z(n9951) );
  AND U19903 ( .A(n9952), .B(p_input[21043]), .Z(o[1043]) );
  AND U19904 ( .A(p_input[11043]), .B(p_input[1043]), .Z(n9952) );
  AND U19905 ( .A(n9953), .B(p_input[21042]), .Z(o[1042]) );
  AND U19906 ( .A(p_input[11042]), .B(p_input[1042]), .Z(n9953) );
  AND U19907 ( .A(n9954), .B(p_input[21041]), .Z(o[1041]) );
  AND U19908 ( .A(p_input[11041]), .B(p_input[1041]), .Z(n9954) );
  AND U19909 ( .A(n9955), .B(p_input[21040]), .Z(o[1040]) );
  AND U19910 ( .A(p_input[11040]), .B(p_input[1040]), .Z(n9955) );
  AND U19911 ( .A(n9956), .B(p_input[20103]), .Z(o[103]) );
  AND U19912 ( .A(p_input[103]), .B(p_input[10103]), .Z(n9956) );
  AND U19913 ( .A(n9957), .B(p_input[21039]), .Z(o[1039]) );
  AND U19914 ( .A(p_input[11039]), .B(p_input[1039]), .Z(n9957) );
  AND U19915 ( .A(n9958), .B(p_input[21038]), .Z(o[1038]) );
  AND U19916 ( .A(p_input[11038]), .B(p_input[1038]), .Z(n9958) );
  AND U19917 ( .A(n9959), .B(p_input[21037]), .Z(o[1037]) );
  AND U19918 ( .A(p_input[11037]), .B(p_input[1037]), .Z(n9959) );
  AND U19919 ( .A(n9960), .B(p_input[21036]), .Z(o[1036]) );
  AND U19920 ( .A(p_input[11036]), .B(p_input[1036]), .Z(n9960) );
  AND U19921 ( .A(n9961), .B(p_input[21035]), .Z(o[1035]) );
  AND U19922 ( .A(p_input[11035]), .B(p_input[1035]), .Z(n9961) );
  AND U19923 ( .A(n9962), .B(p_input[21034]), .Z(o[1034]) );
  AND U19924 ( .A(p_input[11034]), .B(p_input[1034]), .Z(n9962) );
  AND U19925 ( .A(n9963), .B(p_input[21033]), .Z(o[1033]) );
  AND U19926 ( .A(p_input[11033]), .B(p_input[1033]), .Z(n9963) );
  AND U19927 ( .A(n9964), .B(p_input[21032]), .Z(o[1032]) );
  AND U19928 ( .A(p_input[11032]), .B(p_input[1032]), .Z(n9964) );
  AND U19929 ( .A(n9965), .B(p_input[21031]), .Z(o[1031]) );
  AND U19930 ( .A(p_input[11031]), .B(p_input[1031]), .Z(n9965) );
  AND U19931 ( .A(n9966), .B(p_input[21030]), .Z(o[1030]) );
  AND U19932 ( .A(p_input[11030]), .B(p_input[1030]), .Z(n9966) );
  AND U19933 ( .A(n9967), .B(p_input[20102]), .Z(o[102]) );
  AND U19934 ( .A(p_input[102]), .B(p_input[10102]), .Z(n9967) );
  AND U19935 ( .A(n9968), .B(p_input[21029]), .Z(o[1029]) );
  AND U19936 ( .A(p_input[11029]), .B(p_input[1029]), .Z(n9968) );
  AND U19937 ( .A(n9969), .B(p_input[21028]), .Z(o[1028]) );
  AND U19938 ( .A(p_input[11028]), .B(p_input[1028]), .Z(n9969) );
  AND U19939 ( .A(n9970), .B(p_input[21027]), .Z(o[1027]) );
  AND U19940 ( .A(p_input[11027]), .B(p_input[1027]), .Z(n9970) );
  AND U19941 ( .A(n9971), .B(p_input[21026]), .Z(o[1026]) );
  AND U19942 ( .A(p_input[11026]), .B(p_input[1026]), .Z(n9971) );
  AND U19943 ( .A(n9972), .B(p_input[21025]), .Z(o[1025]) );
  AND U19944 ( .A(p_input[11025]), .B(p_input[1025]), .Z(n9972) );
  AND U19945 ( .A(n9973), .B(p_input[21024]), .Z(o[1024]) );
  AND U19946 ( .A(p_input[11024]), .B(p_input[1024]), .Z(n9973) );
  AND U19947 ( .A(n9974), .B(p_input[21023]), .Z(o[1023]) );
  AND U19948 ( .A(p_input[11023]), .B(p_input[1023]), .Z(n9974) );
  AND U19949 ( .A(n9975), .B(p_input[21022]), .Z(o[1022]) );
  AND U19950 ( .A(p_input[11022]), .B(p_input[1022]), .Z(n9975) );
  AND U19951 ( .A(n9976), .B(p_input[21021]), .Z(o[1021]) );
  AND U19952 ( .A(p_input[11021]), .B(p_input[1021]), .Z(n9976) );
  AND U19953 ( .A(n9977), .B(p_input[21020]), .Z(o[1020]) );
  AND U19954 ( .A(p_input[11020]), .B(p_input[1020]), .Z(n9977) );
  AND U19955 ( .A(n9978), .B(p_input[20101]), .Z(o[101]) );
  AND U19956 ( .A(p_input[101]), .B(p_input[10101]), .Z(n9978) );
  AND U19957 ( .A(n9979), .B(p_input[21019]), .Z(o[1019]) );
  AND U19958 ( .A(p_input[11019]), .B(p_input[1019]), .Z(n9979) );
  AND U19959 ( .A(n9980), .B(p_input[21018]), .Z(o[1018]) );
  AND U19960 ( .A(p_input[11018]), .B(p_input[1018]), .Z(n9980) );
  AND U19961 ( .A(n9981), .B(p_input[21017]), .Z(o[1017]) );
  AND U19962 ( .A(p_input[11017]), .B(p_input[1017]), .Z(n9981) );
  AND U19963 ( .A(n9982), .B(p_input[21016]), .Z(o[1016]) );
  AND U19964 ( .A(p_input[11016]), .B(p_input[1016]), .Z(n9982) );
  AND U19965 ( .A(n9983), .B(p_input[21015]), .Z(o[1015]) );
  AND U19966 ( .A(p_input[11015]), .B(p_input[1015]), .Z(n9983) );
  AND U19967 ( .A(n9984), .B(p_input[21014]), .Z(o[1014]) );
  AND U19968 ( .A(p_input[11014]), .B(p_input[1014]), .Z(n9984) );
  AND U19969 ( .A(n9985), .B(p_input[21013]), .Z(o[1013]) );
  AND U19970 ( .A(p_input[11013]), .B(p_input[1013]), .Z(n9985) );
  AND U19971 ( .A(n9986), .B(p_input[21012]), .Z(o[1012]) );
  AND U19972 ( .A(p_input[11012]), .B(p_input[1012]), .Z(n9986) );
  AND U19973 ( .A(n9987), .B(p_input[21011]), .Z(o[1011]) );
  AND U19974 ( .A(p_input[11011]), .B(p_input[1011]), .Z(n9987) );
  AND U19975 ( .A(n9988), .B(p_input[21010]), .Z(o[1010]) );
  AND U19976 ( .A(p_input[11010]), .B(p_input[1010]), .Z(n9988) );
  AND U19977 ( .A(n9989), .B(p_input[20100]), .Z(o[100]) );
  AND U19978 ( .A(p_input[10100]), .B(p_input[100]), .Z(n9989) );
  AND U19979 ( .A(n9990), .B(p_input[21009]), .Z(o[1009]) );
  AND U19980 ( .A(p_input[11009]), .B(p_input[1009]), .Z(n9990) );
  AND U19981 ( .A(n9991), .B(p_input[21008]), .Z(o[1008]) );
  AND U19982 ( .A(p_input[11008]), .B(p_input[1008]), .Z(n9991) );
  AND U19983 ( .A(n9992), .B(p_input[21007]), .Z(o[1007]) );
  AND U19984 ( .A(p_input[11007]), .B(p_input[1007]), .Z(n9992) );
  AND U19985 ( .A(n9993), .B(p_input[21006]), .Z(o[1006]) );
  AND U19986 ( .A(p_input[11006]), .B(p_input[1006]), .Z(n9993) );
  AND U19987 ( .A(n9994), .B(p_input[21005]), .Z(o[1005]) );
  AND U19988 ( .A(p_input[11005]), .B(p_input[1005]), .Z(n9994) );
  AND U19989 ( .A(n9995), .B(p_input[21004]), .Z(o[1004]) );
  AND U19990 ( .A(p_input[11004]), .B(p_input[1004]), .Z(n9995) );
  AND U19991 ( .A(n9996), .B(p_input[21003]), .Z(o[1003]) );
  AND U19992 ( .A(p_input[11003]), .B(p_input[1003]), .Z(n9996) );
  AND U19993 ( .A(n9997), .B(p_input[21002]), .Z(o[1002]) );
  AND U19994 ( .A(p_input[11002]), .B(p_input[1002]), .Z(n9997) );
  AND U19995 ( .A(n9998), .B(p_input[21001]), .Z(o[1001]) );
  AND U19996 ( .A(p_input[11001]), .B(p_input[1001]), .Z(n9998) );
  AND U19997 ( .A(n9999), .B(p_input[21000]), .Z(o[1000]) );
  AND U19998 ( .A(p_input[11000]), .B(p_input[1000]), .Z(n9999) );
  AND U19999 ( .A(n10000), .B(p_input[20000]), .Z(o[0]) );
  AND U20000 ( .A(p_input[10000]), .B(p_input[0]), .Z(n10000) );
endmodule

