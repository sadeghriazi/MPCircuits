
module auction_BMR_N4_W32 ( p_input, o );
  input [511:0] p_input;
  output [35:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464;

  XNOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(o[3]), .B(n3), .Z(n1) );
  XOR U3 ( .A(n2), .B(n4), .Z(n3) );
  XOR U4 ( .A(n5), .B(n6), .Z(o[8]) );
  AND U5 ( .A(o[3]), .B(n7), .Z(n5) );
  XOR U6 ( .A(n8), .B(n9), .Z(n7) );
  XOR U7 ( .A(n10), .B(n11), .Z(o[7]) );
  AND U8 ( .A(o[3]), .B(n12), .Z(n10) );
  XOR U9 ( .A(n13), .B(n14), .Z(n12) );
  XOR U10 ( .A(n15), .B(n16), .Z(o[6]) );
  AND U11 ( .A(o[3]), .B(n17), .Z(n15) );
  XOR U12 ( .A(n18), .B(n19), .Z(n17) );
  XOR U13 ( .A(n20), .B(n21), .Z(o[5]) );
  AND U14 ( .A(o[3]), .B(n22), .Z(n20) );
  XOR U15 ( .A(n23), .B(n24), .Z(n22) );
  XNOR U16 ( .A(n25), .B(n26), .Z(o[4]) );
  AND U17 ( .A(o[3]), .B(n27), .Z(n25) );
  XNOR U18 ( .A(n28), .B(n26), .Z(n27) );
  XOR U19 ( .A(n29), .B(n30), .Z(o[35]) );
  AND U20 ( .A(o[3]), .B(n31), .Z(n29) );
  XOR U21 ( .A(n32), .B(n33), .Z(n31) );
  XOR U22 ( .A(n34), .B(n35), .Z(o[34]) );
  AND U23 ( .A(o[3]), .B(n36), .Z(n34) );
  XOR U24 ( .A(n37), .B(n38), .Z(n36) );
  XOR U25 ( .A(n39), .B(n40), .Z(o[33]) );
  AND U26 ( .A(o[3]), .B(n41), .Z(n39) );
  XOR U27 ( .A(n42), .B(n43), .Z(n41) );
  XOR U28 ( .A(n44), .B(n45), .Z(o[32]) );
  AND U29 ( .A(o[3]), .B(n46), .Z(n44) );
  XOR U30 ( .A(n47), .B(n48), .Z(n46) );
  XOR U31 ( .A(n49), .B(n50), .Z(o[31]) );
  AND U32 ( .A(o[3]), .B(n51), .Z(n49) );
  XOR U33 ( .A(n52), .B(n53), .Z(n51) );
  XOR U34 ( .A(n54), .B(n55), .Z(o[30]) );
  AND U35 ( .A(o[3]), .B(n56), .Z(n54) );
  XOR U36 ( .A(n57), .B(n58), .Z(n56) );
  XOR U37 ( .A(n59), .B(n60), .Z(o[29]) );
  AND U38 ( .A(o[3]), .B(n61), .Z(n59) );
  XOR U39 ( .A(n62), .B(n63), .Z(n61) );
  XOR U40 ( .A(n64), .B(n65), .Z(o[28]) );
  AND U41 ( .A(o[3]), .B(n66), .Z(n64) );
  XOR U42 ( .A(n67), .B(n68), .Z(n66) );
  XOR U43 ( .A(n69), .B(n70), .Z(o[27]) );
  AND U44 ( .A(o[3]), .B(n71), .Z(n69) );
  XOR U45 ( .A(n72), .B(n73), .Z(n71) );
  XOR U46 ( .A(n74), .B(n75), .Z(o[26]) );
  AND U47 ( .A(o[3]), .B(n76), .Z(n74) );
  XOR U48 ( .A(n77), .B(n78), .Z(n76) );
  XOR U49 ( .A(n79), .B(n80), .Z(o[25]) );
  AND U50 ( .A(o[3]), .B(n81), .Z(n79) );
  XOR U51 ( .A(n82), .B(n83), .Z(n81) );
  XOR U52 ( .A(n84), .B(n85), .Z(o[24]) );
  AND U53 ( .A(o[3]), .B(n86), .Z(n84) );
  XOR U54 ( .A(n87), .B(n88), .Z(n86) );
  XOR U55 ( .A(n89), .B(n90), .Z(o[23]) );
  AND U56 ( .A(o[3]), .B(n91), .Z(n89) );
  XOR U57 ( .A(n92), .B(n93), .Z(n91) );
  XOR U58 ( .A(n94), .B(n95), .Z(o[22]) );
  AND U59 ( .A(o[3]), .B(n96), .Z(n94) );
  XOR U60 ( .A(n97), .B(n98), .Z(n96) );
  XOR U61 ( .A(n99), .B(n100), .Z(o[21]) );
  AND U62 ( .A(o[3]), .B(n101), .Z(n99) );
  XOR U63 ( .A(n102), .B(n103), .Z(n101) );
  XOR U64 ( .A(n104), .B(n105), .Z(o[20]) );
  AND U65 ( .A(o[3]), .B(n106), .Z(n104) );
  XOR U66 ( .A(n107), .B(n108), .Z(n106) );
  XOR U67 ( .A(n109), .B(n110), .Z(o[19]) );
  AND U68 ( .A(o[3]), .B(n111), .Z(n109) );
  XOR U69 ( .A(n112), .B(n113), .Z(n111) );
  XOR U70 ( .A(n114), .B(n115), .Z(o[18]) );
  AND U71 ( .A(o[3]), .B(n116), .Z(n114) );
  XOR U72 ( .A(n117), .B(n118), .Z(n116) );
  XOR U73 ( .A(n119), .B(n120), .Z(o[17]) );
  AND U74 ( .A(o[3]), .B(n121), .Z(n119) );
  XOR U75 ( .A(n122), .B(n123), .Z(n121) );
  XOR U76 ( .A(n124), .B(n125), .Z(o[16]) );
  AND U77 ( .A(o[3]), .B(n126), .Z(n124) );
  XOR U78 ( .A(n127), .B(n128), .Z(n126) );
  XOR U79 ( .A(n129), .B(n130), .Z(o[15]) );
  AND U80 ( .A(o[3]), .B(n131), .Z(n129) );
  XOR U81 ( .A(n132), .B(n133), .Z(n131) );
  XOR U82 ( .A(n134), .B(n135), .Z(o[14]) );
  AND U83 ( .A(o[3]), .B(n136), .Z(n134) );
  XOR U84 ( .A(n137), .B(n138), .Z(n136) );
  XOR U85 ( .A(n139), .B(n140), .Z(o[13]) );
  AND U86 ( .A(o[3]), .B(n141), .Z(n139) );
  XOR U87 ( .A(n142), .B(n143), .Z(n141) );
  XOR U88 ( .A(n144), .B(n145), .Z(o[12]) );
  AND U89 ( .A(o[3]), .B(n146), .Z(n144) );
  XOR U90 ( .A(n147), .B(n148), .Z(n146) );
  XOR U91 ( .A(n149), .B(n150), .Z(o[11]) );
  AND U92 ( .A(o[3]), .B(n151), .Z(n149) );
  XOR U93 ( .A(n152), .B(n153), .Z(n151) );
  XOR U94 ( .A(n154), .B(n155), .Z(o[10]) );
  AND U95 ( .A(o[3]), .B(n156), .Z(n154) );
  XOR U96 ( .A(n157), .B(n158), .Z(n156) );
  XOR U97 ( .A(n159), .B(n160), .Z(o[0]) );
  AND U98 ( .A(o[1]), .B(n161), .Z(n160) );
  XNOR U99 ( .A(n162), .B(n163), .Z(n161) );
  XNOR U100 ( .A(n164), .B(n159), .Z(n163) );
  AND U101 ( .A(o[2]), .B(n165), .Z(n164) );
  XNOR U102 ( .A(n162), .B(n166), .Z(n165) );
  XNOR U103 ( .A(n167), .B(n168), .Z(n166) );
  AND U104 ( .A(o[3]), .B(n169), .Z(n167) );
  XOR U105 ( .A(n168), .B(n170), .Z(n169) );
  XOR U106 ( .A(n171), .B(n172), .Z(n162) );
  AND U107 ( .A(o[3]), .B(n173), .Z(n172) );
  XOR U108 ( .A(n171), .B(n174), .Z(n173) );
  XOR U109 ( .A(n175), .B(n176), .Z(o[1]) );
  AND U110 ( .A(o[2]), .B(n177), .Z(n176) );
  XNOR U111 ( .A(n175), .B(n178), .Z(n177) );
  XNOR U112 ( .A(n179), .B(n180), .Z(n178) );
  AND U113 ( .A(o[3]), .B(n181), .Z(n179) );
  XOR U114 ( .A(n180), .B(n182), .Z(n181) );
  XOR U115 ( .A(n183), .B(n184), .Z(n175) );
  AND U116 ( .A(o[3]), .B(n185), .Z(n184) );
  XOR U117 ( .A(n183), .B(n186), .Z(n185) );
  XOR U118 ( .A(n187), .B(n188), .Z(n159) );
  AND U119 ( .A(o[2]), .B(n189), .Z(n188) );
  XNOR U120 ( .A(n187), .B(n190), .Z(n189) );
  XNOR U121 ( .A(n191), .B(n192), .Z(n190) );
  AND U122 ( .A(o[3]), .B(n193), .Z(n191) );
  XOR U123 ( .A(n192), .B(n194), .Z(n193) );
  XOR U124 ( .A(n195), .B(n196), .Z(o[2]) );
  AND U125 ( .A(o[3]), .B(n197), .Z(n196) );
  XOR U126 ( .A(n195), .B(n198), .Z(n197) );
  XOR U127 ( .A(n199), .B(n200), .Z(n187) );
  AND U128 ( .A(o[3]), .B(n201), .Z(n200) );
  XOR U129 ( .A(n199), .B(n202), .Z(n201) );
  XOR U130 ( .A(n203), .B(n204), .Z(o[3]) );
  AND U131 ( .A(n205), .B(n206), .Z(n204) );
  XOR U132 ( .A(n203), .B(n32), .Z(n206) );
  XOR U133 ( .A(n207), .B(n208), .Z(n32) );
  AND U134 ( .A(n198), .B(n209), .Z(n208) );
  XOR U135 ( .A(n210), .B(n207), .Z(n209) );
  XNOR U136 ( .A(n33), .B(n203), .Z(n205) );
  IV U137 ( .A(n30), .Z(n33) );
  XNOR U138 ( .A(n211), .B(n212), .Z(n30) );
  AND U139 ( .A(n195), .B(n213), .Z(n212) );
  XOR U140 ( .A(n214), .B(n211), .Z(n213) );
  XOR U141 ( .A(n215), .B(n216), .Z(n203) );
  AND U142 ( .A(n217), .B(n218), .Z(n216) );
  XOR U143 ( .A(n215), .B(n37), .Z(n218) );
  XOR U144 ( .A(n219), .B(n220), .Z(n37) );
  AND U145 ( .A(n198), .B(n221), .Z(n220) );
  XOR U146 ( .A(n222), .B(n219), .Z(n221) );
  XNOR U147 ( .A(n38), .B(n215), .Z(n217) );
  IV U148 ( .A(n35), .Z(n38) );
  XNOR U149 ( .A(n223), .B(n224), .Z(n35) );
  AND U150 ( .A(n195), .B(n225), .Z(n224) );
  XOR U151 ( .A(n226), .B(n223), .Z(n225) );
  XOR U152 ( .A(n227), .B(n228), .Z(n215) );
  AND U153 ( .A(n229), .B(n230), .Z(n228) );
  XOR U154 ( .A(n227), .B(n42), .Z(n230) );
  XOR U155 ( .A(n231), .B(n232), .Z(n42) );
  AND U156 ( .A(n198), .B(n233), .Z(n232) );
  XOR U157 ( .A(n234), .B(n231), .Z(n233) );
  XNOR U158 ( .A(n43), .B(n227), .Z(n229) );
  IV U159 ( .A(n40), .Z(n43) );
  XNOR U160 ( .A(n235), .B(n236), .Z(n40) );
  AND U161 ( .A(n195), .B(n237), .Z(n236) );
  XOR U162 ( .A(n238), .B(n235), .Z(n237) );
  XOR U163 ( .A(n239), .B(n240), .Z(n227) );
  AND U164 ( .A(n241), .B(n242), .Z(n240) );
  XOR U165 ( .A(n239), .B(n47), .Z(n242) );
  XOR U166 ( .A(n243), .B(n244), .Z(n47) );
  AND U167 ( .A(n198), .B(n245), .Z(n244) );
  XOR U168 ( .A(n246), .B(n243), .Z(n245) );
  XNOR U169 ( .A(n48), .B(n239), .Z(n241) );
  IV U170 ( .A(n45), .Z(n48) );
  XNOR U171 ( .A(n247), .B(n248), .Z(n45) );
  AND U172 ( .A(n195), .B(n249), .Z(n248) );
  XOR U173 ( .A(n250), .B(n247), .Z(n249) );
  XOR U174 ( .A(n251), .B(n252), .Z(n239) );
  AND U175 ( .A(n253), .B(n254), .Z(n252) );
  XOR U176 ( .A(n251), .B(n52), .Z(n254) );
  XOR U177 ( .A(n255), .B(n256), .Z(n52) );
  AND U178 ( .A(n198), .B(n257), .Z(n256) );
  XOR U179 ( .A(n258), .B(n255), .Z(n257) );
  XNOR U180 ( .A(n53), .B(n251), .Z(n253) );
  IV U181 ( .A(n50), .Z(n53) );
  XNOR U182 ( .A(n259), .B(n260), .Z(n50) );
  AND U183 ( .A(n195), .B(n261), .Z(n260) );
  XOR U184 ( .A(n262), .B(n259), .Z(n261) );
  XOR U185 ( .A(n263), .B(n264), .Z(n251) );
  AND U186 ( .A(n265), .B(n266), .Z(n264) );
  XOR U187 ( .A(n263), .B(n57), .Z(n266) );
  XOR U188 ( .A(n267), .B(n268), .Z(n57) );
  AND U189 ( .A(n198), .B(n269), .Z(n268) );
  XOR U190 ( .A(n270), .B(n267), .Z(n269) );
  XNOR U191 ( .A(n58), .B(n263), .Z(n265) );
  IV U192 ( .A(n55), .Z(n58) );
  XNOR U193 ( .A(n271), .B(n272), .Z(n55) );
  AND U194 ( .A(n195), .B(n273), .Z(n272) );
  XOR U195 ( .A(n274), .B(n271), .Z(n273) );
  XOR U196 ( .A(n275), .B(n276), .Z(n263) );
  AND U197 ( .A(n277), .B(n278), .Z(n276) );
  XOR U198 ( .A(n275), .B(n62), .Z(n278) );
  XOR U199 ( .A(n279), .B(n280), .Z(n62) );
  AND U200 ( .A(n198), .B(n281), .Z(n280) );
  XOR U201 ( .A(n282), .B(n279), .Z(n281) );
  XNOR U202 ( .A(n63), .B(n275), .Z(n277) );
  IV U203 ( .A(n60), .Z(n63) );
  XNOR U204 ( .A(n283), .B(n284), .Z(n60) );
  AND U205 ( .A(n195), .B(n285), .Z(n284) );
  XOR U206 ( .A(n286), .B(n283), .Z(n285) );
  XOR U207 ( .A(n287), .B(n288), .Z(n275) );
  AND U208 ( .A(n289), .B(n290), .Z(n288) );
  XOR U209 ( .A(n287), .B(n67), .Z(n290) );
  XOR U210 ( .A(n291), .B(n292), .Z(n67) );
  AND U211 ( .A(n198), .B(n293), .Z(n292) );
  XOR U212 ( .A(n294), .B(n291), .Z(n293) );
  XNOR U213 ( .A(n68), .B(n287), .Z(n289) );
  IV U214 ( .A(n65), .Z(n68) );
  XNOR U215 ( .A(n295), .B(n296), .Z(n65) );
  AND U216 ( .A(n195), .B(n297), .Z(n296) );
  XOR U217 ( .A(n298), .B(n295), .Z(n297) );
  XOR U218 ( .A(n299), .B(n300), .Z(n287) );
  AND U219 ( .A(n301), .B(n302), .Z(n300) );
  XOR U220 ( .A(n299), .B(n72), .Z(n302) );
  XOR U221 ( .A(n303), .B(n304), .Z(n72) );
  AND U222 ( .A(n198), .B(n305), .Z(n304) );
  XOR U223 ( .A(n306), .B(n303), .Z(n305) );
  XNOR U224 ( .A(n73), .B(n299), .Z(n301) );
  IV U225 ( .A(n70), .Z(n73) );
  XNOR U226 ( .A(n307), .B(n308), .Z(n70) );
  AND U227 ( .A(n195), .B(n309), .Z(n308) );
  XOR U228 ( .A(n310), .B(n307), .Z(n309) );
  XOR U229 ( .A(n311), .B(n312), .Z(n299) );
  AND U230 ( .A(n313), .B(n314), .Z(n312) );
  XOR U231 ( .A(n311), .B(n77), .Z(n314) );
  XOR U232 ( .A(n315), .B(n316), .Z(n77) );
  AND U233 ( .A(n198), .B(n317), .Z(n316) );
  XOR U234 ( .A(n318), .B(n315), .Z(n317) );
  XNOR U235 ( .A(n78), .B(n311), .Z(n313) );
  IV U236 ( .A(n75), .Z(n78) );
  XNOR U237 ( .A(n319), .B(n320), .Z(n75) );
  AND U238 ( .A(n195), .B(n321), .Z(n320) );
  XOR U239 ( .A(n322), .B(n319), .Z(n321) );
  XOR U240 ( .A(n323), .B(n324), .Z(n311) );
  AND U241 ( .A(n325), .B(n326), .Z(n324) );
  XOR U242 ( .A(n323), .B(n82), .Z(n326) );
  XOR U243 ( .A(n327), .B(n328), .Z(n82) );
  AND U244 ( .A(n198), .B(n329), .Z(n328) );
  XOR U245 ( .A(n330), .B(n327), .Z(n329) );
  XNOR U246 ( .A(n83), .B(n323), .Z(n325) );
  IV U247 ( .A(n80), .Z(n83) );
  XNOR U248 ( .A(n331), .B(n332), .Z(n80) );
  AND U249 ( .A(n195), .B(n333), .Z(n332) );
  XOR U250 ( .A(n334), .B(n331), .Z(n333) );
  XOR U251 ( .A(n335), .B(n336), .Z(n323) );
  AND U252 ( .A(n337), .B(n338), .Z(n336) );
  XOR U253 ( .A(n335), .B(n87), .Z(n338) );
  XOR U254 ( .A(n339), .B(n340), .Z(n87) );
  AND U255 ( .A(n198), .B(n341), .Z(n340) );
  XOR U256 ( .A(n342), .B(n339), .Z(n341) );
  XNOR U257 ( .A(n88), .B(n335), .Z(n337) );
  IV U258 ( .A(n85), .Z(n88) );
  XNOR U259 ( .A(n343), .B(n344), .Z(n85) );
  AND U260 ( .A(n195), .B(n345), .Z(n344) );
  XOR U261 ( .A(n346), .B(n343), .Z(n345) );
  XOR U262 ( .A(n347), .B(n348), .Z(n335) );
  AND U263 ( .A(n349), .B(n350), .Z(n348) );
  XOR U264 ( .A(n347), .B(n92), .Z(n350) );
  XOR U265 ( .A(n351), .B(n352), .Z(n92) );
  AND U266 ( .A(n198), .B(n353), .Z(n352) );
  XOR U267 ( .A(n354), .B(n351), .Z(n353) );
  XNOR U268 ( .A(n93), .B(n347), .Z(n349) );
  IV U269 ( .A(n90), .Z(n93) );
  XNOR U270 ( .A(n355), .B(n356), .Z(n90) );
  AND U271 ( .A(n195), .B(n357), .Z(n356) );
  XOR U272 ( .A(n358), .B(n355), .Z(n357) );
  XOR U273 ( .A(n359), .B(n360), .Z(n347) );
  AND U274 ( .A(n361), .B(n362), .Z(n360) );
  XOR U275 ( .A(n359), .B(n97), .Z(n362) );
  XOR U276 ( .A(n363), .B(n364), .Z(n97) );
  AND U277 ( .A(n198), .B(n365), .Z(n364) );
  XOR U278 ( .A(n366), .B(n363), .Z(n365) );
  XNOR U279 ( .A(n98), .B(n359), .Z(n361) );
  IV U280 ( .A(n95), .Z(n98) );
  XNOR U281 ( .A(n367), .B(n368), .Z(n95) );
  AND U282 ( .A(n195), .B(n369), .Z(n368) );
  XOR U283 ( .A(n370), .B(n367), .Z(n369) );
  XOR U284 ( .A(n371), .B(n372), .Z(n359) );
  AND U285 ( .A(n373), .B(n374), .Z(n372) );
  XOR U286 ( .A(n371), .B(n102), .Z(n374) );
  XOR U287 ( .A(n375), .B(n376), .Z(n102) );
  AND U288 ( .A(n198), .B(n377), .Z(n376) );
  XOR U289 ( .A(n378), .B(n375), .Z(n377) );
  XNOR U290 ( .A(n103), .B(n371), .Z(n373) );
  IV U291 ( .A(n100), .Z(n103) );
  XNOR U292 ( .A(n379), .B(n380), .Z(n100) );
  AND U293 ( .A(n195), .B(n381), .Z(n380) );
  XOR U294 ( .A(n382), .B(n379), .Z(n381) );
  XOR U295 ( .A(n383), .B(n384), .Z(n371) );
  AND U296 ( .A(n385), .B(n386), .Z(n384) );
  XOR U297 ( .A(n383), .B(n107), .Z(n386) );
  XOR U298 ( .A(n387), .B(n388), .Z(n107) );
  AND U299 ( .A(n198), .B(n389), .Z(n388) );
  XOR U300 ( .A(n390), .B(n387), .Z(n389) );
  XNOR U301 ( .A(n108), .B(n383), .Z(n385) );
  IV U302 ( .A(n105), .Z(n108) );
  XNOR U303 ( .A(n391), .B(n392), .Z(n105) );
  AND U304 ( .A(n195), .B(n393), .Z(n392) );
  XOR U305 ( .A(n394), .B(n391), .Z(n393) );
  XOR U306 ( .A(n395), .B(n396), .Z(n383) );
  AND U307 ( .A(n397), .B(n398), .Z(n396) );
  XOR U308 ( .A(n395), .B(n112), .Z(n398) );
  XOR U309 ( .A(n399), .B(n400), .Z(n112) );
  AND U310 ( .A(n198), .B(n401), .Z(n400) );
  XOR U311 ( .A(n402), .B(n399), .Z(n401) );
  XNOR U312 ( .A(n113), .B(n395), .Z(n397) );
  IV U313 ( .A(n110), .Z(n113) );
  XNOR U314 ( .A(n403), .B(n404), .Z(n110) );
  AND U315 ( .A(n195), .B(n405), .Z(n404) );
  XOR U316 ( .A(n406), .B(n403), .Z(n405) );
  XOR U317 ( .A(n407), .B(n408), .Z(n395) );
  AND U318 ( .A(n409), .B(n410), .Z(n408) );
  XOR U319 ( .A(n407), .B(n117), .Z(n410) );
  XOR U320 ( .A(n411), .B(n412), .Z(n117) );
  AND U321 ( .A(n198), .B(n413), .Z(n412) );
  XOR U322 ( .A(n414), .B(n411), .Z(n413) );
  XNOR U323 ( .A(n118), .B(n407), .Z(n409) );
  IV U324 ( .A(n115), .Z(n118) );
  XNOR U325 ( .A(n415), .B(n416), .Z(n115) );
  AND U326 ( .A(n195), .B(n417), .Z(n416) );
  XOR U327 ( .A(n418), .B(n415), .Z(n417) );
  XOR U328 ( .A(n419), .B(n420), .Z(n407) );
  AND U329 ( .A(n421), .B(n422), .Z(n420) );
  XOR U330 ( .A(n419), .B(n122), .Z(n422) );
  XOR U331 ( .A(n423), .B(n424), .Z(n122) );
  AND U332 ( .A(n198), .B(n425), .Z(n424) );
  XOR U333 ( .A(n426), .B(n423), .Z(n425) );
  XNOR U334 ( .A(n123), .B(n419), .Z(n421) );
  IV U335 ( .A(n120), .Z(n123) );
  XNOR U336 ( .A(n427), .B(n428), .Z(n120) );
  AND U337 ( .A(n195), .B(n429), .Z(n428) );
  XOR U338 ( .A(n430), .B(n427), .Z(n429) );
  XOR U339 ( .A(n431), .B(n432), .Z(n419) );
  AND U340 ( .A(n433), .B(n434), .Z(n432) );
  XOR U341 ( .A(n431), .B(n127), .Z(n434) );
  XOR U342 ( .A(n435), .B(n436), .Z(n127) );
  AND U343 ( .A(n198), .B(n437), .Z(n436) );
  XOR U344 ( .A(n438), .B(n435), .Z(n437) );
  XNOR U345 ( .A(n128), .B(n431), .Z(n433) );
  IV U346 ( .A(n125), .Z(n128) );
  XNOR U347 ( .A(n439), .B(n440), .Z(n125) );
  AND U348 ( .A(n195), .B(n441), .Z(n440) );
  XOR U349 ( .A(n442), .B(n439), .Z(n441) );
  XOR U350 ( .A(n443), .B(n444), .Z(n431) );
  AND U351 ( .A(n445), .B(n446), .Z(n444) );
  XOR U352 ( .A(n443), .B(n132), .Z(n446) );
  XOR U353 ( .A(n447), .B(n448), .Z(n132) );
  AND U354 ( .A(n198), .B(n449), .Z(n448) );
  XOR U355 ( .A(n450), .B(n447), .Z(n449) );
  XNOR U356 ( .A(n133), .B(n443), .Z(n445) );
  IV U357 ( .A(n130), .Z(n133) );
  XNOR U358 ( .A(n451), .B(n452), .Z(n130) );
  AND U359 ( .A(n195), .B(n453), .Z(n452) );
  XOR U360 ( .A(n454), .B(n451), .Z(n453) );
  XOR U361 ( .A(n455), .B(n456), .Z(n443) );
  AND U362 ( .A(n457), .B(n458), .Z(n456) );
  XOR U363 ( .A(n455), .B(n137), .Z(n458) );
  XOR U364 ( .A(n459), .B(n460), .Z(n137) );
  AND U365 ( .A(n198), .B(n461), .Z(n460) );
  XOR U366 ( .A(n462), .B(n459), .Z(n461) );
  XNOR U367 ( .A(n138), .B(n455), .Z(n457) );
  IV U368 ( .A(n135), .Z(n138) );
  XNOR U369 ( .A(n463), .B(n464), .Z(n135) );
  AND U370 ( .A(n195), .B(n465), .Z(n464) );
  XOR U371 ( .A(n466), .B(n463), .Z(n465) );
  XOR U372 ( .A(n467), .B(n468), .Z(n455) );
  AND U373 ( .A(n469), .B(n470), .Z(n468) );
  XOR U374 ( .A(n467), .B(n142), .Z(n470) );
  XOR U375 ( .A(n471), .B(n472), .Z(n142) );
  AND U376 ( .A(n198), .B(n473), .Z(n472) );
  XOR U377 ( .A(n474), .B(n471), .Z(n473) );
  XNOR U378 ( .A(n143), .B(n467), .Z(n469) );
  IV U379 ( .A(n140), .Z(n143) );
  XNOR U380 ( .A(n475), .B(n476), .Z(n140) );
  AND U381 ( .A(n195), .B(n477), .Z(n476) );
  XOR U382 ( .A(n478), .B(n475), .Z(n477) );
  XOR U383 ( .A(n479), .B(n480), .Z(n467) );
  AND U384 ( .A(n481), .B(n482), .Z(n480) );
  XOR U385 ( .A(n479), .B(n147), .Z(n482) );
  XOR U386 ( .A(n483), .B(n484), .Z(n147) );
  AND U387 ( .A(n198), .B(n485), .Z(n484) );
  XOR U388 ( .A(n486), .B(n483), .Z(n485) );
  XNOR U389 ( .A(n148), .B(n479), .Z(n481) );
  IV U390 ( .A(n145), .Z(n148) );
  XNOR U391 ( .A(n487), .B(n488), .Z(n145) );
  AND U392 ( .A(n195), .B(n489), .Z(n488) );
  XOR U393 ( .A(n490), .B(n487), .Z(n489) );
  XOR U394 ( .A(n491), .B(n492), .Z(n479) );
  AND U395 ( .A(n493), .B(n494), .Z(n492) );
  XOR U396 ( .A(n491), .B(n152), .Z(n494) );
  XOR U397 ( .A(n495), .B(n496), .Z(n152) );
  AND U398 ( .A(n198), .B(n497), .Z(n496) );
  XOR U399 ( .A(n498), .B(n495), .Z(n497) );
  XNOR U400 ( .A(n153), .B(n491), .Z(n493) );
  IV U401 ( .A(n150), .Z(n153) );
  XNOR U402 ( .A(n499), .B(n500), .Z(n150) );
  AND U403 ( .A(n195), .B(n501), .Z(n500) );
  XOR U404 ( .A(n502), .B(n499), .Z(n501) );
  XOR U405 ( .A(n503), .B(n504), .Z(n491) );
  AND U406 ( .A(n505), .B(n506), .Z(n504) );
  XOR U407 ( .A(n503), .B(n157), .Z(n506) );
  XOR U408 ( .A(n507), .B(n508), .Z(n157) );
  AND U409 ( .A(n198), .B(n509), .Z(n508) );
  XOR U410 ( .A(n510), .B(n507), .Z(n509) );
  XNOR U411 ( .A(n158), .B(n503), .Z(n505) );
  IV U412 ( .A(n155), .Z(n158) );
  XNOR U413 ( .A(n511), .B(n512), .Z(n155) );
  AND U414 ( .A(n195), .B(n513), .Z(n512) );
  XOR U415 ( .A(n514), .B(n511), .Z(n513) );
  XOR U416 ( .A(n515), .B(n516), .Z(n503) );
  AND U417 ( .A(n517), .B(n518), .Z(n516) );
  XOR U418 ( .A(n4), .B(n515), .Z(n518) );
  XOR U419 ( .A(n519), .B(n520), .Z(n4) );
  AND U420 ( .A(n198), .B(n521), .Z(n520) );
  XOR U421 ( .A(n519), .B(n522), .Z(n521) );
  XNOR U422 ( .A(n515), .B(n2), .Z(n517) );
  XOR U423 ( .A(n523), .B(n524), .Z(n2) );
  AND U424 ( .A(n195), .B(n525), .Z(n524) );
  XOR U425 ( .A(n523), .B(n526), .Z(n525) );
  XOR U426 ( .A(n527), .B(n528), .Z(n515) );
  AND U427 ( .A(n529), .B(n530), .Z(n528) );
  XOR U428 ( .A(n527), .B(n8), .Z(n530) );
  XOR U429 ( .A(n531), .B(n532), .Z(n8) );
  AND U430 ( .A(n198), .B(n533), .Z(n532) );
  XOR U431 ( .A(n534), .B(n531), .Z(n533) );
  XNOR U432 ( .A(n9), .B(n527), .Z(n529) );
  IV U433 ( .A(n6), .Z(n9) );
  XNOR U434 ( .A(n535), .B(n536), .Z(n6) );
  AND U435 ( .A(n195), .B(n537), .Z(n536) );
  XOR U436 ( .A(n538), .B(n535), .Z(n537) );
  XOR U437 ( .A(n539), .B(n540), .Z(n527) );
  AND U438 ( .A(n541), .B(n542), .Z(n540) );
  XOR U439 ( .A(n539), .B(n13), .Z(n542) );
  XOR U440 ( .A(n543), .B(n544), .Z(n13) );
  AND U441 ( .A(n198), .B(n545), .Z(n544) );
  XOR U442 ( .A(n546), .B(n543), .Z(n545) );
  XNOR U443 ( .A(n14), .B(n539), .Z(n541) );
  IV U444 ( .A(n11), .Z(n14) );
  XNOR U445 ( .A(n547), .B(n548), .Z(n11) );
  AND U446 ( .A(n195), .B(n549), .Z(n548) );
  XOR U447 ( .A(n550), .B(n547), .Z(n549) );
  XOR U448 ( .A(n551), .B(n552), .Z(n539) );
  AND U449 ( .A(n553), .B(n554), .Z(n552) );
  XOR U450 ( .A(n551), .B(n18), .Z(n554) );
  XOR U451 ( .A(n555), .B(n556), .Z(n18) );
  AND U452 ( .A(n198), .B(n557), .Z(n556) );
  XOR U453 ( .A(n558), .B(n555), .Z(n557) );
  XNOR U454 ( .A(n19), .B(n551), .Z(n553) );
  IV U455 ( .A(n16), .Z(n19) );
  XNOR U456 ( .A(n559), .B(n560), .Z(n16) );
  AND U457 ( .A(n195), .B(n561), .Z(n560) );
  XOR U458 ( .A(n562), .B(n559), .Z(n561) );
  XNOR U459 ( .A(n563), .B(n564), .Z(n551) );
  AND U460 ( .A(n565), .B(n566), .Z(n564) );
  XNOR U461 ( .A(n563), .B(n23), .Z(n566) );
  XOR U462 ( .A(n567), .B(n568), .Z(n23) );
  AND U463 ( .A(n198), .B(n569), .Z(n568) );
  XOR U464 ( .A(n570), .B(n567), .Z(n569) );
  XOR U465 ( .A(n24), .B(n563), .Z(n565) );
  IV U466 ( .A(n21), .Z(n24) );
  XNOR U467 ( .A(n571), .B(n572), .Z(n21) );
  AND U468 ( .A(n195), .B(n573), .Z(n572) );
  XOR U469 ( .A(n574), .B(n571), .Z(n573) );
  AND U470 ( .A(n26), .B(n28), .Z(n563) );
  XNOR U471 ( .A(n575), .B(n576), .Z(n28) );
  AND U472 ( .A(n198), .B(n577), .Z(n576) );
  XNOR U473 ( .A(n578), .B(n575), .Z(n577) );
  XOR U474 ( .A(n579), .B(n580), .Z(n198) );
  AND U475 ( .A(n581), .B(n582), .Z(n580) );
  XOR U476 ( .A(n579), .B(n210), .Z(n582) );
  XNOR U477 ( .A(n583), .B(n584), .Z(n210) );
  AND U478 ( .A(n585), .B(n182), .Z(n584) );
  AND U479 ( .A(n583), .B(n586), .Z(n585) );
  XNOR U480 ( .A(n207), .B(n579), .Z(n581) );
  XOR U481 ( .A(n587), .B(n588), .Z(n207) );
  AND U482 ( .A(n589), .B(n180), .Z(n588) );
  NOR U483 ( .A(n587), .B(n590), .Z(n589) );
  XOR U484 ( .A(n591), .B(n592), .Z(n579) );
  AND U485 ( .A(n593), .B(n594), .Z(n592) );
  XOR U486 ( .A(n591), .B(n222), .Z(n594) );
  XOR U487 ( .A(n595), .B(n596), .Z(n222) );
  AND U488 ( .A(n182), .B(n597), .Z(n596) );
  XOR U489 ( .A(n598), .B(n595), .Z(n597) );
  XNOR U490 ( .A(n219), .B(n591), .Z(n593) );
  XOR U491 ( .A(n599), .B(n600), .Z(n219) );
  AND U492 ( .A(n180), .B(n601), .Z(n600) );
  XOR U493 ( .A(n602), .B(n599), .Z(n601) );
  XOR U494 ( .A(n603), .B(n604), .Z(n591) );
  AND U495 ( .A(n605), .B(n606), .Z(n604) );
  XOR U496 ( .A(n603), .B(n234), .Z(n606) );
  XOR U497 ( .A(n607), .B(n608), .Z(n234) );
  AND U498 ( .A(n182), .B(n609), .Z(n608) );
  XOR U499 ( .A(n610), .B(n607), .Z(n609) );
  XNOR U500 ( .A(n231), .B(n603), .Z(n605) );
  XOR U501 ( .A(n611), .B(n612), .Z(n231) );
  AND U502 ( .A(n180), .B(n613), .Z(n612) );
  XOR U503 ( .A(n614), .B(n611), .Z(n613) );
  XOR U504 ( .A(n615), .B(n616), .Z(n603) );
  AND U505 ( .A(n617), .B(n618), .Z(n616) );
  XOR U506 ( .A(n615), .B(n246), .Z(n618) );
  XOR U507 ( .A(n619), .B(n620), .Z(n246) );
  AND U508 ( .A(n182), .B(n621), .Z(n620) );
  XOR U509 ( .A(n622), .B(n619), .Z(n621) );
  XNOR U510 ( .A(n243), .B(n615), .Z(n617) );
  XOR U511 ( .A(n623), .B(n624), .Z(n243) );
  AND U512 ( .A(n180), .B(n625), .Z(n624) );
  XOR U513 ( .A(n626), .B(n623), .Z(n625) );
  XOR U514 ( .A(n627), .B(n628), .Z(n615) );
  AND U515 ( .A(n629), .B(n630), .Z(n628) );
  XOR U516 ( .A(n627), .B(n258), .Z(n630) );
  XOR U517 ( .A(n631), .B(n632), .Z(n258) );
  AND U518 ( .A(n182), .B(n633), .Z(n632) );
  XOR U519 ( .A(n634), .B(n631), .Z(n633) );
  XNOR U520 ( .A(n255), .B(n627), .Z(n629) );
  XOR U521 ( .A(n635), .B(n636), .Z(n255) );
  AND U522 ( .A(n180), .B(n637), .Z(n636) );
  XOR U523 ( .A(n638), .B(n635), .Z(n637) );
  XOR U524 ( .A(n639), .B(n640), .Z(n627) );
  AND U525 ( .A(n641), .B(n642), .Z(n640) );
  XOR U526 ( .A(n639), .B(n270), .Z(n642) );
  XOR U527 ( .A(n643), .B(n644), .Z(n270) );
  AND U528 ( .A(n182), .B(n645), .Z(n644) );
  XOR U529 ( .A(n646), .B(n643), .Z(n645) );
  XNOR U530 ( .A(n267), .B(n639), .Z(n641) );
  XOR U531 ( .A(n647), .B(n648), .Z(n267) );
  AND U532 ( .A(n180), .B(n649), .Z(n648) );
  XOR U533 ( .A(n650), .B(n647), .Z(n649) );
  XOR U534 ( .A(n651), .B(n652), .Z(n639) );
  AND U535 ( .A(n653), .B(n654), .Z(n652) );
  XOR U536 ( .A(n651), .B(n282), .Z(n654) );
  XOR U537 ( .A(n655), .B(n656), .Z(n282) );
  AND U538 ( .A(n182), .B(n657), .Z(n656) );
  XOR U539 ( .A(n658), .B(n655), .Z(n657) );
  XNOR U540 ( .A(n279), .B(n651), .Z(n653) );
  XOR U541 ( .A(n659), .B(n660), .Z(n279) );
  AND U542 ( .A(n180), .B(n661), .Z(n660) );
  XOR U543 ( .A(n662), .B(n659), .Z(n661) );
  XOR U544 ( .A(n663), .B(n664), .Z(n651) );
  AND U545 ( .A(n665), .B(n666), .Z(n664) );
  XOR U546 ( .A(n663), .B(n294), .Z(n666) );
  XOR U547 ( .A(n667), .B(n668), .Z(n294) );
  AND U548 ( .A(n182), .B(n669), .Z(n668) );
  XOR U549 ( .A(n670), .B(n667), .Z(n669) );
  XNOR U550 ( .A(n291), .B(n663), .Z(n665) );
  XOR U551 ( .A(n671), .B(n672), .Z(n291) );
  AND U552 ( .A(n180), .B(n673), .Z(n672) );
  XOR U553 ( .A(n674), .B(n671), .Z(n673) );
  XOR U554 ( .A(n675), .B(n676), .Z(n663) );
  AND U555 ( .A(n677), .B(n678), .Z(n676) );
  XOR U556 ( .A(n675), .B(n306), .Z(n678) );
  XOR U557 ( .A(n679), .B(n680), .Z(n306) );
  AND U558 ( .A(n182), .B(n681), .Z(n680) );
  XOR U559 ( .A(n682), .B(n679), .Z(n681) );
  XNOR U560 ( .A(n303), .B(n675), .Z(n677) );
  XOR U561 ( .A(n683), .B(n684), .Z(n303) );
  AND U562 ( .A(n180), .B(n685), .Z(n684) );
  XOR U563 ( .A(n686), .B(n683), .Z(n685) );
  XOR U564 ( .A(n687), .B(n688), .Z(n675) );
  AND U565 ( .A(n689), .B(n690), .Z(n688) );
  XOR U566 ( .A(n687), .B(n318), .Z(n690) );
  XOR U567 ( .A(n691), .B(n692), .Z(n318) );
  AND U568 ( .A(n182), .B(n693), .Z(n692) );
  XOR U569 ( .A(n694), .B(n691), .Z(n693) );
  XNOR U570 ( .A(n315), .B(n687), .Z(n689) );
  XOR U571 ( .A(n695), .B(n696), .Z(n315) );
  AND U572 ( .A(n180), .B(n697), .Z(n696) );
  XOR U573 ( .A(n698), .B(n695), .Z(n697) );
  XOR U574 ( .A(n699), .B(n700), .Z(n687) );
  AND U575 ( .A(n701), .B(n702), .Z(n700) );
  XOR U576 ( .A(n699), .B(n330), .Z(n702) );
  XOR U577 ( .A(n703), .B(n704), .Z(n330) );
  AND U578 ( .A(n182), .B(n705), .Z(n704) );
  XOR U579 ( .A(n706), .B(n703), .Z(n705) );
  XNOR U580 ( .A(n327), .B(n699), .Z(n701) );
  XOR U581 ( .A(n707), .B(n708), .Z(n327) );
  AND U582 ( .A(n180), .B(n709), .Z(n708) );
  XOR U583 ( .A(n710), .B(n707), .Z(n709) );
  XOR U584 ( .A(n711), .B(n712), .Z(n699) );
  AND U585 ( .A(n713), .B(n714), .Z(n712) );
  XOR U586 ( .A(n711), .B(n342), .Z(n714) );
  XOR U587 ( .A(n715), .B(n716), .Z(n342) );
  AND U588 ( .A(n182), .B(n717), .Z(n716) );
  XOR U589 ( .A(n718), .B(n715), .Z(n717) );
  XNOR U590 ( .A(n339), .B(n711), .Z(n713) );
  XOR U591 ( .A(n719), .B(n720), .Z(n339) );
  AND U592 ( .A(n180), .B(n721), .Z(n720) );
  XOR U593 ( .A(n722), .B(n719), .Z(n721) );
  XOR U594 ( .A(n723), .B(n724), .Z(n711) );
  AND U595 ( .A(n725), .B(n726), .Z(n724) );
  XOR U596 ( .A(n723), .B(n354), .Z(n726) );
  XOR U597 ( .A(n727), .B(n728), .Z(n354) );
  AND U598 ( .A(n182), .B(n729), .Z(n728) );
  XOR U599 ( .A(n730), .B(n727), .Z(n729) );
  XNOR U600 ( .A(n351), .B(n723), .Z(n725) );
  XOR U601 ( .A(n731), .B(n732), .Z(n351) );
  AND U602 ( .A(n180), .B(n733), .Z(n732) );
  XOR U603 ( .A(n734), .B(n731), .Z(n733) );
  XOR U604 ( .A(n735), .B(n736), .Z(n723) );
  AND U605 ( .A(n737), .B(n738), .Z(n736) );
  XOR U606 ( .A(n735), .B(n366), .Z(n738) );
  XOR U607 ( .A(n739), .B(n740), .Z(n366) );
  AND U608 ( .A(n182), .B(n741), .Z(n740) );
  XOR U609 ( .A(n742), .B(n739), .Z(n741) );
  XNOR U610 ( .A(n363), .B(n735), .Z(n737) );
  XOR U611 ( .A(n743), .B(n744), .Z(n363) );
  AND U612 ( .A(n180), .B(n745), .Z(n744) );
  XOR U613 ( .A(n746), .B(n743), .Z(n745) );
  XOR U614 ( .A(n747), .B(n748), .Z(n735) );
  AND U615 ( .A(n749), .B(n750), .Z(n748) );
  XOR U616 ( .A(n747), .B(n378), .Z(n750) );
  XOR U617 ( .A(n751), .B(n752), .Z(n378) );
  AND U618 ( .A(n182), .B(n753), .Z(n752) );
  XOR U619 ( .A(n754), .B(n751), .Z(n753) );
  XNOR U620 ( .A(n375), .B(n747), .Z(n749) );
  XOR U621 ( .A(n755), .B(n756), .Z(n375) );
  AND U622 ( .A(n180), .B(n757), .Z(n756) );
  XOR U623 ( .A(n758), .B(n755), .Z(n757) );
  XOR U624 ( .A(n759), .B(n760), .Z(n747) );
  AND U625 ( .A(n761), .B(n762), .Z(n760) );
  XOR U626 ( .A(n759), .B(n390), .Z(n762) );
  XOR U627 ( .A(n763), .B(n764), .Z(n390) );
  AND U628 ( .A(n182), .B(n765), .Z(n764) );
  XOR U629 ( .A(n766), .B(n763), .Z(n765) );
  XNOR U630 ( .A(n387), .B(n759), .Z(n761) );
  XOR U631 ( .A(n767), .B(n768), .Z(n387) );
  AND U632 ( .A(n180), .B(n769), .Z(n768) );
  XOR U633 ( .A(n770), .B(n767), .Z(n769) );
  XOR U634 ( .A(n771), .B(n772), .Z(n759) );
  AND U635 ( .A(n773), .B(n774), .Z(n772) );
  XOR U636 ( .A(n771), .B(n402), .Z(n774) );
  XOR U637 ( .A(n775), .B(n776), .Z(n402) );
  AND U638 ( .A(n182), .B(n777), .Z(n776) );
  XOR U639 ( .A(n778), .B(n775), .Z(n777) );
  XNOR U640 ( .A(n399), .B(n771), .Z(n773) );
  XOR U641 ( .A(n779), .B(n780), .Z(n399) );
  AND U642 ( .A(n180), .B(n781), .Z(n780) );
  XOR U643 ( .A(n782), .B(n779), .Z(n781) );
  XOR U644 ( .A(n783), .B(n784), .Z(n771) );
  AND U645 ( .A(n785), .B(n786), .Z(n784) );
  XOR U646 ( .A(n783), .B(n414), .Z(n786) );
  XOR U647 ( .A(n787), .B(n788), .Z(n414) );
  AND U648 ( .A(n182), .B(n789), .Z(n788) );
  XOR U649 ( .A(n790), .B(n787), .Z(n789) );
  XNOR U650 ( .A(n411), .B(n783), .Z(n785) );
  XOR U651 ( .A(n791), .B(n792), .Z(n411) );
  AND U652 ( .A(n180), .B(n793), .Z(n792) );
  XOR U653 ( .A(n794), .B(n791), .Z(n793) );
  XOR U654 ( .A(n795), .B(n796), .Z(n783) );
  AND U655 ( .A(n797), .B(n798), .Z(n796) );
  XOR U656 ( .A(n795), .B(n426), .Z(n798) );
  XOR U657 ( .A(n799), .B(n800), .Z(n426) );
  AND U658 ( .A(n182), .B(n801), .Z(n800) );
  XOR U659 ( .A(n802), .B(n799), .Z(n801) );
  XNOR U660 ( .A(n423), .B(n795), .Z(n797) );
  XOR U661 ( .A(n803), .B(n804), .Z(n423) );
  AND U662 ( .A(n180), .B(n805), .Z(n804) );
  XOR U663 ( .A(n806), .B(n803), .Z(n805) );
  XOR U664 ( .A(n807), .B(n808), .Z(n795) );
  AND U665 ( .A(n809), .B(n810), .Z(n808) );
  XOR U666 ( .A(n807), .B(n438), .Z(n810) );
  XOR U667 ( .A(n811), .B(n812), .Z(n438) );
  AND U668 ( .A(n182), .B(n813), .Z(n812) );
  XOR U669 ( .A(n814), .B(n811), .Z(n813) );
  XNOR U670 ( .A(n435), .B(n807), .Z(n809) );
  XOR U671 ( .A(n815), .B(n816), .Z(n435) );
  AND U672 ( .A(n180), .B(n817), .Z(n816) );
  XOR U673 ( .A(n818), .B(n815), .Z(n817) );
  XOR U674 ( .A(n819), .B(n820), .Z(n807) );
  AND U675 ( .A(n821), .B(n822), .Z(n820) );
  XOR U676 ( .A(n819), .B(n450), .Z(n822) );
  XOR U677 ( .A(n823), .B(n824), .Z(n450) );
  AND U678 ( .A(n182), .B(n825), .Z(n824) );
  XOR U679 ( .A(n826), .B(n823), .Z(n825) );
  XNOR U680 ( .A(n447), .B(n819), .Z(n821) );
  XOR U681 ( .A(n827), .B(n828), .Z(n447) );
  AND U682 ( .A(n180), .B(n829), .Z(n828) );
  XOR U683 ( .A(n830), .B(n827), .Z(n829) );
  XOR U684 ( .A(n831), .B(n832), .Z(n819) );
  AND U685 ( .A(n833), .B(n834), .Z(n832) );
  XOR U686 ( .A(n831), .B(n462), .Z(n834) );
  XOR U687 ( .A(n835), .B(n836), .Z(n462) );
  AND U688 ( .A(n182), .B(n837), .Z(n836) );
  XOR U689 ( .A(n838), .B(n835), .Z(n837) );
  XNOR U690 ( .A(n459), .B(n831), .Z(n833) );
  XOR U691 ( .A(n839), .B(n840), .Z(n459) );
  AND U692 ( .A(n180), .B(n841), .Z(n840) );
  XOR U693 ( .A(n842), .B(n839), .Z(n841) );
  XOR U694 ( .A(n843), .B(n844), .Z(n831) );
  AND U695 ( .A(n845), .B(n846), .Z(n844) );
  XOR U696 ( .A(n843), .B(n474), .Z(n846) );
  XOR U697 ( .A(n847), .B(n848), .Z(n474) );
  AND U698 ( .A(n182), .B(n849), .Z(n848) );
  XOR U699 ( .A(n850), .B(n847), .Z(n849) );
  XNOR U700 ( .A(n471), .B(n843), .Z(n845) );
  XOR U701 ( .A(n851), .B(n852), .Z(n471) );
  AND U702 ( .A(n180), .B(n853), .Z(n852) );
  XOR U703 ( .A(n854), .B(n851), .Z(n853) );
  XOR U704 ( .A(n855), .B(n856), .Z(n843) );
  AND U705 ( .A(n857), .B(n858), .Z(n856) );
  XOR U706 ( .A(n855), .B(n486), .Z(n858) );
  XOR U707 ( .A(n859), .B(n860), .Z(n486) );
  AND U708 ( .A(n182), .B(n861), .Z(n860) );
  XOR U709 ( .A(n862), .B(n859), .Z(n861) );
  XNOR U710 ( .A(n483), .B(n855), .Z(n857) );
  XOR U711 ( .A(n863), .B(n864), .Z(n483) );
  AND U712 ( .A(n180), .B(n865), .Z(n864) );
  XOR U713 ( .A(n866), .B(n863), .Z(n865) );
  XOR U714 ( .A(n867), .B(n868), .Z(n855) );
  AND U715 ( .A(n869), .B(n870), .Z(n868) );
  XOR U716 ( .A(n867), .B(n498), .Z(n870) );
  XOR U717 ( .A(n871), .B(n872), .Z(n498) );
  AND U718 ( .A(n182), .B(n873), .Z(n872) );
  XOR U719 ( .A(n874), .B(n871), .Z(n873) );
  XNOR U720 ( .A(n495), .B(n867), .Z(n869) );
  XOR U721 ( .A(n875), .B(n876), .Z(n495) );
  AND U722 ( .A(n180), .B(n877), .Z(n876) );
  XOR U723 ( .A(n878), .B(n875), .Z(n877) );
  XOR U724 ( .A(n879), .B(n880), .Z(n867) );
  AND U725 ( .A(n881), .B(n882), .Z(n880) );
  XOR U726 ( .A(n879), .B(n510), .Z(n882) );
  XOR U727 ( .A(n883), .B(n884), .Z(n510) );
  AND U728 ( .A(n182), .B(n885), .Z(n884) );
  XOR U729 ( .A(n886), .B(n883), .Z(n885) );
  XNOR U730 ( .A(n507), .B(n879), .Z(n881) );
  XOR U731 ( .A(n887), .B(n888), .Z(n507) );
  AND U732 ( .A(n180), .B(n889), .Z(n888) );
  XOR U733 ( .A(n890), .B(n887), .Z(n889) );
  XOR U734 ( .A(n891), .B(n892), .Z(n879) );
  AND U735 ( .A(n893), .B(n894), .Z(n892) );
  XOR U736 ( .A(n522), .B(n891), .Z(n894) );
  XOR U737 ( .A(n895), .B(n896), .Z(n522) );
  AND U738 ( .A(n182), .B(n897), .Z(n896) );
  XOR U739 ( .A(n895), .B(n898), .Z(n897) );
  XNOR U740 ( .A(n891), .B(n519), .Z(n893) );
  XOR U741 ( .A(n899), .B(n900), .Z(n519) );
  AND U742 ( .A(n180), .B(n901), .Z(n900) );
  XOR U743 ( .A(n899), .B(n902), .Z(n901) );
  XOR U744 ( .A(n903), .B(n904), .Z(n891) );
  AND U745 ( .A(n905), .B(n906), .Z(n904) );
  XOR U746 ( .A(n903), .B(n534), .Z(n906) );
  XOR U747 ( .A(n907), .B(n908), .Z(n534) );
  AND U748 ( .A(n182), .B(n909), .Z(n908) );
  XOR U749 ( .A(n910), .B(n907), .Z(n909) );
  XNOR U750 ( .A(n531), .B(n903), .Z(n905) );
  XOR U751 ( .A(n911), .B(n912), .Z(n531) );
  AND U752 ( .A(n180), .B(n913), .Z(n912) );
  XOR U753 ( .A(n914), .B(n911), .Z(n913) );
  XOR U754 ( .A(n915), .B(n916), .Z(n903) );
  AND U755 ( .A(n917), .B(n918), .Z(n916) );
  XOR U756 ( .A(n915), .B(n546), .Z(n918) );
  XOR U757 ( .A(n919), .B(n920), .Z(n546) );
  AND U758 ( .A(n182), .B(n921), .Z(n920) );
  XOR U759 ( .A(n922), .B(n919), .Z(n921) );
  XNOR U760 ( .A(n543), .B(n915), .Z(n917) );
  XOR U761 ( .A(n923), .B(n924), .Z(n543) );
  AND U762 ( .A(n180), .B(n925), .Z(n924) );
  XOR U763 ( .A(n926), .B(n923), .Z(n925) );
  XOR U764 ( .A(n927), .B(n928), .Z(n915) );
  AND U765 ( .A(n929), .B(n930), .Z(n928) );
  XOR U766 ( .A(n927), .B(n558), .Z(n930) );
  XOR U767 ( .A(n931), .B(n932), .Z(n558) );
  AND U768 ( .A(n182), .B(n933), .Z(n932) );
  XOR U769 ( .A(n934), .B(n931), .Z(n933) );
  XNOR U770 ( .A(n555), .B(n927), .Z(n929) );
  XOR U771 ( .A(n935), .B(n936), .Z(n555) );
  AND U772 ( .A(n180), .B(n937), .Z(n936) );
  XOR U773 ( .A(n938), .B(n935), .Z(n937) );
  XOR U774 ( .A(n939), .B(n940), .Z(n927) );
  AND U775 ( .A(n941), .B(n942), .Z(n940) );
  XNOR U776 ( .A(n943), .B(n570), .Z(n942) );
  XOR U777 ( .A(n944), .B(n945), .Z(n570) );
  AND U778 ( .A(n182), .B(n946), .Z(n945) );
  XOR U779 ( .A(n947), .B(n944), .Z(n946) );
  XNOR U780 ( .A(n567), .B(n939), .Z(n941) );
  XOR U781 ( .A(n948), .B(n949), .Z(n567) );
  AND U782 ( .A(n180), .B(n950), .Z(n949) );
  XOR U783 ( .A(n951), .B(n948), .Z(n950) );
  IV U784 ( .A(n943), .Z(n939) );
  AND U785 ( .A(n575), .B(n578), .Z(n943) );
  XNOR U786 ( .A(n952), .B(n953), .Z(n578) );
  AND U787 ( .A(n182), .B(n954), .Z(n953) );
  XNOR U788 ( .A(n955), .B(n952), .Z(n954) );
  XOR U789 ( .A(n956), .B(n957), .Z(n182) );
  AND U790 ( .A(n958), .B(n959), .Z(n957) );
  XOR U791 ( .A(n586), .B(n956), .Z(n959) );
  IV U792 ( .A(n960), .Z(n586) );
  AND U793 ( .A(p_input[511]), .B(p_input[479]), .Z(n960) );
  XOR U794 ( .A(n956), .B(n583), .Z(n958) );
  AND U795 ( .A(p_input[415]), .B(p_input[447]), .Z(n583) );
  XOR U796 ( .A(n961), .B(n962), .Z(n956) );
  AND U797 ( .A(n963), .B(n964), .Z(n962) );
  XOR U798 ( .A(n961), .B(n598), .Z(n964) );
  XNOR U799 ( .A(p_input[478]), .B(n965), .Z(n598) );
  AND U800 ( .A(n170), .B(n966), .Z(n965) );
  XOR U801 ( .A(p_input[510]), .B(p_input[478]), .Z(n966) );
  XNOR U802 ( .A(n595), .B(n961), .Z(n963) );
  XOR U803 ( .A(n967), .B(n968), .Z(n595) );
  AND U804 ( .A(n168), .B(n969), .Z(n968) );
  XOR U805 ( .A(p_input[446]), .B(p_input[414]), .Z(n969) );
  XOR U806 ( .A(n970), .B(n971), .Z(n961) );
  AND U807 ( .A(n972), .B(n973), .Z(n971) );
  XOR U808 ( .A(n970), .B(n610), .Z(n973) );
  XNOR U809 ( .A(p_input[477]), .B(n974), .Z(n610) );
  AND U810 ( .A(n170), .B(n975), .Z(n974) );
  XOR U811 ( .A(p_input[509]), .B(p_input[477]), .Z(n975) );
  XNOR U812 ( .A(n607), .B(n970), .Z(n972) );
  XOR U813 ( .A(n976), .B(n977), .Z(n607) );
  AND U814 ( .A(n168), .B(n978), .Z(n977) );
  XOR U815 ( .A(p_input[445]), .B(p_input[413]), .Z(n978) );
  XOR U816 ( .A(n979), .B(n980), .Z(n970) );
  AND U817 ( .A(n981), .B(n982), .Z(n980) );
  XOR U818 ( .A(n979), .B(n622), .Z(n982) );
  XNOR U819 ( .A(p_input[476]), .B(n983), .Z(n622) );
  AND U820 ( .A(n170), .B(n984), .Z(n983) );
  XOR U821 ( .A(p_input[508]), .B(p_input[476]), .Z(n984) );
  XNOR U822 ( .A(n619), .B(n979), .Z(n981) );
  XOR U823 ( .A(n985), .B(n986), .Z(n619) );
  AND U824 ( .A(n168), .B(n987), .Z(n986) );
  XOR U825 ( .A(p_input[444]), .B(p_input[412]), .Z(n987) );
  XOR U826 ( .A(n988), .B(n989), .Z(n979) );
  AND U827 ( .A(n990), .B(n991), .Z(n989) );
  XOR U828 ( .A(n988), .B(n634), .Z(n991) );
  XNOR U829 ( .A(p_input[475]), .B(n992), .Z(n634) );
  AND U830 ( .A(n170), .B(n993), .Z(n992) );
  XOR U831 ( .A(p_input[507]), .B(p_input[475]), .Z(n993) );
  XNOR U832 ( .A(n631), .B(n988), .Z(n990) );
  XOR U833 ( .A(n994), .B(n995), .Z(n631) );
  AND U834 ( .A(n168), .B(n996), .Z(n995) );
  XOR U835 ( .A(p_input[443]), .B(p_input[411]), .Z(n996) );
  XOR U836 ( .A(n997), .B(n998), .Z(n988) );
  AND U837 ( .A(n999), .B(n1000), .Z(n998) );
  XOR U838 ( .A(n997), .B(n646), .Z(n1000) );
  XNOR U839 ( .A(p_input[474]), .B(n1001), .Z(n646) );
  AND U840 ( .A(n170), .B(n1002), .Z(n1001) );
  XOR U841 ( .A(p_input[506]), .B(p_input[474]), .Z(n1002) );
  XNOR U842 ( .A(n643), .B(n997), .Z(n999) );
  XOR U843 ( .A(n1003), .B(n1004), .Z(n643) );
  AND U844 ( .A(n168), .B(n1005), .Z(n1004) );
  XOR U845 ( .A(p_input[442]), .B(p_input[410]), .Z(n1005) );
  XOR U846 ( .A(n1006), .B(n1007), .Z(n997) );
  AND U847 ( .A(n1008), .B(n1009), .Z(n1007) );
  XOR U848 ( .A(n1006), .B(n658), .Z(n1009) );
  XNOR U849 ( .A(p_input[473]), .B(n1010), .Z(n658) );
  AND U850 ( .A(n170), .B(n1011), .Z(n1010) );
  XOR U851 ( .A(p_input[505]), .B(p_input[473]), .Z(n1011) );
  XNOR U852 ( .A(n655), .B(n1006), .Z(n1008) );
  XOR U853 ( .A(n1012), .B(n1013), .Z(n655) );
  AND U854 ( .A(n168), .B(n1014), .Z(n1013) );
  XOR U855 ( .A(p_input[441]), .B(p_input[409]), .Z(n1014) );
  XOR U856 ( .A(n1015), .B(n1016), .Z(n1006) );
  AND U857 ( .A(n1017), .B(n1018), .Z(n1016) );
  XOR U858 ( .A(n1015), .B(n670), .Z(n1018) );
  XNOR U859 ( .A(p_input[472]), .B(n1019), .Z(n670) );
  AND U860 ( .A(n170), .B(n1020), .Z(n1019) );
  XOR U861 ( .A(p_input[504]), .B(p_input[472]), .Z(n1020) );
  XNOR U862 ( .A(n667), .B(n1015), .Z(n1017) );
  XOR U863 ( .A(n1021), .B(n1022), .Z(n667) );
  AND U864 ( .A(n168), .B(n1023), .Z(n1022) );
  XOR U865 ( .A(p_input[440]), .B(p_input[408]), .Z(n1023) );
  XOR U866 ( .A(n1024), .B(n1025), .Z(n1015) );
  AND U867 ( .A(n1026), .B(n1027), .Z(n1025) );
  XOR U868 ( .A(n1024), .B(n682), .Z(n1027) );
  XNOR U869 ( .A(p_input[471]), .B(n1028), .Z(n682) );
  AND U870 ( .A(n170), .B(n1029), .Z(n1028) );
  XOR U871 ( .A(p_input[503]), .B(p_input[471]), .Z(n1029) );
  XNOR U872 ( .A(n679), .B(n1024), .Z(n1026) );
  XOR U873 ( .A(n1030), .B(n1031), .Z(n679) );
  AND U874 ( .A(n168), .B(n1032), .Z(n1031) );
  XOR U875 ( .A(p_input[439]), .B(p_input[407]), .Z(n1032) );
  XOR U876 ( .A(n1033), .B(n1034), .Z(n1024) );
  AND U877 ( .A(n1035), .B(n1036), .Z(n1034) );
  XOR U878 ( .A(n1033), .B(n694), .Z(n1036) );
  XNOR U879 ( .A(p_input[470]), .B(n1037), .Z(n694) );
  AND U880 ( .A(n170), .B(n1038), .Z(n1037) );
  XOR U881 ( .A(p_input[502]), .B(p_input[470]), .Z(n1038) );
  XNOR U882 ( .A(n691), .B(n1033), .Z(n1035) );
  XOR U883 ( .A(n1039), .B(n1040), .Z(n691) );
  AND U884 ( .A(n168), .B(n1041), .Z(n1040) );
  XOR U885 ( .A(p_input[438]), .B(p_input[406]), .Z(n1041) );
  XOR U886 ( .A(n1042), .B(n1043), .Z(n1033) );
  AND U887 ( .A(n1044), .B(n1045), .Z(n1043) );
  XOR U888 ( .A(n1042), .B(n706), .Z(n1045) );
  XNOR U889 ( .A(p_input[469]), .B(n1046), .Z(n706) );
  AND U890 ( .A(n170), .B(n1047), .Z(n1046) );
  XOR U891 ( .A(p_input[501]), .B(p_input[469]), .Z(n1047) );
  XNOR U892 ( .A(n703), .B(n1042), .Z(n1044) );
  XOR U893 ( .A(n1048), .B(n1049), .Z(n703) );
  AND U894 ( .A(n168), .B(n1050), .Z(n1049) );
  XOR U895 ( .A(p_input[437]), .B(p_input[405]), .Z(n1050) );
  XOR U896 ( .A(n1051), .B(n1052), .Z(n1042) );
  AND U897 ( .A(n1053), .B(n1054), .Z(n1052) );
  XOR U898 ( .A(n1051), .B(n718), .Z(n1054) );
  XNOR U899 ( .A(p_input[468]), .B(n1055), .Z(n718) );
  AND U900 ( .A(n170), .B(n1056), .Z(n1055) );
  XOR U901 ( .A(p_input[500]), .B(p_input[468]), .Z(n1056) );
  XNOR U902 ( .A(n715), .B(n1051), .Z(n1053) );
  XOR U903 ( .A(n1057), .B(n1058), .Z(n715) );
  AND U904 ( .A(n168), .B(n1059), .Z(n1058) );
  XOR U905 ( .A(p_input[436]), .B(p_input[404]), .Z(n1059) );
  XOR U906 ( .A(n1060), .B(n1061), .Z(n1051) );
  AND U907 ( .A(n1062), .B(n1063), .Z(n1061) );
  XOR U908 ( .A(n1060), .B(n730), .Z(n1063) );
  XNOR U909 ( .A(p_input[467]), .B(n1064), .Z(n730) );
  AND U910 ( .A(n170), .B(n1065), .Z(n1064) );
  XOR U911 ( .A(p_input[499]), .B(p_input[467]), .Z(n1065) );
  XNOR U912 ( .A(n727), .B(n1060), .Z(n1062) );
  XOR U913 ( .A(n1066), .B(n1067), .Z(n727) );
  AND U914 ( .A(n168), .B(n1068), .Z(n1067) );
  XOR U915 ( .A(p_input[435]), .B(p_input[403]), .Z(n1068) );
  XOR U916 ( .A(n1069), .B(n1070), .Z(n1060) );
  AND U917 ( .A(n1071), .B(n1072), .Z(n1070) );
  XOR U918 ( .A(n1069), .B(n742), .Z(n1072) );
  XNOR U919 ( .A(p_input[466]), .B(n1073), .Z(n742) );
  AND U920 ( .A(n170), .B(n1074), .Z(n1073) );
  XOR U921 ( .A(p_input[498]), .B(p_input[466]), .Z(n1074) );
  XNOR U922 ( .A(n739), .B(n1069), .Z(n1071) );
  XOR U923 ( .A(n1075), .B(n1076), .Z(n739) );
  AND U924 ( .A(n168), .B(n1077), .Z(n1076) );
  XOR U925 ( .A(p_input[434]), .B(p_input[402]), .Z(n1077) );
  XOR U926 ( .A(n1078), .B(n1079), .Z(n1069) );
  AND U927 ( .A(n1080), .B(n1081), .Z(n1079) );
  XOR U928 ( .A(n1078), .B(n754), .Z(n1081) );
  XNOR U929 ( .A(p_input[465]), .B(n1082), .Z(n754) );
  AND U930 ( .A(n170), .B(n1083), .Z(n1082) );
  XOR U931 ( .A(p_input[497]), .B(p_input[465]), .Z(n1083) );
  XNOR U932 ( .A(n751), .B(n1078), .Z(n1080) );
  XOR U933 ( .A(n1084), .B(n1085), .Z(n751) );
  AND U934 ( .A(n168), .B(n1086), .Z(n1085) );
  XOR U935 ( .A(p_input[433]), .B(p_input[401]), .Z(n1086) );
  XOR U936 ( .A(n1087), .B(n1088), .Z(n1078) );
  AND U937 ( .A(n1089), .B(n1090), .Z(n1088) );
  XOR U938 ( .A(n1087), .B(n766), .Z(n1090) );
  XNOR U939 ( .A(p_input[464]), .B(n1091), .Z(n766) );
  AND U940 ( .A(n170), .B(n1092), .Z(n1091) );
  XOR U941 ( .A(p_input[496]), .B(p_input[464]), .Z(n1092) );
  XNOR U942 ( .A(n763), .B(n1087), .Z(n1089) );
  XOR U943 ( .A(n1093), .B(n1094), .Z(n763) );
  AND U944 ( .A(n168), .B(n1095), .Z(n1094) );
  XOR U945 ( .A(p_input[432]), .B(p_input[400]), .Z(n1095) );
  XOR U946 ( .A(n1096), .B(n1097), .Z(n1087) );
  AND U947 ( .A(n1098), .B(n1099), .Z(n1097) );
  XOR U948 ( .A(n1096), .B(n778), .Z(n1099) );
  XNOR U949 ( .A(p_input[463]), .B(n1100), .Z(n778) );
  AND U950 ( .A(n170), .B(n1101), .Z(n1100) );
  XOR U951 ( .A(p_input[495]), .B(p_input[463]), .Z(n1101) );
  XNOR U952 ( .A(n775), .B(n1096), .Z(n1098) );
  XOR U953 ( .A(n1102), .B(n1103), .Z(n775) );
  AND U954 ( .A(n168), .B(n1104), .Z(n1103) );
  XOR U955 ( .A(p_input[431]), .B(p_input[399]), .Z(n1104) );
  XOR U956 ( .A(n1105), .B(n1106), .Z(n1096) );
  AND U957 ( .A(n1107), .B(n1108), .Z(n1106) );
  XOR U958 ( .A(n1105), .B(n790), .Z(n1108) );
  XNOR U959 ( .A(p_input[462]), .B(n1109), .Z(n790) );
  AND U960 ( .A(n170), .B(n1110), .Z(n1109) );
  XOR U961 ( .A(p_input[494]), .B(p_input[462]), .Z(n1110) );
  XNOR U962 ( .A(n787), .B(n1105), .Z(n1107) );
  XOR U963 ( .A(n1111), .B(n1112), .Z(n787) );
  AND U964 ( .A(n168), .B(n1113), .Z(n1112) );
  XOR U965 ( .A(p_input[430]), .B(p_input[398]), .Z(n1113) );
  XOR U966 ( .A(n1114), .B(n1115), .Z(n1105) );
  AND U967 ( .A(n1116), .B(n1117), .Z(n1115) );
  XOR U968 ( .A(n1114), .B(n802), .Z(n1117) );
  XNOR U969 ( .A(p_input[461]), .B(n1118), .Z(n802) );
  AND U970 ( .A(n170), .B(n1119), .Z(n1118) );
  XOR U971 ( .A(p_input[493]), .B(p_input[461]), .Z(n1119) );
  XNOR U972 ( .A(n799), .B(n1114), .Z(n1116) );
  XOR U973 ( .A(n1120), .B(n1121), .Z(n799) );
  AND U974 ( .A(n168), .B(n1122), .Z(n1121) );
  XOR U975 ( .A(p_input[429]), .B(p_input[397]), .Z(n1122) );
  XOR U976 ( .A(n1123), .B(n1124), .Z(n1114) );
  AND U977 ( .A(n1125), .B(n1126), .Z(n1124) );
  XOR U978 ( .A(n1123), .B(n814), .Z(n1126) );
  XNOR U979 ( .A(p_input[460]), .B(n1127), .Z(n814) );
  AND U980 ( .A(n170), .B(n1128), .Z(n1127) );
  XOR U981 ( .A(p_input[492]), .B(p_input[460]), .Z(n1128) );
  XNOR U982 ( .A(n811), .B(n1123), .Z(n1125) );
  XOR U983 ( .A(n1129), .B(n1130), .Z(n811) );
  AND U984 ( .A(n168), .B(n1131), .Z(n1130) );
  XOR U985 ( .A(p_input[428]), .B(p_input[396]), .Z(n1131) );
  XOR U986 ( .A(n1132), .B(n1133), .Z(n1123) );
  AND U987 ( .A(n1134), .B(n1135), .Z(n1133) );
  XOR U988 ( .A(n1132), .B(n826), .Z(n1135) );
  XNOR U989 ( .A(p_input[459]), .B(n1136), .Z(n826) );
  AND U990 ( .A(n170), .B(n1137), .Z(n1136) );
  XOR U991 ( .A(p_input[491]), .B(p_input[459]), .Z(n1137) );
  XNOR U992 ( .A(n823), .B(n1132), .Z(n1134) );
  XOR U993 ( .A(n1138), .B(n1139), .Z(n823) );
  AND U994 ( .A(n168), .B(n1140), .Z(n1139) );
  XOR U995 ( .A(p_input[427]), .B(p_input[395]), .Z(n1140) );
  XOR U996 ( .A(n1141), .B(n1142), .Z(n1132) );
  AND U997 ( .A(n1143), .B(n1144), .Z(n1142) );
  XOR U998 ( .A(n1141), .B(n838), .Z(n1144) );
  XNOR U999 ( .A(p_input[458]), .B(n1145), .Z(n838) );
  AND U1000 ( .A(n170), .B(n1146), .Z(n1145) );
  XOR U1001 ( .A(p_input[490]), .B(p_input[458]), .Z(n1146) );
  XNOR U1002 ( .A(n835), .B(n1141), .Z(n1143) );
  XOR U1003 ( .A(n1147), .B(n1148), .Z(n835) );
  AND U1004 ( .A(n168), .B(n1149), .Z(n1148) );
  XOR U1005 ( .A(p_input[426]), .B(p_input[394]), .Z(n1149) );
  XOR U1006 ( .A(n1150), .B(n1151), .Z(n1141) );
  AND U1007 ( .A(n1152), .B(n1153), .Z(n1151) );
  XOR U1008 ( .A(n1150), .B(n850), .Z(n1153) );
  XNOR U1009 ( .A(p_input[457]), .B(n1154), .Z(n850) );
  AND U1010 ( .A(n170), .B(n1155), .Z(n1154) );
  XOR U1011 ( .A(p_input[489]), .B(p_input[457]), .Z(n1155) );
  XNOR U1012 ( .A(n847), .B(n1150), .Z(n1152) );
  XOR U1013 ( .A(n1156), .B(n1157), .Z(n847) );
  AND U1014 ( .A(n168), .B(n1158), .Z(n1157) );
  XOR U1015 ( .A(p_input[425]), .B(p_input[393]), .Z(n1158) );
  XOR U1016 ( .A(n1159), .B(n1160), .Z(n1150) );
  AND U1017 ( .A(n1161), .B(n1162), .Z(n1160) );
  XOR U1018 ( .A(n1159), .B(n862), .Z(n1162) );
  XNOR U1019 ( .A(p_input[456]), .B(n1163), .Z(n862) );
  AND U1020 ( .A(n170), .B(n1164), .Z(n1163) );
  XOR U1021 ( .A(p_input[488]), .B(p_input[456]), .Z(n1164) );
  XNOR U1022 ( .A(n859), .B(n1159), .Z(n1161) );
  XOR U1023 ( .A(n1165), .B(n1166), .Z(n859) );
  AND U1024 ( .A(n168), .B(n1167), .Z(n1166) );
  XOR U1025 ( .A(p_input[424]), .B(p_input[392]), .Z(n1167) );
  XOR U1026 ( .A(n1168), .B(n1169), .Z(n1159) );
  AND U1027 ( .A(n1170), .B(n1171), .Z(n1169) );
  XOR U1028 ( .A(n1168), .B(n874), .Z(n1171) );
  XNOR U1029 ( .A(p_input[455]), .B(n1172), .Z(n874) );
  AND U1030 ( .A(n170), .B(n1173), .Z(n1172) );
  XOR U1031 ( .A(p_input[487]), .B(p_input[455]), .Z(n1173) );
  XNOR U1032 ( .A(n871), .B(n1168), .Z(n1170) );
  XOR U1033 ( .A(n1174), .B(n1175), .Z(n871) );
  AND U1034 ( .A(n168), .B(n1176), .Z(n1175) );
  XOR U1035 ( .A(p_input[423]), .B(p_input[391]), .Z(n1176) );
  XOR U1036 ( .A(n1177), .B(n1178), .Z(n1168) );
  AND U1037 ( .A(n1179), .B(n1180), .Z(n1178) );
  XOR U1038 ( .A(n1177), .B(n886), .Z(n1180) );
  XNOR U1039 ( .A(p_input[454]), .B(n1181), .Z(n886) );
  AND U1040 ( .A(n170), .B(n1182), .Z(n1181) );
  XOR U1041 ( .A(p_input[486]), .B(p_input[454]), .Z(n1182) );
  XNOR U1042 ( .A(n883), .B(n1177), .Z(n1179) );
  XOR U1043 ( .A(n1183), .B(n1184), .Z(n883) );
  AND U1044 ( .A(n168), .B(n1185), .Z(n1184) );
  XOR U1045 ( .A(p_input[422]), .B(p_input[390]), .Z(n1185) );
  XOR U1046 ( .A(n1186), .B(n1187), .Z(n1177) );
  AND U1047 ( .A(n1188), .B(n1189), .Z(n1187) );
  XOR U1048 ( .A(n898), .B(n1186), .Z(n1189) );
  XNOR U1049 ( .A(p_input[453]), .B(n1190), .Z(n898) );
  AND U1050 ( .A(n170), .B(n1191), .Z(n1190) );
  XOR U1051 ( .A(p_input[485]), .B(p_input[453]), .Z(n1191) );
  XNOR U1052 ( .A(n1186), .B(n895), .Z(n1188) );
  XOR U1053 ( .A(n1192), .B(n1193), .Z(n895) );
  AND U1054 ( .A(n168), .B(n1194), .Z(n1193) );
  XOR U1055 ( .A(p_input[421]), .B(p_input[389]), .Z(n1194) );
  XOR U1056 ( .A(n1195), .B(n1196), .Z(n1186) );
  AND U1057 ( .A(n1197), .B(n1198), .Z(n1196) );
  XOR U1058 ( .A(n1195), .B(n910), .Z(n1198) );
  XNOR U1059 ( .A(p_input[452]), .B(n1199), .Z(n910) );
  AND U1060 ( .A(n170), .B(n1200), .Z(n1199) );
  XOR U1061 ( .A(p_input[484]), .B(p_input[452]), .Z(n1200) );
  XNOR U1062 ( .A(n907), .B(n1195), .Z(n1197) );
  XOR U1063 ( .A(n1201), .B(n1202), .Z(n907) );
  AND U1064 ( .A(n168), .B(n1203), .Z(n1202) );
  XOR U1065 ( .A(p_input[420]), .B(p_input[388]), .Z(n1203) );
  XOR U1066 ( .A(n1204), .B(n1205), .Z(n1195) );
  AND U1067 ( .A(n1206), .B(n1207), .Z(n1205) );
  XOR U1068 ( .A(n1204), .B(n922), .Z(n1207) );
  XNOR U1069 ( .A(p_input[451]), .B(n1208), .Z(n922) );
  AND U1070 ( .A(n170), .B(n1209), .Z(n1208) );
  XOR U1071 ( .A(p_input[483]), .B(p_input[451]), .Z(n1209) );
  XNOR U1072 ( .A(n919), .B(n1204), .Z(n1206) );
  XOR U1073 ( .A(n1210), .B(n1211), .Z(n919) );
  AND U1074 ( .A(n168), .B(n1212), .Z(n1211) );
  XOR U1075 ( .A(p_input[419]), .B(p_input[387]), .Z(n1212) );
  XOR U1076 ( .A(n1213), .B(n1214), .Z(n1204) );
  AND U1077 ( .A(n1215), .B(n1216), .Z(n1214) );
  XOR U1078 ( .A(n1213), .B(n934), .Z(n1216) );
  XNOR U1079 ( .A(p_input[450]), .B(n1217), .Z(n934) );
  AND U1080 ( .A(n170), .B(n1218), .Z(n1217) );
  XOR U1081 ( .A(p_input[482]), .B(p_input[450]), .Z(n1218) );
  XNOR U1082 ( .A(n931), .B(n1213), .Z(n1215) );
  XOR U1083 ( .A(n1219), .B(n1220), .Z(n931) );
  AND U1084 ( .A(n168), .B(n1221), .Z(n1220) );
  XOR U1085 ( .A(p_input[418]), .B(p_input[386]), .Z(n1221) );
  XOR U1086 ( .A(n1222), .B(n1223), .Z(n1213) );
  AND U1087 ( .A(n1224), .B(n1225), .Z(n1223) );
  XNOR U1088 ( .A(n1226), .B(n947), .Z(n1225) );
  XNOR U1089 ( .A(p_input[449]), .B(n1227), .Z(n947) );
  AND U1090 ( .A(n170), .B(n1228), .Z(n1227) );
  XNOR U1091 ( .A(p_input[481]), .B(n1229), .Z(n1228) );
  IV U1092 ( .A(p_input[449]), .Z(n1229) );
  XNOR U1093 ( .A(n944), .B(n1222), .Z(n1224) );
  XNOR U1094 ( .A(p_input[385]), .B(n1230), .Z(n944) );
  AND U1095 ( .A(n168), .B(n1231), .Z(n1230) );
  XOR U1096 ( .A(p_input[417]), .B(p_input[385]), .Z(n1231) );
  IV U1097 ( .A(n1226), .Z(n1222) );
  AND U1098 ( .A(n952), .B(n955), .Z(n1226) );
  XOR U1099 ( .A(p_input[448]), .B(n1232), .Z(n955) );
  AND U1100 ( .A(n170), .B(n1233), .Z(n1232) );
  XOR U1101 ( .A(p_input[480]), .B(p_input[448]), .Z(n1233) );
  XOR U1102 ( .A(n1234), .B(n1235), .Z(n170) );
  AND U1103 ( .A(n1236), .B(n1237), .Z(n1235) );
  XNOR U1104 ( .A(p_input[511]), .B(n1234), .Z(n1237) );
  XOR U1105 ( .A(n1234), .B(p_input[479]), .Z(n1236) );
  XOR U1106 ( .A(n1238), .B(n1239), .Z(n1234) );
  AND U1107 ( .A(n1240), .B(n1241), .Z(n1239) );
  XNOR U1108 ( .A(p_input[510]), .B(n1238), .Z(n1241) );
  XOR U1109 ( .A(n1238), .B(p_input[478]), .Z(n1240) );
  XOR U1110 ( .A(n1242), .B(n1243), .Z(n1238) );
  AND U1111 ( .A(n1244), .B(n1245), .Z(n1243) );
  XNOR U1112 ( .A(p_input[509]), .B(n1242), .Z(n1245) );
  XOR U1113 ( .A(n1242), .B(p_input[477]), .Z(n1244) );
  XOR U1114 ( .A(n1246), .B(n1247), .Z(n1242) );
  AND U1115 ( .A(n1248), .B(n1249), .Z(n1247) );
  XNOR U1116 ( .A(p_input[508]), .B(n1246), .Z(n1249) );
  XOR U1117 ( .A(n1246), .B(p_input[476]), .Z(n1248) );
  XOR U1118 ( .A(n1250), .B(n1251), .Z(n1246) );
  AND U1119 ( .A(n1252), .B(n1253), .Z(n1251) );
  XNOR U1120 ( .A(p_input[507]), .B(n1250), .Z(n1253) );
  XOR U1121 ( .A(n1250), .B(p_input[475]), .Z(n1252) );
  XOR U1122 ( .A(n1254), .B(n1255), .Z(n1250) );
  AND U1123 ( .A(n1256), .B(n1257), .Z(n1255) );
  XNOR U1124 ( .A(p_input[506]), .B(n1254), .Z(n1257) );
  XOR U1125 ( .A(n1254), .B(p_input[474]), .Z(n1256) );
  XOR U1126 ( .A(n1258), .B(n1259), .Z(n1254) );
  AND U1127 ( .A(n1260), .B(n1261), .Z(n1259) );
  XNOR U1128 ( .A(p_input[505]), .B(n1258), .Z(n1261) );
  XOR U1129 ( .A(n1258), .B(p_input[473]), .Z(n1260) );
  XOR U1130 ( .A(n1262), .B(n1263), .Z(n1258) );
  AND U1131 ( .A(n1264), .B(n1265), .Z(n1263) );
  XNOR U1132 ( .A(p_input[504]), .B(n1262), .Z(n1265) );
  XOR U1133 ( .A(n1262), .B(p_input[472]), .Z(n1264) );
  XOR U1134 ( .A(n1266), .B(n1267), .Z(n1262) );
  AND U1135 ( .A(n1268), .B(n1269), .Z(n1267) );
  XNOR U1136 ( .A(p_input[503]), .B(n1266), .Z(n1269) );
  XOR U1137 ( .A(n1266), .B(p_input[471]), .Z(n1268) );
  XOR U1138 ( .A(n1270), .B(n1271), .Z(n1266) );
  AND U1139 ( .A(n1272), .B(n1273), .Z(n1271) );
  XNOR U1140 ( .A(p_input[502]), .B(n1270), .Z(n1273) );
  XOR U1141 ( .A(n1270), .B(p_input[470]), .Z(n1272) );
  XOR U1142 ( .A(n1274), .B(n1275), .Z(n1270) );
  AND U1143 ( .A(n1276), .B(n1277), .Z(n1275) );
  XNOR U1144 ( .A(p_input[501]), .B(n1274), .Z(n1277) );
  XOR U1145 ( .A(n1274), .B(p_input[469]), .Z(n1276) );
  XOR U1146 ( .A(n1278), .B(n1279), .Z(n1274) );
  AND U1147 ( .A(n1280), .B(n1281), .Z(n1279) );
  XNOR U1148 ( .A(p_input[500]), .B(n1278), .Z(n1281) );
  XOR U1149 ( .A(n1278), .B(p_input[468]), .Z(n1280) );
  XOR U1150 ( .A(n1282), .B(n1283), .Z(n1278) );
  AND U1151 ( .A(n1284), .B(n1285), .Z(n1283) );
  XNOR U1152 ( .A(p_input[499]), .B(n1282), .Z(n1285) );
  XOR U1153 ( .A(n1282), .B(p_input[467]), .Z(n1284) );
  XOR U1154 ( .A(n1286), .B(n1287), .Z(n1282) );
  AND U1155 ( .A(n1288), .B(n1289), .Z(n1287) );
  XNOR U1156 ( .A(p_input[498]), .B(n1286), .Z(n1289) );
  XOR U1157 ( .A(n1286), .B(p_input[466]), .Z(n1288) );
  XOR U1158 ( .A(n1290), .B(n1291), .Z(n1286) );
  AND U1159 ( .A(n1292), .B(n1293), .Z(n1291) );
  XNOR U1160 ( .A(p_input[497]), .B(n1290), .Z(n1293) );
  XOR U1161 ( .A(n1290), .B(p_input[465]), .Z(n1292) );
  XOR U1162 ( .A(n1294), .B(n1295), .Z(n1290) );
  AND U1163 ( .A(n1296), .B(n1297), .Z(n1295) );
  XNOR U1164 ( .A(p_input[496]), .B(n1294), .Z(n1297) );
  XOR U1165 ( .A(n1294), .B(p_input[464]), .Z(n1296) );
  XOR U1166 ( .A(n1298), .B(n1299), .Z(n1294) );
  AND U1167 ( .A(n1300), .B(n1301), .Z(n1299) );
  XNOR U1168 ( .A(p_input[495]), .B(n1298), .Z(n1301) );
  XOR U1169 ( .A(n1298), .B(p_input[463]), .Z(n1300) );
  XOR U1170 ( .A(n1302), .B(n1303), .Z(n1298) );
  AND U1171 ( .A(n1304), .B(n1305), .Z(n1303) );
  XNOR U1172 ( .A(p_input[494]), .B(n1302), .Z(n1305) );
  XOR U1173 ( .A(n1302), .B(p_input[462]), .Z(n1304) );
  XOR U1174 ( .A(n1306), .B(n1307), .Z(n1302) );
  AND U1175 ( .A(n1308), .B(n1309), .Z(n1307) );
  XNOR U1176 ( .A(p_input[493]), .B(n1306), .Z(n1309) );
  XOR U1177 ( .A(n1306), .B(p_input[461]), .Z(n1308) );
  XOR U1178 ( .A(n1310), .B(n1311), .Z(n1306) );
  AND U1179 ( .A(n1312), .B(n1313), .Z(n1311) );
  XNOR U1180 ( .A(p_input[492]), .B(n1310), .Z(n1313) );
  XOR U1181 ( .A(n1310), .B(p_input[460]), .Z(n1312) );
  XOR U1182 ( .A(n1314), .B(n1315), .Z(n1310) );
  AND U1183 ( .A(n1316), .B(n1317), .Z(n1315) );
  XNOR U1184 ( .A(p_input[491]), .B(n1314), .Z(n1317) );
  XOR U1185 ( .A(n1314), .B(p_input[459]), .Z(n1316) );
  XOR U1186 ( .A(n1318), .B(n1319), .Z(n1314) );
  AND U1187 ( .A(n1320), .B(n1321), .Z(n1319) );
  XNOR U1188 ( .A(p_input[490]), .B(n1318), .Z(n1321) );
  XOR U1189 ( .A(n1318), .B(p_input[458]), .Z(n1320) );
  XOR U1190 ( .A(n1322), .B(n1323), .Z(n1318) );
  AND U1191 ( .A(n1324), .B(n1325), .Z(n1323) );
  XNOR U1192 ( .A(p_input[489]), .B(n1322), .Z(n1325) );
  XOR U1193 ( .A(n1322), .B(p_input[457]), .Z(n1324) );
  XOR U1194 ( .A(n1326), .B(n1327), .Z(n1322) );
  AND U1195 ( .A(n1328), .B(n1329), .Z(n1327) );
  XNOR U1196 ( .A(p_input[488]), .B(n1326), .Z(n1329) );
  XOR U1197 ( .A(n1326), .B(p_input[456]), .Z(n1328) );
  XOR U1198 ( .A(n1330), .B(n1331), .Z(n1326) );
  AND U1199 ( .A(n1332), .B(n1333), .Z(n1331) );
  XNOR U1200 ( .A(p_input[487]), .B(n1330), .Z(n1333) );
  XOR U1201 ( .A(n1330), .B(p_input[455]), .Z(n1332) );
  XOR U1202 ( .A(n1334), .B(n1335), .Z(n1330) );
  AND U1203 ( .A(n1336), .B(n1337), .Z(n1335) );
  XNOR U1204 ( .A(p_input[486]), .B(n1334), .Z(n1337) );
  XOR U1205 ( .A(n1334), .B(p_input[454]), .Z(n1336) );
  XOR U1206 ( .A(n1338), .B(n1339), .Z(n1334) );
  AND U1207 ( .A(n1340), .B(n1341), .Z(n1339) );
  XNOR U1208 ( .A(p_input[485]), .B(n1338), .Z(n1341) );
  XOR U1209 ( .A(n1338), .B(p_input[453]), .Z(n1340) );
  XOR U1210 ( .A(n1342), .B(n1343), .Z(n1338) );
  AND U1211 ( .A(n1344), .B(n1345), .Z(n1343) );
  XNOR U1212 ( .A(p_input[484]), .B(n1342), .Z(n1345) );
  XOR U1213 ( .A(n1342), .B(p_input[452]), .Z(n1344) );
  XOR U1214 ( .A(n1346), .B(n1347), .Z(n1342) );
  AND U1215 ( .A(n1348), .B(n1349), .Z(n1347) );
  XNOR U1216 ( .A(p_input[483]), .B(n1346), .Z(n1349) );
  XOR U1217 ( .A(n1346), .B(p_input[451]), .Z(n1348) );
  XOR U1218 ( .A(n1350), .B(n1351), .Z(n1346) );
  AND U1219 ( .A(n1352), .B(n1353), .Z(n1351) );
  XNOR U1220 ( .A(p_input[482]), .B(n1350), .Z(n1353) );
  XOR U1221 ( .A(n1350), .B(p_input[450]), .Z(n1352) );
  XNOR U1222 ( .A(n1354), .B(n1355), .Z(n1350) );
  AND U1223 ( .A(n1356), .B(n1357), .Z(n1355) );
  XOR U1224 ( .A(p_input[481]), .B(n1354), .Z(n1357) );
  XNOR U1225 ( .A(p_input[449]), .B(n1354), .Z(n1356) );
  AND U1226 ( .A(p_input[480]), .B(n1358), .Z(n1354) );
  IV U1227 ( .A(p_input[448]), .Z(n1358) );
  XNOR U1228 ( .A(p_input[384]), .B(n1359), .Z(n952) );
  AND U1229 ( .A(n168), .B(n1360), .Z(n1359) );
  XOR U1230 ( .A(p_input[416]), .B(p_input[384]), .Z(n1360) );
  XOR U1231 ( .A(n1361), .B(n1362), .Z(n168) );
  AND U1232 ( .A(n1363), .B(n1364), .Z(n1362) );
  XNOR U1233 ( .A(p_input[447]), .B(n1361), .Z(n1364) );
  XOR U1234 ( .A(n1361), .B(p_input[415]), .Z(n1363) );
  XOR U1235 ( .A(n1365), .B(n1366), .Z(n1361) );
  AND U1236 ( .A(n1367), .B(n1368), .Z(n1366) );
  XNOR U1237 ( .A(p_input[446]), .B(n1365), .Z(n1368) );
  XNOR U1238 ( .A(n1365), .B(n967), .Z(n1367) );
  IV U1239 ( .A(p_input[414]), .Z(n967) );
  XOR U1240 ( .A(n1369), .B(n1370), .Z(n1365) );
  AND U1241 ( .A(n1371), .B(n1372), .Z(n1370) );
  XNOR U1242 ( .A(p_input[445]), .B(n1369), .Z(n1372) );
  XNOR U1243 ( .A(n1369), .B(n976), .Z(n1371) );
  IV U1244 ( .A(p_input[413]), .Z(n976) );
  XOR U1245 ( .A(n1373), .B(n1374), .Z(n1369) );
  AND U1246 ( .A(n1375), .B(n1376), .Z(n1374) );
  XNOR U1247 ( .A(p_input[444]), .B(n1373), .Z(n1376) );
  XNOR U1248 ( .A(n1373), .B(n985), .Z(n1375) );
  IV U1249 ( .A(p_input[412]), .Z(n985) );
  XOR U1250 ( .A(n1377), .B(n1378), .Z(n1373) );
  AND U1251 ( .A(n1379), .B(n1380), .Z(n1378) );
  XNOR U1252 ( .A(p_input[443]), .B(n1377), .Z(n1380) );
  XNOR U1253 ( .A(n1377), .B(n994), .Z(n1379) );
  IV U1254 ( .A(p_input[411]), .Z(n994) );
  XOR U1255 ( .A(n1381), .B(n1382), .Z(n1377) );
  AND U1256 ( .A(n1383), .B(n1384), .Z(n1382) );
  XNOR U1257 ( .A(p_input[442]), .B(n1381), .Z(n1384) );
  XNOR U1258 ( .A(n1381), .B(n1003), .Z(n1383) );
  IV U1259 ( .A(p_input[410]), .Z(n1003) );
  XOR U1260 ( .A(n1385), .B(n1386), .Z(n1381) );
  AND U1261 ( .A(n1387), .B(n1388), .Z(n1386) );
  XNOR U1262 ( .A(p_input[441]), .B(n1385), .Z(n1388) );
  XNOR U1263 ( .A(n1385), .B(n1012), .Z(n1387) );
  IV U1264 ( .A(p_input[409]), .Z(n1012) );
  XOR U1265 ( .A(n1389), .B(n1390), .Z(n1385) );
  AND U1266 ( .A(n1391), .B(n1392), .Z(n1390) );
  XNOR U1267 ( .A(p_input[440]), .B(n1389), .Z(n1392) );
  XNOR U1268 ( .A(n1389), .B(n1021), .Z(n1391) );
  IV U1269 ( .A(p_input[408]), .Z(n1021) );
  XOR U1270 ( .A(n1393), .B(n1394), .Z(n1389) );
  AND U1271 ( .A(n1395), .B(n1396), .Z(n1394) );
  XNOR U1272 ( .A(p_input[439]), .B(n1393), .Z(n1396) );
  XNOR U1273 ( .A(n1393), .B(n1030), .Z(n1395) );
  IV U1274 ( .A(p_input[407]), .Z(n1030) );
  XOR U1275 ( .A(n1397), .B(n1398), .Z(n1393) );
  AND U1276 ( .A(n1399), .B(n1400), .Z(n1398) );
  XNOR U1277 ( .A(p_input[438]), .B(n1397), .Z(n1400) );
  XNOR U1278 ( .A(n1397), .B(n1039), .Z(n1399) );
  IV U1279 ( .A(p_input[406]), .Z(n1039) );
  XOR U1280 ( .A(n1401), .B(n1402), .Z(n1397) );
  AND U1281 ( .A(n1403), .B(n1404), .Z(n1402) );
  XNOR U1282 ( .A(p_input[437]), .B(n1401), .Z(n1404) );
  XNOR U1283 ( .A(n1401), .B(n1048), .Z(n1403) );
  IV U1284 ( .A(p_input[405]), .Z(n1048) );
  XOR U1285 ( .A(n1405), .B(n1406), .Z(n1401) );
  AND U1286 ( .A(n1407), .B(n1408), .Z(n1406) );
  XNOR U1287 ( .A(p_input[436]), .B(n1405), .Z(n1408) );
  XNOR U1288 ( .A(n1405), .B(n1057), .Z(n1407) );
  IV U1289 ( .A(p_input[404]), .Z(n1057) );
  XOR U1290 ( .A(n1409), .B(n1410), .Z(n1405) );
  AND U1291 ( .A(n1411), .B(n1412), .Z(n1410) );
  XNOR U1292 ( .A(p_input[435]), .B(n1409), .Z(n1412) );
  XNOR U1293 ( .A(n1409), .B(n1066), .Z(n1411) );
  IV U1294 ( .A(p_input[403]), .Z(n1066) );
  XOR U1295 ( .A(n1413), .B(n1414), .Z(n1409) );
  AND U1296 ( .A(n1415), .B(n1416), .Z(n1414) );
  XNOR U1297 ( .A(p_input[434]), .B(n1413), .Z(n1416) );
  XNOR U1298 ( .A(n1413), .B(n1075), .Z(n1415) );
  IV U1299 ( .A(p_input[402]), .Z(n1075) );
  XOR U1300 ( .A(n1417), .B(n1418), .Z(n1413) );
  AND U1301 ( .A(n1419), .B(n1420), .Z(n1418) );
  XNOR U1302 ( .A(p_input[433]), .B(n1417), .Z(n1420) );
  XNOR U1303 ( .A(n1417), .B(n1084), .Z(n1419) );
  IV U1304 ( .A(p_input[401]), .Z(n1084) );
  XOR U1305 ( .A(n1421), .B(n1422), .Z(n1417) );
  AND U1306 ( .A(n1423), .B(n1424), .Z(n1422) );
  XNOR U1307 ( .A(p_input[432]), .B(n1421), .Z(n1424) );
  XNOR U1308 ( .A(n1421), .B(n1093), .Z(n1423) );
  IV U1309 ( .A(p_input[400]), .Z(n1093) );
  XOR U1310 ( .A(n1425), .B(n1426), .Z(n1421) );
  AND U1311 ( .A(n1427), .B(n1428), .Z(n1426) );
  XNOR U1312 ( .A(p_input[431]), .B(n1425), .Z(n1428) );
  XNOR U1313 ( .A(n1425), .B(n1102), .Z(n1427) );
  IV U1314 ( .A(p_input[399]), .Z(n1102) );
  XOR U1315 ( .A(n1429), .B(n1430), .Z(n1425) );
  AND U1316 ( .A(n1431), .B(n1432), .Z(n1430) );
  XNOR U1317 ( .A(p_input[430]), .B(n1429), .Z(n1432) );
  XNOR U1318 ( .A(n1429), .B(n1111), .Z(n1431) );
  IV U1319 ( .A(p_input[398]), .Z(n1111) );
  XOR U1320 ( .A(n1433), .B(n1434), .Z(n1429) );
  AND U1321 ( .A(n1435), .B(n1436), .Z(n1434) );
  XNOR U1322 ( .A(p_input[429]), .B(n1433), .Z(n1436) );
  XNOR U1323 ( .A(n1433), .B(n1120), .Z(n1435) );
  IV U1324 ( .A(p_input[397]), .Z(n1120) );
  XOR U1325 ( .A(n1437), .B(n1438), .Z(n1433) );
  AND U1326 ( .A(n1439), .B(n1440), .Z(n1438) );
  XNOR U1327 ( .A(p_input[428]), .B(n1437), .Z(n1440) );
  XNOR U1328 ( .A(n1437), .B(n1129), .Z(n1439) );
  IV U1329 ( .A(p_input[396]), .Z(n1129) );
  XOR U1330 ( .A(n1441), .B(n1442), .Z(n1437) );
  AND U1331 ( .A(n1443), .B(n1444), .Z(n1442) );
  XNOR U1332 ( .A(p_input[427]), .B(n1441), .Z(n1444) );
  XNOR U1333 ( .A(n1441), .B(n1138), .Z(n1443) );
  IV U1334 ( .A(p_input[395]), .Z(n1138) );
  XOR U1335 ( .A(n1445), .B(n1446), .Z(n1441) );
  AND U1336 ( .A(n1447), .B(n1448), .Z(n1446) );
  XNOR U1337 ( .A(p_input[426]), .B(n1445), .Z(n1448) );
  XNOR U1338 ( .A(n1445), .B(n1147), .Z(n1447) );
  IV U1339 ( .A(p_input[394]), .Z(n1147) );
  XOR U1340 ( .A(n1449), .B(n1450), .Z(n1445) );
  AND U1341 ( .A(n1451), .B(n1452), .Z(n1450) );
  XNOR U1342 ( .A(p_input[425]), .B(n1449), .Z(n1452) );
  XNOR U1343 ( .A(n1449), .B(n1156), .Z(n1451) );
  IV U1344 ( .A(p_input[393]), .Z(n1156) );
  XOR U1345 ( .A(n1453), .B(n1454), .Z(n1449) );
  AND U1346 ( .A(n1455), .B(n1456), .Z(n1454) );
  XNOR U1347 ( .A(p_input[424]), .B(n1453), .Z(n1456) );
  XNOR U1348 ( .A(n1453), .B(n1165), .Z(n1455) );
  IV U1349 ( .A(p_input[392]), .Z(n1165) );
  XOR U1350 ( .A(n1457), .B(n1458), .Z(n1453) );
  AND U1351 ( .A(n1459), .B(n1460), .Z(n1458) );
  XNOR U1352 ( .A(p_input[423]), .B(n1457), .Z(n1460) );
  XNOR U1353 ( .A(n1457), .B(n1174), .Z(n1459) );
  IV U1354 ( .A(p_input[391]), .Z(n1174) );
  XOR U1355 ( .A(n1461), .B(n1462), .Z(n1457) );
  AND U1356 ( .A(n1463), .B(n1464), .Z(n1462) );
  XNOR U1357 ( .A(p_input[422]), .B(n1461), .Z(n1464) );
  XNOR U1358 ( .A(n1461), .B(n1183), .Z(n1463) );
  IV U1359 ( .A(p_input[390]), .Z(n1183) );
  XOR U1360 ( .A(n1465), .B(n1466), .Z(n1461) );
  AND U1361 ( .A(n1467), .B(n1468), .Z(n1466) );
  XNOR U1362 ( .A(p_input[421]), .B(n1465), .Z(n1468) );
  XNOR U1363 ( .A(n1465), .B(n1192), .Z(n1467) );
  IV U1364 ( .A(p_input[389]), .Z(n1192) );
  XOR U1365 ( .A(n1469), .B(n1470), .Z(n1465) );
  AND U1366 ( .A(n1471), .B(n1472), .Z(n1470) );
  XNOR U1367 ( .A(p_input[420]), .B(n1469), .Z(n1472) );
  XNOR U1368 ( .A(n1469), .B(n1201), .Z(n1471) );
  IV U1369 ( .A(p_input[388]), .Z(n1201) );
  XOR U1370 ( .A(n1473), .B(n1474), .Z(n1469) );
  AND U1371 ( .A(n1475), .B(n1476), .Z(n1474) );
  XNOR U1372 ( .A(p_input[419]), .B(n1473), .Z(n1476) );
  XNOR U1373 ( .A(n1473), .B(n1210), .Z(n1475) );
  IV U1374 ( .A(p_input[387]), .Z(n1210) );
  XOR U1375 ( .A(n1477), .B(n1478), .Z(n1473) );
  AND U1376 ( .A(n1479), .B(n1480), .Z(n1478) );
  XNOR U1377 ( .A(p_input[418]), .B(n1477), .Z(n1480) );
  XNOR U1378 ( .A(n1477), .B(n1219), .Z(n1479) );
  IV U1379 ( .A(p_input[386]), .Z(n1219) );
  XNOR U1380 ( .A(n1481), .B(n1482), .Z(n1477) );
  AND U1381 ( .A(n1483), .B(n1484), .Z(n1482) );
  XOR U1382 ( .A(p_input[417]), .B(n1481), .Z(n1484) );
  XNOR U1383 ( .A(p_input[385]), .B(n1481), .Z(n1483) );
  AND U1384 ( .A(p_input[416]), .B(n1485), .Z(n1481) );
  IV U1385 ( .A(p_input[384]), .Z(n1485) );
  XOR U1386 ( .A(n1486), .B(n1487), .Z(n575) );
  AND U1387 ( .A(n180), .B(n1488), .Z(n1487) );
  XNOR U1388 ( .A(n1489), .B(n1486), .Z(n1488) );
  XOR U1389 ( .A(n1490), .B(n1491), .Z(n180) );
  AND U1390 ( .A(n1492), .B(n1493), .Z(n1491) );
  XNOR U1391 ( .A(n590), .B(n1490), .Z(n1493) );
  AND U1392 ( .A(p_input[383]), .B(p_input[351]), .Z(n590) );
  XNOR U1393 ( .A(n1490), .B(n587), .Z(n1492) );
  IV U1394 ( .A(n1494), .Z(n587) );
  AND U1395 ( .A(p_input[287]), .B(p_input[319]), .Z(n1494) );
  XOR U1396 ( .A(n1495), .B(n1496), .Z(n1490) );
  AND U1397 ( .A(n1497), .B(n1498), .Z(n1496) );
  XOR U1398 ( .A(n1495), .B(n602), .Z(n1498) );
  XNOR U1399 ( .A(p_input[350]), .B(n1499), .Z(n602) );
  AND U1400 ( .A(n174), .B(n1500), .Z(n1499) );
  XOR U1401 ( .A(p_input[382]), .B(p_input[350]), .Z(n1500) );
  XNOR U1402 ( .A(n599), .B(n1495), .Z(n1497) );
  XOR U1403 ( .A(n1501), .B(n1502), .Z(n599) );
  AND U1404 ( .A(n171), .B(n1503), .Z(n1502) );
  XOR U1405 ( .A(p_input[318]), .B(p_input[286]), .Z(n1503) );
  XOR U1406 ( .A(n1504), .B(n1505), .Z(n1495) );
  AND U1407 ( .A(n1506), .B(n1507), .Z(n1505) );
  XOR U1408 ( .A(n1504), .B(n614), .Z(n1507) );
  XNOR U1409 ( .A(p_input[349]), .B(n1508), .Z(n614) );
  AND U1410 ( .A(n174), .B(n1509), .Z(n1508) );
  XOR U1411 ( .A(p_input[381]), .B(p_input[349]), .Z(n1509) );
  XNOR U1412 ( .A(n611), .B(n1504), .Z(n1506) );
  XOR U1413 ( .A(n1510), .B(n1511), .Z(n611) );
  AND U1414 ( .A(n171), .B(n1512), .Z(n1511) );
  XOR U1415 ( .A(p_input[317]), .B(p_input[285]), .Z(n1512) );
  XOR U1416 ( .A(n1513), .B(n1514), .Z(n1504) );
  AND U1417 ( .A(n1515), .B(n1516), .Z(n1514) );
  XOR U1418 ( .A(n1513), .B(n626), .Z(n1516) );
  XNOR U1419 ( .A(p_input[348]), .B(n1517), .Z(n626) );
  AND U1420 ( .A(n174), .B(n1518), .Z(n1517) );
  XOR U1421 ( .A(p_input[380]), .B(p_input[348]), .Z(n1518) );
  XNOR U1422 ( .A(n623), .B(n1513), .Z(n1515) );
  XOR U1423 ( .A(n1519), .B(n1520), .Z(n623) );
  AND U1424 ( .A(n171), .B(n1521), .Z(n1520) );
  XOR U1425 ( .A(p_input[316]), .B(p_input[284]), .Z(n1521) );
  XOR U1426 ( .A(n1522), .B(n1523), .Z(n1513) );
  AND U1427 ( .A(n1524), .B(n1525), .Z(n1523) );
  XOR U1428 ( .A(n1522), .B(n638), .Z(n1525) );
  XNOR U1429 ( .A(p_input[347]), .B(n1526), .Z(n638) );
  AND U1430 ( .A(n174), .B(n1527), .Z(n1526) );
  XOR U1431 ( .A(p_input[379]), .B(p_input[347]), .Z(n1527) );
  XNOR U1432 ( .A(n635), .B(n1522), .Z(n1524) );
  XOR U1433 ( .A(n1528), .B(n1529), .Z(n635) );
  AND U1434 ( .A(n171), .B(n1530), .Z(n1529) );
  XOR U1435 ( .A(p_input[315]), .B(p_input[283]), .Z(n1530) );
  XOR U1436 ( .A(n1531), .B(n1532), .Z(n1522) );
  AND U1437 ( .A(n1533), .B(n1534), .Z(n1532) );
  XOR U1438 ( .A(n1531), .B(n650), .Z(n1534) );
  XNOR U1439 ( .A(p_input[346]), .B(n1535), .Z(n650) );
  AND U1440 ( .A(n174), .B(n1536), .Z(n1535) );
  XOR U1441 ( .A(p_input[378]), .B(p_input[346]), .Z(n1536) );
  XNOR U1442 ( .A(n647), .B(n1531), .Z(n1533) );
  XOR U1443 ( .A(n1537), .B(n1538), .Z(n647) );
  AND U1444 ( .A(n171), .B(n1539), .Z(n1538) );
  XOR U1445 ( .A(p_input[314]), .B(p_input[282]), .Z(n1539) );
  XOR U1446 ( .A(n1540), .B(n1541), .Z(n1531) );
  AND U1447 ( .A(n1542), .B(n1543), .Z(n1541) );
  XOR U1448 ( .A(n1540), .B(n662), .Z(n1543) );
  XNOR U1449 ( .A(p_input[345]), .B(n1544), .Z(n662) );
  AND U1450 ( .A(n174), .B(n1545), .Z(n1544) );
  XOR U1451 ( .A(p_input[377]), .B(p_input[345]), .Z(n1545) );
  XNOR U1452 ( .A(n659), .B(n1540), .Z(n1542) );
  XOR U1453 ( .A(n1546), .B(n1547), .Z(n659) );
  AND U1454 ( .A(n171), .B(n1548), .Z(n1547) );
  XOR U1455 ( .A(p_input[313]), .B(p_input[281]), .Z(n1548) );
  XOR U1456 ( .A(n1549), .B(n1550), .Z(n1540) );
  AND U1457 ( .A(n1551), .B(n1552), .Z(n1550) );
  XOR U1458 ( .A(n1549), .B(n674), .Z(n1552) );
  XNOR U1459 ( .A(p_input[344]), .B(n1553), .Z(n674) );
  AND U1460 ( .A(n174), .B(n1554), .Z(n1553) );
  XOR U1461 ( .A(p_input[376]), .B(p_input[344]), .Z(n1554) );
  XNOR U1462 ( .A(n671), .B(n1549), .Z(n1551) );
  XOR U1463 ( .A(n1555), .B(n1556), .Z(n671) );
  AND U1464 ( .A(n171), .B(n1557), .Z(n1556) );
  XOR U1465 ( .A(p_input[312]), .B(p_input[280]), .Z(n1557) );
  XOR U1466 ( .A(n1558), .B(n1559), .Z(n1549) );
  AND U1467 ( .A(n1560), .B(n1561), .Z(n1559) );
  XOR U1468 ( .A(n1558), .B(n686), .Z(n1561) );
  XNOR U1469 ( .A(p_input[343]), .B(n1562), .Z(n686) );
  AND U1470 ( .A(n174), .B(n1563), .Z(n1562) );
  XOR U1471 ( .A(p_input[375]), .B(p_input[343]), .Z(n1563) );
  XNOR U1472 ( .A(n683), .B(n1558), .Z(n1560) );
  XOR U1473 ( .A(n1564), .B(n1565), .Z(n683) );
  AND U1474 ( .A(n171), .B(n1566), .Z(n1565) );
  XOR U1475 ( .A(p_input[311]), .B(p_input[279]), .Z(n1566) );
  XOR U1476 ( .A(n1567), .B(n1568), .Z(n1558) );
  AND U1477 ( .A(n1569), .B(n1570), .Z(n1568) );
  XOR U1478 ( .A(n1567), .B(n698), .Z(n1570) );
  XNOR U1479 ( .A(p_input[342]), .B(n1571), .Z(n698) );
  AND U1480 ( .A(n174), .B(n1572), .Z(n1571) );
  XOR U1481 ( .A(p_input[374]), .B(p_input[342]), .Z(n1572) );
  XNOR U1482 ( .A(n695), .B(n1567), .Z(n1569) );
  XOR U1483 ( .A(n1573), .B(n1574), .Z(n695) );
  AND U1484 ( .A(n171), .B(n1575), .Z(n1574) );
  XOR U1485 ( .A(p_input[310]), .B(p_input[278]), .Z(n1575) );
  XOR U1486 ( .A(n1576), .B(n1577), .Z(n1567) );
  AND U1487 ( .A(n1578), .B(n1579), .Z(n1577) );
  XOR U1488 ( .A(n1576), .B(n710), .Z(n1579) );
  XNOR U1489 ( .A(p_input[341]), .B(n1580), .Z(n710) );
  AND U1490 ( .A(n174), .B(n1581), .Z(n1580) );
  XOR U1491 ( .A(p_input[373]), .B(p_input[341]), .Z(n1581) );
  XNOR U1492 ( .A(n707), .B(n1576), .Z(n1578) );
  XOR U1493 ( .A(n1582), .B(n1583), .Z(n707) );
  AND U1494 ( .A(n171), .B(n1584), .Z(n1583) );
  XOR U1495 ( .A(p_input[309]), .B(p_input[277]), .Z(n1584) );
  XOR U1496 ( .A(n1585), .B(n1586), .Z(n1576) );
  AND U1497 ( .A(n1587), .B(n1588), .Z(n1586) );
  XOR U1498 ( .A(n1585), .B(n722), .Z(n1588) );
  XNOR U1499 ( .A(p_input[340]), .B(n1589), .Z(n722) );
  AND U1500 ( .A(n174), .B(n1590), .Z(n1589) );
  XOR U1501 ( .A(p_input[372]), .B(p_input[340]), .Z(n1590) );
  XNOR U1502 ( .A(n719), .B(n1585), .Z(n1587) );
  XOR U1503 ( .A(n1591), .B(n1592), .Z(n719) );
  AND U1504 ( .A(n171), .B(n1593), .Z(n1592) );
  XOR U1505 ( .A(p_input[308]), .B(p_input[276]), .Z(n1593) );
  XOR U1506 ( .A(n1594), .B(n1595), .Z(n1585) );
  AND U1507 ( .A(n1596), .B(n1597), .Z(n1595) );
  XOR U1508 ( .A(n1594), .B(n734), .Z(n1597) );
  XNOR U1509 ( .A(p_input[339]), .B(n1598), .Z(n734) );
  AND U1510 ( .A(n174), .B(n1599), .Z(n1598) );
  XOR U1511 ( .A(p_input[371]), .B(p_input[339]), .Z(n1599) );
  XNOR U1512 ( .A(n731), .B(n1594), .Z(n1596) );
  XOR U1513 ( .A(n1600), .B(n1601), .Z(n731) );
  AND U1514 ( .A(n171), .B(n1602), .Z(n1601) );
  XOR U1515 ( .A(p_input[307]), .B(p_input[275]), .Z(n1602) );
  XOR U1516 ( .A(n1603), .B(n1604), .Z(n1594) );
  AND U1517 ( .A(n1605), .B(n1606), .Z(n1604) );
  XOR U1518 ( .A(n1603), .B(n746), .Z(n1606) );
  XNOR U1519 ( .A(p_input[338]), .B(n1607), .Z(n746) );
  AND U1520 ( .A(n174), .B(n1608), .Z(n1607) );
  XOR U1521 ( .A(p_input[370]), .B(p_input[338]), .Z(n1608) );
  XNOR U1522 ( .A(n743), .B(n1603), .Z(n1605) );
  XOR U1523 ( .A(n1609), .B(n1610), .Z(n743) );
  AND U1524 ( .A(n171), .B(n1611), .Z(n1610) );
  XOR U1525 ( .A(p_input[306]), .B(p_input[274]), .Z(n1611) );
  XOR U1526 ( .A(n1612), .B(n1613), .Z(n1603) );
  AND U1527 ( .A(n1614), .B(n1615), .Z(n1613) );
  XOR U1528 ( .A(n1612), .B(n758), .Z(n1615) );
  XNOR U1529 ( .A(p_input[337]), .B(n1616), .Z(n758) );
  AND U1530 ( .A(n174), .B(n1617), .Z(n1616) );
  XOR U1531 ( .A(p_input[369]), .B(p_input[337]), .Z(n1617) );
  XNOR U1532 ( .A(n755), .B(n1612), .Z(n1614) );
  XOR U1533 ( .A(n1618), .B(n1619), .Z(n755) );
  AND U1534 ( .A(n171), .B(n1620), .Z(n1619) );
  XOR U1535 ( .A(p_input[305]), .B(p_input[273]), .Z(n1620) );
  XOR U1536 ( .A(n1621), .B(n1622), .Z(n1612) );
  AND U1537 ( .A(n1623), .B(n1624), .Z(n1622) );
  XOR U1538 ( .A(n1621), .B(n770), .Z(n1624) );
  XNOR U1539 ( .A(p_input[336]), .B(n1625), .Z(n770) );
  AND U1540 ( .A(n174), .B(n1626), .Z(n1625) );
  XOR U1541 ( .A(p_input[368]), .B(p_input[336]), .Z(n1626) );
  XNOR U1542 ( .A(n767), .B(n1621), .Z(n1623) );
  XOR U1543 ( .A(n1627), .B(n1628), .Z(n767) );
  AND U1544 ( .A(n171), .B(n1629), .Z(n1628) );
  XOR U1545 ( .A(p_input[304]), .B(p_input[272]), .Z(n1629) );
  XOR U1546 ( .A(n1630), .B(n1631), .Z(n1621) );
  AND U1547 ( .A(n1632), .B(n1633), .Z(n1631) );
  XOR U1548 ( .A(n1630), .B(n782), .Z(n1633) );
  XNOR U1549 ( .A(p_input[335]), .B(n1634), .Z(n782) );
  AND U1550 ( .A(n174), .B(n1635), .Z(n1634) );
  XOR U1551 ( .A(p_input[367]), .B(p_input[335]), .Z(n1635) );
  XNOR U1552 ( .A(n779), .B(n1630), .Z(n1632) );
  XOR U1553 ( .A(n1636), .B(n1637), .Z(n779) );
  AND U1554 ( .A(n171), .B(n1638), .Z(n1637) );
  XOR U1555 ( .A(p_input[303]), .B(p_input[271]), .Z(n1638) );
  XOR U1556 ( .A(n1639), .B(n1640), .Z(n1630) );
  AND U1557 ( .A(n1641), .B(n1642), .Z(n1640) );
  XOR U1558 ( .A(n1639), .B(n794), .Z(n1642) );
  XNOR U1559 ( .A(p_input[334]), .B(n1643), .Z(n794) );
  AND U1560 ( .A(n174), .B(n1644), .Z(n1643) );
  XOR U1561 ( .A(p_input[366]), .B(p_input[334]), .Z(n1644) );
  XNOR U1562 ( .A(n791), .B(n1639), .Z(n1641) );
  XOR U1563 ( .A(n1645), .B(n1646), .Z(n791) );
  AND U1564 ( .A(n171), .B(n1647), .Z(n1646) );
  XOR U1565 ( .A(p_input[302]), .B(p_input[270]), .Z(n1647) );
  XOR U1566 ( .A(n1648), .B(n1649), .Z(n1639) );
  AND U1567 ( .A(n1650), .B(n1651), .Z(n1649) );
  XOR U1568 ( .A(n1648), .B(n806), .Z(n1651) );
  XNOR U1569 ( .A(p_input[333]), .B(n1652), .Z(n806) );
  AND U1570 ( .A(n174), .B(n1653), .Z(n1652) );
  XOR U1571 ( .A(p_input[365]), .B(p_input[333]), .Z(n1653) );
  XNOR U1572 ( .A(n803), .B(n1648), .Z(n1650) );
  XOR U1573 ( .A(n1654), .B(n1655), .Z(n803) );
  AND U1574 ( .A(n171), .B(n1656), .Z(n1655) );
  XOR U1575 ( .A(p_input[301]), .B(p_input[269]), .Z(n1656) );
  XOR U1576 ( .A(n1657), .B(n1658), .Z(n1648) );
  AND U1577 ( .A(n1659), .B(n1660), .Z(n1658) );
  XOR U1578 ( .A(n1657), .B(n818), .Z(n1660) );
  XNOR U1579 ( .A(p_input[332]), .B(n1661), .Z(n818) );
  AND U1580 ( .A(n174), .B(n1662), .Z(n1661) );
  XOR U1581 ( .A(p_input[364]), .B(p_input[332]), .Z(n1662) );
  XNOR U1582 ( .A(n815), .B(n1657), .Z(n1659) );
  XOR U1583 ( .A(n1663), .B(n1664), .Z(n815) );
  AND U1584 ( .A(n171), .B(n1665), .Z(n1664) );
  XOR U1585 ( .A(p_input[300]), .B(p_input[268]), .Z(n1665) );
  XOR U1586 ( .A(n1666), .B(n1667), .Z(n1657) );
  AND U1587 ( .A(n1668), .B(n1669), .Z(n1667) );
  XOR U1588 ( .A(n1666), .B(n830), .Z(n1669) );
  XNOR U1589 ( .A(p_input[331]), .B(n1670), .Z(n830) );
  AND U1590 ( .A(n174), .B(n1671), .Z(n1670) );
  XOR U1591 ( .A(p_input[363]), .B(p_input[331]), .Z(n1671) );
  XNOR U1592 ( .A(n827), .B(n1666), .Z(n1668) );
  XOR U1593 ( .A(n1672), .B(n1673), .Z(n827) );
  AND U1594 ( .A(n171), .B(n1674), .Z(n1673) );
  XOR U1595 ( .A(p_input[299]), .B(p_input[267]), .Z(n1674) );
  XOR U1596 ( .A(n1675), .B(n1676), .Z(n1666) );
  AND U1597 ( .A(n1677), .B(n1678), .Z(n1676) );
  XOR U1598 ( .A(n1675), .B(n842), .Z(n1678) );
  XNOR U1599 ( .A(p_input[330]), .B(n1679), .Z(n842) );
  AND U1600 ( .A(n174), .B(n1680), .Z(n1679) );
  XOR U1601 ( .A(p_input[362]), .B(p_input[330]), .Z(n1680) );
  XNOR U1602 ( .A(n839), .B(n1675), .Z(n1677) );
  XOR U1603 ( .A(n1681), .B(n1682), .Z(n839) );
  AND U1604 ( .A(n171), .B(n1683), .Z(n1682) );
  XOR U1605 ( .A(p_input[298]), .B(p_input[266]), .Z(n1683) );
  XOR U1606 ( .A(n1684), .B(n1685), .Z(n1675) );
  AND U1607 ( .A(n1686), .B(n1687), .Z(n1685) );
  XOR U1608 ( .A(n1684), .B(n854), .Z(n1687) );
  XNOR U1609 ( .A(p_input[329]), .B(n1688), .Z(n854) );
  AND U1610 ( .A(n174), .B(n1689), .Z(n1688) );
  XOR U1611 ( .A(p_input[361]), .B(p_input[329]), .Z(n1689) );
  XNOR U1612 ( .A(n851), .B(n1684), .Z(n1686) );
  XOR U1613 ( .A(n1690), .B(n1691), .Z(n851) );
  AND U1614 ( .A(n171), .B(n1692), .Z(n1691) );
  XOR U1615 ( .A(p_input[297]), .B(p_input[265]), .Z(n1692) );
  XOR U1616 ( .A(n1693), .B(n1694), .Z(n1684) );
  AND U1617 ( .A(n1695), .B(n1696), .Z(n1694) );
  XOR U1618 ( .A(n1693), .B(n866), .Z(n1696) );
  XNOR U1619 ( .A(p_input[328]), .B(n1697), .Z(n866) );
  AND U1620 ( .A(n174), .B(n1698), .Z(n1697) );
  XOR U1621 ( .A(p_input[360]), .B(p_input[328]), .Z(n1698) );
  XNOR U1622 ( .A(n863), .B(n1693), .Z(n1695) );
  XOR U1623 ( .A(n1699), .B(n1700), .Z(n863) );
  AND U1624 ( .A(n171), .B(n1701), .Z(n1700) );
  XOR U1625 ( .A(p_input[296]), .B(p_input[264]), .Z(n1701) );
  XOR U1626 ( .A(n1702), .B(n1703), .Z(n1693) );
  AND U1627 ( .A(n1704), .B(n1705), .Z(n1703) );
  XOR U1628 ( .A(n1702), .B(n878), .Z(n1705) );
  XNOR U1629 ( .A(p_input[327]), .B(n1706), .Z(n878) );
  AND U1630 ( .A(n174), .B(n1707), .Z(n1706) );
  XOR U1631 ( .A(p_input[359]), .B(p_input[327]), .Z(n1707) );
  XNOR U1632 ( .A(n875), .B(n1702), .Z(n1704) );
  XOR U1633 ( .A(n1708), .B(n1709), .Z(n875) );
  AND U1634 ( .A(n171), .B(n1710), .Z(n1709) );
  XOR U1635 ( .A(p_input[295]), .B(p_input[263]), .Z(n1710) );
  XOR U1636 ( .A(n1711), .B(n1712), .Z(n1702) );
  AND U1637 ( .A(n1713), .B(n1714), .Z(n1712) );
  XOR U1638 ( .A(n1711), .B(n890), .Z(n1714) );
  XNOR U1639 ( .A(p_input[326]), .B(n1715), .Z(n890) );
  AND U1640 ( .A(n174), .B(n1716), .Z(n1715) );
  XOR U1641 ( .A(p_input[358]), .B(p_input[326]), .Z(n1716) );
  XNOR U1642 ( .A(n887), .B(n1711), .Z(n1713) );
  XOR U1643 ( .A(n1717), .B(n1718), .Z(n887) );
  AND U1644 ( .A(n171), .B(n1719), .Z(n1718) );
  XOR U1645 ( .A(p_input[294]), .B(p_input[262]), .Z(n1719) );
  XOR U1646 ( .A(n1720), .B(n1721), .Z(n1711) );
  AND U1647 ( .A(n1722), .B(n1723), .Z(n1721) );
  XOR U1648 ( .A(n902), .B(n1720), .Z(n1723) );
  XNOR U1649 ( .A(p_input[325]), .B(n1724), .Z(n902) );
  AND U1650 ( .A(n174), .B(n1725), .Z(n1724) );
  XOR U1651 ( .A(p_input[357]), .B(p_input[325]), .Z(n1725) );
  XNOR U1652 ( .A(n1720), .B(n899), .Z(n1722) );
  XOR U1653 ( .A(n1726), .B(n1727), .Z(n899) );
  AND U1654 ( .A(n171), .B(n1728), .Z(n1727) );
  XOR U1655 ( .A(p_input[293]), .B(p_input[261]), .Z(n1728) );
  XOR U1656 ( .A(n1729), .B(n1730), .Z(n1720) );
  AND U1657 ( .A(n1731), .B(n1732), .Z(n1730) );
  XOR U1658 ( .A(n1729), .B(n914), .Z(n1732) );
  XNOR U1659 ( .A(p_input[324]), .B(n1733), .Z(n914) );
  AND U1660 ( .A(n174), .B(n1734), .Z(n1733) );
  XOR U1661 ( .A(p_input[356]), .B(p_input[324]), .Z(n1734) );
  XNOR U1662 ( .A(n911), .B(n1729), .Z(n1731) );
  XOR U1663 ( .A(n1735), .B(n1736), .Z(n911) );
  AND U1664 ( .A(n171), .B(n1737), .Z(n1736) );
  XOR U1665 ( .A(p_input[292]), .B(p_input[260]), .Z(n1737) );
  XOR U1666 ( .A(n1738), .B(n1739), .Z(n1729) );
  AND U1667 ( .A(n1740), .B(n1741), .Z(n1739) );
  XOR U1668 ( .A(n1738), .B(n926), .Z(n1741) );
  XNOR U1669 ( .A(p_input[323]), .B(n1742), .Z(n926) );
  AND U1670 ( .A(n174), .B(n1743), .Z(n1742) );
  XOR U1671 ( .A(p_input[355]), .B(p_input[323]), .Z(n1743) );
  XNOR U1672 ( .A(n923), .B(n1738), .Z(n1740) );
  XOR U1673 ( .A(n1744), .B(n1745), .Z(n923) );
  AND U1674 ( .A(n171), .B(n1746), .Z(n1745) );
  XOR U1675 ( .A(p_input[291]), .B(p_input[259]), .Z(n1746) );
  XOR U1676 ( .A(n1747), .B(n1748), .Z(n1738) );
  AND U1677 ( .A(n1749), .B(n1750), .Z(n1748) );
  XOR U1678 ( .A(n1747), .B(n938), .Z(n1750) );
  XNOR U1679 ( .A(p_input[322]), .B(n1751), .Z(n938) );
  AND U1680 ( .A(n174), .B(n1752), .Z(n1751) );
  XOR U1681 ( .A(p_input[354]), .B(p_input[322]), .Z(n1752) );
  XNOR U1682 ( .A(n935), .B(n1747), .Z(n1749) );
  XOR U1683 ( .A(n1753), .B(n1754), .Z(n935) );
  AND U1684 ( .A(n171), .B(n1755), .Z(n1754) );
  XOR U1685 ( .A(p_input[290]), .B(p_input[258]), .Z(n1755) );
  XOR U1686 ( .A(n1756), .B(n1757), .Z(n1747) );
  AND U1687 ( .A(n1758), .B(n1759), .Z(n1757) );
  XNOR U1688 ( .A(n1760), .B(n951), .Z(n1759) );
  XNOR U1689 ( .A(p_input[321]), .B(n1761), .Z(n951) );
  AND U1690 ( .A(n174), .B(n1762), .Z(n1761) );
  XNOR U1691 ( .A(p_input[353]), .B(n1763), .Z(n1762) );
  IV U1692 ( .A(p_input[321]), .Z(n1763) );
  XNOR U1693 ( .A(n948), .B(n1756), .Z(n1758) );
  XNOR U1694 ( .A(p_input[257]), .B(n1764), .Z(n948) );
  AND U1695 ( .A(n171), .B(n1765), .Z(n1764) );
  XOR U1696 ( .A(p_input[289]), .B(p_input[257]), .Z(n1765) );
  IV U1697 ( .A(n1760), .Z(n1756) );
  AND U1698 ( .A(n1486), .B(n1489), .Z(n1760) );
  XOR U1699 ( .A(p_input[320]), .B(n1766), .Z(n1489) );
  AND U1700 ( .A(n174), .B(n1767), .Z(n1766) );
  XOR U1701 ( .A(p_input[352]), .B(p_input[320]), .Z(n1767) );
  XOR U1702 ( .A(n1768), .B(n1769), .Z(n174) );
  AND U1703 ( .A(n1770), .B(n1771), .Z(n1769) );
  XNOR U1704 ( .A(p_input[383]), .B(n1768), .Z(n1771) );
  XOR U1705 ( .A(n1768), .B(p_input[351]), .Z(n1770) );
  XOR U1706 ( .A(n1772), .B(n1773), .Z(n1768) );
  AND U1707 ( .A(n1774), .B(n1775), .Z(n1773) );
  XNOR U1708 ( .A(p_input[382]), .B(n1772), .Z(n1775) );
  XOR U1709 ( .A(n1772), .B(p_input[350]), .Z(n1774) );
  XOR U1710 ( .A(n1776), .B(n1777), .Z(n1772) );
  AND U1711 ( .A(n1778), .B(n1779), .Z(n1777) );
  XNOR U1712 ( .A(p_input[381]), .B(n1776), .Z(n1779) );
  XOR U1713 ( .A(n1776), .B(p_input[349]), .Z(n1778) );
  XOR U1714 ( .A(n1780), .B(n1781), .Z(n1776) );
  AND U1715 ( .A(n1782), .B(n1783), .Z(n1781) );
  XNOR U1716 ( .A(p_input[380]), .B(n1780), .Z(n1783) );
  XOR U1717 ( .A(n1780), .B(p_input[348]), .Z(n1782) );
  XOR U1718 ( .A(n1784), .B(n1785), .Z(n1780) );
  AND U1719 ( .A(n1786), .B(n1787), .Z(n1785) );
  XNOR U1720 ( .A(p_input[379]), .B(n1784), .Z(n1787) );
  XOR U1721 ( .A(n1784), .B(p_input[347]), .Z(n1786) );
  XOR U1722 ( .A(n1788), .B(n1789), .Z(n1784) );
  AND U1723 ( .A(n1790), .B(n1791), .Z(n1789) );
  XNOR U1724 ( .A(p_input[378]), .B(n1788), .Z(n1791) );
  XOR U1725 ( .A(n1788), .B(p_input[346]), .Z(n1790) );
  XOR U1726 ( .A(n1792), .B(n1793), .Z(n1788) );
  AND U1727 ( .A(n1794), .B(n1795), .Z(n1793) );
  XNOR U1728 ( .A(p_input[377]), .B(n1792), .Z(n1795) );
  XOR U1729 ( .A(n1792), .B(p_input[345]), .Z(n1794) );
  XOR U1730 ( .A(n1796), .B(n1797), .Z(n1792) );
  AND U1731 ( .A(n1798), .B(n1799), .Z(n1797) );
  XNOR U1732 ( .A(p_input[376]), .B(n1796), .Z(n1799) );
  XOR U1733 ( .A(n1796), .B(p_input[344]), .Z(n1798) );
  XOR U1734 ( .A(n1800), .B(n1801), .Z(n1796) );
  AND U1735 ( .A(n1802), .B(n1803), .Z(n1801) );
  XNOR U1736 ( .A(p_input[375]), .B(n1800), .Z(n1803) );
  XOR U1737 ( .A(n1800), .B(p_input[343]), .Z(n1802) );
  XOR U1738 ( .A(n1804), .B(n1805), .Z(n1800) );
  AND U1739 ( .A(n1806), .B(n1807), .Z(n1805) );
  XNOR U1740 ( .A(p_input[374]), .B(n1804), .Z(n1807) );
  XOR U1741 ( .A(n1804), .B(p_input[342]), .Z(n1806) );
  XOR U1742 ( .A(n1808), .B(n1809), .Z(n1804) );
  AND U1743 ( .A(n1810), .B(n1811), .Z(n1809) );
  XNOR U1744 ( .A(p_input[373]), .B(n1808), .Z(n1811) );
  XOR U1745 ( .A(n1808), .B(p_input[341]), .Z(n1810) );
  XOR U1746 ( .A(n1812), .B(n1813), .Z(n1808) );
  AND U1747 ( .A(n1814), .B(n1815), .Z(n1813) );
  XNOR U1748 ( .A(p_input[372]), .B(n1812), .Z(n1815) );
  XOR U1749 ( .A(n1812), .B(p_input[340]), .Z(n1814) );
  XOR U1750 ( .A(n1816), .B(n1817), .Z(n1812) );
  AND U1751 ( .A(n1818), .B(n1819), .Z(n1817) );
  XNOR U1752 ( .A(p_input[371]), .B(n1816), .Z(n1819) );
  XOR U1753 ( .A(n1816), .B(p_input[339]), .Z(n1818) );
  XOR U1754 ( .A(n1820), .B(n1821), .Z(n1816) );
  AND U1755 ( .A(n1822), .B(n1823), .Z(n1821) );
  XNOR U1756 ( .A(p_input[370]), .B(n1820), .Z(n1823) );
  XOR U1757 ( .A(n1820), .B(p_input[338]), .Z(n1822) );
  XOR U1758 ( .A(n1824), .B(n1825), .Z(n1820) );
  AND U1759 ( .A(n1826), .B(n1827), .Z(n1825) );
  XNOR U1760 ( .A(p_input[369]), .B(n1824), .Z(n1827) );
  XOR U1761 ( .A(n1824), .B(p_input[337]), .Z(n1826) );
  XOR U1762 ( .A(n1828), .B(n1829), .Z(n1824) );
  AND U1763 ( .A(n1830), .B(n1831), .Z(n1829) );
  XNOR U1764 ( .A(p_input[368]), .B(n1828), .Z(n1831) );
  XOR U1765 ( .A(n1828), .B(p_input[336]), .Z(n1830) );
  XOR U1766 ( .A(n1832), .B(n1833), .Z(n1828) );
  AND U1767 ( .A(n1834), .B(n1835), .Z(n1833) );
  XNOR U1768 ( .A(p_input[367]), .B(n1832), .Z(n1835) );
  XOR U1769 ( .A(n1832), .B(p_input[335]), .Z(n1834) );
  XOR U1770 ( .A(n1836), .B(n1837), .Z(n1832) );
  AND U1771 ( .A(n1838), .B(n1839), .Z(n1837) );
  XNOR U1772 ( .A(p_input[366]), .B(n1836), .Z(n1839) );
  XOR U1773 ( .A(n1836), .B(p_input[334]), .Z(n1838) );
  XOR U1774 ( .A(n1840), .B(n1841), .Z(n1836) );
  AND U1775 ( .A(n1842), .B(n1843), .Z(n1841) );
  XNOR U1776 ( .A(p_input[365]), .B(n1840), .Z(n1843) );
  XOR U1777 ( .A(n1840), .B(p_input[333]), .Z(n1842) );
  XOR U1778 ( .A(n1844), .B(n1845), .Z(n1840) );
  AND U1779 ( .A(n1846), .B(n1847), .Z(n1845) );
  XNOR U1780 ( .A(p_input[364]), .B(n1844), .Z(n1847) );
  XOR U1781 ( .A(n1844), .B(p_input[332]), .Z(n1846) );
  XOR U1782 ( .A(n1848), .B(n1849), .Z(n1844) );
  AND U1783 ( .A(n1850), .B(n1851), .Z(n1849) );
  XNOR U1784 ( .A(p_input[363]), .B(n1848), .Z(n1851) );
  XOR U1785 ( .A(n1848), .B(p_input[331]), .Z(n1850) );
  XOR U1786 ( .A(n1852), .B(n1853), .Z(n1848) );
  AND U1787 ( .A(n1854), .B(n1855), .Z(n1853) );
  XNOR U1788 ( .A(p_input[362]), .B(n1852), .Z(n1855) );
  XOR U1789 ( .A(n1852), .B(p_input[330]), .Z(n1854) );
  XOR U1790 ( .A(n1856), .B(n1857), .Z(n1852) );
  AND U1791 ( .A(n1858), .B(n1859), .Z(n1857) );
  XNOR U1792 ( .A(p_input[361]), .B(n1856), .Z(n1859) );
  XOR U1793 ( .A(n1856), .B(p_input[329]), .Z(n1858) );
  XOR U1794 ( .A(n1860), .B(n1861), .Z(n1856) );
  AND U1795 ( .A(n1862), .B(n1863), .Z(n1861) );
  XNOR U1796 ( .A(p_input[360]), .B(n1860), .Z(n1863) );
  XOR U1797 ( .A(n1860), .B(p_input[328]), .Z(n1862) );
  XOR U1798 ( .A(n1864), .B(n1865), .Z(n1860) );
  AND U1799 ( .A(n1866), .B(n1867), .Z(n1865) );
  XNOR U1800 ( .A(p_input[359]), .B(n1864), .Z(n1867) );
  XOR U1801 ( .A(n1864), .B(p_input[327]), .Z(n1866) );
  XOR U1802 ( .A(n1868), .B(n1869), .Z(n1864) );
  AND U1803 ( .A(n1870), .B(n1871), .Z(n1869) );
  XNOR U1804 ( .A(p_input[358]), .B(n1868), .Z(n1871) );
  XOR U1805 ( .A(n1868), .B(p_input[326]), .Z(n1870) );
  XOR U1806 ( .A(n1872), .B(n1873), .Z(n1868) );
  AND U1807 ( .A(n1874), .B(n1875), .Z(n1873) );
  XNOR U1808 ( .A(p_input[357]), .B(n1872), .Z(n1875) );
  XOR U1809 ( .A(n1872), .B(p_input[325]), .Z(n1874) );
  XOR U1810 ( .A(n1876), .B(n1877), .Z(n1872) );
  AND U1811 ( .A(n1878), .B(n1879), .Z(n1877) );
  XNOR U1812 ( .A(p_input[356]), .B(n1876), .Z(n1879) );
  XOR U1813 ( .A(n1876), .B(p_input[324]), .Z(n1878) );
  XOR U1814 ( .A(n1880), .B(n1881), .Z(n1876) );
  AND U1815 ( .A(n1882), .B(n1883), .Z(n1881) );
  XNOR U1816 ( .A(p_input[355]), .B(n1880), .Z(n1883) );
  XOR U1817 ( .A(n1880), .B(p_input[323]), .Z(n1882) );
  XOR U1818 ( .A(n1884), .B(n1885), .Z(n1880) );
  AND U1819 ( .A(n1886), .B(n1887), .Z(n1885) );
  XNOR U1820 ( .A(p_input[354]), .B(n1884), .Z(n1887) );
  XOR U1821 ( .A(n1884), .B(p_input[322]), .Z(n1886) );
  XNOR U1822 ( .A(n1888), .B(n1889), .Z(n1884) );
  AND U1823 ( .A(n1890), .B(n1891), .Z(n1889) );
  XOR U1824 ( .A(p_input[353]), .B(n1888), .Z(n1891) );
  XNOR U1825 ( .A(p_input[321]), .B(n1888), .Z(n1890) );
  AND U1826 ( .A(p_input[352]), .B(n1892), .Z(n1888) );
  IV U1827 ( .A(p_input[320]), .Z(n1892) );
  XNOR U1828 ( .A(p_input[256]), .B(n1893), .Z(n1486) );
  AND U1829 ( .A(n171), .B(n1894), .Z(n1893) );
  XOR U1830 ( .A(p_input[288]), .B(p_input[256]), .Z(n1894) );
  XOR U1831 ( .A(n1895), .B(n1896), .Z(n171) );
  AND U1832 ( .A(n1897), .B(n1898), .Z(n1896) );
  XNOR U1833 ( .A(p_input[319]), .B(n1895), .Z(n1898) );
  XOR U1834 ( .A(n1895), .B(p_input[287]), .Z(n1897) );
  XOR U1835 ( .A(n1899), .B(n1900), .Z(n1895) );
  AND U1836 ( .A(n1901), .B(n1902), .Z(n1900) );
  XNOR U1837 ( .A(p_input[318]), .B(n1899), .Z(n1902) );
  XNOR U1838 ( .A(n1899), .B(n1501), .Z(n1901) );
  IV U1839 ( .A(p_input[286]), .Z(n1501) );
  XOR U1840 ( .A(n1903), .B(n1904), .Z(n1899) );
  AND U1841 ( .A(n1905), .B(n1906), .Z(n1904) );
  XNOR U1842 ( .A(p_input[317]), .B(n1903), .Z(n1906) );
  XNOR U1843 ( .A(n1903), .B(n1510), .Z(n1905) );
  IV U1844 ( .A(p_input[285]), .Z(n1510) );
  XOR U1845 ( .A(n1907), .B(n1908), .Z(n1903) );
  AND U1846 ( .A(n1909), .B(n1910), .Z(n1908) );
  XNOR U1847 ( .A(p_input[316]), .B(n1907), .Z(n1910) );
  XNOR U1848 ( .A(n1907), .B(n1519), .Z(n1909) );
  IV U1849 ( .A(p_input[284]), .Z(n1519) );
  XOR U1850 ( .A(n1911), .B(n1912), .Z(n1907) );
  AND U1851 ( .A(n1913), .B(n1914), .Z(n1912) );
  XNOR U1852 ( .A(p_input[315]), .B(n1911), .Z(n1914) );
  XNOR U1853 ( .A(n1911), .B(n1528), .Z(n1913) );
  IV U1854 ( .A(p_input[283]), .Z(n1528) );
  XOR U1855 ( .A(n1915), .B(n1916), .Z(n1911) );
  AND U1856 ( .A(n1917), .B(n1918), .Z(n1916) );
  XNOR U1857 ( .A(p_input[314]), .B(n1915), .Z(n1918) );
  XNOR U1858 ( .A(n1915), .B(n1537), .Z(n1917) );
  IV U1859 ( .A(p_input[282]), .Z(n1537) );
  XOR U1860 ( .A(n1919), .B(n1920), .Z(n1915) );
  AND U1861 ( .A(n1921), .B(n1922), .Z(n1920) );
  XNOR U1862 ( .A(p_input[313]), .B(n1919), .Z(n1922) );
  XNOR U1863 ( .A(n1919), .B(n1546), .Z(n1921) );
  IV U1864 ( .A(p_input[281]), .Z(n1546) );
  XOR U1865 ( .A(n1923), .B(n1924), .Z(n1919) );
  AND U1866 ( .A(n1925), .B(n1926), .Z(n1924) );
  XNOR U1867 ( .A(p_input[312]), .B(n1923), .Z(n1926) );
  XNOR U1868 ( .A(n1923), .B(n1555), .Z(n1925) );
  IV U1869 ( .A(p_input[280]), .Z(n1555) );
  XOR U1870 ( .A(n1927), .B(n1928), .Z(n1923) );
  AND U1871 ( .A(n1929), .B(n1930), .Z(n1928) );
  XNOR U1872 ( .A(p_input[311]), .B(n1927), .Z(n1930) );
  XNOR U1873 ( .A(n1927), .B(n1564), .Z(n1929) );
  IV U1874 ( .A(p_input[279]), .Z(n1564) );
  XOR U1875 ( .A(n1931), .B(n1932), .Z(n1927) );
  AND U1876 ( .A(n1933), .B(n1934), .Z(n1932) );
  XNOR U1877 ( .A(p_input[310]), .B(n1931), .Z(n1934) );
  XNOR U1878 ( .A(n1931), .B(n1573), .Z(n1933) );
  IV U1879 ( .A(p_input[278]), .Z(n1573) );
  XOR U1880 ( .A(n1935), .B(n1936), .Z(n1931) );
  AND U1881 ( .A(n1937), .B(n1938), .Z(n1936) );
  XNOR U1882 ( .A(p_input[309]), .B(n1935), .Z(n1938) );
  XNOR U1883 ( .A(n1935), .B(n1582), .Z(n1937) );
  IV U1884 ( .A(p_input[277]), .Z(n1582) );
  XOR U1885 ( .A(n1939), .B(n1940), .Z(n1935) );
  AND U1886 ( .A(n1941), .B(n1942), .Z(n1940) );
  XNOR U1887 ( .A(p_input[308]), .B(n1939), .Z(n1942) );
  XNOR U1888 ( .A(n1939), .B(n1591), .Z(n1941) );
  IV U1889 ( .A(p_input[276]), .Z(n1591) );
  XOR U1890 ( .A(n1943), .B(n1944), .Z(n1939) );
  AND U1891 ( .A(n1945), .B(n1946), .Z(n1944) );
  XNOR U1892 ( .A(p_input[307]), .B(n1943), .Z(n1946) );
  XNOR U1893 ( .A(n1943), .B(n1600), .Z(n1945) );
  IV U1894 ( .A(p_input[275]), .Z(n1600) );
  XOR U1895 ( .A(n1947), .B(n1948), .Z(n1943) );
  AND U1896 ( .A(n1949), .B(n1950), .Z(n1948) );
  XNOR U1897 ( .A(p_input[306]), .B(n1947), .Z(n1950) );
  XNOR U1898 ( .A(n1947), .B(n1609), .Z(n1949) );
  IV U1899 ( .A(p_input[274]), .Z(n1609) );
  XOR U1900 ( .A(n1951), .B(n1952), .Z(n1947) );
  AND U1901 ( .A(n1953), .B(n1954), .Z(n1952) );
  XNOR U1902 ( .A(p_input[305]), .B(n1951), .Z(n1954) );
  XNOR U1903 ( .A(n1951), .B(n1618), .Z(n1953) );
  IV U1904 ( .A(p_input[273]), .Z(n1618) );
  XOR U1905 ( .A(n1955), .B(n1956), .Z(n1951) );
  AND U1906 ( .A(n1957), .B(n1958), .Z(n1956) );
  XNOR U1907 ( .A(p_input[304]), .B(n1955), .Z(n1958) );
  XNOR U1908 ( .A(n1955), .B(n1627), .Z(n1957) );
  IV U1909 ( .A(p_input[272]), .Z(n1627) );
  XOR U1910 ( .A(n1959), .B(n1960), .Z(n1955) );
  AND U1911 ( .A(n1961), .B(n1962), .Z(n1960) );
  XNOR U1912 ( .A(p_input[303]), .B(n1959), .Z(n1962) );
  XNOR U1913 ( .A(n1959), .B(n1636), .Z(n1961) );
  IV U1914 ( .A(p_input[271]), .Z(n1636) );
  XOR U1915 ( .A(n1963), .B(n1964), .Z(n1959) );
  AND U1916 ( .A(n1965), .B(n1966), .Z(n1964) );
  XNOR U1917 ( .A(p_input[302]), .B(n1963), .Z(n1966) );
  XNOR U1918 ( .A(n1963), .B(n1645), .Z(n1965) );
  IV U1919 ( .A(p_input[270]), .Z(n1645) );
  XOR U1920 ( .A(n1967), .B(n1968), .Z(n1963) );
  AND U1921 ( .A(n1969), .B(n1970), .Z(n1968) );
  XNOR U1922 ( .A(p_input[301]), .B(n1967), .Z(n1970) );
  XNOR U1923 ( .A(n1967), .B(n1654), .Z(n1969) );
  IV U1924 ( .A(p_input[269]), .Z(n1654) );
  XOR U1925 ( .A(n1971), .B(n1972), .Z(n1967) );
  AND U1926 ( .A(n1973), .B(n1974), .Z(n1972) );
  XNOR U1927 ( .A(p_input[300]), .B(n1971), .Z(n1974) );
  XNOR U1928 ( .A(n1971), .B(n1663), .Z(n1973) );
  IV U1929 ( .A(p_input[268]), .Z(n1663) );
  XOR U1930 ( .A(n1975), .B(n1976), .Z(n1971) );
  AND U1931 ( .A(n1977), .B(n1978), .Z(n1976) );
  XNOR U1932 ( .A(p_input[299]), .B(n1975), .Z(n1978) );
  XNOR U1933 ( .A(n1975), .B(n1672), .Z(n1977) );
  IV U1934 ( .A(p_input[267]), .Z(n1672) );
  XOR U1935 ( .A(n1979), .B(n1980), .Z(n1975) );
  AND U1936 ( .A(n1981), .B(n1982), .Z(n1980) );
  XNOR U1937 ( .A(p_input[298]), .B(n1979), .Z(n1982) );
  XNOR U1938 ( .A(n1979), .B(n1681), .Z(n1981) );
  IV U1939 ( .A(p_input[266]), .Z(n1681) );
  XOR U1940 ( .A(n1983), .B(n1984), .Z(n1979) );
  AND U1941 ( .A(n1985), .B(n1986), .Z(n1984) );
  XNOR U1942 ( .A(p_input[297]), .B(n1983), .Z(n1986) );
  XNOR U1943 ( .A(n1983), .B(n1690), .Z(n1985) );
  IV U1944 ( .A(p_input[265]), .Z(n1690) );
  XOR U1945 ( .A(n1987), .B(n1988), .Z(n1983) );
  AND U1946 ( .A(n1989), .B(n1990), .Z(n1988) );
  XNOR U1947 ( .A(p_input[296]), .B(n1987), .Z(n1990) );
  XNOR U1948 ( .A(n1987), .B(n1699), .Z(n1989) );
  IV U1949 ( .A(p_input[264]), .Z(n1699) );
  XOR U1950 ( .A(n1991), .B(n1992), .Z(n1987) );
  AND U1951 ( .A(n1993), .B(n1994), .Z(n1992) );
  XNOR U1952 ( .A(p_input[295]), .B(n1991), .Z(n1994) );
  XNOR U1953 ( .A(n1991), .B(n1708), .Z(n1993) );
  IV U1954 ( .A(p_input[263]), .Z(n1708) );
  XOR U1955 ( .A(n1995), .B(n1996), .Z(n1991) );
  AND U1956 ( .A(n1997), .B(n1998), .Z(n1996) );
  XNOR U1957 ( .A(p_input[294]), .B(n1995), .Z(n1998) );
  XNOR U1958 ( .A(n1995), .B(n1717), .Z(n1997) );
  IV U1959 ( .A(p_input[262]), .Z(n1717) );
  XOR U1960 ( .A(n1999), .B(n2000), .Z(n1995) );
  AND U1961 ( .A(n2001), .B(n2002), .Z(n2000) );
  XNOR U1962 ( .A(p_input[293]), .B(n1999), .Z(n2002) );
  XNOR U1963 ( .A(n1999), .B(n1726), .Z(n2001) );
  IV U1964 ( .A(p_input[261]), .Z(n1726) );
  XOR U1965 ( .A(n2003), .B(n2004), .Z(n1999) );
  AND U1966 ( .A(n2005), .B(n2006), .Z(n2004) );
  XNOR U1967 ( .A(p_input[292]), .B(n2003), .Z(n2006) );
  XNOR U1968 ( .A(n2003), .B(n1735), .Z(n2005) );
  IV U1969 ( .A(p_input[260]), .Z(n1735) );
  XOR U1970 ( .A(n2007), .B(n2008), .Z(n2003) );
  AND U1971 ( .A(n2009), .B(n2010), .Z(n2008) );
  XNOR U1972 ( .A(p_input[291]), .B(n2007), .Z(n2010) );
  XNOR U1973 ( .A(n2007), .B(n1744), .Z(n2009) );
  IV U1974 ( .A(p_input[259]), .Z(n1744) );
  XOR U1975 ( .A(n2011), .B(n2012), .Z(n2007) );
  AND U1976 ( .A(n2013), .B(n2014), .Z(n2012) );
  XNOR U1977 ( .A(p_input[290]), .B(n2011), .Z(n2014) );
  XNOR U1978 ( .A(n2011), .B(n1753), .Z(n2013) );
  IV U1979 ( .A(p_input[258]), .Z(n1753) );
  XNOR U1980 ( .A(n2015), .B(n2016), .Z(n2011) );
  AND U1981 ( .A(n2017), .B(n2018), .Z(n2016) );
  XOR U1982 ( .A(p_input[289]), .B(n2015), .Z(n2018) );
  XNOR U1983 ( .A(p_input[257]), .B(n2015), .Z(n2017) );
  AND U1984 ( .A(p_input[288]), .B(n2019), .Z(n2015) );
  IV U1985 ( .A(p_input[256]), .Z(n2019) );
  XOR U1986 ( .A(n2020), .B(n2021), .Z(n26) );
  AND U1987 ( .A(n195), .B(n2022), .Z(n2021) );
  XNOR U1988 ( .A(n2023), .B(n2020), .Z(n2022) );
  XOR U1989 ( .A(n2024), .B(n2025), .Z(n195) );
  AND U1990 ( .A(n2026), .B(n2027), .Z(n2025) );
  XOR U1991 ( .A(n2024), .B(n214), .Z(n2027) );
  XNOR U1992 ( .A(n2028), .B(n2029), .Z(n214) );
  AND U1993 ( .A(n2030), .B(n186), .Z(n2029) );
  AND U1994 ( .A(n2028), .B(n2031), .Z(n2030) );
  XNOR U1995 ( .A(n211), .B(n2024), .Z(n2026) );
  XOR U1996 ( .A(n2032), .B(n2033), .Z(n211) );
  AND U1997 ( .A(n2034), .B(n183), .Z(n2033) );
  NOR U1998 ( .A(n2032), .B(n2035), .Z(n2034) );
  XOR U1999 ( .A(n2036), .B(n2037), .Z(n2024) );
  AND U2000 ( .A(n2038), .B(n2039), .Z(n2037) );
  XOR U2001 ( .A(n2036), .B(n226), .Z(n2039) );
  XOR U2002 ( .A(n2040), .B(n2041), .Z(n226) );
  AND U2003 ( .A(n186), .B(n2042), .Z(n2041) );
  XOR U2004 ( .A(n2043), .B(n2040), .Z(n2042) );
  XNOR U2005 ( .A(n223), .B(n2036), .Z(n2038) );
  XOR U2006 ( .A(n2044), .B(n2045), .Z(n223) );
  AND U2007 ( .A(n183), .B(n2046), .Z(n2045) );
  XOR U2008 ( .A(n2047), .B(n2044), .Z(n2046) );
  XOR U2009 ( .A(n2048), .B(n2049), .Z(n2036) );
  AND U2010 ( .A(n2050), .B(n2051), .Z(n2049) );
  XOR U2011 ( .A(n2048), .B(n238), .Z(n2051) );
  XOR U2012 ( .A(n2052), .B(n2053), .Z(n238) );
  AND U2013 ( .A(n186), .B(n2054), .Z(n2053) );
  XOR U2014 ( .A(n2055), .B(n2052), .Z(n2054) );
  XNOR U2015 ( .A(n235), .B(n2048), .Z(n2050) );
  XOR U2016 ( .A(n2056), .B(n2057), .Z(n235) );
  AND U2017 ( .A(n183), .B(n2058), .Z(n2057) );
  XOR U2018 ( .A(n2059), .B(n2056), .Z(n2058) );
  XOR U2019 ( .A(n2060), .B(n2061), .Z(n2048) );
  AND U2020 ( .A(n2062), .B(n2063), .Z(n2061) );
  XOR U2021 ( .A(n2060), .B(n250), .Z(n2063) );
  XOR U2022 ( .A(n2064), .B(n2065), .Z(n250) );
  AND U2023 ( .A(n186), .B(n2066), .Z(n2065) );
  XOR U2024 ( .A(n2067), .B(n2064), .Z(n2066) );
  XNOR U2025 ( .A(n247), .B(n2060), .Z(n2062) );
  XOR U2026 ( .A(n2068), .B(n2069), .Z(n247) );
  AND U2027 ( .A(n183), .B(n2070), .Z(n2069) );
  XOR U2028 ( .A(n2071), .B(n2068), .Z(n2070) );
  XOR U2029 ( .A(n2072), .B(n2073), .Z(n2060) );
  AND U2030 ( .A(n2074), .B(n2075), .Z(n2073) );
  XOR U2031 ( .A(n2072), .B(n262), .Z(n2075) );
  XOR U2032 ( .A(n2076), .B(n2077), .Z(n262) );
  AND U2033 ( .A(n186), .B(n2078), .Z(n2077) );
  XOR U2034 ( .A(n2079), .B(n2076), .Z(n2078) );
  XNOR U2035 ( .A(n259), .B(n2072), .Z(n2074) );
  XOR U2036 ( .A(n2080), .B(n2081), .Z(n259) );
  AND U2037 ( .A(n183), .B(n2082), .Z(n2081) );
  XOR U2038 ( .A(n2083), .B(n2080), .Z(n2082) );
  XOR U2039 ( .A(n2084), .B(n2085), .Z(n2072) );
  AND U2040 ( .A(n2086), .B(n2087), .Z(n2085) );
  XOR U2041 ( .A(n2084), .B(n274), .Z(n2087) );
  XOR U2042 ( .A(n2088), .B(n2089), .Z(n274) );
  AND U2043 ( .A(n186), .B(n2090), .Z(n2089) );
  XOR U2044 ( .A(n2091), .B(n2088), .Z(n2090) );
  XNOR U2045 ( .A(n271), .B(n2084), .Z(n2086) );
  XOR U2046 ( .A(n2092), .B(n2093), .Z(n271) );
  AND U2047 ( .A(n183), .B(n2094), .Z(n2093) );
  XOR U2048 ( .A(n2095), .B(n2092), .Z(n2094) );
  XOR U2049 ( .A(n2096), .B(n2097), .Z(n2084) );
  AND U2050 ( .A(n2098), .B(n2099), .Z(n2097) );
  XOR U2051 ( .A(n2096), .B(n286), .Z(n2099) );
  XOR U2052 ( .A(n2100), .B(n2101), .Z(n286) );
  AND U2053 ( .A(n186), .B(n2102), .Z(n2101) );
  XOR U2054 ( .A(n2103), .B(n2100), .Z(n2102) );
  XNOR U2055 ( .A(n283), .B(n2096), .Z(n2098) );
  XOR U2056 ( .A(n2104), .B(n2105), .Z(n283) );
  AND U2057 ( .A(n183), .B(n2106), .Z(n2105) );
  XOR U2058 ( .A(n2107), .B(n2104), .Z(n2106) );
  XOR U2059 ( .A(n2108), .B(n2109), .Z(n2096) );
  AND U2060 ( .A(n2110), .B(n2111), .Z(n2109) );
  XOR U2061 ( .A(n2108), .B(n298), .Z(n2111) );
  XOR U2062 ( .A(n2112), .B(n2113), .Z(n298) );
  AND U2063 ( .A(n186), .B(n2114), .Z(n2113) );
  XOR U2064 ( .A(n2115), .B(n2112), .Z(n2114) );
  XNOR U2065 ( .A(n295), .B(n2108), .Z(n2110) );
  XOR U2066 ( .A(n2116), .B(n2117), .Z(n295) );
  AND U2067 ( .A(n183), .B(n2118), .Z(n2117) );
  XOR U2068 ( .A(n2119), .B(n2116), .Z(n2118) );
  XOR U2069 ( .A(n2120), .B(n2121), .Z(n2108) );
  AND U2070 ( .A(n2122), .B(n2123), .Z(n2121) );
  XOR U2071 ( .A(n2120), .B(n310), .Z(n2123) );
  XOR U2072 ( .A(n2124), .B(n2125), .Z(n310) );
  AND U2073 ( .A(n186), .B(n2126), .Z(n2125) );
  XOR U2074 ( .A(n2127), .B(n2124), .Z(n2126) );
  XNOR U2075 ( .A(n307), .B(n2120), .Z(n2122) );
  XOR U2076 ( .A(n2128), .B(n2129), .Z(n307) );
  AND U2077 ( .A(n183), .B(n2130), .Z(n2129) );
  XOR U2078 ( .A(n2131), .B(n2128), .Z(n2130) );
  XOR U2079 ( .A(n2132), .B(n2133), .Z(n2120) );
  AND U2080 ( .A(n2134), .B(n2135), .Z(n2133) );
  XOR U2081 ( .A(n2132), .B(n322), .Z(n2135) );
  XOR U2082 ( .A(n2136), .B(n2137), .Z(n322) );
  AND U2083 ( .A(n186), .B(n2138), .Z(n2137) );
  XOR U2084 ( .A(n2139), .B(n2136), .Z(n2138) );
  XNOR U2085 ( .A(n319), .B(n2132), .Z(n2134) );
  XOR U2086 ( .A(n2140), .B(n2141), .Z(n319) );
  AND U2087 ( .A(n183), .B(n2142), .Z(n2141) );
  XOR U2088 ( .A(n2143), .B(n2140), .Z(n2142) );
  XOR U2089 ( .A(n2144), .B(n2145), .Z(n2132) );
  AND U2090 ( .A(n2146), .B(n2147), .Z(n2145) );
  XOR U2091 ( .A(n2144), .B(n334), .Z(n2147) );
  XOR U2092 ( .A(n2148), .B(n2149), .Z(n334) );
  AND U2093 ( .A(n186), .B(n2150), .Z(n2149) );
  XOR U2094 ( .A(n2151), .B(n2148), .Z(n2150) );
  XNOR U2095 ( .A(n331), .B(n2144), .Z(n2146) );
  XOR U2096 ( .A(n2152), .B(n2153), .Z(n331) );
  AND U2097 ( .A(n183), .B(n2154), .Z(n2153) );
  XOR U2098 ( .A(n2155), .B(n2152), .Z(n2154) );
  XOR U2099 ( .A(n2156), .B(n2157), .Z(n2144) );
  AND U2100 ( .A(n2158), .B(n2159), .Z(n2157) );
  XOR U2101 ( .A(n2156), .B(n346), .Z(n2159) );
  XOR U2102 ( .A(n2160), .B(n2161), .Z(n346) );
  AND U2103 ( .A(n186), .B(n2162), .Z(n2161) );
  XOR U2104 ( .A(n2163), .B(n2160), .Z(n2162) );
  XNOR U2105 ( .A(n343), .B(n2156), .Z(n2158) );
  XOR U2106 ( .A(n2164), .B(n2165), .Z(n343) );
  AND U2107 ( .A(n183), .B(n2166), .Z(n2165) );
  XOR U2108 ( .A(n2167), .B(n2164), .Z(n2166) );
  XOR U2109 ( .A(n2168), .B(n2169), .Z(n2156) );
  AND U2110 ( .A(n2170), .B(n2171), .Z(n2169) );
  XOR U2111 ( .A(n2168), .B(n358), .Z(n2171) );
  XOR U2112 ( .A(n2172), .B(n2173), .Z(n358) );
  AND U2113 ( .A(n186), .B(n2174), .Z(n2173) );
  XOR U2114 ( .A(n2175), .B(n2172), .Z(n2174) );
  XNOR U2115 ( .A(n355), .B(n2168), .Z(n2170) );
  XOR U2116 ( .A(n2176), .B(n2177), .Z(n355) );
  AND U2117 ( .A(n183), .B(n2178), .Z(n2177) );
  XOR U2118 ( .A(n2179), .B(n2176), .Z(n2178) );
  XOR U2119 ( .A(n2180), .B(n2181), .Z(n2168) );
  AND U2120 ( .A(n2182), .B(n2183), .Z(n2181) );
  XOR U2121 ( .A(n2180), .B(n370), .Z(n2183) );
  XOR U2122 ( .A(n2184), .B(n2185), .Z(n370) );
  AND U2123 ( .A(n186), .B(n2186), .Z(n2185) );
  XOR U2124 ( .A(n2187), .B(n2184), .Z(n2186) );
  XNOR U2125 ( .A(n367), .B(n2180), .Z(n2182) );
  XOR U2126 ( .A(n2188), .B(n2189), .Z(n367) );
  AND U2127 ( .A(n183), .B(n2190), .Z(n2189) );
  XOR U2128 ( .A(n2191), .B(n2188), .Z(n2190) );
  XOR U2129 ( .A(n2192), .B(n2193), .Z(n2180) );
  AND U2130 ( .A(n2194), .B(n2195), .Z(n2193) );
  XOR U2131 ( .A(n2192), .B(n382), .Z(n2195) );
  XOR U2132 ( .A(n2196), .B(n2197), .Z(n382) );
  AND U2133 ( .A(n186), .B(n2198), .Z(n2197) );
  XOR U2134 ( .A(n2199), .B(n2196), .Z(n2198) );
  XNOR U2135 ( .A(n379), .B(n2192), .Z(n2194) );
  XOR U2136 ( .A(n2200), .B(n2201), .Z(n379) );
  AND U2137 ( .A(n183), .B(n2202), .Z(n2201) );
  XOR U2138 ( .A(n2203), .B(n2200), .Z(n2202) );
  XOR U2139 ( .A(n2204), .B(n2205), .Z(n2192) );
  AND U2140 ( .A(n2206), .B(n2207), .Z(n2205) );
  XOR U2141 ( .A(n2204), .B(n394), .Z(n2207) );
  XOR U2142 ( .A(n2208), .B(n2209), .Z(n394) );
  AND U2143 ( .A(n186), .B(n2210), .Z(n2209) );
  XOR U2144 ( .A(n2211), .B(n2208), .Z(n2210) );
  XNOR U2145 ( .A(n391), .B(n2204), .Z(n2206) );
  XOR U2146 ( .A(n2212), .B(n2213), .Z(n391) );
  AND U2147 ( .A(n183), .B(n2214), .Z(n2213) );
  XOR U2148 ( .A(n2215), .B(n2212), .Z(n2214) );
  XOR U2149 ( .A(n2216), .B(n2217), .Z(n2204) );
  AND U2150 ( .A(n2218), .B(n2219), .Z(n2217) );
  XOR U2151 ( .A(n2216), .B(n406), .Z(n2219) );
  XOR U2152 ( .A(n2220), .B(n2221), .Z(n406) );
  AND U2153 ( .A(n186), .B(n2222), .Z(n2221) );
  XOR U2154 ( .A(n2223), .B(n2220), .Z(n2222) );
  XNOR U2155 ( .A(n403), .B(n2216), .Z(n2218) );
  XOR U2156 ( .A(n2224), .B(n2225), .Z(n403) );
  AND U2157 ( .A(n183), .B(n2226), .Z(n2225) );
  XOR U2158 ( .A(n2227), .B(n2224), .Z(n2226) );
  XOR U2159 ( .A(n2228), .B(n2229), .Z(n2216) );
  AND U2160 ( .A(n2230), .B(n2231), .Z(n2229) );
  XOR U2161 ( .A(n2228), .B(n418), .Z(n2231) );
  XOR U2162 ( .A(n2232), .B(n2233), .Z(n418) );
  AND U2163 ( .A(n186), .B(n2234), .Z(n2233) );
  XOR U2164 ( .A(n2235), .B(n2232), .Z(n2234) );
  XNOR U2165 ( .A(n415), .B(n2228), .Z(n2230) );
  XOR U2166 ( .A(n2236), .B(n2237), .Z(n415) );
  AND U2167 ( .A(n183), .B(n2238), .Z(n2237) );
  XOR U2168 ( .A(n2239), .B(n2236), .Z(n2238) );
  XOR U2169 ( .A(n2240), .B(n2241), .Z(n2228) );
  AND U2170 ( .A(n2242), .B(n2243), .Z(n2241) );
  XOR U2171 ( .A(n2240), .B(n430), .Z(n2243) );
  XOR U2172 ( .A(n2244), .B(n2245), .Z(n430) );
  AND U2173 ( .A(n186), .B(n2246), .Z(n2245) );
  XOR U2174 ( .A(n2247), .B(n2244), .Z(n2246) );
  XNOR U2175 ( .A(n427), .B(n2240), .Z(n2242) );
  XOR U2176 ( .A(n2248), .B(n2249), .Z(n427) );
  AND U2177 ( .A(n183), .B(n2250), .Z(n2249) );
  XOR U2178 ( .A(n2251), .B(n2248), .Z(n2250) );
  XOR U2179 ( .A(n2252), .B(n2253), .Z(n2240) );
  AND U2180 ( .A(n2254), .B(n2255), .Z(n2253) );
  XOR U2181 ( .A(n2252), .B(n442), .Z(n2255) );
  XOR U2182 ( .A(n2256), .B(n2257), .Z(n442) );
  AND U2183 ( .A(n186), .B(n2258), .Z(n2257) );
  XOR U2184 ( .A(n2259), .B(n2256), .Z(n2258) );
  XNOR U2185 ( .A(n439), .B(n2252), .Z(n2254) );
  XOR U2186 ( .A(n2260), .B(n2261), .Z(n439) );
  AND U2187 ( .A(n183), .B(n2262), .Z(n2261) );
  XOR U2188 ( .A(n2263), .B(n2260), .Z(n2262) );
  XOR U2189 ( .A(n2264), .B(n2265), .Z(n2252) );
  AND U2190 ( .A(n2266), .B(n2267), .Z(n2265) );
  XOR U2191 ( .A(n2264), .B(n454), .Z(n2267) );
  XOR U2192 ( .A(n2268), .B(n2269), .Z(n454) );
  AND U2193 ( .A(n186), .B(n2270), .Z(n2269) );
  XOR U2194 ( .A(n2271), .B(n2268), .Z(n2270) );
  XNOR U2195 ( .A(n451), .B(n2264), .Z(n2266) );
  XOR U2196 ( .A(n2272), .B(n2273), .Z(n451) );
  AND U2197 ( .A(n183), .B(n2274), .Z(n2273) );
  XOR U2198 ( .A(n2275), .B(n2272), .Z(n2274) );
  XOR U2199 ( .A(n2276), .B(n2277), .Z(n2264) );
  AND U2200 ( .A(n2278), .B(n2279), .Z(n2277) );
  XOR U2201 ( .A(n2276), .B(n466), .Z(n2279) );
  XOR U2202 ( .A(n2280), .B(n2281), .Z(n466) );
  AND U2203 ( .A(n186), .B(n2282), .Z(n2281) );
  XOR U2204 ( .A(n2283), .B(n2280), .Z(n2282) );
  XNOR U2205 ( .A(n463), .B(n2276), .Z(n2278) );
  XOR U2206 ( .A(n2284), .B(n2285), .Z(n463) );
  AND U2207 ( .A(n183), .B(n2286), .Z(n2285) );
  XOR U2208 ( .A(n2287), .B(n2284), .Z(n2286) );
  XOR U2209 ( .A(n2288), .B(n2289), .Z(n2276) );
  AND U2210 ( .A(n2290), .B(n2291), .Z(n2289) );
  XOR U2211 ( .A(n2288), .B(n478), .Z(n2291) );
  XOR U2212 ( .A(n2292), .B(n2293), .Z(n478) );
  AND U2213 ( .A(n186), .B(n2294), .Z(n2293) );
  XOR U2214 ( .A(n2295), .B(n2292), .Z(n2294) );
  XNOR U2215 ( .A(n475), .B(n2288), .Z(n2290) );
  XOR U2216 ( .A(n2296), .B(n2297), .Z(n475) );
  AND U2217 ( .A(n183), .B(n2298), .Z(n2297) );
  XOR U2218 ( .A(n2299), .B(n2296), .Z(n2298) );
  XOR U2219 ( .A(n2300), .B(n2301), .Z(n2288) );
  AND U2220 ( .A(n2302), .B(n2303), .Z(n2301) );
  XOR U2221 ( .A(n2300), .B(n490), .Z(n2303) );
  XOR U2222 ( .A(n2304), .B(n2305), .Z(n490) );
  AND U2223 ( .A(n186), .B(n2306), .Z(n2305) );
  XOR U2224 ( .A(n2307), .B(n2304), .Z(n2306) );
  XNOR U2225 ( .A(n487), .B(n2300), .Z(n2302) );
  XOR U2226 ( .A(n2308), .B(n2309), .Z(n487) );
  AND U2227 ( .A(n183), .B(n2310), .Z(n2309) );
  XOR U2228 ( .A(n2311), .B(n2308), .Z(n2310) );
  XOR U2229 ( .A(n2312), .B(n2313), .Z(n2300) );
  AND U2230 ( .A(n2314), .B(n2315), .Z(n2313) );
  XOR U2231 ( .A(n2312), .B(n502), .Z(n2315) );
  XOR U2232 ( .A(n2316), .B(n2317), .Z(n502) );
  AND U2233 ( .A(n186), .B(n2318), .Z(n2317) );
  XOR U2234 ( .A(n2319), .B(n2316), .Z(n2318) );
  XNOR U2235 ( .A(n499), .B(n2312), .Z(n2314) );
  XOR U2236 ( .A(n2320), .B(n2321), .Z(n499) );
  AND U2237 ( .A(n183), .B(n2322), .Z(n2321) );
  XOR U2238 ( .A(n2323), .B(n2320), .Z(n2322) );
  XOR U2239 ( .A(n2324), .B(n2325), .Z(n2312) );
  AND U2240 ( .A(n2326), .B(n2327), .Z(n2325) );
  XOR U2241 ( .A(n2324), .B(n514), .Z(n2327) );
  XOR U2242 ( .A(n2328), .B(n2329), .Z(n514) );
  AND U2243 ( .A(n186), .B(n2330), .Z(n2329) );
  XOR U2244 ( .A(n2331), .B(n2328), .Z(n2330) );
  XNOR U2245 ( .A(n511), .B(n2324), .Z(n2326) );
  XOR U2246 ( .A(n2332), .B(n2333), .Z(n511) );
  AND U2247 ( .A(n183), .B(n2334), .Z(n2333) );
  XOR U2248 ( .A(n2335), .B(n2332), .Z(n2334) );
  XOR U2249 ( .A(n2336), .B(n2337), .Z(n2324) );
  AND U2250 ( .A(n2338), .B(n2339), .Z(n2337) );
  XOR U2251 ( .A(n526), .B(n2336), .Z(n2339) );
  XOR U2252 ( .A(n2340), .B(n2341), .Z(n526) );
  AND U2253 ( .A(n186), .B(n2342), .Z(n2341) );
  XOR U2254 ( .A(n2340), .B(n2343), .Z(n2342) );
  XNOR U2255 ( .A(n2336), .B(n523), .Z(n2338) );
  XOR U2256 ( .A(n2344), .B(n2345), .Z(n523) );
  AND U2257 ( .A(n183), .B(n2346), .Z(n2345) );
  XOR U2258 ( .A(n2344), .B(n2347), .Z(n2346) );
  XOR U2259 ( .A(n2348), .B(n2349), .Z(n2336) );
  AND U2260 ( .A(n2350), .B(n2351), .Z(n2349) );
  XOR U2261 ( .A(n2348), .B(n538), .Z(n2351) );
  XOR U2262 ( .A(n2352), .B(n2353), .Z(n538) );
  AND U2263 ( .A(n186), .B(n2354), .Z(n2353) );
  XOR U2264 ( .A(n2355), .B(n2352), .Z(n2354) );
  XNOR U2265 ( .A(n535), .B(n2348), .Z(n2350) );
  XOR U2266 ( .A(n2356), .B(n2357), .Z(n535) );
  AND U2267 ( .A(n183), .B(n2358), .Z(n2357) );
  XOR U2268 ( .A(n2359), .B(n2356), .Z(n2358) );
  XOR U2269 ( .A(n2360), .B(n2361), .Z(n2348) );
  AND U2270 ( .A(n2362), .B(n2363), .Z(n2361) );
  XOR U2271 ( .A(n2360), .B(n550), .Z(n2363) );
  XOR U2272 ( .A(n2364), .B(n2365), .Z(n550) );
  AND U2273 ( .A(n186), .B(n2366), .Z(n2365) );
  XOR U2274 ( .A(n2367), .B(n2364), .Z(n2366) );
  XNOR U2275 ( .A(n547), .B(n2360), .Z(n2362) );
  XOR U2276 ( .A(n2368), .B(n2369), .Z(n547) );
  AND U2277 ( .A(n183), .B(n2370), .Z(n2369) );
  XOR U2278 ( .A(n2371), .B(n2368), .Z(n2370) );
  XOR U2279 ( .A(n2372), .B(n2373), .Z(n2360) );
  AND U2280 ( .A(n2374), .B(n2375), .Z(n2373) );
  XOR U2281 ( .A(n2372), .B(n562), .Z(n2375) );
  XOR U2282 ( .A(n2376), .B(n2377), .Z(n562) );
  AND U2283 ( .A(n186), .B(n2378), .Z(n2377) );
  XOR U2284 ( .A(n2379), .B(n2376), .Z(n2378) );
  XNOR U2285 ( .A(n559), .B(n2372), .Z(n2374) );
  XOR U2286 ( .A(n2380), .B(n2381), .Z(n559) );
  AND U2287 ( .A(n183), .B(n2382), .Z(n2381) );
  XOR U2288 ( .A(n2383), .B(n2380), .Z(n2382) );
  XOR U2289 ( .A(n2384), .B(n2385), .Z(n2372) );
  AND U2290 ( .A(n2386), .B(n2387), .Z(n2385) );
  XNOR U2291 ( .A(n2388), .B(n574), .Z(n2387) );
  XOR U2292 ( .A(n2389), .B(n2390), .Z(n574) );
  AND U2293 ( .A(n186), .B(n2391), .Z(n2390) );
  XOR U2294 ( .A(n2392), .B(n2389), .Z(n2391) );
  XNOR U2295 ( .A(n571), .B(n2384), .Z(n2386) );
  XOR U2296 ( .A(n2393), .B(n2394), .Z(n571) );
  AND U2297 ( .A(n183), .B(n2395), .Z(n2394) );
  XOR U2298 ( .A(n2396), .B(n2393), .Z(n2395) );
  IV U2299 ( .A(n2388), .Z(n2384) );
  AND U2300 ( .A(n2020), .B(n2023), .Z(n2388) );
  XNOR U2301 ( .A(n2397), .B(n2398), .Z(n2023) );
  AND U2302 ( .A(n186), .B(n2399), .Z(n2398) );
  XNOR U2303 ( .A(n2400), .B(n2397), .Z(n2399) );
  XOR U2304 ( .A(n2401), .B(n2402), .Z(n186) );
  AND U2305 ( .A(n2403), .B(n2404), .Z(n2402) );
  XOR U2306 ( .A(n2031), .B(n2401), .Z(n2404) );
  IV U2307 ( .A(n2405), .Z(n2031) );
  AND U2308 ( .A(p_input[255]), .B(p_input[223]), .Z(n2405) );
  XOR U2309 ( .A(n2401), .B(n2028), .Z(n2403) );
  AND U2310 ( .A(p_input[159]), .B(p_input[191]), .Z(n2028) );
  XOR U2311 ( .A(n2406), .B(n2407), .Z(n2401) );
  AND U2312 ( .A(n2408), .B(n2409), .Z(n2407) );
  XOR U2313 ( .A(n2406), .B(n2043), .Z(n2409) );
  XNOR U2314 ( .A(p_input[222]), .B(n2410), .Z(n2043) );
  AND U2315 ( .A(n194), .B(n2411), .Z(n2410) );
  XOR U2316 ( .A(p_input[254]), .B(p_input[222]), .Z(n2411) );
  XNOR U2317 ( .A(n2040), .B(n2406), .Z(n2408) );
  XOR U2318 ( .A(n2412), .B(n2413), .Z(n2040) );
  AND U2319 ( .A(n192), .B(n2414), .Z(n2413) );
  XOR U2320 ( .A(p_input[190]), .B(p_input[158]), .Z(n2414) );
  XOR U2321 ( .A(n2415), .B(n2416), .Z(n2406) );
  AND U2322 ( .A(n2417), .B(n2418), .Z(n2416) );
  XOR U2323 ( .A(n2415), .B(n2055), .Z(n2418) );
  XNOR U2324 ( .A(p_input[221]), .B(n2419), .Z(n2055) );
  AND U2325 ( .A(n194), .B(n2420), .Z(n2419) );
  XOR U2326 ( .A(p_input[253]), .B(p_input[221]), .Z(n2420) );
  XNOR U2327 ( .A(n2052), .B(n2415), .Z(n2417) );
  XOR U2328 ( .A(n2421), .B(n2422), .Z(n2052) );
  AND U2329 ( .A(n192), .B(n2423), .Z(n2422) );
  XOR U2330 ( .A(p_input[189]), .B(p_input[157]), .Z(n2423) );
  XOR U2331 ( .A(n2424), .B(n2425), .Z(n2415) );
  AND U2332 ( .A(n2426), .B(n2427), .Z(n2425) );
  XOR U2333 ( .A(n2424), .B(n2067), .Z(n2427) );
  XNOR U2334 ( .A(p_input[220]), .B(n2428), .Z(n2067) );
  AND U2335 ( .A(n194), .B(n2429), .Z(n2428) );
  XOR U2336 ( .A(p_input[252]), .B(p_input[220]), .Z(n2429) );
  XNOR U2337 ( .A(n2064), .B(n2424), .Z(n2426) );
  XOR U2338 ( .A(n2430), .B(n2431), .Z(n2064) );
  AND U2339 ( .A(n192), .B(n2432), .Z(n2431) );
  XOR U2340 ( .A(p_input[188]), .B(p_input[156]), .Z(n2432) );
  XOR U2341 ( .A(n2433), .B(n2434), .Z(n2424) );
  AND U2342 ( .A(n2435), .B(n2436), .Z(n2434) );
  XOR U2343 ( .A(n2433), .B(n2079), .Z(n2436) );
  XNOR U2344 ( .A(p_input[219]), .B(n2437), .Z(n2079) );
  AND U2345 ( .A(n194), .B(n2438), .Z(n2437) );
  XOR U2346 ( .A(p_input[251]), .B(p_input[219]), .Z(n2438) );
  XNOR U2347 ( .A(n2076), .B(n2433), .Z(n2435) );
  XOR U2348 ( .A(n2439), .B(n2440), .Z(n2076) );
  AND U2349 ( .A(n192), .B(n2441), .Z(n2440) );
  XOR U2350 ( .A(p_input[187]), .B(p_input[155]), .Z(n2441) );
  XOR U2351 ( .A(n2442), .B(n2443), .Z(n2433) );
  AND U2352 ( .A(n2444), .B(n2445), .Z(n2443) );
  XOR U2353 ( .A(n2442), .B(n2091), .Z(n2445) );
  XNOR U2354 ( .A(p_input[218]), .B(n2446), .Z(n2091) );
  AND U2355 ( .A(n194), .B(n2447), .Z(n2446) );
  XOR U2356 ( .A(p_input[250]), .B(p_input[218]), .Z(n2447) );
  XNOR U2357 ( .A(n2088), .B(n2442), .Z(n2444) );
  XOR U2358 ( .A(n2448), .B(n2449), .Z(n2088) );
  AND U2359 ( .A(n192), .B(n2450), .Z(n2449) );
  XOR U2360 ( .A(p_input[186]), .B(p_input[154]), .Z(n2450) );
  XOR U2361 ( .A(n2451), .B(n2452), .Z(n2442) );
  AND U2362 ( .A(n2453), .B(n2454), .Z(n2452) );
  XOR U2363 ( .A(n2451), .B(n2103), .Z(n2454) );
  XNOR U2364 ( .A(p_input[217]), .B(n2455), .Z(n2103) );
  AND U2365 ( .A(n194), .B(n2456), .Z(n2455) );
  XOR U2366 ( .A(p_input[249]), .B(p_input[217]), .Z(n2456) );
  XNOR U2367 ( .A(n2100), .B(n2451), .Z(n2453) );
  XOR U2368 ( .A(n2457), .B(n2458), .Z(n2100) );
  AND U2369 ( .A(n192), .B(n2459), .Z(n2458) );
  XOR U2370 ( .A(p_input[185]), .B(p_input[153]), .Z(n2459) );
  XOR U2371 ( .A(n2460), .B(n2461), .Z(n2451) );
  AND U2372 ( .A(n2462), .B(n2463), .Z(n2461) );
  XOR U2373 ( .A(n2460), .B(n2115), .Z(n2463) );
  XNOR U2374 ( .A(p_input[216]), .B(n2464), .Z(n2115) );
  AND U2375 ( .A(n194), .B(n2465), .Z(n2464) );
  XOR U2376 ( .A(p_input[248]), .B(p_input[216]), .Z(n2465) );
  XNOR U2377 ( .A(n2112), .B(n2460), .Z(n2462) );
  XOR U2378 ( .A(n2466), .B(n2467), .Z(n2112) );
  AND U2379 ( .A(n192), .B(n2468), .Z(n2467) );
  XOR U2380 ( .A(p_input[184]), .B(p_input[152]), .Z(n2468) );
  XOR U2381 ( .A(n2469), .B(n2470), .Z(n2460) );
  AND U2382 ( .A(n2471), .B(n2472), .Z(n2470) );
  XOR U2383 ( .A(n2469), .B(n2127), .Z(n2472) );
  XNOR U2384 ( .A(p_input[215]), .B(n2473), .Z(n2127) );
  AND U2385 ( .A(n194), .B(n2474), .Z(n2473) );
  XOR U2386 ( .A(p_input[247]), .B(p_input[215]), .Z(n2474) );
  XNOR U2387 ( .A(n2124), .B(n2469), .Z(n2471) );
  XOR U2388 ( .A(n2475), .B(n2476), .Z(n2124) );
  AND U2389 ( .A(n192), .B(n2477), .Z(n2476) );
  XOR U2390 ( .A(p_input[183]), .B(p_input[151]), .Z(n2477) );
  XOR U2391 ( .A(n2478), .B(n2479), .Z(n2469) );
  AND U2392 ( .A(n2480), .B(n2481), .Z(n2479) );
  XOR U2393 ( .A(n2478), .B(n2139), .Z(n2481) );
  XNOR U2394 ( .A(p_input[214]), .B(n2482), .Z(n2139) );
  AND U2395 ( .A(n194), .B(n2483), .Z(n2482) );
  XOR U2396 ( .A(p_input[246]), .B(p_input[214]), .Z(n2483) );
  XNOR U2397 ( .A(n2136), .B(n2478), .Z(n2480) );
  XOR U2398 ( .A(n2484), .B(n2485), .Z(n2136) );
  AND U2399 ( .A(n192), .B(n2486), .Z(n2485) );
  XOR U2400 ( .A(p_input[182]), .B(p_input[150]), .Z(n2486) );
  XOR U2401 ( .A(n2487), .B(n2488), .Z(n2478) );
  AND U2402 ( .A(n2489), .B(n2490), .Z(n2488) );
  XOR U2403 ( .A(n2487), .B(n2151), .Z(n2490) );
  XNOR U2404 ( .A(p_input[213]), .B(n2491), .Z(n2151) );
  AND U2405 ( .A(n194), .B(n2492), .Z(n2491) );
  XOR U2406 ( .A(p_input[245]), .B(p_input[213]), .Z(n2492) );
  XNOR U2407 ( .A(n2148), .B(n2487), .Z(n2489) );
  XOR U2408 ( .A(n2493), .B(n2494), .Z(n2148) );
  AND U2409 ( .A(n192), .B(n2495), .Z(n2494) );
  XOR U2410 ( .A(p_input[181]), .B(p_input[149]), .Z(n2495) );
  XOR U2411 ( .A(n2496), .B(n2497), .Z(n2487) );
  AND U2412 ( .A(n2498), .B(n2499), .Z(n2497) );
  XOR U2413 ( .A(n2496), .B(n2163), .Z(n2499) );
  XNOR U2414 ( .A(p_input[212]), .B(n2500), .Z(n2163) );
  AND U2415 ( .A(n194), .B(n2501), .Z(n2500) );
  XOR U2416 ( .A(p_input[244]), .B(p_input[212]), .Z(n2501) );
  XNOR U2417 ( .A(n2160), .B(n2496), .Z(n2498) );
  XOR U2418 ( .A(n2502), .B(n2503), .Z(n2160) );
  AND U2419 ( .A(n192), .B(n2504), .Z(n2503) );
  XOR U2420 ( .A(p_input[180]), .B(p_input[148]), .Z(n2504) );
  XOR U2421 ( .A(n2505), .B(n2506), .Z(n2496) );
  AND U2422 ( .A(n2507), .B(n2508), .Z(n2506) );
  XOR U2423 ( .A(n2505), .B(n2175), .Z(n2508) );
  XNOR U2424 ( .A(p_input[211]), .B(n2509), .Z(n2175) );
  AND U2425 ( .A(n194), .B(n2510), .Z(n2509) );
  XOR U2426 ( .A(p_input[243]), .B(p_input[211]), .Z(n2510) );
  XNOR U2427 ( .A(n2172), .B(n2505), .Z(n2507) );
  XOR U2428 ( .A(n2511), .B(n2512), .Z(n2172) );
  AND U2429 ( .A(n192), .B(n2513), .Z(n2512) );
  XOR U2430 ( .A(p_input[179]), .B(p_input[147]), .Z(n2513) );
  XOR U2431 ( .A(n2514), .B(n2515), .Z(n2505) );
  AND U2432 ( .A(n2516), .B(n2517), .Z(n2515) );
  XOR U2433 ( .A(n2514), .B(n2187), .Z(n2517) );
  XNOR U2434 ( .A(p_input[210]), .B(n2518), .Z(n2187) );
  AND U2435 ( .A(n194), .B(n2519), .Z(n2518) );
  XOR U2436 ( .A(p_input[242]), .B(p_input[210]), .Z(n2519) );
  XNOR U2437 ( .A(n2184), .B(n2514), .Z(n2516) );
  XOR U2438 ( .A(n2520), .B(n2521), .Z(n2184) );
  AND U2439 ( .A(n192), .B(n2522), .Z(n2521) );
  XOR U2440 ( .A(p_input[178]), .B(p_input[146]), .Z(n2522) );
  XOR U2441 ( .A(n2523), .B(n2524), .Z(n2514) );
  AND U2442 ( .A(n2525), .B(n2526), .Z(n2524) );
  XOR U2443 ( .A(n2523), .B(n2199), .Z(n2526) );
  XNOR U2444 ( .A(p_input[209]), .B(n2527), .Z(n2199) );
  AND U2445 ( .A(n194), .B(n2528), .Z(n2527) );
  XOR U2446 ( .A(p_input[241]), .B(p_input[209]), .Z(n2528) );
  XNOR U2447 ( .A(n2196), .B(n2523), .Z(n2525) );
  XOR U2448 ( .A(n2529), .B(n2530), .Z(n2196) );
  AND U2449 ( .A(n192), .B(n2531), .Z(n2530) );
  XOR U2450 ( .A(p_input[177]), .B(p_input[145]), .Z(n2531) );
  XOR U2451 ( .A(n2532), .B(n2533), .Z(n2523) );
  AND U2452 ( .A(n2534), .B(n2535), .Z(n2533) );
  XOR U2453 ( .A(n2532), .B(n2211), .Z(n2535) );
  XNOR U2454 ( .A(p_input[208]), .B(n2536), .Z(n2211) );
  AND U2455 ( .A(n194), .B(n2537), .Z(n2536) );
  XOR U2456 ( .A(p_input[240]), .B(p_input[208]), .Z(n2537) );
  XNOR U2457 ( .A(n2208), .B(n2532), .Z(n2534) );
  XOR U2458 ( .A(n2538), .B(n2539), .Z(n2208) );
  AND U2459 ( .A(n192), .B(n2540), .Z(n2539) );
  XOR U2460 ( .A(p_input[176]), .B(p_input[144]), .Z(n2540) );
  XOR U2461 ( .A(n2541), .B(n2542), .Z(n2532) );
  AND U2462 ( .A(n2543), .B(n2544), .Z(n2542) );
  XOR U2463 ( .A(n2541), .B(n2223), .Z(n2544) );
  XNOR U2464 ( .A(p_input[207]), .B(n2545), .Z(n2223) );
  AND U2465 ( .A(n194), .B(n2546), .Z(n2545) );
  XOR U2466 ( .A(p_input[239]), .B(p_input[207]), .Z(n2546) );
  XNOR U2467 ( .A(n2220), .B(n2541), .Z(n2543) );
  XOR U2468 ( .A(n2547), .B(n2548), .Z(n2220) );
  AND U2469 ( .A(n192), .B(n2549), .Z(n2548) );
  XOR U2470 ( .A(p_input[175]), .B(p_input[143]), .Z(n2549) );
  XOR U2471 ( .A(n2550), .B(n2551), .Z(n2541) );
  AND U2472 ( .A(n2552), .B(n2553), .Z(n2551) );
  XOR U2473 ( .A(n2550), .B(n2235), .Z(n2553) );
  XNOR U2474 ( .A(p_input[206]), .B(n2554), .Z(n2235) );
  AND U2475 ( .A(n194), .B(n2555), .Z(n2554) );
  XOR U2476 ( .A(p_input[238]), .B(p_input[206]), .Z(n2555) );
  XNOR U2477 ( .A(n2232), .B(n2550), .Z(n2552) );
  XOR U2478 ( .A(n2556), .B(n2557), .Z(n2232) );
  AND U2479 ( .A(n192), .B(n2558), .Z(n2557) );
  XOR U2480 ( .A(p_input[174]), .B(p_input[142]), .Z(n2558) );
  XOR U2481 ( .A(n2559), .B(n2560), .Z(n2550) );
  AND U2482 ( .A(n2561), .B(n2562), .Z(n2560) );
  XOR U2483 ( .A(n2559), .B(n2247), .Z(n2562) );
  XNOR U2484 ( .A(p_input[205]), .B(n2563), .Z(n2247) );
  AND U2485 ( .A(n194), .B(n2564), .Z(n2563) );
  XOR U2486 ( .A(p_input[237]), .B(p_input[205]), .Z(n2564) );
  XNOR U2487 ( .A(n2244), .B(n2559), .Z(n2561) );
  XOR U2488 ( .A(n2565), .B(n2566), .Z(n2244) );
  AND U2489 ( .A(n192), .B(n2567), .Z(n2566) );
  XOR U2490 ( .A(p_input[173]), .B(p_input[141]), .Z(n2567) );
  XOR U2491 ( .A(n2568), .B(n2569), .Z(n2559) );
  AND U2492 ( .A(n2570), .B(n2571), .Z(n2569) );
  XOR U2493 ( .A(n2568), .B(n2259), .Z(n2571) );
  XNOR U2494 ( .A(p_input[204]), .B(n2572), .Z(n2259) );
  AND U2495 ( .A(n194), .B(n2573), .Z(n2572) );
  XOR U2496 ( .A(p_input[236]), .B(p_input[204]), .Z(n2573) );
  XNOR U2497 ( .A(n2256), .B(n2568), .Z(n2570) );
  XOR U2498 ( .A(n2574), .B(n2575), .Z(n2256) );
  AND U2499 ( .A(n192), .B(n2576), .Z(n2575) );
  XOR U2500 ( .A(p_input[172]), .B(p_input[140]), .Z(n2576) );
  XOR U2501 ( .A(n2577), .B(n2578), .Z(n2568) );
  AND U2502 ( .A(n2579), .B(n2580), .Z(n2578) );
  XOR U2503 ( .A(n2577), .B(n2271), .Z(n2580) );
  XNOR U2504 ( .A(p_input[203]), .B(n2581), .Z(n2271) );
  AND U2505 ( .A(n194), .B(n2582), .Z(n2581) );
  XOR U2506 ( .A(p_input[235]), .B(p_input[203]), .Z(n2582) );
  XNOR U2507 ( .A(n2268), .B(n2577), .Z(n2579) );
  XOR U2508 ( .A(n2583), .B(n2584), .Z(n2268) );
  AND U2509 ( .A(n192), .B(n2585), .Z(n2584) );
  XOR U2510 ( .A(p_input[171]), .B(p_input[139]), .Z(n2585) );
  XOR U2511 ( .A(n2586), .B(n2587), .Z(n2577) );
  AND U2512 ( .A(n2588), .B(n2589), .Z(n2587) );
  XOR U2513 ( .A(n2586), .B(n2283), .Z(n2589) );
  XNOR U2514 ( .A(p_input[202]), .B(n2590), .Z(n2283) );
  AND U2515 ( .A(n194), .B(n2591), .Z(n2590) );
  XOR U2516 ( .A(p_input[234]), .B(p_input[202]), .Z(n2591) );
  XNOR U2517 ( .A(n2280), .B(n2586), .Z(n2588) );
  XOR U2518 ( .A(n2592), .B(n2593), .Z(n2280) );
  AND U2519 ( .A(n192), .B(n2594), .Z(n2593) );
  XOR U2520 ( .A(p_input[170]), .B(p_input[138]), .Z(n2594) );
  XOR U2521 ( .A(n2595), .B(n2596), .Z(n2586) );
  AND U2522 ( .A(n2597), .B(n2598), .Z(n2596) );
  XOR U2523 ( .A(n2595), .B(n2295), .Z(n2598) );
  XNOR U2524 ( .A(p_input[201]), .B(n2599), .Z(n2295) );
  AND U2525 ( .A(n194), .B(n2600), .Z(n2599) );
  XOR U2526 ( .A(p_input[233]), .B(p_input[201]), .Z(n2600) );
  XNOR U2527 ( .A(n2292), .B(n2595), .Z(n2597) );
  XOR U2528 ( .A(n2601), .B(n2602), .Z(n2292) );
  AND U2529 ( .A(n192), .B(n2603), .Z(n2602) );
  XOR U2530 ( .A(p_input[169]), .B(p_input[137]), .Z(n2603) );
  XOR U2531 ( .A(n2604), .B(n2605), .Z(n2595) );
  AND U2532 ( .A(n2606), .B(n2607), .Z(n2605) );
  XOR U2533 ( .A(n2604), .B(n2307), .Z(n2607) );
  XNOR U2534 ( .A(p_input[200]), .B(n2608), .Z(n2307) );
  AND U2535 ( .A(n194), .B(n2609), .Z(n2608) );
  XOR U2536 ( .A(p_input[232]), .B(p_input[200]), .Z(n2609) );
  XNOR U2537 ( .A(n2304), .B(n2604), .Z(n2606) );
  XOR U2538 ( .A(n2610), .B(n2611), .Z(n2304) );
  AND U2539 ( .A(n192), .B(n2612), .Z(n2611) );
  XOR U2540 ( .A(p_input[168]), .B(p_input[136]), .Z(n2612) );
  XOR U2541 ( .A(n2613), .B(n2614), .Z(n2604) );
  AND U2542 ( .A(n2615), .B(n2616), .Z(n2614) );
  XOR U2543 ( .A(n2613), .B(n2319), .Z(n2616) );
  XNOR U2544 ( .A(p_input[199]), .B(n2617), .Z(n2319) );
  AND U2545 ( .A(n194), .B(n2618), .Z(n2617) );
  XOR U2546 ( .A(p_input[231]), .B(p_input[199]), .Z(n2618) );
  XNOR U2547 ( .A(n2316), .B(n2613), .Z(n2615) );
  XOR U2548 ( .A(n2619), .B(n2620), .Z(n2316) );
  AND U2549 ( .A(n192), .B(n2621), .Z(n2620) );
  XOR U2550 ( .A(p_input[167]), .B(p_input[135]), .Z(n2621) );
  XOR U2551 ( .A(n2622), .B(n2623), .Z(n2613) );
  AND U2552 ( .A(n2624), .B(n2625), .Z(n2623) );
  XOR U2553 ( .A(n2622), .B(n2331), .Z(n2625) );
  XNOR U2554 ( .A(p_input[198]), .B(n2626), .Z(n2331) );
  AND U2555 ( .A(n194), .B(n2627), .Z(n2626) );
  XOR U2556 ( .A(p_input[230]), .B(p_input[198]), .Z(n2627) );
  XNOR U2557 ( .A(n2328), .B(n2622), .Z(n2624) );
  XOR U2558 ( .A(n2628), .B(n2629), .Z(n2328) );
  AND U2559 ( .A(n192), .B(n2630), .Z(n2629) );
  XOR U2560 ( .A(p_input[166]), .B(p_input[134]), .Z(n2630) );
  XOR U2561 ( .A(n2631), .B(n2632), .Z(n2622) );
  AND U2562 ( .A(n2633), .B(n2634), .Z(n2632) );
  XOR U2563 ( .A(n2343), .B(n2631), .Z(n2634) );
  XNOR U2564 ( .A(p_input[197]), .B(n2635), .Z(n2343) );
  AND U2565 ( .A(n194), .B(n2636), .Z(n2635) );
  XOR U2566 ( .A(p_input[229]), .B(p_input[197]), .Z(n2636) );
  XNOR U2567 ( .A(n2631), .B(n2340), .Z(n2633) );
  XOR U2568 ( .A(n2637), .B(n2638), .Z(n2340) );
  AND U2569 ( .A(n192), .B(n2639), .Z(n2638) );
  XOR U2570 ( .A(p_input[165]), .B(p_input[133]), .Z(n2639) );
  XOR U2571 ( .A(n2640), .B(n2641), .Z(n2631) );
  AND U2572 ( .A(n2642), .B(n2643), .Z(n2641) );
  XOR U2573 ( .A(n2640), .B(n2355), .Z(n2643) );
  XNOR U2574 ( .A(p_input[196]), .B(n2644), .Z(n2355) );
  AND U2575 ( .A(n194), .B(n2645), .Z(n2644) );
  XOR U2576 ( .A(p_input[228]), .B(p_input[196]), .Z(n2645) );
  XNOR U2577 ( .A(n2352), .B(n2640), .Z(n2642) );
  XOR U2578 ( .A(n2646), .B(n2647), .Z(n2352) );
  AND U2579 ( .A(n192), .B(n2648), .Z(n2647) );
  XOR U2580 ( .A(p_input[164]), .B(p_input[132]), .Z(n2648) );
  XOR U2581 ( .A(n2649), .B(n2650), .Z(n2640) );
  AND U2582 ( .A(n2651), .B(n2652), .Z(n2650) );
  XOR U2583 ( .A(n2649), .B(n2367), .Z(n2652) );
  XNOR U2584 ( .A(p_input[195]), .B(n2653), .Z(n2367) );
  AND U2585 ( .A(n194), .B(n2654), .Z(n2653) );
  XOR U2586 ( .A(p_input[227]), .B(p_input[195]), .Z(n2654) );
  XNOR U2587 ( .A(n2364), .B(n2649), .Z(n2651) );
  XOR U2588 ( .A(n2655), .B(n2656), .Z(n2364) );
  AND U2589 ( .A(n192), .B(n2657), .Z(n2656) );
  XOR U2590 ( .A(p_input[163]), .B(p_input[131]), .Z(n2657) );
  XOR U2591 ( .A(n2658), .B(n2659), .Z(n2649) );
  AND U2592 ( .A(n2660), .B(n2661), .Z(n2659) );
  XOR U2593 ( .A(n2658), .B(n2379), .Z(n2661) );
  XNOR U2594 ( .A(p_input[194]), .B(n2662), .Z(n2379) );
  AND U2595 ( .A(n194), .B(n2663), .Z(n2662) );
  XOR U2596 ( .A(p_input[226]), .B(p_input[194]), .Z(n2663) );
  XNOR U2597 ( .A(n2376), .B(n2658), .Z(n2660) );
  XOR U2598 ( .A(n2664), .B(n2665), .Z(n2376) );
  AND U2599 ( .A(n192), .B(n2666), .Z(n2665) );
  XOR U2600 ( .A(p_input[162]), .B(p_input[130]), .Z(n2666) );
  XOR U2601 ( .A(n2667), .B(n2668), .Z(n2658) );
  AND U2602 ( .A(n2669), .B(n2670), .Z(n2668) );
  XNOR U2603 ( .A(n2671), .B(n2392), .Z(n2670) );
  XNOR U2604 ( .A(p_input[193]), .B(n2672), .Z(n2392) );
  AND U2605 ( .A(n194), .B(n2673), .Z(n2672) );
  XNOR U2606 ( .A(p_input[225]), .B(n2674), .Z(n2673) );
  IV U2607 ( .A(p_input[193]), .Z(n2674) );
  XNOR U2608 ( .A(n2389), .B(n2667), .Z(n2669) );
  XNOR U2609 ( .A(p_input[129]), .B(n2675), .Z(n2389) );
  AND U2610 ( .A(n192), .B(n2676), .Z(n2675) );
  XOR U2611 ( .A(p_input[161]), .B(p_input[129]), .Z(n2676) );
  IV U2612 ( .A(n2671), .Z(n2667) );
  AND U2613 ( .A(n2397), .B(n2400), .Z(n2671) );
  XOR U2614 ( .A(p_input[192]), .B(n2677), .Z(n2400) );
  AND U2615 ( .A(n194), .B(n2678), .Z(n2677) );
  XOR U2616 ( .A(p_input[224]), .B(p_input[192]), .Z(n2678) );
  XOR U2617 ( .A(n2679), .B(n2680), .Z(n194) );
  AND U2618 ( .A(n2681), .B(n2682), .Z(n2680) );
  XNOR U2619 ( .A(p_input[255]), .B(n2679), .Z(n2682) );
  XOR U2620 ( .A(n2679), .B(p_input[223]), .Z(n2681) );
  XOR U2621 ( .A(n2683), .B(n2684), .Z(n2679) );
  AND U2622 ( .A(n2685), .B(n2686), .Z(n2684) );
  XNOR U2623 ( .A(p_input[254]), .B(n2683), .Z(n2686) );
  XOR U2624 ( .A(n2683), .B(p_input[222]), .Z(n2685) );
  XOR U2625 ( .A(n2687), .B(n2688), .Z(n2683) );
  AND U2626 ( .A(n2689), .B(n2690), .Z(n2688) );
  XNOR U2627 ( .A(p_input[253]), .B(n2687), .Z(n2690) );
  XOR U2628 ( .A(n2687), .B(p_input[221]), .Z(n2689) );
  XOR U2629 ( .A(n2691), .B(n2692), .Z(n2687) );
  AND U2630 ( .A(n2693), .B(n2694), .Z(n2692) );
  XNOR U2631 ( .A(p_input[252]), .B(n2691), .Z(n2694) );
  XOR U2632 ( .A(n2691), .B(p_input[220]), .Z(n2693) );
  XOR U2633 ( .A(n2695), .B(n2696), .Z(n2691) );
  AND U2634 ( .A(n2697), .B(n2698), .Z(n2696) );
  XNOR U2635 ( .A(p_input[251]), .B(n2695), .Z(n2698) );
  XOR U2636 ( .A(n2695), .B(p_input[219]), .Z(n2697) );
  XOR U2637 ( .A(n2699), .B(n2700), .Z(n2695) );
  AND U2638 ( .A(n2701), .B(n2702), .Z(n2700) );
  XNOR U2639 ( .A(p_input[250]), .B(n2699), .Z(n2702) );
  XOR U2640 ( .A(n2699), .B(p_input[218]), .Z(n2701) );
  XOR U2641 ( .A(n2703), .B(n2704), .Z(n2699) );
  AND U2642 ( .A(n2705), .B(n2706), .Z(n2704) );
  XNOR U2643 ( .A(p_input[249]), .B(n2703), .Z(n2706) );
  XOR U2644 ( .A(n2703), .B(p_input[217]), .Z(n2705) );
  XOR U2645 ( .A(n2707), .B(n2708), .Z(n2703) );
  AND U2646 ( .A(n2709), .B(n2710), .Z(n2708) );
  XNOR U2647 ( .A(p_input[248]), .B(n2707), .Z(n2710) );
  XOR U2648 ( .A(n2707), .B(p_input[216]), .Z(n2709) );
  XOR U2649 ( .A(n2711), .B(n2712), .Z(n2707) );
  AND U2650 ( .A(n2713), .B(n2714), .Z(n2712) );
  XNOR U2651 ( .A(p_input[247]), .B(n2711), .Z(n2714) );
  XOR U2652 ( .A(n2711), .B(p_input[215]), .Z(n2713) );
  XOR U2653 ( .A(n2715), .B(n2716), .Z(n2711) );
  AND U2654 ( .A(n2717), .B(n2718), .Z(n2716) );
  XNOR U2655 ( .A(p_input[246]), .B(n2715), .Z(n2718) );
  XOR U2656 ( .A(n2715), .B(p_input[214]), .Z(n2717) );
  XOR U2657 ( .A(n2719), .B(n2720), .Z(n2715) );
  AND U2658 ( .A(n2721), .B(n2722), .Z(n2720) );
  XNOR U2659 ( .A(p_input[245]), .B(n2719), .Z(n2722) );
  XOR U2660 ( .A(n2719), .B(p_input[213]), .Z(n2721) );
  XOR U2661 ( .A(n2723), .B(n2724), .Z(n2719) );
  AND U2662 ( .A(n2725), .B(n2726), .Z(n2724) );
  XNOR U2663 ( .A(p_input[244]), .B(n2723), .Z(n2726) );
  XOR U2664 ( .A(n2723), .B(p_input[212]), .Z(n2725) );
  XOR U2665 ( .A(n2727), .B(n2728), .Z(n2723) );
  AND U2666 ( .A(n2729), .B(n2730), .Z(n2728) );
  XNOR U2667 ( .A(p_input[243]), .B(n2727), .Z(n2730) );
  XOR U2668 ( .A(n2727), .B(p_input[211]), .Z(n2729) );
  XOR U2669 ( .A(n2731), .B(n2732), .Z(n2727) );
  AND U2670 ( .A(n2733), .B(n2734), .Z(n2732) );
  XNOR U2671 ( .A(p_input[242]), .B(n2731), .Z(n2734) );
  XOR U2672 ( .A(n2731), .B(p_input[210]), .Z(n2733) );
  XOR U2673 ( .A(n2735), .B(n2736), .Z(n2731) );
  AND U2674 ( .A(n2737), .B(n2738), .Z(n2736) );
  XNOR U2675 ( .A(p_input[241]), .B(n2735), .Z(n2738) );
  XOR U2676 ( .A(n2735), .B(p_input[209]), .Z(n2737) );
  XOR U2677 ( .A(n2739), .B(n2740), .Z(n2735) );
  AND U2678 ( .A(n2741), .B(n2742), .Z(n2740) );
  XNOR U2679 ( .A(p_input[240]), .B(n2739), .Z(n2742) );
  XOR U2680 ( .A(n2739), .B(p_input[208]), .Z(n2741) );
  XOR U2681 ( .A(n2743), .B(n2744), .Z(n2739) );
  AND U2682 ( .A(n2745), .B(n2746), .Z(n2744) );
  XNOR U2683 ( .A(p_input[239]), .B(n2743), .Z(n2746) );
  XOR U2684 ( .A(n2743), .B(p_input[207]), .Z(n2745) );
  XOR U2685 ( .A(n2747), .B(n2748), .Z(n2743) );
  AND U2686 ( .A(n2749), .B(n2750), .Z(n2748) );
  XNOR U2687 ( .A(p_input[238]), .B(n2747), .Z(n2750) );
  XOR U2688 ( .A(n2747), .B(p_input[206]), .Z(n2749) );
  XOR U2689 ( .A(n2751), .B(n2752), .Z(n2747) );
  AND U2690 ( .A(n2753), .B(n2754), .Z(n2752) );
  XNOR U2691 ( .A(p_input[237]), .B(n2751), .Z(n2754) );
  XOR U2692 ( .A(n2751), .B(p_input[205]), .Z(n2753) );
  XOR U2693 ( .A(n2755), .B(n2756), .Z(n2751) );
  AND U2694 ( .A(n2757), .B(n2758), .Z(n2756) );
  XNOR U2695 ( .A(p_input[236]), .B(n2755), .Z(n2758) );
  XOR U2696 ( .A(n2755), .B(p_input[204]), .Z(n2757) );
  XOR U2697 ( .A(n2759), .B(n2760), .Z(n2755) );
  AND U2698 ( .A(n2761), .B(n2762), .Z(n2760) );
  XNOR U2699 ( .A(p_input[235]), .B(n2759), .Z(n2762) );
  XOR U2700 ( .A(n2759), .B(p_input[203]), .Z(n2761) );
  XOR U2701 ( .A(n2763), .B(n2764), .Z(n2759) );
  AND U2702 ( .A(n2765), .B(n2766), .Z(n2764) );
  XNOR U2703 ( .A(p_input[234]), .B(n2763), .Z(n2766) );
  XOR U2704 ( .A(n2763), .B(p_input[202]), .Z(n2765) );
  XOR U2705 ( .A(n2767), .B(n2768), .Z(n2763) );
  AND U2706 ( .A(n2769), .B(n2770), .Z(n2768) );
  XNOR U2707 ( .A(p_input[233]), .B(n2767), .Z(n2770) );
  XOR U2708 ( .A(n2767), .B(p_input[201]), .Z(n2769) );
  XOR U2709 ( .A(n2771), .B(n2772), .Z(n2767) );
  AND U2710 ( .A(n2773), .B(n2774), .Z(n2772) );
  XNOR U2711 ( .A(p_input[232]), .B(n2771), .Z(n2774) );
  XOR U2712 ( .A(n2771), .B(p_input[200]), .Z(n2773) );
  XOR U2713 ( .A(n2775), .B(n2776), .Z(n2771) );
  AND U2714 ( .A(n2777), .B(n2778), .Z(n2776) );
  XNOR U2715 ( .A(p_input[231]), .B(n2775), .Z(n2778) );
  XOR U2716 ( .A(n2775), .B(p_input[199]), .Z(n2777) );
  XOR U2717 ( .A(n2779), .B(n2780), .Z(n2775) );
  AND U2718 ( .A(n2781), .B(n2782), .Z(n2780) );
  XNOR U2719 ( .A(p_input[230]), .B(n2779), .Z(n2782) );
  XOR U2720 ( .A(n2779), .B(p_input[198]), .Z(n2781) );
  XOR U2721 ( .A(n2783), .B(n2784), .Z(n2779) );
  AND U2722 ( .A(n2785), .B(n2786), .Z(n2784) );
  XNOR U2723 ( .A(p_input[229]), .B(n2783), .Z(n2786) );
  XOR U2724 ( .A(n2783), .B(p_input[197]), .Z(n2785) );
  XOR U2725 ( .A(n2787), .B(n2788), .Z(n2783) );
  AND U2726 ( .A(n2789), .B(n2790), .Z(n2788) );
  XNOR U2727 ( .A(p_input[228]), .B(n2787), .Z(n2790) );
  XOR U2728 ( .A(n2787), .B(p_input[196]), .Z(n2789) );
  XOR U2729 ( .A(n2791), .B(n2792), .Z(n2787) );
  AND U2730 ( .A(n2793), .B(n2794), .Z(n2792) );
  XNOR U2731 ( .A(p_input[227]), .B(n2791), .Z(n2794) );
  XOR U2732 ( .A(n2791), .B(p_input[195]), .Z(n2793) );
  XOR U2733 ( .A(n2795), .B(n2796), .Z(n2791) );
  AND U2734 ( .A(n2797), .B(n2798), .Z(n2796) );
  XNOR U2735 ( .A(p_input[226]), .B(n2795), .Z(n2798) );
  XOR U2736 ( .A(n2795), .B(p_input[194]), .Z(n2797) );
  XNOR U2737 ( .A(n2799), .B(n2800), .Z(n2795) );
  AND U2738 ( .A(n2801), .B(n2802), .Z(n2800) );
  XOR U2739 ( .A(p_input[225]), .B(n2799), .Z(n2802) );
  XNOR U2740 ( .A(p_input[193]), .B(n2799), .Z(n2801) );
  AND U2741 ( .A(p_input[224]), .B(n2803), .Z(n2799) );
  IV U2742 ( .A(p_input[192]), .Z(n2803) );
  XNOR U2743 ( .A(p_input[128]), .B(n2804), .Z(n2397) );
  AND U2744 ( .A(n192), .B(n2805), .Z(n2804) );
  XOR U2745 ( .A(p_input[160]), .B(p_input[128]), .Z(n2805) );
  XOR U2746 ( .A(n2806), .B(n2807), .Z(n192) );
  AND U2747 ( .A(n2808), .B(n2809), .Z(n2807) );
  XNOR U2748 ( .A(p_input[191]), .B(n2806), .Z(n2809) );
  XOR U2749 ( .A(n2806), .B(p_input[159]), .Z(n2808) );
  XOR U2750 ( .A(n2810), .B(n2811), .Z(n2806) );
  AND U2751 ( .A(n2812), .B(n2813), .Z(n2811) );
  XNOR U2752 ( .A(p_input[190]), .B(n2810), .Z(n2813) );
  XNOR U2753 ( .A(n2810), .B(n2412), .Z(n2812) );
  IV U2754 ( .A(p_input[158]), .Z(n2412) );
  XOR U2755 ( .A(n2814), .B(n2815), .Z(n2810) );
  AND U2756 ( .A(n2816), .B(n2817), .Z(n2815) );
  XNOR U2757 ( .A(p_input[189]), .B(n2814), .Z(n2817) );
  XNOR U2758 ( .A(n2814), .B(n2421), .Z(n2816) );
  IV U2759 ( .A(p_input[157]), .Z(n2421) );
  XOR U2760 ( .A(n2818), .B(n2819), .Z(n2814) );
  AND U2761 ( .A(n2820), .B(n2821), .Z(n2819) );
  XNOR U2762 ( .A(p_input[188]), .B(n2818), .Z(n2821) );
  XNOR U2763 ( .A(n2818), .B(n2430), .Z(n2820) );
  IV U2764 ( .A(p_input[156]), .Z(n2430) );
  XOR U2765 ( .A(n2822), .B(n2823), .Z(n2818) );
  AND U2766 ( .A(n2824), .B(n2825), .Z(n2823) );
  XNOR U2767 ( .A(p_input[187]), .B(n2822), .Z(n2825) );
  XNOR U2768 ( .A(n2822), .B(n2439), .Z(n2824) );
  IV U2769 ( .A(p_input[155]), .Z(n2439) );
  XOR U2770 ( .A(n2826), .B(n2827), .Z(n2822) );
  AND U2771 ( .A(n2828), .B(n2829), .Z(n2827) );
  XNOR U2772 ( .A(p_input[186]), .B(n2826), .Z(n2829) );
  XNOR U2773 ( .A(n2826), .B(n2448), .Z(n2828) );
  IV U2774 ( .A(p_input[154]), .Z(n2448) );
  XOR U2775 ( .A(n2830), .B(n2831), .Z(n2826) );
  AND U2776 ( .A(n2832), .B(n2833), .Z(n2831) );
  XNOR U2777 ( .A(p_input[185]), .B(n2830), .Z(n2833) );
  XNOR U2778 ( .A(n2830), .B(n2457), .Z(n2832) );
  IV U2779 ( .A(p_input[153]), .Z(n2457) );
  XOR U2780 ( .A(n2834), .B(n2835), .Z(n2830) );
  AND U2781 ( .A(n2836), .B(n2837), .Z(n2835) );
  XNOR U2782 ( .A(p_input[184]), .B(n2834), .Z(n2837) );
  XNOR U2783 ( .A(n2834), .B(n2466), .Z(n2836) );
  IV U2784 ( .A(p_input[152]), .Z(n2466) );
  XOR U2785 ( .A(n2838), .B(n2839), .Z(n2834) );
  AND U2786 ( .A(n2840), .B(n2841), .Z(n2839) );
  XNOR U2787 ( .A(p_input[183]), .B(n2838), .Z(n2841) );
  XNOR U2788 ( .A(n2838), .B(n2475), .Z(n2840) );
  IV U2789 ( .A(p_input[151]), .Z(n2475) );
  XOR U2790 ( .A(n2842), .B(n2843), .Z(n2838) );
  AND U2791 ( .A(n2844), .B(n2845), .Z(n2843) );
  XNOR U2792 ( .A(p_input[182]), .B(n2842), .Z(n2845) );
  XNOR U2793 ( .A(n2842), .B(n2484), .Z(n2844) );
  IV U2794 ( .A(p_input[150]), .Z(n2484) );
  XOR U2795 ( .A(n2846), .B(n2847), .Z(n2842) );
  AND U2796 ( .A(n2848), .B(n2849), .Z(n2847) );
  XNOR U2797 ( .A(p_input[181]), .B(n2846), .Z(n2849) );
  XNOR U2798 ( .A(n2846), .B(n2493), .Z(n2848) );
  IV U2799 ( .A(p_input[149]), .Z(n2493) );
  XOR U2800 ( .A(n2850), .B(n2851), .Z(n2846) );
  AND U2801 ( .A(n2852), .B(n2853), .Z(n2851) );
  XNOR U2802 ( .A(p_input[180]), .B(n2850), .Z(n2853) );
  XNOR U2803 ( .A(n2850), .B(n2502), .Z(n2852) );
  IV U2804 ( .A(p_input[148]), .Z(n2502) );
  XOR U2805 ( .A(n2854), .B(n2855), .Z(n2850) );
  AND U2806 ( .A(n2856), .B(n2857), .Z(n2855) );
  XNOR U2807 ( .A(p_input[179]), .B(n2854), .Z(n2857) );
  XNOR U2808 ( .A(n2854), .B(n2511), .Z(n2856) );
  IV U2809 ( .A(p_input[147]), .Z(n2511) );
  XOR U2810 ( .A(n2858), .B(n2859), .Z(n2854) );
  AND U2811 ( .A(n2860), .B(n2861), .Z(n2859) );
  XNOR U2812 ( .A(p_input[178]), .B(n2858), .Z(n2861) );
  XNOR U2813 ( .A(n2858), .B(n2520), .Z(n2860) );
  IV U2814 ( .A(p_input[146]), .Z(n2520) );
  XOR U2815 ( .A(n2862), .B(n2863), .Z(n2858) );
  AND U2816 ( .A(n2864), .B(n2865), .Z(n2863) );
  XNOR U2817 ( .A(p_input[177]), .B(n2862), .Z(n2865) );
  XNOR U2818 ( .A(n2862), .B(n2529), .Z(n2864) );
  IV U2819 ( .A(p_input[145]), .Z(n2529) );
  XOR U2820 ( .A(n2866), .B(n2867), .Z(n2862) );
  AND U2821 ( .A(n2868), .B(n2869), .Z(n2867) );
  XNOR U2822 ( .A(p_input[176]), .B(n2866), .Z(n2869) );
  XNOR U2823 ( .A(n2866), .B(n2538), .Z(n2868) );
  IV U2824 ( .A(p_input[144]), .Z(n2538) );
  XOR U2825 ( .A(n2870), .B(n2871), .Z(n2866) );
  AND U2826 ( .A(n2872), .B(n2873), .Z(n2871) );
  XNOR U2827 ( .A(p_input[175]), .B(n2870), .Z(n2873) );
  XNOR U2828 ( .A(n2870), .B(n2547), .Z(n2872) );
  IV U2829 ( .A(p_input[143]), .Z(n2547) );
  XOR U2830 ( .A(n2874), .B(n2875), .Z(n2870) );
  AND U2831 ( .A(n2876), .B(n2877), .Z(n2875) );
  XNOR U2832 ( .A(p_input[174]), .B(n2874), .Z(n2877) );
  XNOR U2833 ( .A(n2874), .B(n2556), .Z(n2876) );
  IV U2834 ( .A(p_input[142]), .Z(n2556) );
  XOR U2835 ( .A(n2878), .B(n2879), .Z(n2874) );
  AND U2836 ( .A(n2880), .B(n2881), .Z(n2879) );
  XNOR U2837 ( .A(p_input[173]), .B(n2878), .Z(n2881) );
  XNOR U2838 ( .A(n2878), .B(n2565), .Z(n2880) );
  IV U2839 ( .A(p_input[141]), .Z(n2565) );
  XOR U2840 ( .A(n2882), .B(n2883), .Z(n2878) );
  AND U2841 ( .A(n2884), .B(n2885), .Z(n2883) );
  XNOR U2842 ( .A(p_input[172]), .B(n2882), .Z(n2885) );
  XNOR U2843 ( .A(n2882), .B(n2574), .Z(n2884) );
  IV U2844 ( .A(p_input[140]), .Z(n2574) );
  XOR U2845 ( .A(n2886), .B(n2887), .Z(n2882) );
  AND U2846 ( .A(n2888), .B(n2889), .Z(n2887) );
  XNOR U2847 ( .A(p_input[171]), .B(n2886), .Z(n2889) );
  XNOR U2848 ( .A(n2886), .B(n2583), .Z(n2888) );
  IV U2849 ( .A(p_input[139]), .Z(n2583) );
  XOR U2850 ( .A(n2890), .B(n2891), .Z(n2886) );
  AND U2851 ( .A(n2892), .B(n2893), .Z(n2891) );
  XNOR U2852 ( .A(p_input[170]), .B(n2890), .Z(n2893) );
  XNOR U2853 ( .A(n2890), .B(n2592), .Z(n2892) );
  IV U2854 ( .A(p_input[138]), .Z(n2592) );
  XOR U2855 ( .A(n2894), .B(n2895), .Z(n2890) );
  AND U2856 ( .A(n2896), .B(n2897), .Z(n2895) );
  XNOR U2857 ( .A(p_input[169]), .B(n2894), .Z(n2897) );
  XNOR U2858 ( .A(n2894), .B(n2601), .Z(n2896) );
  IV U2859 ( .A(p_input[137]), .Z(n2601) );
  XOR U2860 ( .A(n2898), .B(n2899), .Z(n2894) );
  AND U2861 ( .A(n2900), .B(n2901), .Z(n2899) );
  XNOR U2862 ( .A(p_input[168]), .B(n2898), .Z(n2901) );
  XNOR U2863 ( .A(n2898), .B(n2610), .Z(n2900) );
  IV U2864 ( .A(p_input[136]), .Z(n2610) );
  XOR U2865 ( .A(n2902), .B(n2903), .Z(n2898) );
  AND U2866 ( .A(n2904), .B(n2905), .Z(n2903) );
  XNOR U2867 ( .A(p_input[167]), .B(n2902), .Z(n2905) );
  XNOR U2868 ( .A(n2902), .B(n2619), .Z(n2904) );
  IV U2869 ( .A(p_input[135]), .Z(n2619) );
  XOR U2870 ( .A(n2906), .B(n2907), .Z(n2902) );
  AND U2871 ( .A(n2908), .B(n2909), .Z(n2907) );
  XNOR U2872 ( .A(p_input[166]), .B(n2906), .Z(n2909) );
  XNOR U2873 ( .A(n2906), .B(n2628), .Z(n2908) );
  IV U2874 ( .A(p_input[134]), .Z(n2628) );
  XOR U2875 ( .A(n2910), .B(n2911), .Z(n2906) );
  AND U2876 ( .A(n2912), .B(n2913), .Z(n2911) );
  XNOR U2877 ( .A(p_input[165]), .B(n2910), .Z(n2913) );
  XNOR U2878 ( .A(n2910), .B(n2637), .Z(n2912) );
  IV U2879 ( .A(p_input[133]), .Z(n2637) );
  XOR U2880 ( .A(n2914), .B(n2915), .Z(n2910) );
  AND U2881 ( .A(n2916), .B(n2917), .Z(n2915) );
  XNOR U2882 ( .A(p_input[164]), .B(n2914), .Z(n2917) );
  XNOR U2883 ( .A(n2914), .B(n2646), .Z(n2916) );
  IV U2884 ( .A(p_input[132]), .Z(n2646) );
  XOR U2885 ( .A(n2918), .B(n2919), .Z(n2914) );
  AND U2886 ( .A(n2920), .B(n2921), .Z(n2919) );
  XNOR U2887 ( .A(p_input[163]), .B(n2918), .Z(n2921) );
  XNOR U2888 ( .A(n2918), .B(n2655), .Z(n2920) );
  IV U2889 ( .A(p_input[131]), .Z(n2655) );
  XOR U2890 ( .A(n2922), .B(n2923), .Z(n2918) );
  AND U2891 ( .A(n2924), .B(n2925), .Z(n2923) );
  XNOR U2892 ( .A(p_input[162]), .B(n2922), .Z(n2925) );
  XNOR U2893 ( .A(n2922), .B(n2664), .Z(n2924) );
  IV U2894 ( .A(p_input[130]), .Z(n2664) );
  XNOR U2895 ( .A(n2926), .B(n2927), .Z(n2922) );
  AND U2896 ( .A(n2928), .B(n2929), .Z(n2927) );
  XOR U2897 ( .A(p_input[161]), .B(n2926), .Z(n2929) );
  XNOR U2898 ( .A(p_input[129]), .B(n2926), .Z(n2928) );
  AND U2899 ( .A(p_input[160]), .B(n2930), .Z(n2926) );
  IV U2900 ( .A(p_input[128]), .Z(n2930) );
  XOR U2901 ( .A(n2931), .B(n2932), .Z(n2020) );
  AND U2902 ( .A(n183), .B(n2933), .Z(n2932) );
  XNOR U2903 ( .A(n2934), .B(n2931), .Z(n2933) );
  XOR U2904 ( .A(n2935), .B(n2936), .Z(n183) );
  AND U2905 ( .A(n2937), .B(n2938), .Z(n2936) );
  XNOR U2906 ( .A(n2035), .B(n2935), .Z(n2938) );
  AND U2907 ( .A(p_input[95]), .B(p_input[127]), .Z(n2035) );
  XNOR U2908 ( .A(n2935), .B(n2032), .Z(n2937) );
  IV U2909 ( .A(n2939), .Z(n2032) );
  AND U2910 ( .A(p_input[31]), .B(p_input[63]), .Z(n2939) );
  XOR U2911 ( .A(n2940), .B(n2941), .Z(n2935) );
  AND U2912 ( .A(n2942), .B(n2943), .Z(n2941) );
  XOR U2913 ( .A(n2940), .B(n2047), .Z(n2943) );
  XNOR U2914 ( .A(p_input[94]), .B(n2944), .Z(n2047) );
  AND U2915 ( .A(n202), .B(n2945), .Z(n2944) );
  XOR U2916 ( .A(p_input[94]), .B(p_input[126]), .Z(n2945) );
  XNOR U2917 ( .A(n2044), .B(n2940), .Z(n2942) );
  XOR U2918 ( .A(n2946), .B(n2947), .Z(n2044) );
  AND U2919 ( .A(n199), .B(n2948), .Z(n2947) );
  XOR U2920 ( .A(p_input[62]), .B(p_input[30]), .Z(n2948) );
  XOR U2921 ( .A(n2949), .B(n2950), .Z(n2940) );
  AND U2922 ( .A(n2951), .B(n2952), .Z(n2950) );
  XOR U2923 ( .A(n2949), .B(n2059), .Z(n2952) );
  XNOR U2924 ( .A(p_input[93]), .B(n2953), .Z(n2059) );
  AND U2925 ( .A(n202), .B(n2954), .Z(n2953) );
  XOR U2926 ( .A(p_input[93]), .B(p_input[125]), .Z(n2954) );
  XNOR U2927 ( .A(n2056), .B(n2949), .Z(n2951) );
  XOR U2928 ( .A(n2955), .B(n2956), .Z(n2056) );
  AND U2929 ( .A(n199), .B(n2957), .Z(n2956) );
  XOR U2930 ( .A(p_input[61]), .B(p_input[29]), .Z(n2957) );
  XOR U2931 ( .A(n2958), .B(n2959), .Z(n2949) );
  AND U2932 ( .A(n2960), .B(n2961), .Z(n2959) );
  XOR U2933 ( .A(n2958), .B(n2071), .Z(n2961) );
  XNOR U2934 ( .A(p_input[92]), .B(n2962), .Z(n2071) );
  AND U2935 ( .A(n202), .B(n2963), .Z(n2962) );
  XOR U2936 ( .A(p_input[92]), .B(p_input[124]), .Z(n2963) );
  XNOR U2937 ( .A(n2068), .B(n2958), .Z(n2960) );
  XOR U2938 ( .A(n2964), .B(n2965), .Z(n2068) );
  AND U2939 ( .A(n199), .B(n2966), .Z(n2965) );
  XOR U2940 ( .A(p_input[60]), .B(p_input[28]), .Z(n2966) );
  XOR U2941 ( .A(n2967), .B(n2968), .Z(n2958) );
  AND U2942 ( .A(n2969), .B(n2970), .Z(n2968) );
  XOR U2943 ( .A(n2967), .B(n2083), .Z(n2970) );
  XNOR U2944 ( .A(p_input[91]), .B(n2971), .Z(n2083) );
  AND U2945 ( .A(n202), .B(n2972), .Z(n2971) );
  XOR U2946 ( .A(p_input[91]), .B(p_input[123]), .Z(n2972) );
  XNOR U2947 ( .A(n2080), .B(n2967), .Z(n2969) );
  XOR U2948 ( .A(n2973), .B(n2974), .Z(n2080) );
  AND U2949 ( .A(n199), .B(n2975), .Z(n2974) );
  XOR U2950 ( .A(p_input[59]), .B(p_input[27]), .Z(n2975) );
  XOR U2951 ( .A(n2976), .B(n2977), .Z(n2967) );
  AND U2952 ( .A(n2978), .B(n2979), .Z(n2977) );
  XOR U2953 ( .A(n2976), .B(n2095), .Z(n2979) );
  XNOR U2954 ( .A(p_input[90]), .B(n2980), .Z(n2095) );
  AND U2955 ( .A(n202), .B(n2981), .Z(n2980) );
  XOR U2956 ( .A(p_input[90]), .B(p_input[122]), .Z(n2981) );
  XNOR U2957 ( .A(n2092), .B(n2976), .Z(n2978) );
  XOR U2958 ( .A(n2982), .B(n2983), .Z(n2092) );
  AND U2959 ( .A(n199), .B(n2984), .Z(n2983) );
  XOR U2960 ( .A(p_input[58]), .B(p_input[26]), .Z(n2984) );
  XOR U2961 ( .A(n2985), .B(n2986), .Z(n2976) );
  AND U2962 ( .A(n2987), .B(n2988), .Z(n2986) );
  XOR U2963 ( .A(n2985), .B(n2107), .Z(n2988) );
  XNOR U2964 ( .A(p_input[89]), .B(n2989), .Z(n2107) );
  AND U2965 ( .A(n202), .B(n2990), .Z(n2989) );
  XOR U2966 ( .A(p_input[89]), .B(p_input[121]), .Z(n2990) );
  XNOR U2967 ( .A(n2104), .B(n2985), .Z(n2987) );
  XOR U2968 ( .A(n2991), .B(n2992), .Z(n2104) );
  AND U2969 ( .A(n199), .B(n2993), .Z(n2992) );
  XOR U2970 ( .A(p_input[57]), .B(p_input[25]), .Z(n2993) );
  XOR U2971 ( .A(n2994), .B(n2995), .Z(n2985) );
  AND U2972 ( .A(n2996), .B(n2997), .Z(n2995) );
  XOR U2973 ( .A(n2994), .B(n2119), .Z(n2997) );
  XNOR U2974 ( .A(p_input[88]), .B(n2998), .Z(n2119) );
  AND U2975 ( .A(n202), .B(n2999), .Z(n2998) );
  XOR U2976 ( .A(p_input[88]), .B(p_input[120]), .Z(n2999) );
  XNOR U2977 ( .A(n2116), .B(n2994), .Z(n2996) );
  XOR U2978 ( .A(n3000), .B(n3001), .Z(n2116) );
  AND U2979 ( .A(n199), .B(n3002), .Z(n3001) );
  XOR U2980 ( .A(p_input[56]), .B(p_input[24]), .Z(n3002) );
  XOR U2981 ( .A(n3003), .B(n3004), .Z(n2994) );
  AND U2982 ( .A(n3005), .B(n3006), .Z(n3004) );
  XOR U2983 ( .A(n3003), .B(n2131), .Z(n3006) );
  XNOR U2984 ( .A(p_input[87]), .B(n3007), .Z(n2131) );
  AND U2985 ( .A(n202), .B(n3008), .Z(n3007) );
  XOR U2986 ( .A(p_input[87]), .B(p_input[119]), .Z(n3008) );
  XNOR U2987 ( .A(n2128), .B(n3003), .Z(n3005) );
  XOR U2988 ( .A(n3009), .B(n3010), .Z(n2128) );
  AND U2989 ( .A(n199), .B(n3011), .Z(n3010) );
  XOR U2990 ( .A(p_input[55]), .B(p_input[23]), .Z(n3011) );
  XOR U2991 ( .A(n3012), .B(n3013), .Z(n3003) );
  AND U2992 ( .A(n3014), .B(n3015), .Z(n3013) );
  XOR U2993 ( .A(n3012), .B(n2143), .Z(n3015) );
  XNOR U2994 ( .A(p_input[86]), .B(n3016), .Z(n2143) );
  AND U2995 ( .A(n202), .B(n3017), .Z(n3016) );
  XOR U2996 ( .A(p_input[86]), .B(p_input[118]), .Z(n3017) );
  XNOR U2997 ( .A(n2140), .B(n3012), .Z(n3014) );
  XOR U2998 ( .A(n3018), .B(n3019), .Z(n2140) );
  AND U2999 ( .A(n199), .B(n3020), .Z(n3019) );
  XOR U3000 ( .A(p_input[54]), .B(p_input[22]), .Z(n3020) );
  XOR U3001 ( .A(n3021), .B(n3022), .Z(n3012) );
  AND U3002 ( .A(n3023), .B(n3024), .Z(n3022) );
  XOR U3003 ( .A(n3021), .B(n2155), .Z(n3024) );
  XNOR U3004 ( .A(p_input[85]), .B(n3025), .Z(n2155) );
  AND U3005 ( .A(n202), .B(n3026), .Z(n3025) );
  XOR U3006 ( .A(p_input[85]), .B(p_input[117]), .Z(n3026) );
  XNOR U3007 ( .A(n2152), .B(n3021), .Z(n3023) );
  XOR U3008 ( .A(n3027), .B(n3028), .Z(n2152) );
  AND U3009 ( .A(n199), .B(n3029), .Z(n3028) );
  XOR U3010 ( .A(p_input[53]), .B(p_input[21]), .Z(n3029) );
  XOR U3011 ( .A(n3030), .B(n3031), .Z(n3021) );
  AND U3012 ( .A(n3032), .B(n3033), .Z(n3031) );
  XOR U3013 ( .A(n3030), .B(n2167), .Z(n3033) );
  XNOR U3014 ( .A(p_input[84]), .B(n3034), .Z(n2167) );
  AND U3015 ( .A(n202), .B(n3035), .Z(n3034) );
  XOR U3016 ( .A(p_input[84]), .B(p_input[116]), .Z(n3035) );
  XNOR U3017 ( .A(n2164), .B(n3030), .Z(n3032) );
  XOR U3018 ( .A(n3036), .B(n3037), .Z(n2164) );
  AND U3019 ( .A(n199), .B(n3038), .Z(n3037) );
  XOR U3020 ( .A(p_input[52]), .B(p_input[20]), .Z(n3038) );
  XOR U3021 ( .A(n3039), .B(n3040), .Z(n3030) );
  AND U3022 ( .A(n3041), .B(n3042), .Z(n3040) );
  XOR U3023 ( .A(n3039), .B(n2179), .Z(n3042) );
  XNOR U3024 ( .A(p_input[83]), .B(n3043), .Z(n2179) );
  AND U3025 ( .A(n202), .B(n3044), .Z(n3043) );
  XOR U3026 ( .A(p_input[83]), .B(p_input[115]), .Z(n3044) );
  XNOR U3027 ( .A(n2176), .B(n3039), .Z(n3041) );
  XOR U3028 ( .A(n3045), .B(n3046), .Z(n2176) );
  AND U3029 ( .A(n199), .B(n3047), .Z(n3046) );
  XOR U3030 ( .A(p_input[51]), .B(p_input[19]), .Z(n3047) );
  XOR U3031 ( .A(n3048), .B(n3049), .Z(n3039) );
  AND U3032 ( .A(n3050), .B(n3051), .Z(n3049) );
  XOR U3033 ( .A(n3048), .B(n2191), .Z(n3051) );
  XNOR U3034 ( .A(p_input[82]), .B(n3052), .Z(n2191) );
  AND U3035 ( .A(n202), .B(n3053), .Z(n3052) );
  XOR U3036 ( .A(p_input[82]), .B(p_input[114]), .Z(n3053) );
  XNOR U3037 ( .A(n2188), .B(n3048), .Z(n3050) );
  XOR U3038 ( .A(n3054), .B(n3055), .Z(n2188) );
  AND U3039 ( .A(n199), .B(n3056), .Z(n3055) );
  XOR U3040 ( .A(p_input[50]), .B(p_input[18]), .Z(n3056) );
  XOR U3041 ( .A(n3057), .B(n3058), .Z(n3048) );
  AND U3042 ( .A(n3059), .B(n3060), .Z(n3058) );
  XOR U3043 ( .A(n3057), .B(n2203), .Z(n3060) );
  XNOR U3044 ( .A(p_input[81]), .B(n3061), .Z(n2203) );
  AND U3045 ( .A(n202), .B(n3062), .Z(n3061) );
  XOR U3046 ( .A(p_input[81]), .B(p_input[113]), .Z(n3062) );
  XNOR U3047 ( .A(n2200), .B(n3057), .Z(n3059) );
  XOR U3048 ( .A(n3063), .B(n3064), .Z(n2200) );
  AND U3049 ( .A(n199), .B(n3065), .Z(n3064) );
  XOR U3050 ( .A(p_input[49]), .B(p_input[17]), .Z(n3065) );
  XOR U3051 ( .A(n3066), .B(n3067), .Z(n3057) );
  AND U3052 ( .A(n3068), .B(n3069), .Z(n3067) );
  XOR U3053 ( .A(n3066), .B(n2215), .Z(n3069) );
  XNOR U3054 ( .A(p_input[80]), .B(n3070), .Z(n2215) );
  AND U3055 ( .A(n202), .B(n3071), .Z(n3070) );
  XOR U3056 ( .A(p_input[80]), .B(p_input[112]), .Z(n3071) );
  XNOR U3057 ( .A(n2212), .B(n3066), .Z(n3068) );
  XOR U3058 ( .A(n3072), .B(n3073), .Z(n2212) );
  AND U3059 ( .A(n199), .B(n3074), .Z(n3073) );
  XOR U3060 ( .A(p_input[48]), .B(p_input[16]), .Z(n3074) );
  XOR U3061 ( .A(n3075), .B(n3076), .Z(n3066) );
  AND U3062 ( .A(n3077), .B(n3078), .Z(n3076) );
  XOR U3063 ( .A(n3075), .B(n2227), .Z(n3078) );
  XNOR U3064 ( .A(p_input[79]), .B(n3079), .Z(n2227) );
  AND U3065 ( .A(n202), .B(n3080), .Z(n3079) );
  XOR U3066 ( .A(p_input[79]), .B(p_input[111]), .Z(n3080) );
  XNOR U3067 ( .A(n2224), .B(n3075), .Z(n3077) );
  XOR U3068 ( .A(n3081), .B(n3082), .Z(n2224) );
  AND U3069 ( .A(n199), .B(n3083), .Z(n3082) );
  XOR U3070 ( .A(p_input[47]), .B(p_input[15]), .Z(n3083) );
  XOR U3071 ( .A(n3084), .B(n3085), .Z(n3075) );
  AND U3072 ( .A(n3086), .B(n3087), .Z(n3085) );
  XOR U3073 ( .A(n3084), .B(n2239), .Z(n3087) );
  XNOR U3074 ( .A(p_input[78]), .B(n3088), .Z(n2239) );
  AND U3075 ( .A(n202), .B(n3089), .Z(n3088) );
  XOR U3076 ( .A(p_input[78]), .B(p_input[110]), .Z(n3089) );
  XNOR U3077 ( .A(n2236), .B(n3084), .Z(n3086) );
  XOR U3078 ( .A(n3090), .B(n3091), .Z(n2236) );
  AND U3079 ( .A(n199), .B(n3092), .Z(n3091) );
  XOR U3080 ( .A(p_input[46]), .B(p_input[14]), .Z(n3092) );
  XOR U3081 ( .A(n3093), .B(n3094), .Z(n3084) );
  AND U3082 ( .A(n3095), .B(n3096), .Z(n3094) );
  XOR U3083 ( .A(n3093), .B(n2251), .Z(n3096) );
  XNOR U3084 ( .A(p_input[77]), .B(n3097), .Z(n2251) );
  AND U3085 ( .A(n202), .B(n3098), .Z(n3097) );
  XOR U3086 ( .A(p_input[77]), .B(p_input[109]), .Z(n3098) );
  XNOR U3087 ( .A(n2248), .B(n3093), .Z(n3095) );
  XOR U3088 ( .A(n3099), .B(n3100), .Z(n2248) );
  AND U3089 ( .A(n199), .B(n3101), .Z(n3100) );
  XOR U3090 ( .A(p_input[45]), .B(p_input[13]), .Z(n3101) );
  XOR U3091 ( .A(n3102), .B(n3103), .Z(n3093) );
  AND U3092 ( .A(n3104), .B(n3105), .Z(n3103) );
  XOR U3093 ( .A(n3102), .B(n2263), .Z(n3105) );
  XNOR U3094 ( .A(p_input[76]), .B(n3106), .Z(n2263) );
  AND U3095 ( .A(n202), .B(n3107), .Z(n3106) );
  XOR U3096 ( .A(p_input[76]), .B(p_input[108]), .Z(n3107) );
  XNOR U3097 ( .A(n2260), .B(n3102), .Z(n3104) );
  XOR U3098 ( .A(n3108), .B(n3109), .Z(n2260) );
  AND U3099 ( .A(n199), .B(n3110), .Z(n3109) );
  XOR U3100 ( .A(p_input[44]), .B(p_input[12]), .Z(n3110) );
  XOR U3101 ( .A(n3111), .B(n3112), .Z(n3102) );
  AND U3102 ( .A(n3113), .B(n3114), .Z(n3112) );
  XOR U3103 ( .A(n3111), .B(n2275), .Z(n3114) );
  XNOR U3104 ( .A(p_input[75]), .B(n3115), .Z(n2275) );
  AND U3105 ( .A(n202), .B(n3116), .Z(n3115) );
  XOR U3106 ( .A(p_input[75]), .B(p_input[107]), .Z(n3116) );
  XNOR U3107 ( .A(n2272), .B(n3111), .Z(n3113) );
  XOR U3108 ( .A(n3117), .B(n3118), .Z(n2272) );
  AND U3109 ( .A(n199), .B(n3119), .Z(n3118) );
  XOR U3110 ( .A(p_input[43]), .B(p_input[11]), .Z(n3119) );
  XOR U3111 ( .A(n3120), .B(n3121), .Z(n3111) );
  AND U3112 ( .A(n3122), .B(n3123), .Z(n3121) );
  XOR U3113 ( .A(n3120), .B(n2287), .Z(n3123) );
  XNOR U3114 ( .A(p_input[74]), .B(n3124), .Z(n2287) );
  AND U3115 ( .A(n202), .B(n3125), .Z(n3124) );
  XOR U3116 ( .A(p_input[74]), .B(p_input[106]), .Z(n3125) );
  XNOR U3117 ( .A(n2284), .B(n3120), .Z(n3122) );
  XOR U3118 ( .A(n3126), .B(n3127), .Z(n2284) );
  AND U3119 ( .A(n199), .B(n3128), .Z(n3127) );
  XOR U3120 ( .A(p_input[42]), .B(p_input[10]), .Z(n3128) );
  XOR U3121 ( .A(n3129), .B(n3130), .Z(n3120) );
  AND U3122 ( .A(n3131), .B(n3132), .Z(n3130) );
  XOR U3123 ( .A(n3129), .B(n2299), .Z(n3132) );
  XNOR U3124 ( .A(p_input[73]), .B(n3133), .Z(n2299) );
  AND U3125 ( .A(n202), .B(n3134), .Z(n3133) );
  XOR U3126 ( .A(p_input[73]), .B(p_input[105]), .Z(n3134) );
  XNOR U3127 ( .A(n2296), .B(n3129), .Z(n3131) );
  XOR U3128 ( .A(n3135), .B(n3136), .Z(n2296) );
  AND U3129 ( .A(n199), .B(n3137), .Z(n3136) );
  XOR U3130 ( .A(p_input[9]), .B(p_input[41]), .Z(n3137) );
  XOR U3131 ( .A(n3138), .B(n3139), .Z(n3129) );
  AND U3132 ( .A(n3140), .B(n3141), .Z(n3139) );
  XOR U3133 ( .A(n3138), .B(n2311), .Z(n3141) );
  XNOR U3134 ( .A(p_input[72]), .B(n3142), .Z(n2311) );
  AND U3135 ( .A(n202), .B(n3143), .Z(n3142) );
  XOR U3136 ( .A(p_input[72]), .B(p_input[104]), .Z(n3143) );
  XNOR U3137 ( .A(n2308), .B(n3138), .Z(n3140) );
  XOR U3138 ( .A(n3144), .B(n3145), .Z(n2308) );
  AND U3139 ( .A(n199), .B(n3146), .Z(n3145) );
  XOR U3140 ( .A(p_input[8]), .B(p_input[40]), .Z(n3146) );
  XOR U3141 ( .A(n3147), .B(n3148), .Z(n3138) );
  AND U3142 ( .A(n3149), .B(n3150), .Z(n3148) );
  XOR U3143 ( .A(n3147), .B(n2323), .Z(n3150) );
  XNOR U3144 ( .A(p_input[71]), .B(n3151), .Z(n2323) );
  AND U3145 ( .A(n202), .B(n3152), .Z(n3151) );
  XOR U3146 ( .A(p_input[71]), .B(p_input[103]), .Z(n3152) );
  XNOR U3147 ( .A(n2320), .B(n3147), .Z(n3149) );
  XOR U3148 ( .A(n3153), .B(n3154), .Z(n2320) );
  AND U3149 ( .A(n199), .B(n3155), .Z(n3154) );
  XOR U3150 ( .A(p_input[7]), .B(p_input[39]), .Z(n3155) );
  XOR U3151 ( .A(n3156), .B(n3157), .Z(n3147) );
  AND U3152 ( .A(n3158), .B(n3159), .Z(n3157) );
  XOR U3153 ( .A(n3156), .B(n2335), .Z(n3159) );
  XNOR U3154 ( .A(p_input[70]), .B(n3160), .Z(n2335) );
  AND U3155 ( .A(n202), .B(n3161), .Z(n3160) );
  XOR U3156 ( .A(p_input[70]), .B(p_input[102]), .Z(n3161) );
  XNOR U3157 ( .A(n2332), .B(n3156), .Z(n3158) );
  XOR U3158 ( .A(n3162), .B(n3163), .Z(n2332) );
  AND U3159 ( .A(n199), .B(n3164), .Z(n3163) );
  XOR U3160 ( .A(p_input[6]), .B(p_input[38]), .Z(n3164) );
  XOR U3161 ( .A(n3165), .B(n3166), .Z(n3156) );
  AND U3162 ( .A(n3167), .B(n3168), .Z(n3166) );
  XOR U3163 ( .A(n2347), .B(n3165), .Z(n3168) );
  XNOR U3164 ( .A(p_input[69]), .B(n3169), .Z(n2347) );
  AND U3165 ( .A(n202), .B(n3170), .Z(n3169) );
  XOR U3166 ( .A(p_input[69]), .B(p_input[101]), .Z(n3170) );
  XNOR U3167 ( .A(n3165), .B(n2344), .Z(n3167) );
  XOR U3168 ( .A(n3171), .B(n3172), .Z(n2344) );
  AND U3169 ( .A(n199), .B(n3173), .Z(n3172) );
  XOR U3170 ( .A(p_input[5]), .B(p_input[37]), .Z(n3173) );
  XOR U3171 ( .A(n3174), .B(n3175), .Z(n3165) );
  AND U3172 ( .A(n3176), .B(n3177), .Z(n3175) );
  XOR U3173 ( .A(n3174), .B(n2359), .Z(n3177) );
  XNOR U3174 ( .A(p_input[68]), .B(n3178), .Z(n2359) );
  AND U3175 ( .A(n202), .B(n3179), .Z(n3178) );
  XOR U3176 ( .A(p_input[68]), .B(p_input[100]), .Z(n3179) );
  XNOR U3177 ( .A(n2356), .B(n3174), .Z(n3176) );
  XOR U3178 ( .A(n3180), .B(n3181), .Z(n2356) );
  AND U3179 ( .A(n199), .B(n3182), .Z(n3181) );
  XOR U3180 ( .A(p_input[4]), .B(p_input[36]), .Z(n3182) );
  XOR U3181 ( .A(n3183), .B(n3184), .Z(n3174) );
  AND U3182 ( .A(n3185), .B(n3186), .Z(n3184) );
  XOR U3183 ( .A(n3183), .B(n2371), .Z(n3186) );
  XNOR U3184 ( .A(p_input[67]), .B(n3187), .Z(n2371) );
  AND U3185 ( .A(n202), .B(n3188), .Z(n3187) );
  XOR U3186 ( .A(p_input[99]), .B(p_input[67]), .Z(n3188) );
  XNOR U3187 ( .A(n2368), .B(n3183), .Z(n3185) );
  XOR U3188 ( .A(n3189), .B(n3190), .Z(n2368) );
  AND U3189 ( .A(n199), .B(n3191), .Z(n3190) );
  XOR U3190 ( .A(p_input[3]), .B(p_input[35]), .Z(n3191) );
  XOR U3191 ( .A(n3192), .B(n3193), .Z(n3183) );
  AND U3192 ( .A(n3194), .B(n3195), .Z(n3193) );
  XOR U3193 ( .A(n3192), .B(n2383), .Z(n3195) );
  XNOR U3194 ( .A(p_input[66]), .B(n3196), .Z(n2383) );
  AND U3195 ( .A(n202), .B(n3197), .Z(n3196) );
  XOR U3196 ( .A(p_input[98]), .B(p_input[66]), .Z(n3197) );
  XNOR U3197 ( .A(n2380), .B(n3192), .Z(n3194) );
  XOR U3198 ( .A(n3198), .B(n3199), .Z(n2380) );
  AND U3199 ( .A(n199), .B(n3200), .Z(n3199) );
  XOR U3200 ( .A(p_input[34]), .B(p_input[2]), .Z(n3200) );
  XOR U3201 ( .A(n3201), .B(n3202), .Z(n3192) );
  AND U3202 ( .A(n3203), .B(n3204), .Z(n3202) );
  XNOR U3203 ( .A(n3205), .B(n2396), .Z(n3204) );
  XNOR U3204 ( .A(p_input[65]), .B(n3206), .Z(n2396) );
  AND U3205 ( .A(n202), .B(n3207), .Z(n3206) );
  XNOR U3206 ( .A(p_input[97]), .B(n3208), .Z(n3207) );
  IV U3207 ( .A(p_input[65]), .Z(n3208) );
  XNOR U3208 ( .A(n2393), .B(n3201), .Z(n3203) );
  XNOR U3209 ( .A(p_input[1]), .B(n3209), .Z(n2393) );
  AND U3210 ( .A(n199), .B(n3210), .Z(n3209) );
  XOR U3211 ( .A(p_input[33]), .B(p_input[1]), .Z(n3210) );
  IV U3212 ( .A(n3205), .Z(n3201) );
  AND U3213 ( .A(n2931), .B(n2934), .Z(n3205) );
  XOR U3214 ( .A(p_input[64]), .B(n3211), .Z(n2934) );
  AND U3215 ( .A(n202), .B(n3212), .Z(n3211) );
  XOR U3216 ( .A(p_input[96]), .B(p_input[64]), .Z(n3212) );
  XOR U3217 ( .A(n3213), .B(n3214), .Z(n202) );
  AND U3218 ( .A(n3215), .B(n3216), .Z(n3214) );
  XNOR U3219 ( .A(p_input[127]), .B(n3213), .Z(n3216) );
  XOR U3220 ( .A(n3213), .B(p_input[95]), .Z(n3215) );
  XOR U3221 ( .A(n3217), .B(n3218), .Z(n3213) );
  AND U3222 ( .A(n3219), .B(n3220), .Z(n3218) );
  XNOR U3223 ( .A(p_input[126]), .B(n3217), .Z(n3220) );
  XOR U3224 ( .A(n3217), .B(p_input[94]), .Z(n3219) );
  XOR U3225 ( .A(n3221), .B(n3222), .Z(n3217) );
  AND U3226 ( .A(n3223), .B(n3224), .Z(n3222) );
  XNOR U3227 ( .A(p_input[125]), .B(n3221), .Z(n3224) );
  XOR U3228 ( .A(n3221), .B(p_input[93]), .Z(n3223) );
  XOR U3229 ( .A(n3225), .B(n3226), .Z(n3221) );
  AND U3230 ( .A(n3227), .B(n3228), .Z(n3226) );
  XNOR U3231 ( .A(p_input[124]), .B(n3225), .Z(n3228) );
  XOR U3232 ( .A(n3225), .B(p_input[92]), .Z(n3227) );
  XOR U3233 ( .A(n3229), .B(n3230), .Z(n3225) );
  AND U3234 ( .A(n3231), .B(n3232), .Z(n3230) );
  XNOR U3235 ( .A(p_input[123]), .B(n3229), .Z(n3232) );
  XOR U3236 ( .A(n3229), .B(p_input[91]), .Z(n3231) );
  XOR U3237 ( .A(n3233), .B(n3234), .Z(n3229) );
  AND U3238 ( .A(n3235), .B(n3236), .Z(n3234) );
  XNOR U3239 ( .A(p_input[122]), .B(n3233), .Z(n3236) );
  XOR U3240 ( .A(n3233), .B(p_input[90]), .Z(n3235) );
  XOR U3241 ( .A(n3237), .B(n3238), .Z(n3233) );
  AND U3242 ( .A(n3239), .B(n3240), .Z(n3238) );
  XNOR U3243 ( .A(p_input[121]), .B(n3237), .Z(n3240) );
  XOR U3244 ( .A(n3237), .B(p_input[89]), .Z(n3239) );
  XOR U3245 ( .A(n3241), .B(n3242), .Z(n3237) );
  AND U3246 ( .A(n3243), .B(n3244), .Z(n3242) );
  XNOR U3247 ( .A(p_input[120]), .B(n3241), .Z(n3244) );
  XOR U3248 ( .A(n3241), .B(p_input[88]), .Z(n3243) );
  XOR U3249 ( .A(n3245), .B(n3246), .Z(n3241) );
  AND U3250 ( .A(n3247), .B(n3248), .Z(n3246) );
  XNOR U3251 ( .A(p_input[119]), .B(n3245), .Z(n3248) );
  XOR U3252 ( .A(n3245), .B(p_input[87]), .Z(n3247) );
  XOR U3253 ( .A(n3249), .B(n3250), .Z(n3245) );
  AND U3254 ( .A(n3251), .B(n3252), .Z(n3250) );
  XNOR U3255 ( .A(p_input[118]), .B(n3249), .Z(n3252) );
  XOR U3256 ( .A(n3249), .B(p_input[86]), .Z(n3251) );
  XOR U3257 ( .A(n3253), .B(n3254), .Z(n3249) );
  AND U3258 ( .A(n3255), .B(n3256), .Z(n3254) );
  XNOR U3259 ( .A(p_input[117]), .B(n3253), .Z(n3256) );
  XOR U3260 ( .A(n3253), .B(p_input[85]), .Z(n3255) );
  XOR U3261 ( .A(n3257), .B(n3258), .Z(n3253) );
  AND U3262 ( .A(n3259), .B(n3260), .Z(n3258) );
  XNOR U3263 ( .A(p_input[116]), .B(n3257), .Z(n3260) );
  XOR U3264 ( .A(n3257), .B(p_input[84]), .Z(n3259) );
  XOR U3265 ( .A(n3261), .B(n3262), .Z(n3257) );
  AND U3266 ( .A(n3263), .B(n3264), .Z(n3262) );
  XNOR U3267 ( .A(p_input[115]), .B(n3261), .Z(n3264) );
  XOR U3268 ( .A(n3261), .B(p_input[83]), .Z(n3263) );
  XOR U3269 ( .A(n3265), .B(n3266), .Z(n3261) );
  AND U3270 ( .A(n3267), .B(n3268), .Z(n3266) );
  XNOR U3271 ( .A(p_input[114]), .B(n3265), .Z(n3268) );
  XOR U3272 ( .A(n3265), .B(p_input[82]), .Z(n3267) );
  XOR U3273 ( .A(n3269), .B(n3270), .Z(n3265) );
  AND U3274 ( .A(n3271), .B(n3272), .Z(n3270) );
  XNOR U3275 ( .A(p_input[113]), .B(n3269), .Z(n3272) );
  XOR U3276 ( .A(n3269), .B(p_input[81]), .Z(n3271) );
  XOR U3277 ( .A(n3273), .B(n3274), .Z(n3269) );
  AND U3278 ( .A(n3275), .B(n3276), .Z(n3274) );
  XNOR U3279 ( .A(p_input[112]), .B(n3273), .Z(n3276) );
  XOR U3280 ( .A(n3273), .B(p_input[80]), .Z(n3275) );
  XOR U3281 ( .A(n3277), .B(n3278), .Z(n3273) );
  AND U3282 ( .A(n3279), .B(n3280), .Z(n3278) );
  XNOR U3283 ( .A(p_input[111]), .B(n3277), .Z(n3280) );
  XOR U3284 ( .A(n3277), .B(p_input[79]), .Z(n3279) );
  XOR U3285 ( .A(n3281), .B(n3282), .Z(n3277) );
  AND U3286 ( .A(n3283), .B(n3284), .Z(n3282) );
  XNOR U3287 ( .A(p_input[110]), .B(n3281), .Z(n3284) );
  XOR U3288 ( .A(n3281), .B(p_input[78]), .Z(n3283) );
  XOR U3289 ( .A(n3285), .B(n3286), .Z(n3281) );
  AND U3290 ( .A(n3287), .B(n3288), .Z(n3286) );
  XNOR U3291 ( .A(p_input[109]), .B(n3285), .Z(n3288) );
  XOR U3292 ( .A(n3285), .B(p_input[77]), .Z(n3287) );
  XOR U3293 ( .A(n3289), .B(n3290), .Z(n3285) );
  AND U3294 ( .A(n3291), .B(n3292), .Z(n3290) );
  XNOR U3295 ( .A(p_input[108]), .B(n3289), .Z(n3292) );
  XOR U3296 ( .A(n3289), .B(p_input[76]), .Z(n3291) );
  XOR U3297 ( .A(n3293), .B(n3294), .Z(n3289) );
  AND U3298 ( .A(n3295), .B(n3296), .Z(n3294) );
  XNOR U3299 ( .A(p_input[107]), .B(n3293), .Z(n3296) );
  XOR U3300 ( .A(n3293), .B(p_input[75]), .Z(n3295) );
  XOR U3301 ( .A(n3297), .B(n3298), .Z(n3293) );
  AND U3302 ( .A(n3299), .B(n3300), .Z(n3298) );
  XNOR U3303 ( .A(p_input[106]), .B(n3297), .Z(n3300) );
  XOR U3304 ( .A(n3297), .B(p_input[74]), .Z(n3299) );
  XOR U3305 ( .A(n3301), .B(n3302), .Z(n3297) );
  AND U3306 ( .A(n3303), .B(n3304), .Z(n3302) );
  XNOR U3307 ( .A(p_input[105]), .B(n3301), .Z(n3304) );
  XOR U3308 ( .A(n3301), .B(p_input[73]), .Z(n3303) );
  XOR U3309 ( .A(n3305), .B(n3306), .Z(n3301) );
  AND U3310 ( .A(n3307), .B(n3308), .Z(n3306) );
  XNOR U3311 ( .A(p_input[104]), .B(n3305), .Z(n3308) );
  XOR U3312 ( .A(n3305), .B(p_input[72]), .Z(n3307) );
  XOR U3313 ( .A(n3309), .B(n3310), .Z(n3305) );
  AND U3314 ( .A(n3311), .B(n3312), .Z(n3310) );
  XNOR U3315 ( .A(p_input[103]), .B(n3309), .Z(n3312) );
  XOR U3316 ( .A(n3309), .B(p_input[71]), .Z(n3311) );
  XOR U3317 ( .A(n3313), .B(n3314), .Z(n3309) );
  AND U3318 ( .A(n3315), .B(n3316), .Z(n3314) );
  XNOR U3319 ( .A(p_input[102]), .B(n3313), .Z(n3316) );
  XOR U3320 ( .A(n3313), .B(p_input[70]), .Z(n3315) );
  XOR U3321 ( .A(n3317), .B(n3318), .Z(n3313) );
  AND U3322 ( .A(n3319), .B(n3320), .Z(n3318) );
  XNOR U3323 ( .A(p_input[101]), .B(n3317), .Z(n3320) );
  XOR U3324 ( .A(n3317), .B(p_input[69]), .Z(n3319) );
  XOR U3325 ( .A(n3321), .B(n3322), .Z(n3317) );
  AND U3326 ( .A(n3323), .B(n3324), .Z(n3322) );
  XNOR U3327 ( .A(p_input[100]), .B(n3321), .Z(n3324) );
  XOR U3328 ( .A(n3321), .B(p_input[68]), .Z(n3323) );
  XOR U3329 ( .A(n3325), .B(n3326), .Z(n3321) );
  AND U3330 ( .A(n3327), .B(n3328), .Z(n3326) );
  XNOR U3331 ( .A(p_input[99]), .B(n3325), .Z(n3328) );
  XOR U3332 ( .A(n3325), .B(p_input[67]), .Z(n3327) );
  XOR U3333 ( .A(n3329), .B(n3330), .Z(n3325) );
  AND U3334 ( .A(n3331), .B(n3332), .Z(n3330) );
  XNOR U3335 ( .A(p_input[98]), .B(n3329), .Z(n3332) );
  XOR U3336 ( .A(n3329), .B(p_input[66]), .Z(n3331) );
  XNOR U3337 ( .A(n3333), .B(n3334), .Z(n3329) );
  AND U3338 ( .A(n3335), .B(n3336), .Z(n3334) );
  XOR U3339 ( .A(p_input[97]), .B(n3333), .Z(n3336) );
  XNOR U3340 ( .A(p_input[65]), .B(n3333), .Z(n3335) );
  AND U3341 ( .A(p_input[96]), .B(n3337), .Z(n3333) );
  IV U3342 ( .A(p_input[64]), .Z(n3337) );
  XNOR U3343 ( .A(p_input[0]), .B(n3338), .Z(n2931) );
  AND U3344 ( .A(n199), .B(n3339), .Z(n3338) );
  XOR U3345 ( .A(p_input[32]), .B(p_input[0]), .Z(n3339) );
  XOR U3346 ( .A(n3340), .B(n3341), .Z(n199) );
  AND U3347 ( .A(n3342), .B(n3343), .Z(n3341) );
  XNOR U3348 ( .A(p_input[63]), .B(n3340), .Z(n3343) );
  XOR U3349 ( .A(n3340), .B(p_input[31]), .Z(n3342) );
  XOR U3350 ( .A(n3344), .B(n3345), .Z(n3340) );
  AND U3351 ( .A(n3346), .B(n3347), .Z(n3345) );
  XNOR U3352 ( .A(p_input[62]), .B(n3344), .Z(n3347) );
  XNOR U3353 ( .A(n3344), .B(n2946), .Z(n3346) );
  IV U3354 ( .A(p_input[30]), .Z(n2946) );
  XOR U3355 ( .A(n3348), .B(n3349), .Z(n3344) );
  AND U3356 ( .A(n3350), .B(n3351), .Z(n3349) );
  XNOR U3357 ( .A(p_input[61]), .B(n3348), .Z(n3351) );
  XNOR U3358 ( .A(n3348), .B(n2955), .Z(n3350) );
  IV U3359 ( .A(p_input[29]), .Z(n2955) );
  XOR U3360 ( .A(n3352), .B(n3353), .Z(n3348) );
  AND U3361 ( .A(n3354), .B(n3355), .Z(n3353) );
  XNOR U3362 ( .A(p_input[60]), .B(n3352), .Z(n3355) );
  XNOR U3363 ( .A(n3352), .B(n2964), .Z(n3354) );
  IV U3364 ( .A(p_input[28]), .Z(n2964) );
  XOR U3365 ( .A(n3356), .B(n3357), .Z(n3352) );
  AND U3366 ( .A(n3358), .B(n3359), .Z(n3357) );
  XNOR U3367 ( .A(p_input[59]), .B(n3356), .Z(n3359) );
  XNOR U3368 ( .A(n3356), .B(n2973), .Z(n3358) );
  IV U3369 ( .A(p_input[27]), .Z(n2973) );
  XOR U3370 ( .A(n3360), .B(n3361), .Z(n3356) );
  AND U3371 ( .A(n3362), .B(n3363), .Z(n3361) );
  XNOR U3372 ( .A(p_input[58]), .B(n3360), .Z(n3363) );
  XNOR U3373 ( .A(n3360), .B(n2982), .Z(n3362) );
  IV U3374 ( .A(p_input[26]), .Z(n2982) );
  XOR U3375 ( .A(n3364), .B(n3365), .Z(n3360) );
  AND U3376 ( .A(n3366), .B(n3367), .Z(n3365) );
  XNOR U3377 ( .A(p_input[57]), .B(n3364), .Z(n3367) );
  XNOR U3378 ( .A(n3364), .B(n2991), .Z(n3366) );
  IV U3379 ( .A(p_input[25]), .Z(n2991) );
  XOR U3380 ( .A(n3368), .B(n3369), .Z(n3364) );
  AND U3381 ( .A(n3370), .B(n3371), .Z(n3369) );
  XNOR U3382 ( .A(p_input[56]), .B(n3368), .Z(n3371) );
  XNOR U3383 ( .A(n3368), .B(n3000), .Z(n3370) );
  IV U3384 ( .A(p_input[24]), .Z(n3000) );
  XOR U3385 ( .A(n3372), .B(n3373), .Z(n3368) );
  AND U3386 ( .A(n3374), .B(n3375), .Z(n3373) );
  XNOR U3387 ( .A(p_input[55]), .B(n3372), .Z(n3375) );
  XNOR U3388 ( .A(n3372), .B(n3009), .Z(n3374) );
  IV U3389 ( .A(p_input[23]), .Z(n3009) );
  XOR U3390 ( .A(n3376), .B(n3377), .Z(n3372) );
  AND U3391 ( .A(n3378), .B(n3379), .Z(n3377) );
  XNOR U3392 ( .A(p_input[54]), .B(n3376), .Z(n3379) );
  XNOR U3393 ( .A(n3376), .B(n3018), .Z(n3378) );
  IV U3394 ( .A(p_input[22]), .Z(n3018) );
  XOR U3395 ( .A(n3380), .B(n3381), .Z(n3376) );
  AND U3396 ( .A(n3382), .B(n3383), .Z(n3381) );
  XNOR U3397 ( .A(p_input[53]), .B(n3380), .Z(n3383) );
  XNOR U3398 ( .A(n3380), .B(n3027), .Z(n3382) );
  IV U3399 ( .A(p_input[21]), .Z(n3027) );
  XOR U3400 ( .A(n3384), .B(n3385), .Z(n3380) );
  AND U3401 ( .A(n3386), .B(n3387), .Z(n3385) );
  XNOR U3402 ( .A(p_input[52]), .B(n3384), .Z(n3387) );
  XNOR U3403 ( .A(n3384), .B(n3036), .Z(n3386) );
  IV U3404 ( .A(p_input[20]), .Z(n3036) );
  XOR U3405 ( .A(n3388), .B(n3389), .Z(n3384) );
  AND U3406 ( .A(n3390), .B(n3391), .Z(n3389) );
  XNOR U3407 ( .A(p_input[51]), .B(n3388), .Z(n3391) );
  XNOR U3408 ( .A(n3388), .B(n3045), .Z(n3390) );
  IV U3409 ( .A(p_input[19]), .Z(n3045) );
  XOR U3410 ( .A(n3392), .B(n3393), .Z(n3388) );
  AND U3411 ( .A(n3394), .B(n3395), .Z(n3393) );
  XNOR U3412 ( .A(p_input[50]), .B(n3392), .Z(n3395) );
  XNOR U3413 ( .A(n3392), .B(n3054), .Z(n3394) );
  IV U3414 ( .A(p_input[18]), .Z(n3054) );
  XOR U3415 ( .A(n3396), .B(n3397), .Z(n3392) );
  AND U3416 ( .A(n3398), .B(n3399), .Z(n3397) );
  XNOR U3417 ( .A(p_input[49]), .B(n3396), .Z(n3399) );
  XNOR U3418 ( .A(n3396), .B(n3063), .Z(n3398) );
  IV U3419 ( .A(p_input[17]), .Z(n3063) );
  XOR U3420 ( .A(n3400), .B(n3401), .Z(n3396) );
  AND U3421 ( .A(n3402), .B(n3403), .Z(n3401) );
  XNOR U3422 ( .A(p_input[48]), .B(n3400), .Z(n3403) );
  XNOR U3423 ( .A(n3400), .B(n3072), .Z(n3402) );
  IV U3424 ( .A(p_input[16]), .Z(n3072) );
  XOR U3425 ( .A(n3404), .B(n3405), .Z(n3400) );
  AND U3426 ( .A(n3406), .B(n3407), .Z(n3405) );
  XNOR U3427 ( .A(p_input[47]), .B(n3404), .Z(n3407) );
  XNOR U3428 ( .A(n3404), .B(n3081), .Z(n3406) );
  IV U3429 ( .A(p_input[15]), .Z(n3081) );
  XOR U3430 ( .A(n3408), .B(n3409), .Z(n3404) );
  AND U3431 ( .A(n3410), .B(n3411), .Z(n3409) );
  XNOR U3432 ( .A(p_input[46]), .B(n3408), .Z(n3411) );
  XNOR U3433 ( .A(n3408), .B(n3090), .Z(n3410) );
  IV U3434 ( .A(p_input[14]), .Z(n3090) );
  XOR U3435 ( .A(n3412), .B(n3413), .Z(n3408) );
  AND U3436 ( .A(n3414), .B(n3415), .Z(n3413) );
  XNOR U3437 ( .A(p_input[45]), .B(n3412), .Z(n3415) );
  XNOR U3438 ( .A(n3412), .B(n3099), .Z(n3414) );
  IV U3439 ( .A(p_input[13]), .Z(n3099) );
  XOR U3440 ( .A(n3416), .B(n3417), .Z(n3412) );
  AND U3441 ( .A(n3418), .B(n3419), .Z(n3417) );
  XNOR U3442 ( .A(p_input[44]), .B(n3416), .Z(n3419) );
  XNOR U3443 ( .A(n3416), .B(n3108), .Z(n3418) );
  IV U3444 ( .A(p_input[12]), .Z(n3108) );
  XOR U3445 ( .A(n3420), .B(n3421), .Z(n3416) );
  AND U3446 ( .A(n3422), .B(n3423), .Z(n3421) );
  XNOR U3447 ( .A(p_input[43]), .B(n3420), .Z(n3423) );
  XNOR U3448 ( .A(n3420), .B(n3117), .Z(n3422) );
  IV U3449 ( .A(p_input[11]), .Z(n3117) );
  XOR U3450 ( .A(n3424), .B(n3425), .Z(n3420) );
  AND U3451 ( .A(n3426), .B(n3427), .Z(n3425) );
  XNOR U3452 ( .A(p_input[42]), .B(n3424), .Z(n3427) );
  XNOR U3453 ( .A(n3424), .B(n3126), .Z(n3426) );
  IV U3454 ( .A(p_input[10]), .Z(n3126) );
  XOR U3455 ( .A(n3428), .B(n3429), .Z(n3424) );
  AND U3456 ( .A(n3430), .B(n3431), .Z(n3429) );
  XNOR U3457 ( .A(p_input[41]), .B(n3428), .Z(n3431) );
  XNOR U3458 ( .A(n3428), .B(n3135), .Z(n3430) );
  IV U3459 ( .A(p_input[9]), .Z(n3135) );
  XOR U3460 ( .A(n3432), .B(n3433), .Z(n3428) );
  AND U3461 ( .A(n3434), .B(n3435), .Z(n3433) );
  XNOR U3462 ( .A(p_input[40]), .B(n3432), .Z(n3435) );
  XNOR U3463 ( .A(n3432), .B(n3144), .Z(n3434) );
  IV U3464 ( .A(p_input[8]), .Z(n3144) );
  XOR U3465 ( .A(n3436), .B(n3437), .Z(n3432) );
  AND U3466 ( .A(n3438), .B(n3439), .Z(n3437) );
  XNOR U3467 ( .A(p_input[39]), .B(n3436), .Z(n3439) );
  XNOR U3468 ( .A(n3436), .B(n3153), .Z(n3438) );
  IV U3469 ( .A(p_input[7]), .Z(n3153) );
  XOR U3470 ( .A(n3440), .B(n3441), .Z(n3436) );
  AND U3471 ( .A(n3442), .B(n3443), .Z(n3441) );
  XNOR U3472 ( .A(p_input[38]), .B(n3440), .Z(n3443) );
  XNOR U3473 ( .A(n3440), .B(n3162), .Z(n3442) );
  IV U3474 ( .A(p_input[6]), .Z(n3162) );
  XOR U3475 ( .A(n3444), .B(n3445), .Z(n3440) );
  AND U3476 ( .A(n3446), .B(n3447), .Z(n3445) );
  XNOR U3477 ( .A(p_input[37]), .B(n3444), .Z(n3447) );
  XNOR U3478 ( .A(n3444), .B(n3171), .Z(n3446) );
  IV U3479 ( .A(p_input[5]), .Z(n3171) );
  XOR U3480 ( .A(n3448), .B(n3449), .Z(n3444) );
  AND U3481 ( .A(n3450), .B(n3451), .Z(n3449) );
  XNOR U3482 ( .A(p_input[36]), .B(n3448), .Z(n3451) );
  XNOR U3483 ( .A(n3448), .B(n3180), .Z(n3450) );
  IV U3484 ( .A(p_input[4]), .Z(n3180) );
  XOR U3485 ( .A(n3452), .B(n3453), .Z(n3448) );
  AND U3486 ( .A(n3454), .B(n3455), .Z(n3453) );
  XNOR U3487 ( .A(p_input[35]), .B(n3452), .Z(n3455) );
  XNOR U3488 ( .A(n3452), .B(n3189), .Z(n3454) );
  IV U3489 ( .A(p_input[3]), .Z(n3189) );
  XOR U3490 ( .A(n3456), .B(n3457), .Z(n3452) );
  AND U3491 ( .A(n3458), .B(n3459), .Z(n3457) );
  XNOR U3492 ( .A(p_input[34]), .B(n3456), .Z(n3459) );
  XNOR U3493 ( .A(n3456), .B(n3198), .Z(n3458) );
  IV U3494 ( .A(p_input[2]), .Z(n3198) );
  XNOR U3495 ( .A(n3460), .B(n3461), .Z(n3456) );
  AND U3496 ( .A(n3462), .B(n3463), .Z(n3461) );
  XOR U3497 ( .A(p_input[33]), .B(n3460), .Z(n3463) );
  XNOR U3498 ( .A(p_input[1]), .B(n3460), .Z(n3462) );
  AND U3499 ( .A(p_input[32]), .B(n3464), .Z(n3460) );
  IV U3500 ( .A(p_input[0]), .Z(n3464) );
endmodule

