
module knn_comb_BMR_W16_K1_N8 ( p_input, o );
  input [143:0] p_input;
  output [15:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] , n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158;
  assign \knn_comb_/min_val_out[0][0]  = p_input[112];
  assign \knn_comb_/min_val_out[0][1]  = p_input[113];
  assign \knn_comb_/min_val_out[0][2]  = p_input[114];
  assign \knn_comb_/min_val_out[0][3]  = p_input[115];
  assign \knn_comb_/min_val_out[0][4]  = p_input[116];
  assign \knn_comb_/min_val_out[0][5]  = p_input[117];
  assign \knn_comb_/min_val_out[0][6]  = p_input[118];
  assign \knn_comb_/min_val_out[0][7]  = p_input[119];
  assign \knn_comb_/min_val_out[0][8]  = p_input[120];
  assign \knn_comb_/min_val_out[0][9]  = p_input[121];
  assign \knn_comb_/min_val_out[0][10]  = p_input[122];
  assign \knn_comb_/min_val_out[0][11]  = p_input[123];
  assign \knn_comb_/min_val_out[0][12]  = p_input[124];
  assign \knn_comb_/min_val_out[0][13]  = p_input[125];
  assign \knn_comb_/min_val_out[0][14]  = p_input[126];
  assign \knn_comb_/min_val_out[0][15]  = p_input[127];

  XNOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(n3), .B(n4), .Z(n1) );
  XNOR U3 ( .A(p_input[9]), .B(n2), .Z(n4) );
  XOR U4 ( .A(n5), .B(n6), .Z(n2) );
  AND U5 ( .A(n7), .B(n8), .Z(n6) );
  XNOR U6 ( .A(p_input[25]), .B(n5), .Z(n8) );
  XOR U7 ( .A(n9), .B(n10), .Z(n5) );
  AND U8 ( .A(n11), .B(n12), .Z(n10) );
  XNOR U9 ( .A(p_input[41]), .B(n9), .Z(n12) );
  XOR U10 ( .A(n13), .B(n14), .Z(n9) );
  AND U11 ( .A(n15), .B(n16), .Z(n14) );
  XNOR U12 ( .A(p_input[57]), .B(n13), .Z(n16) );
  XOR U13 ( .A(n17), .B(n18), .Z(n13) );
  AND U14 ( .A(n19), .B(n20), .Z(n18) );
  XNOR U15 ( .A(p_input[73]), .B(n17), .Z(n20) );
  XNOR U16 ( .A(n21), .B(n22), .Z(n17) );
  AND U17 ( .A(n23), .B(n24), .Z(n22) );
  XOR U18 ( .A(p_input[89]), .B(n21), .Z(n24) );
  XOR U19 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n25), .Z(n21) );
  AND U20 ( .A(n26), .B(n27), .Z(n25) );
  XOR U21 ( .A(p_input[105]), .B(\knn_comb_/min_val_out[0][9] ), .Z(n27) );
  XNOR U22 ( .A(n28), .B(n29), .Z(o[8]) );
  AND U23 ( .A(n3), .B(n30), .Z(n28) );
  XNOR U24 ( .A(p_input[8]), .B(n29), .Z(n30) );
  XOR U25 ( .A(n31), .B(n32), .Z(n29) );
  AND U26 ( .A(n7), .B(n33), .Z(n32) );
  XNOR U27 ( .A(p_input[24]), .B(n31), .Z(n33) );
  XOR U28 ( .A(n34), .B(n35), .Z(n31) );
  AND U29 ( .A(n11), .B(n36), .Z(n35) );
  XNOR U30 ( .A(p_input[40]), .B(n34), .Z(n36) );
  XOR U31 ( .A(n37), .B(n38), .Z(n34) );
  AND U32 ( .A(n15), .B(n39), .Z(n38) );
  XNOR U33 ( .A(p_input[56]), .B(n37), .Z(n39) );
  XOR U34 ( .A(n40), .B(n41), .Z(n37) );
  AND U35 ( .A(n19), .B(n42), .Z(n41) );
  XNOR U36 ( .A(p_input[72]), .B(n40), .Z(n42) );
  XNOR U37 ( .A(n43), .B(n44), .Z(n40) );
  AND U38 ( .A(n23), .B(n45), .Z(n44) );
  XOR U39 ( .A(p_input[88]), .B(n43), .Z(n45) );
  XOR U40 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n46), .Z(n43) );
  AND U41 ( .A(n26), .B(n47), .Z(n46) );
  XOR U42 ( .A(p_input[104]), .B(\knn_comb_/min_val_out[0][8] ), .Z(n47) );
  XNOR U43 ( .A(n48), .B(n49), .Z(o[7]) );
  AND U44 ( .A(n3), .B(n50), .Z(n48) );
  XNOR U45 ( .A(p_input[7]), .B(n49), .Z(n50) );
  XOR U46 ( .A(n51), .B(n52), .Z(n49) );
  AND U47 ( .A(n7), .B(n53), .Z(n52) );
  XNOR U48 ( .A(p_input[23]), .B(n51), .Z(n53) );
  XOR U49 ( .A(n54), .B(n55), .Z(n51) );
  AND U50 ( .A(n11), .B(n56), .Z(n55) );
  XNOR U51 ( .A(p_input[39]), .B(n54), .Z(n56) );
  XOR U52 ( .A(n57), .B(n58), .Z(n54) );
  AND U53 ( .A(n15), .B(n59), .Z(n58) );
  XNOR U54 ( .A(p_input[55]), .B(n57), .Z(n59) );
  XOR U55 ( .A(n60), .B(n61), .Z(n57) );
  AND U56 ( .A(n19), .B(n62), .Z(n61) );
  XNOR U57 ( .A(p_input[71]), .B(n60), .Z(n62) );
  XNOR U58 ( .A(n63), .B(n64), .Z(n60) );
  AND U59 ( .A(n23), .B(n65), .Z(n64) );
  XOR U60 ( .A(p_input[87]), .B(n63), .Z(n65) );
  XOR U61 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n66), .Z(n63) );
  AND U62 ( .A(n26), .B(n67), .Z(n66) );
  XOR U63 ( .A(p_input[103]), .B(\knn_comb_/min_val_out[0][7] ), .Z(n67) );
  XNOR U64 ( .A(n68), .B(n69), .Z(o[6]) );
  AND U65 ( .A(n3), .B(n70), .Z(n68) );
  XNOR U66 ( .A(p_input[6]), .B(n69), .Z(n70) );
  XOR U67 ( .A(n71), .B(n72), .Z(n69) );
  AND U68 ( .A(n7), .B(n73), .Z(n72) );
  XNOR U69 ( .A(p_input[22]), .B(n71), .Z(n73) );
  XOR U70 ( .A(n74), .B(n75), .Z(n71) );
  AND U71 ( .A(n11), .B(n76), .Z(n75) );
  XNOR U72 ( .A(p_input[38]), .B(n74), .Z(n76) );
  XOR U73 ( .A(n77), .B(n78), .Z(n74) );
  AND U74 ( .A(n15), .B(n79), .Z(n78) );
  XNOR U75 ( .A(p_input[54]), .B(n77), .Z(n79) );
  XOR U76 ( .A(n80), .B(n81), .Z(n77) );
  AND U77 ( .A(n19), .B(n82), .Z(n81) );
  XNOR U78 ( .A(p_input[70]), .B(n80), .Z(n82) );
  XNOR U79 ( .A(n83), .B(n84), .Z(n80) );
  AND U80 ( .A(n23), .B(n85), .Z(n84) );
  XOR U81 ( .A(p_input[86]), .B(n83), .Z(n85) );
  XOR U82 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n86), .Z(n83) );
  AND U83 ( .A(n26), .B(n87), .Z(n86) );
  XOR U84 ( .A(p_input[102]), .B(\knn_comb_/min_val_out[0][6] ), .Z(n87) );
  XNOR U85 ( .A(n88), .B(n89), .Z(o[5]) );
  AND U86 ( .A(n3), .B(n90), .Z(n88) );
  XNOR U87 ( .A(p_input[5]), .B(n89), .Z(n90) );
  XOR U88 ( .A(n91), .B(n92), .Z(n89) );
  AND U89 ( .A(n7), .B(n93), .Z(n92) );
  XNOR U90 ( .A(p_input[21]), .B(n91), .Z(n93) );
  XOR U91 ( .A(n94), .B(n95), .Z(n91) );
  AND U92 ( .A(n11), .B(n96), .Z(n95) );
  XNOR U93 ( .A(p_input[37]), .B(n94), .Z(n96) );
  XOR U94 ( .A(n97), .B(n98), .Z(n94) );
  AND U95 ( .A(n15), .B(n99), .Z(n98) );
  XNOR U96 ( .A(p_input[53]), .B(n97), .Z(n99) );
  XOR U97 ( .A(n100), .B(n101), .Z(n97) );
  AND U98 ( .A(n19), .B(n102), .Z(n101) );
  XNOR U99 ( .A(p_input[69]), .B(n100), .Z(n102) );
  XNOR U100 ( .A(n103), .B(n104), .Z(n100) );
  AND U101 ( .A(n23), .B(n105), .Z(n104) );
  XOR U102 ( .A(p_input[85]), .B(n103), .Z(n105) );
  XOR U103 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n106), .Z(n103) );
  AND U104 ( .A(n26), .B(n107), .Z(n106) );
  XOR U105 ( .A(p_input[101]), .B(\knn_comb_/min_val_out[0][5] ), .Z(n107) );
  XNOR U106 ( .A(n108), .B(n109), .Z(o[4]) );
  AND U107 ( .A(n3), .B(n110), .Z(n108) );
  XNOR U108 ( .A(p_input[4]), .B(n109), .Z(n110) );
  XOR U109 ( .A(n111), .B(n112), .Z(n109) );
  AND U110 ( .A(n7), .B(n113), .Z(n112) );
  XNOR U111 ( .A(p_input[20]), .B(n111), .Z(n113) );
  XOR U112 ( .A(n114), .B(n115), .Z(n111) );
  AND U113 ( .A(n11), .B(n116), .Z(n115) );
  XNOR U114 ( .A(p_input[36]), .B(n114), .Z(n116) );
  XOR U115 ( .A(n117), .B(n118), .Z(n114) );
  AND U116 ( .A(n15), .B(n119), .Z(n118) );
  XNOR U117 ( .A(p_input[52]), .B(n117), .Z(n119) );
  XOR U118 ( .A(n120), .B(n121), .Z(n117) );
  AND U119 ( .A(n19), .B(n122), .Z(n121) );
  XNOR U120 ( .A(p_input[68]), .B(n120), .Z(n122) );
  XNOR U121 ( .A(n123), .B(n124), .Z(n120) );
  AND U122 ( .A(n23), .B(n125), .Z(n124) );
  XOR U123 ( .A(p_input[84]), .B(n123), .Z(n125) );
  XOR U124 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n126), .Z(n123) );
  AND U125 ( .A(n26), .B(n127), .Z(n126) );
  XOR U126 ( .A(p_input[100]), .B(\knn_comb_/min_val_out[0][4] ), .Z(n127) );
  XNOR U127 ( .A(n128), .B(n129), .Z(o[3]) );
  AND U128 ( .A(n3), .B(n130), .Z(n128) );
  XNOR U129 ( .A(p_input[3]), .B(n129), .Z(n130) );
  XOR U130 ( .A(n131), .B(n132), .Z(n129) );
  AND U131 ( .A(n7), .B(n133), .Z(n132) );
  XNOR U132 ( .A(p_input[19]), .B(n131), .Z(n133) );
  XOR U133 ( .A(n134), .B(n135), .Z(n131) );
  AND U134 ( .A(n11), .B(n136), .Z(n135) );
  XNOR U135 ( .A(p_input[35]), .B(n134), .Z(n136) );
  XOR U136 ( .A(n137), .B(n138), .Z(n134) );
  AND U137 ( .A(n15), .B(n139), .Z(n138) );
  XNOR U138 ( .A(p_input[51]), .B(n137), .Z(n139) );
  XOR U139 ( .A(n140), .B(n141), .Z(n137) );
  AND U140 ( .A(n19), .B(n142), .Z(n141) );
  XNOR U141 ( .A(p_input[67]), .B(n140), .Z(n142) );
  XNOR U142 ( .A(n143), .B(n144), .Z(n140) );
  AND U143 ( .A(n23), .B(n145), .Z(n144) );
  XOR U144 ( .A(p_input[83]), .B(n143), .Z(n145) );
  XOR U145 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n146), .Z(n143) );
  AND U146 ( .A(n26), .B(n147), .Z(n146) );
  XOR U147 ( .A(p_input[99]), .B(\knn_comb_/min_val_out[0][3] ), .Z(n147) );
  XNOR U148 ( .A(n148), .B(n149), .Z(o[2]) );
  AND U149 ( .A(n3), .B(n150), .Z(n148) );
  XNOR U150 ( .A(p_input[2]), .B(n149), .Z(n150) );
  XOR U151 ( .A(n151), .B(n152), .Z(n149) );
  AND U152 ( .A(n7), .B(n153), .Z(n152) );
  XNOR U153 ( .A(p_input[18]), .B(n151), .Z(n153) );
  XOR U154 ( .A(n154), .B(n155), .Z(n151) );
  AND U155 ( .A(n11), .B(n156), .Z(n155) );
  XNOR U156 ( .A(p_input[34]), .B(n154), .Z(n156) );
  XOR U157 ( .A(n157), .B(n158), .Z(n154) );
  AND U158 ( .A(n15), .B(n159), .Z(n158) );
  XNOR U159 ( .A(p_input[50]), .B(n157), .Z(n159) );
  XOR U160 ( .A(n160), .B(n161), .Z(n157) );
  AND U161 ( .A(n19), .B(n162), .Z(n161) );
  XNOR U162 ( .A(p_input[66]), .B(n160), .Z(n162) );
  XNOR U163 ( .A(n163), .B(n164), .Z(n160) );
  AND U164 ( .A(n23), .B(n165), .Z(n164) );
  XOR U165 ( .A(p_input[82]), .B(n163), .Z(n165) );
  XOR U166 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n166), .Z(n163) );
  AND U167 ( .A(n26), .B(n167), .Z(n166) );
  XOR U168 ( .A(p_input[98]), .B(\knn_comb_/min_val_out[0][2] ), .Z(n167) );
  XNOR U169 ( .A(n168), .B(n169), .Z(o[1]) );
  AND U170 ( .A(n3), .B(n170), .Z(n168) );
  XNOR U171 ( .A(p_input[1]), .B(n169), .Z(n170) );
  XOR U172 ( .A(n171), .B(n172), .Z(n169) );
  AND U173 ( .A(n7), .B(n173), .Z(n172) );
  XNOR U174 ( .A(p_input[17]), .B(n171), .Z(n173) );
  XOR U175 ( .A(n174), .B(n175), .Z(n171) );
  AND U176 ( .A(n11), .B(n176), .Z(n175) );
  XNOR U177 ( .A(p_input[33]), .B(n174), .Z(n176) );
  XOR U178 ( .A(n177), .B(n178), .Z(n174) );
  AND U179 ( .A(n15), .B(n179), .Z(n178) );
  XNOR U180 ( .A(p_input[49]), .B(n177), .Z(n179) );
  XOR U181 ( .A(n180), .B(n181), .Z(n177) );
  AND U182 ( .A(n19), .B(n182), .Z(n181) );
  XNOR U183 ( .A(p_input[65]), .B(n180), .Z(n182) );
  XNOR U184 ( .A(n183), .B(n184), .Z(n180) );
  AND U185 ( .A(n23), .B(n185), .Z(n184) );
  XOR U186 ( .A(p_input[81]), .B(n183), .Z(n185) );
  XOR U187 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n186), .Z(n183) );
  AND U188 ( .A(n26), .B(n187), .Z(n186) );
  XOR U189 ( .A(p_input[97]), .B(\knn_comb_/min_val_out[0][1] ), .Z(n187) );
  XNOR U190 ( .A(n188), .B(n189), .Z(o[15]) );
  AND U191 ( .A(n3), .B(n190), .Z(n188) );
  XNOR U192 ( .A(p_input[15]), .B(n189), .Z(n190) );
  XOR U193 ( .A(n191), .B(n192), .Z(n189) );
  AND U194 ( .A(n7), .B(n193), .Z(n192) );
  XNOR U195 ( .A(p_input[31]), .B(n191), .Z(n193) );
  XOR U196 ( .A(n194), .B(n195), .Z(n191) );
  AND U197 ( .A(n11), .B(n196), .Z(n195) );
  XNOR U198 ( .A(p_input[47]), .B(n194), .Z(n196) );
  XOR U199 ( .A(n197), .B(n198), .Z(n194) );
  AND U200 ( .A(n15), .B(n199), .Z(n198) );
  XNOR U201 ( .A(p_input[63]), .B(n197), .Z(n199) );
  XOR U202 ( .A(n200), .B(n201), .Z(n197) );
  AND U203 ( .A(n19), .B(n202), .Z(n201) );
  XNOR U204 ( .A(p_input[79]), .B(n200), .Z(n202) );
  XNOR U205 ( .A(n203), .B(n204), .Z(n200) );
  AND U206 ( .A(n23), .B(n205), .Z(n204) );
  XOR U207 ( .A(p_input[95]), .B(n203), .Z(n205) );
  XOR U208 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n206), .Z(n203) );
  AND U209 ( .A(n26), .B(n207), .Z(n206) );
  XOR U210 ( .A(p_input[111]), .B(\knn_comb_/min_val_out[0][15] ), .Z(n207) );
  XNOR U211 ( .A(n208), .B(n209), .Z(o[14]) );
  AND U212 ( .A(n3), .B(n210), .Z(n208) );
  XNOR U213 ( .A(p_input[14]), .B(n209), .Z(n210) );
  XOR U214 ( .A(n211), .B(n212), .Z(n209) );
  AND U215 ( .A(n7), .B(n213), .Z(n212) );
  XNOR U216 ( .A(p_input[30]), .B(n211), .Z(n213) );
  XOR U217 ( .A(n214), .B(n215), .Z(n211) );
  AND U218 ( .A(n11), .B(n216), .Z(n215) );
  XNOR U219 ( .A(p_input[46]), .B(n214), .Z(n216) );
  XOR U220 ( .A(n217), .B(n218), .Z(n214) );
  AND U221 ( .A(n15), .B(n219), .Z(n218) );
  XNOR U222 ( .A(p_input[62]), .B(n217), .Z(n219) );
  XOR U223 ( .A(n220), .B(n221), .Z(n217) );
  AND U224 ( .A(n19), .B(n222), .Z(n221) );
  XNOR U225 ( .A(p_input[78]), .B(n220), .Z(n222) );
  XNOR U226 ( .A(n223), .B(n224), .Z(n220) );
  AND U227 ( .A(n23), .B(n225), .Z(n224) );
  XOR U228 ( .A(p_input[94]), .B(n223), .Z(n225) );
  XOR U229 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n226), .Z(n223) );
  AND U230 ( .A(n26), .B(n227), .Z(n226) );
  XOR U231 ( .A(p_input[110]), .B(\knn_comb_/min_val_out[0][14] ), .Z(n227) );
  XNOR U232 ( .A(n228), .B(n229), .Z(o[13]) );
  AND U233 ( .A(n3), .B(n230), .Z(n228) );
  XNOR U234 ( .A(p_input[13]), .B(n229), .Z(n230) );
  XOR U235 ( .A(n231), .B(n232), .Z(n229) );
  AND U236 ( .A(n7), .B(n233), .Z(n232) );
  XNOR U237 ( .A(p_input[29]), .B(n231), .Z(n233) );
  XOR U238 ( .A(n234), .B(n235), .Z(n231) );
  AND U239 ( .A(n11), .B(n236), .Z(n235) );
  XNOR U240 ( .A(p_input[45]), .B(n234), .Z(n236) );
  XOR U241 ( .A(n237), .B(n238), .Z(n234) );
  AND U242 ( .A(n15), .B(n239), .Z(n238) );
  XNOR U243 ( .A(p_input[61]), .B(n237), .Z(n239) );
  XOR U244 ( .A(n240), .B(n241), .Z(n237) );
  AND U245 ( .A(n19), .B(n242), .Z(n241) );
  XNOR U246 ( .A(p_input[77]), .B(n240), .Z(n242) );
  XNOR U247 ( .A(n243), .B(n244), .Z(n240) );
  AND U248 ( .A(n23), .B(n245), .Z(n244) );
  XOR U249 ( .A(p_input[93]), .B(n243), .Z(n245) );
  XOR U250 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n246), .Z(n243) );
  AND U251 ( .A(n26), .B(n247), .Z(n246) );
  XOR U252 ( .A(p_input[109]), .B(\knn_comb_/min_val_out[0][13] ), .Z(n247) );
  XNOR U253 ( .A(n248), .B(n249), .Z(o[12]) );
  AND U254 ( .A(n3), .B(n250), .Z(n248) );
  XNOR U255 ( .A(p_input[12]), .B(n249), .Z(n250) );
  XOR U256 ( .A(n251), .B(n252), .Z(n249) );
  AND U257 ( .A(n7), .B(n253), .Z(n252) );
  XNOR U258 ( .A(p_input[28]), .B(n251), .Z(n253) );
  XOR U259 ( .A(n254), .B(n255), .Z(n251) );
  AND U260 ( .A(n11), .B(n256), .Z(n255) );
  XNOR U261 ( .A(p_input[44]), .B(n254), .Z(n256) );
  XOR U262 ( .A(n257), .B(n258), .Z(n254) );
  AND U263 ( .A(n15), .B(n259), .Z(n258) );
  XNOR U264 ( .A(p_input[60]), .B(n257), .Z(n259) );
  XOR U265 ( .A(n260), .B(n261), .Z(n257) );
  AND U266 ( .A(n19), .B(n262), .Z(n261) );
  XNOR U267 ( .A(p_input[76]), .B(n260), .Z(n262) );
  XNOR U268 ( .A(n263), .B(n264), .Z(n260) );
  AND U269 ( .A(n23), .B(n265), .Z(n264) );
  XOR U270 ( .A(p_input[92]), .B(n263), .Z(n265) );
  XOR U271 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n266), .Z(n263) );
  AND U272 ( .A(n26), .B(n267), .Z(n266) );
  XOR U273 ( .A(p_input[108]), .B(\knn_comb_/min_val_out[0][12] ), .Z(n267) );
  XNOR U274 ( .A(n268), .B(n269), .Z(o[11]) );
  AND U275 ( .A(n3), .B(n270), .Z(n268) );
  XNOR U276 ( .A(p_input[11]), .B(n269), .Z(n270) );
  XOR U277 ( .A(n271), .B(n272), .Z(n269) );
  AND U278 ( .A(n7), .B(n273), .Z(n272) );
  XNOR U279 ( .A(p_input[27]), .B(n271), .Z(n273) );
  XOR U280 ( .A(n274), .B(n275), .Z(n271) );
  AND U281 ( .A(n11), .B(n276), .Z(n275) );
  XNOR U282 ( .A(p_input[43]), .B(n274), .Z(n276) );
  XOR U283 ( .A(n277), .B(n278), .Z(n274) );
  AND U284 ( .A(n15), .B(n279), .Z(n278) );
  XNOR U285 ( .A(p_input[59]), .B(n277), .Z(n279) );
  XOR U286 ( .A(n280), .B(n281), .Z(n277) );
  AND U287 ( .A(n19), .B(n282), .Z(n281) );
  XNOR U288 ( .A(p_input[75]), .B(n280), .Z(n282) );
  XNOR U289 ( .A(n283), .B(n284), .Z(n280) );
  AND U290 ( .A(n23), .B(n285), .Z(n284) );
  XOR U291 ( .A(p_input[91]), .B(n283), .Z(n285) );
  XOR U292 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n286), .Z(n283) );
  AND U293 ( .A(n26), .B(n287), .Z(n286) );
  XOR U294 ( .A(p_input[107]), .B(\knn_comb_/min_val_out[0][11] ), .Z(n287) );
  XNOR U295 ( .A(n288), .B(n289), .Z(o[10]) );
  AND U296 ( .A(n3), .B(n290), .Z(n288) );
  XNOR U297 ( .A(p_input[10]), .B(n289), .Z(n290) );
  XOR U298 ( .A(n291), .B(n292), .Z(n289) );
  AND U299 ( .A(n7), .B(n293), .Z(n292) );
  XNOR U300 ( .A(p_input[26]), .B(n291), .Z(n293) );
  XOR U301 ( .A(n294), .B(n295), .Z(n291) );
  AND U302 ( .A(n11), .B(n296), .Z(n295) );
  XNOR U303 ( .A(p_input[42]), .B(n294), .Z(n296) );
  XOR U304 ( .A(n297), .B(n298), .Z(n294) );
  AND U305 ( .A(n15), .B(n299), .Z(n298) );
  XNOR U306 ( .A(p_input[58]), .B(n297), .Z(n299) );
  XOR U307 ( .A(n300), .B(n301), .Z(n297) );
  AND U308 ( .A(n19), .B(n302), .Z(n301) );
  XNOR U309 ( .A(p_input[74]), .B(n300), .Z(n302) );
  XNOR U310 ( .A(n303), .B(n304), .Z(n300) );
  AND U311 ( .A(n23), .B(n305), .Z(n304) );
  XOR U312 ( .A(p_input[90]), .B(n303), .Z(n305) );
  XOR U313 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n306), .Z(n303) );
  AND U314 ( .A(n26), .B(n307), .Z(n306) );
  XOR U315 ( .A(p_input[106]), .B(\knn_comb_/min_val_out[0][10] ), .Z(n307) );
  XNOR U316 ( .A(n308), .B(n309), .Z(o[0]) );
  AND U317 ( .A(n3), .B(n310), .Z(n308) );
  XNOR U318 ( .A(p_input[0]), .B(n309), .Z(n310) );
  XOR U319 ( .A(n311), .B(n312), .Z(n309) );
  AND U320 ( .A(n7), .B(n313), .Z(n312) );
  XNOR U321 ( .A(p_input[16]), .B(n311), .Z(n313) );
  XOR U322 ( .A(n314), .B(n315), .Z(n311) );
  AND U323 ( .A(n11), .B(n316), .Z(n315) );
  XNOR U324 ( .A(p_input[32]), .B(n314), .Z(n316) );
  XOR U325 ( .A(n317), .B(n318), .Z(n314) );
  AND U326 ( .A(n15), .B(n319), .Z(n318) );
  XNOR U327 ( .A(p_input[48]), .B(n317), .Z(n319) );
  XOR U328 ( .A(n320), .B(n321), .Z(n317) );
  AND U329 ( .A(n19), .B(n322), .Z(n321) );
  XNOR U330 ( .A(p_input[64]), .B(n320), .Z(n322) );
  XNOR U331 ( .A(n323), .B(n324), .Z(n320) );
  AND U332 ( .A(n23), .B(n325), .Z(n324) );
  XOR U333 ( .A(p_input[80]), .B(n323), .Z(n325) );
  XOR U334 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n326), .Z(n323) );
  AND U335 ( .A(n26), .B(n327), .Z(n326) );
  XOR U336 ( .A(p_input[96]), .B(\knn_comb_/min_val_out[0][0] ), .Z(n327) );
  XNOR U337 ( .A(n328), .B(n329), .Z(n3) );
  NOR U338 ( .A(n330), .B(n331), .Z(n329) );
  XOR U339 ( .A(n332), .B(n328), .Z(n331) );
  AND U340 ( .A(n333), .B(n334), .Z(n332) );
  NOR U341 ( .A(n335), .B(n328), .Z(n330) );
  AND U342 ( .A(n336), .B(n337), .Z(n335) );
  XOR U343 ( .A(n338), .B(n339), .Z(n328) );
  AND U344 ( .A(n340), .B(n341), .Z(n339) );
  XNOR U345 ( .A(n338), .B(n336), .Z(n341) );
  XNOR U346 ( .A(n342), .B(n343), .Z(n336) );
  XOR U347 ( .A(n344), .B(n337), .Z(n343) );
  AND U348 ( .A(n345), .B(n346), .Z(n337) );
  AND U349 ( .A(n347), .B(n348), .Z(n344) );
  XOR U350 ( .A(n349), .B(n342), .Z(n347) );
  XOR U351 ( .A(n350), .B(n338), .Z(n340) );
  XNOR U352 ( .A(n351), .B(n352), .Z(n350) );
  AND U353 ( .A(n7), .B(n353), .Z(n352) );
  XOR U354 ( .A(n354), .B(n351), .Z(n353) );
  XOR U355 ( .A(n355), .B(n356), .Z(n338) );
  AND U356 ( .A(n357), .B(n358), .Z(n356) );
  XNOR U357 ( .A(n355), .B(n345), .Z(n358) );
  XOR U358 ( .A(n359), .B(n348), .Z(n345) );
  XNOR U359 ( .A(n360), .B(n342), .Z(n348) );
  XOR U360 ( .A(n361), .B(n362), .Z(n342) );
  AND U361 ( .A(n363), .B(n364), .Z(n362) );
  XOR U362 ( .A(n365), .B(n361), .Z(n363) );
  XNOR U363 ( .A(n366), .B(n367), .Z(n360) );
  AND U364 ( .A(n368), .B(n369), .Z(n367) );
  XOR U365 ( .A(n366), .B(n370), .Z(n368) );
  XNOR U366 ( .A(n349), .B(n346), .Z(n359) );
  AND U367 ( .A(n371), .B(n372), .Z(n346) );
  XOR U368 ( .A(n373), .B(n374), .Z(n349) );
  AND U369 ( .A(n375), .B(n376), .Z(n374) );
  XOR U370 ( .A(n373), .B(n377), .Z(n375) );
  XOR U371 ( .A(n378), .B(n355), .Z(n357) );
  XNOR U372 ( .A(n379), .B(n380), .Z(n378) );
  AND U373 ( .A(n7), .B(n381), .Z(n380) );
  XNOR U374 ( .A(n382), .B(n379), .Z(n381) );
  XOR U375 ( .A(n383), .B(n384), .Z(n355) );
  AND U376 ( .A(n385), .B(n386), .Z(n384) );
  XNOR U377 ( .A(n383), .B(n371), .Z(n386) );
  XOR U378 ( .A(n387), .B(n364), .Z(n371) );
  XNOR U379 ( .A(n388), .B(n370), .Z(n364) );
  XNOR U380 ( .A(n389), .B(n390), .Z(n370) );
  NOR U381 ( .A(n391), .B(n392), .Z(n390) );
  XOR U382 ( .A(n389), .B(n393), .Z(n391) );
  XNOR U383 ( .A(n369), .B(n361), .Z(n388) );
  XOR U384 ( .A(n394), .B(n395), .Z(n361) );
  AND U385 ( .A(n396), .B(n397), .Z(n395) );
  XNOR U386 ( .A(n394), .B(n398), .Z(n396) );
  XNOR U387 ( .A(n399), .B(n366), .Z(n369) );
  XOR U388 ( .A(n400), .B(n401), .Z(n366) );
  AND U389 ( .A(n402), .B(n403), .Z(n401) );
  XOR U390 ( .A(n400), .B(n404), .Z(n402) );
  XNOR U391 ( .A(n405), .B(n406), .Z(n399) );
  NOR U392 ( .A(n407), .B(n408), .Z(n406) );
  XOR U393 ( .A(n405), .B(n409), .Z(n407) );
  XNOR U394 ( .A(n365), .B(n372), .Z(n387) );
  NOR U395 ( .A(n410), .B(n411), .Z(n372) );
  XOR U396 ( .A(n377), .B(n376), .Z(n365) );
  XNOR U397 ( .A(n412), .B(n373), .Z(n376) );
  XOR U398 ( .A(n413), .B(n414), .Z(n373) );
  AND U399 ( .A(n415), .B(n416), .Z(n414) );
  XNOR U400 ( .A(n417), .B(n418), .Z(n415) );
  XNOR U401 ( .A(n419), .B(n420), .Z(n412) );
  NOR U402 ( .A(n421), .B(n422), .Z(n420) );
  XNOR U403 ( .A(n419), .B(n423), .Z(n421) );
  XOR U404 ( .A(n424), .B(n425), .Z(n377) );
  NOR U405 ( .A(n426), .B(n427), .Z(n425) );
  XNOR U406 ( .A(n424), .B(n428), .Z(n426) );
  XNOR U407 ( .A(n429), .B(n430), .Z(n385) );
  XOR U408 ( .A(n383), .B(n431), .Z(n430) );
  AND U409 ( .A(n7), .B(n432), .Z(n431) );
  XOR U410 ( .A(n433), .B(n429), .Z(n432) );
  AND U411 ( .A(n434), .B(n410), .Z(n383) );
  XOR U412 ( .A(n435), .B(n411), .Z(n410) );
  XNOR U413 ( .A(p_input[0]), .B(p_input[128]), .Z(n411) );
  XOR U414 ( .A(n398), .B(n397), .Z(n435) );
  XNOR U415 ( .A(n436), .B(n404), .Z(n397) );
  XNOR U416 ( .A(n393), .B(n392), .Z(n404) );
  XNOR U417 ( .A(n437), .B(n389), .Z(n392) );
  XNOR U418 ( .A(p_input[10]), .B(p_input[138]), .Z(n389) );
  XOR U419 ( .A(p_input[11]), .B(n438), .Z(n437) );
  XOR U420 ( .A(p_input[12]), .B(p_input[140]), .Z(n393) );
  XOR U421 ( .A(n403), .B(n439), .Z(n436) );
  IV U422 ( .A(n394), .Z(n439) );
  XOR U423 ( .A(p_input[129]), .B(p_input[1]), .Z(n394) );
  XOR U424 ( .A(n440), .B(n409), .Z(n403) );
  XNOR U425 ( .A(p_input[143]), .B(p_input[15]), .Z(n409) );
  XOR U426 ( .A(n400), .B(n408), .Z(n440) );
  XOR U427 ( .A(n441), .B(n405), .Z(n408) );
  XOR U428 ( .A(p_input[13]), .B(p_input[141]), .Z(n405) );
  XNOR U429 ( .A(p_input[142]), .B(p_input[14]), .Z(n441) );
  XOR U430 ( .A(p_input[137]), .B(p_input[9]), .Z(n400) );
  XNOR U431 ( .A(n418), .B(n416), .Z(n398) );
  XNOR U432 ( .A(n442), .B(n423), .Z(n416) );
  XOR U433 ( .A(p_input[136]), .B(p_input[8]), .Z(n423) );
  XOR U434 ( .A(n413), .B(n422), .Z(n442) );
  XOR U435 ( .A(n443), .B(n419), .Z(n422) );
  XOR U436 ( .A(p_input[134]), .B(p_input[6]), .Z(n419) );
  XNOR U437 ( .A(p_input[135]), .B(p_input[7]), .Z(n443) );
  IV U438 ( .A(n417), .Z(n413) );
  XNOR U439 ( .A(p_input[130]), .B(p_input[2]), .Z(n417) );
  XNOR U440 ( .A(n428), .B(n427), .Z(n418) );
  XOR U441 ( .A(n444), .B(n424), .Z(n427) );
  XOR U442 ( .A(p_input[131]), .B(p_input[3]), .Z(n424) );
  XNOR U443 ( .A(p_input[132]), .B(p_input[4]), .Z(n444) );
  XOR U444 ( .A(p_input[133]), .B(p_input[5]), .Z(n428) );
  XNOR U445 ( .A(n445), .B(n446), .Z(n434) );
  AND U446 ( .A(n7), .B(n447), .Z(n446) );
  XNOR U447 ( .A(n448), .B(n449), .Z(n447) );
  XNOR U448 ( .A(n450), .B(n451), .Z(n7) );
  MUX U449 ( .IN0(n333), .IN1(n334), .SEL(n450), .F(n451) );
  AND U450 ( .A(n452), .B(n453), .Z(n334) );
  AND U451 ( .A(n454), .B(n455), .Z(n333) );
  XOR U452 ( .A(n456), .B(n457), .Z(n450) );
  AND U453 ( .A(n458), .B(n459), .Z(n457) );
  XNOR U454 ( .A(n456), .B(n454), .Z(n459) );
  IV U455 ( .A(n354), .Z(n454) );
  XOR U456 ( .A(n460), .B(n461), .Z(n354) );
  XOR U457 ( .A(n462), .B(n455), .Z(n461) );
  AND U458 ( .A(n382), .B(n463), .Z(n455) );
  AND U459 ( .A(n464), .B(n465), .Z(n462) );
  XOR U460 ( .A(n466), .B(n460), .Z(n464) );
  XNOR U461 ( .A(n351), .B(n456), .Z(n458) );
  XOR U462 ( .A(n467), .B(n468), .Z(n351) );
  AND U463 ( .A(n11), .B(n469), .Z(n468) );
  XOR U464 ( .A(n470), .B(n467), .Z(n469) );
  XOR U465 ( .A(n471), .B(n472), .Z(n456) );
  AND U466 ( .A(n473), .B(n474), .Z(n472) );
  XNOR U467 ( .A(n471), .B(n382), .Z(n474) );
  XOR U468 ( .A(n475), .B(n465), .Z(n382) );
  XNOR U469 ( .A(n476), .B(n460), .Z(n465) );
  XOR U470 ( .A(n477), .B(n478), .Z(n460) );
  AND U471 ( .A(n479), .B(n480), .Z(n478) );
  XOR U472 ( .A(n481), .B(n477), .Z(n479) );
  XNOR U473 ( .A(n482), .B(n483), .Z(n476) );
  AND U474 ( .A(n484), .B(n485), .Z(n483) );
  XOR U475 ( .A(n482), .B(n486), .Z(n484) );
  XNOR U476 ( .A(n466), .B(n463), .Z(n475) );
  AND U477 ( .A(n487), .B(n488), .Z(n463) );
  XOR U478 ( .A(n489), .B(n490), .Z(n466) );
  AND U479 ( .A(n491), .B(n492), .Z(n490) );
  XOR U480 ( .A(n489), .B(n493), .Z(n491) );
  XNOR U481 ( .A(n379), .B(n471), .Z(n473) );
  XOR U482 ( .A(n494), .B(n495), .Z(n379) );
  AND U483 ( .A(n11), .B(n496), .Z(n495) );
  XNOR U484 ( .A(n497), .B(n494), .Z(n496) );
  XOR U485 ( .A(n498), .B(n499), .Z(n471) );
  AND U486 ( .A(n500), .B(n501), .Z(n499) );
  XNOR U487 ( .A(n498), .B(n487), .Z(n501) );
  IV U488 ( .A(n433), .Z(n487) );
  XNOR U489 ( .A(n502), .B(n480), .Z(n433) );
  XNOR U490 ( .A(n503), .B(n486), .Z(n480) );
  XOR U491 ( .A(n504), .B(n505), .Z(n486) );
  NOR U492 ( .A(n506), .B(n507), .Z(n505) );
  XNOR U493 ( .A(n504), .B(n508), .Z(n506) );
  XNOR U494 ( .A(n485), .B(n477), .Z(n503) );
  XOR U495 ( .A(n509), .B(n510), .Z(n477) );
  AND U496 ( .A(n511), .B(n512), .Z(n510) );
  XNOR U497 ( .A(n509), .B(n513), .Z(n511) );
  XNOR U498 ( .A(n514), .B(n482), .Z(n485) );
  XOR U499 ( .A(n515), .B(n516), .Z(n482) );
  AND U500 ( .A(n517), .B(n518), .Z(n516) );
  XOR U501 ( .A(n515), .B(n519), .Z(n517) );
  XNOR U502 ( .A(n520), .B(n521), .Z(n514) );
  NOR U503 ( .A(n522), .B(n523), .Z(n521) );
  XOR U504 ( .A(n520), .B(n524), .Z(n522) );
  XNOR U505 ( .A(n481), .B(n488), .Z(n502) );
  NOR U506 ( .A(n448), .B(n525), .Z(n488) );
  XOR U507 ( .A(n493), .B(n492), .Z(n481) );
  XNOR U508 ( .A(n526), .B(n489), .Z(n492) );
  XOR U509 ( .A(n527), .B(n528), .Z(n489) );
  AND U510 ( .A(n529), .B(n530), .Z(n528) );
  XOR U511 ( .A(n527), .B(n531), .Z(n529) );
  XNOR U512 ( .A(n532), .B(n533), .Z(n526) );
  NOR U513 ( .A(n534), .B(n535), .Z(n533) );
  XNOR U514 ( .A(n532), .B(n536), .Z(n534) );
  XOR U515 ( .A(n537), .B(n538), .Z(n493) );
  NOR U516 ( .A(n539), .B(n540), .Z(n538) );
  XNOR U517 ( .A(n537), .B(n541), .Z(n539) );
  XNOR U518 ( .A(n429), .B(n498), .Z(n500) );
  XOR U519 ( .A(n542), .B(n543), .Z(n429) );
  AND U520 ( .A(n11), .B(n544), .Z(n543) );
  XOR U521 ( .A(n545), .B(n542), .Z(n544) );
  AND U522 ( .A(n449), .B(n448), .Z(n498) );
  XOR U523 ( .A(n546), .B(n525), .Z(n448) );
  XNOR U524 ( .A(p_input[128]), .B(p_input[16]), .Z(n525) );
  XOR U525 ( .A(n513), .B(n512), .Z(n546) );
  XNOR U526 ( .A(n547), .B(n519), .Z(n512) );
  XNOR U527 ( .A(n508), .B(n507), .Z(n519) );
  XOR U528 ( .A(n548), .B(n504), .Z(n507) );
  XNOR U529 ( .A(n549), .B(p_input[26]), .Z(n504) );
  XNOR U530 ( .A(p_input[139]), .B(p_input[27]), .Z(n548) );
  XOR U531 ( .A(p_input[140]), .B(p_input[28]), .Z(n508) );
  XNOR U532 ( .A(n518), .B(n509), .Z(n547) );
  XNOR U533 ( .A(n550), .B(p_input[17]), .Z(n509) );
  XOR U534 ( .A(n551), .B(n524), .Z(n518) );
  XNOR U535 ( .A(p_input[143]), .B(p_input[31]), .Z(n524) );
  XOR U536 ( .A(n515), .B(n523), .Z(n551) );
  XOR U537 ( .A(n552), .B(n520), .Z(n523) );
  XOR U538 ( .A(p_input[141]), .B(p_input[29]), .Z(n520) );
  XNOR U539 ( .A(p_input[142]), .B(p_input[30]), .Z(n552) );
  XOR U540 ( .A(p_input[137]), .B(p_input[25]), .Z(n515) );
  XNOR U541 ( .A(n531), .B(n530), .Z(n513) );
  XNOR U542 ( .A(n553), .B(n536), .Z(n530) );
  XOR U543 ( .A(p_input[136]), .B(p_input[24]), .Z(n536) );
  XOR U544 ( .A(n527), .B(n535), .Z(n553) );
  XOR U545 ( .A(n554), .B(n532), .Z(n535) );
  XOR U546 ( .A(p_input[134]), .B(p_input[22]), .Z(n532) );
  XNOR U547 ( .A(p_input[135]), .B(p_input[23]), .Z(n554) );
  XOR U548 ( .A(p_input[130]), .B(p_input[18]), .Z(n527) );
  XNOR U549 ( .A(n541), .B(n540), .Z(n531) );
  XOR U550 ( .A(n555), .B(n537), .Z(n540) );
  XOR U551 ( .A(p_input[131]), .B(p_input[19]), .Z(n537) );
  XNOR U552 ( .A(p_input[132]), .B(p_input[20]), .Z(n555) );
  XOR U553 ( .A(p_input[133]), .B(p_input[21]), .Z(n541) );
  IV U554 ( .A(n445), .Z(n449) );
  XNOR U555 ( .A(n556), .B(n557), .Z(n445) );
  AND U556 ( .A(n11), .B(n558), .Z(n557) );
  XNOR U557 ( .A(n559), .B(n556), .Z(n558) );
  XNOR U558 ( .A(n560), .B(n561), .Z(n11) );
  MUX U559 ( .IN0(n452), .IN1(n453), .SEL(n560), .F(n561) );
  AND U560 ( .A(n562), .B(n563), .Z(n453) );
  AND U561 ( .A(n564), .B(n565), .Z(n452) );
  XOR U562 ( .A(n566), .B(n567), .Z(n560) );
  AND U563 ( .A(n568), .B(n569), .Z(n567) );
  XNOR U564 ( .A(n566), .B(n564), .Z(n569) );
  IV U565 ( .A(n470), .Z(n564) );
  XOR U566 ( .A(n570), .B(n571), .Z(n470) );
  XOR U567 ( .A(n572), .B(n565), .Z(n571) );
  AND U568 ( .A(n497), .B(n573), .Z(n565) );
  AND U569 ( .A(n574), .B(n575), .Z(n572) );
  XOR U570 ( .A(n576), .B(n570), .Z(n574) );
  XNOR U571 ( .A(n467), .B(n566), .Z(n568) );
  XOR U572 ( .A(n577), .B(n578), .Z(n467) );
  AND U573 ( .A(n15), .B(n579), .Z(n578) );
  XOR U574 ( .A(n580), .B(n577), .Z(n579) );
  XOR U575 ( .A(n581), .B(n582), .Z(n566) );
  AND U576 ( .A(n583), .B(n584), .Z(n582) );
  XNOR U577 ( .A(n581), .B(n497), .Z(n584) );
  XOR U578 ( .A(n585), .B(n575), .Z(n497) );
  XNOR U579 ( .A(n586), .B(n570), .Z(n575) );
  XOR U580 ( .A(n587), .B(n588), .Z(n570) );
  AND U581 ( .A(n589), .B(n590), .Z(n588) );
  XOR U582 ( .A(n591), .B(n587), .Z(n589) );
  XNOR U583 ( .A(n592), .B(n593), .Z(n586) );
  AND U584 ( .A(n594), .B(n595), .Z(n593) );
  XOR U585 ( .A(n592), .B(n596), .Z(n594) );
  XNOR U586 ( .A(n576), .B(n573), .Z(n585) );
  AND U587 ( .A(n597), .B(n598), .Z(n573) );
  XOR U588 ( .A(n599), .B(n600), .Z(n576) );
  AND U589 ( .A(n601), .B(n602), .Z(n600) );
  XOR U590 ( .A(n599), .B(n603), .Z(n601) );
  XNOR U591 ( .A(n494), .B(n581), .Z(n583) );
  XOR U592 ( .A(n604), .B(n605), .Z(n494) );
  AND U593 ( .A(n15), .B(n606), .Z(n605) );
  XNOR U594 ( .A(n607), .B(n604), .Z(n606) );
  XOR U595 ( .A(n608), .B(n609), .Z(n581) );
  AND U596 ( .A(n610), .B(n611), .Z(n609) );
  XNOR U597 ( .A(n608), .B(n597), .Z(n611) );
  IV U598 ( .A(n545), .Z(n597) );
  XNOR U599 ( .A(n612), .B(n590), .Z(n545) );
  XNOR U600 ( .A(n613), .B(n596), .Z(n590) );
  XOR U601 ( .A(n614), .B(n615), .Z(n596) );
  NOR U602 ( .A(n616), .B(n617), .Z(n615) );
  XNOR U603 ( .A(n614), .B(n618), .Z(n616) );
  XNOR U604 ( .A(n595), .B(n587), .Z(n613) );
  XOR U605 ( .A(n619), .B(n620), .Z(n587) );
  AND U606 ( .A(n621), .B(n622), .Z(n620) );
  XNOR U607 ( .A(n619), .B(n623), .Z(n621) );
  XNOR U608 ( .A(n624), .B(n592), .Z(n595) );
  XOR U609 ( .A(n625), .B(n626), .Z(n592) );
  AND U610 ( .A(n627), .B(n628), .Z(n626) );
  XOR U611 ( .A(n625), .B(n629), .Z(n627) );
  XNOR U612 ( .A(n630), .B(n631), .Z(n624) );
  NOR U613 ( .A(n632), .B(n633), .Z(n631) );
  XOR U614 ( .A(n630), .B(n634), .Z(n632) );
  XNOR U615 ( .A(n591), .B(n598), .Z(n612) );
  NOR U616 ( .A(n559), .B(n635), .Z(n598) );
  XOR U617 ( .A(n603), .B(n602), .Z(n591) );
  XNOR U618 ( .A(n636), .B(n599), .Z(n602) );
  XOR U619 ( .A(n637), .B(n638), .Z(n599) );
  AND U620 ( .A(n639), .B(n640), .Z(n638) );
  XOR U621 ( .A(n637), .B(n641), .Z(n639) );
  XNOR U622 ( .A(n642), .B(n643), .Z(n636) );
  NOR U623 ( .A(n644), .B(n645), .Z(n643) );
  XNOR U624 ( .A(n642), .B(n646), .Z(n644) );
  XOR U625 ( .A(n647), .B(n648), .Z(n603) );
  NOR U626 ( .A(n649), .B(n650), .Z(n648) );
  XNOR U627 ( .A(n647), .B(n651), .Z(n649) );
  XNOR U628 ( .A(n542), .B(n608), .Z(n610) );
  XOR U629 ( .A(n652), .B(n653), .Z(n542) );
  AND U630 ( .A(n15), .B(n654), .Z(n653) );
  XOR U631 ( .A(n655), .B(n652), .Z(n654) );
  AND U632 ( .A(n556), .B(n559), .Z(n608) );
  XOR U633 ( .A(n656), .B(n635), .Z(n559) );
  XNOR U634 ( .A(p_input[128]), .B(p_input[32]), .Z(n635) );
  XOR U635 ( .A(n623), .B(n622), .Z(n656) );
  XNOR U636 ( .A(n657), .B(n629), .Z(n622) );
  XNOR U637 ( .A(n618), .B(n617), .Z(n629) );
  XOR U638 ( .A(n658), .B(n614), .Z(n617) );
  XNOR U639 ( .A(n549), .B(p_input[42]), .Z(n614) );
  XNOR U640 ( .A(p_input[139]), .B(p_input[43]), .Z(n658) );
  XOR U641 ( .A(p_input[140]), .B(p_input[44]), .Z(n618) );
  XNOR U642 ( .A(n628), .B(n619), .Z(n657) );
  XNOR U643 ( .A(n550), .B(p_input[33]), .Z(n619) );
  XOR U644 ( .A(n659), .B(n634), .Z(n628) );
  XNOR U645 ( .A(p_input[143]), .B(p_input[47]), .Z(n634) );
  XOR U646 ( .A(n625), .B(n633), .Z(n659) );
  XOR U647 ( .A(n660), .B(n630), .Z(n633) );
  XOR U648 ( .A(p_input[141]), .B(p_input[45]), .Z(n630) );
  XNOR U649 ( .A(p_input[142]), .B(p_input[46]), .Z(n660) );
  XOR U650 ( .A(p_input[137]), .B(p_input[41]), .Z(n625) );
  XNOR U651 ( .A(n641), .B(n640), .Z(n623) );
  XNOR U652 ( .A(n661), .B(n646), .Z(n640) );
  XOR U653 ( .A(p_input[136]), .B(p_input[40]), .Z(n646) );
  XOR U654 ( .A(n637), .B(n645), .Z(n661) );
  XOR U655 ( .A(n662), .B(n642), .Z(n645) );
  XOR U656 ( .A(p_input[134]), .B(p_input[38]), .Z(n642) );
  XNOR U657 ( .A(p_input[135]), .B(p_input[39]), .Z(n662) );
  XOR U658 ( .A(p_input[130]), .B(p_input[34]), .Z(n637) );
  XNOR U659 ( .A(n651), .B(n650), .Z(n641) );
  XOR U660 ( .A(n663), .B(n647), .Z(n650) );
  XOR U661 ( .A(p_input[131]), .B(p_input[35]), .Z(n647) );
  XNOR U662 ( .A(p_input[132]), .B(p_input[36]), .Z(n663) );
  XOR U663 ( .A(p_input[133]), .B(p_input[37]), .Z(n651) );
  XOR U664 ( .A(n664), .B(n665), .Z(n556) );
  AND U665 ( .A(n15), .B(n666), .Z(n665) );
  XNOR U666 ( .A(n667), .B(n664), .Z(n666) );
  XNOR U667 ( .A(n668), .B(n669), .Z(n15) );
  MUX U668 ( .IN0(n562), .IN1(n563), .SEL(n668), .F(n669) );
  AND U669 ( .A(n670), .B(n671), .Z(n563) );
  AND U670 ( .A(n672), .B(n673), .Z(n562) );
  XOR U671 ( .A(n674), .B(n675), .Z(n668) );
  AND U672 ( .A(n676), .B(n677), .Z(n675) );
  XNOR U673 ( .A(n674), .B(n672), .Z(n677) );
  IV U674 ( .A(n580), .Z(n672) );
  XOR U675 ( .A(n678), .B(n679), .Z(n580) );
  XOR U676 ( .A(n680), .B(n673), .Z(n679) );
  AND U677 ( .A(n607), .B(n681), .Z(n673) );
  AND U678 ( .A(n682), .B(n683), .Z(n680) );
  XOR U679 ( .A(n684), .B(n678), .Z(n682) );
  XNOR U680 ( .A(n577), .B(n674), .Z(n676) );
  XOR U681 ( .A(n685), .B(n686), .Z(n577) );
  AND U682 ( .A(n19), .B(n687), .Z(n686) );
  XOR U683 ( .A(n688), .B(n685), .Z(n687) );
  XOR U684 ( .A(n689), .B(n690), .Z(n674) );
  AND U685 ( .A(n691), .B(n692), .Z(n690) );
  XNOR U686 ( .A(n689), .B(n607), .Z(n692) );
  XOR U687 ( .A(n693), .B(n683), .Z(n607) );
  XNOR U688 ( .A(n694), .B(n678), .Z(n683) );
  XOR U689 ( .A(n695), .B(n696), .Z(n678) );
  AND U690 ( .A(n697), .B(n698), .Z(n696) );
  XOR U691 ( .A(n699), .B(n695), .Z(n697) );
  XNOR U692 ( .A(n700), .B(n701), .Z(n694) );
  AND U693 ( .A(n702), .B(n703), .Z(n701) );
  XOR U694 ( .A(n700), .B(n704), .Z(n702) );
  XNOR U695 ( .A(n684), .B(n681), .Z(n693) );
  AND U696 ( .A(n705), .B(n706), .Z(n681) );
  XOR U697 ( .A(n707), .B(n708), .Z(n684) );
  AND U698 ( .A(n709), .B(n710), .Z(n708) );
  XOR U699 ( .A(n707), .B(n711), .Z(n709) );
  XNOR U700 ( .A(n604), .B(n689), .Z(n691) );
  XOR U701 ( .A(n712), .B(n713), .Z(n604) );
  AND U702 ( .A(n19), .B(n714), .Z(n713) );
  XNOR U703 ( .A(n715), .B(n712), .Z(n714) );
  XOR U704 ( .A(n716), .B(n717), .Z(n689) );
  AND U705 ( .A(n718), .B(n719), .Z(n717) );
  XNOR U706 ( .A(n716), .B(n705), .Z(n719) );
  IV U707 ( .A(n655), .Z(n705) );
  XNOR U708 ( .A(n720), .B(n698), .Z(n655) );
  XNOR U709 ( .A(n721), .B(n704), .Z(n698) );
  XOR U710 ( .A(n722), .B(n723), .Z(n704) );
  NOR U711 ( .A(n724), .B(n725), .Z(n723) );
  XNOR U712 ( .A(n722), .B(n726), .Z(n724) );
  XNOR U713 ( .A(n703), .B(n695), .Z(n721) );
  XOR U714 ( .A(n727), .B(n728), .Z(n695) );
  AND U715 ( .A(n729), .B(n730), .Z(n728) );
  XNOR U716 ( .A(n727), .B(n731), .Z(n729) );
  XNOR U717 ( .A(n732), .B(n700), .Z(n703) );
  XOR U718 ( .A(n733), .B(n734), .Z(n700) );
  AND U719 ( .A(n735), .B(n736), .Z(n734) );
  XOR U720 ( .A(n733), .B(n737), .Z(n735) );
  XNOR U721 ( .A(n738), .B(n739), .Z(n732) );
  NOR U722 ( .A(n740), .B(n741), .Z(n739) );
  XOR U723 ( .A(n738), .B(n742), .Z(n740) );
  XNOR U724 ( .A(n699), .B(n706), .Z(n720) );
  NOR U725 ( .A(n667), .B(n743), .Z(n706) );
  XOR U726 ( .A(n711), .B(n710), .Z(n699) );
  XNOR U727 ( .A(n744), .B(n707), .Z(n710) );
  XOR U728 ( .A(n745), .B(n746), .Z(n707) );
  AND U729 ( .A(n747), .B(n748), .Z(n746) );
  XOR U730 ( .A(n745), .B(n749), .Z(n747) );
  XNOR U731 ( .A(n750), .B(n751), .Z(n744) );
  NOR U732 ( .A(n752), .B(n753), .Z(n751) );
  XNOR U733 ( .A(n750), .B(n754), .Z(n752) );
  XOR U734 ( .A(n755), .B(n756), .Z(n711) );
  NOR U735 ( .A(n757), .B(n758), .Z(n756) );
  XNOR U736 ( .A(n755), .B(n759), .Z(n757) );
  XNOR U737 ( .A(n652), .B(n716), .Z(n718) );
  XOR U738 ( .A(n760), .B(n761), .Z(n652) );
  AND U739 ( .A(n19), .B(n762), .Z(n761) );
  XOR U740 ( .A(n763), .B(n760), .Z(n762) );
  AND U741 ( .A(n664), .B(n667), .Z(n716) );
  XOR U742 ( .A(n764), .B(n743), .Z(n667) );
  XNOR U743 ( .A(p_input[128]), .B(p_input[48]), .Z(n743) );
  XOR U744 ( .A(n731), .B(n730), .Z(n764) );
  XNOR U745 ( .A(n765), .B(n737), .Z(n730) );
  XNOR U746 ( .A(n726), .B(n725), .Z(n737) );
  XOR U747 ( .A(n766), .B(n722), .Z(n725) );
  XNOR U748 ( .A(n549), .B(p_input[58]), .Z(n722) );
  XNOR U749 ( .A(p_input[139]), .B(p_input[59]), .Z(n766) );
  XOR U750 ( .A(p_input[140]), .B(p_input[60]), .Z(n726) );
  XNOR U751 ( .A(n736), .B(n727), .Z(n765) );
  XNOR U752 ( .A(n550), .B(p_input[49]), .Z(n727) );
  XOR U753 ( .A(n767), .B(n742), .Z(n736) );
  XNOR U754 ( .A(p_input[143]), .B(p_input[63]), .Z(n742) );
  XOR U755 ( .A(n733), .B(n741), .Z(n767) );
  XOR U756 ( .A(n768), .B(n738), .Z(n741) );
  XOR U757 ( .A(p_input[141]), .B(p_input[61]), .Z(n738) );
  XNOR U758 ( .A(p_input[142]), .B(p_input[62]), .Z(n768) );
  XOR U759 ( .A(p_input[137]), .B(p_input[57]), .Z(n733) );
  XNOR U760 ( .A(n749), .B(n748), .Z(n731) );
  XNOR U761 ( .A(n769), .B(n754), .Z(n748) );
  XOR U762 ( .A(p_input[136]), .B(p_input[56]), .Z(n754) );
  XOR U763 ( .A(n745), .B(n753), .Z(n769) );
  XOR U764 ( .A(n770), .B(n750), .Z(n753) );
  XOR U765 ( .A(p_input[134]), .B(p_input[54]), .Z(n750) );
  XNOR U766 ( .A(p_input[135]), .B(p_input[55]), .Z(n770) );
  XOR U767 ( .A(p_input[130]), .B(p_input[50]), .Z(n745) );
  XNOR U768 ( .A(n759), .B(n758), .Z(n749) );
  XOR U769 ( .A(n771), .B(n755), .Z(n758) );
  XOR U770 ( .A(p_input[131]), .B(p_input[51]), .Z(n755) );
  XNOR U771 ( .A(p_input[132]), .B(p_input[52]), .Z(n771) );
  XOR U772 ( .A(p_input[133]), .B(p_input[53]), .Z(n759) );
  XOR U773 ( .A(n772), .B(n773), .Z(n664) );
  AND U774 ( .A(n19), .B(n774), .Z(n773) );
  XNOR U775 ( .A(n775), .B(n772), .Z(n774) );
  XNOR U776 ( .A(n776), .B(n777), .Z(n19) );
  MUX U777 ( .IN0(n670), .IN1(n671), .SEL(n776), .F(n777) );
  AND U778 ( .A(n778), .B(n779), .Z(n671) );
  AND U779 ( .A(n780), .B(n781), .Z(n670) );
  XOR U780 ( .A(n782), .B(n783), .Z(n776) );
  AND U781 ( .A(n784), .B(n785), .Z(n783) );
  XNOR U782 ( .A(n782), .B(n780), .Z(n785) );
  IV U783 ( .A(n688), .Z(n780) );
  XOR U784 ( .A(n786), .B(n787), .Z(n688) );
  XOR U785 ( .A(n788), .B(n781), .Z(n787) );
  AND U786 ( .A(n715), .B(n789), .Z(n781) );
  AND U787 ( .A(n790), .B(n791), .Z(n788) );
  XOR U788 ( .A(n792), .B(n786), .Z(n790) );
  XNOR U789 ( .A(n685), .B(n782), .Z(n784) );
  XOR U790 ( .A(n793), .B(n794), .Z(n685) );
  AND U791 ( .A(n23), .B(n795), .Z(n794) );
  XOR U792 ( .A(n796), .B(n793), .Z(n795) );
  XOR U793 ( .A(n797), .B(n798), .Z(n782) );
  AND U794 ( .A(n799), .B(n800), .Z(n798) );
  XNOR U795 ( .A(n797), .B(n715), .Z(n800) );
  XOR U796 ( .A(n801), .B(n791), .Z(n715) );
  XNOR U797 ( .A(n802), .B(n786), .Z(n791) );
  XOR U798 ( .A(n803), .B(n804), .Z(n786) );
  AND U799 ( .A(n805), .B(n806), .Z(n804) );
  XOR U800 ( .A(n807), .B(n803), .Z(n805) );
  XNOR U801 ( .A(n808), .B(n809), .Z(n802) );
  AND U802 ( .A(n810), .B(n811), .Z(n809) );
  XOR U803 ( .A(n808), .B(n812), .Z(n810) );
  XNOR U804 ( .A(n792), .B(n789), .Z(n801) );
  AND U805 ( .A(n813), .B(n814), .Z(n789) );
  XOR U806 ( .A(n815), .B(n816), .Z(n792) );
  AND U807 ( .A(n817), .B(n818), .Z(n816) );
  XOR U808 ( .A(n815), .B(n819), .Z(n817) );
  XNOR U809 ( .A(n712), .B(n797), .Z(n799) );
  XOR U810 ( .A(n820), .B(n821), .Z(n712) );
  AND U811 ( .A(n23), .B(n822), .Z(n821) );
  XNOR U812 ( .A(n823), .B(n820), .Z(n822) );
  XOR U813 ( .A(n824), .B(n825), .Z(n797) );
  AND U814 ( .A(n826), .B(n827), .Z(n825) );
  XNOR U815 ( .A(n824), .B(n813), .Z(n827) );
  IV U816 ( .A(n763), .Z(n813) );
  XNOR U817 ( .A(n828), .B(n806), .Z(n763) );
  XNOR U818 ( .A(n829), .B(n812), .Z(n806) );
  XOR U819 ( .A(n830), .B(n831), .Z(n812) );
  NOR U820 ( .A(n832), .B(n833), .Z(n831) );
  XNOR U821 ( .A(n830), .B(n834), .Z(n832) );
  XNOR U822 ( .A(n811), .B(n803), .Z(n829) );
  XOR U823 ( .A(n835), .B(n836), .Z(n803) );
  AND U824 ( .A(n837), .B(n838), .Z(n836) );
  XNOR U825 ( .A(n835), .B(n839), .Z(n837) );
  XNOR U826 ( .A(n840), .B(n808), .Z(n811) );
  XOR U827 ( .A(n841), .B(n842), .Z(n808) );
  AND U828 ( .A(n843), .B(n844), .Z(n842) );
  XOR U829 ( .A(n841), .B(n845), .Z(n843) );
  XNOR U830 ( .A(n846), .B(n847), .Z(n840) );
  NOR U831 ( .A(n848), .B(n849), .Z(n847) );
  XOR U832 ( .A(n846), .B(n850), .Z(n848) );
  XNOR U833 ( .A(n807), .B(n814), .Z(n828) );
  NOR U834 ( .A(n775), .B(n851), .Z(n814) );
  XOR U835 ( .A(n819), .B(n818), .Z(n807) );
  XNOR U836 ( .A(n852), .B(n815), .Z(n818) );
  XOR U837 ( .A(n853), .B(n854), .Z(n815) );
  AND U838 ( .A(n855), .B(n856), .Z(n854) );
  XOR U839 ( .A(n853), .B(n857), .Z(n855) );
  XNOR U840 ( .A(n858), .B(n859), .Z(n852) );
  NOR U841 ( .A(n860), .B(n861), .Z(n859) );
  XNOR U842 ( .A(n858), .B(n862), .Z(n860) );
  XOR U843 ( .A(n863), .B(n864), .Z(n819) );
  NOR U844 ( .A(n865), .B(n866), .Z(n864) );
  XNOR U845 ( .A(n863), .B(n867), .Z(n865) );
  XNOR U846 ( .A(n760), .B(n824), .Z(n826) );
  XOR U847 ( .A(n868), .B(n869), .Z(n760) );
  AND U848 ( .A(n23), .B(n870), .Z(n869) );
  XOR U849 ( .A(n871), .B(n868), .Z(n870) );
  AND U850 ( .A(n772), .B(n775), .Z(n824) );
  XOR U851 ( .A(n872), .B(n851), .Z(n775) );
  XNOR U852 ( .A(p_input[128]), .B(p_input[64]), .Z(n851) );
  XOR U853 ( .A(n839), .B(n838), .Z(n872) );
  XNOR U854 ( .A(n873), .B(n845), .Z(n838) );
  XNOR U855 ( .A(n834), .B(n833), .Z(n845) );
  XOR U856 ( .A(n874), .B(n830), .Z(n833) );
  XNOR U857 ( .A(n549), .B(p_input[74]), .Z(n830) );
  XNOR U858 ( .A(p_input[139]), .B(p_input[75]), .Z(n874) );
  XOR U859 ( .A(p_input[140]), .B(p_input[76]), .Z(n834) );
  XNOR U860 ( .A(n844), .B(n835), .Z(n873) );
  XNOR U861 ( .A(n550), .B(p_input[65]), .Z(n835) );
  XOR U862 ( .A(n875), .B(n850), .Z(n844) );
  XNOR U863 ( .A(p_input[143]), .B(p_input[79]), .Z(n850) );
  XOR U864 ( .A(n841), .B(n849), .Z(n875) );
  XOR U865 ( .A(n876), .B(n846), .Z(n849) );
  XOR U866 ( .A(p_input[141]), .B(p_input[77]), .Z(n846) );
  XNOR U867 ( .A(p_input[142]), .B(p_input[78]), .Z(n876) );
  XOR U868 ( .A(p_input[137]), .B(p_input[73]), .Z(n841) );
  XNOR U869 ( .A(n857), .B(n856), .Z(n839) );
  XNOR U870 ( .A(n877), .B(n862), .Z(n856) );
  XOR U871 ( .A(p_input[136]), .B(p_input[72]), .Z(n862) );
  XOR U872 ( .A(n853), .B(n861), .Z(n877) );
  XOR U873 ( .A(n878), .B(n858), .Z(n861) );
  XOR U874 ( .A(p_input[134]), .B(p_input[70]), .Z(n858) );
  XNOR U875 ( .A(p_input[135]), .B(p_input[71]), .Z(n878) );
  XOR U876 ( .A(p_input[130]), .B(p_input[66]), .Z(n853) );
  XNOR U877 ( .A(n867), .B(n866), .Z(n857) );
  XOR U878 ( .A(n879), .B(n863), .Z(n866) );
  XOR U879 ( .A(p_input[131]), .B(p_input[67]), .Z(n863) );
  XNOR U880 ( .A(p_input[132]), .B(p_input[68]), .Z(n879) );
  XOR U881 ( .A(p_input[133]), .B(p_input[69]), .Z(n867) );
  XOR U882 ( .A(n880), .B(n881), .Z(n772) );
  AND U883 ( .A(n23), .B(n882), .Z(n881) );
  XNOR U884 ( .A(n883), .B(n880), .Z(n882) );
  XNOR U885 ( .A(n884), .B(n885), .Z(n23) );
  MUX U886 ( .IN0(n778), .IN1(n779), .SEL(n884), .F(n885) );
  AND U887 ( .A(n886), .B(n887), .Z(n779) );
  AND U888 ( .A(n888), .B(n889), .Z(n778) );
  XOR U889 ( .A(n890), .B(n891), .Z(n884) );
  AND U890 ( .A(n892), .B(n893), .Z(n891) );
  XNOR U891 ( .A(n890), .B(n888), .Z(n893) );
  IV U892 ( .A(n796), .Z(n888) );
  XOR U893 ( .A(n894), .B(n895), .Z(n796) );
  XOR U894 ( .A(n896), .B(n889), .Z(n895) );
  AND U895 ( .A(n823), .B(n897), .Z(n889) );
  AND U896 ( .A(n898), .B(n899), .Z(n896) );
  XOR U897 ( .A(n900), .B(n894), .Z(n898) );
  XNOR U898 ( .A(n793), .B(n890), .Z(n892) );
  XNOR U899 ( .A(n901), .B(n902), .Z(n793) );
  AND U900 ( .A(n26), .B(n903), .Z(n902) );
  XNOR U901 ( .A(n904), .B(n901), .Z(n903) );
  XOR U902 ( .A(n905), .B(n906), .Z(n890) );
  AND U903 ( .A(n907), .B(n908), .Z(n906) );
  XNOR U904 ( .A(n905), .B(n823), .Z(n908) );
  XOR U905 ( .A(n909), .B(n899), .Z(n823) );
  XNOR U906 ( .A(n910), .B(n894), .Z(n899) );
  XOR U907 ( .A(n911), .B(n912), .Z(n894) );
  AND U908 ( .A(n913), .B(n914), .Z(n912) );
  XOR U909 ( .A(n915), .B(n911), .Z(n913) );
  XNOR U910 ( .A(n916), .B(n917), .Z(n910) );
  AND U911 ( .A(n918), .B(n919), .Z(n917) );
  XOR U912 ( .A(n916), .B(n920), .Z(n918) );
  XNOR U913 ( .A(n900), .B(n897), .Z(n909) );
  AND U914 ( .A(n921), .B(n922), .Z(n897) );
  XOR U915 ( .A(n923), .B(n924), .Z(n900) );
  AND U916 ( .A(n925), .B(n926), .Z(n924) );
  XOR U917 ( .A(n923), .B(n927), .Z(n925) );
  XNOR U918 ( .A(n820), .B(n905), .Z(n907) );
  XNOR U919 ( .A(n928), .B(n929), .Z(n820) );
  AND U920 ( .A(n26), .B(n930), .Z(n929) );
  XOR U921 ( .A(n931), .B(n928), .Z(n930) );
  XOR U922 ( .A(n932), .B(n933), .Z(n905) );
  AND U923 ( .A(n934), .B(n935), .Z(n933) );
  XNOR U924 ( .A(n932), .B(n921), .Z(n935) );
  IV U925 ( .A(n871), .Z(n921) );
  XNOR U926 ( .A(n936), .B(n914), .Z(n871) );
  XNOR U927 ( .A(n937), .B(n920), .Z(n914) );
  XOR U928 ( .A(n938), .B(n939), .Z(n920) );
  NOR U929 ( .A(n940), .B(n941), .Z(n939) );
  XNOR U930 ( .A(n938), .B(n942), .Z(n940) );
  XNOR U931 ( .A(n919), .B(n911), .Z(n937) );
  XOR U932 ( .A(n943), .B(n944), .Z(n911) );
  AND U933 ( .A(n945), .B(n946), .Z(n944) );
  XNOR U934 ( .A(n943), .B(n947), .Z(n945) );
  XNOR U935 ( .A(n948), .B(n916), .Z(n919) );
  XOR U936 ( .A(n949), .B(n950), .Z(n916) );
  AND U937 ( .A(n951), .B(n952), .Z(n950) );
  XOR U938 ( .A(n949), .B(n953), .Z(n951) );
  XNOR U939 ( .A(n954), .B(n955), .Z(n948) );
  NOR U940 ( .A(n956), .B(n957), .Z(n955) );
  XOR U941 ( .A(n954), .B(n958), .Z(n956) );
  XNOR U942 ( .A(n915), .B(n922), .Z(n936) );
  NOR U943 ( .A(n883), .B(n959), .Z(n922) );
  XOR U944 ( .A(n927), .B(n926), .Z(n915) );
  XNOR U945 ( .A(n960), .B(n923), .Z(n926) );
  XOR U946 ( .A(n961), .B(n962), .Z(n923) );
  AND U947 ( .A(n963), .B(n964), .Z(n962) );
  XOR U948 ( .A(n961), .B(n965), .Z(n963) );
  XNOR U949 ( .A(n966), .B(n967), .Z(n960) );
  NOR U950 ( .A(n968), .B(n969), .Z(n967) );
  XNOR U951 ( .A(n966), .B(n970), .Z(n968) );
  XOR U952 ( .A(n971), .B(n972), .Z(n927) );
  NOR U953 ( .A(n973), .B(n974), .Z(n972) );
  XNOR U954 ( .A(n971), .B(n975), .Z(n973) );
  XNOR U955 ( .A(n868), .B(n932), .Z(n934) );
  XNOR U956 ( .A(n976), .B(n977), .Z(n868) );
  AND U957 ( .A(n26), .B(n978), .Z(n977) );
  XNOR U958 ( .A(n979), .B(n976), .Z(n978) );
  AND U959 ( .A(n880), .B(n883), .Z(n932) );
  XOR U960 ( .A(n980), .B(n959), .Z(n883) );
  XNOR U961 ( .A(p_input[128]), .B(p_input[80]), .Z(n959) );
  XOR U962 ( .A(n947), .B(n946), .Z(n980) );
  XNOR U963 ( .A(n981), .B(n953), .Z(n946) );
  XNOR U964 ( .A(n942), .B(n941), .Z(n953) );
  XOR U965 ( .A(n982), .B(n938), .Z(n941) );
  XNOR U966 ( .A(n549), .B(p_input[90]), .Z(n938) );
  XNOR U967 ( .A(p_input[139]), .B(p_input[91]), .Z(n982) );
  XOR U968 ( .A(p_input[140]), .B(p_input[92]), .Z(n942) );
  XNOR U969 ( .A(n952), .B(n943), .Z(n981) );
  XNOR U970 ( .A(n550), .B(p_input[81]), .Z(n943) );
  XOR U971 ( .A(n983), .B(n958), .Z(n952) );
  XNOR U972 ( .A(p_input[143]), .B(p_input[95]), .Z(n958) );
  XOR U973 ( .A(n949), .B(n957), .Z(n983) );
  XOR U974 ( .A(n984), .B(n954), .Z(n957) );
  XOR U975 ( .A(p_input[141]), .B(p_input[93]), .Z(n954) );
  XNOR U976 ( .A(p_input[142]), .B(p_input[94]), .Z(n984) );
  XOR U977 ( .A(p_input[137]), .B(p_input[89]), .Z(n949) );
  XNOR U978 ( .A(n965), .B(n964), .Z(n947) );
  XNOR U979 ( .A(n985), .B(n970), .Z(n964) );
  XOR U980 ( .A(p_input[136]), .B(p_input[88]), .Z(n970) );
  XOR U981 ( .A(n961), .B(n969), .Z(n985) );
  XOR U982 ( .A(n986), .B(n966), .Z(n969) );
  XOR U983 ( .A(p_input[134]), .B(p_input[86]), .Z(n966) );
  XNOR U984 ( .A(p_input[135]), .B(p_input[87]), .Z(n986) );
  XOR U985 ( .A(p_input[130]), .B(p_input[82]), .Z(n961) );
  XNOR U986 ( .A(n975), .B(n974), .Z(n965) );
  XOR U987 ( .A(n987), .B(n971), .Z(n974) );
  XOR U988 ( .A(p_input[131]), .B(p_input[83]), .Z(n971) );
  XNOR U989 ( .A(p_input[132]), .B(p_input[84]), .Z(n987) );
  XOR U990 ( .A(p_input[133]), .B(p_input[85]), .Z(n975) );
  XOR U991 ( .A(n988), .B(n989), .Z(n880) );
  AND U992 ( .A(n26), .B(n990), .Z(n989) );
  XNOR U993 ( .A(n991), .B(n988), .Z(n990) );
  XNOR U994 ( .A(n992), .B(n993), .Z(n26) );
  MUX U995 ( .IN0(n886), .IN1(n887), .SEL(n992), .F(n993) );
  AND U996 ( .A(n901), .B(n994), .Z(n887) );
  AND U997 ( .A(n995), .B(n996), .Z(n886) );
  XOR U998 ( .A(n997), .B(n998), .Z(n992) );
  AND U999 ( .A(n999), .B(n1000), .Z(n998) );
  XNOR U1000 ( .A(n997), .B(n995), .Z(n1000) );
  IV U1001 ( .A(n904), .Z(n995) );
  XOR U1002 ( .A(n1001), .B(n1002), .Z(n904) );
  XOR U1003 ( .A(n1003), .B(n996), .Z(n1002) );
  AND U1004 ( .A(n931), .B(n1004), .Z(n996) );
  AND U1005 ( .A(n1005), .B(n1006), .Z(n1003) );
  XOR U1006 ( .A(n1007), .B(n1001), .Z(n1005) );
  XNOR U1007 ( .A(n1008), .B(n997), .Z(n999) );
  IV U1008 ( .A(n901), .Z(n1008) );
  XNOR U1009 ( .A(n1009), .B(n1010), .Z(n901) );
  XOR U1010 ( .A(n1011), .B(n994), .Z(n1010) );
  AND U1011 ( .A(n928), .B(n1012), .Z(n994) );
  AND U1012 ( .A(n1013), .B(n1014), .Z(n1011) );
  XNOR U1013 ( .A(n1009), .B(n1015), .Z(n1013) );
  XOR U1014 ( .A(n1016), .B(n1017), .Z(n997) );
  AND U1015 ( .A(n1018), .B(n1019), .Z(n1017) );
  XNOR U1016 ( .A(n1016), .B(n931), .Z(n1019) );
  XOR U1017 ( .A(n1020), .B(n1006), .Z(n931) );
  XNOR U1018 ( .A(n1021), .B(n1001), .Z(n1006) );
  XOR U1019 ( .A(n1022), .B(n1023), .Z(n1001) );
  AND U1020 ( .A(n1024), .B(n1025), .Z(n1023) );
  XOR U1021 ( .A(n1026), .B(n1022), .Z(n1024) );
  XNOR U1022 ( .A(n1027), .B(n1028), .Z(n1021) );
  AND U1023 ( .A(n1029), .B(n1030), .Z(n1028) );
  XOR U1024 ( .A(n1027), .B(n1031), .Z(n1029) );
  XNOR U1025 ( .A(n1007), .B(n1004), .Z(n1020) );
  AND U1026 ( .A(n1032), .B(n1033), .Z(n1004) );
  XOR U1027 ( .A(n1034), .B(n1035), .Z(n1007) );
  AND U1028 ( .A(n1036), .B(n1037), .Z(n1035) );
  XOR U1029 ( .A(n1034), .B(n1038), .Z(n1036) );
  XOR U1030 ( .A(n928), .B(n1016), .Z(n1018) );
  XNOR U1031 ( .A(n1039), .B(n1015), .Z(n928) );
  XNOR U1032 ( .A(n1040), .B(n1041), .Z(n1015) );
  AND U1033 ( .A(n1042), .B(n1043), .Z(n1041) );
  XOR U1034 ( .A(n1040), .B(n1044), .Z(n1042) );
  XNOR U1035 ( .A(n1014), .B(n1012), .Z(n1039) );
  AND U1036 ( .A(n976), .B(n1045), .Z(n1012) );
  XNOR U1037 ( .A(n1046), .B(n1009), .Z(n1014) );
  XOR U1038 ( .A(n1047), .B(n1048), .Z(n1009) );
  AND U1039 ( .A(n1049), .B(n1050), .Z(n1048) );
  XOR U1040 ( .A(n1047), .B(n1051), .Z(n1049) );
  XNOR U1041 ( .A(n1052), .B(n1053), .Z(n1046) );
  AND U1042 ( .A(n1054), .B(n1055), .Z(n1053) );
  XNOR U1043 ( .A(n1052), .B(n1056), .Z(n1054) );
  XOR U1044 ( .A(n1057), .B(n1058), .Z(n1016) );
  AND U1045 ( .A(n1059), .B(n1060), .Z(n1058) );
  XNOR U1046 ( .A(n1057), .B(n1032), .Z(n1060) );
  IV U1047 ( .A(n979), .Z(n1032) );
  XNOR U1048 ( .A(n1061), .B(n1025), .Z(n979) );
  XNOR U1049 ( .A(n1062), .B(n1031), .Z(n1025) );
  XNOR U1050 ( .A(n1063), .B(n1064), .Z(n1031) );
  NOR U1051 ( .A(n1065), .B(n1066), .Z(n1064) );
  XOR U1052 ( .A(n1063), .B(n1067), .Z(n1065) );
  XNOR U1053 ( .A(n1030), .B(n1022), .Z(n1062) );
  XOR U1054 ( .A(n1068), .B(n1069), .Z(n1022) );
  AND U1055 ( .A(n1070), .B(n1071), .Z(n1069) );
  XOR U1056 ( .A(n1068), .B(n1072), .Z(n1070) );
  XNOR U1057 ( .A(n1073), .B(n1027), .Z(n1030) );
  XOR U1058 ( .A(n1074), .B(n1075), .Z(n1027) );
  NOR U1059 ( .A(n1076), .B(n1077), .Z(n1075) );
  XNOR U1060 ( .A(n1074), .B(n1078), .Z(n1076) );
  XNOR U1061 ( .A(n1079), .B(n1080), .Z(n1073) );
  NOR U1062 ( .A(n1081), .B(n1082), .Z(n1080) );
  XNOR U1063 ( .A(n1079), .B(n1083), .Z(n1081) );
  XNOR U1064 ( .A(n1026), .B(n1033), .Z(n1061) );
  NOR U1065 ( .A(n991), .B(n1084), .Z(n1033) );
  XOR U1066 ( .A(n1038), .B(n1037), .Z(n1026) );
  XNOR U1067 ( .A(n1085), .B(n1034), .Z(n1037) );
  XOR U1068 ( .A(n1086), .B(n1087), .Z(n1034) );
  NOR U1069 ( .A(n1088), .B(n1089), .Z(n1087) );
  XNOR U1070 ( .A(n1086), .B(n1090), .Z(n1088) );
  XNOR U1071 ( .A(n1091), .B(n1092), .Z(n1085) );
  NOR U1072 ( .A(n1093), .B(n1094), .Z(n1092) );
  XNOR U1073 ( .A(n1091), .B(n1095), .Z(n1093) );
  XOR U1074 ( .A(n1096), .B(n1097), .Z(n1038) );
  NOR U1075 ( .A(n1098), .B(n1099), .Z(n1097) );
  XNOR U1076 ( .A(n1096), .B(n1100), .Z(n1098) );
  XNOR U1077 ( .A(n1101), .B(n1057), .Z(n1059) );
  IV U1078 ( .A(n976), .Z(n1101) );
  XOR U1079 ( .A(n1102), .B(n1051), .Z(n976) );
  XOR U1080 ( .A(n1044), .B(n1043), .Z(n1051) );
  XNOR U1081 ( .A(n1103), .B(n1040), .Z(n1043) );
  XOR U1082 ( .A(n1104), .B(n1105), .Z(n1040) );
  AND U1083 ( .A(n1106), .B(n1107), .Z(n1105) );
  XNOR U1084 ( .A(n1108), .B(n1109), .Z(n1106) );
  IV U1085 ( .A(n1104), .Z(n1108) );
  XNOR U1086 ( .A(n1110), .B(n1111), .Z(n1103) );
  NOR U1087 ( .A(n1112), .B(n1113), .Z(n1111) );
  XNOR U1088 ( .A(n1110), .B(n1114), .Z(n1112) );
  XOR U1089 ( .A(n1115), .B(n1116), .Z(n1044) );
  AND U1090 ( .A(n1117), .B(n1118), .Z(n1116) );
  XOR U1091 ( .A(n1115), .B(n1119), .Z(n1117) );
  XNOR U1092 ( .A(n1050), .B(n1045), .Z(n1102) );
  AND U1093 ( .A(n988), .B(n1120), .Z(n1045) );
  XOR U1094 ( .A(n1121), .B(n1056), .Z(n1050) );
  XNOR U1095 ( .A(n1122), .B(n1123), .Z(n1056) );
  NOR U1096 ( .A(n1124), .B(n1125), .Z(n1123) );
  XNOR U1097 ( .A(n1122), .B(n1126), .Z(n1124) );
  XNOR U1098 ( .A(n1055), .B(n1047), .Z(n1121) );
  XOR U1099 ( .A(n1127), .B(n1128), .Z(n1047) );
  AND U1100 ( .A(n1129), .B(n1130), .Z(n1128) );
  XOR U1101 ( .A(n1127), .B(n1131), .Z(n1129) );
  XNOR U1102 ( .A(n1132), .B(n1052), .Z(n1055) );
  XOR U1103 ( .A(n1133), .B(n1134), .Z(n1052) );
  AND U1104 ( .A(n1135), .B(n1136), .Z(n1134) );
  XOR U1105 ( .A(n1133), .B(n1137), .Z(n1135) );
  XNOR U1106 ( .A(n1138), .B(n1139), .Z(n1132) );
  NOR U1107 ( .A(n1140), .B(n1141), .Z(n1139) );
  XOR U1108 ( .A(n1138), .B(n1142), .Z(n1140) );
  AND U1109 ( .A(n988), .B(n991), .Z(n1057) );
  XOR U1110 ( .A(n1143), .B(n1084), .Z(n991) );
  XNOR U1111 ( .A(p_input[128]), .B(p_input[96]), .Z(n1084) );
  XNOR U1112 ( .A(n1072), .B(n1071), .Z(n1143) );
  XNOR U1113 ( .A(n1144), .B(n1078), .Z(n1071) );
  XNOR U1114 ( .A(n1067), .B(n1066), .Z(n1078) );
  XNOR U1115 ( .A(n1145), .B(n1063), .Z(n1066) );
  XNOR U1116 ( .A(p_input[106]), .B(p_input[138]), .Z(n1063) );
  XOR U1117 ( .A(p_input[107]), .B(n438), .Z(n1145) );
  XOR U1118 ( .A(p_input[108]), .B(p_input[140]), .Z(n1067) );
  XOR U1119 ( .A(n1077), .B(n1068), .Z(n1144) );
  XNOR U1120 ( .A(n550), .B(p_input[97]), .Z(n1068) );
  IV U1121 ( .A(p_input[129]), .Z(n550) );
  XOR U1122 ( .A(n1146), .B(n1083), .Z(n1077) );
  XOR U1123 ( .A(p_input[111]), .B(p_input[143]), .Z(n1083) );
  XOR U1124 ( .A(n1074), .B(n1082), .Z(n1146) );
  XOR U1125 ( .A(n1147), .B(n1079), .Z(n1082) );
  XOR U1126 ( .A(p_input[109]), .B(p_input[141]), .Z(n1079) );
  XNOR U1127 ( .A(p_input[110]), .B(p_input[142]), .Z(n1147) );
  XOR U1128 ( .A(p_input[105]), .B(p_input[137]), .Z(n1074) );
  XNOR U1129 ( .A(n1090), .B(n1089), .Z(n1072) );
  XOR U1130 ( .A(n1148), .B(n1095), .Z(n1089) );
  XOR U1131 ( .A(p_input[104]), .B(p_input[136]), .Z(n1095) );
  XOR U1132 ( .A(n1086), .B(n1094), .Z(n1148) );
  XOR U1133 ( .A(n1149), .B(n1091), .Z(n1094) );
  XOR U1134 ( .A(p_input[102]), .B(p_input[134]), .Z(n1091) );
  XNOR U1135 ( .A(p_input[103]), .B(p_input[135]), .Z(n1149) );
  XOR U1136 ( .A(p_input[130]), .B(p_input[98]), .Z(n1086) );
  XNOR U1137 ( .A(n1100), .B(n1099), .Z(n1090) );
  XOR U1138 ( .A(n1150), .B(n1096), .Z(n1099) );
  XOR U1139 ( .A(p_input[131]), .B(p_input[99]), .Z(n1096) );
  XNOR U1140 ( .A(p_input[100]), .B(p_input[132]), .Z(n1150) );
  XOR U1141 ( .A(p_input[101]), .B(p_input[133]), .Z(n1100) );
  XOR U1142 ( .A(n1151), .B(n1131), .Z(n988) );
  XOR U1143 ( .A(n1109), .B(n1107), .Z(n1131) );
  XNOR U1144 ( .A(n1152), .B(n1114), .Z(n1107) );
  XOR U1145 ( .A(\knn_comb_/min_val_out[0][8] ), .B(p_input[136]), .Z(n1114)
         );
  XOR U1146 ( .A(n1104), .B(n1113), .Z(n1152) );
  XOR U1147 ( .A(n1153), .B(n1110), .Z(n1113) );
  XOR U1148 ( .A(\knn_comb_/min_val_out[0][6] ), .B(p_input[134]), .Z(n1110)
         );
  XNOR U1149 ( .A(\knn_comb_/min_val_out[0][7] ), .B(p_input[135]), .Z(n1153)
         );
  XOR U1150 ( .A(\knn_comb_/min_val_out[0][2] ), .B(p_input[130]), .Z(n1104)
         );
  XOR U1151 ( .A(n1119), .B(n1118), .Z(n1109) );
  XNOR U1152 ( .A(n1154), .B(n1115), .Z(n1118) );
  XOR U1153 ( .A(\knn_comb_/min_val_out[0][3] ), .B(p_input[131]), .Z(n1115)
         );
  XNOR U1154 ( .A(\knn_comb_/min_val_out[0][4] ), .B(p_input[132]), .Z(n1154)
         );
  XOR U1155 ( .A(\knn_comb_/min_val_out[0][5] ), .B(p_input[133]), .Z(n1119)
         );
  XNOR U1156 ( .A(n1130), .B(n1120), .Z(n1151) );
  XOR U1157 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[128]), .Z(n1120)
         );
  XNOR U1158 ( .A(n1155), .B(n1137), .Z(n1130) );
  XNOR U1159 ( .A(n1126), .B(n1125), .Z(n1137) );
  XOR U1160 ( .A(n1156), .B(n1122), .Z(n1125) );
  XNOR U1161 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n549), .Z(n1122) );
  IV U1162 ( .A(p_input[138]), .Z(n549) );
  XOR U1163 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n438), .Z(n1156) );
  IV U1164 ( .A(p_input[139]), .Z(n438) );
  XOR U1165 ( .A(\knn_comb_/min_val_out[0][12] ), .B(p_input[140]), .Z(n1126)
         );
  XNOR U1166 ( .A(n1136), .B(n1127), .Z(n1155) );
  XOR U1167 ( .A(\knn_comb_/min_val_out[0][1] ), .B(p_input[129]), .Z(n1127)
         );
  XOR U1168 ( .A(n1157), .B(n1142), .Z(n1136) );
  XNOR U1169 ( .A(\knn_comb_/min_val_out[0][15] ), .B(p_input[143]), .Z(n1142)
         );
  XOR U1170 ( .A(n1133), .B(n1141), .Z(n1157) );
  XOR U1171 ( .A(n1158), .B(n1138), .Z(n1141) );
  XOR U1172 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[141]), .Z(n1138)
         );
  XNOR U1173 ( .A(\knn_comb_/min_val_out[0][14] ), .B(p_input[142]), .Z(n1158)
         );
  XOR U1174 ( .A(\knn_comb_/min_val_out[0][9] ), .B(p_input[137]), .Z(n1133)
         );
endmodule

