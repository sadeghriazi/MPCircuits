
module knn_comb_BMR_W32_K2_N4 ( p_input, o );
  input [159:0] p_input;
  output [63:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/min_val_out[0][16] , \knn_comb_/min_val_out[0][17] ,
         \knn_comb_/min_val_out[0][18] , \knn_comb_/min_val_out[0][19] ,
         \knn_comb_/min_val_out[0][20] , \knn_comb_/min_val_out[0][21] ,
         \knn_comb_/min_val_out[0][22] , \knn_comb_/min_val_out[0][23] ,
         \knn_comb_/min_val_out[0][24] , \knn_comb_/min_val_out[0][25] ,
         \knn_comb_/min_val_out[0][26] , \knn_comb_/min_val_out[0][27] ,
         \knn_comb_/min_val_out[0][28] , \knn_comb_/min_val_out[0][29] ,
         \knn_comb_/min_val_out[0][30] , \knn_comb_/min_val_out[0][31] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][31] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547;
  assign \knn_comb_/min_val_out[0][0]  = p_input[96];
  assign \knn_comb_/min_val_out[0][1]  = p_input[97];
  assign \knn_comb_/min_val_out[0][2]  = p_input[98];
  assign \knn_comb_/min_val_out[0][3]  = p_input[99];
  assign \knn_comb_/min_val_out[0][4]  = p_input[100];
  assign \knn_comb_/min_val_out[0][5]  = p_input[101];
  assign \knn_comb_/min_val_out[0][6]  = p_input[102];
  assign \knn_comb_/min_val_out[0][7]  = p_input[103];
  assign \knn_comb_/min_val_out[0][8]  = p_input[104];
  assign \knn_comb_/min_val_out[0][9]  = p_input[105];
  assign \knn_comb_/min_val_out[0][10]  = p_input[106];
  assign \knn_comb_/min_val_out[0][11]  = p_input[107];
  assign \knn_comb_/min_val_out[0][12]  = p_input[108];
  assign \knn_comb_/min_val_out[0][13]  = p_input[109];
  assign \knn_comb_/min_val_out[0][14]  = p_input[110];
  assign \knn_comb_/min_val_out[0][15]  = p_input[111];
  assign \knn_comb_/min_val_out[0][16]  = p_input[112];
  assign \knn_comb_/min_val_out[0][17]  = p_input[113];
  assign \knn_comb_/min_val_out[0][18]  = p_input[114];
  assign \knn_comb_/min_val_out[0][19]  = p_input[115];
  assign \knn_comb_/min_val_out[0][20]  = p_input[116];
  assign \knn_comb_/min_val_out[0][21]  = p_input[117];
  assign \knn_comb_/min_val_out[0][22]  = p_input[118];
  assign \knn_comb_/min_val_out[0][23]  = p_input[119];
  assign \knn_comb_/min_val_out[0][24]  = p_input[120];
  assign \knn_comb_/min_val_out[0][25]  = p_input[121];
  assign \knn_comb_/min_val_out[0][26]  = p_input[122];
  assign \knn_comb_/min_val_out[0][27]  = p_input[123];
  assign \knn_comb_/min_val_out[0][28]  = p_input[124];
  assign \knn_comb_/min_val_out[0][29]  = p_input[125];
  assign \knn_comb_/min_val_out[0][30]  = p_input[126];
  assign \knn_comb_/min_val_out[0][31]  = p_input[127];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][0]  = p_input[64];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][1]  = p_input[65];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][2]  = p_input[66];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][3]  = p_input[67];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][4]  = p_input[68];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][5]  = p_input[69];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][6]  = p_input[70];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][7]  = p_input[71];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][8]  = p_input[72];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][9]  = p_input[73];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][10]  = p_input[74];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][11]  = p_input[75];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][12]  = p_input[76];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][13]  = p_input[77];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][14]  = p_input[78];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][15]  = p_input[79];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][16]  = p_input[80];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][17]  = p_input[81];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][18]  = p_input[82];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][19]  = p_input[83];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][20]  = p_input[84];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][21]  = p_input[85];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][22]  = p_input[86];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][23]  = p_input[87];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][24]  = p_input[88];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][25]  = p_input[89];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][26]  = p_input[90];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][27]  = p_input[91];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][28]  = p_input[92];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][29]  = p_input[93];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][30]  = p_input[94];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][31]  = p_input[95];

  XOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  XOR U2 ( .A(n3), .B(n4), .Z(o[8]) );
  XOR U3 ( .A(n5), .B(n6), .Z(o[7]) );
  XOR U4 ( .A(n7), .B(n8), .Z(o[6]) );
  XOR U5 ( .A(n9), .B(n10), .Z(o[63]) );
  XOR U6 ( .A(n11), .B(n12), .Z(o[62]) );
  XOR U7 ( .A(n13), .B(n14), .Z(o[61]) );
  XOR U8 ( .A(n15), .B(n16), .Z(o[60]) );
  XOR U9 ( .A(n17), .B(n18), .Z(o[5]) );
  XOR U10 ( .A(n19), .B(n20), .Z(o[59]) );
  XOR U11 ( .A(n21), .B(n22), .Z(o[58]) );
  XOR U12 ( .A(n23), .B(n24), .Z(o[57]) );
  XOR U13 ( .A(n25), .B(n26), .Z(o[56]) );
  XOR U14 ( .A(n27), .B(n28), .Z(o[55]) );
  XOR U15 ( .A(n29), .B(n30), .Z(o[54]) );
  XOR U16 ( .A(n31), .B(n32), .Z(o[53]) );
  XOR U17 ( .A(n33), .B(n34), .Z(o[52]) );
  XOR U18 ( .A(n35), .B(n36), .Z(o[51]) );
  XOR U19 ( .A(n37), .B(n38), .Z(o[50]) );
  XOR U20 ( .A(n39), .B(n40), .Z(o[4]) );
  XOR U21 ( .A(n41), .B(n42), .Z(o[49]) );
  XOR U22 ( .A(n43), .B(n44), .Z(o[48]) );
  XOR U23 ( .A(n45), .B(n46), .Z(o[47]) );
  XOR U24 ( .A(n47), .B(n48), .Z(o[46]) );
  XOR U25 ( .A(n49), .B(n50), .Z(o[45]) );
  XOR U26 ( .A(n51), .B(n52), .Z(o[44]) );
  XOR U27 ( .A(n53), .B(n54), .Z(o[43]) );
  XOR U28 ( .A(n55), .B(n56), .Z(o[42]) );
  XOR U29 ( .A(n1), .B(n57), .Z(o[41]) );
  AND U30 ( .A(n58), .B(n59), .Z(n1) );
  XOR U31 ( .A(n2), .B(n57), .Z(n59) );
  XOR U32 ( .A(n60), .B(n61), .Z(n57) );
  AND U33 ( .A(n62), .B(n63), .Z(n61) );
  XOR U34 ( .A(p_input[9]), .B(n60), .Z(n63) );
  XOR U35 ( .A(n64), .B(n65), .Z(n60) );
  AND U36 ( .A(n66), .B(n67), .Z(n65) );
  XNOR U37 ( .A(n68), .B(n69), .Z(n2) );
  AND U38 ( .A(n70), .B(n67), .Z(n69) );
  XOR U39 ( .A(n71), .B(n64), .Z(n67) );
  XOR U40 ( .A(n72), .B(n73), .Z(n64) );
  AND U41 ( .A(n74), .B(n75), .Z(n73) );
  XOR U42 ( .A(p_input[41]), .B(n72), .Z(n75) );
  XOR U43 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .B(n76), .Z(n72) );
  AND U44 ( .A(n77), .B(n78), .Z(n76) );
  IV U45 ( .A(n71), .Z(n68) );
  XOR U46 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n79), .Z(n71) );
  AND U47 ( .A(n80), .B(n78), .Z(n79) );
  XNOR U48 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n81), .Z(n78) );
  IV U49 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .Z(n81) );
  XOR U50 ( .A(n3), .B(n82), .Z(o[40]) );
  AND U51 ( .A(n58), .B(n83), .Z(n3) );
  XOR U52 ( .A(n4), .B(n82), .Z(n83) );
  XOR U53 ( .A(n84), .B(n85), .Z(n82) );
  AND U54 ( .A(n62), .B(n86), .Z(n85) );
  XOR U55 ( .A(p_input[8]), .B(n84), .Z(n86) );
  XOR U56 ( .A(n87), .B(n88), .Z(n84) );
  AND U57 ( .A(n66), .B(n89), .Z(n88) );
  XNOR U58 ( .A(n90), .B(n91), .Z(n4) );
  AND U59 ( .A(n70), .B(n89), .Z(n91) );
  XOR U60 ( .A(n92), .B(n87), .Z(n89) );
  XOR U61 ( .A(n93), .B(n94), .Z(n87) );
  AND U62 ( .A(n74), .B(n95), .Z(n94) );
  XOR U63 ( .A(p_input[40]), .B(n93), .Z(n95) );
  XOR U64 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .B(n96), .Z(n93) );
  AND U65 ( .A(n77), .B(n97), .Z(n96) );
  IV U66 ( .A(n92), .Z(n90) );
  XOR U67 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n98), .Z(n92) );
  AND U68 ( .A(n80), .B(n97), .Z(n98) );
  XOR U69 ( .A(\knn_comb_/min_val_out[0][8] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .Z(n97) );
  XOR U70 ( .A(n99), .B(n100), .Z(o[3]) );
  XOR U71 ( .A(n5), .B(n101), .Z(o[39]) );
  AND U72 ( .A(n58), .B(n102), .Z(n5) );
  XOR U73 ( .A(n6), .B(n101), .Z(n102) );
  XOR U74 ( .A(n103), .B(n104), .Z(n101) );
  AND U75 ( .A(n62), .B(n105), .Z(n104) );
  XOR U76 ( .A(p_input[7]), .B(n103), .Z(n105) );
  XOR U77 ( .A(n106), .B(n107), .Z(n103) );
  AND U78 ( .A(n66), .B(n108), .Z(n107) );
  XNOR U79 ( .A(n109), .B(n110), .Z(n6) );
  AND U80 ( .A(n70), .B(n108), .Z(n110) );
  XOR U81 ( .A(n111), .B(n106), .Z(n108) );
  XOR U82 ( .A(n112), .B(n113), .Z(n106) );
  AND U83 ( .A(n74), .B(n114), .Z(n113) );
  XOR U84 ( .A(p_input[39]), .B(n112), .Z(n114) );
  XOR U85 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(n115), .Z(
        n112) );
  AND U86 ( .A(n77), .B(n116), .Z(n115) );
  IV U87 ( .A(n111), .Z(n109) );
  XOR U88 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n117), .Z(n111) );
  AND U89 ( .A(n80), .B(n116), .Z(n117) );
  XOR U90 ( .A(\knn_comb_/min_val_out[0][7] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .Z(n116) );
  XOR U91 ( .A(n7), .B(n118), .Z(o[38]) );
  AND U92 ( .A(n58), .B(n119), .Z(n7) );
  XOR U93 ( .A(n8), .B(n118), .Z(n119) );
  XOR U94 ( .A(n120), .B(n121), .Z(n118) );
  AND U95 ( .A(n62), .B(n122), .Z(n121) );
  XOR U96 ( .A(p_input[6]), .B(n120), .Z(n122) );
  XOR U97 ( .A(n123), .B(n124), .Z(n120) );
  AND U98 ( .A(n66), .B(n125), .Z(n124) );
  XNOR U99 ( .A(n126), .B(n127), .Z(n8) );
  AND U100 ( .A(n70), .B(n125), .Z(n127) );
  XOR U101 ( .A(n128), .B(n123), .Z(n125) );
  XOR U102 ( .A(n129), .B(n130), .Z(n123) );
  AND U103 ( .A(n74), .B(n131), .Z(n130) );
  XOR U104 ( .A(p_input[38]), .B(n129), .Z(n131) );
  XOR U105 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .B(n132), .Z(
        n129) );
  AND U106 ( .A(n77), .B(n133), .Z(n132) );
  IV U107 ( .A(n128), .Z(n126) );
  XOR U108 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n134), .Z(n128) );
  AND U109 ( .A(n80), .B(n133), .Z(n134) );
  XOR U110 ( .A(\knn_comb_/min_val_out[0][6] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .Z(n133) );
  XOR U111 ( .A(n17), .B(n135), .Z(o[37]) );
  AND U112 ( .A(n58), .B(n136), .Z(n17) );
  XOR U113 ( .A(n18), .B(n135), .Z(n136) );
  XOR U114 ( .A(n137), .B(n138), .Z(n135) );
  AND U115 ( .A(n62), .B(n139), .Z(n138) );
  XOR U116 ( .A(p_input[5]), .B(n137), .Z(n139) );
  XOR U117 ( .A(n140), .B(n141), .Z(n137) );
  AND U118 ( .A(n66), .B(n142), .Z(n141) );
  XNOR U119 ( .A(n143), .B(n144), .Z(n18) );
  AND U120 ( .A(n70), .B(n142), .Z(n144) );
  XOR U121 ( .A(n145), .B(n140), .Z(n142) );
  XOR U122 ( .A(n146), .B(n147), .Z(n140) );
  AND U123 ( .A(n74), .B(n148), .Z(n147) );
  XOR U124 ( .A(p_input[37]), .B(n146), .Z(n148) );
  XOR U125 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(n149), .Z(
        n146) );
  AND U126 ( .A(n77), .B(n150), .Z(n149) );
  IV U127 ( .A(n145), .Z(n143) );
  XOR U128 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n151), .Z(n145) );
  AND U129 ( .A(n80), .B(n150), .Z(n151) );
  XOR U130 ( .A(\knn_comb_/min_val_out[0][5] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .Z(n150) );
  XOR U131 ( .A(n39), .B(n152), .Z(o[36]) );
  AND U132 ( .A(n58), .B(n153), .Z(n39) );
  XOR U133 ( .A(n40), .B(n152), .Z(n153) );
  XOR U134 ( .A(n154), .B(n155), .Z(n152) );
  AND U135 ( .A(n62), .B(n156), .Z(n155) );
  XOR U136 ( .A(p_input[4]), .B(n154), .Z(n156) );
  XOR U137 ( .A(n157), .B(n158), .Z(n154) );
  AND U138 ( .A(n66), .B(n159), .Z(n158) );
  XNOR U139 ( .A(n160), .B(n161), .Z(n40) );
  AND U140 ( .A(n70), .B(n159), .Z(n161) );
  XOR U141 ( .A(n162), .B(n157), .Z(n159) );
  XOR U142 ( .A(n163), .B(n164), .Z(n157) );
  AND U143 ( .A(n74), .B(n165), .Z(n164) );
  XOR U144 ( .A(p_input[36]), .B(n163), .Z(n165) );
  XOR U145 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(n166), .Z(
        n163) );
  AND U146 ( .A(n77), .B(n167), .Z(n166) );
  IV U147 ( .A(n162), .Z(n160) );
  XOR U148 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n168), .Z(n162) );
  AND U149 ( .A(n80), .B(n167), .Z(n168) );
  XOR U150 ( .A(\knn_comb_/min_val_out[0][4] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .Z(n167) );
  XOR U151 ( .A(n99), .B(n169), .Z(o[35]) );
  AND U152 ( .A(n58), .B(n170), .Z(n99) );
  XOR U153 ( .A(n100), .B(n169), .Z(n170) );
  XOR U154 ( .A(n171), .B(n172), .Z(n169) );
  AND U155 ( .A(n62), .B(n173), .Z(n172) );
  XOR U156 ( .A(p_input[3]), .B(n171), .Z(n173) );
  XOR U157 ( .A(n174), .B(n175), .Z(n171) );
  AND U158 ( .A(n66), .B(n176), .Z(n175) );
  XNOR U159 ( .A(n177), .B(n178), .Z(n100) );
  AND U160 ( .A(n70), .B(n176), .Z(n178) );
  XOR U161 ( .A(n179), .B(n174), .Z(n176) );
  XOR U162 ( .A(n180), .B(n181), .Z(n174) );
  AND U163 ( .A(n74), .B(n182), .Z(n181) );
  XOR U164 ( .A(p_input[35]), .B(n180), .Z(n182) );
  XOR U165 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .B(n183), .Z(
        n180) );
  AND U166 ( .A(n77), .B(n184), .Z(n183) );
  IV U167 ( .A(n179), .Z(n177) );
  XOR U168 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n185), .Z(n179) );
  AND U169 ( .A(n80), .B(n184), .Z(n185) );
  XNOR U170 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n186), .Z(n184) );
  IV U171 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .Z(n186) );
  XOR U172 ( .A(n187), .B(n188), .Z(o[34]) );
  XOR U173 ( .A(n189), .B(n190), .Z(o[33]) );
  XOR U174 ( .A(n191), .B(n192), .Z(o[32]) );
  XOR U175 ( .A(n9), .B(n193), .Z(o[31]) );
  AND U176 ( .A(n58), .B(n194), .Z(n9) );
  XOR U177 ( .A(n10), .B(n193), .Z(n194) );
  XOR U178 ( .A(n195), .B(n196), .Z(n193) );
  AND U179 ( .A(n70), .B(n197), .Z(n196) );
  XOR U180 ( .A(n198), .B(n199), .Z(n10) );
  AND U181 ( .A(n62), .B(n200), .Z(n199) );
  XOR U182 ( .A(p_input[31]), .B(n198), .Z(n200) );
  XNOR U183 ( .A(n201), .B(n202), .Z(n198) );
  AND U184 ( .A(n66), .B(n197), .Z(n202) );
  XNOR U185 ( .A(n201), .B(n195), .Z(n197) );
  XNOR U186 ( .A(n203), .B(n204), .Z(n195) );
  AND U187 ( .A(n80), .B(n205), .Z(n204) );
  XNOR U188 ( .A(n206), .B(n207), .Z(n201) );
  AND U189 ( .A(n74), .B(n208), .Z(n207) );
  XOR U190 ( .A(p_input[63]), .B(n206), .Z(n208) );
  XOR U191 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .B(n209), .Z(
        n206) );
  AND U192 ( .A(n77), .B(n205), .Z(n209) );
  XNOR U193 ( .A(\knn_comb_/min_val_out[0][31] ), .B(n210), .Z(n205) );
  IV U194 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .Z(n210) );
  XOR U195 ( .A(n11), .B(n211), .Z(o[30]) );
  AND U196 ( .A(n58), .B(n212), .Z(n11) );
  XOR U197 ( .A(n12), .B(n211), .Z(n212) );
  XOR U198 ( .A(n213), .B(n214), .Z(n211) );
  AND U199 ( .A(n70), .B(n215), .Z(n214) );
  XOR U200 ( .A(n216), .B(n217), .Z(n12) );
  AND U201 ( .A(n62), .B(n218), .Z(n217) );
  XOR U202 ( .A(p_input[30]), .B(n216), .Z(n218) );
  XNOR U203 ( .A(n219), .B(n220), .Z(n216) );
  AND U204 ( .A(n66), .B(n215), .Z(n220) );
  XNOR U205 ( .A(n219), .B(n213), .Z(n215) );
  XNOR U206 ( .A(n221), .B(n222), .Z(n213) );
  AND U207 ( .A(n80), .B(n223), .Z(n222) );
  XNOR U208 ( .A(n224), .B(n225), .Z(n219) );
  AND U209 ( .A(n74), .B(n226), .Z(n225) );
  XOR U210 ( .A(p_input[62]), .B(n224), .Z(n226) );
  XOR U211 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .B(n227), .Z(
        n224) );
  AND U212 ( .A(n77), .B(n223), .Z(n227) );
  XNOR U213 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n228), .Z(n223) );
  XOR U214 ( .A(n187), .B(n229), .Z(o[2]) );
  AND U215 ( .A(n58), .B(n230), .Z(n187) );
  XOR U216 ( .A(n188), .B(n229), .Z(n230) );
  XOR U217 ( .A(n231), .B(n232), .Z(n229) );
  AND U218 ( .A(n70), .B(n233), .Z(n232) );
  XOR U219 ( .A(n234), .B(n235), .Z(n188) );
  AND U220 ( .A(n62), .B(n236), .Z(n235) );
  XOR U221 ( .A(p_input[2]), .B(n234), .Z(n236) );
  XNOR U222 ( .A(n237), .B(n238), .Z(n234) );
  AND U223 ( .A(n66), .B(n233), .Z(n238) );
  XNOR U224 ( .A(n237), .B(n231), .Z(n233) );
  XOR U225 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n239), .Z(n231) );
  AND U226 ( .A(n80), .B(n240), .Z(n239) );
  XNOR U227 ( .A(n241), .B(n242), .Z(n237) );
  AND U228 ( .A(n74), .B(n243), .Z(n242) );
  XOR U229 ( .A(p_input[34]), .B(n241), .Z(n243) );
  XOR U230 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .B(n244), .Z(
        n241) );
  AND U231 ( .A(n77), .B(n240), .Z(n244) );
  XNOR U232 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n245), .Z(n240) );
  XOR U233 ( .A(n13), .B(n246), .Z(o[29]) );
  AND U234 ( .A(n58), .B(n247), .Z(n13) );
  XOR U235 ( .A(n14), .B(n246), .Z(n247) );
  XOR U236 ( .A(n248), .B(n249), .Z(n246) );
  AND U237 ( .A(n70), .B(n250), .Z(n249) );
  XOR U238 ( .A(n251), .B(n252), .Z(n14) );
  AND U239 ( .A(n62), .B(n253), .Z(n252) );
  XOR U240 ( .A(p_input[29]), .B(n251), .Z(n253) );
  XNOR U241 ( .A(n254), .B(n255), .Z(n251) );
  AND U242 ( .A(n66), .B(n250), .Z(n255) );
  XNOR U243 ( .A(n254), .B(n248), .Z(n250) );
  XOR U244 ( .A(\knn_comb_/min_val_out[0][29] ), .B(n256), .Z(n248) );
  AND U245 ( .A(n80), .B(n257), .Z(n256) );
  XNOR U246 ( .A(n258), .B(n259), .Z(n254) );
  AND U247 ( .A(n74), .B(n260), .Z(n259) );
  XOR U248 ( .A(p_input[61]), .B(n258), .Z(n260) );
  XOR U249 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .B(n261), .Z(
        n258) );
  AND U250 ( .A(n77), .B(n257), .Z(n261) );
  XNOR U251 ( .A(\knn_comb_/min_val_out[0][29] ), .B(n262), .Z(n257) );
  XOR U252 ( .A(n15), .B(n263), .Z(o[28]) );
  AND U253 ( .A(n58), .B(n264), .Z(n15) );
  XOR U254 ( .A(n16), .B(n263), .Z(n264) );
  XOR U255 ( .A(n265), .B(n266), .Z(n263) );
  AND U256 ( .A(n70), .B(n267), .Z(n266) );
  XOR U257 ( .A(n268), .B(n269), .Z(n16) );
  AND U258 ( .A(n62), .B(n270), .Z(n269) );
  XOR U259 ( .A(p_input[28]), .B(n268), .Z(n270) );
  XNOR U260 ( .A(n271), .B(n272), .Z(n268) );
  AND U261 ( .A(n66), .B(n267), .Z(n272) );
  XNOR U262 ( .A(n271), .B(n265), .Z(n267) );
  XOR U263 ( .A(\knn_comb_/min_val_out[0][28] ), .B(n273), .Z(n265) );
  AND U264 ( .A(n80), .B(n274), .Z(n273) );
  XNOR U265 ( .A(n275), .B(n276), .Z(n271) );
  AND U266 ( .A(n74), .B(n277), .Z(n276) );
  XOR U267 ( .A(p_input[60]), .B(n275), .Z(n277) );
  XOR U268 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .B(n278), .Z(
        n275) );
  AND U269 ( .A(n77), .B(n274), .Z(n278) );
  XNOR U270 ( .A(\knn_comb_/min_val_out[0][28] ), .B(n279), .Z(n274) );
  XOR U271 ( .A(n19), .B(n280), .Z(o[27]) );
  AND U272 ( .A(n58), .B(n281), .Z(n19) );
  XOR U273 ( .A(n20), .B(n280), .Z(n281) );
  XOR U274 ( .A(n282), .B(n283), .Z(n280) );
  AND U275 ( .A(n70), .B(n284), .Z(n283) );
  XOR U276 ( .A(n285), .B(n286), .Z(n20) );
  AND U277 ( .A(n62), .B(n287), .Z(n286) );
  XOR U278 ( .A(p_input[27]), .B(n285), .Z(n287) );
  XNOR U279 ( .A(n288), .B(n289), .Z(n285) );
  AND U280 ( .A(n66), .B(n284), .Z(n289) );
  XNOR U281 ( .A(n288), .B(n282), .Z(n284) );
  XNOR U282 ( .A(n290), .B(n291), .Z(n282) );
  AND U283 ( .A(n80), .B(n292), .Z(n291) );
  XNOR U284 ( .A(n293), .B(n294), .Z(n288) );
  AND U285 ( .A(n74), .B(n295), .Z(n294) );
  XOR U286 ( .A(p_input[59]), .B(n293), .Z(n295) );
  XOR U287 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .B(n296), .Z(
        n293) );
  AND U288 ( .A(n77), .B(n292), .Z(n296) );
  XNOR U289 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n297), .Z(n292) );
  XOR U290 ( .A(n21), .B(n298), .Z(o[26]) );
  AND U291 ( .A(n58), .B(n299), .Z(n21) );
  XOR U292 ( .A(n22), .B(n298), .Z(n299) );
  XOR U293 ( .A(n300), .B(n301), .Z(n298) );
  AND U294 ( .A(n70), .B(n302), .Z(n301) );
  XOR U295 ( .A(n303), .B(n304), .Z(n22) );
  AND U296 ( .A(n62), .B(n305), .Z(n304) );
  XOR U297 ( .A(p_input[26]), .B(n303), .Z(n305) );
  XNOR U298 ( .A(n306), .B(n307), .Z(n303) );
  AND U299 ( .A(n66), .B(n302), .Z(n307) );
  XNOR U300 ( .A(n306), .B(n300), .Z(n302) );
  XOR U301 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n308), .Z(n300) );
  AND U302 ( .A(n80), .B(n309), .Z(n308) );
  XNOR U303 ( .A(n310), .B(n311), .Z(n306) );
  AND U304 ( .A(n74), .B(n312), .Z(n311) );
  XOR U305 ( .A(p_input[58]), .B(n310), .Z(n312) );
  XOR U306 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .B(n313), .Z(
        n310) );
  AND U307 ( .A(n77), .B(n309), .Z(n313) );
  XNOR U308 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n314), .Z(n309) );
  XOR U309 ( .A(n23), .B(n315), .Z(o[25]) );
  AND U310 ( .A(n58), .B(n316), .Z(n23) );
  XOR U311 ( .A(n24), .B(n315), .Z(n316) );
  XOR U312 ( .A(n317), .B(n318), .Z(n315) );
  AND U313 ( .A(n70), .B(n319), .Z(n318) );
  XOR U314 ( .A(n320), .B(n321), .Z(n24) );
  AND U315 ( .A(n62), .B(n322), .Z(n321) );
  XOR U316 ( .A(p_input[25]), .B(n320), .Z(n322) );
  XNOR U317 ( .A(n323), .B(n324), .Z(n320) );
  AND U318 ( .A(n66), .B(n319), .Z(n324) );
  XNOR U319 ( .A(n323), .B(n317), .Z(n319) );
  XOR U320 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n325), .Z(n317) );
  AND U321 ( .A(n80), .B(n326), .Z(n325) );
  XNOR U322 ( .A(n327), .B(n328), .Z(n323) );
  AND U323 ( .A(n74), .B(n329), .Z(n328) );
  XOR U324 ( .A(p_input[57]), .B(n327), .Z(n329) );
  XOR U325 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .B(n330), .Z(
        n327) );
  AND U326 ( .A(n77), .B(n326), .Z(n330) );
  XNOR U327 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n331), .Z(n326) );
  IV U328 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .Z(n331) );
  XOR U329 ( .A(n25), .B(n332), .Z(o[24]) );
  AND U330 ( .A(n58), .B(n333), .Z(n25) );
  XOR U331 ( .A(n26), .B(n332), .Z(n333) );
  XOR U332 ( .A(n334), .B(n335), .Z(n332) );
  AND U333 ( .A(n70), .B(n336), .Z(n335) );
  XOR U334 ( .A(n337), .B(n338), .Z(n26) );
  AND U335 ( .A(n62), .B(n339), .Z(n338) );
  XOR U336 ( .A(p_input[24]), .B(n337), .Z(n339) );
  XNOR U337 ( .A(n340), .B(n341), .Z(n337) );
  AND U338 ( .A(n66), .B(n336), .Z(n341) );
  XNOR U339 ( .A(n340), .B(n334), .Z(n336) );
  XOR U340 ( .A(\knn_comb_/min_val_out[0][24] ), .B(n342), .Z(n334) );
  AND U341 ( .A(n80), .B(n343), .Z(n342) );
  XNOR U342 ( .A(n344), .B(n345), .Z(n340) );
  AND U343 ( .A(n74), .B(n346), .Z(n345) );
  XOR U344 ( .A(p_input[56]), .B(n344), .Z(n346) );
  XOR U345 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .B(n347), .Z(
        n344) );
  AND U346 ( .A(n77), .B(n343), .Z(n347) );
  XNOR U347 ( .A(\knn_comb_/min_val_out[0][24] ), .B(n348), .Z(n343) );
  IV U348 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .Z(n348) );
  XOR U349 ( .A(n27), .B(n349), .Z(o[23]) );
  AND U350 ( .A(n58), .B(n350), .Z(n27) );
  XOR U351 ( .A(n28), .B(n349), .Z(n350) );
  XOR U352 ( .A(n351), .B(n352), .Z(n349) );
  AND U353 ( .A(n70), .B(n353), .Z(n352) );
  XOR U354 ( .A(n354), .B(n355), .Z(n28) );
  AND U355 ( .A(n62), .B(n356), .Z(n355) );
  XOR U356 ( .A(p_input[23]), .B(n354), .Z(n356) );
  XNOR U357 ( .A(n357), .B(n358), .Z(n354) );
  AND U358 ( .A(n66), .B(n353), .Z(n358) );
  XNOR U359 ( .A(n357), .B(n351), .Z(n353) );
  XNOR U360 ( .A(n359), .B(n360), .Z(n351) );
  AND U361 ( .A(n80), .B(n361), .Z(n360) );
  XNOR U362 ( .A(n362), .B(n363), .Z(n357) );
  AND U363 ( .A(n74), .B(n364), .Z(n363) );
  XOR U364 ( .A(p_input[55]), .B(n362), .Z(n364) );
  XOR U365 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .B(n365), .Z(
        n362) );
  AND U366 ( .A(n77), .B(n361), .Z(n365) );
  XNOR U367 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n366), .Z(n361) );
  XOR U368 ( .A(n29), .B(n367), .Z(o[22]) );
  AND U369 ( .A(n58), .B(n368), .Z(n29) );
  XOR U370 ( .A(n30), .B(n367), .Z(n368) );
  XOR U371 ( .A(n369), .B(n370), .Z(n367) );
  AND U372 ( .A(n70), .B(n371), .Z(n370) );
  XOR U373 ( .A(n372), .B(n373), .Z(n30) );
  AND U374 ( .A(n62), .B(n374), .Z(n373) );
  XOR U375 ( .A(p_input[22]), .B(n372), .Z(n374) );
  XNOR U376 ( .A(n375), .B(n376), .Z(n372) );
  AND U377 ( .A(n66), .B(n371), .Z(n376) );
  XNOR U378 ( .A(n375), .B(n369), .Z(n371) );
  XOR U379 ( .A(\knn_comb_/min_val_out[0][22] ), .B(n377), .Z(n369) );
  AND U380 ( .A(n80), .B(n378), .Z(n377) );
  XNOR U381 ( .A(n379), .B(n380), .Z(n375) );
  AND U382 ( .A(n74), .B(n381), .Z(n380) );
  XOR U383 ( .A(p_input[54]), .B(n379), .Z(n381) );
  XOR U384 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .B(n382), .Z(
        n379) );
  AND U385 ( .A(n77), .B(n378), .Z(n382) );
  XNOR U386 ( .A(\knn_comb_/min_val_out[0][22] ), .B(n383), .Z(n378) );
  XOR U387 ( .A(n31), .B(n384), .Z(o[21]) );
  AND U388 ( .A(n58), .B(n385), .Z(n31) );
  XOR U389 ( .A(n32), .B(n384), .Z(n385) );
  XOR U390 ( .A(n386), .B(n387), .Z(n384) );
  AND U391 ( .A(n70), .B(n388), .Z(n387) );
  XOR U392 ( .A(n389), .B(n390), .Z(n32) );
  AND U393 ( .A(n62), .B(n391), .Z(n390) );
  XOR U394 ( .A(p_input[21]), .B(n389), .Z(n391) );
  XNOR U395 ( .A(n392), .B(n393), .Z(n389) );
  AND U396 ( .A(n66), .B(n388), .Z(n393) );
  XNOR U397 ( .A(n392), .B(n386), .Z(n388) );
  XOR U398 ( .A(\knn_comb_/min_val_out[0][21] ), .B(n394), .Z(n386) );
  AND U399 ( .A(n80), .B(n395), .Z(n394) );
  XNOR U400 ( .A(n396), .B(n397), .Z(n392) );
  AND U401 ( .A(n74), .B(n398), .Z(n397) );
  XOR U402 ( .A(p_input[53]), .B(n396), .Z(n398) );
  XOR U403 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .B(n399), .Z(
        n396) );
  AND U404 ( .A(n77), .B(n395), .Z(n399) );
  XNOR U405 ( .A(\knn_comb_/min_val_out[0][21] ), .B(n400), .Z(n395) );
  XOR U406 ( .A(n33), .B(n401), .Z(o[20]) );
  AND U407 ( .A(n58), .B(n402), .Z(n33) );
  XOR U408 ( .A(n34), .B(n401), .Z(n402) );
  XOR U409 ( .A(n403), .B(n404), .Z(n401) );
  AND U410 ( .A(n70), .B(n405), .Z(n404) );
  XOR U411 ( .A(n406), .B(n407), .Z(n34) );
  AND U412 ( .A(n62), .B(n408), .Z(n407) );
  XOR U413 ( .A(p_input[20]), .B(n406), .Z(n408) );
  XNOR U414 ( .A(n409), .B(n410), .Z(n406) );
  AND U415 ( .A(n66), .B(n405), .Z(n410) );
  XNOR U416 ( .A(n409), .B(n403), .Z(n405) );
  XNOR U417 ( .A(n411), .B(n412), .Z(n403) );
  AND U418 ( .A(n80), .B(n413), .Z(n412) );
  XNOR U419 ( .A(n414), .B(n415), .Z(n409) );
  AND U420 ( .A(n74), .B(n416), .Z(n415) );
  XOR U421 ( .A(p_input[52]), .B(n414), .Z(n416) );
  XOR U422 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .B(n417), .Z(
        n414) );
  AND U423 ( .A(n77), .B(n413), .Z(n417) );
  XNOR U424 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n418), .Z(n413) );
  XOR U425 ( .A(n189), .B(n419), .Z(o[1]) );
  AND U426 ( .A(n58), .B(n420), .Z(n189) );
  XOR U427 ( .A(n190), .B(n419), .Z(n420) );
  XOR U428 ( .A(n421), .B(n422), .Z(n419) );
  AND U429 ( .A(n70), .B(n423), .Z(n422) );
  XOR U430 ( .A(n424), .B(n425), .Z(n190) );
  AND U431 ( .A(n62), .B(n426), .Z(n425) );
  XOR U432 ( .A(p_input[1]), .B(n424), .Z(n426) );
  XNOR U433 ( .A(n427), .B(n428), .Z(n424) );
  AND U434 ( .A(n66), .B(n423), .Z(n428) );
  XNOR U435 ( .A(n427), .B(n421), .Z(n423) );
  XOR U436 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n429), .Z(n421) );
  AND U437 ( .A(n80), .B(n430), .Z(n429) );
  XNOR U438 ( .A(n431), .B(n432), .Z(n427) );
  AND U439 ( .A(n74), .B(n433), .Z(n432) );
  XOR U440 ( .A(p_input[33]), .B(n431), .Z(n433) );
  XOR U441 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(n434), .Z(
        n431) );
  AND U442 ( .A(n77), .B(n430), .Z(n434) );
  XNOR U443 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n435), .Z(n430) );
  XOR U444 ( .A(n35), .B(n436), .Z(o[19]) );
  AND U445 ( .A(n58), .B(n437), .Z(n35) );
  XOR U446 ( .A(n36), .B(n436), .Z(n437) );
  XOR U447 ( .A(n438), .B(n439), .Z(n436) );
  AND U448 ( .A(n70), .B(n440), .Z(n439) );
  XOR U449 ( .A(n441), .B(n442), .Z(n36) );
  AND U450 ( .A(n62), .B(n443), .Z(n442) );
  XOR U451 ( .A(p_input[19]), .B(n441), .Z(n443) );
  XNOR U452 ( .A(n444), .B(n445), .Z(n441) );
  AND U453 ( .A(n66), .B(n440), .Z(n445) );
  XNOR U454 ( .A(n444), .B(n438), .Z(n440) );
  XOR U455 ( .A(\knn_comb_/min_val_out[0][19] ), .B(n446), .Z(n438) );
  AND U456 ( .A(n80), .B(n447), .Z(n446) );
  XNOR U457 ( .A(n448), .B(n449), .Z(n444) );
  AND U458 ( .A(n74), .B(n450), .Z(n449) );
  XOR U459 ( .A(p_input[51]), .B(n448), .Z(n450) );
  XOR U460 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .B(n451), .Z(
        n448) );
  AND U461 ( .A(n77), .B(n447), .Z(n451) );
  XNOR U462 ( .A(\knn_comb_/min_val_out[0][19] ), .B(n452), .Z(n447) );
  XOR U463 ( .A(n37), .B(n453), .Z(o[18]) );
  AND U464 ( .A(n58), .B(n454), .Z(n37) );
  XOR U465 ( .A(n38), .B(n453), .Z(n454) );
  XOR U466 ( .A(n455), .B(n456), .Z(n453) );
  AND U467 ( .A(n70), .B(n457), .Z(n456) );
  XOR U468 ( .A(n458), .B(n459), .Z(n38) );
  AND U469 ( .A(n62), .B(n460), .Z(n459) );
  XOR U470 ( .A(p_input[18]), .B(n458), .Z(n460) );
  XNOR U471 ( .A(n461), .B(n462), .Z(n458) );
  AND U472 ( .A(n66), .B(n457), .Z(n462) );
  XNOR U473 ( .A(n461), .B(n455), .Z(n457) );
  XOR U474 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n463), .Z(n455) );
  AND U475 ( .A(n80), .B(n464), .Z(n463) );
  XNOR U476 ( .A(n465), .B(n466), .Z(n461) );
  AND U477 ( .A(n74), .B(n467), .Z(n466) );
  XOR U478 ( .A(p_input[50]), .B(n465), .Z(n467) );
  XOR U479 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .B(n468), .Z(
        n465) );
  AND U480 ( .A(n77), .B(n464), .Z(n468) );
  XNOR U481 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n469), .Z(n464) );
  IV U482 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .Z(n469) );
  XOR U483 ( .A(n41), .B(n470), .Z(o[17]) );
  AND U484 ( .A(n58), .B(n471), .Z(n41) );
  XOR U485 ( .A(n42), .B(n470), .Z(n471) );
  XOR U486 ( .A(n472), .B(n473), .Z(n470) );
  AND U487 ( .A(n70), .B(n474), .Z(n473) );
  XOR U488 ( .A(n475), .B(n476), .Z(n42) );
  AND U489 ( .A(n62), .B(n477), .Z(n476) );
  XOR U490 ( .A(p_input[17]), .B(n475), .Z(n477) );
  XNOR U491 ( .A(n478), .B(n479), .Z(n475) );
  AND U492 ( .A(n66), .B(n474), .Z(n479) );
  XNOR U493 ( .A(n478), .B(n472), .Z(n474) );
  XOR U494 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n480), .Z(n472) );
  AND U495 ( .A(n80), .B(n481), .Z(n480) );
  XNOR U496 ( .A(n482), .B(n483), .Z(n478) );
  AND U497 ( .A(n74), .B(n484), .Z(n483) );
  XOR U498 ( .A(p_input[49]), .B(n482), .Z(n484) );
  XOR U499 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .B(n485), .Z(
        n482) );
  AND U500 ( .A(n77), .B(n481), .Z(n485) );
  XNOR U501 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n486), .Z(n481) );
  XOR U502 ( .A(n43), .B(n487), .Z(o[16]) );
  AND U503 ( .A(n58), .B(n488), .Z(n43) );
  XOR U504 ( .A(n44), .B(n487), .Z(n488) );
  XOR U505 ( .A(n489), .B(n490), .Z(n487) );
  AND U506 ( .A(n70), .B(n491), .Z(n490) );
  XOR U507 ( .A(n492), .B(n493), .Z(n44) );
  AND U508 ( .A(n62), .B(n494), .Z(n493) );
  XOR U509 ( .A(p_input[16]), .B(n492), .Z(n494) );
  XNOR U510 ( .A(n495), .B(n496), .Z(n492) );
  AND U511 ( .A(n66), .B(n491), .Z(n496) );
  XNOR U512 ( .A(n495), .B(n489), .Z(n491) );
  XNOR U513 ( .A(n497), .B(n498), .Z(n489) );
  AND U514 ( .A(n80), .B(n499), .Z(n498) );
  XNOR U515 ( .A(n500), .B(n501), .Z(n495) );
  AND U516 ( .A(n74), .B(n502), .Z(n501) );
  XOR U517 ( .A(p_input[48]), .B(n500), .Z(n502) );
  XOR U518 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .B(n503), .Z(
        n500) );
  AND U519 ( .A(n77), .B(n499), .Z(n503) );
  XNOR U520 ( .A(\knn_comb_/min_val_out[0][16] ), .B(n504), .Z(n499) );
  IV U521 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .Z(n504) );
  XOR U522 ( .A(n45), .B(n505), .Z(o[15]) );
  AND U523 ( .A(n58), .B(n506), .Z(n45) );
  XOR U524 ( .A(n46), .B(n505), .Z(n506) );
  XOR U525 ( .A(n507), .B(n508), .Z(n505) );
  AND U526 ( .A(n70), .B(n509), .Z(n508) );
  XOR U527 ( .A(n510), .B(n511), .Z(n46) );
  AND U528 ( .A(n62), .B(n512), .Z(n511) );
  XOR U529 ( .A(p_input[15]), .B(n510), .Z(n512) );
  XNOR U530 ( .A(n513), .B(n514), .Z(n510) );
  AND U531 ( .A(n66), .B(n509), .Z(n514) );
  XNOR U532 ( .A(n513), .B(n507), .Z(n509) );
  XNOR U533 ( .A(n515), .B(n516), .Z(n507) );
  AND U534 ( .A(n80), .B(n517), .Z(n516) );
  XNOR U535 ( .A(n518), .B(n519), .Z(n513) );
  AND U536 ( .A(n74), .B(n520), .Z(n519) );
  XOR U537 ( .A(p_input[47]), .B(n518), .Z(n520) );
  XOR U538 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(n521), .Z(
        n518) );
  AND U539 ( .A(n77), .B(n517), .Z(n521) );
  XNOR U540 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n522), .Z(n517) );
  XOR U541 ( .A(n47), .B(n523), .Z(o[14]) );
  AND U542 ( .A(n58), .B(n524), .Z(n47) );
  XOR U543 ( .A(n48), .B(n523), .Z(n524) );
  XOR U544 ( .A(n525), .B(n526), .Z(n523) );
  AND U545 ( .A(n70), .B(n527), .Z(n526) );
  XOR U546 ( .A(n528), .B(n529), .Z(n48) );
  AND U547 ( .A(n62), .B(n530), .Z(n529) );
  XOR U548 ( .A(p_input[14]), .B(n528), .Z(n530) );
  XNOR U549 ( .A(n531), .B(n532), .Z(n528) );
  AND U550 ( .A(n66), .B(n527), .Z(n532) );
  XNOR U551 ( .A(n531), .B(n525), .Z(n527) );
  XOR U552 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n533), .Z(n525) );
  AND U553 ( .A(n80), .B(n534), .Z(n533) );
  XNOR U554 ( .A(n535), .B(n536), .Z(n531) );
  AND U555 ( .A(n74), .B(n537), .Z(n536) );
  XOR U556 ( .A(p_input[46]), .B(n535), .Z(n537) );
  XOR U557 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(n538), .Z(
        n535) );
  AND U558 ( .A(n77), .B(n534), .Z(n538) );
  XNOR U559 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n539), .Z(n534) );
  XOR U560 ( .A(n49), .B(n540), .Z(o[13]) );
  AND U561 ( .A(n58), .B(n541), .Z(n49) );
  XOR U562 ( .A(n50), .B(n540), .Z(n541) );
  XOR U563 ( .A(n542), .B(n543), .Z(n540) );
  AND U564 ( .A(n70), .B(n544), .Z(n543) );
  XOR U565 ( .A(n545), .B(n546), .Z(n50) );
  AND U566 ( .A(n62), .B(n547), .Z(n546) );
  XOR U567 ( .A(p_input[13]), .B(n545), .Z(n547) );
  XNOR U568 ( .A(n548), .B(n549), .Z(n545) );
  AND U569 ( .A(n66), .B(n544), .Z(n549) );
  XNOR U570 ( .A(n548), .B(n542), .Z(n544) );
  XOR U571 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n550), .Z(n542) );
  AND U572 ( .A(n80), .B(n551), .Z(n550) );
  XNOR U573 ( .A(n552), .B(n553), .Z(n548) );
  AND U574 ( .A(n74), .B(n554), .Z(n553) );
  XOR U575 ( .A(p_input[45]), .B(n552), .Z(n554) );
  XOR U576 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(n555), .Z(
        n552) );
  AND U577 ( .A(n77), .B(n551), .Z(n555) );
  XNOR U578 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n556), .Z(n551) );
  IV U579 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n556) );
  XOR U580 ( .A(n51), .B(n557), .Z(o[12]) );
  AND U581 ( .A(n58), .B(n558), .Z(n51) );
  XOR U582 ( .A(n52), .B(n557), .Z(n558) );
  XOR U583 ( .A(n559), .B(n560), .Z(n557) );
  AND U584 ( .A(n70), .B(n561), .Z(n560) );
  XOR U585 ( .A(n562), .B(n563), .Z(n52) );
  AND U586 ( .A(n62), .B(n564), .Z(n563) );
  XOR U587 ( .A(p_input[12]), .B(n562), .Z(n564) );
  XNOR U588 ( .A(n565), .B(n566), .Z(n562) );
  AND U589 ( .A(n66), .B(n561), .Z(n566) );
  XNOR U590 ( .A(n565), .B(n559), .Z(n561) );
  XNOR U591 ( .A(n567), .B(n568), .Z(n559) );
  AND U592 ( .A(n80), .B(n569), .Z(n568) );
  XNOR U593 ( .A(n570), .B(n571), .Z(n565) );
  AND U594 ( .A(n74), .B(n572), .Z(n571) );
  XOR U595 ( .A(p_input[44]), .B(n570), .Z(n572) );
  XOR U596 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(n573), .Z(
        n570) );
  AND U597 ( .A(n77), .B(n569), .Z(n573) );
  XNOR U598 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n574), .Z(n569) );
  XOR U599 ( .A(n53), .B(n575), .Z(o[11]) );
  AND U600 ( .A(n58), .B(n576), .Z(n53) );
  XOR U601 ( .A(n54), .B(n575), .Z(n576) );
  XOR U602 ( .A(n577), .B(n578), .Z(n575) );
  AND U603 ( .A(n70), .B(n579), .Z(n578) );
  XOR U604 ( .A(n580), .B(n581), .Z(n54) );
  AND U605 ( .A(n62), .B(n582), .Z(n581) );
  XOR U606 ( .A(p_input[11]), .B(n580), .Z(n582) );
  XNOR U607 ( .A(n583), .B(n584), .Z(n580) );
  AND U608 ( .A(n66), .B(n579), .Z(n584) );
  XNOR U609 ( .A(n583), .B(n577), .Z(n579) );
  XOR U610 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n585), .Z(n577) );
  AND U611 ( .A(n80), .B(n586), .Z(n585) );
  XNOR U612 ( .A(n587), .B(n588), .Z(n583) );
  AND U613 ( .A(n74), .B(n589), .Z(n588) );
  XOR U614 ( .A(p_input[43]), .B(n587), .Z(n589) );
  XOR U615 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n590), .Z(
        n587) );
  AND U616 ( .A(n77), .B(n586), .Z(n590) );
  XNOR U617 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n591), .Z(n586) );
  IV U618 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n591) );
  XOR U619 ( .A(n55), .B(n592), .Z(o[10]) );
  AND U620 ( .A(n58), .B(n593), .Z(n55) );
  XOR U621 ( .A(n56), .B(n592), .Z(n593) );
  XOR U622 ( .A(n594), .B(n595), .Z(n592) );
  AND U623 ( .A(n70), .B(n596), .Z(n595) );
  XOR U624 ( .A(n597), .B(n598), .Z(n56) );
  AND U625 ( .A(n62), .B(n599), .Z(n598) );
  XOR U626 ( .A(p_input[10]), .B(n597), .Z(n599) );
  XNOR U627 ( .A(n600), .B(n601), .Z(n597) );
  AND U628 ( .A(n66), .B(n596), .Z(n601) );
  XNOR U629 ( .A(n600), .B(n594), .Z(n596) );
  XOR U630 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n602), .Z(n594) );
  AND U631 ( .A(n80), .B(n603), .Z(n602) );
  XNOR U632 ( .A(n604), .B(n605), .Z(n600) );
  AND U633 ( .A(n74), .B(n606), .Z(n605) );
  XOR U634 ( .A(p_input[42]), .B(n604), .Z(n606) );
  XOR U635 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(n607), .Z(
        n604) );
  AND U636 ( .A(n77), .B(n603), .Z(n607) );
  XNOR U637 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n608), .Z(n603) );
  IV U638 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n608) );
  XOR U639 ( .A(n191), .B(n609), .Z(o[0]) );
  AND U640 ( .A(n58), .B(n610), .Z(n191) );
  XOR U641 ( .A(n192), .B(n609), .Z(n610) );
  XOR U642 ( .A(n611), .B(n612), .Z(n609) );
  AND U643 ( .A(n70), .B(n613), .Z(n612) );
  XOR U644 ( .A(n614), .B(n615), .Z(n192) );
  AND U645 ( .A(n62), .B(n616), .Z(n615) );
  XOR U646 ( .A(p_input[0]), .B(n614), .Z(n616) );
  XNOR U647 ( .A(n617), .B(n618), .Z(n614) );
  AND U648 ( .A(n66), .B(n613), .Z(n618) );
  XNOR U649 ( .A(n617), .B(n611), .Z(n613) );
  XOR U650 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n619), .Z(n611) );
  AND U651 ( .A(n80), .B(n620), .Z(n619) );
  XNOR U652 ( .A(n621), .B(n622), .Z(n617) );
  AND U653 ( .A(n74), .B(n623), .Z(n622) );
  XOR U654 ( .A(p_input[32]), .B(n621), .Z(n623) );
  XOR U655 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(n624), .Z(
        n621) );
  AND U656 ( .A(n77), .B(n620), .Z(n624) );
  XNOR U657 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n625), .Z(n620) );
  XNOR U658 ( .A(n626), .B(n627), .Z(n58) );
  NOR U659 ( .A(n628), .B(n629), .Z(n627) );
  XOR U660 ( .A(n630), .B(n626), .Z(n629) );
  AND U661 ( .A(n631), .B(n632), .Z(n630) );
  NOR U662 ( .A(n626), .B(n633), .Z(n628) );
  AND U663 ( .A(n634), .B(n635), .Z(n633) );
  XOR U664 ( .A(n636), .B(n637), .Z(n626) );
  AND U665 ( .A(n638), .B(n639), .Z(n637) );
  XNOR U666 ( .A(n636), .B(n640), .Z(n639) );
  XOR U667 ( .A(n641), .B(n642), .Z(n640) );
  AND U668 ( .A(n62), .B(n643), .Z(n642) );
  XOR U669 ( .A(n641), .B(n644), .Z(n643) );
  XNOR U670 ( .A(n636), .B(n645), .Z(n638) );
  XOR U671 ( .A(n646), .B(n647), .Z(n645) );
  AND U672 ( .A(n70), .B(n648), .Z(n647) );
  XOR U673 ( .A(n649), .B(n650), .Z(n636) );
  AND U674 ( .A(n651), .B(n652), .Z(n650) );
  XOR U675 ( .A(n653), .B(n649), .Z(n652) );
  XOR U676 ( .A(n654), .B(n655), .Z(n653) );
  AND U677 ( .A(n62), .B(n656), .Z(n655) );
  XNOR U678 ( .A(n657), .B(n654), .Z(n656) );
  XNOR U679 ( .A(n649), .B(n658), .Z(n651) );
  XNOR U680 ( .A(n659), .B(n660), .Z(n658) );
  AND U681 ( .A(n70), .B(n661), .Z(n660) );
  XOR U682 ( .A(n662), .B(n663), .Z(n649) );
  AND U683 ( .A(n664), .B(n665), .Z(n663) );
  XOR U684 ( .A(n666), .B(n662), .Z(n665) );
  XOR U685 ( .A(n667), .B(n668), .Z(n666) );
  AND U686 ( .A(n62), .B(n669), .Z(n668) );
  XNOR U687 ( .A(n670), .B(n667), .Z(n669) );
  XNOR U688 ( .A(n662), .B(n671), .Z(n664) );
  XNOR U689 ( .A(n672), .B(n673), .Z(n671) );
  AND U690 ( .A(n70), .B(n674), .Z(n673) );
  XOR U691 ( .A(n675), .B(n676), .Z(n662) );
  AND U692 ( .A(n677), .B(n678), .Z(n676) );
  XOR U693 ( .A(n675), .B(n679), .Z(n678) );
  XOR U694 ( .A(n680), .B(n681), .Z(n679) );
  AND U695 ( .A(n62), .B(n682), .Z(n681) );
  XNOR U696 ( .A(n683), .B(n680), .Z(n682) );
  XNOR U697 ( .A(n684), .B(n675), .Z(n677) );
  XOR U698 ( .A(n685), .B(n686), .Z(n684) );
  AND U699 ( .A(n70), .B(n687), .Z(n686) );
  AND U700 ( .A(n688), .B(n689), .Z(n675) );
  XNOR U701 ( .A(n690), .B(n691), .Z(n689) );
  AND U702 ( .A(n62), .B(n692), .Z(n691) );
  XNOR U703 ( .A(n693), .B(n690), .Z(n692) );
  XNOR U704 ( .A(n694), .B(n695), .Z(n62) );
  NOR U705 ( .A(n696), .B(n697), .Z(n695) );
  XOR U706 ( .A(n694), .B(n634), .Z(n697) );
  IV U707 ( .A(n698), .Z(n634) );
  NOR U708 ( .A(n631), .B(n632), .Z(n698) );
  NOR U709 ( .A(n694), .B(n635), .Z(n696) );
  AND U710 ( .A(n644), .B(n699), .Z(n635) );
  XOR U711 ( .A(n700), .B(n701), .Z(n694) );
  AND U712 ( .A(n702), .B(n703), .Z(n701) );
  XOR U713 ( .A(n700), .B(n704), .Z(n703) );
  IV U714 ( .A(n644), .Z(n704) );
  XNOR U715 ( .A(n705), .B(n706), .Z(n644) );
  XOR U716 ( .A(n707), .B(n699), .Z(n706) );
  AND U717 ( .A(n657), .B(n708), .Z(n699) );
  AND U718 ( .A(n709), .B(n710), .Z(n707) );
  XOR U719 ( .A(n711), .B(n705), .Z(n709) );
  XOR U720 ( .A(n700), .B(n641), .Z(n702) );
  XNOR U721 ( .A(n712), .B(n713), .Z(n641) );
  AND U722 ( .A(n66), .B(n648), .Z(n713) );
  XOR U723 ( .A(n646), .B(n712), .Z(n648) );
  XOR U724 ( .A(n714), .B(n715), .Z(n700) );
  AND U725 ( .A(n716), .B(n717), .Z(n715) );
  XNOR U726 ( .A(n714), .B(n657), .Z(n717) );
  XOR U727 ( .A(n718), .B(n710), .Z(n657) );
  XNOR U728 ( .A(n719), .B(n705), .Z(n710) );
  XOR U729 ( .A(n720), .B(n721), .Z(n705) );
  AND U730 ( .A(n722), .B(n723), .Z(n721) );
  XOR U731 ( .A(n724), .B(n720), .Z(n722) );
  XNOR U732 ( .A(n725), .B(n726), .Z(n719) );
  AND U733 ( .A(n727), .B(n728), .Z(n726) );
  XOR U734 ( .A(n725), .B(n729), .Z(n727) );
  XNOR U735 ( .A(n711), .B(n708), .Z(n718) );
  AND U736 ( .A(n670), .B(n730), .Z(n708) );
  XOR U737 ( .A(n731), .B(n732), .Z(n711) );
  AND U738 ( .A(n733), .B(n734), .Z(n732) );
  XOR U739 ( .A(n731), .B(n735), .Z(n733) );
  XNOR U740 ( .A(n654), .B(n714), .Z(n716) );
  XNOR U741 ( .A(n736), .B(n737), .Z(n654) );
  AND U742 ( .A(n66), .B(n661), .Z(n737) );
  XNOR U743 ( .A(n736), .B(n738), .Z(n661) );
  XOR U744 ( .A(n739), .B(n740), .Z(n714) );
  AND U745 ( .A(n741), .B(n742), .Z(n740) );
  XOR U746 ( .A(n739), .B(n743), .Z(n742) );
  IV U747 ( .A(n670), .Z(n743) );
  XOR U748 ( .A(n744), .B(n723), .Z(n670) );
  XNOR U749 ( .A(n745), .B(n729), .Z(n723) );
  XOR U750 ( .A(n746), .B(n747), .Z(n729) );
  AND U751 ( .A(n748), .B(n749), .Z(n747) );
  XOR U752 ( .A(n746), .B(n750), .Z(n748) );
  XNOR U753 ( .A(n728), .B(n720), .Z(n745) );
  XOR U754 ( .A(n751), .B(n752), .Z(n720) );
  AND U755 ( .A(n753), .B(n754), .Z(n752) );
  XNOR U756 ( .A(n755), .B(n751), .Z(n753) );
  XNOR U757 ( .A(n756), .B(n725), .Z(n728) );
  XOR U758 ( .A(n757), .B(n758), .Z(n725) );
  AND U759 ( .A(n759), .B(n760), .Z(n758) );
  XOR U760 ( .A(n757), .B(n761), .Z(n759) );
  XNOR U761 ( .A(n762), .B(n763), .Z(n756) );
  AND U762 ( .A(n764), .B(n765), .Z(n763) );
  XNOR U763 ( .A(n762), .B(n766), .Z(n764) );
  XNOR U764 ( .A(n724), .B(n730), .Z(n744) );
  AND U765 ( .A(n683), .B(n767), .Z(n730) );
  XOR U766 ( .A(n735), .B(n734), .Z(n724) );
  XNOR U767 ( .A(n768), .B(n731), .Z(n734) );
  XOR U768 ( .A(n769), .B(n770), .Z(n731) );
  AND U769 ( .A(n771), .B(n772), .Z(n770) );
  XOR U770 ( .A(n769), .B(n773), .Z(n771) );
  XNOR U771 ( .A(n774), .B(n775), .Z(n768) );
  AND U772 ( .A(n776), .B(n777), .Z(n775) );
  XOR U773 ( .A(n774), .B(n778), .Z(n776) );
  XOR U774 ( .A(n779), .B(n780), .Z(n735) );
  AND U775 ( .A(n781), .B(n782), .Z(n780) );
  XOR U776 ( .A(n779), .B(n783), .Z(n781) );
  XNOR U777 ( .A(n667), .B(n739), .Z(n741) );
  XNOR U778 ( .A(n784), .B(n785), .Z(n667) );
  AND U779 ( .A(n66), .B(n674), .Z(n785) );
  XNOR U780 ( .A(n784), .B(n786), .Z(n674) );
  XOR U781 ( .A(n787), .B(n788), .Z(n739) );
  AND U782 ( .A(n789), .B(n790), .Z(n788) );
  XNOR U783 ( .A(n787), .B(n683), .Z(n790) );
  XOR U784 ( .A(n791), .B(n754), .Z(n683) );
  XNOR U785 ( .A(n792), .B(n761), .Z(n754) );
  XOR U786 ( .A(n750), .B(n749), .Z(n761) );
  XNOR U787 ( .A(n793), .B(n746), .Z(n749) );
  XOR U788 ( .A(n794), .B(n795), .Z(n746) );
  AND U789 ( .A(n796), .B(n797), .Z(n795) );
  XOR U790 ( .A(n794), .B(n798), .Z(n796) );
  XNOR U791 ( .A(n799), .B(n800), .Z(n793) );
  NOR U792 ( .A(n801), .B(n802), .Z(n800) );
  XNOR U793 ( .A(n799), .B(n803), .Z(n801) );
  XOR U794 ( .A(n804), .B(n805), .Z(n750) );
  NOR U795 ( .A(n806), .B(n807), .Z(n805) );
  XNOR U796 ( .A(n804), .B(n808), .Z(n806) );
  XNOR U797 ( .A(n760), .B(n751), .Z(n792) );
  XOR U798 ( .A(n809), .B(n810), .Z(n751) );
  NOR U799 ( .A(n811), .B(n812), .Z(n810) );
  XNOR U800 ( .A(n809), .B(n813), .Z(n811) );
  XOR U801 ( .A(n814), .B(n766), .Z(n760) );
  XNOR U802 ( .A(n815), .B(n816), .Z(n766) );
  NOR U803 ( .A(n817), .B(n818), .Z(n816) );
  XNOR U804 ( .A(n815), .B(n819), .Z(n817) );
  XNOR U805 ( .A(n765), .B(n757), .Z(n814) );
  XOR U806 ( .A(n820), .B(n821), .Z(n757) );
  AND U807 ( .A(n822), .B(n823), .Z(n821) );
  XOR U808 ( .A(n820), .B(n824), .Z(n822) );
  XNOR U809 ( .A(n825), .B(n762), .Z(n765) );
  XOR U810 ( .A(n826), .B(n827), .Z(n762) );
  AND U811 ( .A(n828), .B(n829), .Z(n827) );
  XOR U812 ( .A(n826), .B(n830), .Z(n828) );
  XNOR U813 ( .A(n831), .B(n832), .Z(n825) );
  NOR U814 ( .A(n833), .B(n834), .Z(n832) );
  XOR U815 ( .A(n831), .B(n835), .Z(n833) );
  XOR U816 ( .A(n755), .B(n767), .Z(n791) );
  NOR U817 ( .A(n693), .B(n836), .Z(n767) );
  XNOR U818 ( .A(n773), .B(n772), .Z(n755) );
  XNOR U819 ( .A(n837), .B(n778), .Z(n772) );
  XOR U820 ( .A(n838), .B(n839), .Z(n778) );
  NOR U821 ( .A(n840), .B(n841), .Z(n839) );
  XNOR U822 ( .A(n838), .B(n842), .Z(n840) );
  XNOR U823 ( .A(n777), .B(n769), .Z(n837) );
  XOR U824 ( .A(n843), .B(n844), .Z(n769) );
  AND U825 ( .A(n845), .B(n846), .Z(n844) );
  XNOR U826 ( .A(n843), .B(n847), .Z(n845) );
  XNOR U827 ( .A(n848), .B(n774), .Z(n777) );
  XNOR U828 ( .A(n849), .B(n850), .Z(n774) );
  AND U829 ( .A(n851), .B(n852), .Z(n850) );
  XOR U830 ( .A(n853), .B(n854), .Z(n851) );
  XNOR U831 ( .A(n855), .B(n856), .Z(n848) );
  NOR U832 ( .A(n857), .B(n858), .Z(n856) );
  XOR U833 ( .A(n855), .B(n859), .Z(n857) );
  XOR U834 ( .A(n783), .B(n782), .Z(n773) );
  XNOR U835 ( .A(n860), .B(n779), .Z(n782) );
  XOR U836 ( .A(n861), .B(n862), .Z(n779) );
  AND U837 ( .A(n863), .B(n864), .Z(n862) );
  XOR U838 ( .A(n861), .B(n865), .Z(n863) );
  XNOR U839 ( .A(n866), .B(n867), .Z(n860) );
  NOR U840 ( .A(n868), .B(n869), .Z(n867) );
  XNOR U841 ( .A(n866), .B(n870), .Z(n868) );
  XOR U842 ( .A(n871), .B(n872), .Z(n783) );
  NOR U843 ( .A(n873), .B(n874), .Z(n872) );
  XNOR U844 ( .A(n871), .B(n875), .Z(n873) );
  XNOR U845 ( .A(n680), .B(n787), .Z(n789) );
  XNOR U846 ( .A(n876), .B(n877), .Z(n680) );
  AND U847 ( .A(n66), .B(n687), .Z(n877) );
  XNOR U848 ( .A(n876), .B(n685), .Z(n687) );
  AND U849 ( .A(n690), .B(n693), .Z(n787) );
  XOR U850 ( .A(n878), .B(n836), .Z(n693) );
  XNOR U851 ( .A(p_input[0]), .B(p_input[128]), .Z(n836) );
  XOR U852 ( .A(n813), .B(n812), .Z(n878) );
  XOR U853 ( .A(n879), .B(n824), .Z(n812) );
  XOR U854 ( .A(n798), .B(n797), .Z(n824) );
  XNOR U855 ( .A(n880), .B(n803), .Z(n797) );
  XOR U856 ( .A(p_input[152]), .B(p_input[24]), .Z(n803) );
  XOR U857 ( .A(n794), .B(n802), .Z(n880) );
  XOR U858 ( .A(n881), .B(n799), .Z(n802) );
  XOR U859 ( .A(p_input[150]), .B(p_input[22]), .Z(n799) );
  XNOR U860 ( .A(p_input[151]), .B(p_input[23]), .Z(n881) );
  XOR U861 ( .A(p_input[146]), .B(p_input[18]), .Z(n794) );
  XNOR U862 ( .A(n808), .B(n807), .Z(n798) );
  XOR U863 ( .A(n882), .B(n804), .Z(n807) );
  XOR U864 ( .A(p_input[147]), .B(p_input[19]), .Z(n804) );
  XNOR U865 ( .A(p_input[148]), .B(p_input[20]), .Z(n882) );
  XOR U866 ( .A(p_input[149]), .B(p_input[21]), .Z(n808) );
  XNOR U867 ( .A(n823), .B(n809), .Z(n879) );
  XOR U868 ( .A(p_input[129]), .B(p_input[1]), .Z(n809) );
  XNOR U869 ( .A(n883), .B(n830), .Z(n823) );
  XNOR U870 ( .A(n819), .B(n818), .Z(n830) );
  XOR U871 ( .A(n884), .B(n815), .Z(n818) );
  XOR U872 ( .A(p_input[154]), .B(p_input[26]), .Z(n815) );
  XNOR U873 ( .A(p_input[155]), .B(p_input[27]), .Z(n884) );
  XOR U874 ( .A(p_input[156]), .B(p_input[28]), .Z(n819) );
  XNOR U875 ( .A(n829), .B(n820), .Z(n883) );
  XOR U876 ( .A(p_input[145]), .B(p_input[17]), .Z(n820) );
  XOR U877 ( .A(n885), .B(n835), .Z(n829) );
  XNOR U878 ( .A(p_input[159]), .B(p_input[31]), .Z(n835) );
  XOR U879 ( .A(n826), .B(n834), .Z(n885) );
  XOR U880 ( .A(n886), .B(n831), .Z(n834) );
  XOR U881 ( .A(p_input[157]), .B(p_input[29]), .Z(n831) );
  XNOR U882 ( .A(p_input[158]), .B(p_input[30]), .Z(n886) );
  XOR U883 ( .A(p_input[153]), .B(p_input[25]), .Z(n826) );
  XNOR U884 ( .A(n847), .B(n846), .Z(n813) );
  XNOR U885 ( .A(n887), .B(n854), .Z(n846) );
  XNOR U886 ( .A(n842), .B(n841), .Z(n854) );
  XNOR U887 ( .A(n888), .B(n889), .Z(n841) );
  IV U888 ( .A(n838), .Z(n889) );
  XOR U889 ( .A(p_input[11]), .B(p_input[139]), .Z(n838) );
  XNOR U890 ( .A(p_input[12]), .B(p_input[140]), .Z(n888) );
  XOR U891 ( .A(p_input[13]), .B(p_input[141]), .Z(n842) );
  XNOR U892 ( .A(n852), .B(n843), .Z(n887) );
  XOR U893 ( .A(p_input[130]), .B(p_input[2]), .Z(n843) );
  XOR U894 ( .A(n890), .B(n859), .Z(n852) );
  XNOR U895 ( .A(p_input[144]), .B(p_input[16]), .Z(n859) );
  XNOR U896 ( .A(n849), .B(n858), .Z(n890) );
  XOR U897 ( .A(n891), .B(n855), .Z(n858) );
  XOR U898 ( .A(p_input[142]), .B(p_input[14]), .Z(n855) );
  XNOR U899 ( .A(p_input[143]), .B(p_input[15]), .Z(n891) );
  IV U900 ( .A(n853), .Z(n849) );
  XOR U901 ( .A(p_input[10]), .B(p_input[138]), .Z(n853) );
  XNOR U902 ( .A(n865), .B(n864), .Z(n847) );
  XNOR U903 ( .A(n892), .B(n870), .Z(n864) );
  XOR U904 ( .A(p_input[137]), .B(p_input[9]), .Z(n870) );
  XOR U905 ( .A(n861), .B(n869), .Z(n892) );
  XOR U906 ( .A(n893), .B(n866), .Z(n869) );
  XOR U907 ( .A(p_input[135]), .B(p_input[7]), .Z(n866) );
  XNOR U908 ( .A(p_input[136]), .B(p_input[8]), .Z(n893) );
  XOR U909 ( .A(p_input[131]), .B(p_input[3]), .Z(n861) );
  XNOR U910 ( .A(n875), .B(n874), .Z(n865) );
  XOR U911 ( .A(n894), .B(n871), .Z(n874) );
  XOR U912 ( .A(p_input[132]), .B(p_input[4]), .Z(n871) );
  XNOR U913 ( .A(p_input[133]), .B(p_input[5]), .Z(n894) );
  XOR U914 ( .A(p_input[134]), .B(p_input[6]), .Z(n875) );
  XNOR U915 ( .A(n895), .B(n896), .Z(n690) );
  AND U916 ( .A(n66), .B(n897), .Z(n896) );
  XNOR U917 ( .A(n898), .B(n899), .Z(n66) );
  NOR U918 ( .A(n900), .B(n901), .Z(n899) );
  XOR U919 ( .A(n632), .B(n898), .Z(n901) );
  NOR U920 ( .A(n898), .B(n631), .Z(n900) );
  XOR U921 ( .A(n902), .B(n903), .Z(n898) );
  AND U922 ( .A(n904), .B(n905), .Z(n903) );
  XOR U923 ( .A(n902), .B(n712), .Z(n905) );
  XNOR U924 ( .A(n902), .B(n646), .Z(n904) );
  XOR U925 ( .A(n906), .B(n907), .Z(n902) );
  AND U926 ( .A(n908), .B(n909), .Z(n907) );
  XNOR U927 ( .A(n736), .B(n906), .Z(n909) );
  XNOR U928 ( .A(n906), .B(n738), .Z(n908) );
  IV U929 ( .A(n659), .Z(n738) );
  XOR U930 ( .A(n910), .B(n911), .Z(n906) );
  AND U931 ( .A(n912), .B(n913), .Z(n911) );
  XNOR U932 ( .A(n910), .B(n786), .Z(n912) );
  XOR U933 ( .A(n914), .B(n915), .Z(n688) );
  AND U934 ( .A(n70), .B(n897), .Z(n915) );
  XNOR U935 ( .A(n895), .B(n914), .Z(n897) );
  XOR U936 ( .A(n916), .B(n917), .Z(n70) );
  NOR U937 ( .A(n918), .B(n919), .Z(n917) );
  XOR U938 ( .A(n632), .B(n920), .Z(n919) );
  AND U939 ( .A(n921), .B(n922), .Z(n632) );
  NOR U940 ( .A(n920), .B(n631), .Z(n918) );
  AND U941 ( .A(n923), .B(n924), .Z(n631) );
  IV U942 ( .A(n916), .Z(n920) );
  XNOR U943 ( .A(n925), .B(n926), .Z(n916) );
  AND U944 ( .A(n927), .B(n928), .Z(n926) );
  XOR U945 ( .A(n712), .B(n925), .Z(n928) );
  XNOR U946 ( .A(n929), .B(n930), .Z(n712) );
  AND U947 ( .A(n74), .B(n931), .Z(n930) );
  XOR U948 ( .A(n932), .B(n929), .Z(n931) );
  XNOR U949 ( .A(n646), .B(n925), .Z(n927) );
  XOR U950 ( .A(n933), .B(n934), .Z(n646) );
  AND U951 ( .A(n80), .B(n935), .Z(n934) );
  XNOR U952 ( .A(n936), .B(n937), .Z(n935) );
  XOR U953 ( .A(n938), .B(n939), .Z(n925) );
  AND U954 ( .A(n940), .B(n941), .Z(n939) );
  XNOR U955 ( .A(n938), .B(n736), .Z(n941) );
  XNOR U956 ( .A(n942), .B(n943), .Z(n736) );
  AND U957 ( .A(n74), .B(n944), .Z(n943) );
  XNOR U958 ( .A(n945), .B(n942), .Z(n944) );
  XOR U959 ( .A(n659), .B(n938), .Z(n940) );
  XOR U960 ( .A(n946), .B(n947), .Z(n659) );
  AND U961 ( .A(n80), .B(n948), .Z(n947) );
  XOR U962 ( .A(n910), .B(n949), .Z(n938) );
  AND U963 ( .A(n950), .B(n913), .Z(n949) );
  XNOR U964 ( .A(n784), .B(n910), .Z(n913) );
  XNOR U965 ( .A(n951), .B(n952), .Z(n784) );
  AND U966 ( .A(n74), .B(n953), .Z(n952) );
  XNOR U967 ( .A(n954), .B(n951), .Z(n953) );
  XOR U968 ( .A(n672), .B(n910), .Z(n950) );
  IV U969 ( .A(n786), .Z(n672) );
  XOR U970 ( .A(n955), .B(n956), .Z(n786) );
  AND U971 ( .A(n80), .B(n957), .Z(n956) );
  XOR U972 ( .A(n958), .B(n959), .Z(n910) );
  AND U973 ( .A(n960), .B(n961), .Z(n959) );
  XNOR U974 ( .A(n958), .B(n876), .Z(n961) );
  XNOR U975 ( .A(n962), .B(n963), .Z(n876) );
  AND U976 ( .A(n74), .B(n964), .Z(n963) );
  XNOR U977 ( .A(n965), .B(n962), .Z(n964) );
  XOR U978 ( .A(n966), .B(n958), .Z(n960) );
  IV U979 ( .A(n685), .Z(n966) );
  XOR U980 ( .A(n967), .B(n968), .Z(n685) );
  AND U981 ( .A(n80), .B(n969), .Z(n968) );
  AND U982 ( .A(n914), .B(n895), .Z(n958) );
  XNOR U983 ( .A(n970), .B(n971), .Z(n895) );
  AND U984 ( .A(n74), .B(n972), .Z(n971) );
  XNOR U985 ( .A(n973), .B(n970), .Z(n972) );
  XNOR U986 ( .A(n974), .B(n975), .Z(n74) );
  NOR U987 ( .A(n976), .B(n977), .Z(n975) );
  XOR U988 ( .A(n974), .B(n923), .Z(n977) );
  IV U989 ( .A(n978), .Z(n923) );
  AND U990 ( .A(n979), .B(n980), .Z(n978) );
  NOR U991 ( .A(n974), .B(n924), .Z(n976) );
  AND U992 ( .A(n932), .B(n981), .Z(n924) );
  XOR U993 ( .A(n982), .B(n983), .Z(n974) );
  AND U994 ( .A(n984), .B(n985), .Z(n983) );
  XNOR U995 ( .A(n982), .B(n932), .Z(n985) );
  XNOR U996 ( .A(n986), .B(n987), .Z(n932) );
  XOR U997 ( .A(n988), .B(n981), .Z(n987) );
  AND U998 ( .A(n945), .B(n989), .Z(n981) );
  AND U999 ( .A(n990), .B(n991), .Z(n988) );
  XOR U1000 ( .A(n992), .B(n986), .Z(n990) );
  XOR U1001 ( .A(n929), .B(n982), .Z(n984) );
  NOR U1002 ( .A(n993), .B(n936), .Z(n929) );
  AND U1003 ( .A(n77), .B(n933), .Z(n993) );
  XOR U1004 ( .A(n994), .B(n995), .Z(n982) );
  AND U1005 ( .A(n996), .B(n997), .Z(n995) );
  XNOR U1006 ( .A(n994), .B(n945), .Z(n997) );
  XOR U1007 ( .A(n998), .B(n991), .Z(n945) );
  XNOR U1008 ( .A(n999), .B(n986), .Z(n991) );
  XOR U1009 ( .A(n1000), .B(n1001), .Z(n986) );
  AND U1010 ( .A(n1002), .B(n1003), .Z(n1001) );
  XOR U1011 ( .A(n1004), .B(n1000), .Z(n1002) );
  XNOR U1012 ( .A(n1005), .B(n1006), .Z(n999) );
  AND U1013 ( .A(n1007), .B(n1008), .Z(n1006) );
  XOR U1014 ( .A(n1005), .B(n1009), .Z(n1007) );
  XNOR U1015 ( .A(n992), .B(n989), .Z(n998) );
  AND U1016 ( .A(n954), .B(n1010), .Z(n989) );
  XOR U1017 ( .A(n1011), .B(n1012), .Z(n992) );
  AND U1018 ( .A(n1013), .B(n1014), .Z(n1012) );
  XOR U1019 ( .A(n1011), .B(n1015), .Z(n1013) );
  XNOR U1020 ( .A(n942), .B(n994), .Z(n996) );
  XNOR U1021 ( .A(n1016), .B(n1017), .Z(n942) );
  AND U1022 ( .A(n77), .B(n948), .Z(n1017) );
  XOR U1023 ( .A(n1016), .B(n946), .Z(n948) );
  XOR U1024 ( .A(n1018), .B(n1019), .Z(n994) );
  AND U1025 ( .A(n1020), .B(n1021), .Z(n1019) );
  XOR U1026 ( .A(n1018), .B(n1022), .Z(n1021) );
  IV U1027 ( .A(n954), .Z(n1022) );
  XOR U1028 ( .A(n1023), .B(n1003), .Z(n954) );
  XNOR U1029 ( .A(n1024), .B(n1009), .Z(n1003) );
  XOR U1030 ( .A(n1025), .B(n1026), .Z(n1009) );
  AND U1031 ( .A(n1027), .B(n1028), .Z(n1026) );
  XOR U1032 ( .A(n1025), .B(n1029), .Z(n1027) );
  XNOR U1033 ( .A(n1008), .B(n1000), .Z(n1024) );
  XOR U1034 ( .A(n1030), .B(n1031), .Z(n1000) );
  AND U1035 ( .A(n1032), .B(n1033), .Z(n1031) );
  XNOR U1036 ( .A(n1034), .B(n1030), .Z(n1032) );
  XNOR U1037 ( .A(n1035), .B(n1005), .Z(n1008) );
  XOR U1038 ( .A(n1036), .B(n1037), .Z(n1005) );
  AND U1039 ( .A(n1038), .B(n1039), .Z(n1037) );
  XOR U1040 ( .A(n1036), .B(n1040), .Z(n1038) );
  XNOR U1041 ( .A(n1041), .B(n1042), .Z(n1035) );
  AND U1042 ( .A(n1043), .B(n1044), .Z(n1042) );
  XNOR U1043 ( .A(n1041), .B(n1045), .Z(n1043) );
  XNOR U1044 ( .A(n1004), .B(n1010), .Z(n1023) );
  AND U1045 ( .A(n965), .B(n1046), .Z(n1010) );
  XOR U1046 ( .A(n1015), .B(n1014), .Z(n1004) );
  XNOR U1047 ( .A(n1047), .B(n1011), .Z(n1014) );
  XOR U1048 ( .A(n1048), .B(n1049), .Z(n1011) );
  AND U1049 ( .A(n1050), .B(n1051), .Z(n1049) );
  XOR U1050 ( .A(n1048), .B(n1052), .Z(n1050) );
  XNOR U1051 ( .A(n1053), .B(n1054), .Z(n1047) );
  AND U1052 ( .A(n1055), .B(n1056), .Z(n1054) );
  XOR U1053 ( .A(n1053), .B(n1057), .Z(n1055) );
  XOR U1054 ( .A(n1058), .B(n1059), .Z(n1015) );
  AND U1055 ( .A(n1060), .B(n1061), .Z(n1059) );
  XOR U1056 ( .A(n1058), .B(n1062), .Z(n1060) );
  XNOR U1057 ( .A(n951), .B(n1018), .Z(n1020) );
  XNOR U1058 ( .A(n1063), .B(n1064), .Z(n951) );
  AND U1059 ( .A(n77), .B(n957), .Z(n1064) );
  XNOR U1060 ( .A(n1063), .B(n955), .Z(n957) );
  XOR U1061 ( .A(n1065), .B(n1066), .Z(n1018) );
  AND U1062 ( .A(n1067), .B(n1068), .Z(n1066) );
  XNOR U1063 ( .A(n1065), .B(n965), .Z(n1068) );
  XOR U1064 ( .A(n1069), .B(n1033), .Z(n965) );
  XNOR U1065 ( .A(n1070), .B(n1040), .Z(n1033) );
  XOR U1066 ( .A(n1029), .B(n1028), .Z(n1040) );
  XNOR U1067 ( .A(n1071), .B(n1025), .Z(n1028) );
  XOR U1068 ( .A(n1072), .B(n1073), .Z(n1025) );
  AND U1069 ( .A(n1074), .B(n1075), .Z(n1073) );
  XOR U1070 ( .A(n1072), .B(n1076), .Z(n1074) );
  XNOR U1071 ( .A(n1077), .B(n1078), .Z(n1071) );
  NOR U1072 ( .A(n1079), .B(n1080), .Z(n1078) );
  XNOR U1073 ( .A(n1077), .B(n1081), .Z(n1079) );
  XOR U1074 ( .A(n1082), .B(n1083), .Z(n1029) );
  NOR U1075 ( .A(n1084), .B(n1085), .Z(n1083) );
  XNOR U1076 ( .A(n1082), .B(n1086), .Z(n1084) );
  XNOR U1077 ( .A(n1039), .B(n1030), .Z(n1070) );
  XOR U1078 ( .A(n1087), .B(n1088), .Z(n1030) );
  NOR U1079 ( .A(n1089), .B(n1090), .Z(n1088) );
  XNOR U1080 ( .A(n1087), .B(n1091), .Z(n1089) );
  XOR U1081 ( .A(n1092), .B(n1045), .Z(n1039) );
  XNOR U1082 ( .A(n1093), .B(n1094), .Z(n1045) );
  NOR U1083 ( .A(n1095), .B(n1096), .Z(n1094) );
  XNOR U1084 ( .A(n1093), .B(n1097), .Z(n1095) );
  XNOR U1085 ( .A(n1044), .B(n1036), .Z(n1092) );
  XOR U1086 ( .A(n1098), .B(n1099), .Z(n1036) );
  AND U1087 ( .A(n1100), .B(n1101), .Z(n1099) );
  XOR U1088 ( .A(n1098), .B(n1102), .Z(n1100) );
  XNOR U1089 ( .A(n1103), .B(n1041), .Z(n1044) );
  XOR U1090 ( .A(n1104), .B(n1105), .Z(n1041) );
  AND U1091 ( .A(n1106), .B(n1107), .Z(n1105) );
  XOR U1092 ( .A(n1104), .B(n1108), .Z(n1106) );
  XNOR U1093 ( .A(n1109), .B(n1110), .Z(n1103) );
  NOR U1094 ( .A(n1111), .B(n1112), .Z(n1110) );
  XOR U1095 ( .A(n1109), .B(n1113), .Z(n1111) );
  XOR U1096 ( .A(n1034), .B(n1046), .Z(n1069) );
  NOR U1097 ( .A(n973), .B(n1114), .Z(n1046) );
  XNOR U1098 ( .A(n1052), .B(n1051), .Z(n1034) );
  XNOR U1099 ( .A(n1115), .B(n1057), .Z(n1051) );
  XOR U1100 ( .A(n1116), .B(n1117), .Z(n1057) );
  NOR U1101 ( .A(n1118), .B(n1119), .Z(n1117) );
  XNOR U1102 ( .A(n1116), .B(n1120), .Z(n1118) );
  XNOR U1103 ( .A(n1056), .B(n1048), .Z(n1115) );
  XOR U1104 ( .A(n1121), .B(n1122), .Z(n1048) );
  AND U1105 ( .A(n1123), .B(n1124), .Z(n1122) );
  XNOR U1106 ( .A(n1121), .B(n1125), .Z(n1123) );
  XNOR U1107 ( .A(n1126), .B(n1053), .Z(n1056) );
  XOR U1108 ( .A(n1127), .B(n1128), .Z(n1053) );
  AND U1109 ( .A(n1129), .B(n1130), .Z(n1128) );
  XOR U1110 ( .A(n1127), .B(n1131), .Z(n1129) );
  XNOR U1111 ( .A(n1132), .B(n1133), .Z(n1126) );
  NOR U1112 ( .A(n1134), .B(n1135), .Z(n1133) );
  XOR U1113 ( .A(n1132), .B(n1136), .Z(n1134) );
  XOR U1114 ( .A(n1062), .B(n1061), .Z(n1052) );
  XNOR U1115 ( .A(n1137), .B(n1058), .Z(n1061) );
  XOR U1116 ( .A(n1138), .B(n1139), .Z(n1058) );
  AND U1117 ( .A(n1140), .B(n1141), .Z(n1139) );
  XOR U1118 ( .A(n1138), .B(n1142), .Z(n1140) );
  XNOR U1119 ( .A(n1143), .B(n1144), .Z(n1137) );
  NOR U1120 ( .A(n1145), .B(n1146), .Z(n1144) );
  XNOR U1121 ( .A(n1143), .B(n1147), .Z(n1145) );
  XOR U1122 ( .A(n1148), .B(n1149), .Z(n1062) );
  NOR U1123 ( .A(n1150), .B(n1151), .Z(n1149) );
  XNOR U1124 ( .A(n1148), .B(n1152), .Z(n1150) );
  XNOR U1125 ( .A(n962), .B(n1065), .Z(n1067) );
  XNOR U1126 ( .A(n1153), .B(n1154), .Z(n962) );
  AND U1127 ( .A(n77), .B(n969), .Z(n1154) );
  XNOR U1128 ( .A(n1153), .B(n967), .Z(n969) );
  AND U1129 ( .A(n970), .B(n973), .Z(n1065) );
  XOR U1130 ( .A(n1155), .B(n1114), .Z(n973) );
  XNOR U1131 ( .A(p_input[128]), .B(p_input[32]), .Z(n1114) );
  XOR U1132 ( .A(n1091), .B(n1090), .Z(n1155) );
  XOR U1133 ( .A(n1156), .B(n1102), .Z(n1090) );
  XOR U1134 ( .A(n1076), .B(n1075), .Z(n1102) );
  XNOR U1135 ( .A(n1157), .B(n1081), .Z(n1075) );
  XOR U1136 ( .A(p_input[152]), .B(p_input[56]), .Z(n1081) );
  XOR U1137 ( .A(n1072), .B(n1080), .Z(n1157) );
  XOR U1138 ( .A(n1158), .B(n1077), .Z(n1080) );
  XOR U1139 ( .A(p_input[150]), .B(p_input[54]), .Z(n1077) );
  XNOR U1140 ( .A(p_input[151]), .B(p_input[55]), .Z(n1158) );
  XOR U1141 ( .A(p_input[146]), .B(p_input[50]), .Z(n1072) );
  XNOR U1142 ( .A(n1086), .B(n1085), .Z(n1076) );
  XOR U1143 ( .A(n1159), .B(n1082), .Z(n1085) );
  XOR U1144 ( .A(p_input[147]), .B(p_input[51]), .Z(n1082) );
  XNOR U1145 ( .A(p_input[148]), .B(p_input[52]), .Z(n1159) );
  XOR U1146 ( .A(p_input[149]), .B(p_input[53]), .Z(n1086) );
  XNOR U1147 ( .A(n1101), .B(n1087), .Z(n1156) );
  XOR U1148 ( .A(p_input[129]), .B(p_input[33]), .Z(n1087) );
  XNOR U1149 ( .A(n1160), .B(n1108), .Z(n1101) );
  XNOR U1150 ( .A(n1097), .B(n1096), .Z(n1108) );
  XOR U1151 ( .A(n1161), .B(n1093), .Z(n1096) );
  XOR U1152 ( .A(p_input[154]), .B(p_input[58]), .Z(n1093) );
  XNOR U1153 ( .A(p_input[155]), .B(p_input[59]), .Z(n1161) );
  XOR U1154 ( .A(p_input[156]), .B(p_input[60]), .Z(n1097) );
  XNOR U1155 ( .A(n1107), .B(n1098), .Z(n1160) );
  XOR U1156 ( .A(p_input[145]), .B(p_input[49]), .Z(n1098) );
  XOR U1157 ( .A(n1162), .B(n1113), .Z(n1107) );
  XNOR U1158 ( .A(p_input[159]), .B(p_input[63]), .Z(n1113) );
  XOR U1159 ( .A(n1104), .B(n1112), .Z(n1162) );
  XOR U1160 ( .A(n1163), .B(n1109), .Z(n1112) );
  XOR U1161 ( .A(p_input[157]), .B(p_input[61]), .Z(n1109) );
  XNOR U1162 ( .A(p_input[158]), .B(p_input[62]), .Z(n1163) );
  XOR U1163 ( .A(p_input[153]), .B(p_input[57]), .Z(n1104) );
  XNOR U1164 ( .A(n1125), .B(n1124), .Z(n1091) );
  XNOR U1165 ( .A(n1164), .B(n1131), .Z(n1124) );
  XNOR U1166 ( .A(n1120), .B(n1119), .Z(n1131) );
  XOR U1167 ( .A(n1165), .B(n1116), .Z(n1119) );
  XOR U1168 ( .A(p_input[139]), .B(p_input[43]), .Z(n1116) );
  XOR U1169 ( .A(n1166), .B(p_input[44]), .Z(n1165) );
  XOR U1170 ( .A(p_input[141]), .B(p_input[45]), .Z(n1120) );
  XNOR U1171 ( .A(n1130), .B(n1121), .Z(n1164) );
  XOR U1172 ( .A(p_input[130]), .B(p_input[34]), .Z(n1121) );
  XOR U1173 ( .A(n1167), .B(n1136), .Z(n1130) );
  XNOR U1174 ( .A(p_input[144]), .B(p_input[48]), .Z(n1136) );
  XOR U1175 ( .A(n1127), .B(n1135), .Z(n1167) );
  XOR U1176 ( .A(n1168), .B(n1132), .Z(n1135) );
  XOR U1177 ( .A(p_input[142]), .B(p_input[46]), .Z(n1132) );
  XNOR U1178 ( .A(p_input[143]), .B(p_input[47]), .Z(n1168) );
  XOR U1179 ( .A(p_input[138]), .B(p_input[42]), .Z(n1127) );
  XNOR U1180 ( .A(n1142), .B(n1141), .Z(n1125) );
  XNOR U1181 ( .A(n1169), .B(n1147), .Z(n1141) );
  XOR U1182 ( .A(p_input[137]), .B(p_input[41]), .Z(n1147) );
  XOR U1183 ( .A(n1138), .B(n1146), .Z(n1169) );
  XOR U1184 ( .A(n1170), .B(n1143), .Z(n1146) );
  XOR U1185 ( .A(p_input[135]), .B(p_input[39]), .Z(n1143) );
  XNOR U1186 ( .A(p_input[136]), .B(p_input[40]), .Z(n1170) );
  XOR U1187 ( .A(p_input[131]), .B(p_input[35]), .Z(n1138) );
  XNOR U1188 ( .A(n1152), .B(n1151), .Z(n1142) );
  XOR U1189 ( .A(n1171), .B(n1148), .Z(n1151) );
  XOR U1190 ( .A(p_input[132]), .B(p_input[36]), .Z(n1148) );
  XNOR U1191 ( .A(p_input[133]), .B(p_input[37]), .Z(n1171) );
  XOR U1192 ( .A(p_input[134]), .B(p_input[38]), .Z(n1152) );
  XOR U1193 ( .A(n1172), .B(n1173), .Z(n970) );
  AND U1194 ( .A(n77), .B(n1174), .Z(n1173) );
  XNOR U1195 ( .A(n1175), .B(n1176), .Z(n77) );
  NOR U1196 ( .A(n1177), .B(n1178), .Z(n1176) );
  XNOR U1197 ( .A(n980), .B(n1175), .Z(n1178) );
  NOR U1198 ( .A(n1175), .B(n921), .Z(n1177) );
  XOR U1199 ( .A(n1179), .B(n1180), .Z(n1175) );
  AND U1200 ( .A(n1181), .B(n1182), .Z(n1180) );
  XOR U1201 ( .A(n936), .B(n1179), .Z(n1182) );
  XNOR U1202 ( .A(n1179), .B(n933), .Z(n1181) );
  XOR U1203 ( .A(n1183), .B(n1184), .Z(n1179) );
  AND U1204 ( .A(n1185), .B(n1186), .Z(n1184) );
  XNOR U1205 ( .A(n1016), .B(n1183), .Z(n1186) );
  XOR U1206 ( .A(n1183), .B(n946), .Z(n1185) );
  XOR U1207 ( .A(n1187), .B(n1188), .Z(n1183) );
  AND U1208 ( .A(n1189), .B(n1190), .Z(n1188) );
  XNOR U1209 ( .A(n1187), .B(n955), .Z(n1189) );
  XOR U1210 ( .A(n1191), .B(n1192), .Z(n914) );
  AND U1211 ( .A(n80), .B(n1174), .Z(n1192) );
  XNOR U1212 ( .A(n1193), .B(n1191), .Z(n1174) );
  XOR U1213 ( .A(n1194), .B(n1195), .Z(n80) );
  MUX U1214 ( .IN0(n979), .IN1(n980), .SEL(n1194), .F(n1195) );
  IV U1215 ( .A(n922), .Z(n980) );
  AND U1216 ( .A(n937), .B(n1196), .Z(n922) );
  IV U1217 ( .A(n921), .Z(n979) );
  AND U1218 ( .A(n1197), .B(n1198), .Z(n921) );
  IV U1219 ( .A(n936), .Z(n1197) );
  XOR U1220 ( .A(n1199), .B(n1200), .Z(n1194) );
  AND U1221 ( .A(n1201), .B(n1202), .Z(n1200) );
  XOR U1222 ( .A(n1199), .B(n936), .Z(n1202) );
  XOR U1223 ( .A(n1203), .B(n1204), .Z(n936) );
  XOR U1224 ( .A(n1205), .B(n1198), .Z(n1204) );
  AND U1225 ( .A(n1016), .B(n1206), .Z(n1198) );
  AND U1226 ( .A(n1207), .B(n1208), .Z(n1205) );
  XOR U1227 ( .A(n1209), .B(n1203), .Z(n1207) );
  XOR U1228 ( .A(n937), .B(n1199), .Z(n1201) );
  IV U1229 ( .A(n933), .Z(n937) );
  XOR U1230 ( .A(n1210), .B(n1211), .Z(n933) );
  XOR U1231 ( .A(n1212), .B(n1196), .Z(n1211) );
  AND U1232 ( .A(n946), .B(n1213), .Z(n1196) );
  AND U1233 ( .A(n1214), .B(n1215), .Z(n1212) );
  XNOR U1234 ( .A(n1210), .B(n1216), .Z(n1214) );
  XOR U1235 ( .A(n1217), .B(n1218), .Z(n1199) );
  AND U1236 ( .A(n1219), .B(n1220), .Z(n1218) );
  XNOR U1237 ( .A(n1217), .B(n1016), .Z(n1220) );
  XOR U1238 ( .A(n1221), .B(n1208), .Z(n1016) );
  XNOR U1239 ( .A(n1222), .B(n1203), .Z(n1208) );
  XOR U1240 ( .A(n1223), .B(n1224), .Z(n1203) );
  AND U1241 ( .A(n1225), .B(n1226), .Z(n1224) );
  XOR U1242 ( .A(n1227), .B(n1223), .Z(n1225) );
  XNOR U1243 ( .A(n1228), .B(n1229), .Z(n1222) );
  AND U1244 ( .A(n1230), .B(n1231), .Z(n1229) );
  XOR U1245 ( .A(n1228), .B(n1232), .Z(n1230) );
  XNOR U1246 ( .A(n1209), .B(n1206), .Z(n1221) );
  AND U1247 ( .A(n1063), .B(n1233), .Z(n1206) );
  XOR U1248 ( .A(n1234), .B(n1235), .Z(n1209) );
  AND U1249 ( .A(n1236), .B(n1237), .Z(n1235) );
  XOR U1250 ( .A(n1234), .B(n1238), .Z(n1236) );
  XOR U1251 ( .A(n946), .B(n1217), .Z(n1219) );
  XNOR U1252 ( .A(n1239), .B(n1216), .Z(n946) );
  XNOR U1253 ( .A(n1240), .B(n1241), .Z(n1216) );
  AND U1254 ( .A(n1242), .B(n1243), .Z(n1241) );
  XOR U1255 ( .A(n1240), .B(n1244), .Z(n1242) );
  XNOR U1256 ( .A(n1215), .B(n1213), .Z(n1239) );
  AND U1257 ( .A(n1245), .B(n1246), .Z(n1213) );
  XNOR U1258 ( .A(n1247), .B(n1210), .Z(n1215) );
  XOR U1259 ( .A(n1248), .B(n1249), .Z(n1210) );
  AND U1260 ( .A(n1250), .B(n1251), .Z(n1249) );
  XOR U1261 ( .A(n1248), .B(n1252), .Z(n1250) );
  XNOR U1262 ( .A(n1253), .B(n1254), .Z(n1247) );
  AND U1263 ( .A(n1255), .B(n1256), .Z(n1254) );
  XNOR U1264 ( .A(n1253), .B(n1257), .Z(n1255) );
  XOR U1265 ( .A(n1187), .B(n1258), .Z(n1217) );
  AND U1266 ( .A(n1259), .B(n1190), .Z(n1258) );
  XNOR U1267 ( .A(n1063), .B(n1187), .Z(n1190) );
  XOR U1268 ( .A(n1260), .B(n1226), .Z(n1063) );
  XNOR U1269 ( .A(n1261), .B(n1232), .Z(n1226) );
  XOR U1270 ( .A(n1262), .B(n1263), .Z(n1232) );
  AND U1271 ( .A(n1264), .B(n1265), .Z(n1263) );
  XOR U1272 ( .A(n1262), .B(n1266), .Z(n1264) );
  XNOR U1273 ( .A(n1231), .B(n1223), .Z(n1261) );
  XOR U1274 ( .A(n1267), .B(n1268), .Z(n1223) );
  AND U1275 ( .A(n1269), .B(n1270), .Z(n1268) );
  XNOR U1276 ( .A(n1271), .B(n1267), .Z(n1269) );
  XNOR U1277 ( .A(n1272), .B(n1228), .Z(n1231) );
  XOR U1278 ( .A(n1273), .B(n1274), .Z(n1228) );
  AND U1279 ( .A(n1275), .B(n1276), .Z(n1274) );
  XOR U1280 ( .A(n1273), .B(n1277), .Z(n1275) );
  XNOR U1281 ( .A(n1278), .B(n1279), .Z(n1272) );
  AND U1282 ( .A(n1280), .B(n1281), .Z(n1279) );
  XNOR U1283 ( .A(n1278), .B(n1282), .Z(n1280) );
  XNOR U1284 ( .A(n1227), .B(n1233), .Z(n1260) );
  AND U1285 ( .A(n1153), .B(n1283), .Z(n1233) );
  XOR U1286 ( .A(n1238), .B(n1237), .Z(n1227) );
  XNOR U1287 ( .A(n1284), .B(n1234), .Z(n1237) );
  XOR U1288 ( .A(n1285), .B(n1286), .Z(n1234) );
  AND U1289 ( .A(n1287), .B(n1288), .Z(n1286) );
  XOR U1290 ( .A(n1285), .B(n1289), .Z(n1287) );
  XNOR U1291 ( .A(n1290), .B(n1291), .Z(n1284) );
  AND U1292 ( .A(n1292), .B(n1293), .Z(n1291) );
  XOR U1293 ( .A(n1290), .B(n1294), .Z(n1292) );
  XOR U1294 ( .A(n1295), .B(n1296), .Z(n1238) );
  AND U1295 ( .A(n1297), .B(n1298), .Z(n1296) );
  XOR U1296 ( .A(n1295), .B(n1299), .Z(n1297) );
  XOR U1297 ( .A(n1245), .B(n1187), .Z(n1259) );
  IV U1298 ( .A(n955), .Z(n1245) );
  XNOR U1299 ( .A(n1300), .B(n1252), .Z(n955) );
  XOR U1300 ( .A(n1244), .B(n1243), .Z(n1252) );
  XNOR U1301 ( .A(n1301), .B(n1240), .Z(n1243) );
  XOR U1302 ( .A(n1302), .B(n1303), .Z(n1240) );
  AND U1303 ( .A(n1304), .B(n1305), .Z(n1303) );
  XOR U1304 ( .A(n1302), .B(n1306), .Z(n1304) );
  XNOR U1305 ( .A(n1307), .B(n1308), .Z(n1301) );
  AND U1306 ( .A(n1309), .B(n1310), .Z(n1308) );
  XOR U1307 ( .A(n1307), .B(n1311), .Z(n1309) );
  XOR U1308 ( .A(n1312), .B(n1313), .Z(n1244) );
  AND U1309 ( .A(n1314), .B(n1315), .Z(n1313) );
  XOR U1310 ( .A(n1312), .B(n1316), .Z(n1314) );
  XNOR U1311 ( .A(n1251), .B(n1246), .Z(n1300) );
  AND U1312 ( .A(n1317), .B(n1318), .Z(n1246) );
  XOR U1313 ( .A(n1319), .B(n1257), .Z(n1251) );
  XNOR U1314 ( .A(n1320), .B(n1321), .Z(n1257) );
  AND U1315 ( .A(n1322), .B(n1323), .Z(n1321) );
  XOR U1316 ( .A(n1320), .B(n1324), .Z(n1322) );
  XNOR U1317 ( .A(n1256), .B(n1248), .Z(n1319) );
  XOR U1318 ( .A(n1325), .B(n1326), .Z(n1248) );
  AND U1319 ( .A(n1327), .B(n1328), .Z(n1326) );
  XOR U1320 ( .A(n1325), .B(n1329), .Z(n1327) );
  XNOR U1321 ( .A(n1330), .B(n1253), .Z(n1256) );
  XOR U1322 ( .A(n1331), .B(n1332), .Z(n1253) );
  AND U1323 ( .A(n1333), .B(n1334), .Z(n1332) );
  XOR U1324 ( .A(n1331), .B(n1335), .Z(n1333) );
  XNOR U1325 ( .A(n1336), .B(n1337), .Z(n1330) );
  AND U1326 ( .A(n1338), .B(n1339), .Z(n1337) );
  XNOR U1327 ( .A(n1336), .B(n1340), .Z(n1338) );
  XOR U1328 ( .A(n1341), .B(n1342), .Z(n1187) );
  AND U1329 ( .A(n1343), .B(n1344), .Z(n1342) );
  XNOR U1330 ( .A(n1341), .B(n1153), .Z(n1344) );
  XOR U1331 ( .A(n1345), .B(n1270), .Z(n1153) );
  XNOR U1332 ( .A(n1346), .B(n1277), .Z(n1270) );
  XOR U1333 ( .A(n1266), .B(n1265), .Z(n1277) );
  XNOR U1334 ( .A(n1347), .B(n1262), .Z(n1265) );
  XNOR U1335 ( .A(n1348), .B(n1349), .Z(n1262) );
  AND U1336 ( .A(n1350), .B(n1351), .Z(n1349) );
  XOR U1337 ( .A(n1352), .B(n1353), .Z(n1350) );
  XNOR U1338 ( .A(n1354), .B(n1355), .Z(n1347) );
  AND U1339 ( .A(n1356), .B(n1357), .Z(n1355) );
  XNOR U1340 ( .A(n1354), .B(n1358), .Z(n1356) );
  XOR U1341 ( .A(n1359), .B(n1360), .Z(n1266) );
  AND U1342 ( .A(n1361), .B(n1362), .Z(n1360) );
  XOR U1343 ( .A(n1359), .B(n1363), .Z(n1361) );
  XNOR U1344 ( .A(n1276), .B(n1267), .Z(n1346) );
  XOR U1345 ( .A(n1364), .B(n1365), .Z(n1267) );
  NOR U1346 ( .A(n1366), .B(n1367), .Z(n1365) );
  XNOR U1347 ( .A(n1364), .B(n1368), .Z(n1366) );
  XOR U1348 ( .A(n1369), .B(n1282), .Z(n1276) );
  XNOR U1349 ( .A(n1370), .B(n1371), .Z(n1282) );
  AND U1350 ( .A(n1372), .B(n1373), .Z(n1371) );
  XOR U1351 ( .A(n1370), .B(n1374), .Z(n1372) );
  XNOR U1352 ( .A(n1281), .B(n1273), .Z(n1369) );
  XOR U1353 ( .A(n1375), .B(n1376), .Z(n1273) );
  AND U1354 ( .A(n1377), .B(n1378), .Z(n1376) );
  XOR U1355 ( .A(n1375), .B(n1379), .Z(n1377) );
  XNOR U1356 ( .A(n1380), .B(n1278), .Z(n1281) );
  XNOR U1357 ( .A(n1381), .B(n1382), .Z(n1278) );
  AND U1358 ( .A(n1383), .B(n1384), .Z(n1382) );
  XOR U1359 ( .A(n1385), .B(n1386), .Z(n1383) );
  XNOR U1360 ( .A(n1387), .B(n1388), .Z(n1380) );
  AND U1361 ( .A(n1389), .B(n1390), .Z(n1388) );
  XNOR U1362 ( .A(n1387), .B(n1391), .Z(n1389) );
  XOR U1363 ( .A(n1271), .B(n1283), .Z(n1345) );
  AND U1364 ( .A(n1172), .B(n1392), .Z(n1283) );
  XNOR U1365 ( .A(n1289), .B(n1288), .Z(n1271) );
  XNOR U1366 ( .A(n1393), .B(n1294), .Z(n1288) );
  XOR U1367 ( .A(n1394), .B(n1395), .Z(n1294) );
  NOR U1368 ( .A(n1396), .B(n1397), .Z(n1395) );
  XNOR U1369 ( .A(n1394), .B(n1398), .Z(n1396) );
  XNOR U1370 ( .A(n1293), .B(n1285), .Z(n1393) );
  XOR U1371 ( .A(n1399), .B(n1400), .Z(n1285) );
  AND U1372 ( .A(n1401), .B(n1402), .Z(n1400) );
  XNOR U1373 ( .A(n1399), .B(n1403), .Z(n1401) );
  XNOR U1374 ( .A(n1404), .B(n1290), .Z(n1293) );
  XOR U1375 ( .A(n1405), .B(n1406), .Z(n1290) );
  AND U1376 ( .A(n1407), .B(n1408), .Z(n1406) );
  XOR U1377 ( .A(n1405), .B(n1409), .Z(n1407) );
  XNOR U1378 ( .A(n1410), .B(n1411), .Z(n1404) );
  AND U1379 ( .A(n1412), .B(n1413), .Z(n1411) );
  XNOR U1380 ( .A(n1410), .B(n1414), .Z(n1412) );
  XOR U1381 ( .A(n1299), .B(n1298), .Z(n1289) );
  XNOR U1382 ( .A(n1415), .B(n1295), .Z(n1298) );
  XNOR U1383 ( .A(n1416), .B(n1417), .Z(n1295) );
  AND U1384 ( .A(n1418), .B(n1419), .Z(n1417) );
  XOR U1385 ( .A(n1420), .B(n1421), .Z(n1418) );
  XNOR U1386 ( .A(n1422), .B(n1423), .Z(n1415) );
  AND U1387 ( .A(n1424), .B(n1425), .Z(n1423) );
  XNOR U1388 ( .A(n1422), .B(n1426), .Z(n1424) );
  XOR U1389 ( .A(n1427), .B(n1428), .Z(n1299) );
  AND U1390 ( .A(n1429), .B(n1430), .Z(n1428) );
  XOR U1391 ( .A(n1427), .B(n1431), .Z(n1429) );
  XOR U1392 ( .A(n1317), .B(n1341), .Z(n1343) );
  IV U1393 ( .A(n967), .Z(n1317) );
  XNOR U1394 ( .A(n1432), .B(n1329), .Z(n967) );
  XOR U1395 ( .A(n1306), .B(n1305), .Z(n1329) );
  XNOR U1396 ( .A(n1433), .B(n1311), .Z(n1305) );
  XOR U1397 ( .A(n1434), .B(n1435), .Z(n1311) );
  NOR U1398 ( .A(n1436), .B(n1437), .Z(n1435) );
  XNOR U1399 ( .A(n1434), .B(n1438), .Z(n1436) );
  XNOR U1400 ( .A(n1310), .B(n1302), .Z(n1433) );
  XOR U1401 ( .A(n1439), .B(n1440), .Z(n1302) );
  AND U1402 ( .A(n1441), .B(n1442), .Z(n1440) );
  XNOR U1403 ( .A(n1439), .B(n1443), .Z(n1441) );
  XNOR U1404 ( .A(n1444), .B(n1307), .Z(n1310) );
  XOR U1405 ( .A(n1445), .B(n1446), .Z(n1307) );
  AND U1406 ( .A(n1447), .B(n1448), .Z(n1446) );
  XOR U1407 ( .A(n1445), .B(n1449), .Z(n1447) );
  XNOR U1408 ( .A(n1450), .B(n1451), .Z(n1444) );
  NOR U1409 ( .A(n1452), .B(n1453), .Z(n1451) );
  XOR U1410 ( .A(n1450), .B(n1454), .Z(n1452) );
  XOR U1411 ( .A(n1316), .B(n1315), .Z(n1306) );
  XNOR U1412 ( .A(n1455), .B(n1312), .Z(n1315) );
  XOR U1413 ( .A(n1456), .B(n1457), .Z(n1312) );
  AND U1414 ( .A(n1458), .B(n1459), .Z(n1457) );
  XOR U1415 ( .A(n1456), .B(n1460), .Z(n1458) );
  XNOR U1416 ( .A(n1461), .B(n1462), .Z(n1455) );
  NOR U1417 ( .A(n1463), .B(n1464), .Z(n1462) );
  XNOR U1418 ( .A(n1461), .B(n1465), .Z(n1463) );
  XOR U1419 ( .A(n1466), .B(n1467), .Z(n1316) );
  NOR U1420 ( .A(n1468), .B(n1469), .Z(n1467) );
  XNOR U1421 ( .A(n1466), .B(n1470), .Z(n1468) );
  XNOR U1422 ( .A(n1328), .B(n1318), .Z(n1432) );
  AND U1423 ( .A(n1191), .B(n1471), .Z(n1318) );
  XNOR U1424 ( .A(n1472), .B(n1335), .Z(n1328) );
  XOR U1425 ( .A(n1324), .B(n1323), .Z(n1335) );
  XNOR U1426 ( .A(n1473), .B(n1320), .Z(n1323) );
  XOR U1427 ( .A(n1474), .B(n1475), .Z(n1320) );
  AND U1428 ( .A(n1476), .B(n1477), .Z(n1475) );
  XOR U1429 ( .A(n1474), .B(n1478), .Z(n1476) );
  XNOR U1430 ( .A(n1479), .B(n1480), .Z(n1473) );
  NOR U1431 ( .A(n1481), .B(n1482), .Z(n1480) );
  XNOR U1432 ( .A(n1479), .B(n1483), .Z(n1481) );
  XOR U1433 ( .A(n1484), .B(n1485), .Z(n1324) );
  NOR U1434 ( .A(n1486), .B(n1487), .Z(n1485) );
  XNOR U1435 ( .A(n1484), .B(n1488), .Z(n1486) );
  XNOR U1436 ( .A(n1334), .B(n1325), .Z(n1472) );
  XOR U1437 ( .A(n1489), .B(n1490), .Z(n1325) );
  NOR U1438 ( .A(n1491), .B(n1492), .Z(n1490) );
  XNOR U1439 ( .A(n1489), .B(n1493), .Z(n1491) );
  XOR U1440 ( .A(n1494), .B(n1340), .Z(n1334) );
  XNOR U1441 ( .A(n1495), .B(n1496), .Z(n1340) );
  NOR U1442 ( .A(n1497), .B(n1498), .Z(n1496) );
  XNOR U1443 ( .A(n1495), .B(n1499), .Z(n1497) );
  XNOR U1444 ( .A(n1339), .B(n1331), .Z(n1494) );
  XOR U1445 ( .A(n1500), .B(n1501), .Z(n1331) );
  AND U1446 ( .A(n1502), .B(n1503), .Z(n1501) );
  XOR U1447 ( .A(n1500), .B(n1504), .Z(n1502) );
  XNOR U1448 ( .A(n1505), .B(n1336), .Z(n1339) );
  XOR U1449 ( .A(n1506), .B(n1507), .Z(n1336) );
  AND U1450 ( .A(n1508), .B(n1509), .Z(n1507) );
  XOR U1451 ( .A(n1506), .B(n1510), .Z(n1508) );
  XNOR U1452 ( .A(n1511), .B(n1512), .Z(n1505) );
  NOR U1453 ( .A(n1513), .B(n1514), .Z(n1512) );
  XOR U1454 ( .A(n1511), .B(n1515), .Z(n1513) );
  AND U1455 ( .A(n1191), .B(n1193), .Z(n1341) );
  IV U1456 ( .A(n1172), .Z(n1193) );
  XOR U1457 ( .A(n1516), .B(n1392), .Z(n1172) );
  XNOR U1458 ( .A(n625), .B(p_input[128]), .Z(n1392) );
  IV U1459 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n625) );
  XOR U1460 ( .A(n1368), .B(n1367), .Z(n1516) );
  XOR U1461 ( .A(n1517), .B(n1379), .Z(n1367) );
  XOR U1462 ( .A(n1353), .B(n1351), .Z(n1379) );
  XOR U1463 ( .A(n1518), .B(n1358), .Z(n1351) );
  XNOR U1464 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .B(
        p_input[152]), .Z(n1358) );
  XOR U1465 ( .A(n1348), .B(n1357), .Z(n1518) );
  XNOR U1466 ( .A(n1519), .B(n1354), .Z(n1357) );
  XNOR U1467 ( .A(n383), .B(p_input[150]), .Z(n1354) );
  IV U1468 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .Z(n383) );
  XOR U1469 ( .A(n366), .B(p_input[151]), .Z(n1519) );
  IV U1470 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .Z(n366) );
  IV U1471 ( .A(n1352), .Z(n1348) );
  XOR U1472 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .B(
        p_input[146]), .Z(n1352) );
  XOR U1473 ( .A(n1363), .B(n1362), .Z(n1353) );
  XNOR U1474 ( .A(n1520), .B(n1359), .Z(n1362) );
  XNOR U1475 ( .A(n452), .B(p_input[147]), .Z(n1359) );
  IV U1476 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .Z(n452) );
  XOR U1477 ( .A(n418), .B(p_input[148]), .Z(n1520) );
  IV U1478 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .Z(n418) );
  XNOR U1479 ( .A(n400), .B(p_input[149]), .Z(n1363) );
  IV U1480 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .Z(n400) );
  XNOR U1481 ( .A(n1378), .B(n1364), .Z(n1517) );
  XNOR U1482 ( .A(n435), .B(p_input[129]), .Z(n1364) );
  IV U1483 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n435) );
  XNOR U1484 ( .A(n1521), .B(n1386), .Z(n1378) );
  XOR U1485 ( .A(n1374), .B(n1373), .Z(n1386) );
  XNOR U1486 ( .A(n1522), .B(n1370), .Z(n1373) );
  XNOR U1487 ( .A(n314), .B(p_input[154]), .Z(n1370) );
  IV U1488 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .Z(n314) );
  XOR U1489 ( .A(n297), .B(p_input[155]), .Z(n1522) );
  IV U1490 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .Z(n297) );
  XNOR U1491 ( .A(n279), .B(p_input[156]), .Z(n1374) );
  IV U1492 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .Z(n279) );
  XNOR U1493 ( .A(n1384), .B(n1375), .Z(n1521) );
  XNOR U1494 ( .A(n486), .B(p_input[145]), .Z(n1375) );
  IV U1495 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .Z(n486) );
  XOR U1496 ( .A(n1523), .B(n1391), .Z(n1384) );
  XNOR U1497 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .B(
        p_input[159]), .Z(n1391) );
  XOR U1498 ( .A(n1381), .B(n1390), .Z(n1523) );
  XNOR U1499 ( .A(n1524), .B(n1387), .Z(n1390) );
  XNOR U1500 ( .A(n262), .B(p_input[157]), .Z(n1387) );
  IV U1501 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .Z(n262) );
  XOR U1502 ( .A(n228), .B(p_input[158]), .Z(n1524) );
  IV U1503 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .Z(n228) );
  IV U1504 ( .A(n1385), .Z(n1381) );
  XOR U1505 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .B(
        p_input[153]), .Z(n1385) );
  XNOR U1506 ( .A(n1403), .B(n1402), .Z(n1368) );
  XNOR U1507 ( .A(n1525), .B(n1409), .Z(n1402) );
  XNOR U1508 ( .A(n1398), .B(n1397), .Z(n1409) );
  XOR U1509 ( .A(n1526), .B(n1394), .Z(n1397) );
  XOR U1510 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(
        p_input[139]), .Z(n1394) );
  XNOR U1511 ( .A(n574), .B(n1166), .Z(n1526) );
  IV U1512 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n574) );
  XOR U1513 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(
        p_input[141]), .Z(n1398) );
  XNOR U1514 ( .A(n1408), .B(n1399), .Z(n1525) );
  XNOR U1515 ( .A(n245), .B(p_input[130]), .Z(n1399) );
  IV U1516 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n245) );
  XOR U1517 ( .A(n1527), .B(n1414), .Z(n1408) );
  XNOR U1518 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .B(
        p_input[144]), .Z(n1414) );
  XNOR U1519 ( .A(n1405), .B(n1413), .Z(n1527) );
  XNOR U1520 ( .A(n1528), .B(n1410), .Z(n1413) );
  XNOR U1521 ( .A(n539), .B(p_input[142]), .Z(n1410) );
  IV U1522 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n539) );
  XOR U1523 ( .A(n522), .B(p_input[143]), .Z(n1528) );
  IV U1524 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .Z(n522) );
  XOR U1525 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(
        p_input[138]), .Z(n1405) );
  XNOR U1526 ( .A(n1421), .B(n1419), .Z(n1403) );
  XOR U1527 ( .A(n1529), .B(n1426), .Z(n1419) );
  XNOR U1528 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .B(
        p_input[137]), .Z(n1426) );
  XOR U1529 ( .A(n1416), .B(n1425), .Z(n1529) );
  XNOR U1530 ( .A(n1530), .B(n1422), .Z(n1425) );
  XOR U1531 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(
        p_input[135]), .Z(n1422) );
  XNOR U1532 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .B(
        p_input[136]), .Z(n1530) );
  IV U1533 ( .A(n1420), .Z(n1416) );
  XOR U1534 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .B(
        p_input[131]), .Z(n1420) );
  XOR U1535 ( .A(n1431), .B(n1430), .Z(n1421) );
  XNOR U1536 ( .A(n1531), .B(n1427), .Z(n1430) );
  XOR U1537 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(
        p_input[132]), .Z(n1427) );
  XNOR U1538 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(
        p_input[133]), .Z(n1531) );
  XOR U1539 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .B(
        p_input[134]), .Z(n1431) );
  XOR U1540 ( .A(n1532), .B(n1493), .Z(n1191) );
  XNOR U1541 ( .A(n1443), .B(n1442), .Z(n1493) );
  XNOR U1542 ( .A(n1533), .B(n1449), .Z(n1442) );
  XNOR U1543 ( .A(n1438), .B(n1437), .Z(n1449) );
  XOR U1544 ( .A(n1534), .B(n1434), .Z(n1437) );
  XOR U1545 ( .A(\knn_comb_/min_val_out[0][11] ), .B(p_input[139]), .Z(n1434)
         );
  XNOR U1546 ( .A(n567), .B(n1166), .Z(n1534) );
  IV U1547 ( .A(p_input[140]), .Z(n1166) );
  IV U1548 ( .A(\knn_comb_/min_val_out[0][12] ), .Z(n567) );
  XOR U1549 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[141]), .Z(n1438)
         );
  XNOR U1550 ( .A(n1448), .B(n1439), .Z(n1533) );
  XOR U1551 ( .A(\knn_comb_/min_val_out[0][2] ), .B(p_input[130]), .Z(n1439)
         );
  XOR U1552 ( .A(n1535), .B(n1454), .Z(n1448) );
  XOR U1553 ( .A(n497), .B(p_input[144]), .Z(n1454) );
  IV U1554 ( .A(\knn_comb_/min_val_out[0][16] ), .Z(n497) );
  XOR U1555 ( .A(n1445), .B(n1453), .Z(n1535) );
  XOR U1556 ( .A(n1536), .B(n1450), .Z(n1453) );
  XOR U1557 ( .A(\knn_comb_/min_val_out[0][14] ), .B(p_input[142]), .Z(n1450)
         );
  XOR U1558 ( .A(n515), .B(p_input[143]), .Z(n1536) );
  IV U1559 ( .A(\knn_comb_/min_val_out[0][15] ), .Z(n515) );
  XOR U1560 ( .A(\knn_comb_/min_val_out[0][10] ), .B(p_input[138]), .Z(n1445)
         );
  XNOR U1561 ( .A(n1460), .B(n1459), .Z(n1443) );
  XNOR U1562 ( .A(n1537), .B(n1465), .Z(n1459) );
  XOR U1563 ( .A(\knn_comb_/min_val_out[0][9] ), .B(p_input[137]), .Z(n1465)
         );
  XOR U1564 ( .A(n1456), .B(n1464), .Z(n1537) );
  XOR U1565 ( .A(n1538), .B(n1461), .Z(n1464) );
  XOR U1566 ( .A(\knn_comb_/min_val_out[0][7] ), .B(p_input[135]), .Z(n1461)
         );
  XNOR U1567 ( .A(\knn_comb_/min_val_out[0][8] ), .B(p_input[136]), .Z(n1538)
         );
  XOR U1568 ( .A(\knn_comb_/min_val_out[0][3] ), .B(p_input[131]), .Z(n1456)
         );
  XNOR U1569 ( .A(n1470), .B(n1469), .Z(n1460) );
  XOR U1570 ( .A(n1539), .B(n1466), .Z(n1469) );
  XOR U1571 ( .A(\knn_comb_/min_val_out[0][4] ), .B(p_input[132]), .Z(n1466)
         );
  XNOR U1572 ( .A(\knn_comb_/min_val_out[0][5] ), .B(p_input[133]), .Z(n1539)
         );
  XOR U1573 ( .A(\knn_comb_/min_val_out[0][6] ), .B(p_input[134]), .Z(n1470)
         );
  XOR U1574 ( .A(n1492), .B(n1471), .Z(n1532) );
  XOR U1575 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[128]), .Z(n1471)
         );
  XOR U1576 ( .A(n1540), .B(n1504), .Z(n1492) );
  XOR U1577 ( .A(n1478), .B(n1477), .Z(n1504) );
  XNOR U1578 ( .A(n1541), .B(n1483), .Z(n1477) );
  XOR U1579 ( .A(\knn_comb_/min_val_out[0][24] ), .B(p_input[152]), .Z(n1483)
         );
  XOR U1580 ( .A(n1474), .B(n1482), .Z(n1541) );
  XOR U1581 ( .A(n1542), .B(n1479), .Z(n1482) );
  XOR U1582 ( .A(\knn_comb_/min_val_out[0][22] ), .B(p_input[150]), .Z(n1479)
         );
  XOR U1583 ( .A(n359), .B(p_input[151]), .Z(n1542) );
  IV U1584 ( .A(\knn_comb_/min_val_out[0][23] ), .Z(n359) );
  XOR U1585 ( .A(\knn_comb_/min_val_out[0][18] ), .B(p_input[146]), .Z(n1474)
         );
  XNOR U1586 ( .A(n1488), .B(n1487), .Z(n1478) );
  XOR U1587 ( .A(n1543), .B(n1484), .Z(n1487) );
  XOR U1588 ( .A(\knn_comb_/min_val_out[0][19] ), .B(p_input[147]), .Z(n1484)
         );
  XOR U1589 ( .A(n411), .B(p_input[148]), .Z(n1543) );
  IV U1590 ( .A(\knn_comb_/min_val_out[0][20] ), .Z(n411) );
  XOR U1591 ( .A(\knn_comb_/min_val_out[0][21] ), .B(p_input[149]), .Z(n1488)
         );
  XNOR U1592 ( .A(n1503), .B(n1489), .Z(n1540) );
  XOR U1593 ( .A(\knn_comb_/min_val_out[0][1] ), .B(p_input[129]), .Z(n1489)
         );
  XNOR U1594 ( .A(n1544), .B(n1510), .Z(n1503) );
  XNOR U1595 ( .A(n1499), .B(n1498), .Z(n1510) );
  XOR U1596 ( .A(n1545), .B(n1495), .Z(n1498) );
  XOR U1597 ( .A(\knn_comb_/min_val_out[0][26] ), .B(p_input[154]), .Z(n1495)
         );
  XOR U1598 ( .A(n290), .B(p_input[155]), .Z(n1545) );
  IV U1599 ( .A(\knn_comb_/min_val_out[0][27] ), .Z(n290) );
  XOR U1600 ( .A(\knn_comb_/min_val_out[0][28] ), .B(p_input[156]), .Z(n1499)
         );
  XNOR U1601 ( .A(n1509), .B(n1500), .Z(n1544) );
  XOR U1602 ( .A(\knn_comb_/min_val_out[0][17] ), .B(p_input[145]), .Z(n1500)
         );
  XOR U1603 ( .A(n1546), .B(n1515), .Z(n1509) );
  XOR U1604 ( .A(n203), .B(p_input[159]), .Z(n1515) );
  IV U1605 ( .A(\knn_comb_/min_val_out[0][31] ), .Z(n203) );
  XOR U1606 ( .A(n1506), .B(n1514), .Z(n1546) );
  XOR U1607 ( .A(n1547), .B(n1511), .Z(n1514) );
  XOR U1608 ( .A(\knn_comb_/min_val_out[0][29] ), .B(p_input[157]), .Z(n1511)
         );
  XOR U1609 ( .A(n221), .B(p_input[158]), .Z(n1547) );
  IV U1610 ( .A(\knn_comb_/min_val_out[0][30] ), .Z(n221) );
  XOR U1611 ( .A(\knn_comb_/min_val_out[0][25] ), .B(p_input[153]), .Z(n1506)
         );
endmodule

