
module knn_comb_BMR_W16_K2_N64 ( p_input, o );
  input [1039:0] p_input;
  output [31:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][15] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604, n11605, n11606, n11607, n11608, n11609, n11610, n11611,
         n11612, n11613, n11614, n11615, n11616, n11617, n11618, n11619,
         n11620, n11621, n11622, n11623, n11624, n11625, n11626, n11627,
         n11628, n11629, n11630, n11631, n11632, n11633, n11634, n11635,
         n11636, n11637, n11638, n11639, n11640, n11641, n11642, n11643,
         n11644, n11645, n11646, n11647, n11648, n11649, n11650, n11651,
         n11652, n11653, n11654, n11655, n11656, n11657, n11658, n11659,
         n11660, n11661, n11662, n11663, n11664, n11665, n11666, n11667,
         n11668, n11669, n11670, n11671, n11672, n11673, n11674, n11675,
         n11676, n11677, n11678, n11679, n11680, n11681, n11682, n11683,
         n11684, n11685, n11686, n11687, n11688, n11689, n11690, n11691,
         n11692, n11693, n11694, n11695, n11696, n11697, n11698, n11699,
         n11700, n11701, n11702, n11703, n11704, n11705, n11706, n11707,
         n11708, n11709, n11710, n11711, n11712, n11713, n11714, n11715,
         n11716, n11717, n11718, n11719, n11720, n11721, n11722, n11723,
         n11724, n11725, n11726, n11727, n11728, n11729, n11730, n11731,
         n11732, n11733, n11734, n11735, n11736, n11737, n11738, n11739,
         n11740, n11741, n11742, n11743, n11744, n11745, n11746, n11747,
         n11748, n11749, n11750, n11751, n11752, n11753, n11754, n11755,
         n11756, n11757, n11758, n11759, n11760, n11761, n11762, n11763,
         n11764, n11765, n11766, n11767, n11768, n11769, n11770, n11771,
         n11772, n11773, n11774, n11775, n11776, n11777, n11778, n11779,
         n11780, n11781, n11782, n11783, n11784, n11785, n11786, n11787,
         n11788, n11789, n11790, n11791, n11792, n11793, n11794, n11795,
         n11796, n11797, n11798, n11799, n11800, n11801, n11802, n11803,
         n11804, n11805, n11806, n11807, n11808, n11809, n11810, n11811,
         n11812, n11813, n11814, n11815, n11816, n11817, n11818, n11819,
         n11820, n11821, n11822, n11823, n11824, n11825, n11826, n11827,
         n11828, n11829, n11830, n11831, n11832, n11833, n11834, n11835,
         n11836, n11837, n11838, n11839, n11840, n11841, n11842, n11843,
         n11844, n11845, n11846, n11847, n11848, n11849, n11850, n11851,
         n11852, n11853, n11854, n11855, n11856, n11857, n11858, n11859,
         n11860, n11861, n11862, n11863, n11864, n11865, n11866, n11867,
         n11868, n11869, n11870, n11871, n11872, n11873, n11874, n11875,
         n11876, n11877, n11878, n11879, n11880, n11881, n11882, n11883,
         n11884, n11885, n11886, n11887, n11888, n11889, n11890, n11891,
         n11892, n11893, n11894, n11895, n11896, n11897, n11898, n11899,
         n11900, n11901, n11902, n11903, n11904, n11905, n11906, n11907,
         n11908, n11909, n11910, n11911, n11912, n11913, n11914, n11915,
         n11916, n11917, n11918, n11919, n11920, n11921, n11922, n11923,
         n11924, n11925, n11926, n11927, n11928, n11929, n11930, n11931,
         n11932, n11933, n11934, n11935, n11936, n11937, n11938, n11939,
         n11940, n11941, n11942, n11943, n11944, n11945, n11946, n11947,
         n11948, n11949, n11950, n11951, n11952, n11953, n11954, n11955,
         n11956, n11957, n11958, n11959, n11960, n11961, n11962, n11963,
         n11964, n11965, n11966, n11967, n11968, n11969, n11970, n11971,
         n11972, n11973, n11974, n11975, n11976, n11977, n11978, n11979,
         n11980, n11981, n11982, n11983, n11984, n11985, n11986, n11987,
         n11988, n11989, n11990, n11991, n11992, n11993, n11994, n11995,
         n11996, n11997, n11998, n11999, n12000, n12001, n12002, n12003,
         n12004, n12005, n12006, n12007, n12008, n12009, n12010, n12011,
         n12012, n12013, n12014, n12015, n12016, n12017, n12018, n12019,
         n12020, n12021, n12022, n12023, n12024, n12025, n12026, n12027,
         n12028, n12029, n12030, n12031, n12032, n12033, n12034, n12035,
         n12036, n12037, n12038, n12039, n12040, n12041, n12042, n12043,
         n12044, n12045, n12046, n12047, n12048, n12049, n12050, n12051,
         n12052, n12053, n12054, n12055, n12056, n12057, n12058, n12059,
         n12060, n12061, n12062, n12063, n12064, n12065, n12066, n12067,
         n12068, n12069, n12070, n12071, n12072, n12073, n12074, n12075,
         n12076, n12077, n12078, n12079, n12080, n12081, n12082, n12083,
         n12084, n12085, n12086, n12087, n12088, n12089, n12090, n12091,
         n12092, n12093, n12094, n12095, n12096, n12097, n12098, n12099,
         n12100, n12101, n12102, n12103, n12104, n12105, n12106, n12107,
         n12108, n12109, n12110, n12111, n12112, n12113, n12114, n12115,
         n12116, n12117, n12118, n12119, n12120, n12121, n12122, n12123,
         n12124, n12125, n12126, n12127, n12128, n12129, n12130, n12131,
         n12132, n12133, n12134, n12135, n12136, n12137, n12138, n12139,
         n12140, n12141, n12142, n12143, n12144, n12145, n12146, n12147,
         n12148, n12149, n12150, n12151, n12152, n12153, n12154, n12155,
         n12156, n12157, n12158, n12159, n12160, n12161, n12162, n12163,
         n12164, n12165, n12166, n12167, n12168, n12169, n12170, n12171,
         n12172, n12173, n12174, n12175, n12176, n12177, n12178, n12179,
         n12180, n12181, n12182, n12183, n12184, n12185, n12186, n12187,
         n12188, n12189, n12190, n12191, n12192, n12193, n12194, n12195,
         n12196, n12197, n12198, n12199, n12200, n12201, n12202, n12203,
         n12204, n12205, n12206, n12207, n12208, n12209, n12210, n12211,
         n12212, n12213, n12214, n12215, n12216, n12217, n12218, n12219,
         n12220, n12221, n12222, n12223, n12224, n12225, n12226, n12227,
         n12228, n12229, n12230, n12231, n12232, n12233, n12234, n12235,
         n12236, n12237, n12238, n12239, n12240, n12241, n12242, n12243,
         n12244, n12245, n12246, n12247, n12248, n12249, n12250, n12251,
         n12252, n12253, n12254, n12255, n12256, n12257, n12258, n12259,
         n12260, n12261, n12262, n12263, n12264, n12265, n12266, n12267,
         n12268, n12269, n12270, n12271, n12272, n12273, n12274, n12275,
         n12276, n12277, n12278, n12279, n12280, n12281, n12282, n12283,
         n12284, n12285, n12286, n12287, n12288, n12289, n12290, n12291,
         n12292, n12293, n12294, n12295, n12296, n12297, n12298, n12299,
         n12300, n12301, n12302, n12303, n12304, n12305, n12306, n12307,
         n12308, n12309, n12310, n12311, n12312, n12313, n12314, n12315,
         n12316, n12317, n12318, n12319, n12320, n12321, n12322, n12323,
         n12324, n12325, n12326, n12327, n12328, n12329, n12330, n12331,
         n12332, n12333, n12334, n12335, n12336, n12337, n12338, n12339,
         n12340, n12341, n12342, n12343, n12344, n12345, n12346, n12347,
         n12348, n12349, n12350, n12351, n12352, n12353, n12354, n12355,
         n12356, n12357, n12358, n12359, n12360, n12361, n12362, n12363,
         n12364, n12365, n12366, n12367, n12368, n12369, n12370, n12371,
         n12372, n12373, n12374, n12375, n12376, n12377, n12378, n12379,
         n12380, n12381, n12382, n12383, n12384, n12385, n12386, n12387,
         n12388, n12389, n12390, n12391, n12392, n12393, n12394, n12395,
         n12396, n12397, n12398, n12399, n12400, n12401, n12402, n12403,
         n12404, n12405, n12406, n12407, n12408, n12409, n12410, n12411,
         n12412, n12413, n12414, n12415, n12416, n12417, n12418, n12419,
         n12420, n12421, n12422, n12423, n12424, n12425, n12426, n12427,
         n12428, n12429, n12430, n12431, n12432, n12433, n12434, n12435,
         n12436, n12437, n12438, n12439, n12440, n12441, n12442, n12443,
         n12444, n12445, n12446, n12447, n12448, n12449, n12450, n12451,
         n12452, n12453, n12454, n12455, n12456, n12457, n12458, n12459,
         n12460, n12461, n12462, n12463, n12464, n12465, n12466, n12467,
         n12468, n12469, n12470, n12471, n12472, n12473, n12474, n12475,
         n12476, n12477, n12478, n12479, n12480, n12481, n12482, n12483,
         n12484, n12485, n12486, n12487, n12488, n12489, n12490, n12491,
         n12492, n12493, n12494, n12495, n12496, n12497, n12498, n12499,
         n12500, n12501, n12502, n12503, n12504, n12505, n12506, n12507,
         n12508, n12509, n12510, n12511, n12512, n12513, n12514, n12515,
         n12516, n12517, n12518, n12519, n12520, n12521, n12522, n12523,
         n12524, n12525, n12526, n12527, n12528, n12529, n12530, n12531,
         n12532, n12533, n12534, n12535, n12536, n12537, n12538, n12539,
         n12540, n12541, n12542, n12543, n12544, n12545, n12546, n12547,
         n12548, n12549, n12550, n12551, n12552, n12553, n12554, n12555,
         n12556, n12557, n12558, n12559, n12560, n12561, n12562, n12563,
         n12564, n12565, n12566, n12567, n12568, n12569, n12570, n12571,
         n12572, n12573, n12574, n12575, n12576, n12577, n12578, n12579,
         n12580, n12581, n12582, n12583, n12584, n12585, n12586, n12587,
         n12588, n12589, n12590, n12591, n12592, n12593, n12594, n12595,
         n12596, n12597, n12598, n12599, n12600, n12601, n12602, n12603,
         n12604, n12605, n12606, n12607, n12608, n12609, n12610, n12611,
         n12612, n12613, n12614, n12615, n12616, n12617, n12618, n12619,
         n12620, n12621, n12622, n12623, n12624, n12625, n12626, n12627,
         n12628, n12629, n12630, n12631, n12632, n12633, n12634, n12635,
         n12636, n12637, n12638, n12639, n12640, n12641, n12642, n12643,
         n12644, n12645, n12646, n12647, n12648, n12649, n12650, n12651,
         n12652, n12653, n12654, n12655, n12656, n12657, n12658, n12659,
         n12660, n12661, n12662, n12663, n12664, n12665, n12666, n12667,
         n12668, n12669, n12670, n12671, n12672, n12673, n12674, n12675,
         n12676, n12677, n12678, n12679, n12680, n12681, n12682, n12683,
         n12684, n12685, n12686, n12687, n12688, n12689, n12690, n12691,
         n12692, n12693, n12694, n12695, n12696, n12697, n12698, n12699,
         n12700, n12701, n12702, n12703, n12704, n12705, n12706, n12707,
         n12708, n12709, n12710, n12711, n12712, n12713, n12714, n12715,
         n12716, n12717, n12718, n12719, n12720, n12721, n12722, n12723,
         n12724, n12725, n12726, n12727, n12728, n12729, n12730, n12731,
         n12732, n12733, n12734, n12735, n12736, n12737, n12738, n12739,
         n12740, n12741, n12742, n12743, n12744, n12745, n12746, n12747,
         n12748, n12749, n12750, n12751, n12752, n12753, n12754, n12755,
         n12756, n12757, n12758, n12759, n12760, n12761, n12762, n12763,
         n12764, n12765, n12766, n12767, n12768, n12769, n12770, n12771,
         n12772, n12773, n12774, n12775, n12776, n12777, n12778, n12779,
         n12780, n12781, n12782, n12783, n12784, n12785, n12786, n12787,
         n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, n12989, n12990, n12991, n12992, n12993, n12994, n12995,
         n12996, n12997, n12998, n12999, n13000, n13001, n13002, n13003,
         n13004, n13005, n13006, n13007, n13008, n13009, n13010, n13011,
         n13012, n13013, n13014, n13015, n13016, n13017, n13018, n13019,
         n13020, n13021, n13022, n13023, n13024, n13025, n13026, n13027,
         n13028, n13029, n13030, n13031, n13032, n13033, n13034, n13035,
         n13036, n13037, n13038, n13039, n13040, n13041, n13042, n13043,
         n13044, n13045, n13046, n13047, n13048, n13049, n13050, n13051,
         n13052, n13053, n13054, n13055, n13056, n13057, n13058, n13059,
         n13060, n13061, n13062, n13063, n13064, n13065, n13066, n13067,
         n13068, n13069, n13070, n13071, n13072, n13073, n13074, n13075,
         n13076, n13077, n13078, n13079, n13080, n13081, n13082, n13083,
         n13084, n13085, n13086, n13087, n13088, n13089, n13090, n13091,
         n13092, n13093, n13094, n13095, n13096, n13097, n13098, n13099,
         n13100, n13101, n13102, n13103, n13104, n13105, n13106, n13107,
         n13108, n13109, n13110, n13111, n13112, n13113, n13114, n13115,
         n13116, n13117, n13118, n13119, n13120, n13121, n13122, n13123,
         n13124, n13125, n13126, n13127, n13128, n13129, n13130, n13131,
         n13132, n13133, n13134, n13135, n13136, n13137, n13138, n13139,
         n13140, n13141, n13142, n13143, n13144, n13145, n13146, n13147,
         n13148, n13149, n13150, n13151, n13152, n13153, n13154, n13155,
         n13156, n13157, n13158, n13159, n13160, n13161, n13162, n13163,
         n13164, n13165, n13166, n13167, n13168, n13169, n13170, n13171,
         n13172, n13173, n13174, n13175, n13176, n13177, n13178, n13179,
         n13180, n13181, n13182, n13183, n13184, n13185, n13186, n13187,
         n13188, n13189, n13190, n13191, n13192, n13193, n13194, n13195,
         n13196, n13197, n13198, n13199, n13200, n13201, n13202, n13203,
         n13204, n13205, n13206, n13207, n13208, n13209, n13210, n13211,
         n13212, n13213, n13214, n13215, n13216, n13217, n13218, n13219,
         n13220, n13221, n13222, n13223, n13224, n13225, n13226, n13227,
         n13228, n13229, n13230, n13231, n13232, n13233, n13234, n13235,
         n13236, n13237, n13238, n13239, n13240, n13241, n13242, n13243,
         n13244, n13245, n13246, n13247, n13248, n13249, n13250, n13251,
         n13252, n13253, n13254, n13255, n13256, n13257, n13258, n13259,
         n13260, n13261, n13262, n13263, n13264, n13265, n13266, n13267,
         n13268, n13269, n13270, n13271, n13272, n13273, n13274, n13275,
         n13276, n13277, n13278, n13279, n13280, n13281, n13282, n13283,
         n13284, n13285, n13286, n13287, n13288, n13289, n13290, n13291,
         n13292, n13293, n13294, n13295, n13296, n13297, n13298, n13299,
         n13300, n13301, n13302, n13303, n13304, n13305, n13306, n13307,
         n13308, n13309, n13310, n13311, n13312, n13313, n13314, n13315,
         n13316, n13317, n13318, n13319, n13320, n13321, n13322, n13323,
         n13324, n13325, n13326, n13327, n13328, n13329, n13330, n13331,
         n13332, n13333, n13334, n13335, n13336, n13337, n13338, n13339,
         n13340, n13341, n13342, n13343, n13344, n13345, n13346, n13347,
         n13348, n13349, n13350, n13351, n13352, n13353, n13354, n13355,
         n13356, n13357, n13358, n13359, n13360, n13361, n13362, n13363,
         n13364, n13365, n13366, n13367, n13368, n13369, n13370, n13371,
         n13372, n13373, n13374, n13375, n13376, n13377, n13378, n13379,
         n13380, n13381, n13382, n13383, n13384, n13385, n13386, n13387,
         n13388, n13389, n13390, n13391, n13392, n13393, n13394, n13395,
         n13396, n13397, n13398, n13399, n13400, n13401, n13402, n13403,
         n13404, n13405, n13406, n13407, n13408, n13409, n13410, n13411,
         n13412, n13413, n13414, n13415, n13416, n13417, n13418, n13419,
         n13420, n13421, n13422, n13423, n13424, n13425, n13426, n13427,
         n13428, n13429, n13430, n13431, n13432, n13433, n13434, n13435,
         n13436, n13437, n13438, n13439, n13440, n13441, n13442, n13443,
         n13444, n13445, n13446, n13447, n13448, n13449, n13450, n13451,
         n13452, n13453, n13454, n13455, n13456, n13457, n13458, n13459,
         n13460, n13461, n13462, n13463, n13464, n13465, n13466, n13467,
         n13468, n13469, n13470, n13471, n13472, n13473, n13474, n13475,
         n13476, n13477, n13478, n13479, n13480, n13481, n13482, n13483,
         n13484, n13485, n13486, n13487, n13488, n13489, n13490, n13491,
         n13492, n13493, n13494, n13495, n13496, n13497, n13498, n13499,
         n13500, n13501, n13502, n13503, n13504, n13505, n13506, n13507,
         n13508, n13509, n13510, n13511, n13512, n13513, n13514, n13515,
         n13516, n13517, n13518, n13519, n13520, n13521, n13522, n13523,
         n13524, n13525, n13526, n13527, n13528, n13529, n13530, n13531,
         n13532, n13533, n13534, n13535, n13536, n13537, n13538, n13539,
         n13540, n13541, n13542, n13543, n13544, n13545, n13546, n13547,
         n13548, n13549, n13550, n13551, n13552, n13553, n13554, n13555,
         n13556, n13557, n13558, n13559, n13560, n13561, n13562, n13563,
         n13564, n13565, n13566, n13567, n13568, n13569, n13570, n13571,
         n13572, n13573, n13574, n13575, n13576, n13577, n13578, n13579,
         n13580, n13581, n13582, n13583, n13584, n13585, n13586, n13587,
         n13588, n13589, n13590, n13591, n13592, n13593, n13594, n13595,
         n13596, n13597, n13598, n13599, n13600, n13601, n13602, n13603,
         n13604, n13605, n13606, n13607, n13608, n13609, n13610, n13611,
         n13612, n13613, n13614, n13615, n13616, n13617, n13618, n13619,
         n13620, n13621, n13622, n13623, n13624, n13625, n13626, n13627,
         n13628, n13629, n13630, n13631, n13632, n13633, n13634, n13635,
         n13636, n13637, n13638, n13639, n13640, n13641, n13642, n13643,
         n13644, n13645, n13646, n13647, n13648, n13649, n13650, n13651,
         n13652, n13653, n13654, n13655, n13656, n13657, n13658, n13659,
         n13660, n13661, n13662, n13663, n13664, n13665, n13666, n13667,
         n13668, n13669, n13670, n13671, n13672, n13673, n13674, n13675,
         n13676, n13677, n13678, n13679, n13680, n13681, n13682, n13683,
         n13684, n13685, n13686, n13687, n13688, n13689, n13690, n13691,
         n13692, n13693, n13694, n13695, n13696, n13697, n13698, n13699,
         n13700, n13701, n13702, n13703, n13704, n13705, n13706, n13707,
         n13708, n13709, n13710, n13711, n13712, n13713, n13714, n13715,
         n13716, n13717, n13718, n13719, n13720, n13721, n13722, n13723,
         n13724, n13725, n13726, n13727, n13728, n13729, n13730, n13731,
         n13732, n13733, n13734, n13735, n13736, n13737, n13738, n13739,
         n13740, n13741, n13742, n13743, n13744, n13745, n13746, n13747,
         n13748, n13749, n13750, n13751, n13752, n13753, n13754, n13755,
         n13756, n13757, n13758, n13759, n13760, n13761, n13762, n13763,
         n13764, n13765, n13766, n13767, n13768, n13769, n13770, n13771,
         n13772, n13773, n13774, n13775, n13776, n13777, n13778, n13779,
         n13780, n13781, n13782, n13783, n13784, n13785, n13786, n13787,
         n13788, n13789, n13790, n13791, n13792, n13793, n13794, n13795,
         n13796, n13797, n13798, n13799, n13800, n13801, n13802, n13803,
         n13804, n13805, n13806, n13807, n13808, n13809, n13810, n13811,
         n13812, n13813, n13814, n13815, n13816, n13817, n13818, n13819,
         n13820, n13821, n13822, n13823, n13824, n13825, n13826, n13827,
         n13828, n13829, n13830, n13831, n13832, n13833, n13834, n13835,
         n13836, n13837, n13838, n13839, n13840, n13841, n13842, n13843,
         n13844, n13845, n13846, n13847, n13848, n13849, n13850, n13851,
         n13852, n13853, n13854, n13855, n13856, n13857, n13858, n13859,
         n13860, n13861, n13862, n13863, n13864, n13865, n13866, n13867,
         n13868, n13869, n13870, n13871, n13872, n13873, n13874, n13875,
         n13876, n13877, n13878, n13879, n13880, n13881, n13882, n13883,
         n13884, n13885, n13886, n13887, n13888, n13889, n13890, n13891,
         n13892, n13893, n13894, n13895, n13896, n13897, n13898, n13899,
         n13900, n13901, n13902, n13903, n13904, n13905, n13906, n13907,
         n13908, n13909, n13910, n13911, n13912, n13913, n13914, n13915,
         n13916, n13917, n13918, n13919, n13920, n13921, n13922, n13923,
         n13924, n13925, n13926, n13927, n13928, n13929, n13930, n13931,
         n13932, n13933, n13934, n13935, n13936, n13937, n13938, n13939,
         n13940, n13941, n13942, n13943, n13944, n13945, n13946, n13947,
         n13948, n13949, n13950, n13951, n13952, n13953, n13954, n13955,
         n13956, n13957, n13958, n13959, n13960, n13961, n13962, n13963,
         n13964, n13965, n13966, n13967, n13968, n13969, n13970, n13971,
         n13972, n13973, n13974, n13975, n13976, n13977, n13978, n13979,
         n13980, n13981, n13982, n13983, n13984, n13985, n13986, n13987,
         n13988, n13989, n13990, n13991, n13992, n13993, n13994, n13995,
         n13996, n13997, n13998, n13999, n14000, n14001, n14002, n14003,
         n14004, n14005, n14006, n14007, n14008, n14009, n14010, n14011,
         n14012, n14013, n14014, n14015, n14016, n14017, n14018, n14019,
         n14020, n14021, n14022, n14023, n14024, n14025, n14026, n14027,
         n14028, n14029, n14030, n14031, n14032, n14033, n14034, n14035,
         n14036, n14037, n14038, n14039, n14040, n14041, n14042, n14043,
         n14044, n14045, n14046, n14047, n14048, n14049, n14050, n14051,
         n14052, n14053, n14054, n14055, n14056, n14057, n14058, n14059,
         n14060, n14061, n14062, n14063, n14064, n14065, n14066, n14067,
         n14068, n14069, n14070, n14071, n14072, n14073, n14074, n14075,
         n14076, n14077, n14078, n14079, n14080, n14081, n14082, n14083,
         n14084, n14085, n14086, n14087, n14088, n14089, n14090, n14091,
         n14092, n14093, n14094, n14095, n14096, n14097, n14098, n14099,
         n14100, n14101, n14102, n14103, n14104, n14105, n14106, n14107,
         n14108, n14109, n14110, n14111, n14112, n14113, n14114, n14115,
         n14116, n14117, n14118, n14119, n14120, n14121, n14122, n14123,
         n14124, n14125, n14126, n14127, n14128, n14129, n14130, n14131,
         n14132, n14133, n14134, n14135, n14136, n14137, n14138, n14139,
         n14140, n14141, n14142, n14143, n14144, n14145, n14146, n14147,
         n14148, n14149, n14150, n14151, n14152, n14153, n14154, n14155,
         n14156, n14157, n14158, n14159, n14160, n14161, n14162, n14163,
         n14164, n14165, n14166, n14167, n14168, n14169, n14170, n14171,
         n14172, n14173, n14174, n14175, n14176, n14177, n14178, n14179,
         n14180, n14181, n14182, n14183, n14184, n14185, n14186, n14187,
         n14188, n14189, n14190, n14191, n14192, n14193, n14194, n14195,
         n14196, n14197, n14198, n14199, n14200, n14201, n14202, n14203,
         n14204, n14205, n14206, n14207, n14208, n14209, n14210, n14211,
         n14212, n14213, n14214, n14215, n14216, n14217, n14218, n14219,
         n14220, n14221, n14222, n14223, n14224, n14225, n14226, n14227,
         n14228, n14229, n14230, n14231, n14232, n14233, n14234, n14235,
         n14236, n14237, n14238, n14239, n14240, n14241, n14242, n14243,
         n14244, n14245, n14246, n14247, n14248, n14249, n14250, n14251,
         n14252, n14253, n14254, n14255, n14256, n14257, n14258, n14259,
         n14260, n14261, n14262, n14263, n14264, n14265, n14266, n14267,
         n14268, n14269, n14270, n14271, n14272, n14273, n14274, n14275,
         n14276, n14277, n14278, n14279, n14280, n14281, n14282, n14283,
         n14284, n14285, n14286, n14287, n14288, n14289, n14290, n14291,
         n14292, n14293, n14294, n14295, n14296, n14297, n14298, n14299,
         n14300, n14301, n14302, n14303, n14304, n14305, n14306, n14307,
         n14308, n14309, n14310, n14311, n14312, n14313, n14314, n14315,
         n14316, n14317, n14318, n14319, n14320, n14321, n14322, n14323,
         n14324, n14325, n14326, n14327, n14328, n14329, n14330, n14331,
         n14332, n14333, n14334, n14335, n14336, n14337, n14338, n14339,
         n14340, n14341, n14342, n14343, n14344, n14345, n14346, n14347,
         n14348, n14349, n14350, n14351, n14352, n14353, n14354, n14355,
         n14356, n14357, n14358, n14359, n14360, n14361, n14362, n14363,
         n14364, n14365, n14366, n14367, n14368, n14369, n14370, n14371,
         n14372, n14373, n14374, n14375, n14376, n14377, n14378, n14379,
         n14380, n14381, n14382, n14383, n14384, n14385, n14386, n14387,
         n14388, n14389, n14390, n14391, n14392, n14393, n14394, n14395,
         n14396, n14397, n14398, n14399, n14400, n14401, n14402, n14403,
         n14404, n14405, n14406, n14407, n14408, n14409, n14410, n14411,
         n14412, n14413, n14414, n14415, n14416, n14417, n14418, n14419,
         n14420, n14421, n14422, n14423, n14424, n14425, n14426, n14427,
         n14428, n14429, n14430, n14431, n14432, n14433, n14434, n14435,
         n14436, n14437, n14438, n14439, n14440, n14441, n14442, n14443,
         n14444, n14445, n14446, n14447, n14448, n14449, n14450, n14451,
         n14452, n14453, n14454, n14455, n14456, n14457, n14458, n14459,
         n14460, n14461, n14462, n14463, n14464, n14465, n14466, n14467,
         n14468, n14469, n14470, n14471, n14472, n14473, n14474, n14475,
         n14476, n14477, n14478, n14479, n14480, n14481, n14482, n14483,
         n14484, n14485, n14486, n14487, n14488, n14489, n14490, n14491,
         n14492, n14493, n14494, n14495, n14496, n14497, n14498, n14499,
         n14500, n14501, n14502, n14503, n14504, n14505, n14506, n14507,
         n14508, n14509, n14510, n14511, n14512, n14513, n14514, n14515,
         n14516, n14517, n14518, n14519, n14520, n14521, n14522, n14523,
         n14524, n14525, n14526, n14527, n14528, n14529, n14530, n14531,
         n14532, n14533, n14534, n14535, n14536, n14537, n14538, n14539,
         n14540, n14541, n14542, n14543, n14544, n14545, n14546, n14547,
         n14548, n14549, n14550, n14551, n14552, n14553, n14554, n14555,
         n14556, n14557, n14558, n14559, n14560, n14561, n14562, n14563,
         n14564, n14565, n14566, n14567, n14568, n14569, n14570, n14571,
         n14572, n14573, n14574, n14575, n14576, n14577, n14578, n14579,
         n14580, n14581, n14582, n14583, n14584, n14585, n14586, n14587,
         n14588, n14589, n14590, n14591, n14592, n14593, n14594, n14595,
         n14596, n14597, n14598, n14599, n14600, n14601, n14602, n14603,
         n14604, n14605, n14606, n14607, n14608, n14609, n14610, n14611,
         n14612, n14613, n14614, n14615, n14616, n14617, n14618, n14619,
         n14620, n14621, n14622, n14623, n14624, n14625, n14626, n14627,
         n14628, n14629, n14630, n14631, n14632, n14633, n14634, n14635,
         n14636, n14637, n14638, n14639, n14640, n14641, n14642, n14643,
         n14644, n14645, n14646, n14647, n14648, n14649, n14650, n14651,
         n14652, n14653, n14654, n14655, n14656, n14657, n14658, n14659,
         n14660, n14661, n14662, n14663, n14664, n14665, n14666, n14667,
         n14668, n14669, n14670, n14671, n14672, n14673, n14674, n14675,
         n14676, n14677, n14678, n14679, n14680, n14681, n14682, n14683,
         n14684, n14685, n14686, n14687, n14688, n14689, n14690, n14691,
         n14692, n14693, n14694, n14695, n14696, n14697, n14698, n14699,
         n14700, n14701, n14702, n14703, n14704, n14705, n14706, n14707,
         n14708, n14709, n14710, n14711, n14712, n14713, n14714, n14715,
         n14716, n14717, n14718, n14719, n14720, n14721, n14722, n14723,
         n14724, n14725, n14726, n14727, n14728, n14729, n14730, n14731,
         n14732, n14733, n14734, n14735, n14736, n14737, n14738, n14739,
         n14740, n14741, n14742, n14743, n14744, n14745, n14746, n14747,
         n14748, n14749, n14750, n14751, n14752, n14753, n14754, n14755,
         n14756, n14757, n14758, n14759, n14760, n14761, n14762, n14763,
         n14764, n14765, n14766, n14767, n14768, n14769, n14770, n14771,
         n14772, n14773, n14774, n14775, n14776, n14777, n14778, n14779,
         n14780, n14781, n14782, n14783, n14784, n14785, n14786, n14787,
         n14788, n14789, n14790, n14791, n14792, n14793, n14794, n14795,
         n14796, n14797, n14798, n14799, n14800, n14801, n14802, n14803,
         n14804, n14805, n14806, n14807, n14808, n14809, n14810, n14811,
         n14812, n14813, n14814, n14815, n14816, n14817, n14818, n14819,
         n14820, n14821, n14822, n14823, n14824, n14825, n14826, n14827,
         n14828, n14829, n14830, n14831, n14832, n14833, n14834, n14835,
         n14836, n14837, n14838, n14839, n14840, n14841, n14842, n14843,
         n14844, n14845, n14846, n14847, n14848, n14849, n14850, n14851,
         n14852, n14853, n14854, n14855, n14856, n14857, n14858, n14859,
         n14860, n14861, n14862, n14863, n14864, n14865, n14866, n14867,
         n14868, n14869, n14870, n14871, n14872, n14873, n14874, n14875,
         n14876, n14877, n14878, n14879, n14880, n14881, n14882, n14883,
         n14884, n14885, n14886, n14887, n14888, n14889, n14890, n14891,
         n14892, n14893, n14894, n14895, n14896, n14897, n14898, n14899,
         n14900, n14901, n14902, n14903, n14904, n14905, n14906, n14907,
         n14908, n14909, n14910, n14911, n14912, n14913, n14914, n14915,
         n14916, n14917, n14918, n14919, n14920, n14921, n14922, n14923,
         n14924, n14925, n14926, n14927, n14928, n14929, n14930, n14931,
         n14932, n14933, n14934, n14935, n14936, n14937, n14938, n14939,
         n14940, n14941, n14942, n14943, n14944, n14945, n14946, n14947,
         n14948, n14949, n14950, n14951, n14952, n14953, n14954, n14955,
         n14956, n14957, n14958, n14959, n14960, n14961, n14962, n14963,
         n14964, n14965, n14966, n14967, n14968, n14969, n14970, n14971,
         n14972, n14973, n14974, n14975, n14976, n14977, n14978, n14979,
         n14980, n14981, n14982, n14983, n14984, n14985, n14986, n14987,
         n14988, n14989, n14990, n14991, n14992, n14993, n14994, n14995,
         n14996, n14997, n14998, n14999, n15000, n15001, n15002, n15003,
         n15004, n15005, n15006, n15007, n15008, n15009, n15010, n15011,
         n15012, n15013, n15014, n15015, n15016, n15017, n15018, n15019,
         n15020, n15021, n15022, n15023, n15024, n15025, n15026, n15027,
         n15028, n15029, n15030, n15031, n15032, n15033, n15034, n15035,
         n15036, n15037, n15038, n15039, n15040, n15041, n15042, n15043,
         n15044, n15045, n15046, n15047, n15048, n15049, n15050, n15051,
         n15052, n15053, n15054, n15055, n15056, n15057, n15058, n15059,
         n15060, n15061, n15062, n15063, n15064, n15065, n15066, n15067,
         n15068, n15069, n15070, n15071, n15072, n15073, n15074, n15075,
         n15076, n15077, n15078, n15079, n15080, n15081, n15082, n15083,
         n15084, n15085, n15086, n15087, n15088, n15089, n15090, n15091,
         n15092, n15093, n15094, n15095, n15096, n15097, n15098, n15099,
         n15100, n15101, n15102, n15103, n15104, n15105, n15106, n15107,
         n15108, n15109, n15110, n15111, n15112, n15113, n15114, n15115,
         n15116, n15117, n15118, n15119, n15120, n15121, n15122, n15123,
         n15124, n15125, n15126, n15127, n15128, n15129, n15130, n15131,
         n15132, n15133, n15134, n15135, n15136, n15137, n15138, n15139,
         n15140, n15141, n15142, n15143, n15144, n15145, n15146, n15147,
         n15148, n15149, n15150, n15151, n15152, n15153, n15154, n15155,
         n15156, n15157, n15158, n15159, n15160, n15161, n15162, n15163,
         n15164, n15165, n15166, n15167, n15168, n15169, n15170, n15171,
         n15172, n15173, n15174, n15175, n15176, n15177, n15178, n15179,
         n15180, n15181, n15182, n15183, n15184, n15185, n15186, n15187,
         n15188, n15189, n15190, n15191, n15192, n15193, n15194, n15195,
         n15196, n15197, n15198, n15199, n15200, n15201, n15202, n15203,
         n15204, n15205, n15206, n15207, n15208, n15209, n15210, n15211,
         n15212, n15213, n15214, n15215, n15216, n15217, n15218, n15219,
         n15220, n15221, n15222, n15223, n15224, n15225, n15226, n15227,
         n15228, n15229, n15230, n15231, n15232, n15233, n15234, n15235,
         n15236, n15237, n15238, n15239, n15240, n15241, n15242, n15243,
         n15244, n15245, n15246, n15247, n15248, n15249, n15250, n15251,
         n15252, n15253, n15254, n15255, n15256, n15257, n15258, n15259,
         n15260, n15261, n15262, n15263, n15264, n15265, n15266, n15267,
         n15268, n15269, n15270, n15271, n15272, n15273, n15274, n15275,
         n15276, n15277, n15278, n15279, n15280, n15281, n15282, n15283,
         n15284, n15285, n15286, n15287, n15288, n15289, n15290, n15291,
         n15292, n15293, n15294, n15295, n15296, n15297, n15298, n15299,
         n15300, n15301, n15302, n15303, n15304, n15305, n15306, n15307,
         n15308, n15309, n15310, n15311, n15312, n15313, n15314, n15315,
         n15316, n15317, n15318, n15319, n15320, n15321, n15322, n15323,
         n15324, n15325, n15326, n15327, n15328, n15329, n15330, n15331,
         n15332, n15333, n15334, n15335, n15336, n15337, n15338, n15339,
         n15340, n15341, n15342, n15343, n15344, n15345, n15346, n15347,
         n15348, n15349, n15350, n15351, n15352, n15353, n15354, n15355,
         n15356, n15357, n15358, n15359, n15360, n15361, n15362, n15363,
         n15364, n15365, n15366, n15367, n15368, n15369, n15370, n15371,
         n15372, n15373, n15374, n15375, n15376, n15377, n15378, n15379,
         n15380, n15381, n15382, n15383, n15384, n15385, n15386, n15387,
         n15388, n15389, n15390, n15391, n15392, n15393, n15394, n15395,
         n15396, n15397, n15398, n15399, n15400, n15401, n15402, n15403,
         n15404, n15405, n15406, n15407, n15408, n15409, n15410, n15411,
         n15412, n15413, n15414, n15415, n15416, n15417, n15418, n15419,
         n15420, n15421, n15422, n15423, n15424, n15425, n15426, n15427,
         n15428, n15429, n15430, n15431, n15432, n15433, n15434, n15435,
         n15436, n15437, n15438, n15439, n15440, n15441, n15442, n15443,
         n15444, n15445, n15446, n15447, n15448, n15449, n15450, n15451,
         n15452, n15453, n15454, n15455, n15456, n15457, n15458, n15459,
         n15460, n15461, n15462, n15463, n15464, n15465, n15466, n15467,
         n15468, n15469, n15470, n15471, n15472, n15473, n15474, n15475,
         n15476, n15477, n15478, n15479, n15480, n15481, n15482, n15483,
         n15484, n15485, n15486, n15487, n15488, n15489, n15490, n15491,
         n15492, n15493, n15494, n15495, n15496, n15497, n15498, n15499,
         n15500, n15501, n15502, n15503, n15504, n15505, n15506, n15507,
         n15508, n15509, n15510, n15511, n15512, n15513, n15514, n15515,
         n15516, n15517, n15518, n15519, n15520, n15521, n15522, n15523,
         n15524, n15525, n15526, n15527, n15528, n15529, n15530, n15531,
         n15532, n15533, n15534, n15535, n15536, n15537, n15538, n15539,
         n15540, n15541, n15542, n15543, n15544, n15545, n15546, n15547,
         n15548, n15549, n15550, n15551, n15552, n15553, n15554, n15555,
         n15556, n15557, n15558, n15559, n15560, n15561, n15562, n15563,
         n15564, n15565, n15566, n15567, n15568, n15569, n15570, n15571,
         n15572, n15573, n15574, n15575, n15576, n15577, n15578, n15579,
         n15580, n15581, n15582, n15583, n15584, n15585, n15586, n15587,
         n15588, n15589, n15590, n15591, n15592, n15593, n15594, n15595,
         n15596, n15597, n15598, n15599, n15600, n15601, n15602, n15603,
         n15604, n15605, n15606, n15607, n15608, n15609, n15610, n15611,
         n15612, n15613, n15614, n15615, n15616, n15617, n15618, n15619,
         n15620, n15621, n15622, n15623, n15624, n15625, n15626, n15627,
         n15628, n15629, n15630, n15631, n15632, n15633, n15634, n15635,
         n15636, n15637, n15638, n15639, n15640, n15641, n15642, n15643,
         n15644, n15645, n15646, n15647, n15648, n15649, n15650, n15651,
         n15652, n15653, n15654, n15655, n15656, n15657, n15658, n15659,
         n15660, n15661, n15662, n15663, n15664, n15665, n15666, n15667,
         n15668, n15669, n15670, n15671, n15672, n15673, n15674, n15675,
         n15676, n15677, n15678, n15679, n15680, n15681, n15682, n15683,
         n15684, n15685, n15686, n15687, n15688, n15689, n15690, n15691,
         n15692, n15693, n15694, n15695, n15696, n15697, n15698, n15699,
         n15700, n15701, n15702, n15703, n15704, n15705, n15706, n15707,
         n15708, n15709, n15710, n15711, n15712, n15713, n15714, n15715,
         n15716, n15717, n15718, n15719, n15720, n15721, n15722, n15723,
         n15724, n15725, n15726, n15727, n15728, n15729, n15730, n15731,
         n15732, n15733, n15734, n15735, n15736, n15737, n15738, n15739,
         n15740, n15741, n15742, n15743, n15744, n15745, n15746, n15747,
         n15748, n15749, n15750, n15751, n15752, n15753, n15754, n15755,
         n15756, n15757, n15758, n15759, n15760, n15761, n15762, n15763,
         n15764, n15765, n15766, n15767, n15768, n15769, n15770, n15771,
         n15772, n15773, n15774, n15775, n15776, n15777, n15778, n15779,
         n15780, n15781, n15782, n15783, n15784, n15785, n15786, n15787,
         n15788, n15789, n15790, n15791, n15792, n15793, n15794, n15795,
         n15796, n15797, n15798, n15799, n15800, n15801, n15802, n15803,
         n15804, n15805, n15806, n15807, n15808, n15809, n15810, n15811,
         n15812, n15813, n15814, n15815, n15816, n15817, n15818, n15819,
         n15820, n15821, n15822, n15823, n15824, n15825, n15826, n15827,
         n15828, n15829, n15830, n15831, n15832, n15833, n15834, n15835,
         n15836, n15837, n15838, n15839, n15840, n15841, n15842, n15843,
         n15844, n15845, n15846, n15847, n15848, n15849, n15850, n15851,
         n15852, n15853, n15854, n15855, n15856, n15857, n15858, n15859,
         n15860, n15861, n15862, n15863, n15864, n15865, n15866, n15867,
         n15868, n15869, n15870, n15871, n15872, n15873, n15874, n15875,
         n15876, n15877, n15878, n15879, n15880, n15881, n15882, n15883,
         n15884, n15885, n15886, n15887, n15888, n15889, n15890, n15891,
         n15892, n15893, n15894, n15895, n15896, n15897, n15898, n15899,
         n15900, n15901, n15902, n15903, n15904, n15905, n15906, n15907,
         n15908, n15909, n15910, n15911, n15912, n15913, n15914, n15915,
         n15916, n15917, n15918, n15919, n15920, n15921, n15922, n15923,
         n15924, n15925, n15926, n15927, n15928, n15929, n15930, n15931,
         n15932, n15933, n15934, n15935, n15936, n15937, n15938, n15939,
         n15940, n15941, n15942, n15943, n15944, n15945, n15946, n15947,
         n15948, n15949, n15950, n15951, n15952, n15953, n15954, n15955,
         n15956, n15957, n15958, n15959, n15960, n15961, n15962, n15963,
         n15964, n15965, n15966, n15967, n15968, n15969, n15970, n15971,
         n15972, n15973, n15974, n15975, n15976, n15977, n15978, n15979,
         n15980, n15981, n15982, n15983, n15984, n15985, n15986, n15987,
         n15988, n15989, n15990, n15991, n15992, n15993, n15994, n15995,
         n15996, n15997, n15998, n15999, n16000, n16001, n16002, n16003,
         n16004, n16005, n16006, n16007, n16008, n16009, n16010, n16011,
         n16012, n16013, n16014, n16015, n16016, n16017, n16018, n16019,
         n16020, n16021, n16022, n16023, n16024, n16025, n16026, n16027,
         n16028, n16029, n16030, n16031, n16032, n16033, n16034, n16035,
         n16036, n16037, n16038, n16039, n16040, n16041, n16042, n16043,
         n16044, n16045, n16046, n16047, n16048, n16049, n16050, n16051,
         n16052, n16053, n16054, n16055, n16056, n16057, n16058, n16059,
         n16060, n16061, n16062, n16063, n16064, n16065, n16066, n16067,
         n16068, n16069, n16070, n16071, n16072, n16073, n16074, n16075,
         n16076, n16077, n16078, n16079, n16080, n16081, n16082, n16083,
         n16084, n16085, n16086, n16087, n16088, n16089, n16090, n16091,
         n16092, n16093, n16094, n16095, n16096, n16097, n16098, n16099,
         n16100, n16101, n16102, n16103, n16104, n16105, n16106, n16107,
         n16108, n16109, n16110, n16111, n16112, n16113, n16114, n16115,
         n16116, n16117, n16118, n16119, n16120, n16121, n16122, n16123,
         n16124, n16125, n16126, n16127, n16128, n16129, n16130, n16131,
         n16132, n16133, n16134, n16135, n16136, n16137, n16138, n16139,
         n16140, n16141, n16142, n16143, n16144, n16145, n16146, n16147,
         n16148, n16149, n16150, n16151, n16152, n16153, n16154, n16155,
         n16156, n16157, n16158, n16159, n16160, n16161, n16162, n16163,
         n16164, n16165, n16166, n16167, n16168, n16169, n16170, n16171,
         n16172, n16173, n16174, n16175, n16176, n16177, n16178, n16179,
         n16180, n16181, n16182, n16183, n16184, n16185, n16186, n16187,
         n16188, n16189, n16190, n16191, n16192, n16193, n16194, n16195,
         n16196, n16197, n16198, n16199, n16200, n16201, n16202, n16203,
         n16204, n16205, n16206, n16207, n16208, n16209, n16210, n16211,
         n16212, n16213, n16214, n16215, n16216, n16217, n16218, n16219,
         n16220, n16221, n16222, n16223, n16224, n16225, n16226, n16227,
         n16228, n16229, n16230, n16231, n16232, n16233, n16234, n16235,
         n16236, n16237, n16238, n16239, n16240, n16241, n16242, n16243,
         n16244, n16245, n16246, n16247, n16248, n16249, n16250, n16251,
         n16252, n16253, n16254, n16255, n16256, n16257, n16258, n16259,
         n16260, n16261, n16262, n16263, n16264, n16265, n16266, n16267,
         n16268, n16269, n16270, n16271, n16272, n16273, n16274, n16275,
         n16276, n16277, n16278, n16279, n16280, n16281, n16282, n16283,
         n16284, n16285, n16286, n16287, n16288, n16289, n16290, n16291,
         n16292, n16293, n16294, n16295, n16296, n16297, n16298, n16299,
         n16300, n16301, n16302, n16303, n16304, n16305, n16306, n16307,
         n16308, n16309, n16310, n16311, n16312, n16313, n16314, n16315,
         n16316, n16317, n16318, n16319, n16320, n16321, n16322, n16323,
         n16324, n16325, n16326, n16327, n16328, n16329, n16330, n16331,
         n16332, n16333, n16334, n16335, n16336, n16337, n16338, n16339,
         n16340, n16341, n16342, n16343, n16344, n16345, n16346, n16347,
         n16348, n16349, n16350, n16351, n16352, n16353, n16354, n16355,
         n16356, n16357, n16358, n16359, n16360, n16361, n16362, n16363,
         n16364, n16365, n16366, n16367, n16368, n16369, n16370, n16371,
         n16372, n16373, n16374, n16375, n16376, n16377, n16378, n16379,
         n16380, n16381, n16382, n16383, n16384, n16385, n16386, n16387,
         n16388, n16389, n16390, n16391, n16392, n16393, n16394, n16395,
         n16396, n16397, n16398, n16399, n16400, n16401, n16402, n16403,
         n16404, n16405, n16406, n16407, n16408, n16409, n16410, n16411,
         n16412, n16413, n16414, n16415, n16416, n16417, n16418, n16419,
         n16420, n16421, n16422, n16423, n16424, n16425, n16426, n16427,
         n16428, n16429, n16430, n16431, n16432, n16433, n16434, n16435,
         n16436, n16437, n16438, n16439, n16440, n16441, n16442, n16443,
         n16444, n16445, n16446, n16447, n16448, n16449, n16450, n16451,
         n16452, n16453, n16454, n16455, n16456, n16457, n16458, n16459,
         n16460, n16461, n16462, n16463, n16464, n16465, n16466, n16467,
         n16468, n16469, n16470, n16471, n16472, n16473, n16474, n16475,
         n16476, n16477, n16478, n16479, n16480, n16481, n16482, n16483,
         n16484, n16485, n16486, n16487, n16488, n16489, n16490, n16491,
         n16492, n16493, n16494, n16495, n16496, n16497, n16498, n16499,
         n16500, n16501, n16502, n16503, n16504, n16505, n16506, n16507,
         n16508, n16509, n16510, n16511, n16512, n16513, n16514, n16515,
         n16516, n16517, n16518, n16519, n16520, n16521, n16522, n16523,
         n16524, n16525, n16526, n16527, n16528, n16529, n16530, n16531,
         n16532, n16533, n16534, n16535, n16536, n16537, n16538, n16539,
         n16540, n16541, n16542, n16543, n16544, n16545, n16546, n16547,
         n16548, n16549, n16550, n16551, n16552, n16553, n16554, n16555,
         n16556, n16557, n16558, n16559, n16560, n16561, n16562, n16563,
         n16564, n16565, n16566, n16567, n16568, n16569, n16570, n16571,
         n16572, n16573, n16574, n16575, n16576, n16577, n16578, n16579,
         n16580, n16581, n16582, n16583, n16584, n16585, n16586, n16587,
         n16588, n16589, n16590, n16591, n16592, n16593, n16594, n16595,
         n16596, n16597, n16598, n16599, n16600, n16601, n16602, n16603,
         n16604, n16605, n16606, n16607, n16608, n16609, n16610, n16611,
         n16612, n16613, n16614, n16615, n16616, n16617, n16618, n16619,
         n16620, n16621, n16622, n16623, n16624, n16625, n16626, n16627,
         n16628, n16629, n16630, n16631, n16632, n16633, n16634, n16635,
         n16636, n16637, n16638, n16639, n16640, n16641, n16642, n16643,
         n16644, n16645, n16646, n16647, n16648, n16649, n16650, n16651,
         n16652, n16653, n16654, n16655, n16656, n16657, n16658, n16659,
         n16660, n16661, n16662, n16663, n16664, n16665, n16666, n16667,
         n16668, n16669, n16670, n16671, n16672, n16673, n16674, n16675,
         n16676, n16677, n16678, n16679, n16680, n16681, n16682, n16683,
         n16684, n16685, n16686, n16687, n16688, n16689, n16690, n16691,
         n16692, n16693, n16694, n16695, n16696, n16697, n16698, n16699,
         n16700, n16701, n16702, n16703, n16704, n16705, n16706, n16707,
         n16708, n16709, n16710, n16711, n16712, n16713, n16714, n16715,
         n16716, n16717, n16718, n16719, n16720, n16721, n16722, n16723,
         n16724, n16725, n16726, n16727, n16728, n16729, n16730, n16731,
         n16732, n16733, n16734, n16735, n16736, n16737, n16738, n16739,
         n16740, n16741, n16742, n16743, n16744, n16745, n16746, n16747,
         n16748, n16749, n16750, n16751, n16752, n16753, n16754, n16755,
         n16756, n16757, n16758, n16759, n16760, n16761, n16762, n16763,
         n16764, n16765, n16766, n16767, n16768, n16769, n16770, n16771,
         n16772, n16773, n16774, n16775, n16776, n16777, n16778, n16779,
         n16780, n16781, n16782, n16783, n16784, n16785, n16786, n16787,
         n16788, n16789, n16790, n16791, n16792, n16793, n16794, n16795,
         n16796, n16797, n16798, n16799, n16800, n16801, n16802, n16803,
         n16804, n16805, n16806, n16807, n16808, n16809, n16810, n16811,
         n16812, n16813, n16814, n16815, n16816, n16817, n16818, n16819,
         n16820, n16821, n16822, n16823, n16824, n16825, n16826, n16827,
         n16828, n16829, n16830, n16831, n16832, n16833, n16834, n16835,
         n16836, n16837, n16838, n16839, n16840, n16841, n16842, n16843,
         n16844, n16845, n16846, n16847, n16848, n16849, n16850, n16851,
         n16852, n16853, n16854, n16855, n16856, n16857, n16858, n16859,
         n16860, n16861, n16862, n16863, n16864, n16865, n16866, n16867,
         n16868, n16869, n16870, n16871, n16872, n16873, n16874, n16875,
         n16876, n16877, n16878, n16879, n16880, n16881, n16882, n16883,
         n16884, n16885, n16886, n16887, n16888, n16889, n16890, n16891,
         n16892, n16893, n16894, n16895, n16896, n16897, n16898, n16899,
         n16900, n16901, n16902, n16903, n16904, n16905, n16906, n16907,
         n16908, n16909, n16910, n16911, n16912, n16913, n16914, n16915,
         n16916, n16917, n16918, n16919, n16920, n16921, n16922, n16923,
         n16924, n16925, n16926, n16927, n16928, n16929, n16930, n16931,
         n16932, n16933, n16934, n16935, n16936, n16937, n16938, n16939,
         n16940, n16941, n16942, n16943, n16944, n16945, n16946, n16947,
         n16948, n16949, n16950, n16951, n16952, n16953, n16954, n16955,
         n16956, n16957, n16958, n16959, n16960, n16961, n16962, n16963,
         n16964, n16965, n16966, n16967, n16968, n16969, n16970, n16971,
         n16972, n16973, n16974, n16975, n16976, n16977, n16978, n16979,
         n16980, n16981, n16982, n16983, n16984, n16985, n16986, n16987,
         n16988, n16989, n16990, n16991, n16992, n16993, n16994, n16995,
         n16996, n16997, n16998, n16999, n17000, n17001, n17002, n17003,
         n17004, n17005, n17006, n17007, n17008, n17009, n17010, n17011,
         n17012, n17013, n17014, n17015, n17016, n17017, n17018, n17019,
         n17020, n17021, n17022, n17023, n17024, n17025, n17026, n17027,
         n17028, n17029, n17030, n17031, n17032, n17033, n17034, n17035,
         n17036, n17037, n17038, n17039, n17040, n17041, n17042, n17043,
         n17044, n17045, n17046, n17047, n17048, n17049, n17050, n17051,
         n17052, n17053, n17054, n17055, n17056, n17057, n17058, n17059,
         n17060, n17061, n17062, n17063, n17064, n17065, n17066, n17067,
         n17068, n17069, n17070, n17071, n17072, n17073, n17074, n17075,
         n17076, n17077, n17078, n17079, n17080, n17081, n17082, n17083,
         n17084, n17085, n17086, n17087, n17088, n17089, n17090, n17091,
         n17092, n17093, n17094, n17095, n17096, n17097, n17098, n17099,
         n17100, n17101, n17102, n17103, n17104, n17105, n17106, n17107,
         n17108, n17109, n17110, n17111, n17112, n17113, n17114, n17115,
         n17116, n17117, n17118, n17119, n17120, n17121, n17122, n17123,
         n17124, n17125, n17126, n17127, n17128, n17129, n17130, n17131,
         n17132, n17133, n17134, n17135, n17136, n17137, n17138, n17139,
         n17140, n17141, n17142, n17143, n17144, n17145, n17146, n17147,
         n17148, n17149, n17150, n17151, n17152, n17153, n17154, n17155,
         n17156, n17157, n17158, n17159, n17160, n17161, n17162, n17163,
         n17164, n17165, n17166, n17167, n17168, n17169, n17170, n17171,
         n17172, n17173, n17174, n17175, n17176, n17177, n17178, n17179,
         n17180, n17181, n17182, n17183, n17184, n17185, n17186, n17187,
         n17188, n17189, n17190, n17191, n17192, n17193, n17194, n17195,
         n17196, n17197, n17198, n17199, n17200, n17201, n17202, n17203,
         n17204, n17205, n17206, n17207, n17208, n17209, n17210, n17211,
         n17212, n17213, n17214, n17215, n17216, n17217, n17218, n17219,
         n17220, n17221, n17222, n17223, n17224, n17225, n17226, n17227,
         n17228, n17229, n17230, n17231, n17232, n17233, n17234, n17235,
         n17236, n17237, n17238, n17239, n17240, n17241, n17242, n17243,
         n17244, n17245, n17246, n17247, n17248, n17249, n17250, n17251,
         n17252, n17253, n17254, n17255, n17256, n17257, n17258, n17259,
         n17260, n17261, n17262, n17263, n17264, n17265, n17266, n17267,
         n17268, n17269, n17270, n17271, n17272, n17273, n17274, n17275,
         n17276, n17277, n17278, n17279, n17280, n17281, n17282, n17283,
         n17284, n17285, n17286, n17287, n17288, n17289, n17290, n17291,
         n17292, n17293, n17294, n17295, n17296, n17297, n17298, n17299,
         n17300, n17301, n17302, n17303, n17304, n17305, n17306, n17307,
         n17308, n17309, n17310, n17311, n17312, n17313, n17314, n17315,
         n17316, n17317, n17318, n17319, n17320, n17321, n17322, n17323,
         n17324, n17325, n17326, n17327, n17328, n17329, n17330, n17331,
         n17332, n17333, n17334, n17335, n17336, n17337, n17338, n17339,
         n17340, n17341, n17342, n17343, n17344, n17345, n17346, n17347,
         n17348, n17349, n17350, n17351, n17352, n17353, n17354, n17355,
         n17356, n17357, n17358, n17359, n17360, n17361, n17362, n17363,
         n17364, n17365, n17366, n17367, n17368, n17369, n17370, n17371,
         n17372, n17373, n17374, n17375, n17376, n17377, n17378, n17379,
         n17380, n17381, n17382, n17383, n17384, n17385, n17386, n17387,
         n17388, n17389, n17390, n17391, n17392, n17393, n17394, n17395,
         n17396, n17397, n17398, n17399, n17400, n17401, n17402, n17403,
         n17404, n17405, n17406, n17407, n17408, n17409, n17410, n17411,
         n17412, n17413, n17414, n17415, n17416, n17417, n17418, n17419,
         n17420, n17421, n17422, n17423, n17424, n17425, n17426, n17427,
         n17428, n17429, n17430, n17431, n17432, n17433, n17434, n17435,
         n17436, n17437, n17438, n17439, n17440, n17441, n17442, n17443,
         n17444, n17445, n17446, n17447, n17448, n17449, n17450, n17451,
         n17452, n17453, n17454, n17455, n17456, n17457, n17458, n17459,
         n17460, n17461, n17462, n17463, n17464, n17465, n17466, n17467,
         n17468, n17469, n17470, n17471, n17472, n17473, n17474, n17475,
         n17476, n17477, n17478, n17479, n17480, n17481, n17482, n17483,
         n17484, n17485, n17486, n17487, n17488, n17489, n17490, n17491,
         n17492, n17493, n17494, n17495, n17496, n17497, n17498, n17499,
         n17500, n17501, n17502, n17503, n17504, n17505, n17506, n17507,
         n17508, n17509, n17510, n17511, n17512, n17513, n17514, n17515,
         n17516, n17517, n17518, n17519, n17520, n17521, n17522, n17523,
         n17524, n17525, n17526, n17527, n17528, n17529, n17530, n17531,
         n17532, n17533, n17534, n17535, n17536, n17537, n17538, n17539,
         n17540, n17541, n17542, n17543, n17544, n17545, n17546, n17547,
         n17548, n17549, n17550, n17551, n17552, n17553, n17554, n17555,
         n17556, n17557, n17558, n17559, n17560, n17561, n17562, n17563,
         n17564, n17565, n17566, n17567, n17568, n17569, n17570, n17571,
         n17572, n17573, n17574, n17575, n17576, n17577, n17578, n17579,
         n17580, n17581, n17582, n17583, n17584, n17585, n17586, n17587,
         n17588, n17589, n17590, n17591, n17592, n17593, n17594, n17595,
         n17596, n17597, n17598, n17599, n17600, n17601, n17602, n17603,
         n17604, n17605, n17606, n17607, n17608, n17609, n17610, n17611,
         n17612, n17613, n17614, n17615, n17616, n17617, n17618, n17619,
         n17620, n17621, n17622, n17623, n17624, n17625, n17626, n17627,
         n17628, n17629, n17630, n17631, n17632, n17633, n17634, n17635,
         n17636, n17637, n17638, n17639, n17640, n17641, n17642, n17643,
         n17644, n17645, n17646, n17647, n17648, n17649, n17650, n17651,
         n17652, n17653, n17654, n17655, n17656, n17657, n17658, n17659,
         n17660, n17661, n17662, n17663, n17664, n17665, n17666, n17667,
         n17668, n17669, n17670, n17671, n17672, n17673, n17674, n17675,
         n17676, n17677, n17678, n17679, n17680, n17681, n17682, n17683,
         n17684, n17685, n17686, n17687, n17688, n17689, n17690, n17691,
         n17692, n17693, n17694, n17695, n17696, n17697, n17698, n17699,
         n17700, n17701, n17702, n17703, n17704, n17705, n17706, n17707,
         n17708, n17709, n17710, n17711, n17712, n17713, n17714, n17715,
         n17716, n17717, n17718, n17719, n17720, n17721, n17722, n17723,
         n17724, n17725, n17726, n17727, n17728, n17729, n17730, n17731,
         n17732, n17733, n17734, n17735, n17736, n17737, n17738, n17739,
         n17740, n17741, n17742, n17743, n17744, n17745, n17746, n17747,
         n17748, n17749, n17750, n17751, n17752, n17753, n17754, n17755,
         n17756, n17757, n17758, n17759, n17760, n17761, n17762, n17763,
         n17764, n17765, n17766, n17767, n17768, n17769, n17770, n17771,
         n17772, n17773, n17774, n17775, n17776, n17777, n17778, n17779,
         n17780, n17781, n17782, n17783, n17784, n17785, n17786, n17787,
         n17788, n17789, n17790, n17791, n17792, n17793, n17794, n17795,
         n17796, n17797, n17798, n17799, n17800, n17801, n17802, n17803,
         n17804, n17805, n17806, n17807, n17808, n17809, n17810, n17811,
         n17812, n17813, n17814, n17815, n17816, n17817, n17818, n17819,
         n17820, n17821, n17822, n17823, n17824, n17825, n17826, n17827,
         n17828, n17829, n17830, n17831, n17832, n17833, n17834, n17835,
         n17836, n17837, n17838, n17839, n17840, n17841, n17842, n17843,
         n17844, n17845, n17846, n17847, n17848, n17849, n17850, n17851,
         n17852, n17853, n17854, n17855, n17856, n17857, n17858, n17859,
         n17860, n17861, n17862, n17863, n17864, n17865, n17866, n17867,
         n17868, n17869, n17870, n17871, n17872, n17873, n17874, n17875,
         n17876, n17877, n17878, n17879, n17880, n17881, n17882, n17883,
         n17884, n17885, n17886, n17887, n17888, n17889, n17890, n17891,
         n17892, n17893, n17894, n17895, n17896, n17897, n17898, n17899,
         n17900, n17901, n17902, n17903, n17904, n17905, n17906, n17907,
         n17908, n17909, n17910, n17911, n17912, n17913, n17914, n17915,
         n17916, n17917, n17918, n17919, n17920, n17921, n17922, n17923,
         n17924, n17925, n17926, n17927, n17928, n17929, n17930, n17931,
         n17932, n17933, n17934, n17935, n17936, n17937, n17938, n17939,
         n17940, n17941, n17942, n17943, n17944, n17945, n17946, n17947,
         n17948, n17949, n17950, n17951, n17952, n17953, n17954, n17955,
         n17956, n17957, n17958, n17959, n17960, n17961, n17962, n17963,
         n17964, n17965, n17966, n17967, n17968, n17969, n17970, n17971,
         n17972, n17973, n17974, n17975, n17976, n17977, n17978, n17979,
         n17980, n17981, n17982, n17983, n17984, n17985, n17986, n17987,
         n17988, n17989, n17990, n17991, n17992, n17993, n17994, n17995,
         n17996, n17997, n17998, n17999, n18000, n18001, n18002, n18003,
         n18004, n18005, n18006, n18007, n18008, n18009, n18010, n18011,
         n18012, n18013, n18014, n18015, n18016, n18017, n18018, n18019,
         n18020, n18021, n18022, n18023, n18024, n18025, n18026, n18027,
         n18028, n18029, n18030, n18031, n18032, n18033, n18034, n18035,
         n18036, n18037, n18038, n18039, n18040, n18041, n18042, n18043,
         n18044, n18045, n18046, n18047, n18048, n18049, n18050, n18051,
         n18052, n18053, n18054, n18055, n18056, n18057, n18058, n18059,
         n18060, n18061, n18062, n18063, n18064, n18065, n18066, n18067,
         n18068, n18069, n18070, n18071, n18072, n18073, n18074, n18075,
         n18076, n18077, n18078, n18079, n18080, n18081, n18082, n18083,
         n18084, n18085, n18086, n18087, n18088, n18089, n18090, n18091,
         n18092, n18093, n18094, n18095, n18096, n18097, n18098, n18099,
         n18100, n18101, n18102, n18103, n18104, n18105, n18106, n18107,
         n18108, n18109, n18110, n18111, n18112, n18113, n18114, n18115,
         n18116, n18117, n18118, n18119, n18120, n18121, n18122, n18123,
         n18124, n18125, n18126, n18127, n18128, n18129, n18130, n18131,
         n18132, n18133, n18134, n18135, n18136, n18137, n18138, n18139,
         n18140, n18141, n18142, n18143, n18144, n18145, n18146, n18147,
         n18148, n18149, n18150, n18151, n18152, n18153, n18154, n18155,
         n18156, n18157, n18158, n18159, n18160, n18161, n18162, n18163,
         n18164, n18165, n18166, n18167, n18168, n18169, n18170, n18171,
         n18172, n18173, n18174, n18175, n18176, n18177, n18178, n18179,
         n18180, n18181, n18182, n18183, n18184, n18185, n18186, n18187,
         n18188, n18189, n18190, n18191, n18192, n18193, n18194, n18195,
         n18196, n18197, n18198, n18199, n18200, n18201, n18202, n18203,
         n18204, n18205, n18206, n18207, n18208, n18209, n18210, n18211,
         n18212, n18213, n18214, n18215, n18216, n18217, n18218, n18219,
         n18220, n18221, n18222, n18223, n18224, n18225, n18226, n18227,
         n18228, n18229, n18230, n18231, n18232, n18233, n18234, n18235,
         n18236, n18237, n18238, n18239, n18240, n18241, n18242, n18243,
         n18244, n18245, n18246, n18247, n18248, n18249, n18250, n18251,
         n18252, n18253, n18254, n18255, n18256, n18257, n18258, n18259,
         n18260, n18261, n18262, n18263, n18264, n18265, n18266, n18267,
         n18268, n18269, n18270, n18271, n18272, n18273, n18274, n18275,
         n18276, n18277, n18278, n18279, n18280, n18281, n18282, n18283,
         n18284, n18285, n18286, n18287, n18288, n18289, n18290, n18291,
         n18292, n18293, n18294, n18295, n18296, n18297, n18298, n18299,
         n18300, n18301, n18302, n18303, n18304, n18305, n18306, n18307,
         n18308, n18309, n18310, n18311, n18312, n18313, n18314, n18315,
         n18316, n18317, n18318, n18319, n18320, n18321, n18322, n18323,
         n18324, n18325, n18326, n18327, n18328, n18329, n18330, n18331,
         n18332, n18333, n18334, n18335, n18336, n18337, n18338, n18339,
         n18340, n18341, n18342, n18343, n18344, n18345, n18346, n18347,
         n18348, n18349, n18350, n18351, n18352, n18353, n18354, n18355,
         n18356, n18357, n18358, n18359, n18360, n18361, n18362, n18363,
         n18364, n18365, n18366, n18367, n18368, n18369, n18370, n18371,
         n18372, n18373, n18374, n18375, n18376, n18377, n18378, n18379,
         n18380, n18381, n18382, n18383, n18384, n18385, n18386, n18387,
         n18388, n18389, n18390, n18391, n18392, n18393, n18394, n18395,
         n18396, n18397, n18398, n18399, n18400, n18401;
  assign \knn_comb_/min_val_out[0][0]  = p_input[1008];
  assign \knn_comb_/min_val_out[0][1]  = p_input[1009];
  assign \knn_comb_/min_val_out[0][2]  = p_input[1010];
  assign \knn_comb_/min_val_out[0][3]  = p_input[1011];
  assign \knn_comb_/min_val_out[0][4]  = p_input[1012];
  assign \knn_comb_/min_val_out[0][5]  = p_input[1013];
  assign \knn_comb_/min_val_out[0][6]  = p_input[1014];
  assign \knn_comb_/min_val_out[0][7]  = p_input[1015];
  assign \knn_comb_/min_val_out[0][8]  = p_input[1016];
  assign \knn_comb_/min_val_out[0][9]  = p_input[1017];
  assign \knn_comb_/min_val_out[0][10]  = p_input[1018];
  assign \knn_comb_/min_val_out[0][11]  = p_input[1019];
  assign \knn_comb_/min_val_out[0][12]  = p_input[1020];
  assign \knn_comb_/min_val_out[0][13]  = p_input[1021];
  assign \knn_comb_/min_val_out[0][14]  = p_input[1022];
  assign \knn_comb_/min_val_out[0][15]  = p_input[1023];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][0]  = p_input[992];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][1]  = p_input[993];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][2]  = p_input[994];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][3]  = p_input[995];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][4]  = p_input[996];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][5]  = p_input[997];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][6]  = p_input[998];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][7]  = p_input[999];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][8]  = p_input[1000];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][9]  = p_input[1001];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][10]  = p_input[1002];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][11]  = p_input[1003];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][12]  = p_input[1004];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][13]  = p_input[1005];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][14]  = p_input[1006];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][15]  = p_input[1007];

  XOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  XOR U2 ( .A(n3), .B(n4), .Z(o[8]) );
  XOR U3 ( .A(n5), .B(n6), .Z(o[7]) );
  XOR U4 ( .A(n7), .B(n8), .Z(o[6]) );
  XOR U5 ( .A(n9), .B(n10), .Z(o[5]) );
  XOR U6 ( .A(n11), .B(n12), .Z(o[4]) );
  XOR U7 ( .A(n13), .B(n14), .Z(o[3]) );
  XOR U8 ( .A(n15), .B(n16), .Z(o[31]) );
  XOR U9 ( .A(n17), .B(n18), .Z(o[30]) );
  XOR U10 ( .A(n19), .B(n20), .Z(o[2]) );
  XOR U11 ( .A(n21), .B(n22), .Z(o[29]) );
  XOR U12 ( .A(n23), .B(n24), .Z(o[28]) );
  XOR U13 ( .A(n25), .B(n26), .Z(o[27]) );
  XOR U14 ( .A(n27), .B(n28), .Z(o[26]) );
  XOR U15 ( .A(n1), .B(n29), .Z(o[25]) );
  AND U16 ( .A(n30), .B(n31), .Z(n1) );
  XOR U17 ( .A(n2), .B(n29), .Z(n31) );
  XOR U18 ( .A(n32), .B(n33), .Z(n29) );
  AND U19 ( .A(n34), .B(n35), .Z(n33) );
  XOR U20 ( .A(p_input[9]), .B(n32), .Z(n35) );
  XOR U21 ( .A(n36), .B(n37), .Z(n32) );
  AND U22 ( .A(n38), .B(n39), .Z(n37) );
  XOR U23 ( .A(n40), .B(n41), .Z(n2) );
  AND U24 ( .A(n42), .B(n39), .Z(n41) );
  XNOR U25 ( .A(n43), .B(n36), .Z(n39) );
  XOR U26 ( .A(n44), .B(n45), .Z(n36) );
  AND U27 ( .A(n46), .B(n47), .Z(n45) );
  XOR U28 ( .A(p_input[25]), .B(n44), .Z(n47) );
  XOR U29 ( .A(n48), .B(n49), .Z(n44) );
  AND U30 ( .A(n50), .B(n51), .Z(n49) );
  IV U31 ( .A(n40), .Z(n43) );
  XNOR U32 ( .A(n52), .B(n53), .Z(n40) );
  AND U33 ( .A(n54), .B(n51), .Z(n53) );
  XNOR U34 ( .A(n52), .B(n48), .Z(n51) );
  XOR U35 ( .A(n55), .B(n56), .Z(n48) );
  AND U36 ( .A(n57), .B(n58), .Z(n56) );
  XOR U37 ( .A(p_input[41]), .B(n55), .Z(n58) );
  XOR U38 ( .A(n59), .B(n60), .Z(n55) );
  AND U39 ( .A(n61), .B(n62), .Z(n60) );
  XOR U40 ( .A(n63), .B(n64), .Z(n52) );
  AND U41 ( .A(n65), .B(n62), .Z(n64) );
  XNOR U42 ( .A(n63), .B(n59), .Z(n62) );
  XOR U43 ( .A(n66), .B(n67), .Z(n59) );
  AND U44 ( .A(n68), .B(n69), .Z(n67) );
  XOR U45 ( .A(p_input[57]), .B(n66), .Z(n69) );
  XOR U46 ( .A(n70), .B(n71), .Z(n66) );
  AND U47 ( .A(n72), .B(n73), .Z(n71) );
  XOR U48 ( .A(n74), .B(n75), .Z(n63) );
  AND U49 ( .A(n76), .B(n73), .Z(n75) );
  XNOR U50 ( .A(n74), .B(n70), .Z(n73) );
  XOR U51 ( .A(n77), .B(n78), .Z(n70) );
  AND U52 ( .A(n79), .B(n80), .Z(n78) );
  XOR U53 ( .A(p_input[73]), .B(n77), .Z(n80) );
  XOR U54 ( .A(n81), .B(n82), .Z(n77) );
  AND U55 ( .A(n83), .B(n84), .Z(n82) );
  XOR U56 ( .A(n85), .B(n86), .Z(n74) );
  AND U57 ( .A(n87), .B(n84), .Z(n86) );
  XNOR U58 ( .A(n85), .B(n81), .Z(n84) );
  XOR U59 ( .A(n88), .B(n89), .Z(n81) );
  AND U60 ( .A(n90), .B(n91), .Z(n89) );
  XOR U61 ( .A(p_input[89]), .B(n88), .Z(n91) );
  XOR U62 ( .A(n92), .B(n93), .Z(n88) );
  AND U63 ( .A(n94), .B(n95), .Z(n93) );
  XOR U64 ( .A(n96), .B(n97), .Z(n85) );
  AND U65 ( .A(n98), .B(n95), .Z(n97) );
  XNOR U66 ( .A(n96), .B(n92), .Z(n95) );
  XOR U67 ( .A(n99), .B(n100), .Z(n92) );
  AND U68 ( .A(n101), .B(n102), .Z(n100) );
  XOR U69 ( .A(p_input[105]), .B(n99), .Z(n102) );
  XOR U70 ( .A(n103), .B(n104), .Z(n99) );
  AND U71 ( .A(n105), .B(n106), .Z(n104) );
  XOR U72 ( .A(n107), .B(n108), .Z(n96) );
  AND U73 ( .A(n109), .B(n106), .Z(n108) );
  XNOR U74 ( .A(n107), .B(n103), .Z(n106) );
  XOR U75 ( .A(n110), .B(n111), .Z(n103) );
  AND U76 ( .A(n112), .B(n113), .Z(n111) );
  XOR U77 ( .A(p_input[121]), .B(n110), .Z(n113) );
  XOR U78 ( .A(n114), .B(n115), .Z(n110) );
  AND U79 ( .A(n116), .B(n117), .Z(n115) );
  XOR U80 ( .A(n118), .B(n119), .Z(n107) );
  AND U81 ( .A(n120), .B(n117), .Z(n119) );
  XNOR U82 ( .A(n118), .B(n114), .Z(n117) );
  XOR U83 ( .A(n121), .B(n122), .Z(n114) );
  AND U84 ( .A(n123), .B(n124), .Z(n122) );
  XOR U85 ( .A(p_input[137]), .B(n121), .Z(n124) );
  XOR U86 ( .A(n125), .B(n126), .Z(n121) );
  AND U87 ( .A(n127), .B(n128), .Z(n126) );
  XOR U88 ( .A(n129), .B(n130), .Z(n118) );
  AND U89 ( .A(n131), .B(n128), .Z(n130) );
  XNOR U90 ( .A(n129), .B(n125), .Z(n128) );
  XOR U91 ( .A(n132), .B(n133), .Z(n125) );
  AND U92 ( .A(n134), .B(n135), .Z(n133) );
  XOR U93 ( .A(p_input[153]), .B(n132), .Z(n135) );
  XOR U94 ( .A(n136), .B(n137), .Z(n132) );
  AND U95 ( .A(n138), .B(n139), .Z(n137) );
  XOR U96 ( .A(n140), .B(n141), .Z(n129) );
  AND U97 ( .A(n142), .B(n139), .Z(n141) );
  XNOR U98 ( .A(n140), .B(n136), .Z(n139) );
  XOR U99 ( .A(n143), .B(n144), .Z(n136) );
  AND U100 ( .A(n145), .B(n146), .Z(n144) );
  XOR U101 ( .A(p_input[169]), .B(n143), .Z(n146) );
  XOR U102 ( .A(n147), .B(n148), .Z(n143) );
  AND U103 ( .A(n149), .B(n150), .Z(n148) );
  XOR U104 ( .A(n151), .B(n152), .Z(n140) );
  AND U105 ( .A(n153), .B(n150), .Z(n152) );
  XNOR U106 ( .A(n151), .B(n147), .Z(n150) );
  XOR U107 ( .A(n154), .B(n155), .Z(n147) );
  AND U108 ( .A(n156), .B(n157), .Z(n155) );
  XOR U109 ( .A(p_input[185]), .B(n154), .Z(n157) );
  XOR U110 ( .A(n158), .B(n159), .Z(n154) );
  AND U111 ( .A(n160), .B(n161), .Z(n159) );
  XOR U112 ( .A(n162), .B(n163), .Z(n151) );
  AND U113 ( .A(n164), .B(n161), .Z(n163) );
  XNOR U114 ( .A(n162), .B(n158), .Z(n161) );
  XOR U115 ( .A(n165), .B(n166), .Z(n158) );
  AND U116 ( .A(n167), .B(n168), .Z(n166) );
  XOR U117 ( .A(p_input[201]), .B(n165), .Z(n168) );
  XOR U118 ( .A(n169), .B(n170), .Z(n165) );
  AND U119 ( .A(n171), .B(n172), .Z(n170) );
  XOR U120 ( .A(n173), .B(n174), .Z(n162) );
  AND U121 ( .A(n175), .B(n172), .Z(n174) );
  XNOR U122 ( .A(n173), .B(n169), .Z(n172) );
  XOR U123 ( .A(n176), .B(n177), .Z(n169) );
  AND U124 ( .A(n178), .B(n179), .Z(n177) );
  XOR U125 ( .A(p_input[217]), .B(n176), .Z(n179) );
  XOR U126 ( .A(n180), .B(n181), .Z(n176) );
  AND U127 ( .A(n182), .B(n183), .Z(n181) );
  XOR U128 ( .A(n184), .B(n185), .Z(n173) );
  AND U129 ( .A(n186), .B(n183), .Z(n185) );
  XNOR U130 ( .A(n184), .B(n180), .Z(n183) );
  XOR U131 ( .A(n187), .B(n188), .Z(n180) );
  AND U132 ( .A(n189), .B(n190), .Z(n188) );
  XOR U133 ( .A(p_input[233]), .B(n187), .Z(n190) );
  XOR U134 ( .A(n191), .B(n192), .Z(n187) );
  AND U135 ( .A(n193), .B(n194), .Z(n192) );
  XOR U136 ( .A(n195), .B(n196), .Z(n184) );
  AND U137 ( .A(n197), .B(n194), .Z(n196) );
  XNOR U138 ( .A(n195), .B(n191), .Z(n194) );
  XOR U139 ( .A(n198), .B(n199), .Z(n191) );
  AND U140 ( .A(n200), .B(n201), .Z(n199) );
  XOR U141 ( .A(p_input[249]), .B(n198), .Z(n201) );
  XOR U142 ( .A(n202), .B(n203), .Z(n198) );
  AND U143 ( .A(n204), .B(n205), .Z(n203) );
  XOR U144 ( .A(n206), .B(n207), .Z(n195) );
  AND U145 ( .A(n208), .B(n205), .Z(n207) );
  XNOR U146 ( .A(n206), .B(n202), .Z(n205) );
  XOR U147 ( .A(n209), .B(n210), .Z(n202) );
  AND U148 ( .A(n211), .B(n212), .Z(n210) );
  XOR U149 ( .A(p_input[265]), .B(n209), .Z(n212) );
  XOR U150 ( .A(n213), .B(n214), .Z(n209) );
  AND U151 ( .A(n215), .B(n216), .Z(n214) );
  XOR U152 ( .A(n217), .B(n218), .Z(n206) );
  AND U153 ( .A(n219), .B(n216), .Z(n218) );
  XNOR U154 ( .A(n217), .B(n213), .Z(n216) );
  XOR U155 ( .A(n220), .B(n221), .Z(n213) );
  AND U156 ( .A(n222), .B(n223), .Z(n221) );
  XOR U157 ( .A(p_input[281]), .B(n220), .Z(n223) );
  XOR U158 ( .A(n224), .B(n225), .Z(n220) );
  AND U159 ( .A(n226), .B(n227), .Z(n225) );
  XOR U160 ( .A(n228), .B(n229), .Z(n217) );
  AND U161 ( .A(n230), .B(n227), .Z(n229) );
  XNOR U162 ( .A(n228), .B(n224), .Z(n227) );
  XOR U163 ( .A(n231), .B(n232), .Z(n224) );
  AND U164 ( .A(n233), .B(n234), .Z(n232) );
  XOR U165 ( .A(p_input[297]), .B(n231), .Z(n234) );
  XOR U166 ( .A(n235), .B(n236), .Z(n231) );
  AND U167 ( .A(n237), .B(n238), .Z(n236) );
  XOR U168 ( .A(n239), .B(n240), .Z(n228) );
  AND U169 ( .A(n241), .B(n238), .Z(n240) );
  XNOR U170 ( .A(n239), .B(n235), .Z(n238) );
  XOR U171 ( .A(n242), .B(n243), .Z(n235) );
  AND U172 ( .A(n244), .B(n245), .Z(n243) );
  XOR U173 ( .A(p_input[313]), .B(n242), .Z(n245) );
  XOR U174 ( .A(n246), .B(n247), .Z(n242) );
  AND U175 ( .A(n248), .B(n249), .Z(n247) );
  XOR U176 ( .A(n250), .B(n251), .Z(n239) );
  AND U177 ( .A(n252), .B(n249), .Z(n251) );
  XNOR U178 ( .A(n250), .B(n246), .Z(n249) );
  XOR U179 ( .A(n253), .B(n254), .Z(n246) );
  AND U180 ( .A(n255), .B(n256), .Z(n254) );
  XOR U181 ( .A(p_input[329]), .B(n253), .Z(n256) );
  XOR U182 ( .A(n257), .B(n258), .Z(n253) );
  AND U183 ( .A(n259), .B(n260), .Z(n258) );
  XOR U184 ( .A(n261), .B(n262), .Z(n250) );
  AND U185 ( .A(n263), .B(n260), .Z(n262) );
  XNOR U186 ( .A(n261), .B(n257), .Z(n260) );
  XOR U187 ( .A(n264), .B(n265), .Z(n257) );
  AND U188 ( .A(n266), .B(n267), .Z(n265) );
  XOR U189 ( .A(p_input[345]), .B(n264), .Z(n267) );
  XOR U190 ( .A(n268), .B(n269), .Z(n264) );
  AND U191 ( .A(n270), .B(n271), .Z(n269) );
  XOR U192 ( .A(n272), .B(n273), .Z(n261) );
  AND U193 ( .A(n274), .B(n271), .Z(n273) );
  XNOR U194 ( .A(n272), .B(n268), .Z(n271) );
  XOR U195 ( .A(n275), .B(n276), .Z(n268) );
  AND U196 ( .A(n277), .B(n278), .Z(n276) );
  XOR U197 ( .A(p_input[361]), .B(n275), .Z(n278) );
  XOR U198 ( .A(n279), .B(n280), .Z(n275) );
  AND U199 ( .A(n281), .B(n282), .Z(n280) );
  XOR U200 ( .A(n283), .B(n284), .Z(n272) );
  AND U201 ( .A(n285), .B(n282), .Z(n284) );
  XNOR U202 ( .A(n283), .B(n279), .Z(n282) );
  XOR U203 ( .A(n286), .B(n287), .Z(n279) );
  AND U204 ( .A(n288), .B(n289), .Z(n287) );
  XOR U205 ( .A(p_input[377]), .B(n286), .Z(n289) );
  XOR U206 ( .A(n290), .B(n291), .Z(n286) );
  AND U207 ( .A(n292), .B(n293), .Z(n291) );
  XOR U208 ( .A(n294), .B(n295), .Z(n283) );
  AND U209 ( .A(n296), .B(n293), .Z(n295) );
  XNOR U210 ( .A(n294), .B(n290), .Z(n293) );
  XOR U211 ( .A(n297), .B(n298), .Z(n290) );
  AND U212 ( .A(n299), .B(n300), .Z(n298) );
  XOR U213 ( .A(p_input[393]), .B(n297), .Z(n300) );
  XOR U214 ( .A(n301), .B(n302), .Z(n297) );
  AND U215 ( .A(n303), .B(n304), .Z(n302) );
  XOR U216 ( .A(n305), .B(n306), .Z(n294) );
  AND U217 ( .A(n307), .B(n304), .Z(n306) );
  XNOR U218 ( .A(n305), .B(n301), .Z(n304) );
  XOR U219 ( .A(n308), .B(n309), .Z(n301) );
  AND U220 ( .A(n310), .B(n311), .Z(n309) );
  XOR U221 ( .A(p_input[409]), .B(n308), .Z(n311) );
  XOR U222 ( .A(n312), .B(n313), .Z(n308) );
  AND U223 ( .A(n314), .B(n315), .Z(n313) );
  XOR U224 ( .A(n316), .B(n317), .Z(n305) );
  AND U225 ( .A(n318), .B(n315), .Z(n317) );
  XNOR U226 ( .A(n316), .B(n312), .Z(n315) );
  XOR U227 ( .A(n319), .B(n320), .Z(n312) );
  AND U228 ( .A(n321), .B(n322), .Z(n320) );
  XOR U229 ( .A(p_input[425]), .B(n319), .Z(n322) );
  XOR U230 ( .A(n323), .B(n324), .Z(n319) );
  AND U231 ( .A(n325), .B(n326), .Z(n324) );
  XOR U232 ( .A(n327), .B(n328), .Z(n316) );
  AND U233 ( .A(n329), .B(n326), .Z(n328) );
  XNOR U234 ( .A(n327), .B(n323), .Z(n326) );
  XOR U235 ( .A(n330), .B(n331), .Z(n323) );
  AND U236 ( .A(n332), .B(n333), .Z(n331) );
  XOR U237 ( .A(p_input[441]), .B(n330), .Z(n333) );
  XOR U238 ( .A(n334), .B(n335), .Z(n330) );
  AND U239 ( .A(n336), .B(n337), .Z(n335) );
  XOR U240 ( .A(n338), .B(n339), .Z(n327) );
  AND U241 ( .A(n340), .B(n337), .Z(n339) );
  XNOR U242 ( .A(n338), .B(n334), .Z(n337) );
  XOR U243 ( .A(n341), .B(n342), .Z(n334) );
  AND U244 ( .A(n343), .B(n344), .Z(n342) );
  XOR U245 ( .A(p_input[457]), .B(n341), .Z(n344) );
  XOR U246 ( .A(n345), .B(n346), .Z(n341) );
  AND U247 ( .A(n347), .B(n348), .Z(n346) );
  XOR U248 ( .A(n349), .B(n350), .Z(n338) );
  AND U249 ( .A(n351), .B(n348), .Z(n350) );
  XNOR U250 ( .A(n349), .B(n345), .Z(n348) );
  XOR U251 ( .A(n352), .B(n353), .Z(n345) );
  AND U252 ( .A(n354), .B(n355), .Z(n353) );
  XOR U253 ( .A(p_input[473]), .B(n352), .Z(n355) );
  XOR U254 ( .A(n356), .B(n357), .Z(n352) );
  AND U255 ( .A(n358), .B(n359), .Z(n357) );
  XOR U256 ( .A(n360), .B(n361), .Z(n349) );
  AND U257 ( .A(n362), .B(n359), .Z(n361) );
  XNOR U258 ( .A(n360), .B(n356), .Z(n359) );
  XOR U259 ( .A(n363), .B(n364), .Z(n356) );
  AND U260 ( .A(n365), .B(n366), .Z(n364) );
  XOR U261 ( .A(p_input[489]), .B(n363), .Z(n366) );
  XOR U262 ( .A(n367), .B(n368), .Z(n363) );
  AND U263 ( .A(n369), .B(n370), .Z(n368) );
  XOR U264 ( .A(n371), .B(n372), .Z(n360) );
  AND U265 ( .A(n373), .B(n370), .Z(n372) );
  XNOR U266 ( .A(n371), .B(n367), .Z(n370) );
  XOR U267 ( .A(n374), .B(n375), .Z(n367) );
  AND U268 ( .A(n376), .B(n377), .Z(n375) );
  XOR U269 ( .A(p_input[505]), .B(n374), .Z(n377) );
  XOR U270 ( .A(n378), .B(n379), .Z(n374) );
  AND U271 ( .A(n380), .B(n381), .Z(n379) );
  XOR U272 ( .A(n382), .B(n383), .Z(n371) );
  AND U273 ( .A(n384), .B(n381), .Z(n383) );
  XNOR U274 ( .A(n382), .B(n378), .Z(n381) );
  XOR U275 ( .A(n385), .B(n386), .Z(n378) );
  AND U276 ( .A(n387), .B(n388), .Z(n386) );
  XOR U277 ( .A(p_input[521]), .B(n385), .Z(n388) );
  XOR U278 ( .A(n389), .B(n390), .Z(n385) );
  AND U279 ( .A(n391), .B(n392), .Z(n390) );
  XOR U280 ( .A(n393), .B(n394), .Z(n382) );
  AND U281 ( .A(n395), .B(n392), .Z(n394) );
  XNOR U282 ( .A(n393), .B(n389), .Z(n392) );
  XOR U283 ( .A(n396), .B(n397), .Z(n389) );
  AND U284 ( .A(n398), .B(n399), .Z(n397) );
  XOR U285 ( .A(p_input[537]), .B(n396), .Z(n399) );
  XOR U286 ( .A(n400), .B(n401), .Z(n396) );
  AND U287 ( .A(n402), .B(n403), .Z(n401) );
  XOR U288 ( .A(n404), .B(n405), .Z(n393) );
  AND U289 ( .A(n406), .B(n403), .Z(n405) );
  XNOR U290 ( .A(n404), .B(n400), .Z(n403) );
  XOR U291 ( .A(n407), .B(n408), .Z(n400) );
  AND U292 ( .A(n409), .B(n410), .Z(n408) );
  XOR U293 ( .A(p_input[553]), .B(n407), .Z(n410) );
  XOR U294 ( .A(n411), .B(n412), .Z(n407) );
  AND U295 ( .A(n413), .B(n414), .Z(n412) );
  XOR U296 ( .A(n415), .B(n416), .Z(n404) );
  AND U297 ( .A(n417), .B(n414), .Z(n416) );
  XNOR U298 ( .A(n415), .B(n411), .Z(n414) );
  XOR U299 ( .A(n418), .B(n419), .Z(n411) );
  AND U300 ( .A(n420), .B(n421), .Z(n419) );
  XOR U301 ( .A(p_input[569]), .B(n418), .Z(n421) );
  XOR U302 ( .A(n422), .B(n423), .Z(n418) );
  AND U303 ( .A(n424), .B(n425), .Z(n423) );
  XOR U304 ( .A(n426), .B(n427), .Z(n415) );
  AND U305 ( .A(n428), .B(n425), .Z(n427) );
  XNOR U306 ( .A(n426), .B(n422), .Z(n425) );
  XOR U307 ( .A(n429), .B(n430), .Z(n422) );
  AND U308 ( .A(n431), .B(n432), .Z(n430) );
  XOR U309 ( .A(p_input[585]), .B(n429), .Z(n432) );
  XOR U310 ( .A(n433), .B(n434), .Z(n429) );
  AND U311 ( .A(n435), .B(n436), .Z(n434) );
  XOR U312 ( .A(n437), .B(n438), .Z(n426) );
  AND U313 ( .A(n439), .B(n436), .Z(n438) );
  XNOR U314 ( .A(n437), .B(n433), .Z(n436) );
  XOR U315 ( .A(n440), .B(n441), .Z(n433) );
  AND U316 ( .A(n442), .B(n443), .Z(n441) );
  XOR U317 ( .A(p_input[601]), .B(n440), .Z(n443) );
  XOR U318 ( .A(n444), .B(n445), .Z(n440) );
  AND U319 ( .A(n446), .B(n447), .Z(n445) );
  XOR U320 ( .A(n448), .B(n449), .Z(n437) );
  AND U321 ( .A(n450), .B(n447), .Z(n449) );
  XNOR U322 ( .A(n448), .B(n444), .Z(n447) );
  XOR U323 ( .A(n451), .B(n452), .Z(n444) );
  AND U324 ( .A(n453), .B(n454), .Z(n452) );
  XOR U325 ( .A(p_input[617]), .B(n451), .Z(n454) );
  XOR U326 ( .A(n455), .B(n456), .Z(n451) );
  AND U327 ( .A(n457), .B(n458), .Z(n456) );
  XOR U328 ( .A(n459), .B(n460), .Z(n448) );
  AND U329 ( .A(n461), .B(n458), .Z(n460) );
  XNOR U330 ( .A(n459), .B(n455), .Z(n458) );
  XOR U331 ( .A(n462), .B(n463), .Z(n455) );
  AND U332 ( .A(n464), .B(n465), .Z(n463) );
  XOR U333 ( .A(p_input[633]), .B(n462), .Z(n465) );
  XOR U334 ( .A(n466), .B(n467), .Z(n462) );
  AND U335 ( .A(n468), .B(n469), .Z(n467) );
  XOR U336 ( .A(n470), .B(n471), .Z(n459) );
  AND U337 ( .A(n472), .B(n469), .Z(n471) );
  XNOR U338 ( .A(n470), .B(n466), .Z(n469) );
  XOR U339 ( .A(n473), .B(n474), .Z(n466) );
  AND U340 ( .A(n475), .B(n476), .Z(n474) );
  XOR U341 ( .A(p_input[649]), .B(n473), .Z(n476) );
  XOR U342 ( .A(n477), .B(n478), .Z(n473) );
  AND U343 ( .A(n479), .B(n480), .Z(n478) );
  XOR U344 ( .A(n481), .B(n482), .Z(n470) );
  AND U345 ( .A(n483), .B(n480), .Z(n482) );
  XNOR U346 ( .A(n481), .B(n477), .Z(n480) );
  XOR U347 ( .A(n484), .B(n485), .Z(n477) );
  AND U348 ( .A(n486), .B(n487), .Z(n485) );
  XOR U349 ( .A(p_input[665]), .B(n484), .Z(n487) );
  XOR U350 ( .A(n488), .B(n489), .Z(n484) );
  AND U351 ( .A(n490), .B(n491), .Z(n489) );
  XOR U352 ( .A(n492), .B(n493), .Z(n481) );
  AND U353 ( .A(n494), .B(n491), .Z(n493) );
  XNOR U354 ( .A(n492), .B(n488), .Z(n491) );
  XOR U355 ( .A(n495), .B(n496), .Z(n488) );
  AND U356 ( .A(n497), .B(n498), .Z(n496) );
  XOR U357 ( .A(p_input[681]), .B(n495), .Z(n498) );
  XOR U358 ( .A(n499), .B(n500), .Z(n495) );
  AND U359 ( .A(n501), .B(n502), .Z(n500) );
  XOR U360 ( .A(n503), .B(n504), .Z(n492) );
  AND U361 ( .A(n505), .B(n502), .Z(n504) );
  XNOR U362 ( .A(n503), .B(n499), .Z(n502) );
  XOR U363 ( .A(n506), .B(n507), .Z(n499) );
  AND U364 ( .A(n508), .B(n509), .Z(n507) );
  XOR U365 ( .A(p_input[697]), .B(n506), .Z(n509) );
  XOR U366 ( .A(n510), .B(n511), .Z(n506) );
  AND U367 ( .A(n512), .B(n513), .Z(n511) );
  XOR U368 ( .A(n514), .B(n515), .Z(n503) );
  AND U369 ( .A(n516), .B(n513), .Z(n515) );
  XNOR U370 ( .A(n514), .B(n510), .Z(n513) );
  XOR U371 ( .A(n517), .B(n518), .Z(n510) );
  AND U372 ( .A(n519), .B(n520), .Z(n518) );
  XOR U373 ( .A(p_input[713]), .B(n517), .Z(n520) );
  XOR U374 ( .A(n521), .B(n522), .Z(n517) );
  AND U375 ( .A(n523), .B(n524), .Z(n522) );
  XOR U376 ( .A(n525), .B(n526), .Z(n514) );
  AND U377 ( .A(n527), .B(n524), .Z(n526) );
  XNOR U378 ( .A(n525), .B(n521), .Z(n524) );
  XOR U379 ( .A(n528), .B(n529), .Z(n521) );
  AND U380 ( .A(n530), .B(n531), .Z(n529) );
  XOR U381 ( .A(p_input[729]), .B(n528), .Z(n531) );
  XOR U382 ( .A(n532), .B(n533), .Z(n528) );
  AND U383 ( .A(n534), .B(n535), .Z(n533) );
  XOR U384 ( .A(n536), .B(n537), .Z(n525) );
  AND U385 ( .A(n538), .B(n535), .Z(n537) );
  XNOR U386 ( .A(n536), .B(n532), .Z(n535) );
  XOR U387 ( .A(n539), .B(n540), .Z(n532) );
  AND U388 ( .A(n541), .B(n542), .Z(n540) );
  XOR U389 ( .A(p_input[745]), .B(n539), .Z(n542) );
  XOR U390 ( .A(n543), .B(n544), .Z(n539) );
  AND U391 ( .A(n545), .B(n546), .Z(n544) );
  XOR U392 ( .A(n547), .B(n548), .Z(n536) );
  AND U393 ( .A(n549), .B(n546), .Z(n548) );
  XNOR U394 ( .A(n547), .B(n543), .Z(n546) );
  XOR U395 ( .A(n550), .B(n551), .Z(n543) );
  AND U396 ( .A(n552), .B(n553), .Z(n551) );
  XOR U397 ( .A(p_input[761]), .B(n550), .Z(n553) );
  XOR U398 ( .A(n554), .B(n555), .Z(n550) );
  AND U399 ( .A(n556), .B(n557), .Z(n555) );
  XOR U400 ( .A(n558), .B(n559), .Z(n547) );
  AND U401 ( .A(n560), .B(n557), .Z(n559) );
  XNOR U402 ( .A(n558), .B(n554), .Z(n557) );
  XOR U403 ( .A(n561), .B(n562), .Z(n554) );
  AND U404 ( .A(n563), .B(n564), .Z(n562) );
  XOR U405 ( .A(p_input[777]), .B(n561), .Z(n564) );
  XOR U406 ( .A(n565), .B(n566), .Z(n561) );
  AND U407 ( .A(n567), .B(n568), .Z(n566) );
  XOR U408 ( .A(n569), .B(n570), .Z(n558) );
  AND U409 ( .A(n571), .B(n568), .Z(n570) );
  XNOR U410 ( .A(n569), .B(n565), .Z(n568) );
  XOR U411 ( .A(n572), .B(n573), .Z(n565) );
  AND U412 ( .A(n574), .B(n575), .Z(n573) );
  XOR U413 ( .A(p_input[793]), .B(n572), .Z(n575) );
  XOR U414 ( .A(n576), .B(n577), .Z(n572) );
  AND U415 ( .A(n578), .B(n579), .Z(n577) );
  XOR U416 ( .A(n580), .B(n581), .Z(n569) );
  AND U417 ( .A(n582), .B(n579), .Z(n581) );
  XNOR U418 ( .A(n580), .B(n576), .Z(n579) );
  XOR U419 ( .A(n583), .B(n584), .Z(n576) );
  AND U420 ( .A(n585), .B(n586), .Z(n584) );
  XOR U421 ( .A(p_input[809]), .B(n583), .Z(n586) );
  XOR U422 ( .A(n587), .B(n588), .Z(n583) );
  AND U423 ( .A(n589), .B(n590), .Z(n588) );
  XOR U424 ( .A(n591), .B(n592), .Z(n580) );
  AND U425 ( .A(n593), .B(n590), .Z(n592) );
  XNOR U426 ( .A(n591), .B(n587), .Z(n590) );
  XOR U427 ( .A(n594), .B(n595), .Z(n587) );
  AND U428 ( .A(n596), .B(n597), .Z(n595) );
  XOR U429 ( .A(p_input[825]), .B(n594), .Z(n597) );
  XOR U430 ( .A(n598), .B(n599), .Z(n594) );
  AND U431 ( .A(n600), .B(n601), .Z(n599) );
  XOR U432 ( .A(n602), .B(n603), .Z(n591) );
  AND U433 ( .A(n604), .B(n601), .Z(n603) );
  XNOR U434 ( .A(n602), .B(n598), .Z(n601) );
  XOR U435 ( .A(n605), .B(n606), .Z(n598) );
  AND U436 ( .A(n607), .B(n608), .Z(n606) );
  XOR U437 ( .A(p_input[841]), .B(n605), .Z(n608) );
  XOR U438 ( .A(n609), .B(n610), .Z(n605) );
  AND U439 ( .A(n611), .B(n612), .Z(n610) );
  XOR U440 ( .A(n613), .B(n614), .Z(n602) );
  AND U441 ( .A(n615), .B(n612), .Z(n614) );
  XNOR U442 ( .A(n613), .B(n609), .Z(n612) );
  XOR U443 ( .A(n616), .B(n617), .Z(n609) );
  AND U444 ( .A(n618), .B(n619), .Z(n617) );
  XOR U445 ( .A(p_input[857]), .B(n616), .Z(n619) );
  XOR U446 ( .A(n620), .B(n621), .Z(n616) );
  AND U447 ( .A(n622), .B(n623), .Z(n621) );
  XOR U448 ( .A(n624), .B(n625), .Z(n613) );
  AND U449 ( .A(n626), .B(n623), .Z(n625) );
  XNOR U450 ( .A(n624), .B(n620), .Z(n623) );
  XOR U451 ( .A(n627), .B(n628), .Z(n620) );
  AND U452 ( .A(n629), .B(n630), .Z(n628) );
  XOR U453 ( .A(p_input[873]), .B(n627), .Z(n630) );
  XOR U454 ( .A(n631), .B(n632), .Z(n627) );
  AND U455 ( .A(n633), .B(n634), .Z(n632) );
  XOR U456 ( .A(n635), .B(n636), .Z(n624) );
  AND U457 ( .A(n637), .B(n634), .Z(n636) );
  XNOR U458 ( .A(n635), .B(n631), .Z(n634) );
  XOR U459 ( .A(n638), .B(n639), .Z(n631) );
  AND U460 ( .A(n640), .B(n641), .Z(n639) );
  XOR U461 ( .A(p_input[889]), .B(n638), .Z(n641) );
  XOR U462 ( .A(n642), .B(n643), .Z(n638) );
  AND U463 ( .A(n644), .B(n645), .Z(n643) );
  XOR U464 ( .A(n646), .B(n647), .Z(n635) );
  AND U465 ( .A(n648), .B(n645), .Z(n647) );
  XNOR U466 ( .A(n646), .B(n642), .Z(n645) );
  XOR U467 ( .A(n649), .B(n650), .Z(n642) );
  AND U468 ( .A(n651), .B(n652), .Z(n650) );
  XOR U469 ( .A(p_input[905]), .B(n649), .Z(n652) );
  XOR U470 ( .A(n653), .B(n654), .Z(n649) );
  AND U471 ( .A(n655), .B(n656), .Z(n654) );
  XOR U472 ( .A(n657), .B(n658), .Z(n646) );
  AND U473 ( .A(n659), .B(n656), .Z(n658) );
  XNOR U474 ( .A(n657), .B(n653), .Z(n656) );
  XOR U475 ( .A(n660), .B(n661), .Z(n653) );
  AND U476 ( .A(n662), .B(n663), .Z(n661) );
  XOR U477 ( .A(p_input[921]), .B(n660), .Z(n663) );
  XOR U478 ( .A(n664), .B(n665), .Z(n660) );
  AND U479 ( .A(n666), .B(n667), .Z(n665) );
  XOR U480 ( .A(n668), .B(n669), .Z(n657) );
  AND U481 ( .A(n670), .B(n667), .Z(n669) );
  XNOR U482 ( .A(n668), .B(n664), .Z(n667) );
  XOR U483 ( .A(n671), .B(n672), .Z(n664) );
  AND U484 ( .A(n673), .B(n674), .Z(n672) );
  XOR U485 ( .A(p_input[937]), .B(n671), .Z(n674) );
  XOR U486 ( .A(n675), .B(n676), .Z(n671) );
  AND U487 ( .A(n677), .B(n678), .Z(n676) );
  XOR U488 ( .A(n679), .B(n680), .Z(n668) );
  AND U489 ( .A(n681), .B(n678), .Z(n680) );
  XNOR U490 ( .A(n679), .B(n675), .Z(n678) );
  XOR U491 ( .A(n682), .B(n683), .Z(n675) );
  AND U492 ( .A(n684), .B(n685), .Z(n683) );
  XOR U493 ( .A(p_input[953]), .B(n682), .Z(n685) );
  XOR U494 ( .A(n686), .B(n687), .Z(n682) );
  AND U495 ( .A(n688), .B(n689), .Z(n687) );
  XOR U496 ( .A(n690), .B(n691), .Z(n679) );
  AND U497 ( .A(n692), .B(n689), .Z(n691) );
  XNOR U498 ( .A(n690), .B(n686), .Z(n689) );
  XOR U499 ( .A(n693), .B(n694), .Z(n686) );
  AND U500 ( .A(n695), .B(n696), .Z(n694) );
  XOR U501 ( .A(p_input[969]), .B(n693), .Z(n696) );
  XOR U502 ( .A(n697), .B(n698), .Z(n693) );
  AND U503 ( .A(n699), .B(n700), .Z(n698) );
  XOR U504 ( .A(n701), .B(n702), .Z(n690) );
  AND U505 ( .A(n703), .B(n700), .Z(n702) );
  XNOR U506 ( .A(n701), .B(n697), .Z(n700) );
  XOR U507 ( .A(n704), .B(n705), .Z(n697) );
  AND U508 ( .A(n706), .B(n707), .Z(n705) );
  XOR U509 ( .A(p_input[985]), .B(n704), .Z(n707) );
  XNOR U510 ( .A(n708), .B(n709), .Z(n704) );
  AND U511 ( .A(n710), .B(n711), .Z(n709) );
  XNOR U512 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n712), .Z(n701) );
  AND U513 ( .A(n713), .B(n711), .Z(n712) );
  XOR U514 ( .A(n714), .B(n708), .Z(n711) );
  XOR U515 ( .A(n3), .B(n715), .Z(o[24]) );
  AND U516 ( .A(n30), .B(n716), .Z(n3) );
  XOR U517 ( .A(n4), .B(n715), .Z(n716) );
  XOR U518 ( .A(n717), .B(n718), .Z(n715) );
  AND U519 ( .A(n34), .B(n719), .Z(n718) );
  XOR U520 ( .A(p_input[8]), .B(n717), .Z(n719) );
  XOR U521 ( .A(n720), .B(n721), .Z(n717) );
  AND U522 ( .A(n38), .B(n722), .Z(n721) );
  XOR U523 ( .A(n723), .B(n724), .Z(n4) );
  AND U524 ( .A(n42), .B(n722), .Z(n724) );
  XNOR U525 ( .A(n725), .B(n720), .Z(n722) );
  XOR U526 ( .A(n726), .B(n727), .Z(n720) );
  AND U527 ( .A(n46), .B(n728), .Z(n727) );
  XOR U528 ( .A(p_input[24]), .B(n726), .Z(n728) );
  XOR U529 ( .A(n729), .B(n730), .Z(n726) );
  AND U530 ( .A(n50), .B(n731), .Z(n730) );
  IV U531 ( .A(n723), .Z(n725) );
  XNOR U532 ( .A(n732), .B(n733), .Z(n723) );
  AND U533 ( .A(n54), .B(n731), .Z(n733) );
  XNOR U534 ( .A(n732), .B(n729), .Z(n731) );
  XOR U535 ( .A(n734), .B(n735), .Z(n729) );
  AND U536 ( .A(n57), .B(n736), .Z(n735) );
  XOR U537 ( .A(p_input[40]), .B(n734), .Z(n736) );
  XOR U538 ( .A(n737), .B(n738), .Z(n734) );
  AND U539 ( .A(n61), .B(n739), .Z(n738) );
  XOR U540 ( .A(n740), .B(n741), .Z(n732) );
  AND U541 ( .A(n65), .B(n739), .Z(n741) );
  XNOR U542 ( .A(n740), .B(n737), .Z(n739) );
  XOR U543 ( .A(n742), .B(n743), .Z(n737) );
  AND U544 ( .A(n68), .B(n744), .Z(n743) );
  XOR U545 ( .A(p_input[56]), .B(n742), .Z(n744) );
  XOR U546 ( .A(n745), .B(n746), .Z(n742) );
  AND U547 ( .A(n72), .B(n747), .Z(n746) );
  XOR U548 ( .A(n748), .B(n749), .Z(n740) );
  AND U549 ( .A(n76), .B(n747), .Z(n749) );
  XNOR U550 ( .A(n748), .B(n745), .Z(n747) );
  XOR U551 ( .A(n750), .B(n751), .Z(n745) );
  AND U552 ( .A(n79), .B(n752), .Z(n751) );
  XOR U553 ( .A(p_input[72]), .B(n750), .Z(n752) );
  XOR U554 ( .A(n753), .B(n754), .Z(n750) );
  AND U555 ( .A(n83), .B(n755), .Z(n754) );
  XOR U556 ( .A(n756), .B(n757), .Z(n748) );
  AND U557 ( .A(n87), .B(n755), .Z(n757) );
  XNOR U558 ( .A(n756), .B(n753), .Z(n755) );
  XOR U559 ( .A(n758), .B(n759), .Z(n753) );
  AND U560 ( .A(n90), .B(n760), .Z(n759) );
  XOR U561 ( .A(p_input[88]), .B(n758), .Z(n760) );
  XOR U562 ( .A(n761), .B(n762), .Z(n758) );
  AND U563 ( .A(n94), .B(n763), .Z(n762) );
  XOR U564 ( .A(n764), .B(n765), .Z(n756) );
  AND U565 ( .A(n98), .B(n763), .Z(n765) );
  XNOR U566 ( .A(n764), .B(n761), .Z(n763) );
  XOR U567 ( .A(n766), .B(n767), .Z(n761) );
  AND U568 ( .A(n101), .B(n768), .Z(n767) );
  XOR U569 ( .A(p_input[104]), .B(n766), .Z(n768) );
  XOR U570 ( .A(n769), .B(n770), .Z(n766) );
  AND U571 ( .A(n105), .B(n771), .Z(n770) );
  XOR U572 ( .A(n772), .B(n773), .Z(n764) );
  AND U573 ( .A(n109), .B(n771), .Z(n773) );
  XNOR U574 ( .A(n772), .B(n769), .Z(n771) );
  XOR U575 ( .A(n774), .B(n775), .Z(n769) );
  AND U576 ( .A(n112), .B(n776), .Z(n775) );
  XOR U577 ( .A(p_input[120]), .B(n774), .Z(n776) );
  XOR U578 ( .A(n777), .B(n778), .Z(n774) );
  AND U579 ( .A(n116), .B(n779), .Z(n778) );
  XOR U580 ( .A(n780), .B(n781), .Z(n772) );
  AND U581 ( .A(n120), .B(n779), .Z(n781) );
  XNOR U582 ( .A(n780), .B(n777), .Z(n779) );
  XOR U583 ( .A(n782), .B(n783), .Z(n777) );
  AND U584 ( .A(n123), .B(n784), .Z(n783) );
  XOR U585 ( .A(p_input[136]), .B(n782), .Z(n784) );
  XOR U586 ( .A(n785), .B(n786), .Z(n782) );
  AND U587 ( .A(n127), .B(n787), .Z(n786) );
  XOR U588 ( .A(n788), .B(n789), .Z(n780) );
  AND U589 ( .A(n131), .B(n787), .Z(n789) );
  XNOR U590 ( .A(n788), .B(n785), .Z(n787) );
  XOR U591 ( .A(n790), .B(n791), .Z(n785) );
  AND U592 ( .A(n134), .B(n792), .Z(n791) );
  XOR U593 ( .A(p_input[152]), .B(n790), .Z(n792) );
  XOR U594 ( .A(n793), .B(n794), .Z(n790) );
  AND U595 ( .A(n138), .B(n795), .Z(n794) );
  XOR U596 ( .A(n796), .B(n797), .Z(n788) );
  AND U597 ( .A(n142), .B(n795), .Z(n797) );
  XNOR U598 ( .A(n796), .B(n793), .Z(n795) );
  XOR U599 ( .A(n798), .B(n799), .Z(n793) );
  AND U600 ( .A(n145), .B(n800), .Z(n799) );
  XOR U601 ( .A(p_input[168]), .B(n798), .Z(n800) );
  XOR U602 ( .A(n801), .B(n802), .Z(n798) );
  AND U603 ( .A(n149), .B(n803), .Z(n802) );
  XOR U604 ( .A(n804), .B(n805), .Z(n796) );
  AND U605 ( .A(n153), .B(n803), .Z(n805) );
  XNOR U606 ( .A(n804), .B(n801), .Z(n803) );
  XOR U607 ( .A(n806), .B(n807), .Z(n801) );
  AND U608 ( .A(n156), .B(n808), .Z(n807) );
  XOR U609 ( .A(p_input[184]), .B(n806), .Z(n808) );
  XOR U610 ( .A(n809), .B(n810), .Z(n806) );
  AND U611 ( .A(n160), .B(n811), .Z(n810) );
  XOR U612 ( .A(n812), .B(n813), .Z(n804) );
  AND U613 ( .A(n164), .B(n811), .Z(n813) );
  XNOR U614 ( .A(n812), .B(n809), .Z(n811) );
  XOR U615 ( .A(n814), .B(n815), .Z(n809) );
  AND U616 ( .A(n167), .B(n816), .Z(n815) );
  XOR U617 ( .A(p_input[200]), .B(n814), .Z(n816) );
  XOR U618 ( .A(n817), .B(n818), .Z(n814) );
  AND U619 ( .A(n171), .B(n819), .Z(n818) );
  XOR U620 ( .A(n820), .B(n821), .Z(n812) );
  AND U621 ( .A(n175), .B(n819), .Z(n821) );
  XNOR U622 ( .A(n820), .B(n817), .Z(n819) );
  XOR U623 ( .A(n822), .B(n823), .Z(n817) );
  AND U624 ( .A(n178), .B(n824), .Z(n823) );
  XOR U625 ( .A(p_input[216]), .B(n822), .Z(n824) );
  XOR U626 ( .A(n825), .B(n826), .Z(n822) );
  AND U627 ( .A(n182), .B(n827), .Z(n826) );
  XOR U628 ( .A(n828), .B(n829), .Z(n820) );
  AND U629 ( .A(n186), .B(n827), .Z(n829) );
  XNOR U630 ( .A(n828), .B(n825), .Z(n827) );
  XOR U631 ( .A(n830), .B(n831), .Z(n825) );
  AND U632 ( .A(n189), .B(n832), .Z(n831) );
  XOR U633 ( .A(p_input[232]), .B(n830), .Z(n832) );
  XOR U634 ( .A(n833), .B(n834), .Z(n830) );
  AND U635 ( .A(n193), .B(n835), .Z(n834) );
  XOR U636 ( .A(n836), .B(n837), .Z(n828) );
  AND U637 ( .A(n197), .B(n835), .Z(n837) );
  XNOR U638 ( .A(n836), .B(n833), .Z(n835) );
  XOR U639 ( .A(n838), .B(n839), .Z(n833) );
  AND U640 ( .A(n200), .B(n840), .Z(n839) );
  XOR U641 ( .A(p_input[248]), .B(n838), .Z(n840) );
  XOR U642 ( .A(n841), .B(n842), .Z(n838) );
  AND U643 ( .A(n204), .B(n843), .Z(n842) );
  XOR U644 ( .A(n844), .B(n845), .Z(n836) );
  AND U645 ( .A(n208), .B(n843), .Z(n845) );
  XNOR U646 ( .A(n844), .B(n841), .Z(n843) );
  XOR U647 ( .A(n846), .B(n847), .Z(n841) );
  AND U648 ( .A(n211), .B(n848), .Z(n847) );
  XOR U649 ( .A(p_input[264]), .B(n846), .Z(n848) );
  XOR U650 ( .A(n849), .B(n850), .Z(n846) );
  AND U651 ( .A(n215), .B(n851), .Z(n850) );
  XOR U652 ( .A(n852), .B(n853), .Z(n844) );
  AND U653 ( .A(n219), .B(n851), .Z(n853) );
  XNOR U654 ( .A(n852), .B(n849), .Z(n851) );
  XOR U655 ( .A(n854), .B(n855), .Z(n849) );
  AND U656 ( .A(n222), .B(n856), .Z(n855) );
  XOR U657 ( .A(p_input[280]), .B(n854), .Z(n856) );
  XOR U658 ( .A(n857), .B(n858), .Z(n854) );
  AND U659 ( .A(n226), .B(n859), .Z(n858) );
  XOR U660 ( .A(n860), .B(n861), .Z(n852) );
  AND U661 ( .A(n230), .B(n859), .Z(n861) );
  XNOR U662 ( .A(n860), .B(n857), .Z(n859) );
  XOR U663 ( .A(n862), .B(n863), .Z(n857) );
  AND U664 ( .A(n233), .B(n864), .Z(n863) );
  XOR U665 ( .A(p_input[296]), .B(n862), .Z(n864) );
  XOR U666 ( .A(n865), .B(n866), .Z(n862) );
  AND U667 ( .A(n237), .B(n867), .Z(n866) );
  XOR U668 ( .A(n868), .B(n869), .Z(n860) );
  AND U669 ( .A(n241), .B(n867), .Z(n869) );
  XNOR U670 ( .A(n868), .B(n865), .Z(n867) );
  XOR U671 ( .A(n870), .B(n871), .Z(n865) );
  AND U672 ( .A(n244), .B(n872), .Z(n871) );
  XOR U673 ( .A(p_input[312]), .B(n870), .Z(n872) );
  XOR U674 ( .A(n873), .B(n874), .Z(n870) );
  AND U675 ( .A(n248), .B(n875), .Z(n874) );
  XOR U676 ( .A(n876), .B(n877), .Z(n868) );
  AND U677 ( .A(n252), .B(n875), .Z(n877) );
  XNOR U678 ( .A(n876), .B(n873), .Z(n875) );
  XOR U679 ( .A(n878), .B(n879), .Z(n873) );
  AND U680 ( .A(n255), .B(n880), .Z(n879) );
  XOR U681 ( .A(p_input[328]), .B(n878), .Z(n880) );
  XOR U682 ( .A(n881), .B(n882), .Z(n878) );
  AND U683 ( .A(n259), .B(n883), .Z(n882) );
  XOR U684 ( .A(n884), .B(n885), .Z(n876) );
  AND U685 ( .A(n263), .B(n883), .Z(n885) );
  XNOR U686 ( .A(n884), .B(n881), .Z(n883) );
  XOR U687 ( .A(n886), .B(n887), .Z(n881) );
  AND U688 ( .A(n266), .B(n888), .Z(n887) );
  XOR U689 ( .A(p_input[344]), .B(n886), .Z(n888) );
  XOR U690 ( .A(n889), .B(n890), .Z(n886) );
  AND U691 ( .A(n270), .B(n891), .Z(n890) );
  XOR U692 ( .A(n892), .B(n893), .Z(n884) );
  AND U693 ( .A(n274), .B(n891), .Z(n893) );
  XNOR U694 ( .A(n892), .B(n889), .Z(n891) );
  XOR U695 ( .A(n894), .B(n895), .Z(n889) );
  AND U696 ( .A(n277), .B(n896), .Z(n895) );
  XOR U697 ( .A(p_input[360]), .B(n894), .Z(n896) );
  XOR U698 ( .A(n897), .B(n898), .Z(n894) );
  AND U699 ( .A(n281), .B(n899), .Z(n898) );
  XOR U700 ( .A(n900), .B(n901), .Z(n892) );
  AND U701 ( .A(n285), .B(n899), .Z(n901) );
  XNOR U702 ( .A(n900), .B(n897), .Z(n899) );
  XOR U703 ( .A(n902), .B(n903), .Z(n897) );
  AND U704 ( .A(n288), .B(n904), .Z(n903) );
  XOR U705 ( .A(p_input[376]), .B(n902), .Z(n904) );
  XOR U706 ( .A(n905), .B(n906), .Z(n902) );
  AND U707 ( .A(n292), .B(n907), .Z(n906) );
  XOR U708 ( .A(n908), .B(n909), .Z(n900) );
  AND U709 ( .A(n296), .B(n907), .Z(n909) );
  XNOR U710 ( .A(n908), .B(n905), .Z(n907) );
  XOR U711 ( .A(n910), .B(n911), .Z(n905) );
  AND U712 ( .A(n299), .B(n912), .Z(n911) );
  XOR U713 ( .A(p_input[392]), .B(n910), .Z(n912) );
  XOR U714 ( .A(n913), .B(n914), .Z(n910) );
  AND U715 ( .A(n303), .B(n915), .Z(n914) );
  XOR U716 ( .A(n916), .B(n917), .Z(n908) );
  AND U717 ( .A(n307), .B(n915), .Z(n917) );
  XNOR U718 ( .A(n916), .B(n913), .Z(n915) );
  XOR U719 ( .A(n918), .B(n919), .Z(n913) );
  AND U720 ( .A(n310), .B(n920), .Z(n919) );
  XOR U721 ( .A(p_input[408]), .B(n918), .Z(n920) );
  XOR U722 ( .A(n921), .B(n922), .Z(n918) );
  AND U723 ( .A(n314), .B(n923), .Z(n922) );
  XOR U724 ( .A(n924), .B(n925), .Z(n916) );
  AND U725 ( .A(n318), .B(n923), .Z(n925) );
  XNOR U726 ( .A(n924), .B(n921), .Z(n923) );
  XOR U727 ( .A(n926), .B(n927), .Z(n921) );
  AND U728 ( .A(n321), .B(n928), .Z(n927) );
  XOR U729 ( .A(p_input[424]), .B(n926), .Z(n928) );
  XOR U730 ( .A(n929), .B(n930), .Z(n926) );
  AND U731 ( .A(n325), .B(n931), .Z(n930) );
  XOR U732 ( .A(n932), .B(n933), .Z(n924) );
  AND U733 ( .A(n329), .B(n931), .Z(n933) );
  XNOR U734 ( .A(n932), .B(n929), .Z(n931) );
  XOR U735 ( .A(n934), .B(n935), .Z(n929) );
  AND U736 ( .A(n332), .B(n936), .Z(n935) );
  XOR U737 ( .A(p_input[440]), .B(n934), .Z(n936) );
  XOR U738 ( .A(n937), .B(n938), .Z(n934) );
  AND U739 ( .A(n336), .B(n939), .Z(n938) );
  XOR U740 ( .A(n940), .B(n941), .Z(n932) );
  AND U741 ( .A(n340), .B(n939), .Z(n941) );
  XNOR U742 ( .A(n940), .B(n937), .Z(n939) );
  XOR U743 ( .A(n942), .B(n943), .Z(n937) );
  AND U744 ( .A(n343), .B(n944), .Z(n943) );
  XOR U745 ( .A(p_input[456]), .B(n942), .Z(n944) );
  XOR U746 ( .A(n945), .B(n946), .Z(n942) );
  AND U747 ( .A(n347), .B(n947), .Z(n946) );
  XOR U748 ( .A(n948), .B(n949), .Z(n940) );
  AND U749 ( .A(n351), .B(n947), .Z(n949) );
  XNOR U750 ( .A(n948), .B(n945), .Z(n947) );
  XOR U751 ( .A(n950), .B(n951), .Z(n945) );
  AND U752 ( .A(n354), .B(n952), .Z(n951) );
  XOR U753 ( .A(p_input[472]), .B(n950), .Z(n952) );
  XOR U754 ( .A(n953), .B(n954), .Z(n950) );
  AND U755 ( .A(n358), .B(n955), .Z(n954) );
  XOR U756 ( .A(n956), .B(n957), .Z(n948) );
  AND U757 ( .A(n362), .B(n955), .Z(n957) );
  XNOR U758 ( .A(n956), .B(n953), .Z(n955) );
  XOR U759 ( .A(n958), .B(n959), .Z(n953) );
  AND U760 ( .A(n365), .B(n960), .Z(n959) );
  XOR U761 ( .A(p_input[488]), .B(n958), .Z(n960) );
  XOR U762 ( .A(n961), .B(n962), .Z(n958) );
  AND U763 ( .A(n369), .B(n963), .Z(n962) );
  XOR U764 ( .A(n964), .B(n965), .Z(n956) );
  AND U765 ( .A(n373), .B(n963), .Z(n965) );
  XNOR U766 ( .A(n964), .B(n961), .Z(n963) );
  XOR U767 ( .A(n966), .B(n967), .Z(n961) );
  AND U768 ( .A(n376), .B(n968), .Z(n967) );
  XOR U769 ( .A(p_input[504]), .B(n966), .Z(n968) );
  XOR U770 ( .A(n969), .B(n970), .Z(n966) );
  AND U771 ( .A(n380), .B(n971), .Z(n970) );
  XOR U772 ( .A(n972), .B(n973), .Z(n964) );
  AND U773 ( .A(n384), .B(n971), .Z(n973) );
  XNOR U774 ( .A(n972), .B(n969), .Z(n971) );
  XOR U775 ( .A(n974), .B(n975), .Z(n969) );
  AND U776 ( .A(n387), .B(n976), .Z(n975) );
  XOR U777 ( .A(p_input[520]), .B(n974), .Z(n976) );
  XOR U778 ( .A(n977), .B(n978), .Z(n974) );
  AND U779 ( .A(n391), .B(n979), .Z(n978) );
  XOR U780 ( .A(n980), .B(n981), .Z(n972) );
  AND U781 ( .A(n395), .B(n979), .Z(n981) );
  XNOR U782 ( .A(n980), .B(n977), .Z(n979) );
  XOR U783 ( .A(n982), .B(n983), .Z(n977) );
  AND U784 ( .A(n398), .B(n984), .Z(n983) );
  XOR U785 ( .A(p_input[536]), .B(n982), .Z(n984) );
  XOR U786 ( .A(n985), .B(n986), .Z(n982) );
  AND U787 ( .A(n402), .B(n987), .Z(n986) );
  XOR U788 ( .A(n988), .B(n989), .Z(n980) );
  AND U789 ( .A(n406), .B(n987), .Z(n989) );
  XNOR U790 ( .A(n988), .B(n985), .Z(n987) );
  XOR U791 ( .A(n990), .B(n991), .Z(n985) );
  AND U792 ( .A(n409), .B(n992), .Z(n991) );
  XOR U793 ( .A(p_input[552]), .B(n990), .Z(n992) );
  XOR U794 ( .A(n993), .B(n994), .Z(n990) );
  AND U795 ( .A(n413), .B(n995), .Z(n994) );
  XOR U796 ( .A(n996), .B(n997), .Z(n988) );
  AND U797 ( .A(n417), .B(n995), .Z(n997) );
  XNOR U798 ( .A(n996), .B(n993), .Z(n995) );
  XOR U799 ( .A(n998), .B(n999), .Z(n993) );
  AND U800 ( .A(n420), .B(n1000), .Z(n999) );
  XOR U801 ( .A(p_input[568]), .B(n998), .Z(n1000) );
  XOR U802 ( .A(n1001), .B(n1002), .Z(n998) );
  AND U803 ( .A(n424), .B(n1003), .Z(n1002) );
  XOR U804 ( .A(n1004), .B(n1005), .Z(n996) );
  AND U805 ( .A(n428), .B(n1003), .Z(n1005) );
  XNOR U806 ( .A(n1004), .B(n1001), .Z(n1003) );
  XOR U807 ( .A(n1006), .B(n1007), .Z(n1001) );
  AND U808 ( .A(n431), .B(n1008), .Z(n1007) );
  XOR U809 ( .A(p_input[584]), .B(n1006), .Z(n1008) );
  XOR U810 ( .A(n1009), .B(n1010), .Z(n1006) );
  AND U811 ( .A(n435), .B(n1011), .Z(n1010) );
  XOR U812 ( .A(n1012), .B(n1013), .Z(n1004) );
  AND U813 ( .A(n439), .B(n1011), .Z(n1013) );
  XNOR U814 ( .A(n1012), .B(n1009), .Z(n1011) );
  XOR U815 ( .A(n1014), .B(n1015), .Z(n1009) );
  AND U816 ( .A(n442), .B(n1016), .Z(n1015) );
  XOR U817 ( .A(p_input[600]), .B(n1014), .Z(n1016) );
  XOR U818 ( .A(n1017), .B(n1018), .Z(n1014) );
  AND U819 ( .A(n446), .B(n1019), .Z(n1018) );
  XOR U820 ( .A(n1020), .B(n1021), .Z(n1012) );
  AND U821 ( .A(n450), .B(n1019), .Z(n1021) );
  XNOR U822 ( .A(n1020), .B(n1017), .Z(n1019) );
  XOR U823 ( .A(n1022), .B(n1023), .Z(n1017) );
  AND U824 ( .A(n453), .B(n1024), .Z(n1023) );
  XOR U825 ( .A(p_input[616]), .B(n1022), .Z(n1024) );
  XOR U826 ( .A(n1025), .B(n1026), .Z(n1022) );
  AND U827 ( .A(n457), .B(n1027), .Z(n1026) );
  XOR U828 ( .A(n1028), .B(n1029), .Z(n1020) );
  AND U829 ( .A(n461), .B(n1027), .Z(n1029) );
  XNOR U830 ( .A(n1028), .B(n1025), .Z(n1027) );
  XOR U831 ( .A(n1030), .B(n1031), .Z(n1025) );
  AND U832 ( .A(n464), .B(n1032), .Z(n1031) );
  XOR U833 ( .A(p_input[632]), .B(n1030), .Z(n1032) );
  XOR U834 ( .A(n1033), .B(n1034), .Z(n1030) );
  AND U835 ( .A(n468), .B(n1035), .Z(n1034) );
  XOR U836 ( .A(n1036), .B(n1037), .Z(n1028) );
  AND U837 ( .A(n472), .B(n1035), .Z(n1037) );
  XNOR U838 ( .A(n1036), .B(n1033), .Z(n1035) );
  XOR U839 ( .A(n1038), .B(n1039), .Z(n1033) );
  AND U840 ( .A(n475), .B(n1040), .Z(n1039) );
  XOR U841 ( .A(p_input[648]), .B(n1038), .Z(n1040) );
  XOR U842 ( .A(n1041), .B(n1042), .Z(n1038) );
  AND U843 ( .A(n479), .B(n1043), .Z(n1042) );
  XOR U844 ( .A(n1044), .B(n1045), .Z(n1036) );
  AND U845 ( .A(n483), .B(n1043), .Z(n1045) );
  XNOR U846 ( .A(n1044), .B(n1041), .Z(n1043) );
  XOR U847 ( .A(n1046), .B(n1047), .Z(n1041) );
  AND U848 ( .A(n486), .B(n1048), .Z(n1047) );
  XOR U849 ( .A(p_input[664]), .B(n1046), .Z(n1048) );
  XOR U850 ( .A(n1049), .B(n1050), .Z(n1046) );
  AND U851 ( .A(n490), .B(n1051), .Z(n1050) );
  XOR U852 ( .A(n1052), .B(n1053), .Z(n1044) );
  AND U853 ( .A(n494), .B(n1051), .Z(n1053) );
  XNOR U854 ( .A(n1052), .B(n1049), .Z(n1051) );
  XOR U855 ( .A(n1054), .B(n1055), .Z(n1049) );
  AND U856 ( .A(n497), .B(n1056), .Z(n1055) );
  XOR U857 ( .A(p_input[680]), .B(n1054), .Z(n1056) );
  XOR U858 ( .A(n1057), .B(n1058), .Z(n1054) );
  AND U859 ( .A(n501), .B(n1059), .Z(n1058) );
  XOR U860 ( .A(n1060), .B(n1061), .Z(n1052) );
  AND U861 ( .A(n505), .B(n1059), .Z(n1061) );
  XNOR U862 ( .A(n1060), .B(n1057), .Z(n1059) );
  XOR U863 ( .A(n1062), .B(n1063), .Z(n1057) );
  AND U864 ( .A(n508), .B(n1064), .Z(n1063) );
  XOR U865 ( .A(p_input[696]), .B(n1062), .Z(n1064) );
  XOR U866 ( .A(n1065), .B(n1066), .Z(n1062) );
  AND U867 ( .A(n512), .B(n1067), .Z(n1066) );
  XOR U868 ( .A(n1068), .B(n1069), .Z(n1060) );
  AND U869 ( .A(n516), .B(n1067), .Z(n1069) );
  XNOR U870 ( .A(n1068), .B(n1065), .Z(n1067) );
  XOR U871 ( .A(n1070), .B(n1071), .Z(n1065) );
  AND U872 ( .A(n519), .B(n1072), .Z(n1071) );
  XOR U873 ( .A(p_input[712]), .B(n1070), .Z(n1072) );
  XOR U874 ( .A(n1073), .B(n1074), .Z(n1070) );
  AND U875 ( .A(n523), .B(n1075), .Z(n1074) );
  XOR U876 ( .A(n1076), .B(n1077), .Z(n1068) );
  AND U877 ( .A(n527), .B(n1075), .Z(n1077) );
  XNOR U878 ( .A(n1076), .B(n1073), .Z(n1075) );
  XOR U879 ( .A(n1078), .B(n1079), .Z(n1073) );
  AND U880 ( .A(n530), .B(n1080), .Z(n1079) );
  XOR U881 ( .A(p_input[728]), .B(n1078), .Z(n1080) );
  XOR U882 ( .A(n1081), .B(n1082), .Z(n1078) );
  AND U883 ( .A(n534), .B(n1083), .Z(n1082) );
  XOR U884 ( .A(n1084), .B(n1085), .Z(n1076) );
  AND U885 ( .A(n538), .B(n1083), .Z(n1085) );
  XNOR U886 ( .A(n1084), .B(n1081), .Z(n1083) );
  XOR U887 ( .A(n1086), .B(n1087), .Z(n1081) );
  AND U888 ( .A(n541), .B(n1088), .Z(n1087) );
  XOR U889 ( .A(p_input[744]), .B(n1086), .Z(n1088) );
  XOR U890 ( .A(n1089), .B(n1090), .Z(n1086) );
  AND U891 ( .A(n545), .B(n1091), .Z(n1090) );
  XOR U892 ( .A(n1092), .B(n1093), .Z(n1084) );
  AND U893 ( .A(n549), .B(n1091), .Z(n1093) );
  XNOR U894 ( .A(n1092), .B(n1089), .Z(n1091) );
  XOR U895 ( .A(n1094), .B(n1095), .Z(n1089) );
  AND U896 ( .A(n552), .B(n1096), .Z(n1095) );
  XOR U897 ( .A(p_input[760]), .B(n1094), .Z(n1096) );
  XOR U898 ( .A(n1097), .B(n1098), .Z(n1094) );
  AND U899 ( .A(n556), .B(n1099), .Z(n1098) );
  XOR U900 ( .A(n1100), .B(n1101), .Z(n1092) );
  AND U901 ( .A(n560), .B(n1099), .Z(n1101) );
  XNOR U902 ( .A(n1100), .B(n1097), .Z(n1099) );
  XOR U903 ( .A(n1102), .B(n1103), .Z(n1097) );
  AND U904 ( .A(n563), .B(n1104), .Z(n1103) );
  XOR U905 ( .A(p_input[776]), .B(n1102), .Z(n1104) );
  XOR U906 ( .A(n1105), .B(n1106), .Z(n1102) );
  AND U907 ( .A(n567), .B(n1107), .Z(n1106) );
  XOR U908 ( .A(n1108), .B(n1109), .Z(n1100) );
  AND U909 ( .A(n571), .B(n1107), .Z(n1109) );
  XNOR U910 ( .A(n1108), .B(n1105), .Z(n1107) );
  XOR U911 ( .A(n1110), .B(n1111), .Z(n1105) );
  AND U912 ( .A(n574), .B(n1112), .Z(n1111) );
  XOR U913 ( .A(p_input[792]), .B(n1110), .Z(n1112) );
  XOR U914 ( .A(n1113), .B(n1114), .Z(n1110) );
  AND U915 ( .A(n578), .B(n1115), .Z(n1114) );
  XOR U916 ( .A(n1116), .B(n1117), .Z(n1108) );
  AND U917 ( .A(n582), .B(n1115), .Z(n1117) );
  XNOR U918 ( .A(n1116), .B(n1113), .Z(n1115) );
  XOR U919 ( .A(n1118), .B(n1119), .Z(n1113) );
  AND U920 ( .A(n585), .B(n1120), .Z(n1119) );
  XOR U921 ( .A(p_input[808]), .B(n1118), .Z(n1120) );
  XOR U922 ( .A(n1121), .B(n1122), .Z(n1118) );
  AND U923 ( .A(n589), .B(n1123), .Z(n1122) );
  XOR U924 ( .A(n1124), .B(n1125), .Z(n1116) );
  AND U925 ( .A(n593), .B(n1123), .Z(n1125) );
  XNOR U926 ( .A(n1124), .B(n1121), .Z(n1123) );
  XOR U927 ( .A(n1126), .B(n1127), .Z(n1121) );
  AND U928 ( .A(n596), .B(n1128), .Z(n1127) );
  XOR U929 ( .A(p_input[824]), .B(n1126), .Z(n1128) );
  XOR U930 ( .A(n1129), .B(n1130), .Z(n1126) );
  AND U931 ( .A(n600), .B(n1131), .Z(n1130) );
  XOR U932 ( .A(n1132), .B(n1133), .Z(n1124) );
  AND U933 ( .A(n604), .B(n1131), .Z(n1133) );
  XNOR U934 ( .A(n1132), .B(n1129), .Z(n1131) );
  XOR U935 ( .A(n1134), .B(n1135), .Z(n1129) );
  AND U936 ( .A(n607), .B(n1136), .Z(n1135) );
  XOR U937 ( .A(p_input[840]), .B(n1134), .Z(n1136) );
  XOR U938 ( .A(n1137), .B(n1138), .Z(n1134) );
  AND U939 ( .A(n611), .B(n1139), .Z(n1138) );
  XOR U940 ( .A(n1140), .B(n1141), .Z(n1132) );
  AND U941 ( .A(n615), .B(n1139), .Z(n1141) );
  XNOR U942 ( .A(n1140), .B(n1137), .Z(n1139) );
  XOR U943 ( .A(n1142), .B(n1143), .Z(n1137) );
  AND U944 ( .A(n618), .B(n1144), .Z(n1143) );
  XOR U945 ( .A(p_input[856]), .B(n1142), .Z(n1144) );
  XOR U946 ( .A(n1145), .B(n1146), .Z(n1142) );
  AND U947 ( .A(n622), .B(n1147), .Z(n1146) );
  XOR U948 ( .A(n1148), .B(n1149), .Z(n1140) );
  AND U949 ( .A(n626), .B(n1147), .Z(n1149) );
  XNOR U950 ( .A(n1148), .B(n1145), .Z(n1147) );
  XOR U951 ( .A(n1150), .B(n1151), .Z(n1145) );
  AND U952 ( .A(n629), .B(n1152), .Z(n1151) );
  XOR U953 ( .A(p_input[872]), .B(n1150), .Z(n1152) );
  XOR U954 ( .A(n1153), .B(n1154), .Z(n1150) );
  AND U955 ( .A(n633), .B(n1155), .Z(n1154) );
  XOR U956 ( .A(n1156), .B(n1157), .Z(n1148) );
  AND U957 ( .A(n637), .B(n1155), .Z(n1157) );
  XNOR U958 ( .A(n1156), .B(n1153), .Z(n1155) );
  XOR U959 ( .A(n1158), .B(n1159), .Z(n1153) );
  AND U960 ( .A(n640), .B(n1160), .Z(n1159) );
  XOR U961 ( .A(p_input[888]), .B(n1158), .Z(n1160) );
  XOR U962 ( .A(n1161), .B(n1162), .Z(n1158) );
  AND U963 ( .A(n644), .B(n1163), .Z(n1162) );
  XOR U964 ( .A(n1164), .B(n1165), .Z(n1156) );
  AND U965 ( .A(n648), .B(n1163), .Z(n1165) );
  XNOR U966 ( .A(n1164), .B(n1161), .Z(n1163) );
  XOR U967 ( .A(n1166), .B(n1167), .Z(n1161) );
  AND U968 ( .A(n651), .B(n1168), .Z(n1167) );
  XOR U969 ( .A(p_input[904]), .B(n1166), .Z(n1168) );
  XOR U970 ( .A(n1169), .B(n1170), .Z(n1166) );
  AND U971 ( .A(n655), .B(n1171), .Z(n1170) );
  XOR U972 ( .A(n1172), .B(n1173), .Z(n1164) );
  AND U973 ( .A(n659), .B(n1171), .Z(n1173) );
  XNOR U974 ( .A(n1172), .B(n1169), .Z(n1171) );
  XOR U975 ( .A(n1174), .B(n1175), .Z(n1169) );
  AND U976 ( .A(n662), .B(n1176), .Z(n1175) );
  XOR U977 ( .A(p_input[920]), .B(n1174), .Z(n1176) );
  XOR U978 ( .A(n1177), .B(n1178), .Z(n1174) );
  AND U979 ( .A(n666), .B(n1179), .Z(n1178) );
  XOR U980 ( .A(n1180), .B(n1181), .Z(n1172) );
  AND U981 ( .A(n670), .B(n1179), .Z(n1181) );
  XNOR U982 ( .A(n1180), .B(n1177), .Z(n1179) );
  XOR U983 ( .A(n1182), .B(n1183), .Z(n1177) );
  AND U984 ( .A(n673), .B(n1184), .Z(n1183) );
  XOR U985 ( .A(p_input[936]), .B(n1182), .Z(n1184) );
  XOR U986 ( .A(n1185), .B(n1186), .Z(n1182) );
  AND U987 ( .A(n677), .B(n1187), .Z(n1186) );
  XOR U988 ( .A(n1188), .B(n1189), .Z(n1180) );
  AND U989 ( .A(n681), .B(n1187), .Z(n1189) );
  XNOR U990 ( .A(n1188), .B(n1185), .Z(n1187) );
  XOR U991 ( .A(n1190), .B(n1191), .Z(n1185) );
  AND U992 ( .A(n684), .B(n1192), .Z(n1191) );
  XOR U993 ( .A(p_input[952]), .B(n1190), .Z(n1192) );
  XOR U994 ( .A(n1193), .B(n1194), .Z(n1190) );
  AND U995 ( .A(n688), .B(n1195), .Z(n1194) );
  XOR U996 ( .A(n1196), .B(n1197), .Z(n1188) );
  AND U997 ( .A(n692), .B(n1195), .Z(n1197) );
  XNOR U998 ( .A(n1196), .B(n1193), .Z(n1195) );
  XOR U999 ( .A(n1198), .B(n1199), .Z(n1193) );
  AND U1000 ( .A(n695), .B(n1200), .Z(n1199) );
  XOR U1001 ( .A(p_input[968]), .B(n1198), .Z(n1200) );
  XOR U1002 ( .A(n1201), .B(n1202), .Z(n1198) );
  AND U1003 ( .A(n699), .B(n1203), .Z(n1202) );
  XOR U1004 ( .A(n1204), .B(n1205), .Z(n1196) );
  AND U1005 ( .A(n703), .B(n1203), .Z(n1205) );
  XNOR U1006 ( .A(n1204), .B(n1201), .Z(n1203) );
  XOR U1007 ( .A(n1206), .B(n1207), .Z(n1201) );
  AND U1008 ( .A(n706), .B(n1208), .Z(n1207) );
  XOR U1009 ( .A(p_input[984]), .B(n1206), .Z(n1208) );
  XNOR U1010 ( .A(n1209), .B(n1210), .Z(n1206) );
  AND U1011 ( .A(n710), .B(n1211), .Z(n1210) );
  XNOR U1012 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n1212), .Z(n1204) );
  AND U1013 ( .A(n713), .B(n1211), .Z(n1212) );
  XOR U1014 ( .A(n1213), .B(n1209), .Z(n1211) );
  XOR U1015 ( .A(n5), .B(n1214), .Z(o[23]) );
  AND U1016 ( .A(n30), .B(n1215), .Z(n5) );
  XOR U1017 ( .A(n6), .B(n1214), .Z(n1215) );
  XOR U1018 ( .A(n1216), .B(n1217), .Z(n1214) );
  AND U1019 ( .A(n34), .B(n1218), .Z(n1217) );
  XOR U1020 ( .A(p_input[7]), .B(n1216), .Z(n1218) );
  XOR U1021 ( .A(n1219), .B(n1220), .Z(n1216) );
  AND U1022 ( .A(n38), .B(n1221), .Z(n1220) );
  XOR U1023 ( .A(n1222), .B(n1223), .Z(n6) );
  AND U1024 ( .A(n42), .B(n1221), .Z(n1223) );
  XNOR U1025 ( .A(n1224), .B(n1219), .Z(n1221) );
  XOR U1026 ( .A(n1225), .B(n1226), .Z(n1219) );
  AND U1027 ( .A(n46), .B(n1227), .Z(n1226) );
  XOR U1028 ( .A(p_input[23]), .B(n1225), .Z(n1227) );
  XOR U1029 ( .A(n1228), .B(n1229), .Z(n1225) );
  AND U1030 ( .A(n50), .B(n1230), .Z(n1229) );
  IV U1031 ( .A(n1222), .Z(n1224) );
  XNOR U1032 ( .A(n1231), .B(n1232), .Z(n1222) );
  AND U1033 ( .A(n54), .B(n1230), .Z(n1232) );
  XNOR U1034 ( .A(n1231), .B(n1228), .Z(n1230) );
  XOR U1035 ( .A(n1233), .B(n1234), .Z(n1228) );
  AND U1036 ( .A(n57), .B(n1235), .Z(n1234) );
  XOR U1037 ( .A(p_input[39]), .B(n1233), .Z(n1235) );
  XOR U1038 ( .A(n1236), .B(n1237), .Z(n1233) );
  AND U1039 ( .A(n61), .B(n1238), .Z(n1237) );
  XOR U1040 ( .A(n1239), .B(n1240), .Z(n1231) );
  AND U1041 ( .A(n65), .B(n1238), .Z(n1240) );
  XNOR U1042 ( .A(n1239), .B(n1236), .Z(n1238) );
  XOR U1043 ( .A(n1241), .B(n1242), .Z(n1236) );
  AND U1044 ( .A(n68), .B(n1243), .Z(n1242) );
  XOR U1045 ( .A(p_input[55]), .B(n1241), .Z(n1243) );
  XOR U1046 ( .A(n1244), .B(n1245), .Z(n1241) );
  AND U1047 ( .A(n72), .B(n1246), .Z(n1245) );
  XOR U1048 ( .A(n1247), .B(n1248), .Z(n1239) );
  AND U1049 ( .A(n76), .B(n1246), .Z(n1248) );
  XNOR U1050 ( .A(n1247), .B(n1244), .Z(n1246) );
  XOR U1051 ( .A(n1249), .B(n1250), .Z(n1244) );
  AND U1052 ( .A(n79), .B(n1251), .Z(n1250) );
  XOR U1053 ( .A(p_input[71]), .B(n1249), .Z(n1251) );
  XOR U1054 ( .A(n1252), .B(n1253), .Z(n1249) );
  AND U1055 ( .A(n83), .B(n1254), .Z(n1253) );
  XOR U1056 ( .A(n1255), .B(n1256), .Z(n1247) );
  AND U1057 ( .A(n87), .B(n1254), .Z(n1256) );
  XNOR U1058 ( .A(n1255), .B(n1252), .Z(n1254) );
  XOR U1059 ( .A(n1257), .B(n1258), .Z(n1252) );
  AND U1060 ( .A(n90), .B(n1259), .Z(n1258) );
  XOR U1061 ( .A(p_input[87]), .B(n1257), .Z(n1259) );
  XOR U1062 ( .A(n1260), .B(n1261), .Z(n1257) );
  AND U1063 ( .A(n94), .B(n1262), .Z(n1261) );
  XOR U1064 ( .A(n1263), .B(n1264), .Z(n1255) );
  AND U1065 ( .A(n98), .B(n1262), .Z(n1264) );
  XNOR U1066 ( .A(n1263), .B(n1260), .Z(n1262) );
  XOR U1067 ( .A(n1265), .B(n1266), .Z(n1260) );
  AND U1068 ( .A(n101), .B(n1267), .Z(n1266) );
  XOR U1069 ( .A(p_input[103]), .B(n1265), .Z(n1267) );
  XOR U1070 ( .A(n1268), .B(n1269), .Z(n1265) );
  AND U1071 ( .A(n105), .B(n1270), .Z(n1269) );
  XOR U1072 ( .A(n1271), .B(n1272), .Z(n1263) );
  AND U1073 ( .A(n109), .B(n1270), .Z(n1272) );
  XNOR U1074 ( .A(n1271), .B(n1268), .Z(n1270) );
  XOR U1075 ( .A(n1273), .B(n1274), .Z(n1268) );
  AND U1076 ( .A(n112), .B(n1275), .Z(n1274) );
  XOR U1077 ( .A(p_input[119]), .B(n1273), .Z(n1275) );
  XOR U1078 ( .A(n1276), .B(n1277), .Z(n1273) );
  AND U1079 ( .A(n116), .B(n1278), .Z(n1277) );
  XOR U1080 ( .A(n1279), .B(n1280), .Z(n1271) );
  AND U1081 ( .A(n120), .B(n1278), .Z(n1280) );
  XNOR U1082 ( .A(n1279), .B(n1276), .Z(n1278) );
  XOR U1083 ( .A(n1281), .B(n1282), .Z(n1276) );
  AND U1084 ( .A(n123), .B(n1283), .Z(n1282) );
  XOR U1085 ( .A(p_input[135]), .B(n1281), .Z(n1283) );
  XOR U1086 ( .A(n1284), .B(n1285), .Z(n1281) );
  AND U1087 ( .A(n127), .B(n1286), .Z(n1285) );
  XOR U1088 ( .A(n1287), .B(n1288), .Z(n1279) );
  AND U1089 ( .A(n131), .B(n1286), .Z(n1288) );
  XNOR U1090 ( .A(n1287), .B(n1284), .Z(n1286) );
  XOR U1091 ( .A(n1289), .B(n1290), .Z(n1284) );
  AND U1092 ( .A(n134), .B(n1291), .Z(n1290) );
  XOR U1093 ( .A(p_input[151]), .B(n1289), .Z(n1291) );
  XOR U1094 ( .A(n1292), .B(n1293), .Z(n1289) );
  AND U1095 ( .A(n138), .B(n1294), .Z(n1293) );
  XOR U1096 ( .A(n1295), .B(n1296), .Z(n1287) );
  AND U1097 ( .A(n142), .B(n1294), .Z(n1296) );
  XNOR U1098 ( .A(n1295), .B(n1292), .Z(n1294) );
  XOR U1099 ( .A(n1297), .B(n1298), .Z(n1292) );
  AND U1100 ( .A(n145), .B(n1299), .Z(n1298) );
  XOR U1101 ( .A(p_input[167]), .B(n1297), .Z(n1299) );
  XOR U1102 ( .A(n1300), .B(n1301), .Z(n1297) );
  AND U1103 ( .A(n149), .B(n1302), .Z(n1301) );
  XOR U1104 ( .A(n1303), .B(n1304), .Z(n1295) );
  AND U1105 ( .A(n153), .B(n1302), .Z(n1304) );
  XNOR U1106 ( .A(n1303), .B(n1300), .Z(n1302) );
  XOR U1107 ( .A(n1305), .B(n1306), .Z(n1300) );
  AND U1108 ( .A(n156), .B(n1307), .Z(n1306) );
  XOR U1109 ( .A(p_input[183]), .B(n1305), .Z(n1307) );
  XOR U1110 ( .A(n1308), .B(n1309), .Z(n1305) );
  AND U1111 ( .A(n160), .B(n1310), .Z(n1309) );
  XOR U1112 ( .A(n1311), .B(n1312), .Z(n1303) );
  AND U1113 ( .A(n164), .B(n1310), .Z(n1312) );
  XNOR U1114 ( .A(n1311), .B(n1308), .Z(n1310) );
  XOR U1115 ( .A(n1313), .B(n1314), .Z(n1308) );
  AND U1116 ( .A(n167), .B(n1315), .Z(n1314) );
  XOR U1117 ( .A(p_input[199]), .B(n1313), .Z(n1315) );
  XOR U1118 ( .A(n1316), .B(n1317), .Z(n1313) );
  AND U1119 ( .A(n171), .B(n1318), .Z(n1317) );
  XOR U1120 ( .A(n1319), .B(n1320), .Z(n1311) );
  AND U1121 ( .A(n175), .B(n1318), .Z(n1320) );
  XNOR U1122 ( .A(n1319), .B(n1316), .Z(n1318) );
  XOR U1123 ( .A(n1321), .B(n1322), .Z(n1316) );
  AND U1124 ( .A(n178), .B(n1323), .Z(n1322) );
  XOR U1125 ( .A(p_input[215]), .B(n1321), .Z(n1323) );
  XOR U1126 ( .A(n1324), .B(n1325), .Z(n1321) );
  AND U1127 ( .A(n182), .B(n1326), .Z(n1325) );
  XOR U1128 ( .A(n1327), .B(n1328), .Z(n1319) );
  AND U1129 ( .A(n186), .B(n1326), .Z(n1328) );
  XNOR U1130 ( .A(n1327), .B(n1324), .Z(n1326) );
  XOR U1131 ( .A(n1329), .B(n1330), .Z(n1324) );
  AND U1132 ( .A(n189), .B(n1331), .Z(n1330) );
  XOR U1133 ( .A(p_input[231]), .B(n1329), .Z(n1331) );
  XOR U1134 ( .A(n1332), .B(n1333), .Z(n1329) );
  AND U1135 ( .A(n193), .B(n1334), .Z(n1333) );
  XOR U1136 ( .A(n1335), .B(n1336), .Z(n1327) );
  AND U1137 ( .A(n197), .B(n1334), .Z(n1336) );
  XNOR U1138 ( .A(n1335), .B(n1332), .Z(n1334) );
  XOR U1139 ( .A(n1337), .B(n1338), .Z(n1332) );
  AND U1140 ( .A(n200), .B(n1339), .Z(n1338) );
  XOR U1141 ( .A(p_input[247]), .B(n1337), .Z(n1339) );
  XOR U1142 ( .A(n1340), .B(n1341), .Z(n1337) );
  AND U1143 ( .A(n204), .B(n1342), .Z(n1341) );
  XOR U1144 ( .A(n1343), .B(n1344), .Z(n1335) );
  AND U1145 ( .A(n208), .B(n1342), .Z(n1344) );
  XNOR U1146 ( .A(n1343), .B(n1340), .Z(n1342) );
  XOR U1147 ( .A(n1345), .B(n1346), .Z(n1340) );
  AND U1148 ( .A(n211), .B(n1347), .Z(n1346) );
  XOR U1149 ( .A(p_input[263]), .B(n1345), .Z(n1347) );
  XOR U1150 ( .A(n1348), .B(n1349), .Z(n1345) );
  AND U1151 ( .A(n215), .B(n1350), .Z(n1349) );
  XOR U1152 ( .A(n1351), .B(n1352), .Z(n1343) );
  AND U1153 ( .A(n219), .B(n1350), .Z(n1352) );
  XNOR U1154 ( .A(n1351), .B(n1348), .Z(n1350) );
  XOR U1155 ( .A(n1353), .B(n1354), .Z(n1348) );
  AND U1156 ( .A(n222), .B(n1355), .Z(n1354) );
  XOR U1157 ( .A(p_input[279]), .B(n1353), .Z(n1355) );
  XOR U1158 ( .A(n1356), .B(n1357), .Z(n1353) );
  AND U1159 ( .A(n226), .B(n1358), .Z(n1357) );
  XOR U1160 ( .A(n1359), .B(n1360), .Z(n1351) );
  AND U1161 ( .A(n230), .B(n1358), .Z(n1360) );
  XNOR U1162 ( .A(n1359), .B(n1356), .Z(n1358) );
  XOR U1163 ( .A(n1361), .B(n1362), .Z(n1356) );
  AND U1164 ( .A(n233), .B(n1363), .Z(n1362) );
  XOR U1165 ( .A(p_input[295]), .B(n1361), .Z(n1363) );
  XOR U1166 ( .A(n1364), .B(n1365), .Z(n1361) );
  AND U1167 ( .A(n237), .B(n1366), .Z(n1365) );
  XOR U1168 ( .A(n1367), .B(n1368), .Z(n1359) );
  AND U1169 ( .A(n241), .B(n1366), .Z(n1368) );
  XNOR U1170 ( .A(n1367), .B(n1364), .Z(n1366) );
  XOR U1171 ( .A(n1369), .B(n1370), .Z(n1364) );
  AND U1172 ( .A(n244), .B(n1371), .Z(n1370) );
  XOR U1173 ( .A(p_input[311]), .B(n1369), .Z(n1371) );
  XOR U1174 ( .A(n1372), .B(n1373), .Z(n1369) );
  AND U1175 ( .A(n248), .B(n1374), .Z(n1373) );
  XOR U1176 ( .A(n1375), .B(n1376), .Z(n1367) );
  AND U1177 ( .A(n252), .B(n1374), .Z(n1376) );
  XNOR U1178 ( .A(n1375), .B(n1372), .Z(n1374) );
  XOR U1179 ( .A(n1377), .B(n1378), .Z(n1372) );
  AND U1180 ( .A(n255), .B(n1379), .Z(n1378) );
  XOR U1181 ( .A(p_input[327]), .B(n1377), .Z(n1379) );
  XOR U1182 ( .A(n1380), .B(n1381), .Z(n1377) );
  AND U1183 ( .A(n259), .B(n1382), .Z(n1381) );
  XOR U1184 ( .A(n1383), .B(n1384), .Z(n1375) );
  AND U1185 ( .A(n263), .B(n1382), .Z(n1384) );
  XNOR U1186 ( .A(n1383), .B(n1380), .Z(n1382) );
  XOR U1187 ( .A(n1385), .B(n1386), .Z(n1380) );
  AND U1188 ( .A(n266), .B(n1387), .Z(n1386) );
  XOR U1189 ( .A(p_input[343]), .B(n1385), .Z(n1387) );
  XOR U1190 ( .A(n1388), .B(n1389), .Z(n1385) );
  AND U1191 ( .A(n270), .B(n1390), .Z(n1389) );
  XOR U1192 ( .A(n1391), .B(n1392), .Z(n1383) );
  AND U1193 ( .A(n274), .B(n1390), .Z(n1392) );
  XNOR U1194 ( .A(n1391), .B(n1388), .Z(n1390) );
  XOR U1195 ( .A(n1393), .B(n1394), .Z(n1388) );
  AND U1196 ( .A(n277), .B(n1395), .Z(n1394) );
  XOR U1197 ( .A(p_input[359]), .B(n1393), .Z(n1395) );
  XOR U1198 ( .A(n1396), .B(n1397), .Z(n1393) );
  AND U1199 ( .A(n281), .B(n1398), .Z(n1397) );
  XOR U1200 ( .A(n1399), .B(n1400), .Z(n1391) );
  AND U1201 ( .A(n285), .B(n1398), .Z(n1400) );
  XNOR U1202 ( .A(n1399), .B(n1396), .Z(n1398) );
  XOR U1203 ( .A(n1401), .B(n1402), .Z(n1396) );
  AND U1204 ( .A(n288), .B(n1403), .Z(n1402) );
  XOR U1205 ( .A(p_input[375]), .B(n1401), .Z(n1403) );
  XOR U1206 ( .A(n1404), .B(n1405), .Z(n1401) );
  AND U1207 ( .A(n292), .B(n1406), .Z(n1405) );
  XOR U1208 ( .A(n1407), .B(n1408), .Z(n1399) );
  AND U1209 ( .A(n296), .B(n1406), .Z(n1408) );
  XNOR U1210 ( .A(n1407), .B(n1404), .Z(n1406) );
  XOR U1211 ( .A(n1409), .B(n1410), .Z(n1404) );
  AND U1212 ( .A(n299), .B(n1411), .Z(n1410) );
  XOR U1213 ( .A(p_input[391]), .B(n1409), .Z(n1411) );
  XOR U1214 ( .A(n1412), .B(n1413), .Z(n1409) );
  AND U1215 ( .A(n303), .B(n1414), .Z(n1413) );
  XOR U1216 ( .A(n1415), .B(n1416), .Z(n1407) );
  AND U1217 ( .A(n307), .B(n1414), .Z(n1416) );
  XNOR U1218 ( .A(n1415), .B(n1412), .Z(n1414) );
  XOR U1219 ( .A(n1417), .B(n1418), .Z(n1412) );
  AND U1220 ( .A(n310), .B(n1419), .Z(n1418) );
  XOR U1221 ( .A(p_input[407]), .B(n1417), .Z(n1419) );
  XOR U1222 ( .A(n1420), .B(n1421), .Z(n1417) );
  AND U1223 ( .A(n314), .B(n1422), .Z(n1421) );
  XOR U1224 ( .A(n1423), .B(n1424), .Z(n1415) );
  AND U1225 ( .A(n318), .B(n1422), .Z(n1424) );
  XNOR U1226 ( .A(n1423), .B(n1420), .Z(n1422) );
  XOR U1227 ( .A(n1425), .B(n1426), .Z(n1420) );
  AND U1228 ( .A(n321), .B(n1427), .Z(n1426) );
  XOR U1229 ( .A(p_input[423]), .B(n1425), .Z(n1427) );
  XOR U1230 ( .A(n1428), .B(n1429), .Z(n1425) );
  AND U1231 ( .A(n325), .B(n1430), .Z(n1429) );
  XOR U1232 ( .A(n1431), .B(n1432), .Z(n1423) );
  AND U1233 ( .A(n329), .B(n1430), .Z(n1432) );
  XNOR U1234 ( .A(n1431), .B(n1428), .Z(n1430) );
  XOR U1235 ( .A(n1433), .B(n1434), .Z(n1428) );
  AND U1236 ( .A(n332), .B(n1435), .Z(n1434) );
  XOR U1237 ( .A(p_input[439]), .B(n1433), .Z(n1435) );
  XOR U1238 ( .A(n1436), .B(n1437), .Z(n1433) );
  AND U1239 ( .A(n336), .B(n1438), .Z(n1437) );
  XOR U1240 ( .A(n1439), .B(n1440), .Z(n1431) );
  AND U1241 ( .A(n340), .B(n1438), .Z(n1440) );
  XNOR U1242 ( .A(n1439), .B(n1436), .Z(n1438) );
  XOR U1243 ( .A(n1441), .B(n1442), .Z(n1436) );
  AND U1244 ( .A(n343), .B(n1443), .Z(n1442) );
  XOR U1245 ( .A(p_input[455]), .B(n1441), .Z(n1443) );
  XOR U1246 ( .A(n1444), .B(n1445), .Z(n1441) );
  AND U1247 ( .A(n347), .B(n1446), .Z(n1445) );
  XOR U1248 ( .A(n1447), .B(n1448), .Z(n1439) );
  AND U1249 ( .A(n351), .B(n1446), .Z(n1448) );
  XNOR U1250 ( .A(n1447), .B(n1444), .Z(n1446) );
  XOR U1251 ( .A(n1449), .B(n1450), .Z(n1444) );
  AND U1252 ( .A(n354), .B(n1451), .Z(n1450) );
  XOR U1253 ( .A(p_input[471]), .B(n1449), .Z(n1451) );
  XOR U1254 ( .A(n1452), .B(n1453), .Z(n1449) );
  AND U1255 ( .A(n358), .B(n1454), .Z(n1453) );
  XOR U1256 ( .A(n1455), .B(n1456), .Z(n1447) );
  AND U1257 ( .A(n362), .B(n1454), .Z(n1456) );
  XNOR U1258 ( .A(n1455), .B(n1452), .Z(n1454) );
  XOR U1259 ( .A(n1457), .B(n1458), .Z(n1452) );
  AND U1260 ( .A(n365), .B(n1459), .Z(n1458) );
  XOR U1261 ( .A(p_input[487]), .B(n1457), .Z(n1459) );
  XOR U1262 ( .A(n1460), .B(n1461), .Z(n1457) );
  AND U1263 ( .A(n369), .B(n1462), .Z(n1461) );
  XOR U1264 ( .A(n1463), .B(n1464), .Z(n1455) );
  AND U1265 ( .A(n373), .B(n1462), .Z(n1464) );
  XNOR U1266 ( .A(n1463), .B(n1460), .Z(n1462) );
  XOR U1267 ( .A(n1465), .B(n1466), .Z(n1460) );
  AND U1268 ( .A(n376), .B(n1467), .Z(n1466) );
  XOR U1269 ( .A(p_input[503]), .B(n1465), .Z(n1467) );
  XOR U1270 ( .A(n1468), .B(n1469), .Z(n1465) );
  AND U1271 ( .A(n380), .B(n1470), .Z(n1469) );
  XOR U1272 ( .A(n1471), .B(n1472), .Z(n1463) );
  AND U1273 ( .A(n384), .B(n1470), .Z(n1472) );
  XNOR U1274 ( .A(n1471), .B(n1468), .Z(n1470) );
  XOR U1275 ( .A(n1473), .B(n1474), .Z(n1468) );
  AND U1276 ( .A(n387), .B(n1475), .Z(n1474) );
  XOR U1277 ( .A(p_input[519]), .B(n1473), .Z(n1475) );
  XOR U1278 ( .A(n1476), .B(n1477), .Z(n1473) );
  AND U1279 ( .A(n391), .B(n1478), .Z(n1477) );
  XOR U1280 ( .A(n1479), .B(n1480), .Z(n1471) );
  AND U1281 ( .A(n395), .B(n1478), .Z(n1480) );
  XNOR U1282 ( .A(n1479), .B(n1476), .Z(n1478) );
  XOR U1283 ( .A(n1481), .B(n1482), .Z(n1476) );
  AND U1284 ( .A(n398), .B(n1483), .Z(n1482) );
  XOR U1285 ( .A(p_input[535]), .B(n1481), .Z(n1483) );
  XOR U1286 ( .A(n1484), .B(n1485), .Z(n1481) );
  AND U1287 ( .A(n402), .B(n1486), .Z(n1485) );
  XOR U1288 ( .A(n1487), .B(n1488), .Z(n1479) );
  AND U1289 ( .A(n406), .B(n1486), .Z(n1488) );
  XNOR U1290 ( .A(n1487), .B(n1484), .Z(n1486) );
  XOR U1291 ( .A(n1489), .B(n1490), .Z(n1484) );
  AND U1292 ( .A(n409), .B(n1491), .Z(n1490) );
  XOR U1293 ( .A(p_input[551]), .B(n1489), .Z(n1491) );
  XOR U1294 ( .A(n1492), .B(n1493), .Z(n1489) );
  AND U1295 ( .A(n413), .B(n1494), .Z(n1493) );
  XOR U1296 ( .A(n1495), .B(n1496), .Z(n1487) );
  AND U1297 ( .A(n417), .B(n1494), .Z(n1496) );
  XNOR U1298 ( .A(n1495), .B(n1492), .Z(n1494) );
  XOR U1299 ( .A(n1497), .B(n1498), .Z(n1492) );
  AND U1300 ( .A(n420), .B(n1499), .Z(n1498) );
  XOR U1301 ( .A(p_input[567]), .B(n1497), .Z(n1499) );
  XOR U1302 ( .A(n1500), .B(n1501), .Z(n1497) );
  AND U1303 ( .A(n424), .B(n1502), .Z(n1501) );
  XOR U1304 ( .A(n1503), .B(n1504), .Z(n1495) );
  AND U1305 ( .A(n428), .B(n1502), .Z(n1504) );
  XNOR U1306 ( .A(n1503), .B(n1500), .Z(n1502) );
  XOR U1307 ( .A(n1505), .B(n1506), .Z(n1500) );
  AND U1308 ( .A(n431), .B(n1507), .Z(n1506) );
  XOR U1309 ( .A(p_input[583]), .B(n1505), .Z(n1507) );
  XOR U1310 ( .A(n1508), .B(n1509), .Z(n1505) );
  AND U1311 ( .A(n435), .B(n1510), .Z(n1509) );
  XOR U1312 ( .A(n1511), .B(n1512), .Z(n1503) );
  AND U1313 ( .A(n439), .B(n1510), .Z(n1512) );
  XNOR U1314 ( .A(n1511), .B(n1508), .Z(n1510) );
  XOR U1315 ( .A(n1513), .B(n1514), .Z(n1508) );
  AND U1316 ( .A(n442), .B(n1515), .Z(n1514) );
  XOR U1317 ( .A(p_input[599]), .B(n1513), .Z(n1515) );
  XOR U1318 ( .A(n1516), .B(n1517), .Z(n1513) );
  AND U1319 ( .A(n446), .B(n1518), .Z(n1517) );
  XOR U1320 ( .A(n1519), .B(n1520), .Z(n1511) );
  AND U1321 ( .A(n450), .B(n1518), .Z(n1520) );
  XNOR U1322 ( .A(n1519), .B(n1516), .Z(n1518) );
  XOR U1323 ( .A(n1521), .B(n1522), .Z(n1516) );
  AND U1324 ( .A(n453), .B(n1523), .Z(n1522) );
  XOR U1325 ( .A(p_input[615]), .B(n1521), .Z(n1523) );
  XOR U1326 ( .A(n1524), .B(n1525), .Z(n1521) );
  AND U1327 ( .A(n457), .B(n1526), .Z(n1525) );
  XOR U1328 ( .A(n1527), .B(n1528), .Z(n1519) );
  AND U1329 ( .A(n461), .B(n1526), .Z(n1528) );
  XNOR U1330 ( .A(n1527), .B(n1524), .Z(n1526) );
  XOR U1331 ( .A(n1529), .B(n1530), .Z(n1524) );
  AND U1332 ( .A(n464), .B(n1531), .Z(n1530) );
  XOR U1333 ( .A(p_input[631]), .B(n1529), .Z(n1531) );
  XOR U1334 ( .A(n1532), .B(n1533), .Z(n1529) );
  AND U1335 ( .A(n468), .B(n1534), .Z(n1533) );
  XOR U1336 ( .A(n1535), .B(n1536), .Z(n1527) );
  AND U1337 ( .A(n472), .B(n1534), .Z(n1536) );
  XNOR U1338 ( .A(n1535), .B(n1532), .Z(n1534) );
  XOR U1339 ( .A(n1537), .B(n1538), .Z(n1532) );
  AND U1340 ( .A(n475), .B(n1539), .Z(n1538) );
  XOR U1341 ( .A(p_input[647]), .B(n1537), .Z(n1539) );
  XOR U1342 ( .A(n1540), .B(n1541), .Z(n1537) );
  AND U1343 ( .A(n479), .B(n1542), .Z(n1541) );
  XOR U1344 ( .A(n1543), .B(n1544), .Z(n1535) );
  AND U1345 ( .A(n483), .B(n1542), .Z(n1544) );
  XNOR U1346 ( .A(n1543), .B(n1540), .Z(n1542) );
  XOR U1347 ( .A(n1545), .B(n1546), .Z(n1540) );
  AND U1348 ( .A(n486), .B(n1547), .Z(n1546) );
  XOR U1349 ( .A(p_input[663]), .B(n1545), .Z(n1547) );
  XOR U1350 ( .A(n1548), .B(n1549), .Z(n1545) );
  AND U1351 ( .A(n490), .B(n1550), .Z(n1549) );
  XOR U1352 ( .A(n1551), .B(n1552), .Z(n1543) );
  AND U1353 ( .A(n494), .B(n1550), .Z(n1552) );
  XNOR U1354 ( .A(n1551), .B(n1548), .Z(n1550) );
  XOR U1355 ( .A(n1553), .B(n1554), .Z(n1548) );
  AND U1356 ( .A(n497), .B(n1555), .Z(n1554) );
  XOR U1357 ( .A(p_input[679]), .B(n1553), .Z(n1555) );
  XOR U1358 ( .A(n1556), .B(n1557), .Z(n1553) );
  AND U1359 ( .A(n501), .B(n1558), .Z(n1557) );
  XOR U1360 ( .A(n1559), .B(n1560), .Z(n1551) );
  AND U1361 ( .A(n505), .B(n1558), .Z(n1560) );
  XNOR U1362 ( .A(n1559), .B(n1556), .Z(n1558) );
  XOR U1363 ( .A(n1561), .B(n1562), .Z(n1556) );
  AND U1364 ( .A(n508), .B(n1563), .Z(n1562) );
  XOR U1365 ( .A(p_input[695]), .B(n1561), .Z(n1563) );
  XOR U1366 ( .A(n1564), .B(n1565), .Z(n1561) );
  AND U1367 ( .A(n512), .B(n1566), .Z(n1565) );
  XOR U1368 ( .A(n1567), .B(n1568), .Z(n1559) );
  AND U1369 ( .A(n516), .B(n1566), .Z(n1568) );
  XNOR U1370 ( .A(n1567), .B(n1564), .Z(n1566) );
  XOR U1371 ( .A(n1569), .B(n1570), .Z(n1564) );
  AND U1372 ( .A(n519), .B(n1571), .Z(n1570) );
  XOR U1373 ( .A(p_input[711]), .B(n1569), .Z(n1571) );
  XOR U1374 ( .A(n1572), .B(n1573), .Z(n1569) );
  AND U1375 ( .A(n523), .B(n1574), .Z(n1573) );
  XOR U1376 ( .A(n1575), .B(n1576), .Z(n1567) );
  AND U1377 ( .A(n527), .B(n1574), .Z(n1576) );
  XNOR U1378 ( .A(n1575), .B(n1572), .Z(n1574) );
  XOR U1379 ( .A(n1577), .B(n1578), .Z(n1572) );
  AND U1380 ( .A(n530), .B(n1579), .Z(n1578) );
  XOR U1381 ( .A(p_input[727]), .B(n1577), .Z(n1579) );
  XOR U1382 ( .A(n1580), .B(n1581), .Z(n1577) );
  AND U1383 ( .A(n534), .B(n1582), .Z(n1581) );
  XOR U1384 ( .A(n1583), .B(n1584), .Z(n1575) );
  AND U1385 ( .A(n538), .B(n1582), .Z(n1584) );
  XNOR U1386 ( .A(n1583), .B(n1580), .Z(n1582) );
  XOR U1387 ( .A(n1585), .B(n1586), .Z(n1580) );
  AND U1388 ( .A(n541), .B(n1587), .Z(n1586) );
  XOR U1389 ( .A(p_input[743]), .B(n1585), .Z(n1587) );
  XOR U1390 ( .A(n1588), .B(n1589), .Z(n1585) );
  AND U1391 ( .A(n545), .B(n1590), .Z(n1589) );
  XOR U1392 ( .A(n1591), .B(n1592), .Z(n1583) );
  AND U1393 ( .A(n549), .B(n1590), .Z(n1592) );
  XNOR U1394 ( .A(n1591), .B(n1588), .Z(n1590) );
  XOR U1395 ( .A(n1593), .B(n1594), .Z(n1588) );
  AND U1396 ( .A(n552), .B(n1595), .Z(n1594) );
  XOR U1397 ( .A(p_input[759]), .B(n1593), .Z(n1595) );
  XOR U1398 ( .A(n1596), .B(n1597), .Z(n1593) );
  AND U1399 ( .A(n556), .B(n1598), .Z(n1597) );
  XOR U1400 ( .A(n1599), .B(n1600), .Z(n1591) );
  AND U1401 ( .A(n560), .B(n1598), .Z(n1600) );
  XNOR U1402 ( .A(n1599), .B(n1596), .Z(n1598) );
  XOR U1403 ( .A(n1601), .B(n1602), .Z(n1596) );
  AND U1404 ( .A(n563), .B(n1603), .Z(n1602) );
  XOR U1405 ( .A(p_input[775]), .B(n1601), .Z(n1603) );
  XOR U1406 ( .A(n1604), .B(n1605), .Z(n1601) );
  AND U1407 ( .A(n567), .B(n1606), .Z(n1605) );
  XOR U1408 ( .A(n1607), .B(n1608), .Z(n1599) );
  AND U1409 ( .A(n571), .B(n1606), .Z(n1608) );
  XNOR U1410 ( .A(n1607), .B(n1604), .Z(n1606) );
  XOR U1411 ( .A(n1609), .B(n1610), .Z(n1604) );
  AND U1412 ( .A(n574), .B(n1611), .Z(n1610) );
  XOR U1413 ( .A(p_input[791]), .B(n1609), .Z(n1611) );
  XOR U1414 ( .A(n1612), .B(n1613), .Z(n1609) );
  AND U1415 ( .A(n578), .B(n1614), .Z(n1613) );
  XOR U1416 ( .A(n1615), .B(n1616), .Z(n1607) );
  AND U1417 ( .A(n582), .B(n1614), .Z(n1616) );
  XNOR U1418 ( .A(n1615), .B(n1612), .Z(n1614) );
  XOR U1419 ( .A(n1617), .B(n1618), .Z(n1612) );
  AND U1420 ( .A(n585), .B(n1619), .Z(n1618) );
  XOR U1421 ( .A(p_input[807]), .B(n1617), .Z(n1619) );
  XOR U1422 ( .A(n1620), .B(n1621), .Z(n1617) );
  AND U1423 ( .A(n589), .B(n1622), .Z(n1621) );
  XOR U1424 ( .A(n1623), .B(n1624), .Z(n1615) );
  AND U1425 ( .A(n593), .B(n1622), .Z(n1624) );
  XNOR U1426 ( .A(n1623), .B(n1620), .Z(n1622) );
  XOR U1427 ( .A(n1625), .B(n1626), .Z(n1620) );
  AND U1428 ( .A(n596), .B(n1627), .Z(n1626) );
  XOR U1429 ( .A(p_input[823]), .B(n1625), .Z(n1627) );
  XOR U1430 ( .A(n1628), .B(n1629), .Z(n1625) );
  AND U1431 ( .A(n600), .B(n1630), .Z(n1629) );
  XOR U1432 ( .A(n1631), .B(n1632), .Z(n1623) );
  AND U1433 ( .A(n604), .B(n1630), .Z(n1632) );
  XNOR U1434 ( .A(n1631), .B(n1628), .Z(n1630) );
  XOR U1435 ( .A(n1633), .B(n1634), .Z(n1628) );
  AND U1436 ( .A(n607), .B(n1635), .Z(n1634) );
  XOR U1437 ( .A(p_input[839]), .B(n1633), .Z(n1635) );
  XOR U1438 ( .A(n1636), .B(n1637), .Z(n1633) );
  AND U1439 ( .A(n611), .B(n1638), .Z(n1637) );
  XOR U1440 ( .A(n1639), .B(n1640), .Z(n1631) );
  AND U1441 ( .A(n615), .B(n1638), .Z(n1640) );
  XNOR U1442 ( .A(n1639), .B(n1636), .Z(n1638) );
  XOR U1443 ( .A(n1641), .B(n1642), .Z(n1636) );
  AND U1444 ( .A(n618), .B(n1643), .Z(n1642) );
  XOR U1445 ( .A(p_input[855]), .B(n1641), .Z(n1643) );
  XOR U1446 ( .A(n1644), .B(n1645), .Z(n1641) );
  AND U1447 ( .A(n622), .B(n1646), .Z(n1645) );
  XOR U1448 ( .A(n1647), .B(n1648), .Z(n1639) );
  AND U1449 ( .A(n626), .B(n1646), .Z(n1648) );
  XNOR U1450 ( .A(n1647), .B(n1644), .Z(n1646) );
  XOR U1451 ( .A(n1649), .B(n1650), .Z(n1644) );
  AND U1452 ( .A(n629), .B(n1651), .Z(n1650) );
  XOR U1453 ( .A(p_input[871]), .B(n1649), .Z(n1651) );
  XOR U1454 ( .A(n1652), .B(n1653), .Z(n1649) );
  AND U1455 ( .A(n633), .B(n1654), .Z(n1653) );
  XOR U1456 ( .A(n1655), .B(n1656), .Z(n1647) );
  AND U1457 ( .A(n637), .B(n1654), .Z(n1656) );
  XNOR U1458 ( .A(n1655), .B(n1652), .Z(n1654) );
  XOR U1459 ( .A(n1657), .B(n1658), .Z(n1652) );
  AND U1460 ( .A(n640), .B(n1659), .Z(n1658) );
  XOR U1461 ( .A(p_input[887]), .B(n1657), .Z(n1659) );
  XOR U1462 ( .A(n1660), .B(n1661), .Z(n1657) );
  AND U1463 ( .A(n644), .B(n1662), .Z(n1661) );
  XOR U1464 ( .A(n1663), .B(n1664), .Z(n1655) );
  AND U1465 ( .A(n648), .B(n1662), .Z(n1664) );
  XNOR U1466 ( .A(n1663), .B(n1660), .Z(n1662) );
  XOR U1467 ( .A(n1665), .B(n1666), .Z(n1660) );
  AND U1468 ( .A(n651), .B(n1667), .Z(n1666) );
  XOR U1469 ( .A(p_input[903]), .B(n1665), .Z(n1667) );
  XOR U1470 ( .A(n1668), .B(n1669), .Z(n1665) );
  AND U1471 ( .A(n655), .B(n1670), .Z(n1669) );
  XOR U1472 ( .A(n1671), .B(n1672), .Z(n1663) );
  AND U1473 ( .A(n659), .B(n1670), .Z(n1672) );
  XNOR U1474 ( .A(n1671), .B(n1668), .Z(n1670) );
  XOR U1475 ( .A(n1673), .B(n1674), .Z(n1668) );
  AND U1476 ( .A(n662), .B(n1675), .Z(n1674) );
  XOR U1477 ( .A(p_input[919]), .B(n1673), .Z(n1675) );
  XOR U1478 ( .A(n1676), .B(n1677), .Z(n1673) );
  AND U1479 ( .A(n666), .B(n1678), .Z(n1677) );
  XOR U1480 ( .A(n1679), .B(n1680), .Z(n1671) );
  AND U1481 ( .A(n670), .B(n1678), .Z(n1680) );
  XNOR U1482 ( .A(n1679), .B(n1676), .Z(n1678) );
  XOR U1483 ( .A(n1681), .B(n1682), .Z(n1676) );
  AND U1484 ( .A(n673), .B(n1683), .Z(n1682) );
  XOR U1485 ( .A(p_input[935]), .B(n1681), .Z(n1683) );
  XOR U1486 ( .A(n1684), .B(n1685), .Z(n1681) );
  AND U1487 ( .A(n677), .B(n1686), .Z(n1685) );
  XOR U1488 ( .A(n1687), .B(n1688), .Z(n1679) );
  AND U1489 ( .A(n681), .B(n1686), .Z(n1688) );
  XNOR U1490 ( .A(n1687), .B(n1684), .Z(n1686) );
  XOR U1491 ( .A(n1689), .B(n1690), .Z(n1684) );
  AND U1492 ( .A(n684), .B(n1691), .Z(n1690) );
  XOR U1493 ( .A(p_input[951]), .B(n1689), .Z(n1691) );
  XOR U1494 ( .A(n1692), .B(n1693), .Z(n1689) );
  AND U1495 ( .A(n688), .B(n1694), .Z(n1693) );
  XOR U1496 ( .A(n1695), .B(n1696), .Z(n1687) );
  AND U1497 ( .A(n692), .B(n1694), .Z(n1696) );
  XNOR U1498 ( .A(n1695), .B(n1692), .Z(n1694) );
  XOR U1499 ( .A(n1697), .B(n1698), .Z(n1692) );
  AND U1500 ( .A(n695), .B(n1699), .Z(n1698) );
  XOR U1501 ( .A(p_input[967]), .B(n1697), .Z(n1699) );
  XOR U1502 ( .A(n1700), .B(n1701), .Z(n1697) );
  AND U1503 ( .A(n699), .B(n1702), .Z(n1701) );
  XOR U1504 ( .A(n1703), .B(n1704), .Z(n1695) );
  AND U1505 ( .A(n703), .B(n1702), .Z(n1704) );
  XNOR U1506 ( .A(n1703), .B(n1700), .Z(n1702) );
  XOR U1507 ( .A(n1705), .B(n1706), .Z(n1700) );
  AND U1508 ( .A(n706), .B(n1707), .Z(n1706) );
  XOR U1509 ( .A(p_input[983]), .B(n1705), .Z(n1707) );
  XNOR U1510 ( .A(n1708), .B(n1709), .Z(n1705) );
  AND U1511 ( .A(n710), .B(n1710), .Z(n1709) );
  XNOR U1512 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n1711), .Z(n1703) );
  AND U1513 ( .A(n713), .B(n1710), .Z(n1711) );
  XOR U1514 ( .A(n1712), .B(n1708), .Z(n1710) );
  IV U1515 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .Z(n1708) );
  IV U1516 ( .A(\knn_comb_/min_val_out[0][7] ), .Z(n1712) );
  XOR U1517 ( .A(n7), .B(n1713), .Z(o[22]) );
  AND U1518 ( .A(n30), .B(n1714), .Z(n7) );
  XOR U1519 ( .A(n8), .B(n1713), .Z(n1714) );
  XOR U1520 ( .A(n1715), .B(n1716), .Z(n1713) );
  AND U1521 ( .A(n34), .B(n1717), .Z(n1716) );
  XOR U1522 ( .A(p_input[6]), .B(n1715), .Z(n1717) );
  XOR U1523 ( .A(n1718), .B(n1719), .Z(n1715) );
  AND U1524 ( .A(n38), .B(n1720), .Z(n1719) );
  XOR U1525 ( .A(n1721), .B(n1722), .Z(n8) );
  AND U1526 ( .A(n42), .B(n1720), .Z(n1722) );
  XNOR U1527 ( .A(n1723), .B(n1718), .Z(n1720) );
  XOR U1528 ( .A(n1724), .B(n1725), .Z(n1718) );
  AND U1529 ( .A(n46), .B(n1726), .Z(n1725) );
  XOR U1530 ( .A(p_input[22]), .B(n1724), .Z(n1726) );
  XOR U1531 ( .A(n1727), .B(n1728), .Z(n1724) );
  AND U1532 ( .A(n50), .B(n1729), .Z(n1728) );
  IV U1533 ( .A(n1721), .Z(n1723) );
  XNOR U1534 ( .A(n1730), .B(n1731), .Z(n1721) );
  AND U1535 ( .A(n54), .B(n1729), .Z(n1731) );
  XNOR U1536 ( .A(n1730), .B(n1727), .Z(n1729) );
  XOR U1537 ( .A(n1732), .B(n1733), .Z(n1727) );
  AND U1538 ( .A(n57), .B(n1734), .Z(n1733) );
  XOR U1539 ( .A(p_input[38]), .B(n1732), .Z(n1734) );
  XOR U1540 ( .A(n1735), .B(n1736), .Z(n1732) );
  AND U1541 ( .A(n61), .B(n1737), .Z(n1736) );
  XOR U1542 ( .A(n1738), .B(n1739), .Z(n1730) );
  AND U1543 ( .A(n65), .B(n1737), .Z(n1739) );
  XNOR U1544 ( .A(n1738), .B(n1735), .Z(n1737) );
  XOR U1545 ( .A(n1740), .B(n1741), .Z(n1735) );
  AND U1546 ( .A(n68), .B(n1742), .Z(n1741) );
  XOR U1547 ( .A(p_input[54]), .B(n1740), .Z(n1742) );
  XOR U1548 ( .A(n1743), .B(n1744), .Z(n1740) );
  AND U1549 ( .A(n72), .B(n1745), .Z(n1744) );
  XOR U1550 ( .A(n1746), .B(n1747), .Z(n1738) );
  AND U1551 ( .A(n76), .B(n1745), .Z(n1747) );
  XNOR U1552 ( .A(n1746), .B(n1743), .Z(n1745) );
  XOR U1553 ( .A(n1748), .B(n1749), .Z(n1743) );
  AND U1554 ( .A(n79), .B(n1750), .Z(n1749) );
  XOR U1555 ( .A(p_input[70]), .B(n1748), .Z(n1750) );
  XOR U1556 ( .A(n1751), .B(n1752), .Z(n1748) );
  AND U1557 ( .A(n83), .B(n1753), .Z(n1752) );
  XOR U1558 ( .A(n1754), .B(n1755), .Z(n1746) );
  AND U1559 ( .A(n87), .B(n1753), .Z(n1755) );
  XNOR U1560 ( .A(n1754), .B(n1751), .Z(n1753) );
  XOR U1561 ( .A(n1756), .B(n1757), .Z(n1751) );
  AND U1562 ( .A(n90), .B(n1758), .Z(n1757) );
  XOR U1563 ( .A(p_input[86]), .B(n1756), .Z(n1758) );
  XOR U1564 ( .A(n1759), .B(n1760), .Z(n1756) );
  AND U1565 ( .A(n94), .B(n1761), .Z(n1760) );
  XOR U1566 ( .A(n1762), .B(n1763), .Z(n1754) );
  AND U1567 ( .A(n98), .B(n1761), .Z(n1763) );
  XNOR U1568 ( .A(n1762), .B(n1759), .Z(n1761) );
  XOR U1569 ( .A(n1764), .B(n1765), .Z(n1759) );
  AND U1570 ( .A(n101), .B(n1766), .Z(n1765) );
  XOR U1571 ( .A(p_input[102]), .B(n1764), .Z(n1766) );
  XOR U1572 ( .A(n1767), .B(n1768), .Z(n1764) );
  AND U1573 ( .A(n105), .B(n1769), .Z(n1768) );
  XOR U1574 ( .A(n1770), .B(n1771), .Z(n1762) );
  AND U1575 ( .A(n109), .B(n1769), .Z(n1771) );
  XNOR U1576 ( .A(n1770), .B(n1767), .Z(n1769) );
  XOR U1577 ( .A(n1772), .B(n1773), .Z(n1767) );
  AND U1578 ( .A(n112), .B(n1774), .Z(n1773) );
  XOR U1579 ( .A(p_input[118]), .B(n1772), .Z(n1774) );
  XOR U1580 ( .A(n1775), .B(n1776), .Z(n1772) );
  AND U1581 ( .A(n116), .B(n1777), .Z(n1776) );
  XOR U1582 ( .A(n1778), .B(n1779), .Z(n1770) );
  AND U1583 ( .A(n120), .B(n1777), .Z(n1779) );
  XNOR U1584 ( .A(n1778), .B(n1775), .Z(n1777) );
  XOR U1585 ( .A(n1780), .B(n1781), .Z(n1775) );
  AND U1586 ( .A(n123), .B(n1782), .Z(n1781) );
  XOR U1587 ( .A(p_input[134]), .B(n1780), .Z(n1782) );
  XOR U1588 ( .A(n1783), .B(n1784), .Z(n1780) );
  AND U1589 ( .A(n127), .B(n1785), .Z(n1784) );
  XOR U1590 ( .A(n1786), .B(n1787), .Z(n1778) );
  AND U1591 ( .A(n131), .B(n1785), .Z(n1787) );
  XNOR U1592 ( .A(n1786), .B(n1783), .Z(n1785) );
  XOR U1593 ( .A(n1788), .B(n1789), .Z(n1783) );
  AND U1594 ( .A(n134), .B(n1790), .Z(n1789) );
  XOR U1595 ( .A(p_input[150]), .B(n1788), .Z(n1790) );
  XOR U1596 ( .A(n1791), .B(n1792), .Z(n1788) );
  AND U1597 ( .A(n138), .B(n1793), .Z(n1792) );
  XOR U1598 ( .A(n1794), .B(n1795), .Z(n1786) );
  AND U1599 ( .A(n142), .B(n1793), .Z(n1795) );
  XNOR U1600 ( .A(n1794), .B(n1791), .Z(n1793) );
  XOR U1601 ( .A(n1796), .B(n1797), .Z(n1791) );
  AND U1602 ( .A(n145), .B(n1798), .Z(n1797) );
  XOR U1603 ( .A(p_input[166]), .B(n1796), .Z(n1798) );
  XOR U1604 ( .A(n1799), .B(n1800), .Z(n1796) );
  AND U1605 ( .A(n149), .B(n1801), .Z(n1800) );
  XOR U1606 ( .A(n1802), .B(n1803), .Z(n1794) );
  AND U1607 ( .A(n153), .B(n1801), .Z(n1803) );
  XNOR U1608 ( .A(n1802), .B(n1799), .Z(n1801) );
  XOR U1609 ( .A(n1804), .B(n1805), .Z(n1799) );
  AND U1610 ( .A(n156), .B(n1806), .Z(n1805) );
  XOR U1611 ( .A(p_input[182]), .B(n1804), .Z(n1806) );
  XOR U1612 ( .A(n1807), .B(n1808), .Z(n1804) );
  AND U1613 ( .A(n160), .B(n1809), .Z(n1808) );
  XOR U1614 ( .A(n1810), .B(n1811), .Z(n1802) );
  AND U1615 ( .A(n164), .B(n1809), .Z(n1811) );
  XNOR U1616 ( .A(n1810), .B(n1807), .Z(n1809) );
  XOR U1617 ( .A(n1812), .B(n1813), .Z(n1807) );
  AND U1618 ( .A(n167), .B(n1814), .Z(n1813) );
  XOR U1619 ( .A(p_input[198]), .B(n1812), .Z(n1814) );
  XOR U1620 ( .A(n1815), .B(n1816), .Z(n1812) );
  AND U1621 ( .A(n171), .B(n1817), .Z(n1816) );
  XOR U1622 ( .A(n1818), .B(n1819), .Z(n1810) );
  AND U1623 ( .A(n175), .B(n1817), .Z(n1819) );
  XNOR U1624 ( .A(n1818), .B(n1815), .Z(n1817) );
  XOR U1625 ( .A(n1820), .B(n1821), .Z(n1815) );
  AND U1626 ( .A(n178), .B(n1822), .Z(n1821) );
  XOR U1627 ( .A(p_input[214]), .B(n1820), .Z(n1822) );
  XOR U1628 ( .A(n1823), .B(n1824), .Z(n1820) );
  AND U1629 ( .A(n182), .B(n1825), .Z(n1824) );
  XOR U1630 ( .A(n1826), .B(n1827), .Z(n1818) );
  AND U1631 ( .A(n186), .B(n1825), .Z(n1827) );
  XNOR U1632 ( .A(n1826), .B(n1823), .Z(n1825) );
  XOR U1633 ( .A(n1828), .B(n1829), .Z(n1823) );
  AND U1634 ( .A(n189), .B(n1830), .Z(n1829) );
  XOR U1635 ( .A(p_input[230]), .B(n1828), .Z(n1830) );
  XOR U1636 ( .A(n1831), .B(n1832), .Z(n1828) );
  AND U1637 ( .A(n193), .B(n1833), .Z(n1832) );
  XOR U1638 ( .A(n1834), .B(n1835), .Z(n1826) );
  AND U1639 ( .A(n197), .B(n1833), .Z(n1835) );
  XNOR U1640 ( .A(n1834), .B(n1831), .Z(n1833) );
  XOR U1641 ( .A(n1836), .B(n1837), .Z(n1831) );
  AND U1642 ( .A(n200), .B(n1838), .Z(n1837) );
  XOR U1643 ( .A(p_input[246]), .B(n1836), .Z(n1838) );
  XOR U1644 ( .A(n1839), .B(n1840), .Z(n1836) );
  AND U1645 ( .A(n204), .B(n1841), .Z(n1840) );
  XOR U1646 ( .A(n1842), .B(n1843), .Z(n1834) );
  AND U1647 ( .A(n208), .B(n1841), .Z(n1843) );
  XNOR U1648 ( .A(n1842), .B(n1839), .Z(n1841) );
  XOR U1649 ( .A(n1844), .B(n1845), .Z(n1839) );
  AND U1650 ( .A(n211), .B(n1846), .Z(n1845) );
  XOR U1651 ( .A(p_input[262]), .B(n1844), .Z(n1846) );
  XOR U1652 ( .A(n1847), .B(n1848), .Z(n1844) );
  AND U1653 ( .A(n215), .B(n1849), .Z(n1848) );
  XOR U1654 ( .A(n1850), .B(n1851), .Z(n1842) );
  AND U1655 ( .A(n219), .B(n1849), .Z(n1851) );
  XNOR U1656 ( .A(n1850), .B(n1847), .Z(n1849) );
  XOR U1657 ( .A(n1852), .B(n1853), .Z(n1847) );
  AND U1658 ( .A(n222), .B(n1854), .Z(n1853) );
  XOR U1659 ( .A(p_input[278]), .B(n1852), .Z(n1854) );
  XOR U1660 ( .A(n1855), .B(n1856), .Z(n1852) );
  AND U1661 ( .A(n226), .B(n1857), .Z(n1856) );
  XOR U1662 ( .A(n1858), .B(n1859), .Z(n1850) );
  AND U1663 ( .A(n230), .B(n1857), .Z(n1859) );
  XNOR U1664 ( .A(n1858), .B(n1855), .Z(n1857) );
  XOR U1665 ( .A(n1860), .B(n1861), .Z(n1855) );
  AND U1666 ( .A(n233), .B(n1862), .Z(n1861) );
  XOR U1667 ( .A(p_input[294]), .B(n1860), .Z(n1862) );
  XOR U1668 ( .A(n1863), .B(n1864), .Z(n1860) );
  AND U1669 ( .A(n237), .B(n1865), .Z(n1864) );
  XOR U1670 ( .A(n1866), .B(n1867), .Z(n1858) );
  AND U1671 ( .A(n241), .B(n1865), .Z(n1867) );
  XNOR U1672 ( .A(n1866), .B(n1863), .Z(n1865) );
  XOR U1673 ( .A(n1868), .B(n1869), .Z(n1863) );
  AND U1674 ( .A(n244), .B(n1870), .Z(n1869) );
  XOR U1675 ( .A(p_input[310]), .B(n1868), .Z(n1870) );
  XOR U1676 ( .A(n1871), .B(n1872), .Z(n1868) );
  AND U1677 ( .A(n248), .B(n1873), .Z(n1872) );
  XOR U1678 ( .A(n1874), .B(n1875), .Z(n1866) );
  AND U1679 ( .A(n252), .B(n1873), .Z(n1875) );
  XNOR U1680 ( .A(n1874), .B(n1871), .Z(n1873) );
  XOR U1681 ( .A(n1876), .B(n1877), .Z(n1871) );
  AND U1682 ( .A(n255), .B(n1878), .Z(n1877) );
  XOR U1683 ( .A(p_input[326]), .B(n1876), .Z(n1878) );
  XOR U1684 ( .A(n1879), .B(n1880), .Z(n1876) );
  AND U1685 ( .A(n259), .B(n1881), .Z(n1880) );
  XOR U1686 ( .A(n1882), .B(n1883), .Z(n1874) );
  AND U1687 ( .A(n263), .B(n1881), .Z(n1883) );
  XNOR U1688 ( .A(n1882), .B(n1879), .Z(n1881) );
  XOR U1689 ( .A(n1884), .B(n1885), .Z(n1879) );
  AND U1690 ( .A(n266), .B(n1886), .Z(n1885) );
  XOR U1691 ( .A(p_input[342]), .B(n1884), .Z(n1886) );
  XOR U1692 ( .A(n1887), .B(n1888), .Z(n1884) );
  AND U1693 ( .A(n270), .B(n1889), .Z(n1888) );
  XOR U1694 ( .A(n1890), .B(n1891), .Z(n1882) );
  AND U1695 ( .A(n274), .B(n1889), .Z(n1891) );
  XNOR U1696 ( .A(n1890), .B(n1887), .Z(n1889) );
  XOR U1697 ( .A(n1892), .B(n1893), .Z(n1887) );
  AND U1698 ( .A(n277), .B(n1894), .Z(n1893) );
  XOR U1699 ( .A(p_input[358]), .B(n1892), .Z(n1894) );
  XOR U1700 ( .A(n1895), .B(n1896), .Z(n1892) );
  AND U1701 ( .A(n281), .B(n1897), .Z(n1896) );
  XOR U1702 ( .A(n1898), .B(n1899), .Z(n1890) );
  AND U1703 ( .A(n285), .B(n1897), .Z(n1899) );
  XNOR U1704 ( .A(n1898), .B(n1895), .Z(n1897) );
  XOR U1705 ( .A(n1900), .B(n1901), .Z(n1895) );
  AND U1706 ( .A(n288), .B(n1902), .Z(n1901) );
  XOR U1707 ( .A(p_input[374]), .B(n1900), .Z(n1902) );
  XOR U1708 ( .A(n1903), .B(n1904), .Z(n1900) );
  AND U1709 ( .A(n292), .B(n1905), .Z(n1904) );
  XOR U1710 ( .A(n1906), .B(n1907), .Z(n1898) );
  AND U1711 ( .A(n296), .B(n1905), .Z(n1907) );
  XNOR U1712 ( .A(n1906), .B(n1903), .Z(n1905) );
  XOR U1713 ( .A(n1908), .B(n1909), .Z(n1903) );
  AND U1714 ( .A(n299), .B(n1910), .Z(n1909) );
  XOR U1715 ( .A(p_input[390]), .B(n1908), .Z(n1910) );
  XOR U1716 ( .A(n1911), .B(n1912), .Z(n1908) );
  AND U1717 ( .A(n303), .B(n1913), .Z(n1912) );
  XOR U1718 ( .A(n1914), .B(n1915), .Z(n1906) );
  AND U1719 ( .A(n307), .B(n1913), .Z(n1915) );
  XNOR U1720 ( .A(n1914), .B(n1911), .Z(n1913) );
  XOR U1721 ( .A(n1916), .B(n1917), .Z(n1911) );
  AND U1722 ( .A(n310), .B(n1918), .Z(n1917) );
  XOR U1723 ( .A(p_input[406]), .B(n1916), .Z(n1918) );
  XOR U1724 ( .A(n1919), .B(n1920), .Z(n1916) );
  AND U1725 ( .A(n314), .B(n1921), .Z(n1920) );
  XOR U1726 ( .A(n1922), .B(n1923), .Z(n1914) );
  AND U1727 ( .A(n318), .B(n1921), .Z(n1923) );
  XNOR U1728 ( .A(n1922), .B(n1919), .Z(n1921) );
  XOR U1729 ( .A(n1924), .B(n1925), .Z(n1919) );
  AND U1730 ( .A(n321), .B(n1926), .Z(n1925) );
  XOR U1731 ( .A(p_input[422]), .B(n1924), .Z(n1926) );
  XOR U1732 ( .A(n1927), .B(n1928), .Z(n1924) );
  AND U1733 ( .A(n325), .B(n1929), .Z(n1928) );
  XOR U1734 ( .A(n1930), .B(n1931), .Z(n1922) );
  AND U1735 ( .A(n329), .B(n1929), .Z(n1931) );
  XNOR U1736 ( .A(n1930), .B(n1927), .Z(n1929) );
  XOR U1737 ( .A(n1932), .B(n1933), .Z(n1927) );
  AND U1738 ( .A(n332), .B(n1934), .Z(n1933) );
  XOR U1739 ( .A(p_input[438]), .B(n1932), .Z(n1934) );
  XOR U1740 ( .A(n1935), .B(n1936), .Z(n1932) );
  AND U1741 ( .A(n336), .B(n1937), .Z(n1936) );
  XOR U1742 ( .A(n1938), .B(n1939), .Z(n1930) );
  AND U1743 ( .A(n340), .B(n1937), .Z(n1939) );
  XNOR U1744 ( .A(n1938), .B(n1935), .Z(n1937) );
  XOR U1745 ( .A(n1940), .B(n1941), .Z(n1935) );
  AND U1746 ( .A(n343), .B(n1942), .Z(n1941) );
  XOR U1747 ( .A(p_input[454]), .B(n1940), .Z(n1942) );
  XOR U1748 ( .A(n1943), .B(n1944), .Z(n1940) );
  AND U1749 ( .A(n347), .B(n1945), .Z(n1944) );
  XOR U1750 ( .A(n1946), .B(n1947), .Z(n1938) );
  AND U1751 ( .A(n351), .B(n1945), .Z(n1947) );
  XNOR U1752 ( .A(n1946), .B(n1943), .Z(n1945) );
  XOR U1753 ( .A(n1948), .B(n1949), .Z(n1943) );
  AND U1754 ( .A(n354), .B(n1950), .Z(n1949) );
  XOR U1755 ( .A(p_input[470]), .B(n1948), .Z(n1950) );
  XOR U1756 ( .A(n1951), .B(n1952), .Z(n1948) );
  AND U1757 ( .A(n358), .B(n1953), .Z(n1952) );
  XOR U1758 ( .A(n1954), .B(n1955), .Z(n1946) );
  AND U1759 ( .A(n362), .B(n1953), .Z(n1955) );
  XNOR U1760 ( .A(n1954), .B(n1951), .Z(n1953) );
  XOR U1761 ( .A(n1956), .B(n1957), .Z(n1951) );
  AND U1762 ( .A(n365), .B(n1958), .Z(n1957) );
  XOR U1763 ( .A(p_input[486]), .B(n1956), .Z(n1958) );
  XOR U1764 ( .A(n1959), .B(n1960), .Z(n1956) );
  AND U1765 ( .A(n369), .B(n1961), .Z(n1960) );
  XOR U1766 ( .A(n1962), .B(n1963), .Z(n1954) );
  AND U1767 ( .A(n373), .B(n1961), .Z(n1963) );
  XNOR U1768 ( .A(n1962), .B(n1959), .Z(n1961) );
  XOR U1769 ( .A(n1964), .B(n1965), .Z(n1959) );
  AND U1770 ( .A(n376), .B(n1966), .Z(n1965) );
  XOR U1771 ( .A(p_input[502]), .B(n1964), .Z(n1966) );
  XOR U1772 ( .A(n1967), .B(n1968), .Z(n1964) );
  AND U1773 ( .A(n380), .B(n1969), .Z(n1968) );
  XOR U1774 ( .A(n1970), .B(n1971), .Z(n1962) );
  AND U1775 ( .A(n384), .B(n1969), .Z(n1971) );
  XNOR U1776 ( .A(n1970), .B(n1967), .Z(n1969) );
  XOR U1777 ( .A(n1972), .B(n1973), .Z(n1967) );
  AND U1778 ( .A(n387), .B(n1974), .Z(n1973) );
  XOR U1779 ( .A(p_input[518]), .B(n1972), .Z(n1974) );
  XOR U1780 ( .A(n1975), .B(n1976), .Z(n1972) );
  AND U1781 ( .A(n391), .B(n1977), .Z(n1976) );
  XOR U1782 ( .A(n1978), .B(n1979), .Z(n1970) );
  AND U1783 ( .A(n395), .B(n1977), .Z(n1979) );
  XNOR U1784 ( .A(n1978), .B(n1975), .Z(n1977) );
  XOR U1785 ( .A(n1980), .B(n1981), .Z(n1975) );
  AND U1786 ( .A(n398), .B(n1982), .Z(n1981) );
  XOR U1787 ( .A(p_input[534]), .B(n1980), .Z(n1982) );
  XOR U1788 ( .A(n1983), .B(n1984), .Z(n1980) );
  AND U1789 ( .A(n402), .B(n1985), .Z(n1984) );
  XOR U1790 ( .A(n1986), .B(n1987), .Z(n1978) );
  AND U1791 ( .A(n406), .B(n1985), .Z(n1987) );
  XNOR U1792 ( .A(n1986), .B(n1983), .Z(n1985) );
  XOR U1793 ( .A(n1988), .B(n1989), .Z(n1983) );
  AND U1794 ( .A(n409), .B(n1990), .Z(n1989) );
  XOR U1795 ( .A(p_input[550]), .B(n1988), .Z(n1990) );
  XOR U1796 ( .A(n1991), .B(n1992), .Z(n1988) );
  AND U1797 ( .A(n413), .B(n1993), .Z(n1992) );
  XOR U1798 ( .A(n1994), .B(n1995), .Z(n1986) );
  AND U1799 ( .A(n417), .B(n1993), .Z(n1995) );
  XNOR U1800 ( .A(n1994), .B(n1991), .Z(n1993) );
  XOR U1801 ( .A(n1996), .B(n1997), .Z(n1991) );
  AND U1802 ( .A(n420), .B(n1998), .Z(n1997) );
  XOR U1803 ( .A(p_input[566]), .B(n1996), .Z(n1998) );
  XOR U1804 ( .A(n1999), .B(n2000), .Z(n1996) );
  AND U1805 ( .A(n424), .B(n2001), .Z(n2000) );
  XOR U1806 ( .A(n2002), .B(n2003), .Z(n1994) );
  AND U1807 ( .A(n428), .B(n2001), .Z(n2003) );
  XNOR U1808 ( .A(n2002), .B(n1999), .Z(n2001) );
  XOR U1809 ( .A(n2004), .B(n2005), .Z(n1999) );
  AND U1810 ( .A(n431), .B(n2006), .Z(n2005) );
  XOR U1811 ( .A(p_input[582]), .B(n2004), .Z(n2006) );
  XOR U1812 ( .A(n2007), .B(n2008), .Z(n2004) );
  AND U1813 ( .A(n435), .B(n2009), .Z(n2008) );
  XOR U1814 ( .A(n2010), .B(n2011), .Z(n2002) );
  AND U1815 ( .A(n439), .B(n2009), .Z(n2011) );
  XNOR U1816 ( .A(n2010), .B(n2007), .Z(n2009) );
  XOR U1817 ( .A(n2012), .B(n2013), .Z(n2007) );
  AND U1818 ( .A(n442), .B(n2014), .Z(n2013) );
  XOR U1819 ( .A(p_input[598]), .B(n2012), .Z(n2014) );
  XOR U1820 ( .A(n2015), .B(n2016), .Z(n2012) );
  AND U1821 ( .A(n446), .B(n2017), .Z(n2016) );
  XOR U1822 ( .A(n2018), .B(n2019), .Z(n2010) );
  AND U1823 ( .A(n450), .B(n2017), .Z(n2019) );
  XNOR U1824 ( .A(n2018), .B(n2015), .Z(n2017) );
  XOR U1825 ( .A(n2020), .B(n2021), .Z(n2015) );
  AND U1826 ( .A(n453), .B(n2022), .Z(n2021) );
  XOR U1827 ( .A(p_input[614]), .B(n2020), .Z(n2022) );
  XOR U1828 ( .A(n2023), .B(n2024), .Z(n2020) );
  AND U1829 ( .A(n457), .B(n2025), .Z(n2024) );
  XOR U1830 ( .A(n2026), .B(n2027), .Z(n2018) );
  AND U1831 ( .A(n461), .B(n2025), .Z(n2027) );
  XNOR U1832 ( .A(n2026), .B(n2023), .Z(n2025) );
  XOR U1833 ( .A(n2028), .B(n2029), .Z(n2023) );
  AND U1834 ( .A(n464), .B(n2030), .Z(n2029) );
  XOR U1835 ( .A(p_input[630]), .B(n2028), .Z(n2030) );
  XOR U1836 ( .A(n2031), .B(n2032), .Z(n2028) );
  AND U1837 ( .A(n468), .B(n2033), .Z(n2032) );
  XOR U1838 ( .A(n2034), .B(n2035), .Z(n2026) );
  AND U1839 ( .A(n472), .B(n2033), .Z(n2035) );
  XNOR U1840 ( .A(n2034), .B(n2031), .Z(n2033) );
  XOR U1841 ( .A(n2036), .B(n2037), .Z(n2031) );
  AND U1842 ( .A(n475), .B(n2038), .Z(n2037) );
  XOR U1843 ( .A(p_input[646]), .B(n2036), .Z(n2038) );
  XOR U1844 ( .A(n2039), .B(n2040), .Z(n2036) );
  AND U1845 ( .A(n479), .B(n2041), .Z(n2040) );
  XOR U1846 ( .A(n2042), .B(n2043), .Z(n2034) );
  AND U1847 ( .A(n483), .B(n2041), .Z(n2043) );
  XNOR U1848 ( .A(n2042), .B(n2039), .Z(n2041) );
  XOR U1849 ( .A(n2044), .B(n2045), .Z(n2039) );
  AND U1850 ( .A(n486), .B(n2046), .Z(n2045) );
  XOR U1851 ( .A(p_input[662]), .B(n2044), .Z(n2046) );
  XOR U1852 ( .A(n2047), .B(n2048), .Z(n2044) );
  AND U1853 ( .A(n490), .B(n2049), .Z(n2048) );
  XOR U1854 ( .A(n2050), .B(n2051), .Z(n2042) );
  AND U1855 ( .A(n494), .B(n2049), .Z(n2051) );
  XNOR U1856 ( .A(n2050), .B(n2047), .Z(n2049) );
  XOR U1857 ( .A(n2052), .B(n2053), .Z(n2047) );
  AND U1858 ( .A(n497), .B(n2054), .Z(n2053) );
  XOR U1859 ( .A(p_input[678]), .B(n2052), .Z(n2054) );
  XOR U1860 ( .A(n2055), .B(n2056), .Z(n2052) );
  AND U1861 ( .A(n501), .B(n2057), .Z(n2056) );
  XOR U1862 ( .A(n2058), .B(n2059), .Z(n2050) );
  AND U1863 ( .A(n505), .B(n2057), .Z(n2059) );
  XNOR U1864 ( .A(n2058), .B(n2055), .Z(n2057) );
  XOR U1865 ( .A(n2060), .B(n2061), .Z(n2055) );
  AND U1866 ( .A(n508), .B(n2062), .Z(n2061) );
  XOR U1867 ( .A(p_input[694]), .B(n2060), .Z(n2062) );
  XOR U1868 ( .A(n2063), .B(n2064), .Z(n2060) );
  AND U1869 ( .A(n512), .B(n2065), .Z(n2064) );
  XOR U1870 ( .A(n2066), .B(n2067), .Z(n2058) );
  AND U1871 ( .A(n516), .B(n2065), .Z(n2067) );
  XNOR U1872 ( .A(n2066), .B(n2063), .Z(n2065) );
  XOR U1873 ( .A(n2068), .B(n2069), .Z(n2063) );
  AND U1874 ( .A(n519), .B(n2070), .Z(n2069) );
  XOR U1875 ( .A(p_input[710]), .B(n2068), .Z(n2070) );
  XOR U1876 ( .A(n2071), .B(n2072), .Z(n2068) );
  AND U1877 ( .A(n523), .B(n2073), .Z(n2072) );
  XOR U1878 ( .A(n2074), .B(n2075), .Z(n2066) );
  AND U1879 ( .A(n527), .B(n2073), .Z(n2075) );
  XNOR U1880 ( .A(n2074), .B(n2071), .Z(n2073) );
  XOR U1881 ( .A(n2076), .B(n2077), .Z(n2071) );
  AND U1882 ( .A(n530), .B(n2078), .Z(n2077) );
  XOR U1883 ( .A(p_input[726]), .B(n2076), .Z(n2078) );
  XOR U1884 ( .A(n2079), .B(n2080), .Z(n2076) );
  AND U1885 ( .A(n534), .B(n2081), .Z(n2080) );
  XOR U1886 ( .A(n2082), .B(n2083), .Z(n2074) );
  AND U1887 ( .A(n538), .B(n2081), .Z(n2083) );
  XNOR U1888 ( .A(n2082), .B(n2079), .Z(n2081) );
  XOR U1889 ( .A(n2084), .B(n2085), .Z(n2079) );
  AND U1890 ( .A(n541), .B(n2086), .Z(n2085) );
  XOR U1891 ( .A(p_input[742]), .B(n2084), .Z(n2086) );
  XOR U1892 ( .A(n2087), .B(n2088), .Z(n2084) );
  AND U1893 ( .A(n545), .B(n2089), .Z(n2088) );
  XOR U1894 ( .A(n2090), .B(n2091), .Z(n2082) );
  AND U1895 ( .A(n549), .B(n2089), .Z(n2091) );
  XNOR U1896 ( .A(n2090), .B(n2087), .Z(n2089) );
  XOR U1897 ( .A(n2092), .B(n2093), .Z(n2087) );
  AND U1898 ( .A(n552), .B(n2094), .Z(n2093) );
  XOR U1899 ( .A(p_input[758]), .B(n2092), .Z(n2094) );
  XOR U1900 ( .A(n2095), .B(n2096), .Z(n2092) );
  AND U1901 ( .A(n556), .B(n2097), .Z(n2096) );
  XOR U1902 ( .A(n2098), .B(n2099), .Z(n2090) );
  AND U1903 ( .A(n560), .B(n2097), .Z(n2099) );
  XNOR U1904 ( .A(n2098), .B(n2095), .Z(n2097) );
  XOR U1905 ( .A(n2100), .B(n2101), .Z(n2095) );
  AND U1906 ( .A(n563), .B(n2102), .Z(n2101) );
  XOR U1907 ( .A(p_input[774]), .B(n2100), .Z(n2102) );
  XOR U1908 ( .A(n2103), .B(n2104), .Z(n2100) );
  AND U1909 ( .A(n567), .B(n2105), .Z(n2104) );
  XOR U1910 ( .A(n2106), .B(n2107), .Z(n2098) );
  AND U1911 ( .A(n571), .B(n2105), .Z(n2107) );
  XNOR U1912 ( .A(n2106), .B(n2103), .Z(n2105) );
  XOR U1913 ( .A(n2108), .B(n2109), .Z(n2103) );
  AND U1914 ( .A(n574), .B(n2110), .Z(n2109) );
  XOR U1915 ( .A(p_input[790]), .B(n2108), .Z(n2110) );
  XOR U1916 ( .A(n2111), .B(n2112), .Z(n2108) );
  AND U1917 ( .A(n578), .B(n2113), .Z(n2112) );
  XOR U1918 ( .A(n2114), .B(n2115), .Z(n2106) );
  AND U1919 ( .A(n582), .B(n2113), .Z(n2115) );
  XNOR U1920 ( .A(n2114), .B(n2111), .Z(n2113) );
  XOR U1921 ( .A(n2116), .B(n2117), .Z(n2111) );
  AND U1922 ( .A(n585), .B(n2118), .Z(n2117) );
  XOR U1923 ( .A(p_input[806]), .B(n2116), .Z(n2118) );
  XOR U1924 ( .A(n2119), .B(n2120), .Z(n2116) );
  AND U1925 ( .A(n589), .B(n2121), .Z(n2120) );
  XOR U1926 ( .A(n2122), .B(n2123), .Z(n2114) );
  AND U1927 ( .A(n593), .B(n2121), .Z(n2123) );
  XNOR U1928 ( .A(n2122), .B(n2119), .Z(n2121) );
  XOR U1929 ( .A(n2124), .B(n2125), .Z(n2119) );
  AND U1930 ( .A(n596), .B(n2126), .Z(n2125) );
  XOR U1931 ( .A(p_input[822]), .B(n2124), .Z(n2126) );
  XOR U1932 ( .A(n2127), .B(n2128), .Z(n2124) );
  AND U1933 ( .A(n600), .B(n2129), .Z(n2128) );
  XOR U1934 ( .A(n2130), .B(n2131), .Z(n2122) );
  AND U1935 ( .A(n604), .B(n2129), .Z(n2131) );
  XNOR U1936 ( .A(n2130), .B(n2127), .Z(n2129) );
  XOR U1937 ( .A(n2132), .B(n2133), .Z(n2127) );
  AND U1938 ( .A(n607), .B(n2134), .Z(n2133) );
  XOR U1939 ( .A(p_input[838]), .B(n2132), .Z(n2134) );
  XOR U1940 ( .A(n2135), .B(n2136), .Z(n2132) );
  AND U1941 ( .A(n611), .B(n2137), .Z(n2136) );
  XOR U1942 ( .A(n2138), .B(n2139), .Z(n2130) );
  AND U1943 ( .A(n615), .B(n2137), .Z(n2139) );
  XNOR U1944 ( .A(n2138), .B(n2135), .Z(n2137) );
  XOR U1945 ( .A(n2140), .B(n2141), .Z(n2135) );
  AND U1946 ( .A(n618), .B(n2142), .Z(n2141) );
  XOR U1947 ( .A(p_input[854]), .B(n2140), .Z(n2142) );
  XOR U1948 ( .A(n2143), .B(n2144), .Z(n2140) );
  AND U1949 ( .A(n622), .B(n2145), .Z(n2144) );
  XOR U1950 ( .A(n2146), .B(n2147), .Z(n2138) );
  AND U1951 ( .A(n626), .B(n2145), .Z(n2147) );
  XNOR U1952 ( .A(n2146), .B(n2143), .Z(n2145) );
  XOR U1953 ( .A(n2148), .B(n2149), .Z(n2143) );
  AND U1954 ( .A(n629), .B(n2150), .Z(n2149) );
  XOR U1955 ( .A(p_input[870]), .B(n2148), .Z(n2150) );
  XOR U1956 ( .A(n2151), .B(n2152), .Z(n2148) );
  AND U1957 ( .A(n633), .B(n2153), .Z(n2152) );
  XOR U1958 ( .A(n2154), .B(n2155), .Z(n2146) );
  AND U1959 ( .A(n637), .B(n2153), .Z(n2155) );
  XNOR U1960 ( .A(n2154), .B(n2151), .Z(n2153) );
  XOR U1961 ( .A(n2156), .B(n2157), .Z(n2151) );
  AND U1962 ( .A(n640), .B(n2158), .Z(n2157) );
  XOR U1963 ( .A(p_input[886]), .B(n2156), .Z(n2158) );
  XOR U1964 ( .A(n2159), .B(n2160), .Z(n2156) );
  AND U1965 ( .A(n644), .B(n2161), .Z(n2160) );
  XOR U1966 ( .A(n2162), .B(n2163), .Z(n2154) );
  AND U1967 ( .A(n648), .B(n2161), .Z(n2163) );
  XNOR U1968 ( .A(n2162), .B(n2159), .Z(n2161) );
  XOR U1969 ( .A(n2164), .B(n2165), .Z(n2159) );
  AND U1970 ( .A(n651), .B(n2166), .Z(n2165) );
  XOR U1971 ( .A(p_input[902]), .B(n2164), .Z(n2166) );
  XOR U1972 ( .A(n2167), .B(n2168), .Z(n2164) );
  AND U1973 ( .A(n655), .B(n2169), .Z(n2168) );
  XOR U1974 ( .A(n2170), .B(n2171), .Z(n2162) );
  AND U1975 ( .A(n659), .B(n2169), .Z(n2171) );
  XNOR U1976 ( .A(n2170), .B(n2167), .Z(n2169) );
  XOR U1977 ( .A(n2172), .B(n2173), .Z(n2167) );
  AND U1978 ( .A(n662), .B(n2174), .Z(n2173) );
  XOR U1979 ( .A(p_input[918]), .B(n2172), .Z(n2174) );
  XOR U1980 ( .A(n2175), .B(n2176), .Z(n2172) );
  AND U1981 ( .A(n666), .B(n2177), .Z(n2176) );
  XOR U1982 ( .A(n2178), .B(n2179), .Z(n2170) );
  AND U1983 ( .A(n670), .B(n2177), .Z(n2179) );
  XNOR U1984 ( .A(n2178), .B(n2175), .Z(n2177) );
  XOR U1985 ( .A(n2180), .B(n2181), .Z(n2175) );
  AND U1986 ( .A(n673), .B(n2182), .Z(n2181) );
  XOR U1987 ( .A(p_input[934]), .B(n2180), .Z(n2182) );
  XOR U1988 ( .A(n2183), .B(n2184), .Z(n2180) );
  AND U1989 ( .A(n677), .B(n2185), .Z(n2184) );
  XOR U1990 ( .A(n2186), .B(n2187), .Z(n2178) );
  AND U1991 ( .A(n681), .B(n2185), .Z(n2187) );
  XNOR U1992 ( .A(n2186), .B(n2183), .Z(n2185) );
  XOR U1993 ( .A(n2188), .B(n2189), .Z(n2183) );
  AND U1994 ( .A(n684), .B(n2190), .Z(n2189) );
  XOR U1995 ( .A(p_input[950]), .B(n2188), .Z(n2190) );
  XOR U1996 ( .A(n2191), .B(n2192), .Z(n2188) );
  AND U1997 ( .A(n688), .B(n2193), .Z(n2192) );
  XOR U1998 ( .A(n2194), .B(n2195), .Z(n2186) );
  AND U1999 ( .A(n692), .B(n2193), .Z(n2195) );
  XNOR U2000 ( .A(n2194), .B(n2191), .Z(n2193) );
  XOR U2001 ( .A(n2196), .B(n2197), .Z(n2191) );
  AND U2002 ( .A(n695), .B(n2198), .Z(n2197) );
  XOR U2003 ( .A(p_input[966]), .B(n2196), .Z(n2198) );
  XOR U2004 ( .A(n2199), .B(n2200), .Z(n2196) );
  AND U2005 ( .A(n699), .B(n2201), .Z(n2200) );
  XOR U2006 ( .A(n2202), .B(n2203), .Z(n2194) );
  AND U2007 ( .A(n703), .B(n2201), .Z(n2203) );
  XNOR U2008 ( .A(n2202), .B(n2199), .Z(n2201) );
  XOR U2009 ( .A(n2204), .B(n2205), .Z(n2199) );
  AND U2010 ( .A(n706), .B(n2206), .Z(n2205) );
  XOR U2011 ( .A(p_input[982]), .B(n2204), .Z(n2206) );
  XNOR U2012 ( .A(n2207), .B(n2208), .Z(n2204) );
  AND U2013 ( .A(n710), .B(n2209), .Z(n2208) );
  XNOR U2014 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n2210), .Z(n2202) );
  AND U2015 ( .A(n713), .B(n2209), .Z(n2210) );
  XOR U2016 ( .A(n2211), .B(n2207), .Z(n2209) );
  XOR U2017 ( .A(n9), .B(n2212), .Z(o[21]) );
  AND U2018 ( .A(n30), .B(n2213), .Z(n9) );
  XOR U2019 ( .A(n10), .B(n2212), .Z(n2213) );
  XOR U2020 ( .A(n2214), .B(n2215), .Z(n2212) );
  AND U2021 ( .A(n34), .B(n2216), .Z(n2215) );
  XOR U2022 ( .A(p_input[5]), .B(n2214), .Z(n2216) );
  XOR U2023 ( .A(n2217), .B(n2218), .Z(n2214) );
  AND U2024 ( .A(n38), .B(n2219), .Z(n2218) );
  XOR U2025 ( .A(n2220), .B(n2221), .Z(n10) );
  AND U2026 ( .A(n42), .B(n2219), .Z(n2221) );
  XNOR U2027 ( .A(n2222), .B(n2217), .Z(n2219) );
  XOR U2028 ( .A(n2223), .B(n2224), .Z(n2217) );
  AND U2029 ( .A(n46), .B(n2225), .Z(n2224) );
  XOR U2030 ( .A(p_input[21]), .B(n2223), .Z(n2225) );
  XOR U2031 ( .A(n2226), .B(n2227), .Z(n2223) );
  AND U2032 ( .A(n50), .B(n2228), .Z(n2227) );
  IV U2033 ( .A(n2220), .Z(n2222) );
  XNOR U2034 ( .A(n2229), .B(n2230), .Z(n2220) );
  AND U2035 ( .A(n54), .B(n2228), .Z(n2230) );
  XNOR U2036 ( .A(n2229), .B(n2226), .Z(n2228) );
  XOR U2037 ( .A(n2231), .B(n2232), .Z(n2226) );
  AND U2038 ( .A(n57), .B(n2233), .Z(n2232) );
  XOR U2039 ( .A(p_input[37]), .B(n2231), .Z(n2233) );
  XOR U2040 ( .A(n2234), .B(n2235), .Z(n2231) );
  AND U2041 ( .A(n61), .B(n2236), .Z(n2235) );
  XOR U2042 ( .A(n2237), .B(n2238), .Z(n2229) );
  AND U2043 ( .A(n65), .B(n2236), .Z(n2238) );
  XNOR U2044 ( .A(n2237), .B(n2234), .Z(n2236) );
  XOR U2045 ( .A(n2239), .B(n2240), .Z(n2234) );
  AND U2046 ( .A(n68), .B(n2241), .Z(n2240) );
  XOR U2047 ( .A(p_input[53]), .B(n2239), .Z(n2241) );
  XOR U2048 ( .A(n2242), .B(n2243), .Z(n2239) );
  AND U2049 ( .A(n72), .B(n2244), .Z(n2243) );
  XOR U2050 ( .A(n2245), .B(n2246), .Z(n2237) );
  AND U2051 ( .A(n76), .B(n2244), .Z(n2246) );
  XNOR U2052 ( .A(n2245), .B(n2242), .Z(n2244) );
  XOR U2053 ( .A(n2247), .B(n2248), .Z(n2242) );
  AND U2054 ( .A(n79), .B(n2249), .Z(n2248) );
  XOR U2055 ( .A(p_input[69]), .B(n2247), .Z(n2249) );
  XOR U2056 ( .A(n2250), .B(n2251), .Z(n2247) );
  AND U2057 ( .A(n83), .B(n2252), .Z(n2251) );
  XOR U2058 ( .A(n2253), .B(n2254), .Z(n2245) );
  AND U2059 ( .A(n87), .B(n2252), .Z(n2254) );
  XNOR U2060 ( .A(n2253), .B(n2250), .Z(n2252) );
  XOR U2061 ( .A(n2255), .B(n2256), .Z(n2250) );
  AND U2062 ( .A(n90), .B(n2257), .Z(n2256) );
  XOR U2063 ( .A(p_input[85]), .B(n2255), .Z(n2257) );
  XOR U2064 ( .A(n2258), .B(n2259), .Z(n2255) );
  AND U2065 ( .A(n94), .B(n2260), .Z(n2259) );
  XOR U2066 ( .A(n2261), .B(n2262), .Z(n2253) );
  AND U2067 ( .A(n98), .B(n2260), .Z(n2262) );
  XNOR U2068 ( .A(n2261), .B(n2258), .Z(n2260) );
  XOR U2069 ( .A(n2263), .B(n2264), .Z(n2258) );
  AND U2070 ( .A(n101), .B(n2265), .Z(n2264) );
  XOR U2071 ( .A(p_input[101]), .B(n2263), .Z(n2265) );
  XOR U2072 ( .A(n2266), .B(n2267), .Z(n2263) );
  AND U2073 ( .A(n105), .B(n2268), .Z(n2267) );
  XOR U2074 ( .A(n2269), .B(n2270), .Z(n2261) );
  AND U2075 ( .A(n109), .B(n2268), .Z(n2270) );
  XNOR U2076 ( .A(n2269), .B(n2266), .Z(n2268) );
  XOR U2077 ( .A(n2271), .B(n2272), .Z(n2266) );
  AND U2078 ( .A(n112), .B(n2273), .Z(n2272) );
  XOR U2079 ( .A(p_input[117]), .B(n2271), .Z(n2273) );
  XOR U2080 ( .A(n2274), .B(n2275), .Z(n2271) );
  AND U2081 ( .A(n116), .B(n2276), .Z(n2275) );
  XOR U2082 ( .A(n2277), .B(n2278), .Z(n2269) );
  AND U2083 ( .A(n120), .B(n2276), .Z(n2278) );
  XNOR U2084 ( .A(n2277), .B(n2274), .Z(n2276) );
  XOR U2085 ( .A(n2279), .B(n2280), .Z(n2274) );
  AND U2086 ( .A(n123), .B(n2281), .Z(n2280) );
  XOR U2087 ( .A(p_input[133]), .B(n2279), .Z(n2281) );
  XOR U2088 ( .A(n2282), .B(n2283), .Z(n2279) );
  AND U2089 ( .A(n127), .B(n2284), .Z(n2283) );
  XOR U2090 ( .A(n2285), .B(n2286), .Z(n2277) );
  AND U2091 ( .A(n131), .B(n2284), .Z(n2286) );
  XNOR U2092 ( .A(n2285), .B(n2282), .Z(n2284) );
  XOR U2093 ( .A(n2287), .B(n2288), .Z(n2282) );
  AND U2094 ( .A(n134), .B(n2289), .Z(n2288) );
  XOR U2095 ( .A(p_input[149]), .B(n2287), .Z(n2289) );
  XOR U2096 ( .A(n2290), .B(n2291), .Z(n2287) );
  AND U2097 ( .A(n138), .B(n2292), .Z(n2291) );
  XOR U2098 ( .A(n2293), .B(n2294), .Z(n2285) );
  AND U2099 ( .A(n142), .B(n2292), .Z(n2294) );
  XNOR U2100 ( .A(n2293), .B(n2290), .Z(n2292) );
  XOR U2101 ( .A(n2295), .B(n2296), .Z(n2290) );
  AND U2102 ( .A(n145), .B(n2297), .Z(n2296) );
  XOR U2103 ( .A(p_input[165]), .B(n2295), .Z(n2297) );
  XOR U2104 ( .A(n2298), .B(n2299), .Z(n2295) );
  AND U2105 ( .A(n149), .B(n2300), .Z(n2299) );
  XOR U2106 ( .A(n2301), .B(n2302), .Z(n2293) );
  AND U2107 ( .A(n153), .B(n2300), .Z(n2302) );
  XNOR U2108 ( .A(n2301), .B(n2298), .Z(n2300) );
  XOR U2109 ( .A(n2303), .B(n2304), .Z(n2298) );
  AND U2110 ( .A(n156), .B(n2305), .Z(n2304) );
  XOR U2111 ( .A(p_input[181]), .B(n2303), .Z(n2305) );
  XOR U2112 ( .A(n2306), .B(n2307), .Z(n2303) );
  AND U2113 ( .A(n160), .B(n2308), .Z(n2307) );
  XOR U2114 ( .A(n2309), .B(n2310), .Z(n2301) );
  AND U2115 ( .A(n164), .B(n2308), .Z(n2310) );
  XNOR U2116 ( .A(n2309), .B(n2306), .Z(n2308) );
  XOR U2117 ( .A(n2311), .B(n2312), .Z(n2306) );
  AND U2118 ( .A(n167), .B(n2313), .Z(n2312) );
  XOR U2119 ( .A(p_input[197]), .B(n2311), .Z(n2313) );
  XOR U2120 ( .A(n2314), .B(n2315), .Z(n2311) );
  AND U2121 ( .A(n171), .B(n2316), .Z(n2315) );
  XOR U2122 ( .A(n2317), .B(n2318), .Z(n2309) );
  AND U2123 ( .A(n175), .B(n2316), .Z(n2318) );
  XNOR U2124 ( .A(n2317), .B(n2314), .Z(n2316) );
  XOR U2125 ( .A(n2319), .B(n2320), .Z(n2314) );
  AND U2126 ( .A(n178), .B(n2321), .Z(n2320) );
  XOR U2127 ( .A(p_input[213]), .B(n2319), .Z(n2321) );
  XOR U2128 ( .A(n2322), .B(n2323), .Z(n2319) );
  AND U2129 ( .A(n182), .B(n2324), .Z(n2323) );
  XOR U2130 ( .A(n2325), .B(n2326), .Z(n2317) );
  AND U2131 ( .A(n186), .B(n2324), .Z(n2326) );
  XNOR U2132 ( .A(n2325), .B(n2322), .Z(n2324) );
  XOR U2133 ( .A(n2327), .B(n2328), .Z(n2322) );
  AND U2134 ( .A(n189), .B(n2329), .Z(n2328) );
  XOR U2135 ( .A(p_input[229]), .B(n2327), .Z(n2329) );
  XOR U2136 ( .A(n2330), .B(n2331), .Z(n2327) );
  AND U2137 ( .A(n193), .B(n2332), .Z(n2331) );
  XOR U2138 ( .A(n2333), .B(n2334), .Z(n2325) );
  AND U2139 ( .A(n197), .B(n2332), .Z(n2334) );
  XNOR U2140 ( .A(n2333), .B(n2330), .Z(n2332) );
  XOR U2141 ( .A(n2335), .B(n2336), .Z(n2330) );
  AND U2142 ( .A(n200), .B(n2337), .Z(n2336) );
  XOR U2143 ( .A(p_input[245]), .B(n2335), .Z(n2337) );
  XOR U2144 ( .A(n2338), .B(n2339), .Z(n2335) );
  AND U2145 ( .A(n204), .B(n2340), .Z(n2339) );
  XOR U2146 ( .A(n2341), .B(n2342), .Z(n2333) );
  AND U2147 ( .A(n208), .B(n2340), .Z(n2342) );
  XNOR U2148 ( .A(n2341), .B(n2338), .Z(n2340) );
  XOR U2149 ( .A(n2343), .B(n2344), .Z(n2338) );
  AND U2150 ( .A(n211), .B(n2345), .Z(n2344) );
  XOR U2151 ( .A(p_input[261]), .B(n2343), .Z(n2345) );
  XOR U2152 ( .A(n2346), .B(n2347), .Z(n2343) );
  AND U2153 ( .A(n215), .B(n2348), .Z(n2347) );
  XOR U2154 ( .A(n2349), .B(n2350), .Z(n2341) );
  AND U2155 ( .A(n219), .B(n2348), .Z(n2350) );
  XNOR U2156 ( .A(n2349), .B(n2346), .Z(n2348) );
  XOR U2157 ( .A(n2351), .B(n2352), .Z(n2346) );
  AND U2158 ( .A(n222), .B(n2353), .Z(n2352) );
  XOR U2159 ( .A(p_input[277]), .B(n2351), .Z(n2353) );
  XOR U2160 ( .A(n2354), .B(n2355), .Z(n2351) );
  AND U2161 ( .A(n226), .B(n2356), .Z(n2355) );
  XOR U2162 ( .A(n2357), .B(n2358), .Z(n2349) );
  AND U2163 ( .A(n230), .B(n2356), .Z(n2358) );
  XNOR U2164 ( .A(n2357), .B(n2354), .Z(n2356) );
  XOR U2165 ( .A(n2359), .B(n2360), .Z(n2354) );
  AND U2166 ( .A(n233), .B(n2361), .Z(n2360) );
  XOR U2167 ( .A(p_input[293]), .B(n2359), .Z(n2361) );
  XOR U2168 ( .A(n2362), .B(n2363), .Z(n2359) );
  AND U2169 ( .A(n237), .B(n2364), .Z(n2363) );
  XOR U2170 ( .A(n2365), .B(n2366), .Z(n2357) );
  AND U2171 ( .A(n241), .B(n2364), .Z(n2366) );
  XNOR U2172 ( .A(n2365), .B(n2362), .Z(n2364) );
  XOR U2173 ( .A(n2367), .B(n2368), .Z(n2362) );
  AND U2174 ( .A(n244), .B(n2369), .Z(n2368) );
  XOR U2175 ( .A(p_input[309]), .B(n2367), .Z(n2369) );
  XOR U2176 ( .A(n2370), .B(n2371), .Z(n2367) );
  AND U2177 ( .A(n248), .B(n2372), .Z(n2371) );
  XOR U2178 ( .A(n2373), .B(n2374), .Z(n2365) );
  AND U2179 ( .A(n252), .B(n2372), .Z(n2374) );
  XNOR U2180 ( .A(n2373), .B(n2370), .Z(n2372) );
  XOR U2181 ( .A(n2375), .B(n2376), .Z(n2370) );
  AND U2182 ( .A(n255), .B(n2377), .Z(n2376) );
  XOR U2183 ( .A(p_input[325]), .B(n2375), .Z(n2377) );
  XOR U2184 ( .A(n2378), .B(n2379), .Z(n2375) );
  AND U2185 ( .A(n259), .B(n2380), .Z(n2379) );
  XOR U2186 ( .A(n2381), .B(n2382), .Z(n2373) );
  AND U2187 ( .A(n263), .B(n2380), .Z(n2382) );
  XNOR U2188 ( .A(n2381), .B(n2378), .Z(n2380) );
  XOR U2189 ( .A(n2383), .B(n2384), .Z(n2378) );
  AND U2190 ( .A(n266), .B(n2385), .Z(n2384) );
  XOR U2191 ( .A(p_input[341]), .B(n2383), .Z(n2385) );
  XOR U2192 ( .A(n2386), .B(n2387), .Z(n2383) );
  AND U2193 ( .A(n270), .B(n2388), .Z(n2387) );
  XOR U2194 ( .A(n2389), .B(n2390), .Z(n2381) );
  AND U2195 ( .A(n274), .B(n2388), .Z(n2390) );
  XNOR U2196 ( .A(n2389), .B(n2386), .Z(n2388) );
  XOR U2197 ( .A(n2391), .B(n2392), .Z(n2386) );
  AND U2198 ( .A(n277), .B(n2393), .Z(n2392) );
  XOR U2199 ( .A(p_input[357]), .B(n2391), .Z(n2393) );
  XOR U2200 ( .A(n2394), .B(n2395), .Z(n2391) );
  AND U2201 ( .A(n281), .B(n2396), .Z(n2395) );
  XOR U2202 ( .A(n2397), .B(n2398), .Z(n2389) );
  AND U2203 ( .A(n285), .B(n2396), .Z(n2398) );
  XNOR U2204 ( .A(n2397), .B(n2394), .Z(n2396) );
  XOR U2205 ( .A(n2399), .B(n2400), .Z(n2394) );
  AND U2206 ( .A(n288), .B(n2401), .Z(n2400) );
  XOR U2207 ( .A(p_input[373]), .B(n2399), .Z(n2401) );
  XOR U2208 ( .A(n2402), .B(n2403), .Z(n2399) );
  AND U2209 ( .A(n292), .B(n2404), .Z(n2403) );
  XOR U2210 ( .A(n2405), .B(n2406), .Z(n2397) );
  AND U2211 ( .A(n296), .B(n2404), .Z(n2406) );
  XNOR U2212 ( .A(n2405), .B(n2402), .Z(n2404) );
  XOR U2213 ( .A(n2407), .B(n2408), .Z(n2402) );
  AND U2214 ( .A(n299), .B(n2409), .Z(n2408) );
  XOR U2215 ( .A(p_input[389]), .B(n2407), .Z(n2409) );
  XOR U2216 ( .A(n2410), .B(n2411), .Z(n2407) );
  AND U2217 ( .A(n303), .B(n2412), .Z(n2411) );
  XOR U2218 ( .A(n2413), .B(n2414), .Z(n2405) );
  AND U2219 ( .A(n307), .B(n2412), .Z(n2414) );
  XNOR U2220 ( .A(n2413), .B(n2410), .Z(n2412) );
  XOR U2221 ( .A(n2415), .B(n2416), .Z(n2410) );
  AND U2222 ( .A(n310), .B(n2417), .Z(n2416) );
  XOR U2223 ( .A(p_input[405]), .B(n2415), .Z(n2417) );
  XOR U2224 ( .A(n2418), .B(n2419), .Z(n2415) );
  AND U2225 ( .A(n314), .B(n2420), .Z(n2419) );
  XOR U2226 ( .A(n2421), .B(n2422), .Z(n2413) );
  AND U2227 ( .A(n318), .B(n2420), .Z(n2422) );
  XNOR U2228 ( .A(n2421), .B(n2418), .Z(n2420) );
  XOR U2229 ( .A(n2423), .B(n2424), .Z(n2418) );
  AND U2230 ( .A(n321), .B(n2425), .Z(n2424) );
  XOR U2231 ( .A(p_input[421]), .B(n2423), .Z(n2425) );
  XOR U2232 ( .A(n2426), .B(n2427), .Z(n2423) );
  AND U2233 ( .A(n325), .B(n2428), .Z(n2427) );
  XOR U2234 ( .A(n2429), .B(n2430), .Z(n2421) );
  AND U2235 ( .A(n329), .B(n2428), .Z(n2430) );
  XNOR U2236 ( .A(n2429), .B(n2426), .Z(n2428) );
  XOR U2237 ( .A(n2431), .B(n2432), .Z(n2426) );
  AND U2238 ( .A(n332), .B(n2433), .Z(n2432) );
  XOR U2239 ( .A(p_input[437]), .B(n2431), .Z(n2433) );
  XOR U2240 ( .A(n2434), .B(n2435), .Z(n2431) );
  AND U2241 ( .A(n336), .B(n2436), .Z(n2435) );
  XOR U2242 ( .A(n2437), .B(n2438), .Z(n2429) );
  AND U2243 ( .A(n340), .B(n2436), .Z(n2438) );
  XNOR U2244 ( .A(n2437), .B(n2434), .Z(n2436) );
  XOR U2245 ( .A(n2439), .B(n2440), .Z(n2434) );
  AND U2246 ( .A(n343), .B(n2441), .Z(n2440) );
  XOR U2247 ( .A(p_input[453]), .B(n2439), .Z(n2441) );
  XOR U2248 ( .A(n2442), .B(n2443), .Z(n2439) );
  AND U2249 ( .A(n347), .B(n2444), .Z(n2443) );
  XOR U2250 ( .A(n2445), .B(n2446), .Z(n2437) );
  AND U2251 ( .A(n351), .B(n2444), .Z(n2446) );
  XNOR U2252 ( .A(n2445), .B(n2442), .Z(n2444) );
  XOR U2253 ( .A(n2447), .B(n2448), .Z(n2442) );
  AND U2254 ( .A(n354), .B(n2449), .Z(n2448) );
  XOR U2255 ( .A(p_input[469]), .B(n2447), .Z(n2449) );
  XOR U2256 ( .A(n2450), .B(n2451), .Z(n2447) );
  AND U2257 ( .A(n358), .B(n2452), .Z(n2451) );
  XOR U2258 ( .A(n2453), .B(n2454), .Z(n2445) );
  AND U2259 ( .A(n362), .B(n2452), .Z(n2454) );
  XNOR U2260 ( .A(n2453), .B(n2450), .Z(n2452) );
  XOR U2261 ( .A(n2455), .B(n2456), .Z(n2450) );
  AND U2262 ( .A(n365), .B(n2457), .Z(n2456) );
  XOR U2263 ( .A(p_input[485]), .B(n2455), .Z(n2457) );
  XOR U2264 ( .A(n2458), .B(n2459), .Z(n2455) );
  AND U2265 ( .A(n369), .B(n2460), .Z(n2459) );
  XOR U2266 ( .A(n2461), .B(n2462), .Z(n2453) );
  AND U2267 ( .A(n373), .B(n2460), .Z(n2462) );
  XNOR U2268 ( .A(n2461), .B(n2458), .Z(n2460) );
  XOR U2269 ( .A(n2463), .B(n2464), .Z(n2458) );
  AND U2270 ( .A(n376), .B(n2465), .Z(n2464) );
  XOR U2271 ( .A(p_input[501]), .B(n2463), .Z(n2465) );
  XOR U2272 ( .A(n2466), .B(n2467), .Z(n2463) );
  AND U2273 ( .A(n380), .B(n2468), .Z(n2467) );
  XOR U2274 ( .A(n2469), .B(n2470), .Z(n2461) );
  AND U2275 ( .A(n384), .B(n2468), .Z(n2470) );
  XNOR U2276 ( .A(n2469), .B(n2466), .Z(n2468) );
  XOR U2277 ( .A(n2471), .B(n2472), .Z(n2466) );
  AND U2278 ( .A(n387), .B(n2473), .Z(n2472) );
  XOR U2279 ( .A(p_input[517]), .B(n2471), .Z(n2473) );
  XOR U2280 ( .A(n2474), .B(n2475), .Z(n2471) );
  AND U2281 ( .A(n391), .B(n2476), .Z(n2475) );
  XOR U2282 ( .A(n2477), .B(n2478), .Z(n2469) );
  AND U2283 ( .A(n395), .B(n2476), .Z(n2478) );
  XNOR U2284 ( .A(n2477), .B(n2474), .Z(n2476) );
  XOR U2285 ( .A(n2479), .B(n2480), .Z(n2474) );
  AND U2286 ( .A(n398), .B(n2481), .Z(n2480) );
  XOR U2287 ( .A(p_input[533]), .B(n2479), .Z(n2481) );
  XOR U2288 ( .A(n2482), .B(n2483), .Z(n2479) );
  AND U2289 ( .A(n402), .B(n2484), .Z(n2483) );
  XOR U2290 ( .A(n2485), .B(n2486), .Z(n2477) );
  AND U2291 ( .A(n406), .B(n2484), .Z(n2486) );
  XNOR U2292 ( .A(n2485), .B(n2482), .Z(n2484) );
  XOR U2293 ( .A(n2487), .B(n2488), .Z(n2482) );
  AND U2294 ( .A(n409), .B(n2489), .Z(n2488) );
  XOR U2295 ( .A(p_input[549]), .B(n2487), .Z(n2489) );
  XOR U2296 ( .A(n2490), .B(n2491), .Z(n2487) );
  AND U2297 ( .A(n413), .B(n2492), .Z(n2491) );
  XOR U2298 ( .A(n2493), .B(n2494), .Z(n2485) );
  AND U2299 ( .A(n417), .B(n2492), .Z(n2494) );
  XNOR U2300 ( .A(n2493), .B(n2490), .Z(n2492) );
  XOR U2301 ( .A(n2495), .B(n2496), .Z(n2490) );
  AND U2302 ( .A(n420), .B(n2497), .Z(n2496) );
  XOR U2303 ( .A(p_input[565]), .B(n2495), .Z(n2497) );
  XOR U2304 ( .A(n2498), .B(n2499), .Z(n2495) );
  AND U2305 ( .A(n424), .B(n2500), .Z(n2499) );
  XOR U2306 ( .A(n2501), .B(n2502), .Z(n2493) );
  AND U2307 ( .A(n428), .B(n2500), .Z(n2502) );
  XNOR U2308 ( .A(n2501), .B(n2498), .Z(n2500) );
  XOR U2309 ( .A(n2503), .B(n2504), .Z(n2498) );
  AND U2310 ( .A(n431), .B(n2505), .Z(n2504) );
  XOR U2311 ( .A(p_input[581]), .B(n2503), .Z(n2505) );
  XOR U2312 ( .A(n2506), .B(n2507), .Z(n2503) );
  AND U2313 ( .A(n435), .B(n2508), .Z(n2507) );
  XOR U2314 ( .A(n2509), .B(n2510), .Z(n2501) );
  AND U2315 ( .A(n439), .B(n2508), .Z(n2510) );
  XNOR U2316 ( .A(n2509), .B(n2506), .Z(n2508) );
  XOR U2317 ( .A(n2511), .B(n2512), .Z(n2506) );
  AND U2318 ( .A(n442), .B(n2513), .Z(n2512) );
  XOR U2319 ( .A(p_input[597]), .B(n2511), .Z(n2513) );
  XOR U2320 ( .A(n2514), .B(n2515), .Z(n2511) );
  AND U2321 ( .A(n446), .B(n2516), .Z(n2515) );
  XOR U2322 ( .A(n2517), .B(n2518), .Z(n2509) );
  AND U2323 ( .A(n450), .B(n2516), .Z(n2518) );
  XNOR U2324 ( .A(n2517), .B(n2514), .Z(n2516) );
  XOR U2325 ( .A(n2519), .B(n2520), .Z(n2514) );
  AND U2326 ( .A(n453), .B(n2521), .Z(n2520) );
  XOR U2327 ( .A(p_input[613]), .B(n2519), .Z(n2521) );
  XOR U2328 ( .A(n2522), .B(n2523), .Z(n2519) );
  AND U2329 ( .A(n457), .B(n2524), .Z(n2523) );
  XOR U2330 ( .A(n2525), .B(n2526), .Z(n2517) );
  AND U2331 ( .A(n461), .B(n2524), .Z(n2526) );
  XNOR U2332 ( .A(n2525), .B(n2522), .Z(n2524) );
  XOR U2333 ( .A(n2527), .B(n2528), .Z(n2522) );
  AND U2334 ( .A(n464), .B(n2529), .Z(n2528) );
  XOR U2335 ( .A(p_input[629]), .B(n2527), .Z(n2529) );
  XOR U2336 ( .A(n2530), .B(n2531), .Z(n2527) );
  AND U2337 ( .A(n468), .B(n2532), .Z(n2531) );
  XOR U2338 ( .A(n2533), .B(n2534), .Z(n2525) );
  AND U2339 ( .A(n472), .B(n2532), .Z(n2534) );
  XNOR U2340 ( .A(n2533), .B(n2530), .Z(n2532) );
  XOR U2341 ( .A(n2535), .B(n2536), .Z(n2530) );
  AND U2342 ( .A(n475), .B(n2537), .Z(n2536) );
  XOR U2343 ( .A(p_input[645]), .B(n2535), .Z(n2537) );
  XOR U2344 ( .A(n2538), .B(n2539), .Z(n2535) );
  AND U2345 ( .A(n479), .B(n2540), .Z(n2539) );
  XOR U2346 ( .A(n2541), .B(n2542), .Z(n2533) );
  AND U2347 ( .A(n483), .B(n2540), .Z(n2542) );
  XNOR U2348 ( .A(n2541), .B(n2538), .Z(n2540) );
  XOR U2349 ( .A(n2543), .B(n2544), .Z(n2538) );
  AND U2350 ( .A(n486), .B(n2545), .Z(n2544) );
  XOR U2351 ( .A(p_input[661]), .B(n2543), .Z(n2545) );
  XOR U2352 ( .A(n2546), .B(n2547), .Z(n2543) );
  AND U2353 ( .A(n490), .B(n2548), .Z(n2547) );
  XOR U2354 ( .A(n2549), .B(n2550), .Z(n2541) );
  AND U2355 ( .A(n494), .B(n2548), .Z(n2550) );
  XNOR U2356 ( .A(n2549), .B(n2546), .Z(n2548) );
  XOR U2357 ( .A(n2551), .B(n2552), .Z(n2546) );
  AND U2358 ( .A(n497), .B(n2553), .Z(n2552) );
  XOR U2359 ( .A(p_input[677]), .B(n2551), .Z(n2553) );
  XOR U2360 ( .A(n2554), .B(n2555), .Z(n2551) );
  AND U2361 ( .A(n501), .B(n2556), .Z(n2555) );
  XOR U2362 ( .A(n2557), .B(n2558), .Z(n2549) );
  AND U2363 ( .A(n505), .B(n2556), .Z(n2558) );
  XNOR U2364 ( .A(n2557), .B(n2554), .Z(n2556) );
  XOR U2365 ( .A(n2559), .B(n2560), .Z(n2554) );
  AND U2366 ( .A(n508), .B(n2561), .Z(n2560) );
  XOR U2367 ( .A(p_input[693]), .B(n2559), .Z(n2561) );
  XOR U2368 ( .A(n2562), .B(n2563), .Z(n2559) );
  AND U2369 ( .A(n512), .B(n2564), .Z(n2563) );
  XOR U2370 ( .A(n2565), .B(n2566), .Z(n2557) );
  AND U2371 ( .A(n516), .B(n2564), .Z(n2566) );
  XNOR U2372 ( .A(n2565), .B(n2562), .Z(n2564) );
  XOR U2373 ( .A(n2567), .B(n2568), .Z(n2562) );
  AND U2374 ( .A(n519), .B(n2569), .Z(n2568) );
  XOR U2375 ( .A(p_input[709]), .B(n2567), .Z(n2569) );
  XOR U2376 ( .A(n2570), .B(n2571), .Z(n2567) );
  AND U2377 ( .A(n523), .B(n2572), .Z(n2571) );
  XOR U2378 ( .A(n2573), .B(n2574), .Z(n2565) );
  AND U2379 ( .A(n527), .B(n2572), .Z(n2574) );
  XNOR U2380 ( .A(n2573), .B(n2570), .Z(n2572) );
  XOR U2381 ( .A(n2575), .B(n2576), .Z(n2570) );
  AND U2382 ( .A(n530), .B(n2577), .Z(n2576) );
  XOR U2383 ( .A(p_input[725]), .B(n2575), .Z(n2577) );
  XOR U2384 ( .A(n2578), .B(n2579), .Z(n2575) );
  AND U2385 ( .A(n534), .B(n2580), .Z(n2579) );
  XOR U2386 ( .A(n2581), .B(n2582), .Z(n2573) );
  AND U2387 ( .A(n538), .B(n2580), .Z(n2582) );
  XNOR U2388 ( .A(n2581), .B(n2578), .Z(n2580) );
  XOR U2389 ( .A(n2583), .B(n2584), .Z(n2578) );
  AND U2390 ( .A(n541), .B(n2585), .Z(n2584) );
  XOR U2391 ( .A(p_input[741]), .B(n2583), .Z(n2585) );
  XOR U2392 ( .A(n2586), .B(n2587), .Z(n2583) );
  AND U2393 ( .A(n545), .B(n2588), .Z(n2587) );
  XOR U2394 ( .A(n2589), .B(n2590), .Z(n2581) );
  AND U2395 ( .A(n549), .B(n2588), .Z(n2590) );
  XNOR U2396 ( .A(n2589), .B(n2586), .Z(n2588) );
  XOR U2397 ( .A(n2591), .B(n2592), .Z(n2586) );
  AND U2398 ( .A(n552), .B(n2593), .Z(n2592) );
  XOR U2399 ( .A(p_input[757]), .B(n2591), .Z(n2593) );
  XOR U2400 ( .A(n2594), .B(n2595), .Z(n2591) );
  AND U2401 ( .A(n556), .B(n2596), .Z(n2595) );
  XOR U2402 ( .A(n2597), .B(n2598), .Z(n2589) );
  AND U2403 ( .A(n560), .B(n2596), .Z(n2598) );
  XNOR U2404 ( .A(n2597), .B(n2594), .Z(n2596) );
  XOR U2405 ( .A(n2599), .B(n2600), .Z(n2594) );
  AND U2406 ( .A(n563), .B(n2601), .Z(n2600) );
  XOR U2407 ( .A(p_input[773]), .B(n2599), .Z(n2601) );
  XOR U2408 ( .A(n2602), .B(n2603), .Z(n2599) );
  AND U2409 ( .A(n567), .B(n2604), .Z(n2603) );
  XOR U2410 ( .A(n2605), .B(n2606), .Z(n2597) );
  AND U2411 ( .A(n571), .B(n2604), .Z(n2606) );
  XNOR U2412 ( .A(n2605), .B(n2602), .Z(n2604) );
  XOR U2413 ( .A(n2607), .B(n2608), .Z(n2602) );
  AND U2414 ( .A(n574), .B(n2609), .Z(n2608) );
  XOR U2415 ( .A(p_input[789]), .B(n2607), .Z(n2609) );
  XOR U2416 ( .A(n2610), .B(n2611), .Z(n2607) );
  AND U2417 ( .A(n578), .B(n2612), .Z(n2611) );
  XOR U2418 ( .A(n2613), .B(n2614), .Z(n2605) );
  AND U2419 ( .A(n582), .B(n2612), .Z(n2614) );
  XNOR U2420 ( .A(n2613), .B(n2610), .Z(n2612) );
  XOR U2421 ( .A(n2615), .B(n2616), .Z(n2610) );
  AND U2422 ( .A(n585), .B(n2617), .Z(n2616) );
  XOR U2423 ( .A(p_input[805]), .B(n2615), .Z(n2617) );
  XOR U2424 ( .A(n2618), .B(n2619), .Z(n2615) );
  AND U2425 ( .A(n589), .B(n2620), .Z(n2619) );
  XOR U2426 ( .A(n2621), .B(n2622), .Z(n2613) );
  AND U2427 ( .A(n593), .B(n2620), .Z(n2622) );
  XNOR U2428 ( .A(n2621), .B(n2618), .Z(n2620) );
  XOR U2429 ( .A(n2623), .B(n2624), .Z(n2618) );
  AND U2430 ( .A(n596), .B(n2625), .Z(n2624) );
  XOR U2431 ( .A(p_input[821]), .B(n2623), .Z(n2625) );
  XOR U2432 ( .A(n2626), .B(n2627), .Z(n2623) );
  AND U2433 ( .A(n600), .B(n2628), .Z(n2627) );
  XOR U2434 ( .A(n2629), .B(n2630), .Z(n2621) );
  AND U2435 ( .A(n604), .B(n2628), .Z(n2630) );
  XNOR U2436 ( .A(n2629), .B(n2626), .Z(n2628) );
  XOR U2437 ( .A(n2631), .B(n2632), .Z(n2626) );
  AND U2438 ( .A(n607), .B(n2633), .Z(n2632) );
  XOR U2439 ( .A(p_input[837]), .B(n2631), .Z(n2633) );
  XOR U2440 ( .A(n2634), .B(n2635), .Z(n2631) );
  AND U2441 ( .A(n611), .B(n2636), .Z(n2635) );
  XOR U2442 ( .A(n2637), .B(n2638), .Z(n2629) );
  AND U2443 ( .A(n615), .B(n2636), .Z(n2638) );
  XNOR U2444 ( .A(n2637), .B(n2634), .Z(n2636) );
  XOR U2445 ( .A(n2639), .B(n2640), .Z(n2634) );
  AND U2446 ( .A(n618), .B(n2641), .Z(n2640) );
  XOR U2447 ( .A(p_input[853]), .B(n2639), .Z(n2641) );
  XOR U2448 ( .A(n2642), .B(n2643), .Z(n2639) );
  AND U2449 ( .A(n622), .B(n2644), .Z(n2643) );
  XOR U2450 ( .A(n2645), .B(n2646), .Z(n2637) );
  AND U2451 ( .A(n626), .B(n2644), .Z(n2646) );
  XNOR U2452 ( .A(n2645), .B(n2642), .Z(n2644) );
  XOR U2453 ( .A(n2647), .B(n2648), .Z(n2642) );
  AND U2454 ( .A(n629), .B(n2649), .Z(n2648) );
  XOR U2455 ( .A(p_input[869]), .B(n2647), .Z(n2649) );
  XOR U2456 ( .A(n2650), .B(n2651), .Z(n2647) );
  AND U2457 ( .A(n633), .B(n2652), .Z(n2651) );
  XOR U2458 ( .A(n2653), .B(n2654), .Z(n2645) );
  AND U2459 ( .A(n637), .B(n2652), .Z(n2654) );
  XNOR U2460 ( .A(n2653), .B(n2650), .Z(n2652) );
  XOR U2461 ( .A(n2655), .B(n2656), .Z(n2650) );
  AND U2462 ( .A(n640), .B(n2657), .Z(n2656) );
  XOR U2463 ( .A(p_input[885]), .B(n2655), .Z(n2657) );
  XOR U2464 ( .A(n2658), .B(n2659), .Z(n2655) );
  AND U2465 ( .A(n644), .B(n2660), .Z(n2659) );
  XOR U2466 ( .A(n2661), .B(n2662), .Z(n2653) );
  AND U2467 ( .A(n648), .B(n2660), .Z(n2662) );
  XNOR U2468 ( .A(n2661), .B(n2658), .Z(n2660) );
  XOR U2469 ( .A(n2663), .B(n2664), .Z(n2658) );
  AND U2470 ( .A(n651), .B(n2665), .Z(n2664) );
  XOR U2471 ( .A(p_input[901]), .B(n2663), .Z(n2665) );
  XOR U2472 ( .A(n2666), .B(n2667), .Z(n2663) );
  AND U2473 ( .A(n655), .B(n2668), .Z(n2667) );
  XOR U2474 ( .A(n2669), .B(n2670), .Z(n2661) );
  AND U2475 ( .A(n659), .B(n2668), .Z(n2670) );
  XNOR U2476 ( .A(n2669), .B(n2666), .Z(n2668) );
  XOR U2477 ( .A(n2671), .B(n2672), .Z(n2666) );
  AND U2478 ( .A(n662), .B(n2673), .Z(n2672) );
  XOR U2479 ( .A(p_input[917]), .B(n2671), .Z(n2673) );
  XOR U2480 ( .A(n2674), .B(n2675), .Z(n2671) );
  AND U2481 ( .A(n666), .B(n2676), .Z(n2675) );
  XOR U2482 ( .A(n2677), .B(n2678), .Z(n2669) );
  AND U2483 ( .A(n670), .B(n2676), .Z(n2678) );
  XNOR U2484 ( .A(n2677), .B(n2674), .Z(n2676) );
  XOR U2485 ( .A(n2679), .B(n2680), .Z(n2674) );
  AND U2486 ( .A(n673), .B(n2681), .Z(n2680) );
  XOR U2487 ( .A(p_input[933]), .B(n2679), .Z(n2681) );
  XOR U2488 ( .A(n2682), .B(n2683), .Z(n2679) );
  AND U2489 ( .A(n677), .B(n2684), .Z(n2683) );
  XOR U2490 ( .A(n2685), .B(n2686), .Z(n2677) );
  AND U2491 ( .A(n681), .B(n2684), .Z(n2686) );
  XNOR U2492 ( .A(n2685), .B(n2682), .Z(n2684) );
  XOR U2493 ( .A(n2687), .B(n2688), .Z(n2682) );
  AND U2494 ( .A(n684), .B(n2689), .Z(n2688) );
  XOR U2495 ( .A(p_input[949]), .B(n2687), .Z(n2689) );
  XOR U2496 ( .A(n2690), .B(n2691), .Z(n2687) );
  AND U2497 ( .A(n688), .B(n2692), .Z(n2691) );
  XOR U2498 ( .A(n2693), .B(n2694), .Z(n2685) );
  AND U2499 ( .A(n692), .B(n2692), .Z(n2694) );
  XNOR U2500 ( .A(n2693), .B(n2690), .Z(n2692) );
  XOR U2501 ( .A(n2695), .B(n2696), .Z(n2690) );
  AND U2502 ( .A(n695), .B(n2697), .Z(n2696) );
  XOR U2503 ( .A(p_input[965]), .B(n2695), .Z(n2697) );
  XOR U2504 ( .A(n2698), .B(n2699), .Z(n2695) );
  AND U2505 ( .A(n699), .B(n2700), .Z(n2699) );
  XOR U2506 ( .A(n2701), .B(n2702), .Z(n2693) );
  AND U2507 ( .A(n703), .B(n2700), .Z(n2702) );
  XNOR U2508 ( .A(n2701), .B(n2698), .Z(n2700) );
  XOR U2509 ( .A(n2703), .B(n2704), .Z(n2698) );
  AND U2510 ( .A(n706), .B(n2705), .Z(n2704) );
  XOR U2511 ( .A(p_input[981]), .B(n2703), .Z(n2705) );
  XNOR U2512 ( .A(n2706), .B(n2707), .Z(n2703) );
  AND U2513 ( .A(n710), .B(n2708), .Z(n2707) );
  XNOR U2514 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n2709), .Z(n2701) );
  AND U2515 ( .A(n713), .B(n2708), .Z(n2709) );
  XOR U2516 ( .A(n2710), .B(n2706), .Z(n2708) );
  XOR U2517 ( .A(n11), .B(n2711), .Z(o[20]) );
  AND U2518 ( .A(n30), .B(n2712), .Z(n11) );
  XOR U2519 ( .A(n12), .B(n2711), .Z(n2712) );
  XOR U2520 ( .A(n2713), .B(n2714), .Z(n2711) );
  AND U2521 ( .A(n34), .B(n2715), .Z(n2714) );
  XOR U2522 ( .A(p_input[4]), .B(n2713), .Z(n2715) );
  XOR U2523 ( .A(n2716), .B(n2717), .Z(n2713) );
  AND U2524 ( .A(n38), .B(n2718), .Z(n2717) );
  XOR U2525 ( .A(n2719), .B(n2720), .Z(n12) );
  AND U2526 ( .A(n42), .B(n2718), .Z(n2720) );
  XNOR U2527 ( .A(n2721), .B(n2716), .Z(n2718) );
  XOR U2528 ( .A(n2722), .B(n2723), .Z(n2716) );
  AND U2529 ( .A(n46), .B(n2724), .Z(n2723) );
  XOR U2530 ( .A(p_input[20]), .B(n2722), .Z(n2724) );
  XOR U2531 ( .A(n2725), .B(n2726), .Z(n2722) );
  AND U2532 ( .A(n50), .B(n2727), .Z(n2726) );
  IV U2533 ( .A(n2719), .Z(n2721) );
  XNOR U2534 ( .A(n2728), .B(n2729), .Z(n2719) );
  AND U2535 ( .A(n54), .B(n2727), .Z(n2729) );
  XNOR U2536 ( .A(n2728), .B(n2725), .Z(n2727) );
  XOR U2537 ( .A(n2730), .B(n2731), .Z(n2725) );
  AND U2538 ( .A(n57), .B(n2732), .Z(n2731) );
  XOR U2539 ( .A(p_input[36]), .B(n2730), .Z(n2732) );
  XOR U2540 ( .A(n2733), .B(n2734), .Z(n2730) );
  AND U2541 ( .A(n61), .B(n2735), .Z(n2734) );
  XOR U2542 ( .A(n2736), .B(n2737), .Z(n2728) );
  AND U2543 ( .A(n65), .B(n2735), .Z(n2737) );
  XNOR U2544 ( .A(n2736), .B(n2733), .Z(n2735) );
  XOR U2545 ( .A(n2738), .B(n2739), .Z(n2733) );
  AND U2546 ( .A(n68), .B(n2740), .Z(n2739) );
  XOR U2547 ( .A(p_input[52]), .B(n2738), .Z(n2740) );
  XOR U2548 ( .A(n2741), .B(n2742), .Z(n2738) );
  AND U2549 ( .A(n72), .B(n2743), .Z(n2742) );
  XOR U2550 ( .A(n2744), .B(n2745), .Z(n2736) );
  AND U2551 ( .A(n76), .B(n2743), .Z(n2745) );
  XNOR U2552 ( .A(n2744), .B(n2741), .Z(n2743) );
  XOR U2553 ( .A(n2746), .B(n2747), .Z(n2741) );
  AND U2554 ( .A(n79), .B(n2748), .Z(n2747) );
  XOR U2555 ( .A(p_input[68]), .B(n2746), .Z(n2748) );
  XOR U2556 ( .A(n2749), .B(n2750), .Z(n2746) );
  AND U2557 ( .A(n83), .B(n2751), .Z(n2750) );
  XOR U2558 ( .A(n2752), .B(n2753), .Z(n2744) );
  AND U2559 ( .A(n87), .B(n2751), .Z(n2753) );
  XNOR U2560 ( .A(n2752), .B(n2749), .Z(n2751) );
  XOR U2561 ( .A(n2754), .B(n2755), .Z(n2749) );
  AND U2562 ( .A(n90), .B(n2756), .Z(n2755) );
  XOR U2563 ( .A(p_input[84]), .B(n2754), .Z(n2756) );
  XOR U2564 ( .A(n2757), .B(n2758), .Z(n2754) );
  AND U2565 ( .A(n94), .B(n2759), .Z(n2758) );
  XOR U2566 ( .A(n2760), .B(n2761), .Z(n2752) );
  AND U2567 ( .A(n98), .B(n2759), .Z(n2761) );
  XNOR U2568 ( .A(n2760), .B(n2757), .Z(n2759) );
  XOR U2569 ( .A(n2762), .B(n2763), .Z(n2757) );
  AND U2570 ( .A(n101), .B(n2764), .Z(n2763) );
  XOR U2571 ( .A(p_input[100]), .B(n2762), .Z(n2764) );
  XOR U2572 ( .A(n2765), .B(n2766), .Z(n2762) );
  AND U2573 ( .A(n105), .B(n2767), .Z(n2766) );
  XOR U2574 ( .A(n2768), .B(n2769), .Z(n2760) );
  AND U2575 ( .A(n109), .B(n2767), .Z(n2769) );
  XNOR U2576 ( .A(n2768), .B(n2765), .Z(n2767) );
  XOR U2577 ( .A(n2770), .B(n2771), .Z(n2765) );
  AND U2578 ( .A(n112), .B(n2772), .Z(n2771) );
  XOR U2579 ( .A(p_input[116]), .B(n2770), .Z(n2772) );
  XOR U2580 ( .A(n2773), .B(n2774), .Z(n2770) );
  AND U2581 ( .A(n116), .B(n2775), .Z(n2774) );
  XOR U2582 ( .A(n2776), .B(n2777), .Z(n2768) );
  AND U2583 ( .A(n120), .B(n2775), .Z(n2777) );
  XNOR U2584 ( .A(n2776), .B(n2773), .Z(n2775) );
  XOR U2585 ( .A(n2778), .B(n2779), .Z(n2773) );
  AND U2586 ( .A(n123), .B(n2780), .Z(n2779) );
  XOR U2587 ( .A(p_input[132]), .B(n2778), .Z(n2780) );
  XOR U2588 ( .A(n2781), .B(n2782), .Z(n2778) );
  AND U2589 ( .A(n127), .B(n2783), .Z(n2782) );
  XOR U2590 ( .A(n2784), .B(n2785), .Z(n2776) );
  AND U2591 ( .A(n131), .B(n2783), .Z(n2785) );
  XNOR U2592 ( .A(n2784), .B(n2781), .Z(n2783) );
  XOR U2593 ( .A(n2786), .B(n2787), .Z(n2781) );
  AND U2594 ( .A(n134), .B(n2788), .Z(n2787) );
  XOR U2595 ( .A(p_input[148]), .B(n2786), .Z(n2788) );
  XOR U2596 ( .A(n2789), .B(n2790), .Z(n2786) );
  AND U2597 ( .A(n138), .B(n2791), .Z(n2790) );
  XOR U2598 ( .A(n2792), .B(n2793), .Z(n2784) );
  AND U2599 ( .A(n142), .B(n2791), .Z(n2793) );
  XNOR U2600 ( .A(n2792), .B(n2789), .Z(n2791) );
  XOR U2601 ( .A(n2794), .B(n2795), .Z(n2789) );
  AND U2602 ( .A(n145), .B(n2796), .Z(n2795) );
  XOR U2603 ( .A(p_input[164]), .B(n2794), .Z(n2796) );
  XOR U2604 ( .A(n2797), .B(n2798), .Z(n2794) );
  AND U2605 ( .A(n149), .B(n2799), .Z(n2798) );
  XOR U2606 ( .A(n2800), .B(n2801), .Z(n2792) );
  AND U2607 ( .A(n153), .B(n2799), .Z(n2801) );
  XNOR U2608 ( .A(n2800), .B(n2797), .Z(n2799) );
  XOR U2609 ( .A(n2802), .B(n2803), .Z(n2797) );
  AND U2610 ( .A(n156), .B(n2804), .Z(n2803) );
  XOR U2611 ( .A(p_input[180]), .B(n2802), .Z(n2804) );
  XOR U2612 ( .A(n2805), .B(n2806), .Z(n2802) );
  AND U2613 ( .A(n160), .B(n2807), .Z(n2806) );
  XOR U2614 ( .A(n2808), .B(n2809), .Z(n2800) );
  AND U2615 ( .A(n164), .B(n2807), .Z(n2809) );
  XNOR U2616 ( .A(n2808), .B(n2805), .Z(n2807) );
  XOR U2617 ( .A(n2810), .B(n2811), .Z(n2805) );
  AND U2618 ( .A(n167), .B(n2812), .Z(n2811) );
  XOR U2619 ( .A(p_input[196]), .B(n2810), .Z(n2812) );
  XOR U2620 ( .A(n2813), .B(n2814), .Z(n2810) );
  AND U2621 ( .A(n171), .B(n2815), .Z(n2814) );
  XOR U2622 ( .A(n2816), .B(n2817), .Z(n2808) );
  AND U2623 ( .A(n175), .B(n2815), .Z(n2817) );
  XNOR U2624 ( .A(n2816), .B(n2813), .Z(n2815) );
  XOR U2625 ( .A(n2818), .B(n2819), .Z(n2813) );
  AND U2626 ( .A(n178), .B(n2820), .Z(n2819) );
  XOR U2627 ( .A(p_input[212]), .B(n2818), .Z(n2820) );
  XOR U2628 ( .A(n2821), .B(n2822), .Z(n2818) );
  AND U2629 ( .A(n182), .B(n2823), .Z(n2822) );
  XOR U2630 ( .A(n2824), .B(n2825), .Z(n2816) );
  AND U2631 ( .A(n186), .B(n2823), .Z(n2825) );
  XNOR U2632 ( .A(n2824), .B(n2821), .Z(n2823) );
  XOR U2633 ( .A(n2826), .B(n2827), .Z(n2821) );
  AND U2634 ( .A(n189), .B(n2828), .Z(n2827) );
  XOR U2635 ( .A(p_input[228]), .B(n2826), .Z(n2828) );
  XOR U2636 ( .A(n2829), .B(n2830), .Z(n2826) );
  AND U2637 ( .A(n193), .B(n2831), .Z(n2830) );
  XOR U2638 ( .A(n2832), .B(n2833), .Z(n2824) );
  AND U2639 ( .A(n197), .B(n2831), .Z(n2833) );
  XNOR U2640 ( .A(n2832), .B(n2829), .Z(n2831) );
  XOR U2641 ( .A(n2834), .B(n2835), .Z(n2829) );
  AND U2642 ( .A(n200), .B(n2836), .Z(n2835) );
  XOR U2643 ( .A(p_input[244]), .B(n2834), .Z(n2836) );
  XOR U2644 ( .A(n2837), .B(n2838), .Z(n2834) );
  AND U2645 ( .A(n204), .B(n2839), .Z(n2838) );
  XOR U2646 ( .A(n2840), .B(n2841), .Z(n2832) );
  AND U2647 ( .A(n208), .B(n2839), .Z(n2841) );
  XNOR U2648 ( .A(n2840), .B(n2837), .Z(n2839) );
  XOR U2649 ( .A(n2842), .B(n2843), .Z(n2837) );
  AND U2650 ( .A(n211), .B(n2844), .Z(n2843) );
  XOR U2651 ( .A(p_input[260]), .B(n2842), .Z(n2844) );
  XOR U2652 ( .A(n2845), .B(n2846), .Z(n2842) );
  AND U2653 ( .A(n215), .B(n2847), .Z(n2846) );
  XOR U2654 ( .A(n2848), .B(n2849), .Z(n2840) );
  AND U2655 ( .A(n219), .B(n2847), .Z(n2849) );
  XNOR U2656 ( .A(n2848), .B(n2845), .Z(n2847) );
  XOR U2657 ( .A(n2850), .B(n2851), .Z(n2845) );
  AND U2658 ( .A(n222), .B(n2852), .Z(n2851) );
  XOR U2659 ( .A(p_input[276]), .B(n2850), .Z(n2852) );
  XOR U2660 ( .A(n2853), .B(n2854), .Z(n2850) );
  AND U2661 ( .A(n226), .B(n2855), .Z(n2854) );
  XOR U2662 ( .A(n2856), .B(n2857), .Z(n2848) );
  AND U2663 ( .A(n230), .B(n2855), .Z(n2857) );
  XNOR U2664 ( .A(n2856), .B(n2853), .Z(n2855) );
  XOR U2665 ( .A(n2858), .B(n2859), .Z(n2853) );
  AND U2666 ( .A(n233), .B(n2860), .Z(n2859) );
  XOR U2667 ( .A(p_input[292]), .B(n2858), .Z(n2860) );
  XOR U2668 ( .A(n2861), .B(n2862), .Z(n2858) );
  AND U2669 ( .A(n237), .B(n2863), .Z(n2862) );
  XOR U2670 ( .A(n2864), .B(n2865), .Z(n2856) );
  AND U2671 ( .A(n241), .B(n2863), .Z(n2865) );
  XNOR U2672 ( .A(n2864), .B(n2861), .Z(n2863) );
  XOR U2673 ( .A(n2866), .B(n2867), .Z(n2861) );
  AND U2674 ( .A(n244), .B(n2868), .Z(n2867) );
  XOR U2675 ( .A(p_input[308]), .B(n2866), .Z(n2868) );
  XOR U2676 ( .A(n2869), .B(n2870), .Z(n2866) );
  AND U2677 ( .A(n248), .B(n2871), .Z(n2870) );
  XOR U2678 ( .A(n2872), .B(n2873), .Z(n2864) );
  AND U2679 ( .A(n252), .B(n2871), .Z(n2873) );
  XNOR U2680 ( .A(n2872), .B(n2869), .Z(n2871) );
  XOR U2681 ( .A(n2874), .B(n2875), .Z(n2869) );
  AND U2682 ( .A(n255), .B(n2876), .Z(n2875) );
  XOR U2683 ( .A(p_input[324]), .B(n2874), .Z(n2876) );
  XOR U2684 ( .A(n2877), .B(n2878), .Z(n2874) );
  AND U2685 ( .A(n259), .B(n2879), .Z(n2878) );
  XOR U2686 ( .A(n2880), .B(n2881), .Z(n2872) );
  AND U2687 ( .A(n263), .B(n2879), .Z(n2881) );
  XNOR U2688 ( .A(n2880), .B(n2877), .Z(n2879) );
  XOR U2689 ( .A(n2882), .B(n2883), .Z(n2877) );
  AND U2690 ( .A(n266), .B(n2884), .Z(n2883) );
  XOR U2691 ( .A(p_input[340]), .B(n2882), .Z(n2884) );
  XOR U2692 ( .A(n2885), .B(n2886), .Z(n2882) );
  AND U2693 ( .A(n270), .B(n2887), .Z(n2886) );
  XOR U2694 ( .A(n2888), .B(n2889), .Z(n2880) );
  AND U2695 ( .A(n274), .B(n2887), .Z(n2889) );
  XNOR U2696 ( .A(n2888), .B(n2885), .Z(n2887) );
  XOR U2697 ( .A(n2890), .B(n2891), .Z(n2885) );
  AND U2698 ( .A(n277), .B(n2892), .Z(n2891) );
  XOR U2699 ( .A(p_input[356]), .B(n2890), .Z(n2892) );
  XOR U2700 ( .A(n2893), .B(n2894), .Z(n2890) );
  AND U2701 ( .A(n281), .B(n2895), .Z(n2894) );
  XOR U2702 ( .A(n2896), .B(n2897), .Z(n2888) );
  AND U2703 ( .A(n285), .B(n2895), .Z(n2897) );
  XNOR U2704 ( .A(n2896), .B(n2893), .Z(n2895) );
  XOR U2705 ( .A(n2898), .B(n2899), .Z(n2893) );
  AND U2706 ( .A(n288), .B(n2900), .Z(n2899) );
  XOR U2707 ( .A(p_input[372]), .B(n2898), .Z(n2900) );
  XOR U2708 ( .A(n2901), .B(n2902), .Z(n2898) );
  AND U2709 ( .A(n292), .B(n2903), .Z(n2902) );
  XOR U2710 ( .A(n2904), .B(n2905), .Z(n2896) );
  AND U2711 ( .A(n296), .B(n2903), .Z(n2905) );
  XNOR U2712 ( .A(n2904), .B(n2901), .Z(n2903) );
  XOR U2713 ( .A(n2906), .B(n2907), .Z(n2901) );
  AND U2714 ( .A(n299), .B(n2908), .Z(n2907) );
  XOR U2715 ( .A(p_input[388]), .B(n2906), .Z(n2908) );
  XOR U2716 ( .A(n2909), .B(n2910), .Z(n2906) );
  AND U2717 ( .A(n303), .B(n2911), .Z(n2910) );
  XOR U2718 ( .A(n2912), .B(n2913), .Z(n2904) );
  AND U2719 ( .A(n307), .B(n2911), .Z(n2913) );
  XNOR U2720 ( .A(n2912), .B(n2909), .Z(n2911) );
  XOR U2721 ( .A(n2914), .B(n2915), .Z(n2909) );
  AND U2722 ( .A(n310), .B(n2916), .Z(n2915) );
  XOR U2723 ( .A(p_input[404]), .B(n2914), .Z(n2916) );
  XOR U2724 ( .A(n2917), .B(n2918), .Z(n2914) );
  AND U2725 ( .A(n314), .B(n2919), .Z(n2918) );
  XOR U2726 ( .A(n2920), .B(n2921), .Z(n2912) );
  AND U2727 ( .A(n318), .B(n2919), .Z(n2921) );
  XNOR U2728 ( .A(n2920), .B(n2917), .Z(n2919) );
  XOR U2729 ( .A(n2922), .B(n2923), .Z(n2917) );
  AND U2730 ( .A(n321), .B(n2924), .Z(n2923) );
  XOR U2731 ( .A(p_input[420]), .B(n2922), .Z(n2924) );
  XOR U2732 ( .A(n2925), .B(n2926), .Z(n2922) );
  AND U2733 ( .A(n325), .B(n2927), .Z(n2926) );
  XOR U2734 ( .A(n2928), .B(n2929), .Z(n2920) );
  AND U2735 ( .A(n329), .B(n2927), .Z(n2929) );
  XNOR U2736 ( .A(n2928), .B(n2925), .Z(n2927) );
  XOR U2737 ( .A(n2930), .B(n2931), .Z(n2925) );
  AND U2738 ( .A(n332), .B(n2932), .Z(n2931) );
  XOR U2739 ( .A(p_input[436]), .B(n2930), .Z(n2932) );
  XOR U2740 ( .A(n2933), .B(n2934), .Z(n2930) );
  AND U2741 ( .A(n336), .B(n2935), .Z(n2934) );
  XOR U2742 ( .A(n2936), .B(n2937), .Z(n2928) );
  AND U2743 ( .A(n340), .B(n2935), .Z(n2937) );
  XNOR U2744 ( .A(n2936), .B(n2933), .Z(n2935) );
  XOR U2745 ( .A(n2938), .B(n2939), .Z(n2933) );
  AND U2746 ( .A(n343), .B(n2940), .Z(n2939) );
  XOR U2747 ( .A(p_input[452]), .B(n2938), .Z(n2940) );
  XOR U2748 ( .A(n2941), .B(n2942), .Z(n2938) );
  AND U2749 ( .A(n347), .B(n2943), .Z(n2942) );
  XOR U2750 ( .A(n2944), .B(n2945), .Z(n2936) );
  AND U2751 ( .A(n351), .B(n2943), .Z(n2945) );
  XNOR U2752 ( .A(n2944), .B(n2941), .Z(n2943) );
  XOR U2753 ( .A(n2946), .B(n2947), .Z(n2941) );
  AND U2754 ( .A(n354), .B(n2948), .Z(n2947) );
  XOR U2755 ( .A(p_input[468]), .B(n2946), .Z(n2948) );
  XOR U2756 ( .A(n2949), .B(n2950), .Z(n2946) );
  AND U2757 ( .A(n358), .B(n2951), .Z(n2950) );
  XOR U2758 ( .A(n2952), .B(n2953), .Z(n2944) );
  AND U2759 ( .A(n362), .B(n2951), .Z(n2953) );
  XNOR U2760 ( .A(n2952), .B(n2949), .Z(n2951) );
  XOR U2761 ( .A(n2954), .B(n2955), .Z(n2949) );
  AND U2762 ( .A(n365), .B(n2956), .Z(n2955) );
  XOR U2763 ( .A(p_input[484]), .B(n2954), .Z(n2956) );
  XOR U2764 ( .A(n2957), .B(n2958), .Z(n2954) );
  AND U2765 ( .A(n369), .B(n2959), .Z(n2958) );
  XOR U2766 ( .A(n2960), .B(n2961), .Z(n2952) );
  AND U2767 ( .A(n373), .B(n2959), .Z(n2961) );
  XNOR U2768 ( .A(n2960), .B(n2957), .Z(n2959) );
  XOR U2769 ( .A(n2962), .B(n2963), .Z(n2957) );
  AND U2770 ( .A(n376), .B(n2964), .Z(n2963) );
  XOR U2771 ( .A(p_input[500]), .B(n2962), .Z(n2964) );
  XOR U2772 ( .A(n2965), .B(n2966), .Z(n2962) );
  AND U2773 ( .A(n380), .B(n2967), .Z(n2966) );
  XOR U2774 ( .A(n2968), .B(n2969), .Z(n2960) );
  AND U2775 ( .A(n384), .B(n2967), .Z(n2969) );
  XNOR U2776 ( .A(n2968), .B(n2965), .Z(n2967) );
  XOR U2777 ( .A(n2970), .B(n2971), .Z(n2965) );
  AND U2778 ( .A(n387), .B(n2972), .Z(n2971) );
  XOR U2779 ( .A(p_input[516]), .B(n2970), .Z(n2972) );
  XOR U2780 ( .A(n2973), .B(n2974), .Z(n2970) );
  AND U2781 ( .A(n391), .B(n2975), .Z(n2974) );
  XOR U2782 ( .A(n2976), .B(n2977), .Z(n2968) );
  AND U2783 ( .A(n395), .B(n2975), .Z(n2977) );
  XNOR U2784 ( .A(n2976), .B(n2973), .Z(n2975) );
  XOR U2785 ( .A(n2978), .B(n2979), .Z(n2973) );
  AND U2786 ( .A(n398), .B(n2980), .Z(n2979) );
  XOR U2787 ( .A(p_input[532]), .B(n2978), .Z(n2980) );
  XOR U2788 ( .A(n2981), .B(n2982), .Z(n2978) );
  AND U2789 ( .A(n402), .B(n2983), .Z(n2982) );
  XOR U2790 ( .A(n2984), .B(n2985), .Z(n2976) );
  AND U2791 ( .A(n406), .B(n2983), .Z(n2985) );
  XNOR U2792 ( .A(n2984), .B(n2981), .Z(n2983) );
  XOR U2793 ( .A(n2986), .B(n2987), .Z(n2981) );
  AND U2794 ( .A(n409), .B(n2988), .Z(n2987) );
  XOR U2795 ( .A(p_input[548]), .B(n2986), .Z(n2988) );
  XOR U2796 ( .A(n2989), .B(n2990), .Z(n2986) );
  AND U2797 ( .A(n413), .B(n2991), .Z(n2990) );
  XOR U2798 ( .A(n2992), .B(n2993), .Z(n2984) );
  AND U2799 ( .A(n417), .B(n2991), .Z(n2993) );
  XNOR U2800 ( .A(n2992), .B(n2989), .Z(n2991) );
  XOR U2801 ( .A(n2994), .B(n2995), .Z(n2989) );
  AND U2802 ( .A(n420), .B(n2996), .Z(n2995) );
  XOR U2803 ( .A(p_input[564]), .B(n2994), .Z(n2996) );
  XOR U2804 ( .A(n2997), .B(n2998), .Z(n2994) );
  AND U2805 ( .A(n424), .B(n2999), .Z(n2998) );
  XOR U2806 ( .A(n3000), .B(n3001), .Z(n2992) );
  AND U2807 ( .A(n428), .B(n2999), .Z(n3001) );
  XNOR U2808 ( .A(n3000), .B(n2997), .Z(n2999) );
  XOR U2809 ( .A(n3002), .B(n3003), .Z(n2997) );
  AND U2810 ( .A(n431), .B(n3004), .Z(n3003) );
  XOR U2811 ( .A(p_input[580]), .B(n3002), .Z(n3004) );
  XOR U2812 ( .A(n3005), .B(n3006), .Z(n3002) );
  AND U2813 ( .A(n435), .B(n3007), .Z(n3006) );
  XOR U2814 ( .A(n3008), .B(n3009), .Z(n3000) );
  AND U2815 ( .A(n439), .B(n3007), .Z(n3009) );
  XNOR U2816 ( .A(n3008), .B(n3005), .Z(n3007) );
  XOR U2817 ( .A(n3010), .B(n3011), .Z(n3005) );
  AND U2818 ( .A(n442), .B(n3012), .Z(n3011) );
  XOR U2819 ( .A(p_input[596]), .B(n3010), .Z(n3012) );
  XOR U2820 ( .A(n3013), .B(n3014), .Z(n3010) );
  AND U2821 ( .A(n446), .B(n3015), .Z(n3014) );
  XOR U2822 ( .A(n3016), .B(n3017), .Z(n3008) );
  AND U2823 ( .A(n450), .B(n3015), .Z(n3017) );
  XNOR U2824 ( .A(n3016), .B(n3013), .Z(n3015) );
  XOR U2825 ( .A(n3018), .B(n3019), .Z(n3013) );
  AND U2826 ( .A(n453), .B(n3020), .Z(n3019) );
  XOR U2827 ( .A(p_input[612]), .B(n3018), .Z(n3020) );
  XOR U2828 ( .A(n3021), .B(n3022), .Z(n3018) );
  AND U2829 ( .A(n457), .B(n3023), .Z(n3022) );
  XOR U2830 ( .A(n3024), .B(n3025), .Z(n3016) );
  AND U2831 ( .A(n461), .B(n3023), .Z(n3025) );
  XNOR U2832 ( .A(n3024), .B(n3021), .Z(n3023) );
  XOR U2833 ( .A(n3026), .B(n3027), .Z(n3021) );
  AND U2834 ( .A(n464), .B(n3028), .Z(n3027) );
  XOR U2835 ( .A(p_input[628]), .B(n3026), .Z(n3028) );
  XOR U2836 ( .A(n3029), .B(n3030), .Z(n3026) );
  AND U2837 ( .A(n468), .B(n3031), .Z(n3030) );
  XOR U2838 ( .A(n3032), .B(n3033), .Z(n3024) );
  AND U2839 ( .A(n472), .B(n3031), .Z(n3033) );
  XNOR U2840 ( .A(n3032), .B(n3029), .Z(n3031) );
  XOR U2841 ( .A(n3034), .B(n3035), .Z(n3029) );
  AND U2842 ( .A(n475), .B(n3036), .Z(n3035) );
  XOR U2843 ( .A(p_input[644]), .B(n3034), .Z(n3036) );
  XOR U2844 ( .A(n3037), .B(n3038), .Z(n3034) );
  AND U2845 ( .A(n479), .B(n3039), .Z(n3038) );
  XOR U2846 ( .A(n3040), .B(n3041), .Z(n3032) );
  AND U2847 ( .A(n483), .B(n3039), .Z(n3041) );
  XNOR U2848 ( .A(n3040), .B(n3037), .Z(n3039) );
  XOR U2849 ( .A(n3042), .B(n3043), .Z(n3037) );
  AND U2850 ( .A(n486), .B(n3044), .Z(n3043) );
  XOR U2851 ( .A(p_input[660]), .B(n3042), .Z(n3044) );
  XOR U2852 ( .A(n3045), .B(n3046), .Z(n3042) );
  AND U2853 ( .A(n490), .B(n3047), .Z(n3046) );
  XOR U2854 ( .A(n3048), .B(n3049), .Z(n3040) );
  AND U2855 ( .A(n494), .B(n3047), .Z(n3049) );
  XNOR U2856 ( .A(n3048), .B(n3045), .Z(n3047) );
  XOR U2857 ( .A(n3050), .B(n3051), .Z(n3045) );
  AND U2858 ( .A(n497), .B(n3052), .Z(n3051) );
  XOR U2859 ( .A(p_input[676]), .B(n3050), .Z(n3052) );
  XOR U2860 ( .A(n3053), .B(n3054), .Z(n3050) );
  AND U2861 ( .A(n501), .B(n3055), .Z(n3054) );
  XOR U2862 ( .A(n3056), .B(n3057), .Z(n3048) );
  AND U2863 ( .A(n505), .B(n3055), .Z(n3057) );
  XNOR U2864 ( .A(n3056), .B(n3053), .Z(n3055) );
  XOR U2865 ( .A(n3058), .B(n3059), .Z(n3053) );
  AND U2866 ( .A(n508), .B(n3060), .Z(n3059) );
  XOR U2867 ( .A(p_input[692]), .B(n3058), .Z(n3060) );
  XOR U2868 ( .A(n3061), .B(n3062), .Z(n3058) );
  AND U2869 ( .A(n512), .B(n3063), .Z(n3062) );
  XOR U2870 ( .A(n3064), .B(n3065), .Z(n3056) );
  AND U2871 ( .A(n516), .B(n3063), .Z(n3065) );
  XNOR U2872 ( .A(n3064), .B(n3061), .Z(n3063) );
  XOR U2873 ( .A(n3066), .B(n3067), .Z(n3061) );
  AND U2874 ( .A(n519), .B(n3068), .Z(n3067) );
  XOR U2875 ( .A(p_input[708]), .B(n3066), .Z(n3068) );
  XOR U2876 ( .A(n3069), .B(n3070), .Z(n3066) );
  AND U2877 ( .A(n523), .B(n3071), .Z(n3070) );
  XOR U2878 ( .A(n3072), .B(n3073), .Z(n3064) );
  AND U2879 ( .A(n527), .B(n3071), .Z(n3073) );
  XNOR U2880 ( .A(n3072), .B(n3069), .Z(n3071) );
  XOR U2881 ( .A(n3074), .B(n3075), .Z(n3069) );
  AND U2882 ( .A(n530), .B(n3076), .Z(n3075) );
  XOR U2883 ( .A(p_input[724]), .B(n3074), .Z(n3076) );
  XOR U2884 ( .A(n3077), .B(n3078), .Z(n3074) );
  AND U2885 ( .A(n534), .B(n3079), .Z(n3078) );
  XOR U2886 ( .A(n3080), .B(n3081), .Z(n3072) );
  AND U2887 ( .A(n538), .B(n3079), .Z(n3081) );
  XNOR U2888 ( .A(n3080), .B(n3077), .Z(n3079) );
  XOR U2889 ( .A(n3082), .B(n3083), .Z(n3077) );
  AND U2890 ( .A(n541), .B(n3084), .Z(n3083) );
  XOR U2891 ( .A(p_input[740]), .B(n3082), .Z(n3084) );
  XOR U2892 ( .A(n3085), .B(n3086), .Z(n3082) );
  AND U2893 ( .A(n545), .B(n3087), .Z(n3086) );
  XOR U2894 ( .A(n3088), .B(n3089), .Z(n3080) );
  AND U2895 ( .A(n549), .B(n3087), .Z(n3089) );
  XNOR U2896 ( .A(n3088), .B(n3085), .Z(n3087) );
  XOR U2897 ( .A(n3090), .B(n3091), .Z(n3085) );
  AND U2898 ( .A(n552), .B(n3092), .Z(n3091) );
  XOR U2899 ( .A(p_input[756]), .B(n3090), .Z(n3092) );
  XOR U2900 ( .A(n3093), .B(n3094), .Z(n3090) );
  AND U2901 ( .A(n556), .B(n3095), .Z(n3094) );
  XOR U2902 ( .A(n3096), .B(n3097), .Z(n3088) );
  AND U2903 ( .A(n560), .B(n3095), .Z(n3097) );
  XNOR U2904 ( .A(n3096), .B(n3093), .Z(n3095) );
  XOR U2905 ( .A(n3098), .B(n3099), .Z(n3093) );
  AND U2906 ( .A(n563), .B(n3100), .Z(n3099) );
  XOR U2907 ( .A(p_input[772]), .B(n3098), .Z(n3100) );
  XOR U2908 ( .A(n3101), .B(n3102), .Z(n3098) );
  AND U2909 ( .A(n567), .B(n3103), .Z(n3102) );
  XOR U2910 ( .A(n3104), .B(n3105), .Z(n3096) );
  AND U2911 ( .A(n571), .B(n3103), .Z(n3105) );
  XNOR U2912 ( .A(n3104), .B(n3101), .Z(n3103) );
  XOR U2913 ( .A(n3106), .B(n3107), .Z(n3101) );
  AND U2914 ( .A(n574), .B(n3108), .Z(n3107) );
  XOR U2915 ( .A(p_input[788]), .B(n3106), .Z(n3108) );
  XOR U2916 ( .A(n3109), .B(n3110), .Z(n3106) );
  AND U2917 ( .A(n578), .B(n3111), .Z(n3110) );
  XOR U2918 ( .A(n3112), .B(n3113), .Z(n3104) );
  AND U2919 ( .A(n582), .B(n3111), .Z(n3113) );
  XNOR U2920 ( .A(n3112), .B(n3109), .Z(n3111) );
  XOR U2921 ( .A(n3114), .B(n3115), .Z(n3109) );
  AND U2922 ( .A(n585), .B(n3116), .Z(n3115) );
  XOR U2923 ( .A(p_input[804]), .B(n3114), .Z(n3116) );
  XOR U2924 ( .A(n3117), .B(n3118), .Z(n3114) );
  AND U2925 ( .A(n589), .B(n3119), .Z(n3118) );
  XOR U2926 ( .A(n3120), .B(n3121), .Z(n3112) );
  AND U2927 ( .A(n593), .B(n3119), .Z(n3121) );
  XNOR U2928 ( .A(n3120), .B(n3117), .Z(n3119) );
  XOR U2929 ( .A(n3122), .B(n3123), .Z(n3117) );
  AND U2930 ( .A(n596), .B(n3124), .Z(n3123) );
  XOR U2931 ( .A(p_input[820]), .B(n3122), .Z(n3124) );
  XOR U2932 ( .A(n3125), .B(n3126), .Z(n3122) );
  AND U2933 ( .A(n600), .B(n3127), .Z(n3126) );
  XOR U2934 ( .A(n3128), .B(n3129), .Z(n3120) );
  AND U2935 ( .A(n604), .B(n3127), .Z(n3129) );
  XNOR U2936 ( .A(n3128), .B(n3125), .Z(n3127) );
  XOR U2937 ( .A(n3130), .B(n3131), .Z(n3125) );
  AND U2938 ( .A(n607), .B(n3132), .Z(n3131) );
  XOR U2939 ( .A(p_input[836]), .B(n3130), .Z(n3132) );
  XOR U2940 ( .A(n3133), .B(n3134), .Z(n3130) );
  AND U2941 ( .A(n611), .B(n3135), .Z(n3134) );
  XOR U2942 ( .A(n3136), .B(n3137), .Z(n3128) );
  AND U2943 ( .A(n615), .B(n3135), .Z(n3137) );
  XNOR U2944 ( .A(n3136), .B(n3133), .Z(n3135) );
  XOR U2945 ( .A(n3138), .B(n3139), .Z(n3133) );
  AND U2946 ( .A(n618), .B(n3140), .Z(n3139) );
  XOR U2947 ( .A(p_input[852]), .B(n3138), .Z(n3140) );
  XOR U2948 ( .A(n3141), .B(n3142), .Z(n3138) );
  AND U2949 ( .A(n622), .B(n3143), .Z(n3142) );
  XOR U2950 ( .A(n3144), .B(n3145), .Z(n3136) );
  AND U2951 ( .A(n626), .B(n3143), .Z(n3145) );
  XNOR U2952 ( .A(n3144), .B(n3141), .Z(n3143) );
  XOR U2953 ( .A(n3146), .B(n3147), .Z(n3141) );
  AND U2954 ( .A(n629), .B(n3148), .Z(n3147) );
  XOR U2955 ( .A(p_input[868]), .B(n3146), .Z(n3148) );
  XOR U2956 ( .A(n3149), .B(n3150), .Z(n3146) );
  AND U2957 ( .A(n633), .B(n3151), .Z(n3150) );
  XOR U2958 ( .A(n3152), .B(n3153), .Z(n3144) );
  AND U2959 ( .A(n637), .B(n3151), .Z(n3153) );
  XNOR U2960 ( .A(n3152), .B(n3149), .Z(n3151) );
  XOR U2961 ( .A(n3154), .B(n3155), .Z(n3149) );
  AND U2962 ( .A(n640), .B(n3156), .Z(n3155) );
  XOR U2963 ( .A(p_input[884]), .B(n3154), .Z(n3156) );
  XOR U2964 ( .A(n3157), .B(n3158), .Z(n3154) );
  AND U2965 ( .A(n644), .B(n3159), .Z(n3158) );
  XOR U2966 ( .A(n3160), .B(n3161), .Z(n3152) );
  AND U2967 ( .A(n648), .B(n3159), .Z(n3161) );
  XNOR U2968 ( .A(n3160), .B(n3157), .Z(n3159) );
  XOR U2969 ( .A(n3162), .B(n3163), .Z(n3157) );
  AND U2970 ( .A(n651), .B(n3164), .Z(n3163) );
  XOR U2971 ( .A(p_input[900]), .B(n3162), .Z(n3164) );
  XOR U2972 ( .A(n3165), .B(n3166), .Z(n3162) );
  AND U2973 ( .A(n655), .B(n3167), .Z(n3166) );
  XOR U2974 ( .A(n3168), .B(n3169), .Z(n3160) );
  AND U2975 ( .A(n659), .B(n3167), .Z(n3169) );
  XNOR U2976 ( .A(n3168), .B(n3165), .Z(n3167) );
  XOR U2977 ( .A(n3170), .B(n3171), .Z(n3165) );
  AND U2978 ( .A(n662), .B(n3172), .Z(n3171) );
  XOR U2979 ( .A(p_input[916]), .B(n3170), .Z(n3172) );
  XOR U2980 ( .A(n3173), .B(n3174), .Z(n3170) );
  AND U2981 ( .A(n666), .B(n3175), .Z(n3174) );
  XOR U2982 ( .A(n3176), .B(n3177), .Z(n3168) );
  AND U2983 ( .A(n670), .B(n3175), .Z(n3177) );
  XNOR U2984 ( .A(n3176), .B(n3173), .Z(n3175) );
  XOR U2985 ( .A(n3178), .B(n3179), .Z(n3173) );
  AND U2986 ( .A(n673), .B(n3180), .Z(n3179) );
  XOR U2987 ( .A(p_input[932]), .B(n3178), .Z(n3180) );
  XOR U2988 ( .A(n3181), .B(n3182), .Z(n3178) );
  AND U2989 ( .A(n677), .B(n3183), .Z(n3182) );
  XOR U2990 ( .A(n3184), .B(n3185), .Z(n3176) );
  AND U2991 ( .A(n681), .B(n3183), .Z(n3185) );
  XNOR U2992 ( .A(n3184), .B(n3181), .Z(n3183) );
  XOR U2993 ( .A(n3186), .B(n3187), .Z(n3181) );
  AND U2994 ( .A(n684), .B(n3188), .Z(n3187) );
  XOR U2995 ( .A(p_input[948]), .B(n3186), .Z(n3188) );
  XOR U2996 ( .A(n3189), .B(n3190), .Z(n3186) );
  AND U2997 ( .A(n688), .B(n3191), .Z(n3190) );
  XOR U2998 ( .A(n3192), .B(n3193), .Z(n3184) );
  AND U2999 ( .A(n692), .B(n3191), .Z(n3193) );
  XNOR U3000 ( .A(n3192), .B(n3189), .Z(n3191) );
  XOR U3001 ( .A(n3194), .B(n3195), .Z(n3189) );
  AND U3002 ( .A(n695), .B(n3196), .Z(n3195) );
  XOR U3003 ( .A(p_input[964]), .B(n3194), .Z(n3196) );
  XOR U3004 ( .A(n3197), .B(n3198), .Z(n3194) );
  AND U3005 ( .A(n699), .B(n3199), .Z(n3198) );
  XOR U3006 ( .A(n3200), .B(n3201), .Z(n3192) );
  AND U3007 ( .A(n703), .B(n3199), .Z(n3201) );
  XNOR U3008 ( .A(n3200), .B(n3197), .Z(n3199) );
  XOR U3009 ( .A(n3202), .B(n3203), .Z(n3197) );
  AND U3010 ( .A(n706), .B(n3204), .Z(n3203) );
  XOR U3011 ( .A(p_input[980]), .B(n3202), .Z(n3204) );
  XNOR U3012 ( .A(n3205), .B(n3206), .Z(n3202) );
  AND U3013 ( .A(n710), .B(n3207), .Z(n3206) );
  XNOR U3014 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n3208), .Z(n3200) );
  AND U3015 ( .A(n713), .B(n3207), .Z(n3208) );
  XOR U3016 ( .A(n3209), .B(n3205), .Z(n3207) );
  IV U3017 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .Z(n3205) );
  IV U3018 ( .A(\knn_comb_/min_val_out[0][4] ), .Z(n3209) );
  XOR U3019 ( .A(n3210), .B(n3211), .Z(o[1]) );
  XOR U3020 ( .A(n13), .B(n3212), .Z(o[19]) );
  AND U3021 ( .A(n30), .B(n3213), .Z(n13) );
  XOR U3022 ( .A(n14), .B(n3212), .Z(n3213) );
  XOR U3023 ( .A(n3214), .B(n3215), .Z(n3212) );
  AND U3024 ( .A(n34), .B(n3216), .Z(n3215) );
  XOR U3025 ( .A(p_input[3]), .B(n3214), .Z(n3216) );
  XOR U3026 ( .A(n3217), .B(n3218), .Z(n3214) );
  AND U3027 ( .A(n38), .B(n3219), .Z(n3218) );
  XOR U3028 ( .A(n3220), .B(n3221), .Z(n14) );
  AND U3029 ( .A(n42), .B(n3219), .Z(n3221) );
  XNOR U3030 ( .A(n3222), .B(n3217), .Z(n3219) );
  XOR U3031 ( .A(n3223), .B(n3224), .Z(n3217) );
  AND U3032 ( .A(n46), .B(n3225), .Z(n3224) );
  XOR U3033 ( .A(p_input[19]), .B(n3223), .Z(n3225) );
  XOR U3034 ( .A(n3226), .B(n3227), .Z(n3223) );
  AND U3035 ( .A(n50), .B(n3228), .Z(n3227) );
  IV U3036 ( .A(n3220), .Z(n3222) );
  XNOR U3037 ( .A(n3229), .B(n3230), .Z(n3220) );
  AND U3038 ( .A(n54), .B(n3228), .Z(n3230) );
  XNOR U3039 ( .A(n3229), .B(n3226), .Z(n3228) );
  XOR U3040 ( .A(n3231), .B(n3232), .Z(n3226) );
  AND U3041 ( .A(n57), .B(n3233), .Z(n3232) );
  XOR U3042 ( .A(p_input[35]), .B(n3231), .Z(n3233) );
  XOR U3043 ( .A(n3234), .B(n3235), .Z(n3231) );
  AND U3044 ( .A(n61), .B(n3236), .Z(n3235) );
  XOR U3045 ( .A(n3237), .B(n3238), .Z(n3229) );
  AND U3046 ( .A(n65), .B(n3236), .Z(n3238) );
  XNOR U3047 ( .A(n3237), .B(n3234), .Z(n3236) );
  XOR U3048 ( .A(n3239), .B(n3240), .Z(n3234) );
  AND U3049 ( .A(n68), .B(n3241), .Z(n3240) );
  XOR U3050 ( .A(p_input[51]), .B(n3239), .Z(n3241) );
  XOR U3051 ( .A(n3242), .B(n3243), .Z(n3239) );
  AND U3052 ( .A(n72), .B(n3244), .Z(n3243) );
  XOR U3053 ( .A(n3245), .B(n3246), .Z(n3237) );
  AND U3054 ( .A(n76), .B(n3244), .Z(n3246) );
  XNOR U3055 ( .A(n3245), .B(n3242), .Z(n3244) );
  XOR U3056 ( .A(n3247), .B(n3248), .Z(n3242) );
  AND U3057 ( .A(n79), .B(n3249), .Z(n3248) );
  XOR U3058 ( .A(p_input[67]), .B(n3247), .Z(n3249) );
  XOR U3059 ( .A(n3250), .B(n3251), .Z(n3247) );
  AND U3060 ( .A(n83), .B(n3252), .Z(n3251) );
  XOR U3061 ( .A(n3253), .B(n3254), .Z(n3245) );
  AND U3062 ( .A(n87), .B(n3252), .Z(n3254) );
  XNOR U3063 ( .A(n3253), .B(n3250), .Z(n3252) );
  XOR U3064 ( .A(n3255), .B(n3256), .Z(n3250) );
  AND U3065 ( .A(n90), .B(n3257), .Z(n3256) );
  XOR U3066 ( .A(p_input[83]), .B(n3255), .Z(n3257) );
  XOR U3067 ( .A(n3258), .B(n3259), .Z(n3255) );
  AND U3068 ( .A(n94), .B(n3260), .Z(n3259) );
  XOR U3069 ( .A(n3261), .B(n3262), .Z(n3253) );
  AND U3070 ( .A(n98), .B(n3260), .Z(n3262) );
  XNOR U3071 ( .A(n3261), .B(n3258), .Z(n3260) );
  XOR U3072 ( .A(n3263), .B(n3264), .Z(n3258) );
  AND U3073 ( .A(n101), .B(n3265), .Z(n3264) );
  XOR U3074 ( .A(p_input[99]), .B(n3263), .Z(n3265) );
  XOR U3075 ( .A(n3266), .B(n3267), .Z(n3263) );
  AND U3076 ( .A(n105), .B(n3268), .Z(n3267) );
  XOR U3077 ( .A(n3269), .B(n3270), .Z(n3261) );
  AND U3078 ( .A(n109), .B(n3268), .Z(n3270) );
  XNOR U3079 ( .A(n3269), .B(n3266), .Z(n3268) );
  XOR U3080 ( .A(n3271), .B(n3272), .Z(n3266) );
  AND U3081 ( .A(n112), .B(n3273), .Z(n3272) );
  XOR U3082 ( .A(p_input[115]), .B(n3271), .Z(n3273) );
  XOR U3083 ( .A(n3274), .B(n3275), .Z(n3271) );
  AND U3084 ( .A(n116), .B(n3276), .Z(n3275) );
  XOR U3085 ( .A(n3277), .B(n3278), .Z(n3269) );
  AND U3086 ( .A(n120), .B(n3276), .Z(n3278) );
  XNOR U3087 ( .A(n3277), .B(n3274), .Z(n3276) );
  XOR U3088 ( .A(n3279), .B(n3280), .Z(n3274) );
  AND U3089 ( .A(n123), .B(n3281), .Z(n3280) );
  XOR U3090 ( .A(p_input[131]), .B(n3279), .Z(n3281) );
  XOR U3091 ( .A(n3282), .B(n3283), .Z(n3279) );
  AND U3092 ( .A(n127), .B(n3284), .Z(n3283) );
  XOR U3093 ( .A(n3285), .B(n3286), .Z(n3277) );
  AND U3094 ( .A(n131), .B(n3284), .Z(n3286) );
  XNOR U3095 ( .A(n3285), .B(n3282), .Z(n3284) );
  XOR U3096 ( .A(n3287), .B(n3288), .Z(n3282) );
  AND U3097 ( .A(n134), .B(n3289), .Z(n3288) );
  XOR U3098 ( .A(p_input[147]), .B(n3287), .Z(n3289) );
  XOR U3099 ( .A(n3290), .B(n3291), .Z(n3287) );
  AND U3100 ( .A(n138), .B(n3292), .Z(n3291) );
  XOR U3101 ( .A(n3293), .B(n3294), .Z(n3285) );
  AND U3102 ( .A(n142), .B(n3292), .Z(n3294) );
  XNOR U3103 ( .A(n3293), .B(n3290), .Z(n3292) );
  XOR U3104 ( .A(n3295), .B(n3296), .Z(n3290) );
  AND U3105 ( .A(n145), .B(n3297), .Z(n3296) );
  XOR U3106 ( .A(p_input[163]), .B(n3295), .Z(n3297) );
  XOR U3107 ( .A(n3298), .B(n3299), .Z(n3295) );
  AND U3108 ( .A(n149), .B(n3300), .Z(n3299) );
  XOR U3109 ( .A(n3301), .B(n3302), .Z(n3293) );
  AND U3110 ( .A(n153), .B(n3300), .Z(n3302) );
  XNOR U3111 ( .A(n3301), .B(n3298), .Z(n3300) );
  XOR U3112 ( .A(n3303), .B(n3304), .Z(n3298) );
  AND U3113 ( .A(n156), .B(n3305), .Z(n3304) );
  XOR U3114 ( .A(p_input[179]), .B(n3303), .Z(n3305) );
  XOR U3115 ( .A(n3306), .B(n3307), .Z(n3303) );
  AND U3116 ( .A(n160), .B(n3308), .Z(n3307) );
  XOR U3117 ( .A(n3309), .B(n3310), .Z(n3301) );
  AND U3118 ( .A(n164), .B(n3308), .Z(n3310) );
  XNOR U3119 ( .A(n3309), .B(n3306), .Z(n3308) );
  XOR U3120 ( .A(n3311), .B(n3312), .Z(n3306) );
  AND U3121 ( .A(n167), .B(n3313), .Z(n3312) );
  XOR U3122 ( .A(p_input[195]), .B(n3311), .Z(n3313) );
  XOR U3123 ( .A(n3314), .B(n3315), .Z(n3311) );
  AND U3124 ( .A(n171), .B(n3316), .Z(n3315) );
  XOR U3125 ( .A(n3317), .B(n3318), .Z(n3309) );
  AND U3126 ( .A(n175), .B(n3316), .Z(n3318) );
  XNOR U3127 ( .A(n3317), .B(n3314), .Z(n3316) );
  XOR U3128 ( .A(n3319), .B(n3320), .Z(n3314) );
  AND U3129 ( .A(n178), .B(n3321), .Z(n3320) );
  XOR U3130 ( .A(p_input[211]), .B(n3319), .Z(n3321) );
  XOR U3131 ( .A(n3322), .B(n3323), .Z(n3319) );
  AND U3132 ( .A(n182), .B(n3324), .Z(n3323) );
  XOR U3133 ( .A(n3325), .B(n3326), .Z(n3317) );
  AND U3134 ( .A(n186), .B(n3324), .Z(n3326) );
  XNOR U3135 ( .A(n3325), .B(n3322), .Z(n3324) );
  XOR U3136 ( .A(n3327), .B(n3328), .Z(n3322) );
  AND U3137 ( .A(n189), .B(n3329), .Z(n3328) );
  XOR U3138 ( .A(p_input[227]), .B(n3327), .Z(n3329) );
  XOR U3139 ( .A(n3330), .B(n3331), .Z(n3327) );
  AND U3140 ( .A(n193), .B(n3332), .Z(n3331) );
  XOR U3141 ( .A(n3333), .B(n3334), .Z(n3325) );
  AND U3142 ( .A(n197), .B(n3332), .Z(n3334) );
  XNOR U3143 ( .A(n3333), .B(n3330), .Z(n3332) );
  XOR U3144 ( .A(n3335), .B(n3336), .Z(n3330) );
  AND U3145 ( .A(n200), .B(n3337), .Z(n3336) );
  XOR U3146 ( .A(p_input[243]), .B(n3335), .Z(n3337) );
  XOR U3147 ( .A(n3338), .B(n3339), .Z(n3335) );
  AND U3148 ( .A(n204), .B(n3340), .Z(n3339) );
  XOR U3149 ( .A(n3341), .B(n3342), .Z(n3333) );
  AND U3150 ( .A(n208), .B(n3340), .Z(n3342) );
  XNOR U3151 ( .A(n3341), .B(n3338), .Z(n3340) );
  XOR U3152 ( .A(n3343), .B(n3344), .Z(n3338) );
  AND U3153 ( .A(n211), .B(n3345), .Z(n3344) );
  XOR U3154 ( .A(p_input[259]), .B(n3343), .Z(n3345) );
  XOR U3155 ( .A(n3346), .B(n3347), .Z(n3343) );
  AND U3156 ( .A(n215), .B(n3348), .Z(n3347) );
  XOR U3157 ( .A(n3349), .B(n3350), .Z(n3341) );
  AND U3158 ( .A(n219), .B(n3348), .Z(n3350) );
  XNOR U3159 ( .A(n3349), .B(n3346), .Z(n3348) );
  XOR U3160 ( .A(n3351), .B(n3352), .Z(n3346) );
  AND U3161 ( .A(n222), .B(n3353), .Z(n3352) );
  XOR U3162 ( .A(p_input[275]), .B(n3351), .Z(n3353) );
  XOR U3163 ( .A(n3354), .B(n3355), .Z(n3351) );
  AND U3164 ( .A(n226), .B(n3356), .Z(n3355) );
  XOR U3165 ( .A(n3357), .B(n3358), .Z(n3349) );
  AND U3166 ( .A(n230), .B(n3356), .Z(n3358) );
  XNOR U3167 ( .A(n3357), .B(n3354), .Z(n3356) );
  XOR U3168 ( .A(n3359), .B(n3360), .Z(n3354) );
  AND U3169 ( .A(n233), .B(n3361), .Z(n3360) );
  XOR U3170 ( .A(p_input[291]), .B(n3359), .Z(n3361) );
  XOR U3171 ( .A(n3362), .B(n3363), .Z(n3359) );
  AND U3172 ( .A(n237), .B(n3364), .Z(n3363) );
  XOR U3173 ( .A(n3365), .B(n3366), .Z(n3357) );
  AND U3174 ( .A(n241), .B(n3364), .Z(n3366) );
  XNOR U3175 ( .A(n3365), .B(n3362), .Z(n3364) );
  XOR U3176 ( .A(n3367), .B(n3368), .Z(n3362) );
  AND U3177 ( .A(n244), .B(n3369), .Z(n3368) );
  XOR U3178 ( .A(p_input[307]), .B(n3367), .Z(n3369) );
  XOR U3179 ( .A(n3370), .B(n3371), .Z(n3367) );
  AND U3180 ( .A(n248), .B(n3372), .Z(n3371) );
  XOR U3181 ( .A(n3373), .B(n3374), .Z(n3365) );
  AND U3182 ( .A(n252), .B(n3372), .Z(n3374) );
  XNOR U3183 ( .A(n3373), .B(n3370), .Z(n3372) );
  XOR U3184 ( .A(n3375), .B(n3376), .Z(n3370) );
  AND U3185 ( .A(n255), .B(n3377), .Z(n3376) );
  XOR U3186 ( .A(p_input[323]), .B(n3375), .Z(n3377) );
  XOR U3187 ( .A(n3378), .B(n3379), .Z(n3375) );
  AND U3188 ( .A(n259), .B(n3380), .Z(n3379) );
  XOR U3189 ( .A(n3381), .B(n3382), .Z(n3373) );
  AND U3190 ( .A(n263), .B(n3380), .Z(n3382) );
  XNOR U3191 ( .A(n3381), .B(n3378), .Z(n3380) );
  XOR U3192 ( .A(n3383), .B(n3384), .Z(n3378) );
  AND U3193 ( .A(n266), .B(n3385), .Z(n3384) );
  XOR U3194 ( .A(p_input[339]), .B(n3383), .Z(n3385) );
  XOR U3195 ( .A(n3386), .B(n3387), .Z(n3383) );
  AND U3196 ( .A(n270), .B(n3388), .Z(n3387) );
  XOR U3197 ( .A(n3389), .B(n3390), .Z(n3381) );
  AND U3198 ( .A(n274), .B(n3388), .Z(n3390) );
  XNOR U3199 ( .A(n3389), .B(n3386), .Z(n3388) );
  XOR U3200 ( .A(n3391), .B(n3392), .Z(n3386) );
  AND U3201 ( .A(n277), .B(n3393), .Z(n3392) );
  XOR U3202 ( .A(p_input[355]), .B(n3391), .Z(n3393) );
  XOR U3203 ( .A(n3394), .B(n3395), .Z(n3391) );
  AND U3204 ( .A(n281), .B(n3396), .Z(n3395) );
  XOR U3205 ( .A(n3397), .B(n3398), .Z(n3389) );
  AND U3206 ( .A(n285), .B(n3396), .Z(n3398) );
  XNOR U3207 ( .A(n3397), .B(n3394), .Z(n3396) );
  XOR U3208 ( .A(n3399), .B(n3400), .Z(n3394) );
  AND U3209 ( .A(n288), .B(n3401), .Z(n3400) );
  XOR U3210 ( .A(p_input[371]), .B(n3399), .Z(n3401) );
  XOR U3211 ( .A(n3402), .B(n3403), .Z(n3399) );
  AND U3212 ( .A(n292), .B(n3404), .Z(n3403) );
  XOR U3213 ( .A(n3405), .B(n3406), .Z(n3397) );
  AND U3214 ( .A(n296), .B(n3404), .Z(n3406) );
  XNOR U3215 ( .A(n3405), .B(n3402), .Z(n3404) );
  XOR U3216 ( .A(n3407), .B(n3408), .Z(n3402) );
  AND U3217 ( .A(n299), .B(n3409), .Z(n3408) );
  XOR U3218 ( .A(p_input[387]), .B(n3407), .Z(n3409) );
  XOR U3219 ( .A(n3410), .B(n3411), .Z(n3407) );
  AND U3220 ( .A(n303), .B(n3412), .Z(n3411) );
  XOR U3221 ( .A(n3413), .B(n3414), .Z(n3405) );
  AND U3222 ( .A(n307), .B(n3412), .Z(n3414) );
  XNOR U3223 ( .A(n3413), .B(n3410), .Z(n3412) );
  XOR U3224 ( .A(n3415), .B(n3416), .Z(n3410) );
  AND U3225 ( .A(n310), .B(n3417), .Z(n3416) );
  XOR U3226 ( .A(p_input[403]), .B(n3415), .Z(n3417) );
  XOR U3227 ( .A(n3418), .B(n3419), .Z(n3415) );
  AND U3228 ( .A(n314), .B(n3420), .Z(n3419) );
  XOR U3229 ( .A(n3421), .B(n3422), .Z(n3413) );
  AND U3230 ( .A(n318), .B(n3420), .Z(n3422) );
  XNOR U3231 ( .A(n3421), .B(n3418), .Z(n3420) );
  XOR U3232 ( .A(n3423), .B(n3424), .Z(n3418) );
  AND U3233 ( .A(n321), .B(n3425), .Z(n3424) );
  XOR U3234 ( .A(p_input[419]), .B(n3423), .Z(n3425) );
  XOR U3235 ( .A(n3426), .B(n3427), .Z(n3423) );
  AND U3236 ( .A(n325), .B(n3428), .Z(n3427) );
  XOR U3237 ( .A(n3429), .B(n3430), .Z(n3421) );
  AND U3238 ( .A(n329), .B(n3428), .Z(n3430) );
  XNOR U3239 ( .A(n3429), .B(n3426), .Z(n3428) );
  XOR U3240 ( .A(n3431), .B(n3432), .Z(n3426) );
  AND U3241 ( .A(n332), .B(n3433), .Z(n3432) );
  XOR U3242 ( .A(p_input[435]), .B(n3431), .Z(n3433) );
  XOR U3243 ( .A(n3434), .B(n3435), .Z(n3431) );
  AND U3244 ( .A(n336), .B(n3436), .Z(n3435) );
  XOR U3245 ( .A(n3437), .B(n3438), .Z(n3429) );
  AND U3246 ( .A(n340), .B(n3436), .Z(n3438) );
  XNOR U3247 ( .A(n3437), .B(n3434), .Z(n3436) );
  XOR U3248 ( .A(n3439), .B(n3440), .Z(n3434) );
  AND U3249 ( .A(n343), .B(n3441), .Z(n3440) );
  XOR U3250 ( .A(p_input[451]), .B(n3439), .Z(n3441) );
  XOR U3251 ( .A(n3442), .B(n3443), .Z(n3439) );
  AND U3252 ( .A(n347), .B(n3444), .Z(n3443) );
  XOR U3253 ( .A(n3445), .B(n3446), .Z(n3437) );
  AND U3254 ( .A(n351), .B(n3444), .Z(n3446) );
  XNOR U3255 ( .A(n3445), .B(n3442), .Z(n3444) );
  XOR U3256 ( .A(n3447), .B(n3448), .Z(n3442) );
  AND U3257 ( .A(n354), .B(n3449), .Z(n3448) );
  XOR U3258 ( .A(p_input[467]), .B(n3447), .Z(n3449) );
  XOR U3259 ( .A(n3450), .B(n3451), .Z(n3447) );
  AND U3260 ( .A(n358), .B(n3452), .Z(n3451) );
  XOR U3261 ( .A(n3453), .B(n3454), .Z(n3445) );
  AND U3262 ( .A(n362), .B(n3452), .Z(n3454) );
  XNOR U3263 ( .A(n3453), .B(n3450), .Z(n3452) );
  XOR U3264 ( .A(n3455), .B(n3456), .Z(n3450) );
  AND U3265 ( .A(n365), .B(n3457), .Z(n3456) );
  XOR U3266 ( .A(p_input[483]), .B(n3455), .Z(n3457) );
  XOR U3267 ( .A(n3458), .B(n3459), .Z(n3455) );
  AND U3268 ( .A(n369), .B(n3460), .Z(n3459) );
  XOR U3269 ( .A(n3461), .B(n3462), .Z(n3453) );
  AND U3270 ( .A(n373), .B(n3460), .Z(n3462) );
  XNOR U3271 ( .A(n3461), .B(n3458), .Z(n3460) );
  XOR U3272 ( .A(n3463), .B(n3464), .Z(n3458) );
  AND U3273 ( .A(n376), .B(n3465), .Z(n3464) );
  XOR U3274 ( .A(p_input[499]), .B(n3463), .Z(n3465) );
  XOR U3275 ( .A(n3466), .B(n3467), .Z(n3463) );
  AND U3276 ( .A(n380), .B(n3468), .Z(n3467) );
  XOR U3277 ( .A(n3469), .B(n3470), .Z(n3461) );
  AND U3278 ( .A(n384), .B(n3468), .Z(n3470) );
  XNOR U3279 ( .A(n3469), .B(n3466), .Z(n3468) );
  XOR U3280 ( .A(n3471), .B(n3472), .Z(n3466) );
  AND U3281 ( .A(n387), .B(n3473), .Z(n3472) );
  XOR U3282 ( .A(p_input[515]), .B(n3471), .Z(n3473) );
  XOR U3283 ( .A(n3474), .B(n3475), .Z(n3471) );
  AND U3284 ( .A(n391), .B(n3476), .Z(n3475) );
  XOR U3285 ( .A(n3477), .B(n3478), .Z(n3469) );
  AND U3286 ( .A(n395), .B(n3476), .Z(n3478) );
  XNOR U3287 ( .A(n3477), .B(n3474), .Z(n3476) );
  XOR U3288 ( .A(n3479), .B(n3480), .Z(n3474) );
  AND U3289 ( .A(n398), .B(n3481), .Z(n3480) );
  XOR U3290 ( .A(p_input[531]), .B(n3479), .Z(n3481) );
  XOR U3291 ( .A(n3482), .B(n3483), .Z(n3479) );
  AND U3292 ( .A(n402), .B(n3484), .Z(n3483) );
  XOR U3293 ( .A(n3485), .B(n3486), .Z(n3477) );
  AND U3294 ( .A(n406), .B(n3484), .Z(n3486) );
  XNOR U3295 ( .A(n3485), .B(n3482), .Z(n3484) );
  XOR U3296 ( .A(n3487), .B(n3488), .Z(n3482) );
  AND U3297 ( .A(n409), .B(n3489), .Z(n3488) );
  XOR U3298 ( .A(p_input[547]), .B(n3487), .Z(n3489) );
  XOR U3299 ( .A(n3490), .B(n3491), .Z(n3487) );
  AND U3300 ( .A(n413), .B(n3492), .Z(n3491) );
  XOR U3301 ( .A(n3493), .B(n3494), .Z(n3485) );
  AND U3302 ( .A(n417), .B(n3492), .Z(n3494) );
  XNOR U3303 ( .A(n3493), .B(n3490), .Z(n3492) );
  XOR U3304 ( .A(n3495), .B(n3496), .Z(n3490) );
  AND U3305 ( .A(n420), .B(n3497), .Z(n3496) );
  XOR U3306 ( .A(p_input[563]), .B(n3495), .Z(n3497) );
  XOR U3307 ( .A(n3498), .B(n3499), .Z(n3495) );
  AND U3308 ( .A(n424), .B(n3500), .Z(n3499) );
  XOR U3309 ( .A(n3501), .B(n3502), .Z(n3493) );
  AND U3310 ( .A(n428), .B(n3500), .Z(n3502) );
  XNOR U3311 ( .A(n3501), .B(n3498), .Z(n3500) );
  XOR U3312 ( .A(n3503), .B(n3504), .Z(n3498) );
  AND U3313 ( .A(n431), .B(n3505), .Z(n3504) );
  XOR U3314 ( .A(p_input[579]), .B(n3503), .Z(n3505) );
  XOR U3315 ( .A(n3506), .B(n3507), .Z(n3503) );
  AND U3316 ( .A(n435), .B(n3508), .Z(n3507) );
  XOR U3317 ( .A(n3509), .B(n3510), .Z(n3501) );
  AND U3318 ( .A(n439), .B(n3508), .Z(n3510) );
  XNOR U3319 ( .A(n3509), .B(n3506), .Z(n3508) );
  XOR U3320 ( .A(n3511), .B(n3512), .Z(n3506) );
  AND U3321 ( .A(n442), .B(n3513), .Z(n3512) );
  XOR U3322 ( .A(p_input[595]), .B(n3511), .Z(n3513) );
  XOR U3323 ( .A(n3514), .B(n3515), .Z(n3511) );
  AND U3324 ( .A(n446), .B(n3516), .Z(n3515) );
  XOR U3325 ( .A(n3517), .B(n3518), .Z(n3509) );
  AND U3326 ( .A(n450), .B(n3516), .Z(n3518) );
  XNOR U3327 ( .A(n3517), .B(n3514), .Z(n3516) );
  XOR U3328 ( .A(n3519), .B(n3520), .Z(n3514) );
  AND U3329 ( .A(n453), .B(n3521), .Z(n3520) );
  XOR U3330 ( .A(p_input[611]), .B(n3519), .Z(n3521) );
  XOR U3331 ( .A(n3522), .B(n3523), .Z(n3519) );
  AND U3332 ( .A(n457), .B(n3524), .Z(n3523) );
  XOR U3333 ( .A(n3525), .B(n3526), .Z(n3517) );
  AND U3334 ( .A(n461), .B(n3524), .Z(n3526) );
  XNOR U3335 ( .A(n3525), .B(n3522), .Z(n3524) );
  XOR U3336 ( .A(n3527), .B(n3528), .Z(n3522) );
  AND U3337 ( .A(n464), .B(n3529), .Z(n3528) );
  XOR U3338 ( .A(p_input[627]), .B(n3527), .Z(n3529) );
  XOR U3339 ( .A(n3530), .B(n3531), .Z(n3527) );
  AND U3340 ( .A(n468), .B(n3532), .Z(n3531) );
  XOR U3341 ( .A(n3533), .B(n3534), .Z(n3525) );
  AND U3342 ( .A(n472), .B(n3532), .Z(n3534) );
  XNOR U3343 ( .A(n3533), .B(n3530), .Z(n3532) );
  XOR U3344 ( .A(n3535), .B(n3536), .Z(n3530) );
  AND U3345 ( .A(n475), .B(n3537), .Z(n3536) );
  XOR U3346 ( .A(p_input[643]), .B(n3535), .Z(n3537) );
  XOR U3347 ( .A(n3538), .B(n3539), .Z(n3535) );
  AND U3348 ( .A(n479), .B(n3540), .Z(n3539) );
  XOR U3349 ( .A(n3541), .B(n3542), .Z(n3533) );
  AND U3350 ( .A(n483), .B(n3540), .Z(n3542) );
  XNOR U3351 ( .A(n3541), .B(n3538), .Z(n3540) );
  XOR U3352 ( .A(n3543), .B(n3544), .Z(n3538) );
  AND U3353 ( .A(n486), .B(n3545), .Z(n3544) );
  XOR U3354 ( .A(p_input[659]), .B(n3543), .Z(n3545) );
  XOR U3355 ( .A(n3546), .B(n3547), .Z(n3543) );
  AND U3356 ( .A(n490), .B(n3548), .Z(n3547) );
  XOR U3357 ( .A(n3549), .B(n3550), .Z(n3541) );
  AND U3358 ( .A(n494), .B(n3548), .Z(n3550) );
  XNOR U3359 ( .A(n3549), .B(n3546), .Z(n3548) );
  XOR U3360 ( .A(n3551), .B(n3552), .Z(n3546) );
  AND U3361 ( .A(n497), .B(n3553), .Z(n3552) );
  XOR U3362 ( .A(p_input[675]), .B(n3551), .Z(n3553) );
  XOR U3363 ( .A(n3554), .B(n3555), .Z(n3551) );
  AND U3364 ( .A(n501), .B(n3556), .Z(n3555) );
  XOR U3365 ( .A(n3557), .B(n3558), .Z(n3549) );
  AND U3366 ( .A(n505), .B(n3556), .Z(n3558) );
  XNOR U3367 ( .A(n3557), .B(n3554), .Z(n3556) );
  XOR U3368 ( .A(n3559), .B(n3560), .Z(n3554) );
  AND U3369 ( .A(n508), .B(n3561), .Z(n3560) );
  XOR U3370 ( .A(p_input[691]), .B(n3559), .Z(n3561) );
  XOR U3371 ( .A(n3562), .B(n3563), .Z(n3559) );
  AND U3372 ( .A(n512), .B(n3564), .Z(n3563) );
  XOR U3373 ( .A(n3565), .B(n3566), .Z(n3557) );
  AND U3374 ( .A(n516), .B(n3564), .Z(n3566) );
  XNOR U3375 ( .A(n3565), .B(n3562), .Z(n3564) );
  XOR U3376 ( .A(n3567), .B(n3568), .Z(n3562) );
  AND U3377 ( .A(n519), .B(n3569), .Z(n3568) );
  XOR U3378 ( .A(p_input[707]), .B(n3567), .Z(n3569) );
  XOR U3379 ( .A(n3570), .B(n3571), .Z(n3567) );
  AND U3380 ( .A(n523), .B(n3572), .Z(n3571) );
  XOR U3381 ( .A(n3573), .B(n3574), .Z(n3565) );
  AND U3382 ( .A(n527), .B(n3572), .Z(n3574) );
  XNOR U3383 ( .A(n3573), .B(n3570), .Z(n3572) );
  XOR U3384 ( .A(n3575), .B(n3576), .Z(n3570) );
  AND U3385 ( .A(n530), .B(n3577), .Z(n3576) );
  XOR U3386 ( .A(p_input[723]), .B(n3575), .Z(n3577) );
  XOR U3387 ( .A(n3578), .B(n3579), .Z(n3575) );
  AND U3388 ( .A(n534), .B(n3580), .Z(n3579) );
  XOR U3389 ( .A(n3581), .B(n3582), .Z(n3573) );
  AND U3390 ( .A(n538), .B(n3580), .Z(n3582) );
  XNOR U3391 ( .A(n3581), .B(n3578), .Z(n3580) );
  XOR U3392 ( .A(n3583), .B(n3584), .Z(n3578) );
  AND U3393 ( .A(n541), .B(n3585), .Z(n3584) );
  XOR U3394 ( .A(p_input[739]), .B(n3583), .Z(n3585) );
  XOR U3395 ( .A(n3586), .B(n3587), .Z(n3583) );
  AND U3396 ( .A(n545), .B(n3588), .Z(n3587) );
  XOR U3397 ( .A(n3589), .B(n3590), .Z(n3581) );
  AND U3398 ( .A(n549), .B(n3588), .Z(n3590) );
  XNOR U3399 ( .A(n3589), .B(n3586), .Z(n3588) );
  XOR U3400 ( .A(n3591), .B(n3592), .Z(n3586) );
  AND U3401 ( .A(n552), .B(n3593), .Z(n3592) );
  XOR U3402 ( .A(p_input[755]), .B(n3591), .Z(n3593) );
  XOR U3403 ( .A(n3594), .B(n3595), .Z(n3591) );
  AND U3404 ( .A(n556), .B(n3596), .Z(n3595) );
  XOR U3405 ( .A(n3597), .B(n3598), .Z(n3589) );
  AND U3406 ( .A(n560), .B(n3596), .Z(n3598) );
  XNOR U3407 ( .A(n3597), .B(n3594), .Z(n3596) );
  XOR U3408 ( .A(n3599), .B(n3600), .Z(n3594) );
  AND U3409 ( .A(n563), .B(n3601), .Z(n3600) );
  XOR U3410 ( .A(p_input[771]), .B(n3599), .Z(n3601) );
  XOR U3411 ( .A(n3602), .B(n3603), .Z(n3599) );
  AND U3412 ( .A(n567), .B(n3604), .Z(n3603) );
  XOR U3413 ( .A(n3605), .B(n3606), .Z(n3597) );
  AND U3414 ( .A(n571), .B(n3604), .Z(n3606) );
  XNOR U3415 ( .A(n3605), .B(n3602), .Z(n3604) );
  XOR U3416 ( .A(n3607), .B(n3608), .Z(n3602) );
  AND U3417 ( .A(n574), .B(n3609), .Z(n3608) );
  XOR U3418 ( .A(p_input[787]), .B(n3607), .Z(n3609) );
  XOR U3419 ( .A(n3610), .B(n3611), .Z(n3607) );
  AND U3420 ( .A(n578), .B(n3612), .Z(n3611) );
  XOR U3421 ( .A(n3613), .B(n3614), .Z(n3605) );
  AND U3422 ( .A(n582), .B(n3612), .Z(n3614) );
  XNOR U3423 ( .A(n3613), .B(n3610), .Z(n3612) );
  XOR U3424 ( .A(n3615), .B(n3616), .Z(n3610) );
  AND U3425 ( .A(n585), .B(n3617), .Z(n3616) );
  XOR U3426 ( .A(p_input[803]), .B(n3615), .Z(n3617) );
  XOR U3427 ( .A(n3618), .B(n3619), .Z(n3615) );
  AND U3428 ( .A(n589), .B(n3620), .Z(n3619) );
  XOR U3429 ( .A(n3621), .B(n3622), .Z(n3613) );
  AND U3430 ( .A(n593), .B(n3620), .Z(n3622) );
  XNOR U3431 ( .A(n3621), .B(n3618), .Z(n3620) );
  XOR U3432 ( .A(n3623), .B(n3624), .Z(n3618) );
  AND U3433 ( .A(n596), .B(n3625), .Z(n3624) );
  XOR U3434 ( .A(p_input[819]), .B(n3623), .Z(n3625) );
  XOR U3435 ( .A(n3626), .B(n3627), .Z(n3623) );
  AND U3436 ( .A(n600), .B(n3628), .Z(n3627) );
  XOR U3437 ( .A(n3629), .B(n3630), .Z(n3621) );
  AND U3438 ( .A(n604), .B(n3628), .Z(n3630) );
  XNOR U3439 ( .A(n3629), .B(n3626), .Z(n3628) );
  XOR U3440 ( .A(n3631), .B(n3632), .Z(n3626) );
  AND U3441 ( .A(n607), .B(n3633), .Z(n3632) );
  XOR U3442 ( .A(p_input[835]), .B(n3631), .Z(n3633) );
  XOR U3443 ( .A(n3634), .B(n3635), .Z(n3631) );
  AND U3444 ( .A(n611), .B(n3636), .Z(n3635) );
  XOR U3445 ( .A(n3637), .B(n3638), .Z(n3629) );
  AND U3446 ( .A(n615), .B(n3636), .Z(n3638) );
  XNOR U3447 ( .A(n3637), .B(n3634), .Z(n3636) );
  XOR U3448 ( .A(n3639), .B(n3640), .Z(n3634) );
  AND U3449 ( .A(n618), .B(n3641), .Z(n3640) );
  XOR U3450 ( .A(p_input[851]), .B(n3639), .Z(n3641) );
  XOR U3451 ( .A(n3642), .B(n3643), .Z(n3639) );
  AND U3452 ( .A(n622), .B(n3644), .Z(n3643) );
  XOR U3453 ( .A(n3645), .B(n3646), .Z(n3637) );
  AND U3454 ( .A(n626), .B(n3644), .Z(n3646) );
  XNOR U3455 ( .A(n3645), .B(n3642), .Z(n3644) );
  XOR U3456 ( .A(n3647), .B(n3648), .Z(n3642) );
  AND U3457 ( .A(n629), .B(n3649), .Z(n3648) );
  XOR U3458 ( .A(p_input[867]), .B(n3647), .Z(n3649) );
  XOR U3459 ( .A(n3650), .B(n3651), .Z(n3647) );
  AND U3460 ( .A(n633), .B(n3652), .Z(n3651) );
  XOR U3461 ( .A(n3653), .B(n3654), .Z(n3645) );
  AND U3462 ( .A(n637), .B(n3652), .Z(n3654) );
  XNOR U3463 ( .A(n3653), .B(n3650), .Z(n3652) );
  XOR U3464 ( .A(n3655), .B(n3656), .Z(n3650) );
  AND U3465 ( .A(n640), .B(n3657), .Z(n3656) );
  XOR U3466 ( .A(p_input[883]), .B(n3655), .Z(n3657) );
  XOR U3467 ( .A(n3658), .B(n3659), .Z(n3655) );
  AND U3468 ( .A(n644), .B(n3660), .Z(n3659) );
  XOR U3469 ( .A(n3661), .B(n3662), .Z(n3653) );
  AND U3470 ( .A(n648), .B(n3660), .Z(n3662) );
  XNOR U3471 ( .A(n3661), .B(n3658), .Z(n3660) );
  XOR U3472 ( .A(n3663), .B(n3664), .Z(n3658) );
  AND U3473 ( .A(n651), .B(n3665), .Z(n3664) );
  XOR U3474 ( .A(p_input[899]), .B(n3663), .Z(n3665) );
  XOR U3475 ( .A(n3666), .B(n3667), .Z(n3663) );
  AND U3476 ( .A(n655), .B(n3668), .Z(n3667) );
  XOR U3477 ( .A(n3669), .B(n3670), .Z(n3661) );
  AND U3478 ( .A(n659), .B(n3668), .Z(n3670) );
  XNOR U3479 ( .A(n3669), .B(n3666), .Z(n3668) );
  XOR U3480 ( .A(n3671), .B(n3672), .Z(n3666) );
  AND U3481 ( .A(n662), .B(n3673), .Z(n3672) );
  XOR U3482 ( .A(p_input[915]), .B(n3671), .Z(n3673) );
  XOR U3483 ( .A(n3674), .B(n3675), .Z(n3671) );
  AND U3484 ( .A(n666), .B(n3676), .Z(n3675) );
  XOR U3485 ( .A(n3677), .B(n3678), .Z(n3669) );
  AND U3486 ( .A(n670), .B(n3676), .Z(n3678) );
  XNOR U3487 ( .A(n3677), .B(n3674), .Z(n3676) );
  XOR U3488 ( .A(n3679), .B(n3680), .Z(n3674) );
  AND U3489 ( .A(n673), .B(n3681), .Z(n3680) );
  XOR U3490 ( .A(p_input[931]), .B(n3679), .Z(n3681) );
  XOR U3491 ( .A(n3682), .B(n3683), .Z(n3679) );
  AND U3492 ( .A(n677), .B(n3684), .Z(n3683) );
  XOR U3493 ( .A(n3685), .B(n3686), .Z(n3677) );
  AND U3494 ( .A(n681), .B(n3684), .Z(n3686) );
  XNOR U3495 ( .A(n3685), .B(n3682), .Z(n3684) );
  XOR U3496 ( .A(n3687), .B(n3688), .Z(n3682) );
  AND U3497 ( .A(n684), .B(n3689), .Z(n3688) );
  XOR U3498 ( .A(p_input[947]), .B(n3687), .Z(n3689) );
  XOR U3499 ( .A(n3690), .B(n3691), .Z(n3687) );
  AND U3500 ( .A(n688), .B(n3692), .Z(n3691) );
  XOR U3501 ( .A(n3693), .B(n3694), .Z(n3685) );
  AND U3502 ( .A(n692), .B(n3692), .Z(n3694) );
  XNOR U3503 ( .A(n3693), .B(n3690), .Z(n3692) );
  XOR U3504 ( .A(n3695), .B(n3696), .Z(n3690) );
  AND U3505 ( .A(n695), .B(n3697), .Z(n3696) );
  XOR U3506 ( .A(p_input[963]), .B(n3695), .Z(n3697) );
  XOR U3507 ( .A(n3698), .B(n3699), .Z(n3695) );
  AND U3508 ( .A(n699), .B(n3700), .Z(n3699) );
  XOR U3509 ( .A(n3701), .B(n3702), .Z(n3693) );
  AND U3510 ( .A(n703), .B(n3700), .Z(n3702) );
  XNOR U3511 ( .A(n3701), .B(n3698), .Z(n3700) );
  XOR U3512 ( .A(n3703), .B(n3704), .Z(n3698) );
  AND U3513 ( .A(n706), .B(n3705), .Z(n3704) );
  XOR U3514 ( .A(p_input[979]), .B(n3703), .Z(n3705) );
  XNOR U3515 ( .A(n3706), .B(n3707), .Z(n3703) );
  AND U3516 ( .A(n710), .B(n3708), .Z(n3707) );
  XNOR U3517 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n3709), .Z(n3701) );
  AND U3518 ( .A(n713), .B(n3708), .Z(n3709) );
  XOR U3519 ( .A(n3710), .B(n3706), .Z(n3708) );
  IV U3520 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .Z(n3706) );
  XOR U3521 ( .A(n19), .B(n3711), .Z(o[18]) );
  AND U3522 ( .A(n30), .B(n3712), .Z(n19) );
  XOR U3523 ( .A(n20), .B(n3711), .Z(n3712) );
  XOR U3524 ( .A(n3713), .B(n3714), .Z(n3711) );
  AND U3525 ( .A(n34), .B(n3715), .Z(n3714) );
  XOR U3526 ( .A(p_input[2]), .B(n3713), .Z(n3715) );
  XOR U3527 ( .A(n3716), .B(n3717), .Z(n3713) );
  AND U3528 ( .A(n38), .B(n3718), .Z(n3717) );
  XOR U3529 ( .A(n3719), .B(n3720), .Z(n20) );
  AND U3530 ( .A(n42), .B(n3718), .Z(n3720) );
  XNOR U3531 ( .A(n3721), .B(n3716), .Z(n3718) );
  XOR U3532 ( .A(n3722), .B(n3723), .Z(n3716) );
  AND U3533 ( .A(n46), .B(n3724), .Z(n3723) );
  XOR U3534 ( .A(p_input[18]), .B(n3722), .Z(n3724) );
  XOR U3535 ( .A(n3725), .B(n3726), .Z(n3722) );
  AND U3536 ( .A(n50), .B(n3727), .Z(n3726) );
  IV U3537 ( .A(n3719), .Z(n3721) );
  XNOR U3538 ( .A(n3728), .B(n3729), .Z(n3719) );
  AND U3539 ( .A(n54), .B(n3727), .Z(n3729) );
  XNOR U3540 ( .A(n3728), .B(n3725), .Z(n3727) );
  XOR U3541 ( .A(n3730), .B(n3731), .Z(n3725) );
  AND U3542 ( .A(n57), .B(n3732), .Z(n3731) );
  XOR U3543 ( .A(p_input[34]), .B(n3730), .Z(n3732) );
  XOR U3544 ( .A(n3733), .B(n3734), .Z(n3730) );
  AND U3545 ( .A(n61), .B(n3735), .Z(n3734) );
  XOR U3546 ( .A(n3736), .B(n3737), .Z(n3728) );
  AND U3547 ( .A(n65), .B(n3735), .Z(n3737) );
  XNOR U3548 ( .A(n3736), .B(n3733), .Z(n3735) );
  XOR U3549 ( .A(n3738), .B(n3739), .Z(n3733) );
  AND U3550 ( .A(n68), .B(n3740), .Z(n3739) );
  XOR U3551 ( .A(p_input[50]), .B(n3738), .Z(n3740) );
  XOR U3552 ( .A(n3741), .B(n3742), .Z(n3738) );
  AND U3553 ( .A(n72), .B(n3743), .Z(n3742) );
  XOR U3554 ( .A(n3744), .B(n3745), .Z(n3736) );
  AND U3555 ( .A(n76), .B(n3743), .Z(n3745) );
  XNOR U3556 ( .A(n3744), .B(n3741), .Z(n3743) );
  XOR U3557 ( .A(n3746), .B(n3747), .Z(n3741) );
  AND U3558 ( .A(n79), .B(n3748), .Z(n3747) );
  XOR U3559 ( .A(p_input[66]), .B(n3746), .Z(n3748) );
  XOR U3560 ( .A(n3749), .B(n3750), .Z(n3746) );
  AND U3561 ( .A(n83), .B(n3751), .Z(n3750) );
  XOR U3562 ( .A(n3752), .B(n3753), .Z(n3744) );
  AND U3563 ( .A(n87), .B(n3751), .Z(n3753) );
  XNOR U3564 ( .A(n3752), .B(n3749), .Z(n3751) );
  XOR U3565 ( .A(n3754), .B(n3755), .Z(n3749) );
  AND U3566 ( .A(n90), .B(n3756), .Z(n3755) );
  XOR U3567 ( .A(p_input[82]), .B(n3754), .Z(n3756) );
  XOR U3568 ( .A(n3757), .B(n3758), .Z(n3754) );
  AND U3569 ( .A(n94), .B(n3759), .Z(n3758) );
  XOR U3570 ( .A(n3760), .B(n3761), .Z(n3752) );
  AND U3571 ( .A(n98), .B(n3759), .Z(n3761) );
  XNOR U3572 ( .A(n3760), .B(n3757), .Z(n3759) );
  XOR U3573 ( .A(n3762), .B(n3763), .Z(n3757) );
  AND U3574 ( .A(n101), .B(n3764), .Z(n3763) );
  XOR U3575 ( .A(p_input[98]), .B(n3762), .Z(n3764) );
  XOR U3576 ( .A(n3765), .B(n3766), .Z(n3762) );
  AND U3577 ( .A(n105), .B(n3767), .Z(n3766) );
  XOR U3578 ( .A(n3768), .B(n3769), .Z(n3760) );
  AND U3579 ( .A(n109), .B(n3767), .Z(n3769) );
  XNOR U3580 ( .A(n3768), .B(n3765), .Z(n3767) );
  XOR U3581 ( .A(n3770), .B(n3771), .Z(n3765) );
  AND U3582 ( .A(n112), .B(n3772), .Z(n3771) );
  XOR U3583 ( .A(p_input[114]), .B(n3770), .Z(n3772) );
  XOR U3584 ( .A(n3773), .B(n3774), .Z(n3770) );
  AND U3585 ( .A(n116), .B(n3775), .Z(n3774) );
  XOR U3586 ( .A(n3776), .B(n3777), .Z(n3768) );
  AND U3587 ( .A(n120), .B(n3775), .Z(n3777) );
  XNOR U3588 ( .A(n3776), .B(n3773), .Z(n3775) );
  XOR U3589 ( .A(n3778), .B(n3779), .Z(n3773) );
  AND U3590 ( .A(n123), .B(n3780), .Z(n3779) );
  XOR U3591 ( .A(p_input[130]), .B(n3778), .Z(n3780) );
  XOR U3592 ( .A(n3781), .B(n3782), .Z(n3778) );
  AND U3593 ( .A(n127), .B(n3783), .Z(n3782) );
  XOR U3594 ( .A(n3784), .B(n3785), .Z(n3776) );
  AND U3595 ( .A(n131), .B(n3783), .Z(n3785) );
  XNOR U3596 ( .A(n3784), .B(n3781), .Z(n3783) );
  XOR U3597 ( .A(n3786), .B(n3787), .Z(n3781) );
  AND U3598 ( .A(n134), .B(n3788), .Z(n3787) );
  XOR U3599 ( .A(p_input[146]), .B(n3786), .Z(n3788) );
  XOR U3600 ( .A(n3789), .B(n3790), .Z(n3786) );
  AND U3601 ( .A(n138), .B(n3791), .Z(n3790) );
  XOR U3602 ( .A(n3792), .B(n3793), .Z(n3784) );
  AND U3603 ( .A(n142), .B(n3791), .Z(n3793) );
  XNOR U3604 ( .A(n3792), .B(n3789), .Z(n3791) );
  XOR U3605 ( .A(n3794), .B(n3795), .Z(n3789) );
  AND U3606 ( .A(n145), .B(n3796), .Z(n3795) );
  XOR U3607 ( .A(p_input[162]), .B(n3794), .Z(n3796) );
  XOR U3608 ( .A(n3797), .B(n3798), .Z(n3794) );
  AND U3609 ( .A(n149), .B(n3799), .Z(n3798) );
  XOR U3610 ( .A(n3800), .B(n3801), .Z(n3792) );
  AND U3611 ( .A(n153), .B(n3799), .Z(n3801) );
  XNOR U3612 ( .A(n3800), .B(n3797), .Z(n3799) );
  XOR U3613 ( .A(n3802), .B(n3803), .Z(n3797) );
  AND U3614 ( .A(n156), .B(n3804), .Z(n3803) );
  XOR U3615 ( .A(p_input[178]), .B(n3802), .Z(n3804) );
  XOR U3616 ( .A(n3805), .B(n3806), .Z(n3802) );
  AND U3617 ( .A(n160), .B(n3807), .Z(n3806) );
  XOR U3618 ( .A(n3808), .B(n3809), .Z(n3800) );
  AND U3619 ( .A(n164), .B(n3807), .Z(n3809) );
  XNOR U3620 ( .A(n3808), .B(n3805), .Z(n3807) );
  XOR U3621 ( .A(n3810), .B(n3811), .Z(n3805) );
  AND U3622 ( .A(n167), .B(n3812), .Z(n3811) );
  XOR U3623 ( .A(p_input[194]), .B(n3810), .Z(n3812) );
  XOR U3624 ( .A(n3813), .B(n3814), .Z(n3810) );
  AND U3625 ( .A(n171), .B(n3815), .Z(n3814) );
  XOR U3626 ( .A(n3816), .B(n3817), .Z(n3808) );
  AND U3627 ( .A(n175), .B(n3815), .Z(n3817) );
  XNOR U3628 ( .A(n3816), .B(n3813), .Z(n3815) );
  XOR U3629 ( .A(n3818), .B(n3819), .Z(n3813) );
  AND U3630 ( .A(n178), .B(n3820), .Z(n3819) );
  XOR U3631 ( .A(p_input[210]), .B(n3818), .Z(n3820) );
  XOR U3632 ( .A(n3821), .B(n3822), .Z(n3818) );
  AND U3633 ( .A(n182), .B(n3823), .Z(n3822) );
  XOR U3634 ( .A(n3824), .B(n3825), .Z(n3816) );
  AND U3635 ( .A(n186), .B(n3823), .Z(n3825) );
  XNOR U3636 ( .A(n3824), .B(n3821), .Z(n3823) );
  XOR U3637 ( .A(n3826), .B(n3827), .Z(n3821) );
  AND U3638 ( .A(n189), .B(n3828), .Z(n3827) );
  XOR U3639 ( .A(p_input[226]), .B(n3826), .Z(n3828) );
  XOR U3640 ( .A(n3829), .B(n3830), .Z(n3826) );
  AND U3641 ( .A(n193), .B(n3831), .Z(n3830) );
  XOR U3642 ( .A(n3832), .B(n3833), .Z(n3824) );
  AND U3643 ( .A(n197), .B(n3831), .Z(n3833) );
  XNOR U3644 ( .A(n3832), .B(n3829), .Z(n3831) );
  XOR U3645 ( .A(n3834), .B(n3835), .Z(n3829) );
  AND U3646 ( .A(n200), .B(n3836), .Z(n3835) );
  XOR U3647 ( .A(p_input[242]), .B(n3834), .Z(n3836) );
  XOR U3648 ( .A(n3837), .B(n3838), .Z(n3834) );
  AND U3649 ( .A(n204), .B(n3839), .Z(n3838) );
  XOR U3650 ( .A(n3840), .B(n3841), .Z(n3832) );
  AND U3651 ( .A(n208), .B(n3839), .Z(n3841) );
  XNOR U3652 ( .A(n3840), .B(n3837), .Z(n3839) );
  XOR U3653 ( .A(n3842), .B(n3843), .Z(n3837) );
  AND U3654 ( .A(n211), .B(n3844), .Z(n3843) );
  XOR U3655 ( .A(p_input[258]), .B(n3842), .Z(n3844) );
  XOR U3656 ( .A(n3845), .B(n3846), .Z(n3842) );
  AND U3657 ( .A(n215), .B(n3847), .Z(n3846) );
  XOR U3658 ( .A(n3848), .B(n3849), .Z(n3840) );
  AND U3659 ( .A(n219), .B(n3847), .Z(n3849) );
  XNOR U3660 ( .A(n3848), .B(n3845), .Z(n3847) );
  XOR U3661 ( .A(n3850), .B(n3851), .Z(n3845) );
  AND U3662 ( .A(n222), .B(n3852), .Z(n3851) );
  XOR U3663 ( .A(p_input[274]), .B(n3850), .Z(n3852) );
  XOR U3664 ( .A(n3853), .B(n3854), .Z(n3850) );
  AND U3665 ( .A(n226), .B(n3855), .Z(n3854) );
  XOR U3666 ( .A(n3856), .B(n3857), .Z(n3848) );
  AND U3667 ( .A(n230), .B(n3855), .Z(n3857) );
  XNOR U3668 ( .A(n3856), .B(n3853), .Z(n3855) );
  XOR U3669 ( .A(n3858), .B(n3859), .Z(n3853) );
  AND U3670 ( .A(n233), .B(n3860), .Z(n3859) );
  XOR U3671 ( .A(p_input[290]), .B(n3858), .Z(n3860) );
  XOR U3672 ( .A(n3861), .B(n3862), .Z(n3858) );
  AND U3673 ( .A(n237), .B(n3863), .Z(n3862) );
  XOR U3674 ( .A(n3864), .B(n3865), .Z(n3856) );
  AND U3675 ( .A(n241), .B(n3863), .Z(n3865) );
  XNOR U3676 ( .A(n3864), .B(n3861), .Z(n3863) );
  XOR U3677 ( .A(n3866), .B(n3867), .Z(n3861) );
  AND U3678 ( .A(n244), .B(n3868), .Z(n3867) );
  XOR U3679 ( .A(p_input[306]), .B(n3866), .Z(n3868) );
  XOR U3680 ( .A(n3869), .B(n3870), .Z(n3866) );
  AND U3681 ( .A(n248), .B(n3871), .Z(n3870) );
  XOR U3682 ( .A(n3872), .B(n3873), .Z(n3864) );
  AND U3683 ( .A(n252), .B(n3871), .Z(n3873) );
  XNOR U3684 ( .A(n3872), .B(n3869), .Z(n3871) );
  XOR U3685 ( .A(n3874), .B(n3875), .Z(n3869) );
  AND U3686 ( .A(n255), .B(n3876), .Z(n3875) );
  XOR U3687 ( .A(p_input[322]), .B(n3874), .Z(n3876) );
  XOR U3688 ( .A(n3877), .B(n3878), .Z(n3874) );
  AND U3689 ( .A(n259), .B(n3879), .Z(n3878) );
  XOR U3690 ( .A(n3880), .B(n3881), .Z(n3872) );
  AND U3691 ( .A(n263), .B(n3879), .Z(n3881) );
  XNOR U3692 ( .A(n3880), .B(n3877), .Z(n3879) );
  XOR U3693 ( .A(n3882), .B(n3883), .Z(n3877) );
  AND U3694 ( .A(n266), .B(n3884), .Z(n3883) );
  XOR U3695 ( .A(p_input[338]), .B(n3882), .Z(n3884) );
  XOR U3696 ( .A(n3885), .B(n3886), .Z(n3882) );
  AND U3697 ( .A(n270), .B(n3887), .Z(n3886) );
  XOR U3698 ( .A(n3888), .B(n3889), .Z(n3880) );
  AND U3699 ( .A(n274), .B(n3887), .Z(n3889) );
  XNOR U3700 ( .A(n3888), .B(n3885), .Z(n3887) );
  XOR U3701 ( .A(n3890), .B(n3891), .Z(n3885) );
  AND U3702 ( .A(n277), .B(n3892), .Z(n3891) );
  XOR U3703 ( .A(p_input[354]), .B(n3890), .Z(n3892) );
  XOR U3704 ( .A(n3893), .B(n3894), .Z(n3890) );
  AND U3705 ( .A(n281), .B(n3895), .Z(n3894) );
  XOR U3706 ( .A(n3896), .B(n3897), .Z(n3888) );
  AND U3707 ( .A(n285), .B(n3895), .Z(n3897) );
  XNOR U3708 ( .A(n3896), .B(n3893), .Z(n3895) );
  XOR U3709 ( .A(n3898), .B(n3899), .Z(n3893) );
  AND U3710 ( .A(n288), .B(n3900), .Z(n3899) );
  XOR U3711 ( .A(p_input[370]), .B(n3898), .Z(n3900) );
  XOR U3712 ( .A(n3901), .B(n3902), .Z(n3898) );
  AND U3713 ( .A(n292), .B(n3903), .Z(n3902) );
  XOR U3714 ( .A(n3904), .B(n3905), .Z(n3896) );
  AND U3715 ( .A(n296), .B(n3903), .Z(n3905) );
  XNOR U3716 ( .A(n3904), .B(n3901), .Z(n3903) );
  XOR U3717 ( .A(n3906), .B(n3907), .Z(n3901) );
  AND U3718 ( .A(n299), .B(n3908), .Z(n3907) );
  XOR U3719 ( .A(p_input[386]), .B(n3906), .Z(n3908) );
  XOR U3720 ( .A(n3909), .B(n3910), .Z(n3906) );
  AND U3721 ( .A(n303), .B(n3911), .Z(n3910) );
  XOR U3722 ( .A(n3912), .B(n3913), .Z(n3904) );
  AND U3723 ( .A(n307), .B(n3911), .Z(n3913) );
  XNOR U3724 ( .A(n3912), .B(n3909), .Z(n3911) );
  XOR U3725 ( .A(n3914), .B(n3915), .Z(n3909) );
  AND U3726 ( .A(n310), .B(n3916), .Z(n3915) );
  XOR U3727 ( .A(p_input[402]), .B(n3914), .Z(n3916) );
  XOR U3728 ( .A(n3917), .B(n3918), .Z(n3914) );
  AND U3729 ( .A(n314), .B(n3919), .Z(n3918) );
  XOR U3730 ( .A(n3920), .B(n3921), .Z(n3912) );
  AND U3731 ( .A(n318), .B(n3919), .Z(n3921) );
  XNOR U3732 ( .A(n3920), .B(n3917), .Z(n3919) );
  XOR U3733 ( .A(n3922), .B(n3923), .Z(n3917) );
  AND U3734 ( .A(n321), .B(n3924), .Z(n3923) );
  XOR U3735 ( .A(p_input[418]), .B(n3922), .Z(n3924) );
  XOR U3736 ( .A(n3925), .B(n3926), .Z(n3922) );
  AND U3737 ( .A(n325), .B(n3927), .Z(n3926) );
  XOR U3738 ( .A(n3928), .B(n3929), .Z(n3920) );
  AND U3739 ( .A(n329), .B(n3927), .Z(n3929) );
  XNOR U3740 ( .A(n3928), .B(n3925), .Z(n3927) );
  XOR U3741 ( .A(n3930), .B(n3931), .Z(n3925) );
  AND U3742 ( .A(n332), .B(n3932), .Z(n3931) );
  XOR U3743 ( .A(p_input[434]), .B(n3930), .Z(n3932) );
  XOR U3744 ( .A(n3933), .B(n3934), .Z(n3930) );
  AND U3745 ( .A(n336), .B(n3935), .Z(n3934) );
  XOR U3746 ( .A(n3936), .B(n3937), .Z(n3928) );
  AND U3747 ( .A(n340), .B(n3935), .Z(n3937) );
  XNOR U3748 ( .A(n3936), .B(n3933), .Z(n3935) );
  XOR U3749 ( .A(n3938), .B(n3939), .Z(n3933) );
  AND U3750 ( .A(n343), .B(n3940), .Z(n3939) );
  XOR U3751 ( .A(p_input[450]), .B(n3938), .Z(n3940) );
  XOR U3752 ( .A(n3941), .B(n3942), .Z(n3938) );
  AND U3753 ( .A(n347), .B(n3943), .Z(n3942) );
  XOR U3754 ( .A(n3944), .B(n3945), .Z(n3936) );
  AND U3755 ( .A(n351), .B(n3943), .Z(n3945) );
  XNOR U3756 ( .A(n3944), .B(n3941), .Z(n3943) );
  XOR U3757 ( .A(n3946), .B(n3947), .Z(n3941) );
  AND U3758 ( .A(n354), .B(n3948), .Z(n3947) );
  XOR U3759 ( .A(p_input[466]), .B(n3946), .Z(n3948) );
  XOR U3760 ( .A(n3949), .B(n3950), .Z(n3946) );
  AND U3761 ( .A(n358), .B(n3951), .Z(n3950) );
  XOR U3762 ( .A(n3952), .B(n3953), .Z(n3944) );
  AND U3763 ( .A(n362), .B(n3951), .Z(n3953) );
  XNOR U3764 ( .A(n3952), .B(n3949), .Z(n3951) );
  XOR U3765 ( .A(n3954), .B(n3955), .Z(n3949) );
  AND U3766 ( .A(n365), .B(n3956), .Z(n3955) );
  XOR U3767 ( .A(p_input[482]), .B(n3954), .Z(n3956) );
  XOR U3768 ( .A(n3957), .B(n3958), .Z(n3954) );
  AND U3769 ( .A(n369), .B(n3959), .Z(n3958) );
  XOR U3770 ( .A(n3960), .B(n3961), .Z(n3952) );
  AND U3771 ( .A(n373), .B(n3959), .Z(n3961) );
  XNOR U3772 ( .A(n3960), .B(n3957), .Z(n3959) );
  XOR U3773 ( .A(n3962), .B(n3963), .Z(n3957) );
  AND U3774 ( .A(n376), .B(n3964), .Z(n3963) );
  XOR U3775 ( .A(p_input[498]), .B(n3962), .Z(n3964) );
  XOR U3776 ( .A(n3965), .B(n3966), .Z(n3962) );
  AND U3777 ( .A(n380), .B(n3967), .Z(n3966) );
  XOR U3778 ( .A(n3968), .B(n3969), .Z(n3960) );
  AND U3779 ( .A(n384), .B(n3967), .Z(n3969) );
  XNOR U3780 ( .A(n3968), .B(n3965), .Z(n3967) );
  XOR U3781 ( .A(n3970), .B(n3971), .Z(n3965) );
  AND U3782 ( .A(n387), .B(n3972), .Z(n3971) );
  XOR U3783 ( .A(p_input[514]), .B(n3970), .Z(n3972) );
  XOR U3784 ( .A(n3973), .B(n3974), .Z(n3970) );
  AND U3785 ( .A(n391), .B(n3975), .Z(n3974) );
  XOR U3786 ( .A(n3976), .B(n3977), .Z(n3968) );
  AND U3787 ( .A(n395), .B(n3975), .Z(n3977) );
  XNOR U3788 ( .A(n3976), .B(n3973), .Z(n3975) );
  XOR U3789 ( .A(n3978), .B(n3979), .Z(n3973) );
  AND U3790 ( .A(n398), .B(n3980), .Z(n3979) );
  XOR U3791 ( .A(p_input[530]), .B(n3978), .Z(n3980) );
  XOR U3792 ( .A(n3981), .B(n3982), .Z(n3978) );
  AND U3793 ( .A(n402), .B(n3983), .Z(n3982) );
  XOR U3794 ( .A(n3984), .B(n3985), .Z(n3976) );
  AND U3795 ( .A(n406), .B(n3983), .Z(n3985) );
  XNOR U3796 ( .A(n3984), .B(n3981), .Z(n3983) );
  XOR U3797 ( .A(n3986), .B(n3987), .Z(n3981) );
  AND U3798 ( .A(n409), .B(n3988), .Z(n3987) );
  XOR U3799 ( .A(p_input[546]), .B(n3986), .Z(n3988) );
  XOR U3800 ( .A(n3989), .B(n3990), .Z(n3986) );
  AND U3801 ( .A(n413), .B(n3991), .Z(n3990) );
  XOR U3802 ( .A(n3992), .B(n3993), .Z(n3984) );
  AND U3803 ( .A(n417), .B(n3991), .Z(n3993) );
  XNOR U3804 ( .A(n3992), .B(n3989), .Z(n3991) );
  XOR U3805 ( .A(n3994), .B(n3995), .Z(n3989) );
  AND U3806 ( .A(n420), .B(n3996), .Z(n3995) );
  XOR U3807 ( .A(p_input[562]), .B(n3994), .Z(n3996) );
  XOR U3808 ( .A(n3997), .B(n3998), .Z(n3994) );
  AND U3809 ( .A(n424), .B(n3999), .Z(n3998) );
  XOR U3810 ( .A(n4000), .B(n4001), .Z(n3992) );
  AND U3811 ( .A(n428), .B(n3999), .Z(n4001) );
  XNOR U3812 ( .A(n4000), .B(n3997), .Z(n3999) );
  XOR U3813 ( .A(n4002), .B(n4003), .Z(n3997) );
  AND U3814 ( .A(n431), .B(n4004), .Z(n4003) );
  XOR U3815 ( .A(p_input[578]), .B(n4002), .Z(n4004) );
  XOR U3816 ( .A(n4005), .B(n4006), .Z(n4002) );
  AND U3817 ( .A(n435), .B(n4007), .Z(n4006) );
  XOR U3818 ( .A(n4008), .B(n4009), .Z(n4000) );
  AND U3819 ( .A(n439), .B(n4007), .Z(n4009) );
  XNOR U3820 ( .A(n4008), .B(n4005), .Z(n4007) );
  XOR U3821 ( .A(n4010), .B(n4011), .Z(n4005) );
  AND U3822 ( .A(n442), .B(n4012), .Z(n4011) );
  XOR U3823 ( .A(p_input[594]), .B(n4010), .Z(n4012) );
  XOR U3824 ( .A(n4013), .B(n4014), .Z(n4010) );
  AND U3825 ( .A(n446), .B(n4015), .Z(n4014) );
  XOR U3826 ( .A(n4016), .B(n4017), .Z(n4008) );
  AND U3827 ( .A(n450), .B(n4015), .Z(n4017) );
  XNOR U3828 ( .A(n4016), .B(n4013), .Z(n4015) );
  XOR U3829 ( .A(n4018), .B(n4019), .Z(n4013) );
  AND U3830 ( .A(n453), .B(n4020), .Z(n4019) );
  XOR U3831 ( .A(p_input[610]), .B(n4018), .Z(n4020) );
  XOR U3832 ( .A(n4021), .B(n4022), .Z(n4018) );
  AND U3833 ( .A(n457), .B(n4023), .Z(n4022) );
  XOR U3834 ( .A(n4024), .B(n4025), .Z(n4016) );
  AND U3835 ( .A(n461), .B(n4023), .Z(n4025) );
  XNOR U3836 ( .A(n4024), .B(n4021), .Z(n4023) );
  XOR U3837 ( .A(n4026), .B(n4027), .Z(n4021) );
  AND U3838 ( .A(n464), .B(n4028), .Z(n4027) );
  XOR U3839 ( .A(p_input[626]), .B(n4026), .Z(n4028) );
  XOR U3840 ( .A(n4029), .B(n4030), .Z(n4026) );
  AND U3841 ( .A(n468), .B(n4031), .Z(n4030) );
  XOR U3842 ( .A(n4032), .B(n4033), .Z(n4024) );
  AND U3843 ( .A(n472), .B(n4031), .Z(n4033) );
  XNOR U3844 ( .A(n4032), .B(n4029), .Z(n4031) );
  XOR U3845 ( .A(n4034), .B(n4035), .Z(n4029) );
  AND U3846 ( .A(n475), .B(n4036), .Z(n4035) );
  XOR U3847 ( .A(p_input[642]), .B(n4034), .Z(n4036) );
  XOR U3848 ( .A(n4037), .B(n4038), .Z(n4034) );
  AND U3849 ( .A(n479), .B(n4039), .Z(n4038) );
  XOR U3850 ( .A(n4040), .B(n4041), .Z(n4032) );
  AND U3851 ( .A(n483), .B(n4039), .Z(n4041) );
  XNOR U3852 ( .A(n4040), .B(n4037), .Z(n4039) );
  XOR U3853 ( .A(n4042), .B(n4043), .Z(n4037) );
  AND U3854 ( .A(n486), .B(n4044), .Z(n4043) );
  XOR U3855 ( .A(p_input[658]), .B(n4042), .Z(n4044) );
  XOR U3856 ( .A(n4045), .B(n4046), .Z(n4042) );
  AND U3857 ( .A(n490), .B(n4047), .Z(n4046) );
  XOR U3858 ( .A(n4048), .B(n4049), .Z(n4040) );
  AND U3859 ( .A(n494), .B(n4047), .Z(n4049) );
  XNOR U3860 ( .A(n4048), .B(n4045), .Z(n4047) );
  XOR U3861 ( .A(n4050), .B(n4051), .Z(n4045) );
  AND U3862 ( .A(n497), .B(n4052), .Z(n4051) );
  XOR U3863 ( .A(p_input[674]), .B(n4050), .Z(n4052) );
  XOR U3864 ( .A(n4053), .B(n4054), .Z(n4050) );
  AND U3865 ( .A(n501), .B(n4055), .Z(n4054) );
  XOR U3866 ( .A(n4056), .B(n4057), .Z(n4048) );
  AND U3867 ( .A(n505), .B(n4055), .Z(n4057) );
  XNOR U3868 ( .A(n4056), .B(n4053), .Z(n4055) );
  XOR U3869 ( .A(n4058), .B(n4059), .Z(n4053) );
  AND U3870 ( .A(n508), .B(n4060), .Z(n4059) );
  XOR U3871 ( .A(p_input[690]), .B(n4058), .Z(n4060) );
  XOR U3872 ( .A(n4061), .B(n4062), .Z(n4058) );
  AND U3873 ( .A(n512), .B(n4063), .Z(n4062) );
  XOR U3874 ( .A(n4064), .B(n4065), .Z(n4056) );
  AND U3875 ( .A(n516), .B(n4063), .Z(n4065) );
  XNOR U3876 ( .A(n4064), .B(n4061), .Z(n4063) );
  XOR U3877 ( .A(n4066), .B(n4067), .Z(n4061) );
  AND U3878 ( .A(n519), .B(n4068), .Z(n4067) );
  XOR U3879 ( .A(p_input[706]), .B(n4066), .Z(n4068) );
  XOR U3880 ( .A(n4069), .B(n4070), .Z(n4066) );
  AND U3881 ( .A(n523), .B(n4071), .Z(n4070) );
  XOR U3882 ( .A(n4072), .B(n4073), .Z(n4064) );
  AND U3883 ( .A(n527), .B(n4071), .Z(n4073) );
  XNOR U3884 ( .A(n4072), .B(n4069), .Z(n4071) );
  XOR U3885 ( .A(n4074), .B(n4075), .Z(n4069) );
  AND U3886 ( .A(n530), .B(n4076), .Z(n4075) );
  XOR U3887 ( .A(p_input[722]), .B(n4074), .Z(n4076) );
  XOR U3888 ( .A(n4077), .B(n4078), .Z(n4074) );
  AND U3889 ( .A(n534), .B(n4079), .Z(n4078) );
  XOR U3890 ( .A(n4080), .B(n4081), .Z(n4072) );
  AND U3891 ( .A(n538), .B(n4079), .Z(n4081) );
  XNOR U3892 ( .A(n4080), .B(n4077), .Z(n4079) );
  XOR U3893 ( .A(n4082), .B(n4083), .Z(n4077) );
  AND U3894 ( .A(n541), .B(n4084), .Z(n4083) );
  XOR U3895 ( .A(p_input[738]), .B(n4082), .Z(n4084) );
  XOR U3896 ( .A(n4085), .B(n4086), .Z(n4082) );
  AND U3897 ( .A(n545), .B(n4087), .Z(n4086) );
  XOR U3898 ( .A(n4088), .B(n4089), .Z(n4080) );
  AND U3899 ( .A(n549), .B(n4087), .Z(n4089) );
  XNOR U3900 ( .A(n4088), .B(n4085), .Z(n4087) );
  XOR U3901 ( .A(n4090), .B(n4091), .Z(n4085) );
  AND U3902 ( .A(n552), .B(n4092), .Z(n4091) );
  XOR U3903 ( .A(p_input[754]), .B(n4090), .Z(n4092) );
  XOR U3904 ( .A(n4093), .B(n4094), .Z(n4090) );
  AND U3905 ( .A(n556), .B(n4095), .Z(n4094) );
  XOR U3906 ( .A(n4096), .B(n4097), .Z(n4088) );
  AND U3907 ( .A(n560), .B(n4095), .Z(n4097) );
  XNOR U3908 ( .A(n4096), .B(n4093), .Z(n4095) );
  XOR U3909 ( .A(n4098), .B(n4099), .Z(n4093) );
  AND U3910 ( .A(n563), .B(n4100), .Z(n4099) );
  XOR U3911 ( .A(p_input[770]), .B(n4098), .Z(n4100) );
  XOR U3912 ( .A(n4101), .B(n4102), .Z(n4098) );
  AND U3913 ( .A(n567), .B(n4103), .Z(n4102) );
  XOR U3914 ( .A(n4104), .B(n4105), .Z(n4096) );
  AND U3915 ( .A(n571), .B(n4103), .Z(n4105) );
  XNOR U3916 ( .A(n4104), .B(n4101), .Z(n4103) );
  XOR U3917 ( .A(n4106), .B(n4107), .Z(n4101) );
  AND U3918 ( .A(n574), .B(n4108), .Z(n4107) );
  XOR U3919 ( .A(p_input[786]), .B(n4106), .Z(n4108) );
  XOR U3920 ( .A(n4109), .B(n4110), .Z(n4106) );
  AND U3921 ( .A(n578), .B(n4111), .Z(n4110) );
  XOR U3922 ( .A(n4112), .B(n4113), .Z(n4104) );
  AND U3923 ( .A(n582), .B(n4111), .Z(n4113) );
  XNOR U3924 ( .A(n4112), .B(n4109), .Z(n4111) );
  XOR U3925 ( .A(n4114), .B(n4115), .Z(n4109) );
  AND U3926 ( .A(n585), .B(n4116), .Z(n4115) );
  XOR U3927 ( .A(p_input[802]), .B(n4114), .Z(n4116) );
  XOR U3928 ( .A(n4117), .B(n4118), .Z(n4114) );
  AND U3929 ( .A(n589), .B(n4119), .Z(n4118) );
  XOR U3930 ( .A(n4120), .B(n4121), .Z(n4112) );
  AND U3931 ( .A(n593), .B(n4119), .Z(n4121) );
  XNOR U3932 ( .A(n4120), .B(n4117), .Z(n4119) );
  XOR U3933 ( .A(n4122), .B(n4123), .Z(n4117) );
  AND U3934 ( .A(n596), .B(n4124), .Z(n4123) );
  XOR U3935 ( .A(p_input[818]), .B(n4122), .Z(n4124) );
  XOR U3936 ( .A(n4125), .B(n4126), .Z(n4122) );
  AND U3937 ( .A(n600), .B(n4127), .Z(n4126) );
  XOR U3938 ( .A(n4128), .B(n4129), .Z(n4120) );
  AND U3939 ( .A(n604), .B(n4127), .Z(n4129) );
  XNOR U3940 ( .A(n4128), .B(n4125), .Z(n4127) );
  XOR U3941 ( .A(n4130), .B(n4131), .Z(n4125) );
  AND U3942 ( .A(n607), .B(n4132), .Z(n4131) );
  XOR U3943 ( .A(p_input[834]), .B(n4130), .Z(n4132) );
  XOR U3944 ( .A(n4133), .B(n4134), .Z(n4130) );
  AND U3945 ( .A(n611), .B(n4135), .Z(n4134) );
  XOR U3946 ( .A(n4136), .B(n4137), .Z(n4128) );
  AND U3947 ( .A(n615), .B(n4135), .Z(n4137) );
  XNOR U3948 ( .A(n4136), .B(n4133), .Z(n4135) );
  XOR U3949 ( .A(n4138), .B(n4139), .Z(n4133) );
  AND U3950 ( .A(n618), .B(n4140), .Z(n4139) );
  XOR U3951 ( .A(p_input[850]), .B(n4138), .Z(n4140) );
  XOR U3952 ( .A(n4141), .B(n4142), .Z(n4138) );
  AND U3953 ( .A(n622), .B(n4143), .Z(n4142) );
  XOR U3954 ( .A(n4144), .B(n4145), .Z(n4136) );
  AND U3955 ( .A(n626), .B(n4143), .Z(n4145) );
  XNOR U3956 ( .A(n4144), .B(n4141), .Z(n4143) );
  XOR U3957 ( .A(n4146), .B(n4147), .Z(n4141) );
  AND U3958 ( .A(n629), .B(n4148), .Z(n4147) );
  XOR U3959 ( .A(p_input[866]), .B(n4146), .Z(n4148) );
  XOR U3960 ( .A(n4149), .B(n4150), .Z(n4146) );
  AND U3961 ( .A(n633), .B(n4151), .Z(n4150) );
  XOR U3962 ( .A(n4152), .B(n4153), .Z(n4144) );
  AND U3963 ( .A(n637), .B(n4151), .Z(n4153) );
  XNOR U3964 ( .A(n4152), .B(n4149), .Z(n4151) );
  XOR U3965 ( .A(n4154), .B(n4155), .Z(n4149) );
  AND U3966 ( .A(n640), .B(n4156), .Z(n4155) );
  XOR U3967 ( .A(p_input[882]), .B(n4154), .Z(n4156) );
  XOR U3968 ( .A(n4157), .B(n4158), .Z(n4154) );
  AND U3969 ( .A(n644), .B(n4159), .Z(n4158) );
  XOR U3970 ( .A(n4160), .B(n4161), .Z(n4152) );
  AND U3971 ( .A(n648), .B(n4159), .Z(n4161) );
  XNOR U3972 ( .A(n4160), .B(n4157), .Z(n4159) );
  XOR U3973 ( .A(n4162), .B(n4163), .Z(n4157) );
  AND U3974 ( .A(n651), .B(n4164), .Z(n4163) );
  XOR U3975 ( .A(p_input[898]), .B(n4162), .Z(n4164) );
  XOR U3976 ( .A(n4165), .B(n4166), .Z(n4162) );
  AND U3977 ( .A(n655), .B(n4167), .Z(n4166) );
  XOR U3978 ( .A(n4168), .B(n4169), .Z(n4160) );
  AND U3979 ( .A(n659), .B(n4167), .Z(n4169) );
  XNOR U3980 ( .A(n4168), .B(n4165), .Z(n4167) );
  XOR U3981 ( .A(n4170), .B(n4171), .Z(n4165) );
  AND U3982 ( .A(n662), .B(n4172), .Z(n4171) );
  XOR U3983 ( .A(p_input[914]), .B(n4170), .Z(n4172) );
  XOR U3984 ( .A(n4173), .B(n4174), .Z(n4170) );
  AND U3985 ( .A(n666), .B(n4175), .Z(n4174) );
  XOR U3986 ( .A(n4176), .B(n4177), .Z(n4168) );
  AND U3987 ( .A(n670), .B(n4175), .Z(n4177) );
  XNOR U3988 ( .A(n4176), .B(n4173), .Z(n4175) );
  XOR U3989 ( .A(n4178), .B(n4179), .Z(n4173) );
  AND U3990 ( .A(n673), .B(n4180), .Z(n4179) );
  XOR U3991 ( .A(p_input[930]), .B(n4178), .Z(n4180) );
  XOR U3992 ( .A(n4181), .B(n4182), .Z(n4178) );
  AND U3993 ( .A(n677), .B(n4183), .Z(n4182) );
  XOR U3994 ( .A(n4184), .B(n4185), .Z(n4176) );
  AND U3995 ( .A(n681), .B(n4183), .Z(n4185) );
  XNOR U3996 ( .A(n4184), .B(n4181), .Z(n4183) );
  XOR U3997 ( .A(n4186), .B(n4187), .Z(n4181) );
  AND U3998 ( .A(n684), .B(n4188), .Z(n4187) );
  XOR U3999 ( .A(p_input[946]), .B(n4186), .Z(n4188) );
  XOR U4000 ( .A(n4189), .B(n4190), .Z(n4186) );
  AND U4001 ( .A(n688), .B(n4191), .Z(n4190) );
  XOR U4002 ( .A(n4192), .B(n4193), .Z(n4184) );
  AND U4003 ( .A(n692), .B(n4191), .Z(n4193) );
  XNOR U4004 ( .A(n4192), .B(n4189), .Z(n4191) );
  XOR U4005 ( .A(n4194), .B(n4195), .Z(n4189) );
  AND U4006 ( .A(n695), .B(n4196), .Z(n4195) );
  XOR U4007 ( .A(p_input[962]), .B(n4194), .Z(n4196) );
  XOR U4008 ( .A(n4197), .B(n4198), .Z(n4194) );
  AND U4009 ( .A(n699), .B(n4199), .Z(n4198) );
  XOR U4010 ( .A(n4200), .B(n4201), .Z(n4192) );
  AND U4011 ( .A(n703), .B(n4199), .Z(n4201) );
  XNOR U4012 ( .A(n4200), .B(n4197), .Z(n4199) );
  XOR U4013 ( .A(n4202), .B(n4203), .Z(n4197) );
  AND U4014 ( .A(n706), .B(n4204), .Z(n4203) );
  XOR U4015 ( .A(p_input[978]), .B(n4202), .Z(n4204) );
  XNOR U4016 ( .A(n4205), .B(n4206), .Z(n4202) );
  AND U4017 ( .A(n710), .B(n4207), .Z(n4206) );
  XNOR U4018 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n4208), .Z(n4200) );
  AND U4019 ( .A(n713), .B(n4207), .Z(n4208) );
  XOR U4020 ( .A(n4209), .B(n4205), .Z(n4207) );
  XOR U4021 ( .A(n3210), .B(n4210), .Z(o[17]) );
  AND U4022 ( .A(n30), .B(n4211), .Z(n3210) );
  XOR U4023 ( .A(n3211), .B(n4210), .Z(n4211) );
  XOR U4024 ( .A(n4212), .B(n4213), .Z(n4210) );
  AND U4025 ( .A(n34), .B(n4214), .Z(n4213) );
  XOR U4026 ( .A(p_input[1]), .B(n4212), .Z(n4214) );
  XOR U4027 ( .A(n4215), .B(n4216), .Z(n4212) );
  AND U4028 ( .A(n38), .B(n4217), .Z(n4216) );
  XOR U4029 ( .A(n4218), .B(n4219), .Z(n3211) );
  AND U4030 ( .A(n42), .B(n4217), .Z(n4219) );
  XNOR U4031 ( .A(n4220), .B(n4215), .Z(n4217) );
  XOR U4032 ( .A(n4221), .B(n4222), .Z(n4215) );
  AND U4033 ( .A(n46), .B(n4223), .Z(n4222) );
  XOR U4034 ( .A(p_input[17]), .B(n4221), .Z(n4223) );
  XOR U4035 ( .A(n4224), .B(n4225), .Z(n4221) );
  AND U4036 ( .A(n50), .B(n4226), .Z(n4225) );
  IV U4037 ( .A(n4218), .Z(n4220) );
  XNOR U4038 ( .A(n4227), .B(n4228), .Z(n4218) );
  AND U4039 ( .A(n54), .B(n4226), .Z(n4228) );
  XNOR U4040 ( .A(n4227), .B(n4224), .Z(n4226) );
  XOR U4041 ( .A(n4229), .B(n4230), .Z(n4224) );
  AND U4042 ( .A(n57), .B(n4231), .Z(n4230) );
  XOR U4043 ( .A(p_input[33]), .B(n4229), .Z(n4231) );
  XOR U4044 ( .A(n4232), .B(n4233), .Z(n4229) );
  AND U4045 ( .A(n61), .B(n4234), .Z(n4233) );
  XOR U4046 ( .A(n4235), .B(n4236), .Z(n4227) );
  AND U4047 ( .A(n65), .B(n4234), .Z(n4236) );
  XNOR U4048 ( .A(n4235), .B(n4232), .Z(n4234) );
  XOR U4049 ( .A(n4237), .B(n4238), .Z(n4232) );
  AND U4050 ( .A(n68), .B(n4239), .Z(n4238) );
  XOR U4051 ( .A(p_input[49]), .B(n4237), .Z(n4239) );
  XOR U4052 ( .A(n4240), .B(n4241), .Z(n4237) );
  AND U4053 ( .A(n72), .B(n4242), .Z(n4241) );
  XOR U4054 ( .A(n4243), .B(n4244), .Z(n4235) );
  AND U4055 ( .A(n76), .B(n4242), .Z(n4244) );
  XNOR U4056 ( .A(n4243), .B(n4240), .Z(n4242) );
  XOR U4057 ( .A(n4245), .B(n4246), .Z(n4240) );
  AND U4058 ( .A(n79), .B(n4247), .Z(n4246) );
  XOR U4059 ( .A(p_input[65]), .B(n4245), .Z(n4247) );
  XOR U4060 ( .A(n4248), .B(n4249), .Z(n4245) );
  AND U4061 ( .A(n83), .B(n4250), .Z(n4249) );
  XOR U4062 ( .A(n4251), .B(n4252), .Z(n4243) );
  AND U4063 ( .A(n87), .B(n4250), .Z(n4252) );
  XNOR U4064 ( .A(n4251), .B(n4248), .Z(n4250) );
  XOR U4065 ( .A(n4253), .B(n4254), .Z(n4248) );
  AND U4066 ( .A(n90), .B(n4255), .Z(n4254) );
  XOR U4067 ( .A(p_input[81]), .B(n4253), .Z(n4255) );
  XOR U4068 ( .A(n4256), .B(n4257), .Z(n4253) );
  AND U4069 ( .A(n94), .B(n4258), .Z(n4257) );
  XOR U4070 ( .A(n4259), .B(n4260), .Z(n4251) );
  AND U4071 ( .A(n98), .B(n4258), .Z(n4260) );
  XNOR U4072 ( .A(n4259), .B(n4256), .Z(n4258) );
  XOR U4073 ( .A(n4261), .B(n4262), .Z(n4256) );
  AND U4074 ( .A(n101), .B(n4263), .Z(n4262) );
  XOR U4075 ( .A(p_input[97]), .B(n4261), .Z(n4263) );
  XOR U4076 ( .A(n4264), .B(n4265), .Z(n4261) );
  AND U4077 ( .A(n105), .B(n4266), .Z(n4265) );
  XOR U4078 ( .A(n4267), .B(n4268), .Z(n4259) );
  AND U4079 ( .A(n109), .B(n4266), .Z(n4268) );
  XNOR U4080 ( .A(n4267), .B(n4264), .Z(n4266) );
  XOR U4081 ( .A(n4269), .B(n4270), .Z(n4264) );
  AND U4082 ( .A(n112), .B(n4271), .Z(n4270) );
  XOR U4083 ( .A(p_input[113]), .B(n4269), .Z(n4271) );
  XOR U4084 ( .A(n4272), .B(n4273), .Z(n4269) );
  AND U4085 ( .A(n116), .B(n4274), .Z(n4273) );
  XOR U4086 ( .A(n4275), .B(n4276), .Z(n4267) );
  AND U4087 ( .A(n120), .B(n4274), .Z(n4276) );
  XNOR U4088 ( .A(n4275), .B(n4272), .Z(n4274) );
  XOR U4089 ( .A(n4277), .B(n4278), .Z(n4272) );
  AND U4090 ( .A(n123), .B(n4279), .Z(n4278) );
  XOR U4091 ( .A(p_input[129]), .B(n4277), .Z(n4279) );
  XOR U4092 ( .A(n4280), .B(n4281), .Z(n4277) );
  AND U4093 ( .A(n127), .B(n4282), .Z(n4281) );
  XOR U4094 ( .A(n4283), .B(n4284), .Z(n4275) );
  AND U4095 ( .A(n131), .B(n4282), .Z(n4284) );
  XNOR U4096 ( .A(n4283), .B(n4280), .Z(n4282) );
  XOR U4097 ( .A(n4285), .B(n4286), .Z(n4280) );
  AND U4098 ( .A(n134), .B(n4287), .Z(n4286) );
  XOR U4099 ( .A(p_input[145]), .B(n4285), .Z(n4287) );
  XOR U4100 ( .A(n4288), .B(n4289), .Z(n4285) );
  AND U4101 ( .A(n138), .B(n4290), .Z(n4289) );
  XOR U4102 ( .A(n4291), .B(n4292), .Z(n4283) );
  AND U4103 ( .A(n142), .B(n4290), .Z(n4292) );
  XNOR U4104 ( .A(n4291), .B(n4288), .Z(n4290) );
  XOR U4105 ( .A(n4293), .B(n4294), .Z(n4288) );
  AND U4106 ( .A(n145), .B(n4295), .Z(n4294) );
  XOR U4107 ( .A(p_input[161]), .B(n4293), .Z(n4295) );
  XOR U4108 ( .A(n4296), .B(n4297), .Z(n4293) );
  AND U4109 ( .A(n149), .B(n4298), .Z(n4297) );
  XOR U4110 ( .A(n4299), .B(n4300), .Z(n4291) );
  AND U4111 ( .A(n153), .B(n4298), .Z(n4300) );
  XNOR U4112 ( .A(n4299), .B(n4296), .Z(n4298) );
  XOR U4113 ( .A(n4301), .B(n4302), .Z(n4296) );
  AND U4114 ( .A(n156), .B(n4303), .Z(n4302) );
  XOR U4115 ( .A(p_input[177]), .B(n4301), .Z(n4303) );
  XOR U4116 ( .A(n4304), .B(n4305), .Z(n4301) );
  AND U4117 ( .A(n160), .B(n4306), .Z(n4305) );
  XOR U4118 ( .A(n4307), .B(n4308), .Z(n4299) );
  AND U4119 ( .A(n164), .B(n4306), .Z(n4308) );
  XNOR U4120 ( .A(n4307), .B(n4304), .Z(n4306) );
  XOR U4121 ( .A(n4309), .B(n4310), .Z(n4304) );
  AND U4122 ( .A(n167), .B(n4311), .Z(n4310) );
  XOR U4123 ( .A(p_input[193]), .B(n4309), .Z(n4311) );
  XOR U4124 ( .A(n4312), .B(n4313), .Z(n4309) );
  AND U4125 ( .A(n171), .B(n4314), .Z(n4313) );
  XOR U4126 ( .A(n4315), .B(n4316), .Z(n4307) );
  AND U4127 ( .A(n175), .B(n4314), .Z(n4316) );
  XNOR U4128 ( .A(n4315), .B(n4312), .Z(n4314) );
  XOR U4129 ( .A(n4317), .B(n4318), .Z(n4312) );
  AND U4130 ( .A(n178), .B(n4319), .Z(n4318) );
  XOR U4131 ( .A(p_input[209]), .B(n4317), .Z(n4319) );
  XOR U4132 ( .A(n4320), .B(n4321), .Z(n4317) );
  AND U4133 ( .A(n182), .B(n4322), .Z(n4321) );
  XOR U4134 ( .A(n4323), .B(n4324), .Z(n4315) );
  AND U4135 ( .A(n186), .B(n4322), .Z(n4324) );
  XNOR U4136 ( .A(n4323), .B(n4320), .Z(n4322) );
  XOR U4137 ( .A(n4325), .B(n4326), .Z(n4320) );
  AND U4138 ( .A(n189), .B(n4327), .Z(n4326) );
  XOR U4139 ( .A(p_input[225]), .B(n4325), .Z(n4327) );
  XOR U4140 ( .A(n4328), .B(n4329), .Z(n4325) );
  AND U4141 ( .A(n193), .B(n4330), .Z(n4329) );
  XOR U4142 ( .A(n4331), .B(n4332), .Z(n4323) );
  AND U4143 ( .A(n197), .B(n4330), .Z(n4332) );
  XNOR U4144 ( .A(n4331), .B(n4328), .Z(n4330) );
  XOR U4145 ( .A(n4333), .B(n4334), .Z(n4328) );
  AND U4146 ( .A(n200), .B(n4335), .Z(n4334) );
  XOR U4147 ( .A(p_input[241]), .B(n4333), .Z(n4335) );
  XOR U4148 ( .A(n4336), .B(n4337), .Z(n4333) );
  AND U4149 ( .A(n204), .B(n4338), .Z(n4337) );
  XOR U4150 ( .A(n4339), .B(n4340), .Z(n4331) );
  AND U4151 ( .A(n208), .B(n4338), .Z(n4340) );
  XNOR U4152 ( .A(n4339), .B(n4336), .Z(n4338) );
  XOR U4153 ( .A(n4341), .B(n4342), .Z(n4336) );
  AND U4154 ( .A(n211), .B(n4343), .Z(n4342) );
  XOR U4155 ( .A(p_input[257]), .B(n4341), .Z(n4343) );
  XOR U4156 ( .A(n4344), .B(n4345), .Z(n4341) );
  AND U4157 ( .A(n215), .B(n4346), .Z(n4345) );
  XOR U4158 ( .A(n4347), .B(n4348), .Z(n4339) );
  AND U4159 ( .A(n219), .B(n4346), .Z(n4348) );
  XNOR U4160 ( .A(n4347), .B(n4344), .Z(n4346) );
  XOR U4161 ( .A(n4349), .B(n4350), .Z(n4344) );
  AND U4162 ( .A(n222), .B(n4351), .Z(n4350) );
  XOR U4163 ( .A(p_input[273]), .B(n4349), .Z(n4351) );
  XOR U4164 ( .A(n4352), .B(n4353), .Z(n4349) );
  AND U4165 ( .A(n226), .B(n4354), .Z(n4353) );
  XOR U4166 ( .A(n4355), .B(n4356), .Z(n4347) );
  AND U4167 ( .A(n230), .B(n4354), .Z(n4356) );
  XNOR U4168 ( .A(n4355), .B(n4352), .Z(n4354) );
  XOR U4169 ( .A(n4357), .B(n4358), .Z(n4352) );
  AND U4170 ( .A(n233), .B(n4359), .Z(n4358) );
  XOR U4171 ( .A(p_input[289]), .B(n4357), .Z(n4359) );
  XOR U4172 ( .A(n4360), .B(n4361), .Z(n4357) );
  AND U4173 ( .A(n237), .B(n4362), .Z(n4361) );
  XOR U4174 ( .A(n4363), .B(n4364), .Z(n4355) );
  AND U4175 ( .A(n241), .B(n4362), .Z(n4364) );
  XNOR U4176 ( .A(n4363), .B(n4360), .Z(n4362) );
  XOR U4177 ( .A(n4365), .B(n4366), .Z(n4360) );
  AND U4178 ( .A(n244), .B(n4367), .Z(n4366) );
  XOR U4179 ( .A(p_input[305]), .B(n4365), .Z(n4367) );
  XOR U4180 ( .A(n4368), .B(n4369), .Z(n4365) );
  AND U4181 ( .A(n248), .B(n4370), .Z(n4369) );
  XOR U4182 ( .A(n4371), .B(n4372), .Z(n4363) );
  AND U4183 ( .A(n252), .B(n4370), .Z(n4372) );
  XNOR U4184 ( .A(n4371), .B(n4368), .Z(n4370) );
  XOR U4185 ( .A(n4373), .B(n4374), .Z(n4368) );
  AND U4186 ( .A(n255), .B(n4375), .Z(n4374) );
  XOR U4187 ( .A(p_input[321]), .B(n4373), .Z(n4375) );
  XOR U4188 ( .A(n4376), .B(n4377), .Z(n4373) );
  AND U4189 ( .A(n259), .B(n4378), .Z(n4377) );
  XOR U4190 ( .A(n4379), .B(n4380), .Z(n4371) );
  AND U4191 ( .A(n263), .B(n4378), .Z(n4380) );
  XNOR U4192 ( .A(n4379), .B(n4376), .Z(n4378) );
  XOR U4193 ( .A(n4381), .B(n4382), .Z(n4376) );
  AND U4194 ( .A(n266), .B(n4383), .Z(n4382) );
  XOR U4195 ( .A(p_input[337]), .B(n4381), .Z(n4383) );
  XOR U4196 ( .A(n4384), .B(n4385), .Z(n4381) );
  AND U4197 ( .A(n270), .B(n4386), .Z(n4385) );
  XOR U4198 ( .A(n4387), .B(n4388), .Z(n4379) );
  AND U4199 ( .A(n274), .B(n4386), .Z(n4388) );
  XNOR U4200 ( .A(n4387), .B(n4384), .Z(n4386) );
  XOR U4201 ( .A(n4389), .B(n4390), .Z(n4384) );
  AND U4202 ( .A(n277), .B(n4391), .Z(n4390) );
  XOR U4203 ( .A(p_input[353]), .B(n4389), .Z(n4391) );
  XOR U4204 ( .A(n4392), .B(n4393), .Z(n4389) );
  AND U4205 ( .A(n281), .B(n4394), .Z(n4393) );
  XOR U4206 ( .A(n4395), .B(n4396), .Z(n4387) );
  AND U4207 ( .A(n285), .B(n4394), .Z(n4396) );
  XNOR U4208 ( .A(n4395), .B(n4392), .Z(n4394) );
  XOR U4209 ( .A(n4397), .B(n4398), .Z(n4392) );
  AND U4210 ( .A(n288), .B(n4399), .Z(n4398) );
  XOR U4211 ( .A(p_input[369]), .B(n4397), .Z(n4399) );
  XOR U4212 ( .A(n4400), .B(n4401), .Z(n4397) );
  AND U4213 ( .A(n292), .B(n4402), .Z(n4401) );
  XOR U4214 ( .A(n4403), .B(n4404), .Z(n4395) );
  AND U4215 ( .A(n296), .B(n4402), .Z(n4404) );
  XNOR U4216 ( .A(n4403), .B(n4400), .Z(n4402) );
  XOR U4217 ( .A(n4405), .B(n4406), .Z(n4400) );
  AND U4218 ( .A(n299), .B(n4407), .Z(n4406) );
  XOR U4219 ( .A(p_input[385]), .B(n4405), .Z(n4407) );
  XOR U4220 ( .A(n4408), .B(n4409), .Z(n4405) );
  AND U4221 ( .A(n303), .B(n4410), .Z(n4409) );
  XOR U4222 ( .A(n4411), .B(n4412), .Z(n4403) );
  AND U4223 ( .A(n307), .B(n4410), .Z(n4412) );
  XNOR U4224 ( .A(n4411), .B(n4408), .Z(n4410) );
  XOR U4225 ( .A(n4413), .B(n4414), .Z(n4408) );
  AND U4226 ( .A(n310), .B(n4415), .Z(n4414) );
  XOR U4227 ( .A(p_input[401]), .B(n4413), .Z(n4415) );
  XOR U4228 ( .A(n4416), .B(n4417), .Z(n4413) );
  AND U4229 ( .A(n314), .B(n4418), .Z(n4417) );
  XOR U4230 ( .A(n4419), .B(n4420), .Z(n4411) );
  AND U4231 ( .A(n318), .B(n4418), .Z(n4420) );
  XNOR U4232 ( .A(n4419), .B(n4416), .Z(n4418) );
  XOR U4233 ( .A(n4421), .B(n4422), .Z(n4416) );
  AND U4234 ( .A(n321), .B(n4423), .Z(n4422) );
  XOR U4235 ( .A(p_input[417]), .B(n4421), .Z(n4423) );
  XOR U4236 ( .A(n4424), .B(n4425), .Z(n4421) );
  AND U4237 ( .A(n325), .B(n4426), .Z(n4425) );
  XOR U4238 ( .A(n4427), .B(n4428), .Z(n4419) );
  AND U4239 ( .A(n329), .B(n4426), .Z(n4428) );
  XNOR U4240 ( .A(n4427), .B(n4424), .Z(n4426) );
  XOR U4241 ( .A(n4429), .B(n4430), .Z(n4424) );
  AND U4242 ( .A(n332), .B(n4431), .Z(n4430) );
  XOR U4243 ( .A(p_input[433]), .B(n4429), .Z(n4431) );
  XOR U4244 ( .A(n4432), .B(n4433), .Z(n4429) );
  AND U4245 ( .A(n336), .B(n4434), .Z(n4433) );
  XOR U4246 ( .A(n4435), .B(n4436), .Z(n4427) );
  AND U4247 ( .A(n340), .B(n4434), .Z(n4436) );
  XNOR U4248 ( .A(n4435), .B(n4432), .Z(n4434) );
  XOR U4249 ( .A(n4437), .B(n4438), .Z(n4432) );
  AND U4250 ( .A(n343), .B(n4439), .Z(n4438) );
  XOR U4251 ( .A(p_input[449]), .B(n4437), .Z(n4439) );
  XOR U4252 ( .A(n4440), .B(n4441), .Z(n4437) );
  AND U4253 ( .A(n347), .B(n4442), .Z(n4441) );
  XOR U4254 ( .A(n4443), .B(n4444), .Z(n4435) );
  AND U4255 ( .A(n351), .B(n4442), .Z(n4444) );
  XNOR U4256 ( .A(n4443), .B(n4440), .Z(n4442) );
  XOR U4257 ( .A(n4445), .B(n4446), .Z(n4440) );
  AND U4258 ( .A(n354), .B(n4447), .Z(n4446) );
  XOR U4259 ( .A(p_input[465]), .B(n4445), .Z(n4447) );
  XOR U4260 ( .A(n4448), .B(n4449), .Z(n4445) );
  AND U4261 ( .A(n358), .B(n4450), .Z(n4449) );
  XOR U4262 ( .A(n4451), .B(n4452), .Z(n4443) );
  AND U4263 ( .A(n362), .B(n4450), .Z(n4452) );
  XNOR U4264 ( .A(n4451), .B(n4448), .Z(n4450) );
  XOR U4265 ( .A(n4453), .B(n4454), .Z(n4448) );
  AND U4266 ( .A(n365), .B(n4455), .Z(n4454) );
  XOR U4267 ( .A(p_input[481]), .B(n4453), .Z(n4455) );
  XOR U4268 ( .A(n4456), .B(n4457), .Z(n4453) );
  AND U4269 ( .A(n369), .B(n4458), .Z(n4457) );
  XOR U4270 ( .A(n4459), .B(n4460), .Z(n4451) );
  AND U4271 ( .A(n373), .B(n4458), .Z(n4460) );
  XNOR U4272 ( .A(n4459), .B(n4456), .Z(n4458) );
  XOR U4273 ( .A(n4461), .B(n4462), .Z(n4456) );
  AND U4274 ( .A(n376), .B(n4463), .Z(n4462) );
  XOR U4275 ( .A(p_input[497]), .B(n4461), .Z(n4463) );
  XOR U4276 ( .A(n4464), .B(n4465), .Z(n4461) );
  AND U4277 ( .A(n380), .B(n4466), .Z(n4465) );
  XOR U4278 ( .A(n4467), .B(n4468), .Z(n4459) );
  AND U4279 ( .A(n384), .B(n4466), .Z(n4468) );
  XNOR U4280 ( .A(n4467), .B(n4464), .Z(n4466) );
  XOR U4281 ( .A(n4469), .B(n4470), .Z(n4464) );
  AND U4282 ( .A(n387), .B(n4471), .Z(n4470) );
  XOR U4283 ( .A(p_input[513]), .B(n4469), .Z(n4471) );
  XOR U4284 ( .A(n4472), .B(n4473), .Z(n4469) );
  AND U4285 ( .A(n391), .B(n4474), .Z(n4473) );
  XOR U4286 ( .A(n4475), .B(n4476), .Z(n4467) );
  AND U4287 ( .A(n395), .B(n4474), .Z(n4476) );
  XNOR U4288 ( .A(n4475), .B(n4472), .Z(n4474) );
  XOR U4289 ( .A(n4477), .B(n4478), .Z(n4472) );
  AND U4290 ( .A(n398), .B(n4479), .Z(n4478) );
  XOR U4291 ( .A(p_input[529]), .B(n4477), .Z(n4479) );
  XOR U4292 ( .A(n4480), .B(n4481), .Z(n4477) );
  AND U4293 ( .A(n402), .B(n4482), .Z(n4481) );
  XOR U4294 ( .A(n4483), .B(n4484), .Z(n4475) );
  AND U4295 ( .A(n406), .B(n4482), .Z(n4484) );
  XNOR U4296 ( .A(n4483), .B(n4480), .Z(n4482) );
  XOR U4297 ( .A(n4485), .B(n4486), .Z(n4480) );
  AND U4298 ( .A(n409), .B(n4487), .Z(n4486) );
  XOR U4299 ( .A(p_input[545]), .B(n4485), .Z(n4487) );
  XOR U4300 ( .A(n4488), .B(n4489), .Z(n4485) );
  AND U4301 ( .A(n413), .B(n4490), .Z(n4489) );
  XOR U4302 ( .A(n4491), .B(n4492), .Z(n4483) );
  AND U4303 ( .A(n417), .B(n4490), .Z(n4492) );
  XNOR U4304 ( .A(n4491), .B(n4488), .Z(n4490) );
  XOR U4305 ( .A(n4493), .B(n4494), .Z(n4488) );
  AND U4306 ( .A(n420), .B(n4495), .Z(n4494) );
  XOR U4307 ( .A(p_input[561]), .B(n4493), .Z(n4495) );
  XOR U4308 ( .A(n4496), .B(n4497), .Z(n4493) );
  AND U4309 ( .A(n424), .B(n4498), .Z(n4497) );
  XOR U4310 ( .A(n4499), .B(n4500), .Z(n4491) );
  AND U4311 ( .A(n428), .B(n4498), .Z(n4500) );
  XNOR U4312 ( .A(n4499), .B(n4496), .Z(n4498) );
  XOR U4313 ( .A(n4501), .B(n4502), .Z(n4496) );
  AND U4314 ( .A(n431), .B(n4503), .Z(n4502) );
  XOR U4315 ( .A(p_input[577]), .B(n4501), .Z(n4503) );
  XOR U4316 ( .A(n4504), .B(n4505), .Z(n4501) );
  AND U4317 ( .A(n435), .B(n4506), .Z(n4505) );
  XOR U4318 ( .A(n4507), .B(n4508), .Z(n4499) );
  AND U4319 ( .A(n439), .B(n4506), .Z(n4508) );
  XNOR U4320 ( .A(n4507), .B(n4504), .Z(n4506) );
  XOR U4321 ( .A(n4509), .B(n4510), .Z(n4504) );
  AND U4322 ( .A(n442), .B(n4511), .Z(n4510) );
  XOR U4323 ( .A(p_input[593]), .B(n4509), .Z(n4511) );
  XOR U4324 ( .A(n4512), .B(n4513), .Z(n4509) );
  AND U4325 ( .A(n446), .B(n4514), .Z(n4513) );
  XOR U4326 ( .A(n4515), .B(n4516), .Z(n4507) );
  AND U4327 ( .A(n450), .B(n4514), .Z(n4516) );
  XNOR U4328 ( .A(n4515), .B(n4512), .Z(n4514) );
  XOR U4329 ( .A(n4517), .B(n4518), .Z(n4512) );
  AND U4330 ( .A(n453), .B(n4519), .Z(n4518) );
  XOR U4331 ( .A(p_input[609]), .B(n4517), .Z(n4519) );
  XOR U4332 ( .A(n4520), .B(n4521), .Z(n4517) );
  AND U4333 ( .A(n457), .B(n4522), .Z(n4521) );
  XOR U4334 ( .A(n4523), .B(n4524), .Z(n4515) );
  AND U4335 ( .A(n461), .B(n4522), .Z(n4524) );
  XNOR U4336 ( .A(n4523), .B(n4520), .Z(n4522) );
  XOR U4337 ( .A(n4525), .B(n4526), .Z(n4520) );
  AND U4338 ( .A(n464), .B(n4527), .Z(n4526) );
  XOR U4339 ( .A(p_input[625]), .B(n4525), .Z(n4527) );
  XOR U4340 ( .A(n4528), .B(n4529), .Z(n4525) );
  AND U4341 ( .A(n468), .B(n4530), .Z(n4529) );
  XOR U4342 ( .A(n4531), .B(n4532), .Z(n4523) );
  AND U4343 ( .A(n472), .B(n4530), .Z(n4532) );
  XNOR U4344 ( .A(n4531), .B(n4528), .Z(n4530) );
  XOR U4345 ( .A(n4533), .B(n4534), .Z(n4528) );
  AND U4346 ( .A(n475), .B(n4535), .Z(n4534) );
  XOR U4347 ( .A(p_input[641]), .B(n4533), .Z(n4535) );
  XOR U4348 ( .A(n4536), .B(n4537), .Z(n4533) );
  AND U4349 ( .A(n479), .B(n4538), .Z(n4537) );
  XOR U4350 ( .A(n4539), .B(n4540), .Z(n4531) );
  AND U4351 ( .A(n483), .B(n4538), .Z(n4540) );
  XNOR U4352 ( .A(n4539), .B(n4536), .Z(n4538) );
  XOR U4353 ( .A(n4541), .B(n4542), .Z(n4536) );
  AND U4354 ( .A(n486), .B(n4543), .Z(n4542) );
  XOR U4355 ( .A(p_input[657]), .B(n4541), .Z(n4543) );
  XOR U4356 ( .A(n4544), .B(n4545), .Z(n4541) );
  AND U4357 ( .A(n490), .B(n4546), .Z(n4545) );
  XOR U4358 ( .A(n4547), .B(n4548), .Z(n4539) );
  AND U4359 ( .A(n494), .B(n4546), .Z(n4548) );
  XNOR U4360 ( .A(n4547), .B(n4544), .Z(n4546) );
  XOR U4361 ( .A(n4549), .B(n4550), .Z(n4544) );
  AND U4362 ( .A(n497), .B(n4551), .Z(n4550) );
  XOR U4363 ( .A(p_input[673]), .B(n4549), .Z(n4551) );
  XOR U4364 ( .A(n4552), .B(n4553), .Z(n4549) );
  AND U4365 ( .A(n501), .B(n4554), .Z(n4553) );
  XOR U4366 ( .A(n4555), .B(n4556), .Z(n4547) );
  AND U4367 ( .A(n505), .B(n4554), .Z(n4556) );
  XNOR U4368 ( .A(n4555), .B(n4552), .Z(n4554) );
  XOR U4369 ( .A(n4557), .B(n4558), .Z(n4552) );
  AND U4370 ( .A(n508), .B(n4559), .Z(n4558) );
  XOR U4371 ( .A(p_input[689]), .B(n4557), .Z(n4559) );
  XOR U4372 ( .A(n4560), .B(n4561), .Z(n4557) );
  AND U4373 ( .A(n512), .B(n4562), .Z(n4561) );
  XOR U4374 ( .A(n4563), .B(n4564), .Z(n4555) );
  AND U4375 ( .A(n516), .B(n4562), .Z(n4564) );
  XNOR U4376 ( .A(n4563), .B(n4560), .Z(n4562) );
  XOR U4377 ( .A(n4565), .B(n4566), .Z(n4560) );
  AND U4378 ( .A(n519), .B(n4567), .Z(n4566) );
  XOR U4379 ( .A(p_input[705]), .B(n4565), .Z(n4567) );
  XOR U4380 ( .A(n4568), .B(n4569), .Z(n4565) );
  AND U4381 ( .A(n523), .B(n4570), .Z(n4569) );
  XOR U4382 ( .A(n4571), .B(n4572), .Z(n4563) );
  AND U4383 ( .A(n527), .B(n4570), .Z(n4572) );
  XNOR U4384 ( .A(n4571), .B(n4568), .Z(n4570) );
  XOR U4385 ( .A(n4573), .B(n4574), .Z(n4568) );
  AND U4386 ( .A(n530), .B(n4575), .Z(n4574) );
  XOR U4387 ( .A(p_input[721]), .B(n4573), .Z(n4575) );
  XOR U4388 ( .A(n4576), .B(n4577), .Z(n4573) );
  AND U4389 ( .A(n534), .B(n4578), .Z(n4577) );
  XOR U4390 ( .A(n4579), .B(n4580), .Z(n4571) );
  AND U4391 ( .A(n538), .B(n4578), .Z(n4580) );
  XNOR U4392 ( .A(n4579), .B(n4576), .Z(n4578) );
  XOR U4393 ( .A(n4581), .B(n4582), .Z(n4576) );
  AND U4394 ( .A(n541), .B(n4583), .Z(n4582) );
  XOR U4395 ( .A(p_input[737]), .B(n4581), .Z(n4583) );
  XOR U4396 ( .A(n4584), .B(n4585), .Z(n4581) );
  AND U4397 ( .A(n545), .B(n4586), .Z(n4585) );
  XOR U4398 ( .A(n4587), .B(n4588), .Z(n4579) );
  AND U4399 ( .A(n549), .B(n4586), .Z(n4588) );
  XNOR U4400 ( .A(n4587), .B(n4584), .Z(n4586) );
  XOR U4401 ( .A(n4589), .B(n4590), .Z(n4584) );
  AND U4402 ( .A(n552), .B(n4591), .Z(n4590) );
  XOR U4403 ( .A(p_input[753]), .B(n4589), .Z(n4591) );
  XOR U4404 ( .A(n4592), .B(n4593), .Z(n4589) );
  AND U4405 ( .A(n556), .B(n4594), .Z(n4593) );
  XOR U4406 ( .A(n4595), .B(n4596), .Z(n4587) );
  AND U4407 ( .A(n560), .B(n4594), .Z(n4596) );
  XNOR U4408 ( .A(n4595), .B(n4592), .Z(n4594) );
  XOR U4409 ( .A(n4597), .B(n4598), .Z(n4592) );
  AND U4410 ( .A(n563), .B(n4599), .Z(n4598) );
  XOR U4411 ( .A(p_input[769]), .B(n4597), .Z(n4599) );
  XOR U4412 ( .A(n4600), .B(n4601), .Z(n4597) );
  AND U4413 ( .A(n567), .B(n4602), .Z(n4601) );
  XOR U4414 ( .A(n4603), .B(n4604), .Z(n4595) );
  AND U4415 ( .A(n571), .B(n4602), .Z(n4604) );
  XNOR U4416 ( .A(n4603), .B(n4600), .Z(n4602) );
  XOR U4417 ( .A(n4605), .B(n4606), .Z(n4600) );
  AND U4418 ( .A(n574), .B(n4607), .Z(n4606) );
  XOR U4419 ( .A(p_input[785]), .B(n4605), .Z(n4607) );
  XOR U4420 ( .A(n4608), .B(n4609), .Z(n4605) );
  AND U4421 ( .A(n578), .B(n4610), .Z(n4609) );
  XOR U4422 ( .A(n4611), .B(n4612), .Z(n4603) );
  AND U4423 ( .A(n582), .B(n4610), .Z(n4612) );
  XNOR U4424 ( .A(n4611), .B(n4608), .Z(n4610) );
  XOR U4425 ( .A(n4613), .B(n4614), .Z(n4608) );
  AND U4426 ( .A(n585), .B(n4615), .Z(n4614) );
  XOR U4427 ( .A(p_input[801]), .B(n4613), .Z(n4615) );
  XOR U4428 ( .A(n4616), .B(n4617), .Z(n4613) );
  AND U4429 ( .A(n589), .B(n4618), .Z(n4617) );
  XOR U4430 ( .A(n4619), .B(n4620), .Z(n4611) );
  AND U4431 ( .A(n593), .B(n4618), .Z(n4620) );
  XNOR U4432 ( .A(n4619), .B(n4616), .Z(n4618) );
  XOR U4433 ( .A(n4621), .B(n4622), .Z(n4616) );
  AND U4434 ( .A(n596), .B(n4623), .Z(n4622) );
  XOR U4435 ( .A(p_input[817]), .B(n4621), .Z(n4623) );
  XOR U4436 ( .A(n4624), .B(n4625), .Z(n4621) );
  AND U4437 ( .A(n600), .B(n4626), .Z(n4625) );
  XOR U4438 ( .A(n4627), .B(n4628), .Z(n4619) );
  AND U4439 ( .A(n604), .B(n4626), .Z(n4628) );
  XNOR U4440 ( .A(n4627), .B(n4624), .Z(n4626) );
  XOR U4441 ( .A(n4629), .B(n4630), .Z(n4624) );
  AND U4442 ( .A(n607), .B(n4631), .Z(n4630) );
  XOR U4443 ( .A(p_input[833]), .B(n4629), .Z(n4631) );
  XOR U4444 ( .A(n4632), .B(n4633), .Z(n4629) );
  AND U4445 ( .A(n611), .B(n4634), .Z(n4633) );
  XOR U4446 ( .A(n4635), .B(n4636), .Z(n4627) );
  AND U4447 ( .A(n615), .B(n4634), .Z(n4636) );
  XNOR U4448 ( .A(n4635), .B(n4632), .Z(n4634) );
  XOR U4449 ( .A(n4637), .B(n4638), .Z(n4632) );
  AND U4450 ( .A(n618), .B(n4639), .Z(n4638) );
  XOR U4451 ( .A(p_input[849]), .B(n4637), .Z(n4639) );
  XOR U4452 ( .A(n4640), .B(n4641), .Z(n4637) );
  AND U4453 ( .A(n622), .B(n4642), .Z(n4641) );
  XOR U4454 ( .A(n4643), .B(n4644), .Z(n4635) );
  AND U4455 ( .A(n626), .B(n4642), .Z(n4644) );
  XNOR U4456 ( .A(n4643), .B(n4640), .Z(n4642) );
  XOR U4457 ( .A(n4645), .B(n4646), .Z(n4640) );
  AND U4458 ( .A(n629), .B(n4647), .Z(n4646) );
  XOR U4459 ( .A(p_input[865]), .B(n4645), .Z(n4647) );
  XOR U4460 ( .A(n4648), .B(n4649), .Z(n4645) );
  AND U4461 ( .A(n633), .B(n4650), .Z(n4649) );
  XOR U4462 ( .A(n4651), .B(n4652), .Z(n4643) );
  AND U4463 ( .A(n637), .B(n4650), .Z(n4652) );
  XNOR U4464 ( .A(n4651), .B(n4648), .Z(n4650) );
  XOR U4465 ( .A(n4653), .B(n4654), .Z(n4648) );
  AND U4466 ( .A(n640), .B(n4655), .Z(n4654) );
  XOR U4467 ( .A(p_input[881]), .B(n4653), .Z(n4655) );
  XOR U4468 ( .A(n4656), .B(n4657), .Z(n4653) );
  AND U4469 ( .A(n644), .B(n4658), .Z(n4657) );
  XOR U4470 ( .A(n4659), .B(n4660), .Z(n4651) );
  AND U4471 ( .A(n648), .B(n4658), .Z(n4660) );
  XNOR U4472 ( .A(n4659), .B(n4656), .Z(n4658) );
  XOR U4473 ( .A(n4661), .B(n4662), .Z(n4656) );
  AND U4474 ( .A(n651), .B(n4663), .Z(n4662) );
  XOR U4475 ( .A(p_input[897]), .B(n4661), .Z(n4663) );
  XOR U4476 ( .A(n4664), .B(n4665), .Z(n4661) );
  AND U4477 ( .A(n655), .B(n4666), .Z(n4665) );
  XOR U4478 ( .A(n4667), .B(n4668), .Z(n4659) );
  AND U4479 ( .A(n659), .B(n4666), .Z(n4668) );
  XNOR U4480 ( .A(n4667), .B(n4664), .Z(n4666) );
  XOR U4481 ( .A(n4669), .B(n4670), .Z(n4664) );
  AND U4482 ( .A(n662), .B(n4671), .Z(n4670) );
  XOR U4483 ( .A(p_input[913]), .B(n4669), .Z(n4671) );
  XOR U4484 ( .A(n4672), .B(n4673), .Z(n4669) );
  AND U4485 ( .A(n666), .B(n4674), .Z(n4673) );
  XOR U4486 ( .A(n4675), .B(n4676), .Z(n4667) );
  AND U4487 ( .A(n670), .B(n4674), .Z(n4676) );
  XNOR U4488 ( .A(n4675), .B(n4672), .Z(n4674) );
  XOR U4489 ( .A(n4677), .B(n4678), .Z(n4672) );
  AND U4490 ( .A(n673), .B(n4679), .Z(n4678) );
  XOR U4491 ( .A(p_input[929]), .B(n4677), .Z(n4679) );
  XOR U4492 ( .A(n4680), .B(n4681), .Z(n4677) );
  AND U4493 ( .A(n677), .B(n4682), .Z(n4681) );
  XOR U4494 ( .A(n4683), .B(n4684), .Z(n4675) );
  AND U4495 ( .A(n681), .B(n4682), .Z(n4684) );
  XNOR U4496 ( .A(n4683), .B(n4680), .Z(n4682) );
  XOR U4497 ( .A(n4685), .B(n4686), .Z(n4680) );
  AND U4498 ( .A(n684), .B(n4687), .Z(n4686) );
  XOR U4499 ( .A(p_input[945]), .B(n4685), .Z(n4687) );
  XOR U4500 ( .A(n4688), .B(n4689), .Z(n4685) );
  AND U4501 ( .A(n688), .B(n4690), .Z(n4689) );
  XOR U4502 ( .A(n4691), .B(n4692), .Z(n4683) );
  AND U4503 ( .A(n692), .B(n4690), .Z(n4692) );
  XNOR U4504 ( .A(n4691), .B(n4688), .Z(n4690) );
  XOR U4505 ( .A(n4693), .B(n4694), .Z(n4688) );
  AND U4506 ( .A(n695), .B(n4695), .Z(n4694) );
  XOR U4507 ( .A(p_input[961]), .B(n4693), .Z(n4695) );
  XOR U4508 ( .A(n4696), .B(n4697), .Z(n4693) );
  AND U4509 ( .A(n699), .B(n4698), .Z(n4697) );
  XOR U4510 ( .A(n4699), .B(n4700), .Z(n4691) );
  AND U4511 ( .A(n703), .B(n4698), .Z(n4700) );
  XNOR U4512 ( .A(n4699), .B(n4696), .Z(n4698) );
  XOR U4513 ( .A(n4701), .B(n4702), .Z(n4696) );
  AND U4514 ( .A(n706), .B(n4703), .Z(n4702) );
  XOR U4515 ( .A(p_input[977]), .B(n4701), .Z(n4703) );
  XNOR U4516 ( .A(n4704), .B(n4705), .Z(n4701) );
  AND U4517 ( .A(n710), .B(n4706), .Z(n4705) );
  XNOR U4518 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n4707), .Z(n4699) );
  AND U4519 ( .A(n713), .B(n4706), .Z(n4707) );
  XOR U4520 ( .A(n4708), .B(n4704), .Z(n4706) );
  IV U4521 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n4704) );
  XOR U4522 ( .A(n4709), .B(n4710), .Z(o[16]) );
  XOR U4523 ( .A(n15), .B(n4711), .Z(o[15]) );
  AND U4524 ( .A(n30), .B(n4712), .Z(n15) );
  XOR U4525 ( .A(n16), .B(n4711), .Z(n4712) );
  XOR U4526 ( .A(n4713), .B(n4714), .Z(n4711) );
  AND U4527 ( .A(n42), .B(n4715), .Z(n4714) );
  XOR U4528 ( .A(n4716), .B(n4717), .Z(n16) );
  AND U4529 ( .A(n34), .B(n4718), .Z(n4717) );
  XOR U4530 ( .A(p_input[15]), .B(n4716), .Z(n4718) );
  XNOR U4531 ( .A(n4719), .B(n4720), .Z(n4716) );
  AND U4532 ( .A(n38), .B(n4715), .Z(n4720) );
  XNOR U4533 ( .A(n4719), .B(n4713), .Z(n4715) );
  XOR U4534 ( .A(n4721), .B(n4722), .Z(n4713) );
  AND U4535 ( .A(n54), .B(n4723), .Z(n4722) );
  XNOR U4536 ( .A(n4724), .B(n4725), .Z(n4719) );
  AND U4537 ( .A(n46), .B(n4726), .Z(n4725) );
  XOR U4538 ( .A(p_input[31]), .B(n4724), .Z(n4726) );
  XNOR U4539 ( .A(n4727), .B(n4728), .Z(n4724) );
  AND U4540 ( .A(n50), .B(n4723), .Z(n4728) );
  XNOR U4541 ( .A(n4727), .B(n4721), .Z(n4723) );
  XOR U4542 ( .A(n4729), .B(n4730), .Z(n4721) );
  AND U4543 ( .A(n65), .B(n4731), .Z(n4730) );
  XNOR U4544 ( .A(n4732), .B(n4733), .Z(n4727) );
  AND U4545 ( .A(n57), .B(n4734), .Z(n4733) );
  XOR U4546 ( .A(p_input[47]), .B(n4732), .Z(n4734) );
  XNOR U4547 ( .A(n4735), .B(n4736), .Z(n4732) );
  AND U4548 ( .A(n61), .B(n4731), .Z(n4736) );
  XNOR U4549 ( .A(n4735), .B(n4729), .Z(n4731) );
  XOR U4550 ( .A(n4737), .B(n4738), .Z(n4729) );
  AND U4551 ( .A(n76), .B(n4739), .Z(n4738) );
  XNOR U4552 ( .A(n4740), .B(n4741), .Z(n4735) );
  AND U4553 ( .A(n68), .B(n4742), .Z(n4741) );
  XOR U4554 ( .A(p_input[63]), .B(n4740), .Z(n4742) );
  XNOR U4555 ( .A(n4743), .B(n4744), .Z(n4740) );
  AND U4556 ( .A(n72), .B(n4739), .Z(n4744) );
  XNOR U4557 ( .A(n4743), .B(n4737), .Z(n4739) );
  XOR U4558 ( .A(n4745), .B(n4746), .Z(n4737) );
  AND U4559 ( .A(n87), .B(n4747), .Z(n4746) );
  XNOR U4560 ( .A(n4748), .B(n4749), .Z(n4743) );
  AND U4561 ( .A(n79), .B(n4750), .Z(n4749) );
  XOR U4562 ( .A(p_input[79]), .B(n4748), .Z(n4750) );
  XNOR U4563 ( .A(n4751), .B(n4752), .Z(n4748) );
  AND U4564 ( .A(n83), .B(n4747), .Z(n4752) );
  XNOR U4565 ( .A(n4751), .B(n4745), .Z(n4747) );
  XOR U4566 ( .A(n4753), .B(n4754), .Z(n4745) );
  AND U4567 ( .A(n98), .B(n4755), .Z(n4754) );
  XNOR U4568 ( .A(n4756), .B(n4757), .Z(n4751) );
  AND U4569 ( .A(n90), .B(n4758), .Z(n4757) );
  XOR U4570 ( .A(p_input[95]), .B(n4756), .Z(n4758) );
  XNOR U4571 ( .A(n4759), .B(n4760), .Z(n4756) );
  AND U4572 ( .A(n94), .B(n4755), .Z(n4760) );
  XNOR U4573 ( .A(n4759), .B(n4753), .Z(n4755) );
  XOR U4574 ( .A(n4761), .B(n4762), .Z(n4753) );
  AND U4575 ( .A(n109), .B(n4763), .Z(n4762) );
  XNOR U4576 ( .A(n4764), .B(n4765), .Z(n4759) );
  AND U4577 ( .A(n101), .B(n4766), .Z(n4765) );
  XOR U4578 ( .A(p_input[111]), .B(n4764), .Z(n4766) );
  XNOR U4579 ( .A(n4767), .B(n4768), .Z(n4764) );
  AND U4580 ( .A(n105), .B(n4763), .Z(n4768) );
  XNOR U4581 ( .A(n4767), .B(n4761), .Z(n4763) );
  XOR U4582 ( .A(n4769), .B(n4770), .Z(n4761) );
  AND U4583 ( .A(n120), .B(n4771), .Z(n4770) );
  XNOR U4584 ( .A(n4772), .B(n4773), .Z(n4767) );
  AND U4585 ( .A(n112), .B(n4774), .Z(n4773) );
  XOR U4586 ( .A(p_input[127]), .B(n4772), .Z(n4774) );
  XNOR U4587 ( .A(n4775), .B(n4776), .Z(n4772) );
  AND U4588 ( .A(n116), .B(n4771), .Z(n4776) );
  XNOR U4589 ( .A(n4775), .B(n4769), .Z(n4771) );
  XOR U4590 ( .A(n4777), .B(n4778), .Z(n4769) );
  AND U4591 ( .A(n131), .B(n4779), .Z(n4778) );
  XNOR U4592 ( .A(n4780), .B(n4781), .Z(n4775) );
  AND U4593 ( .A(n123), .B(n4782), .Z(n4781) );
  XOR U4594 ( .A(p_input[143]), .B(n4780), .Z(n4782) );
  XNOR U4595 ( .A(n4783), .B(n4784), .Z(n4780) );
  AND U4596 ( .A(n127), .B(n4779), .Z(n4784) );
  XNOR U4597 ( .A(n4783), .B(n4777), .Z(n4779) );
  XOR U4598 ( .A(n4785), .B(n4786), .Z(n4777) );
  AND U4599 ( .A(n142), .B(n4787), .Z(n4786) );
  XNOR U4600 ( .A(n4788), .B(n4789), .Z(n4783) );
  AND U4601 ( .A(n134), .B(n4790), .Z(n4789) );
  XOR U4602 ( .A(p_input[159]), .B(n4788), .Z(n4790) );
  XNOR U4603 ( .A(n4791), .B(n4792), .Z(n4788) );
  AND U4604 ( .A(n138), .B(n4787), .Z(n4792) );
  XNOR U4605 ( .A(n4791), .B(n4785), .Z(n4787) );
  XOR U4606 ( .A(n4793), .B(n4794), .Z(n4785) );
  AND U4607 ( .A(n153), .B(n4795), .Z(n4794) );
  XNOR U4608 ( .A(n4796), .B(n4797), .Z(n4791) );
  AND U4609 ( .A(n145), .B(n4798), .Z(n4797) );
  XOR U4610 ( .A(p_input[175]), .B(n4796), .Z(n4798) );
  XNOR U4611 ( .A(n4799), .B(n4800), .Z(n4796) );
  AND U4612 ( .A(n149), .B(n4795), .Z(n4800) );
  XNOR U4613 ( .A(n4799), .B(n4793), .Z(n4795) );
  XOR U4614 ( .A(n4801), .B(n4802), .Z(n4793) );
  AND U4615 ( .A(n164), .B(n4803), .Z(n4802) );
  XNOR U4616 ( .A(n4804), .B(n4805), .Z(n4799) );
  AND U4617 ( .A(n156), .B(n4806), .Z(n4805) );
  XOR U4618 ( .A(p_input[191]), .B(n4804), .Z(n4806) );
  XNOR U4619 ( .A(n4807), .B(n4808), .Z(n4804) );
  AND U4620 ( .A(n160), .B(n4803), .Z(n4808) );
  XNOR U4621 ( .A(n4807), .B(n4801), .Z(n4803) );
  XOR U4622 ( .A(n4809), .B(n4810), .Z(n4801) );
  AND U4623 ( .A(n175), .B(n4811), .Z(n4810) );
  XNOR U4624 ( .A(n4812), .B(n4813), .Z(n4807) );
  AND U4625 ( .A(n167), .B(n4814), .Z(n4813) );
  XOR U4626 ( .A(p_input[207]), .B(n4812), .Z(n4814) );
  XNOR U4627 ( .A(n4815), .B(n4816), .Z(n4812) );
  AND U4628 ( .A(n171), .B(n4811), .Z(n4816) );
  XNOR U4629 ( .A(n4815), .B(n4809), .Z(n4811) );
  XOR U4630 ( .A(n4817), .B(n4818), .Z(n4809) );
  AND U4631 ( .A(n186), .B(n4819), .Z(n4818) );
  XNOR U4632 ( .A(n4820), .B(n4821), .Z(n4815) );
  AND U4633 ( .A(n178), .B(n4822), .Z(n4821) );
  XOR U4634 ( .A(p_input[223]), .B(n4820), .Z(n4822) );
  XNOR U4635 ( .A(n4823), .B(n4824), .Z(n4820) );
  AND U4636 ( .A(n182), .B(n4819), .Z(n4824) );
  XNOR U4637 ( .A(n4823), .B(n4817), .Z(n4819) );
  XOR U4638 ( .A(n4825), .B(n4826), .Z(n4817) );
  AND U4639 ( .A(n197), .B(n4827), .Z(n4826) );
  XNOR U4640 ( .A(n4828), .B(n4829), .Z(n4823) );
  AND U4641 ( .A(n189), .B(n4830), .Z(n4829) );
  XOR U4642 ( .A(p_input[239]), .B(n4828), .Z(n4830) );
  XNOR U4643 ( .A(n4831), .B(n4832), .Z(n4828) );
  AND U4644 ( .A(n193), .B(n4827), .Z(n4832) );
  XNOR U4645 ( .A(n4831), .B(n4825), .Z(n4827) );
  XOR U4646 ( .A(n4833), .B(n4834), .Z(n4825) );
  AND U4647 ( .A(n208), .B(n4835), .Z(n4834) );
  XNOR U4648 ( .A(n4836), .B(n4837), .Z(n4831) );
  AND U4649 ( .A(n200), .B(n4838), .Z(n4837) );
  XOR U4650 ( .A(p_input[255]), .B(n4836), .Z(n4838) );
  XNOR U4651 ( .A(n4839), .B(n4840), .Z(n4836) );
  AND U4652 ( .A(n204), .B(n4835), .Z(n4840) );
  XNOR U4653 ( .A(n4839), .B(n4833), .Z(n4835) );
  XOR U4654 ( .A(n4841), .B(n4842), .Z(n4833) );
  AND U4655 ( .A(n219), .B(n4843), .Z(n4842) );
  XNOR U4656 ( .A(n4844), .B(n4845), .Z(n4839) );
  AND U4657 ( .A(n211), .B(n4846), .Z(n4845) );
  XOR U4658 ( .A(p_input[271]), .B(n4844), .Z(n4846) );
  XNOR U4659 ( .A(n4847), .B(n4848), .Z(n4844) );
  AND U4660 ( .A(n215), .B(n4843), .Z(n4848) );
  XNOR U4661 ( .A(n4847), .B(n4841), .Z(n4843) );
  XOR U4662 ( .A(n4849), .B(n4850), .Z(n4841) );
  AND U4663 ( .A(n230), .B(n4851), .Z(n4850) );
  XNOR U4664 ( .A(n4852), .B(n4853), .Z(n4847) );
  AND U4665 ( .A(n222), .B(n4854), .Z(n4853) );
  XOR U4666 ( .A(p_input[287]), .B(n4852), .Z(n4854) );
  XNOR U4667 ( .A(n4855), .B(n4856), .Z(n4852) );
  AND U4668 ( .A(n226), .B(n4851), .Z(n4856) );
  XNOR U4669 ( .A(n4855), .B(n4849), .Z(n4851) );
  XOR U4670 ( .A(n4857), .B(n4858), .Z(n4849) );
  AND U4671 ( .A(n241), .B(n4859), .Z(n4858) );
  XNOR U4672 ( .A(n4860), .B(n4861), .Z(n4855) );
  AND U4673 ( .A(n233), .B(n4862), .Z(n4861) );
  XOR U4674 ( .A(p_input[303]), .B(n4860), .Z(n4862) );
  XNOR U4675 ( .A(n4863), .B(n4864), .Z(n4860) );
  AND U4676 ( .A(n237), .B(n4859), .Z(n4864) );
  XNOR U4677 ( .A(n4863), .B(n4857), .Z(n4859) );
  XOR U4678 ( .A(n4865), .B(n4866), .Z(n4857) );
  AND U4679 ( .A(n252), .B(n4867), .Z(n4866) );
  XNOR U4680 ( .A(n4868), .B(n4869), .Z(n4863) );
  AND U4681 ( .A(n244), .B(n4870), .Z(n4869) );
  XOR U4682 ( .A(p_input[319]), .B(n4868), .Z(n4870) );
  XNOR U4683 ( .A(n4871), .B(n4872), .Z(n4868) );
  AND U4684 ( .A(n248), .B(n4867), .Z(n4872) );
  XNOR U4685 ( .A(n4871), .B(n4865), .Z(n4867) );
  XOR U4686 ( .A(n4873), .B(n4874), .Z(n4865) );
  AND U4687 ( .A(n263), .B(n4875), .Z(n4874) );
  XNOR U4688 ( .A(n4876), .B(n4877), .Z(n4871) );
  AND U4689 ( .A(n255), .B(n4878), .Z(n4877) );
  XOR U4690 ( .A(p_input[335]), .B(n4876), .Z(n4878) );
  XNOR U4691 ( .A(n4879), .B(n4880), .Z(n4876) );
  AND U4692 ( .A(n259), .B(n4875), .Z(n4880) );
  XNOR U4693 ( .A(n4879), .B(n4873), .Z(n4875) );
  XOR U4694 ( .A(n4881), .B(n4882), .Z(n4873) );
  AND U4695 ( .A(n274), .B(n4883), .Z(n4882) );
  XNOR U4696 ( .A(n4884), .B(n4885), .Z(n4879) );
  AND U4697 ( .A(n266), .B(n4886), .Z(n4885) );
  XOR U4698 ( .A(p_input[351]), .B(n4884), .Z(n4886) );
  XNOR U4699 ( .A(n4887), .B(n4888), .Z(n4884) );
  AND U4700 ( .A(n270), .B(n4883), .Z(n4888) );
  XNOR U4701 ( .A(n4887), .B(n4881), .Z(n4883) );
  XOR U4702 ( .A(n4889), .B(n4890), .Z(n4881) );
  AND U4703 ( .A(n285), .B(n4891), .Z(n4890) );
  XNOR U4704 ( .A(n4892), .B(n4893), .Z(n4887) );
  AND U4705 ( .A(n277), .B(n4894), .Z(n4893) );
  XOR U4706 ( .A(p_input[367]), .B(n4892), .Z(n4894) );
  XNOR U4707 ( .A(n4895), .B(n4896), .Z(n4892) );
  AND U4708 ( .A(n281), .B(n4891), .Z(n4896) );
  XNOR U4709 ( .A(n4895), .B(n4889), .Z(n4891) );
  XOR U4710 ( .A(n4897), .B(n4898), .Z(n4889) );
  AND U4711 ( .A(n296), .B(n4899), .Z(n4898) );
  XNOR U4712 ( .A(n4900), .B(n4901), .Z(n4895) );
  AND U4713 ( .A(n288), .B(n4902), .Z(n4901) );
  XOR U4714 ( .A(p_input[383]), .B(n4900), .Z(n4902) );
  XNOR U4715 ( .A(n4903), .B(n4904), .Z(n4900) );
  AND U4716 ( .A(n292), .B(n4899), .Z(n4904) );
  XNOR U4717 ( .A(n4903), .B(n4897), .Z(n4899) );
  XOR U4718 ( .A(n4905), .B(n4906), .Z(n4897) );
  AND U4719 ( .A(n307), .B(n4907), .Z(n4906) );
  XNOR U4720 ( .A(n4908), .B(n4909), .Z(n4903) );
  AND U4721 ( .A(n299), .B(n4910), .Z(n4909) );
  XOR U4722 ( .A(p_input[399]), .B(n4908), .Z(n4910) );
  XNOR U4723 ( .A(n4911), .B(n4912), .Z(n4908) );
  AND U4724 ( .A(n303), .B(n4907), .Z(n4912) );
  XNOR U4725 ( .A(n4911), .B(n4905), .Z(n4907) );
  XOR U4726 ( .A(n4913), .B(n4914), .Z(n4905) );
  AND U4727 ( .A(n318), .B(n4915), .Z(n4914) );
  XNOR U4728 ( .A(n4916), .B(n4917), .Z(n4911) );
  AND U4729 ( .A(n310), .B(n4918), .Z(n4917) );
  XOR U4730 ( .A(p_input[415]), .B(n4916), .Z(n4918) );
  XNOR U4731 ( .A(n4919), .B(n4920), .Z(n4916) );
  AND U4732 ( .A(n314), .B(n4915), .Z(n4920) );
  XNOR U4733 ( .A(n4919), .B(n4913), .Z(n4915) );
  XOR U4734 ( .A(n4921), .B(n4922), .Z(n4913) );
  AND U4735 ( .A(n329), .B(n4923), .Z(n4922) );
  XNOR U4736 ( .A(n4924), .B(n4925), .Z(n4919) );
  AND U4737 ( .A(n321), .B(n4926), .Z(n4925) );
  XOR U4738 ( .A(p_input[431]), .B(n4924), .Z(n4926) );
  XNOR U4739 ( .A(n4927), .B(n4928), .Z(n4924) );
  AND U4740 ( .A(n325), .B(n4923), .Z(n4928) );
  XNOR U4741 ( .A(n4927), .B(n4921), .Z(n4923) );
  XOR U4742 ( .A(n4929), .B(n4930), .Z(n4921) );
  AND U4743 ( .A(n340), .B(n4931), .Z(n4930) );
  XNOR U4744 ( .A(n4932), .B(n4933), .Z(n4927) );
  AND U4745 ( .A(n332), .B(n4934), .Z(n4933) );
  XOR U4746 ( .A(p_input[447]), .B(n4932), .Z(n4934) );
  XNOR U4747 ( .A(n4935), .B(n4936), .Z(n4932) );
  AND U4748 ( .A(n336), .B(n4931), .Z(n4936) );
  XNOR U4749 ( .A(n4935), .B(n4929), .Z(n4931) );
  XOR U4750 ( .A(n4937), .B(n4938), .Z(n4929) );
  AND U4751 ( .A(n351), .B(n4939), .Z(n4938) );
  XNOR U4752 ( .A(n4940), .B(n4941), .Z(n4935) );
  AND U4753 ( .A(n343), .B(n4942), .Z(n4941) );
  XOR U4754 ( .A(p_input[463]), .B(n4940), .Z(n4942) );
  XNOR U4755 ( .A(n4943), .B(n4944), .Z(n4940) );
  AND U4756 ( .A(n347), .B(n4939), .Z(n4944) );
  XNOR U4757 ( .A(n4943), .B(n4937), .Z(n4939) );
  XOR U4758 ( .A(n4945), .B(n4946), .Z(n4937) );
  AND U4759 ( .A(n362), .B(n4947), .Z(n4946) );
  XNOR U4760 ( .A(n4948), .B(n4949), .Z(n4943) );
  AND U4761 ( .A(n354), .B(n4950), .Z(n4949) );
  XOR U4762 ( .A(p_input[479]), .B(n4948), .Z(n4950) );
  XNOR U4763 ( .A(n4951), .B(n4952), .Z(n4948) );
  AND U4764 ( .A(n358), .B(n4947), .Z(n4952) );
  XNOR U4765 ( .A(n4951), .B(n4945), .Z(n4947) );
  XOR U4766 ( .A(n4953), .B(n4954), .Z(n4945) );
  AND U4767 ( .A(n373), .B(n4955), .Z(n4954) );
  XNOR U4768 ( .A(n4956), .B(n4957), .Z(n4951) );
  AND U4769 ( .A(n365), .B(n4958), .Z(n4957) );
  XOR U4770 ( .A(p_input[495]), .B(n4956), .Z(n4958) );
  XNOR U4771 ( .A(n4959), .B(n4960), .Z(n4956) );
  AND U4772 ( .A(n369), .B(n4955), .Z(n4960) );
  XNOR U4773 ( .A(n4959), .B(n4953), .Z(n4955) );
  XOR U4774 ( .A(n4961), .B(n4962), .Z(n4953) );
  AND U4775 ( .A(n384), .B(n4963), .Z(n4962) );
  XNOR U4776 ( .A(n4964), .B(n4965), .Z(n4959) );
  AND U4777 ( .A(n376), .B(n4966), .Z(n4965) );
  XOR U4778 ( .A(p_input[511]), .B(n4964), .Z(n4966) );
  XNOR U4779 ( .A(n4967), .B(n4968), .Z(n4964) );
  AND U4780 ( .A(n380), .B(n4963), .Z(n4968) );
  XNOR U4781 ( .A(n4967), .B(n4961), .Z(n4963) );
  XOR U4782 ( .A(n4969), .B(n4970), .Z(n4961) );
  AND U4783 ( .A(n395), .B(n4971), .Z(n4970) );
  XNOR U4784 ( .A(n4972), .B(n4973), .Z(n4967) );
  AND U4785 ( .A(n387), .B(n4974), .Z(n4973) );
  XOR U4786 ( .A(p_input[527]), .B(n4972), .Z(n4974) );
  XNOR U4787 ( .A(n4975), .B(n4976), .Z(n4972) );
  AND U4788 ( .A(n391), .B(n4971), .Z(n4976) );
  XNOR U4789 ( .A(n4975), .B(n4969), .Z(n4971) );
  XOR U4790 ( .A(n4977), .B(n4978), .Z(n4969) );
  AND U4791 ( .A(n406), .B(n4979), .Z(n4978) );
  XNOR U4792 ( .A(n4980), .B(n4981), .Z(n4975) );
  AND U4793 ( .A(n398), .B(n4982), .Z(n4981) );
  XOR U4794 ( .A(p_input[543]), .B(n4980), .Z(n4982) );
  XNOR U4795 ( .A(n4983), .B(n4984), .Z(n4980) );
  AND U4796 ( .A(n402), .B(n4979), .Z(n4984) );
  XNOR U4797 ( .A(n4983), .B(n4977), .Z(n4979) );
  XOR U4798 ( .A(n4985), .B(n4986), .Z(n4977) );
  AND U4799 ( .A(n417), .B(n4987), .Z(n4986) );
  XNOR U4800 ( .A(n4988), .B(n4989), .Z(n4983) );
  AND U4801 ( .A(n409), .B(n4990), .Z(n4989) );
  XOR U4802 ( .A(p_input[559]), .B(n4988), .Z(n4990) );
  XNOR U4803 ( .A(n4991), .B(n4992), .Z(n4988) );
  AND U4804 ( .A(n413), .B(n4987), .Z(n4992) );
  XNOR U4805 ( .A(n4991), .B(n4985), .Z(n4987) );
  XOR U4806 ( .A(n4993), .B(n4994), .Z(n4985) );
  AND U4807 ( .A(n428), .B(n4995), .Z(n4994) );
  XNOR U4808 ( .A(n4996), .B(n4997), .Z(n4991) );
  AND U4809 ( .A(n420), .B(n4998), .Z(n4997) );
  XOR U4810 ( .A(p_input[575]), .B(n4996), .Z(n4998) );
  XNOR U4811 ( .A(n4999), .B(n5000), .Z(n4996) );
  AND U4812 ( .A(n424), .B(n4995), .Z(n5000) );
  XNOR U4813 ( .A(n4999), .B(n4993), .Z(n4995) );
  XOR U4814 ( .A(n5001), .B(n5002), .Z(n4993) );
  AND U4815 ( .A(n439), .B(n5003), .Z(n5002) );
  XNOR U4816 ( .A(n5004), .B(n5005), .Z(n4999) );
  AND U4817 ( .A(n431), .B(n5006), .Z(n5005) );
  XOR U4818 ( .A(p_input[591]), .B(n5004), .Z(n5006) );
  XNOR U4819 ( .A(n5007), .B(n5008), .Z(n5004) );
  AND U4820 ( .A(n435), .B(n5003), .Z(n5008) );
  XNOR U4821 ( .A(n5007), .B(n5001), .Z(n5003) );
  XOR U4822 ( .A(n5009), .B(n5010), .Z(n5001) );
  AND U4823 ( .A(n450), .B(n5011), .Z(n5010) );
  XNOR U4824 ( .A(n5012), .B(n5013), .Z(n5007) );
  AND U4825 ( .A(n442), .B(n5014), .Z(n5013) );
  XOR U4826 ( .A(p_input[607]), .B(n5012), .Z(n5014) );
  XNOR U4827 ( .A(n5015), .B(n5016), .Z(n5012) );
  AND U4828 ( .A(n446), .B(n5011), .Z(n5016) );
  XNOR U4829 ( .A(n5015), .B(n5009), .Z(n5011) );
  XOR U4830 ( .A(n5017), .B(n5018), .Z(n5009) );
  AND U4831 ( .A(n461), .B(n5019), .Z(n5018) );
  XNOR U4832 ( .A(n5020), .B(n5021), .Z(n5015) );
  AND U4833 ( .A(n453), .B(n5022), .Z(n5021) );
  XOR U4834 ( .A(p_input[623]), .B(n5020), .Z(n5022) );
  XNOR U4835 ( .A(n5023), .B(n5024), .Z(n5020) );
  AND U4836 ( .A(n457), .B(n5019), .Z(n5024) );
  XNOR U4837 ( .A(n5023), .B(n5017), .Z(n5019) );
  XOR U4838 ( .A(n5025), .B(n5026), .Z(n5017) );
  AND U4839 ( .A(n472), .B(n5027), .Z(n5026) );
  XNOR U4840 ( .A(n5028), .B(n5029), .Z(n5023) );
  AND U4841 ( .A(n464), .B(n5030), .Z(n5029) );
  XOR U4842 ( .A(p_input[639]), .B(n5028), .Z(n5030) );
  XNOR U4843 ( .A(n5031), .B(n5032), .Z(n5028) );
  AND U4844 ( .A(n468), .B(n5027), .Z(n5032) );
  XNOR U4845 ( .A(n5031), .B(n5025), .Z(n5027) );
  XOR U4846 ( .A(n5033), .B(n5034), .Z(n5025) );
  AND U4847 ( .A(n483), .B(n5035), .Z(n5034) );
  XNOR U4848 ( .A(n5036), .B(n5037), .Z(n5031) );
  AND U4849 ( .A(n475), .B(n5038), .Z(n5037) );
  XOR U4850 ( .A(p_input[655]), .B(n5036), .Z(n5038) );
  XNOR U4851 ( .A(n5039), .B(n5040), .Z(n5036) );
  AND U4852 ( .A(n479), .B(n5035), .Z(n5040) );
  XNOR U4853 ( .A(n5039), .B(n5033), .Z(n5035) );
  XOR U4854 ( .A(n5041), .B(n5042), .Z(n5033) );
  AND U4855 ( .A(n494), .B(n5043), .Z(n5042) );
  XNOR U4856 ( .A(n5044), .B(n5045), .Z(n5039) );
  AND U4857 ( .A(n486), .B(n5046), .Z(n5045) );
  XOR U4858 ( .A(p_input[671]), .B(n5044), .Z(n5046) );
  XNOR U4859 ( .A(n5047), .B(n5048), .Z(n5044) );
  AND U4860 ( .A(n490), .B(n5043), .Z(n5048) );
  XNOR U4861 ( .A(n5047), .B(n5041), .Z(n5043) );
  XOR U4862 ( .A(n5049), .B(n5050), .Z(n5041) );
  AND U4863 ( .A(n505), .B(n5051), .Z(n5050) );
  XNOR U4864 ( .A(n5052), .B(n5053), .Z(n5047) );
  AND U4865 ( .A(n497), .B(n5054), .Z(n5053) );
  XOR U4866 ( .A(p_input[687]), .B(n5052), .Z(n5054) );
  XNOR U4867 ( .A(n5055), .B(n5056), .Z(n5052) );
  AND U4868 ( .A(n501), .B(n5051), .Z(n5056) );
  XNOR U4869 ( .A(n5055), .B(n5049), .Z(n5051) );
  XOR U4870 ( .A(n5057), .B(n5058), .Z(n5049) );
  AND U4871 ( .A(n516), .B(n5059), .Z(n5058) );
  XNOR U4872 ( .A(n5060), .B(n5061), .Z(n5055) );
  AND U4873 ( .A(n508), .B(n5062), .Z(n5061) );
  XOR U4874 ( .A(p_input[703]), .B(n5060), .Z(n5062) );
  XNOR U4875 ( .A(n5063), .B(n5064), .Z(n5060) );
  AND U4876 ( .A(n512), .B(n5059), .Z(n5064) );
  XNOR U4877 ( .A(n5063), .B(n5057), .Z(n5059) );
  XOR U4878 ( .A(n5065), .B(n5066), .Z(n5057) );
  AND U4879 ( .A(n527), .B(n5067), .Z(n5066) );
  XNOR U4880 ( .A(n5068), .B(n5069), .Z(n5063) );
  AND U4881 ( .A(n519), .B(n5070), .Z(n5069) );
  XOR U4882 ( .A(p_input[719]), .B(n5068), .Z(n5070) );
  XNOR U4883 ( .A(n5071), .B(n5072), .Z(n5068) );
  AND U4884 ( .A(n523), .B(n5067), .Z(n5072) );
  XNOR U4885 ( .A(n5071), .B(n5065), .Z(n5067) );
  XOR U4886 ( .A(n5073), .B(n5074), .Z(n5065) );
  AND U4887 ( .A(n538), .B(n5075), .Z(n5074) );
  XNOR U4888 ( .A(n5076), .B(n5077), .Z(n5071) );
  AND U4889 ( .A(n530), .B(n5078), .Z(n5077) );
  XOR U4890 ( .A(p_input[735]), .B(n5076), .Z(n5078) );
  XNOR U4891 ( .A(n5079), .B(n5080), .Z(n5076) );
  AND U4892 ( .A(n534), .B(n5075), .Z(n5080) );
  XNOR U4893 ( .A(n5079), .B(n5073), .Z(n5075) );
  XOR U4894 ( .A(n5081), .B(n5082), .Z(n5073) );
  AND U4895 ( .A(n549), .B(n5083), .Z(n5082) );
  XNOR U4896 ( .A(n5084), .B(n5085), .Z(n5079) );
  AND U4897 ( .A(n541), .B(n5086), .Z(n5085) );
  XOR U4898 ( .A(p_input[751]), .B(n5084), .Z(n5086) );
  XNOR U4899 ( .A(n5087), .B(n5088), .Z(n5084) );
  AND U4900 ( .A(n545), .B(n5083), .Z(n5088) );
  XNOR U4901 ( .A(n5087), .B(n5081), .Z(n5083) );
  XOR U4902 ( .A(n5089), .B(n5090), .Z(n5081) );
  AND U4903 ( .A(n560), .B(n5091), .Z(n5090) );
  XNOR U4904 ( .A(n5092), .B(n5093), .Z(n5087) );
  AND U4905 ( .A(n552), .B(n5094), .Z(n5093) );
  XOR U4906 ( .A(p_input[767]), .B(n5092), .Z(n5094) );
  XNOR U4907 ( .A(n5095), .B(n5096), .Z(n5092) );
  AND U4908 ( .A(n556), .B(n5091), .Z(n5096) );
  XNOR U4909 ( .A(n5095), .B(n5089), .Z(n5091) );
  XOR U4910 ( .A(n5097), .B(n5098), .Z(n5089) );
  AND U4911 ( .A(n571), .B(n5099), .Z(n5098) );
  XNOR U4912 ( .A(n5100), .B(n5101), .Z(n5095) );
  AND U4913 ( .A(n563), .B(n5102), .Z(n5101) );
  XOR U4914 ( .A(p_input[783]), .B(n5100), .Z(n5102) );
  XNOR U4915 ( .A(n5103), .B(n5104), .Z(n5100) );
  AND U4916 ( .A(n567), .B(n5099), .Z(n5104) );
  XNOR U4917 ( .A(n5103), .B(n5097), .Z(n5099) );
  XOR U4918 ( .A(n5105), .B(n5106), .Z(n5097) );
  AND U4919 ( .A(n582), .B(n5107), .Z(n5106) );
  XNOR U4920 ( .A(n5108), .B(n5109), .Z(n5103) );
  AND U4921 ( .A(n574), .B(n5110), .Z(n5109) );
  XOR U4922 ( .A(p_input[799]), .B(n5108), .Z(n5110) );
  XNOR U4923 ( .A(n5111), .B(n5112), .Z(n5108) );
  AND U4924 ( .A(n578), .B(n5107), .Z(n5112) );
  XNOR U4925 ( .A(n5111), .B(n5105), .Z(n5107) );
  XOR U4926 ( .A(n5113), .B(n5114), .Z(n5105) );
  AND U4927 ( .A(n593), .B(n5115), .Z(n5114) );
  XNOR U4928 ( .A(n5116), .B(n5117), .Z(n5111) );
  AND U4929 ( .A(n585), .B(n5118), .Z(n5117) );
  XOR U4930 ( .A(p_input[815]), .B(n5116), .Z(n5118) );
  XNOR U4931 ( .A(n5119), .B(n5120), .Z(n5116) );
  AND U4932 ( .A(n589), .B(n5115), .Z(n5120) );
  XNOR U4933 ( .A(n5119), .B(n5113), .Z(n5115) );
  XOR U4934 ( .A(n5121), .B(n5122), .Z(n5113) );
  AND U4935 ( .A(n604), .B(n5123), .Z(n5122) );
  XNOR U4936 ( .A(n5124), .B(n5125), .Z(n5119) );
  AND U4937 ( .A(n596), .B(n5126), .Z(n5125) );
  XOR U4938 ( .A(p_input[831]), .B(n5124), .Z(n5126) );
  XNOR U4939 ( .A(n5127), .B(n5128), .Z(n5124) );
  AND U4940 ( .A(n600), .B(n5123), .Z(n5128) );
  XNOR U4941 ( .A(n5127), .B(n5121), .Z(n5123) );
  XOR U4942 ( .A(n5129), .B(n5130), .Z(n5121) );
  AND U4943 ( .A(n615), .B(n5131), .Z(n5130) );
  XNOR U4944 ( .A(n5132), .B(n5133), .Z(n5127) );
  AND U4945 ( .A(n607), .B(n5134), .Z(n5133) );
  XOR U4946 ( .A(p_input[847]), .B(n5132), .Z(n5134) );
  XNOR U4947 ( .A(n5135), .B(n5136), .Z(n5132) );
  AND U4948 ( .A(n611), .B(n5131), .Z(n5136) );
  XNOR U4949 ( .A(n5135), .B(n5129), .Z(n5131) );
  XOR U4950 ( .A(n5137), .B(n5138), .Z(n5129) );
  AND U4951 ( .A(n626), .B(n5139), .Z(n5138) );
  XNOR U4952 ( .A(n5140), .B(n5141), .Z(n5135) );
  AND U4953 ( .A(n618), .B(n5142), .Z(n5141) );
  XOR U4954 ( .A(p_input[863]), .B(n5140), .Z(n5142) );
  XNOR U4955 ( .A(n5143), .B(n5144), .Z(n5140) );
  AND U4956 ( .A(n622), .B(n5139), .Z(n5144) );
  XNOR U4957 ( .A(n5143), .B(n5137), .Z(n5139) );
  XOR U4958 ( .A(n5145), .B(n5146), .Z(n5137) );
  AND U4959 ( .A(n637), .B(n5147), .Z(n5146) );
  XNOR U4960 ( .A(n5148), .B(n5149), .Z(n5143) );
  AND U4961 ( .A(n629), .B(n5150), .Z(n5149) );
  XOR U4962 ( .A(p_input[879]), .B(n5148), .Z(n5150) );
  XNOR U4963 ( .A(n5151), .B(n5152), .Z(n5148) );
  AND U4964 ( .A(n633), .B(n5147), .Z(n5152) );
  XNOR U4965 ( .A(n5151), .B(n5145), .Z(n5147) );
  XOR U4966 ( .A(n5153), .B(n5154), .Z(n5145) );
  AND U4967 ( .A(n648), .B(n5155), .Z(n5154) );
  XNOR U4968 ( .A(n5156), .B(n5157), .Z(n5151) );
  AND U4969 ( .A(n640), .B(n5158), .Z(n5157) );
  XOR U4970 ( .A(p_input[895]), .B(n5156), .Z(n5158) );
  XNOR U4971 ( .A(n5159), .B(n5160), .Z(n5156) );
  AND U4972 ( .A(n644), .B(n5155), .Z(n5160) );
  XNOR U4973 ( .A(n5159), .B(n5153), .Z(n5155) );
  XOR U4974 ( .A(n5161), .B(n5162), .Z(n5153) );
  AND U4975 ( .A(n659), .B(n5163), .Z(n5162) );
  XNOR U4976 ( .A(n5164), .B(n5165), .Z(n5159) );
  AND U4977 ( .A(n651), .B(n5166), .Z(n5165) );
  XOR U4978 ( .A(p_input[911]), .B(n5164), .Z(n5166) );
  XNOR U4979 ( .A(n5167), .B(n5168), .Z(n5164) );
  AND U4980 ( .A(n655), .B(n5163), .Z(n5168) );
  XNOR U4981 ( .A(n5167), .B(n5161), .Z(n5163) );
  XOR U4982 ( .A(n5169), .B(n5170), .Z(n5161) );
  AND U4983 ( .A(n670), .B(n5171), .Z(n5170) );
  XNOR U4984 ( .A(n5172), .B(n5173), .Z(n5167) );
  AND U4985 ( .A(n662), .B(n5174), .Z(n5173) );
  XOR U4986 ( .A(p_input[927]), .B(n5172), .Z(n5174) );
  XNOR U4987 ( .A(n5175), .B(n5176), .Z(n5172) );
  AND U4988 ( .A(n666), .B(n5171), .Z(n5176) );
  XNOR U4989 ( .A(n5175), .B(n5169), .Z(n5171) );
  XOR U4990 ( .A(n5177), .B(n5178), .Z(n5169) );
  AND U4991 ( .A(n681), .B(n5179), .Z(n5178) );
  XNOR U4992 ( .A(n5180), .B(n5181), .Z(n5175) );
  AND U4993 ( .A(n673), .B(n5182), .Z(n5181) );
  XOR U4994 ( .A(p_input[943]), .B(n5180), .Z(n5182) );
  XNOR U4995 ( .A(n5183), .B(n5184), .Z(n5180) );
  AND U4996 ( .A(n677), .B(n5179), .Z(n5184) );
  XNOR U4997 ( .A(n5183), .B(n5177), .Z(n5179) );
  XOR U4998 ( .A(n5185), .B(n5186), .Z(n5177) );
  AND U4999 ( .A(n692), .B(n5187), .Z(n5186) );
  XNOR U5000 ( .A(n5188), .B(n5189), .Z(n5183) );
  AND U5001 ( .A(n684), .B(n5190), .Z(n5189) );
  XOR U5002 ( .A(p_input[959]), .B(n5188), .Z(n5190) );
  XNOR U5003 ( .A(n5191), .B(n5192), .Z(n5188) );
  AND U5004 ( .A(n688), .B(n5187), .Z(n5192) );
  XNOR U5005 ( .A(n5191), .B(n5185), .Z(n5187) );
  XOR U5006 ( .A(n5193), .B(n5194), .Z(n5185) );
  AND U5007 ( .A(n703), .B(n5195), .Z(n5194) );
  XNOR U5008 ( .A(n5196), .B(n5197), .Z(n5191) );
  AND U5009 ( .A(n695), .B(n5198), .Z(n5197) );
  XOR U5010 ( .A(p_input[975]), .B(n5196), .Z(n5198) );
  XNOR U5011 ( .A(n5199), .B(n5200), .Z(n5196) );
  AND U5012 ( .A(n699), .B(n5195), .Z(n5200) );
  XNOR U5013 ( .A(n5199), .B(n5193), .Z(n5195) );
  XOR U5014 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n5201), .Z(n5193) );
  AND U5015 ( .A(n713), .B(n5202), .Z(n5201) );
  XNOR U5016 ( .A(n5203), .B(n5204), .Z(n5199) );
  AND U5017 ( .A(n706), .B(n5205), .Z(n5204) );
  XOR U5018 ( .A(p_input[991]), .B(n5203), .Z(n5205) );
  XNOR U5019 ( .A(n5206), .B(n5207), .Z(n5203) );
  AND U5020 ( .A(n710), .B(n5202), .Z(n5207) );
  XOR U5021 ( .A(n5208), .B(n5206), .Z(n5202) );
  IV U5022 ( .A(\knn_comb_/min_val_out[0][15] ), .Z(n5208) );
  XOR U5023 ( .A(n17), .B(n5209), .Z(o[14]) );
  AND U5024 ( .A(n30), .B(n5210), .Z(n17) );
  XOR U5025 ( .A(n18), .B(n5209), .Z(n5210) );
  XOR U5026 ( .A(n5211), .B(n5212), .Z(n5209) );
  AND U5027 ( .A(n42), .B(n5213), .Z(n5212) );
  XOR U5028 ( .A(n5214), .B(n5215), .Z(n18) );
  AND U5029 ( .A(n34), .B(n5216), .Z(n5215) );
  XOR U5030 ( .A(p_input[14]), .B(n5214), .Z(n5216) );
  XNOR U5031 ( .A(n5217), .B(n5218), .Z(n5214) );
  AND U5032 ( .A(n38), .B(n5213), .Z(n5218) );
  XNOR U5033 ( .A(n5217), .B(n5211), .Z(n5213) );
  XOR U5034 ( .A(n5219), .B(n5220), .Z(n5211) );
  AND U5035 ( .A(n54), .B(n5221), .Z(n5220) );
  XNOR U5036 ( .A(n5222), .B(n5223), .Z(n5217) );
  AND U5037 ( .A(n46), .B(n5224), .Z(n5223) );
  XOR U5038 ( .A(p_input[30]), .B(n5222), .Z(n5224) );
  XNOR U5039 ( .A(n5225), .B(n5226), .Z(n5222) );
  AND U5040 ( .A(n50), .B(n5221), .Z(n5226) );
  XNOR U5041 ( .A(n5225), .B(n5219), .Z(n5221) );
  XOR U5042 ( .A(n5227), .B(n5228), .Z(n5219) );
  AND U5043 ( .A(n65), .B(n5229), .Z(n5228) );
  XNOR U5044 ( .A(n5230), .B(n5231), .Z(n5225) );
  AND U5045 ( .A(n57), .B(n5232), .Z(n5231) );
  XOR U5046 ( .A(p_input[46]), .B(n5230), .Z(n5232) );
  XNOR U5047 ( .A(n5233), .B(n5234), .Z(n5230) );
  AND U5048 ( .A(n61), .B(n5229), .Z(n5234) );
  XNOR U5049 ( .A(n5233), .B(n5227), .Z(n5229) );
  XOR U5050 ( .A(n5235), .B(n5236), .Z(n5227) );
  AND U5051 ( .A(n76), .B(n5237), .Z(n5236) );
  XNOR U5052 ( .A(n5238), .B(n5239), .Z(n5233) );
  AND U5053 ( .A(n68), .B(n5240), .Z(n5239) );
  XOR U5054 ( .A(p_input[62]), .B(n5238), .Z(n5240) );
  XNOR U5055 ( .A(n5241), .B(n5242), .Z(n5238) );
  AND U5056 ( .A(n72), .B(n5237), .Z(n5242) );
  XNOR U5057 ( .A(n5241), .B(n5235), .Z(n5237) );
  XOR U5058 ( .A(n5243), .B(n5244), .Z(n5235) );
  AND U5059 ( .A(n87), .B(n5245), .Z(n5244) );
  XNOR U5060 ( .A(n5246), .B(n5247), .Z(n5241) );
  AND U5061 ( .A(n79), .B(n5248), .Z(n5247) );
  XOR U5062 ( .A(p_input[78]), .B(n5246), .Z(n5248) );
  XNOR U5063 ( .A(n5249), .B(n5250), .Z(n5246) );
  AND U5064 ( .A(n83), .B(n5245), .Z(n5250) );
  XNOR U5065 ( .A(n5249), .B(n5243), .Z(n5245) );
  XOR U5066 ( .A(n5251), .B(n5252), .Z(n5243) );
  AND U5067 ( .A(n98), .B(n5253), .Z(n5252) );
  XNOR U5068 ( .A(n5254), .B(n5255), .Z(n5249) );
  AND U5069 ( .A(n90), .B(n5256), .Z(n5255) );
  XOR U5070 ( .A(p_input[94]), .B(n5254), .Z(n5256) );
  XNOR U5071 ( .A(n5257), .B(n5258), .Z(n5254) );
  AND U5072 ( .A(n94), .B(n5253), .Z(n5258) );
  XNOR U5073 ( .A(n5257), .B(n5251), .Z(n5253) );
  XOR U5074 ( .A(n5259), .B(n5260), .Z(n5251) );
  AND U5075 ( .A(n109), .B(n5261), .Z(n5260) );
  XNOR U5076 ( .A(n5262), .B(n5263), .Z(n5257) );
  AND U5077 ( .A(n101), .B(n5264), .Z(n5263) );
  XOR U5078 ( .A(p_input[110]), .B(n5262), .Z(n5264) );
  XNOR U5079 ( .A(n5265), .B(n5266), .Z(n5262) );
  AND U5080 ( .A(n105), .B(n5261), .Z(n5266) );
  XNOR U5081 ( .A(n5265), .B(n5259), .Z(n5261) );
  XOR U5082 ( .A(n5267), .B(n5268), .Z(n5259) );
  AND U5083 ( .A(n120), .B(n5269), .Z(n5268) );
  XNOR U5084 ( .A(n5270), .B(n5271), .Z(n5265) );
  AND U5085 ( .A(n112), .B(n5272), .Z(n5271) );
  XOR U5086 ( .A(p_input[126]), .B(n5270), .Z(n5272) );
  XNOR U5087 ( .A(n5273), .B(n5274), .Z(n5270) );
  AND U5088 ( .A(n116), .B(n5269), .Z(n5274) );
  XNOR U5089 ( .A(n5273), .B(n5267), .Z(n5269) );
  XOR U5090 ( .A(n5275), .B(n5276), .Z(n5267) );
  AND U5091 ( .A(n131), .B(n5277), .Z(n5276) );
  XNOR U5092 ( .A(n5278), .B(n5279), .Z(n5273) );
  AND U5093 ( .A(n123), .B(n5280), .Z(n5279) );
  XOR U5094 ( .A(p_input[142]), .B(n5278), .Z(n5280) );
  XNOR U5095 ( .A(n5281), .B(n5282), .Z(n5278) );
  AND U5096 ( .A(n127), .B(n5277), .Z(n5282) );
  XNOR U5097 ( .A(n5281), .B(n5275), .Z(n5277) );
  XOR U5098 ( .A(n5283), .B(n5284), .Z(n5275) );
  AND U5099 ( .A(n142), .B(n5285), .Z(n5284) );
  XNOR U5100 ( .A(n5286), .B(n5287), .Z(n5281) );
  AND U5101 ( .A(n134), .B(n5288), .Z(n5287) );
  XOR U5102 ( .A(p_input[158]), .B(n5286), .Z(n5288) );
  XNOR U5103 ( .A(n5289), .B(n5290), .Z(n5286) );
  AND U5104 ( .A(n138), .B(n5285), .Z(n5290) );
  XNOR U5105 ( .A(n5289), .B(n5283), .Z(n5285) );
  XOR U5106 ( .A(n5291), .B(n5292), .Z(n5283) );
  AND U5107 ( .A(n153), .B(n5293), .Z(n5292) );
  XNOR U5108 ( .A(n5294), .B(n5295), .Z(n5289) );
  AND U5109 ( .A(n145), .B(n5296), .Z(n5295) );
  XOR U5110 ( .A(p_input[174]), .B(n5294), .Z(n5296) );
  XNOR U5111 ( .A(n5297), .B(n5298), .Z(n5294) );
  AND U5112 ( .A(n149), .B(n5293), .Z(n5298) );
  XNOR U5113 ( .A(n5297), .B(n5291), .Z(n5293) );
  XOR U5114 ( .A(n5299), .B(n5300), .Z(n5291) );
  AND U5115 ( .A(n164), .B(n5301), .Z(n5300) );
  XNOR U5116 ( .A(n5302), .B(n5303), .Z(n5297) );
  AND U5117 ( .A(n156), .B(n5304), .Z(n5303) );
  XOR U5118 ( .A(p_input[190]), .B(n5302), .Z(n5304) );
  XNOR U5119 ( .A(n5305), .B(n5306), .Z(n5302) );
  AND U5120 ( .A(n160), .B(n5301), .Z(n5306) );
  XNOR U5121 ( .A(n5305), .B(n5299), .Z(n5301) );
  XOR U5122 ( .A(n5307), .B(n5308), .Z(n5299) );
  AND U5123 ( .A(n175), .B(n5309), .Z(n5308) );
  XNOR U5124 ( .A(n5310), .B(n5311), .Z(n5305) );
  AND U5125 ( .A(n167), .B(n5312), .Z(n5311) );
  XOR U5126 ( .A(p_input[206]), .B(n5310), .Z(n5312) );
  XNOR U5127 ( .A(n5313), .B(n5314), .Z(n5310) );
  AND U5128 ( .A(n171), .B(n5309), .Z(n5314) );
  XNOR U5129 ( .A(n5313), .B(n5307), .Z(n5309) );
  XOR U5130 ( .A(n5315), .B(n5316), .Z(n5307) );
  AND U5131 ( .A(n186), .B(n5317), .Z(n5316) );
  XNOR U5132 ( .A(n5318), .B(n5319), .Z(n5313) );
  AND U5133 ( .A(n178), .B(n5320), .Z(n5319) );
  XOR U5134 ( .A(p_input[222]), .B(n5318), .Z(n5320) );
  XNOR U5135 ( .A(n5321), .B(n5322), .Z(n5318) );
  AND U5136 ( .A(n182), .B(n5317), .Z(n5322) );
  XNOR U5137 ( .A(n5321), .B(n5315), .Z(n5317) );
  XOR U5138 ( .A(n5323), .B(n5324), .Z(n5315) );
  AND U5139 ( .A(n197), .B(n5325), .Z(n5324) );
  XNOR U5140 ( .A(n5326), .B(n5327), .Z(n5321) );
  AND U5141 ( .A(n189), .B(n5328), .Z(n5327) );
  XOR U5142 ( .A(p_input[238]), .B(n5326), .Z(n5328) );
  XNOR U5143 ( .A(n5329), .B(n5330), .Z(n5326) );
  AND U5144 ( .A(n193), .B(n5325), .Z(n5330) );
  XNOR U5145 ( .A(n5329), .B(n5323), .Z(n5325) );
  XOR U5146 ( .A(n5331), .B(n5332), .Z(n5323) );
  AND U5147 ( .A(n208), .B(n5333), .Z(n5332) );
  XNOR U5148 ( .A(n5334), .B(n5335), .Z(n5329) );
  AND U5149 ( .A(n200), .B(n5336), .Z(n5335) );
  XOR U5150 ( .A(p_input[254]), .B(n5334), .Z(n5336) );
  XNOR U5151 ( .A(n5337), .B(n5338), .Z(n5334) );
  AND U5152 ( .A(n204), .B(n5333), .Z(n5338) );
  XNOR U5153 ( .A(n5337), .B(n5331), .Z(n5333) );
  XOR U5154 ( .A(n5339), .B(n5340), .Z(n5331) );
  AND U5155 ( .A(n219), .B(n5341), .Z(n5340) );
  XNOR U5156 ( .A(n5342), .B(n5343), .Z(n5337) );
  AND U5157 ( .A(n211), .B(n5344), .Z(n5343) );
  XOR U5158 ( .A(p_input[270]), .B(n5342), .Z(n5344) );
  XNOR U5159 ( .A(n5345), .B(n5346), .Z(n5342) );
  AND U5160 ( .A(n215), .B(n5341), .Z(n5346) );
  XNOR U5161 ( .A(n5345), .B(n5339), .Z(n5341) );
  XOR U5162 ( .A(n5347), .B(n5348), .Z(n5339) );
  AND U5163 ( .A(n230), .B(n5349), .Z(n5348) );
  XNOR U5164 ( .A(n5350), .B(n5351), .Z(n5345) );
  AND U5165 ( .A(n222), .B(n5352), .Z(n5351) );
  XOR U5166 ( .A(p_input[286]), .B(n5350), .Z(n5352) );
  XNOR U5167 ( .A(n5353), .B(n5354), .Z(n5350) );
  AND U5168 ( .A(n226), .B(n5349), .Z(n5354) );
  XNOR U5169 ( .A(n5353), .B(n5347), .Z(n5349) );
  XOR U5170 ( .A(n5355), .B(n5356), .Z(n5347) );
  AND U5171 ( .A(n241), .B(n5357), .Z(n5356) );
  XNOR U5172 ( .A(n5358), .B(n5359), .Z(n5353) );
  AND U5173 ( .A(n233), .B(n5360), .Z(n5359) );
  XOR U5174 ( .A(p_input[302]), .B(n5358), .Z(n5360) );
  XNOR U5175 ( .A(n5361), .B(n5362), .Z(n5358) );
  AND U5176 ( .A(n237), .B(n5357), .Z(n5362) );
  XNOR U5177 ( .A(n5361), .B(n5355), .Z(n5357) );
  XOR U5178 ( .A(n5363), .B(n5364), .Z(n5355) );
  AND U5179 ( .A(n252), .B(n5365), .Z(n5364) );
  XNOR U5180 ( .A(n5366), .B(n5367), .Z(n5361) );
  AND U5181 ( .A(n244), .B(n5368), .Z(n5367) );
  XOR U5182 ( .A(p_input[318]), .B(n5366), .Z(n5368) );
  XNOR U5183 ( .A(n5369), .B(n5370), .Z(n5366) );
  AND U5184 ( .A(n248), .B(n5365), .Z(n5370) );
  XNOR U5185 ( .A(n5369), .B(n5363), .Z(n5365) );
  XOR U5186 ( .A(n5371), .B(n5372), .Z(n5363) );
  AND U5187 ( .A(n263), .B(n5373), .Z(n5372) );
  XNOR U5188 ( .A(n5374), .B(n5375), .Z(n5369) );
  AND U5189 ( .A(n255), .B(n5376), .Z(n5375) );
  XOR U5190 ( .A(p_input[334]), .B(n5374), .Z(n5376) );
  XNOR U5191 ( .A(n5377), .B(n5378), .Z(n5374) );
  AND U5192 ( .A(n259), .B(n5373), .Z(n5378) );
  XNOR U5193 ( .A(n5377), .B(n5371), .Z(n5373) );
  XOR U5194 ( .A(n5379), .B(n5380), .Z(n5371) );
  AND U5195 ( .A(n274), .B(n5381), .Z(n5380) );
  XNOR U5196 ( .A(n5382), .B(n5383), .Z(n5377) );
  AND U5197 ( .A(n266), .B(n5384), .Z(n5383) );
  XOR U5198 ( .A(p_input[350]), .B(n5382), .Z(n5384) );
  XNOR U5199 ( .A(n5385), .B(n5386), .Z(n5382) );
  AND U5200 ( .A(n270), .B(n5381), .Z(n5386) );
  XNOR U5201 ( .A(n5385), .B(n5379), .Z(n5381) );
  XOR U5202 ( .A(n5387), .B(n5388), .Z(n5379) );
  AND U5203 ( .A(n285), .B(n5389), .Z(n5388) );
  XNOR U5204 ( .A(n5390), .B(n5391), .Z(n5385) );
  AND U5205 ( .A(n277), .B(n5392), .Z(n5391) );
  XOR U5206 ( .A(p_input[366]), .B(n5390), .Z(n5392) );
  XNOR U5207 ( .A(n5393), .B(n5394), .Z(n5390) );
  AND U5208 ( .A(n281), .B(n5389), .Z(n5394) );
  XNOR U5209 ( .A(n5393), .B(n5387), .Z(n5389) );
  XOR U5210 ( .A(n5395), .B(n5396), .Z(n5387) );
  AND U5211 ( .A(n296), .B(n5397), .Z(n5396) );
  XNOR U5212 ( .A(n5398), .B(n5399), .Z(n5393) );
  AND U5213 ( .A(n288), .B(n5400), .Z(n5399) );
  XOR U5214 ( .A(p_input[382]), .B(n5398), .Z(n5400) );
  XNOR U5215 ( .A(n5401), .B(n5402), .Z(n5398) );
  AND U5216 ( .A(n292), .B(n5397), .Z(n5402) );
  XNOR U5217 ( .A(n5401), .B(n5395), .Z(n5397) );
  XOR U5218 ( .A(n5403), .B(n5404), .Z(n5395) );
  AND U5219 ( .A(n307), .B(n5405), .Z(n5404) );
  XNOR U5220 ( .A(n5406), .B(n5407), .Z(n5401) );
  AND U5221 ( .A(n299), .B(n5408), .Z(n5407) );
  XOR U5222 ( .A(p_input[398]), .B(n5406), .Z(n5408) );
  XNOR U5223 ( .A(n5409), .B(n5410), .Z(n5406) );
  AND U5224 ( .A(n303), .B(n5405), .Z(n5410) );
  XNOR U5225 ( .A(n5409), .B(n5403), .Z(n5405) );
  XOR U5226 ( .A(n5411), .B(n5412), .Z(n5403) );
  AND U5227 ( .A(n318), .B(n5413), .Z(n5412) );
  XNOR U5228 ( .A(n5414), .B(n5415), .Z(n5409) );
  AND U5229 ( .A(n310), .B(n5416), .Z(n5415) );
  XOR U5230 ( .A(p_input[414]), .B(n5414), .Z(n5416) );
  XNOR U5231 ( .A(n5417), .B(n5418), .Z(n5414) );
  AND U5232 ( .A(n314), .B(n5413), .Z(n5418) );
  XNOR U5233 ( .A(n5417), .B(n5411), .Z(n5413) );
  XOR U5234 ( .A(n5419), .B(n5420), .Z(n5411) );
  AND U5235 ( .A(n329), .B(n5421), .Z(n5420) );
  XNOR U5236 ( .A(n5422), .B(n5423), .Z(n5417) );
  AND U5237 ( .A(n321), .B(n5424), .Z(n5423) );
  XOR U5238 ( .A(p_input[430]), .B(n5422), .Z(n5424) );
  XNOR U5239 ( .A(n5425), .B(n5426), .Z(n5422) );
  AND U5240 ( .A(n325), .B(n5421), .Z(n5426) );
  XNOR U5241 ( .A(n5425), .B(n5419), .Z(n5421) );
  XOR U5242 ( .A(n5427), .B(n5428), .Z(n5419) );
  AND U5243 ( .A(n340), .B(n5429), .Z(n5428) );
  XNOR U5244 ( .A(n5430), .B(n5431), .Z(n5425) );
  AND U5245 ( .A(n332), .B(n5432), .Z(n5431) );
  XOR U5246 ( .A(p_input[446]), .B(n5430), .Z(n5432) );
  XNOR U5247 ( .A(n5433), .B(n5434), .Z(n5430) );
  AND U5248 ( .A(n336), .B(n5429), .Z(n5434) );
  XNOR U5249 ( .A(n5433), .B(n5427), .Z(n5429) );
  XOR U5250 ( .A(n5435), .B(n5436), .Z(n5427) );
  AND U5251 ( .A(n351), .B(n5437), .Z(n5436) );
  XNOR U5252 ( .A(n5438), .B(n5439), .Z(n5433) );
  AND U5253 ( .A(n343), .B(n5440), .Z(n5439) );
  XOR U5254 ( .A(p_input[462]), .B(n5438), .Z(n5440) );
  XNOR U5255 ( .A(n5441), .B(n5442), .Z(n5438) );
  AND U5256 ( .A(n347), .B(n5437), .Z(n5442) );
  XNOR U5257 ( .A(n5441), .B(n5435), .Z(n5437) );
  XOR U5258 ( .A(n5443), .B(n5444), .Z(n5435) );
  AND U5259 ( .A(n362), .B(n5445), .Z(n5444) );
  XNOR U5260 ( .A(n5446), .B(n5447), .Z(n5441) );
  AND U5261 ( .A(n354), .B(n5448), .Z(n5447) );
  XOR U5262 ( .A(p_input[478]), .B(n5446), .Z(n5448) );
  XNOR U5263 ( .A(n5449), .B(n5450), .Z(n5446) );
  AND U5264 ( .A(n358), .B(n5445), .Z(n5450) );
  XNOR U5265 ( .A(n5449), .B(n5443), .Z(n5445) );
  XOR U5266 ( .A(n5451), .B(n5452), .Z(n5443) );
  AND U5267 ( .A(n373), .B(n5453), .Z(n5452) );
  XNOR U5268 ( .A(n5454), .B(n5455), .Z(n5449) );
  AND U5269 ( .A(n365), .B(n5456), .Z(n5455) );
  XOR U5270 ( .A(p_input[494]), .B(n5454), .Z(n5456) );
  XNOR U5271 ( .A(n5457), .B(n5458), .Z(n5454) );
  AND U5272 ( .A(n369), .B(n5453), .Z(n5458) );
  XNOR U5273 ( .A(n5457), .B(n5451), .Z(n5453) );
  XOR U5274 ( .A(n5459), .B(n5460), .Z(n5451) );
  AND U5275 ( .A(n384), .B(n5461), .Z(n5460) );
  XNOR U5276 ( .A(n5462), .B(n5463), .Z(n5457) );
  AND U5277 ( .A(n376), .B(n5464), .Z(n5463) );
  XOR U5278 ( .A(p_input[510]), .B(n5462), .Z(n5464) );
  XNOR U5279 ( .A(n5465), .B(n5466), .Z(n5462) );
  AND U5280 ( .A(n380), .B(n5461), .Z(n5466) );
  XNOR U5281 ( .A(n5465), .B(n5459), .Z(n5461) );
  XOR U5282 ( .A(n5467), .B(n5468), .Z(n5459) );
  AND U5283 ( .A(n395), .B(n5469), .Z(n5468) );
  XNOR U5284 ( .A(n5470), .B(n5471), .Z(n5465) );
  AND U5285 ( .A(n387), .B(n5472), .Z(n5471) );
  XOR U5286 ( .A(p_input[526]), .B(n5470), .Z(n5472) );
  XNOR U5287 ( .A(n5473), .B(n5474), .Z(n5470) );
  AND U5288 ( .A(n391), .B(n5469), .Z(n5474) );
  XNOR U5289 ( .A(n5473), .B(n5467), .Z(n5469) );
  XOR U5290 ( .A(n5475), .B(n5476), .Z(n5467) );
  AND U5291 ( .A(n406), .B(n5477), .Z(n5476) );
  XNOR U5292 ( .A(n5478), .B(n5479), .Z(n5473) );
  AND U5293 ( .A(n398), .B(n5480), .Z(n5479) );
  XOR U5294 ( .A(p_input[542]), .B(n5478), .Z(n5480) );
  XNOR U5295 ( .A(n5481), .B(n5482), .Z(n5478) );
  AND U5296 ( .A(n402), .B(n5477), .Z(n5482) );
  XNOR U5297 ( .A(n5481), .B(n5475), .Z(n5477) );
  XOR U5298 ( .A(n5483), .B(n5484), .Z(n5475) );
  AND U5299 ( .A(n417), .B(n5485), .Z(n5484) );
  XNOR U5300 ( .A(n5486), .B(n5487), .Z(n5481) );
  AND U5301 ( .A(n409), .B(n5488), .Z(n5487) );
  XOR U5302 ( .A(p_input[558]), .B(n5486), .Z(n5488) );
  XNOR U5303 ( .A(n5489), .B(n5490), .Z(n5486) );
  AND U5304 ( .A(n413), .B(n5485), .Z(n5490) );
  XNOR U5305 ( .A(n5489), .B(n5483), .Z(n5485) );
  XOR U5306 ( .A(n5491), .B(n5492), .Z(n5483) );
  AND U5307 ( .A(n428), .B(n5493), .Z(n5492) );
  XNOR U5308 ( .A(n5494), .B(n5495), .Z(n5489) );
  AND U5309 ( .A(n420), .B(n5496), .Z(n5495) );
  XOR U5310 ( .A(p_input[574]), .B(n5494), .Z(n5496) );
  XNOR U5311 ( .A(n5497), .B(n5498), .Z(n5494) );
  AND U5312 ( .A(n424), .B(n5493), .Z(n5498) );
  XNOR U5313 ( .A(n5497), .B(n5491), .Z(n5493) );
  XOR U5314 ( .A(n5499), .B(n5500), .Z(n5491) );
  AND U5315 ( .A(n439), .B(n5501), .Z(n5500) );
  XNOR U5316 ( .A(n5502), .B(n5503), .Z(n5497) );
  AND U5317 ( .A(n431), .B(n5504), .Z(n5503) );
  XOR U5318 ( .A(p_input[590]), .B(n5502), .Z(n5504) );
  XNOR U5319 ( .A(n5505), .B(n5506), .Z(n5502) );
  AND U5320 ( .A(n435), .B(n5501), .Z(n5506) );
  XNOR U5321 ( .A(n5505), .B(n5499), .Z(n5501) );
  XOR U5322 ( .A(n5507), .B(n5508), .Z(n5499) );
  AND U5323 ( .A(n450), .B(n5509), .Z(n5508) );
  XNOR U5324 ( .A(n5510), .B(n5511), .Z(n5505) );
  AND U5325 ( .A(n442), .B(n5512), .Z(n5511) );
  XOR U5326 ( .A(p_input[606]), .B(n5510), .Z(n5512) );
  XNOR U5327 ( .A(n5513), .B(n5514), .Z(n5510) );
  AND U5328 ( .A(n446), .B(n5509), .Z(n5514) );
  XNOR U5329 ( .A(n5513), .B(n5507), .Z(n5509) );
  XOR U5330 ( .A(n5515), .B(n5516), .Z(n5507) );
  AND U5331 ( .A(n461), .B(n5517), .Z(n5516) );
  XNOR U5332 ( .A(n5518), .B(n5519), .Z(n5513) );
  AND U5333 ( .A(n453), .B(n5520), .Z(n5519) );
  XOR U5334 ( .A(p_input[622]), .B(n5518), .Z(n5520) );
  XNOR U5335 ( .A(n5521), .B(n5522), .Z(n5518) );
  AND U5336 ( .A(n457), .B(n5517), .Z(n5522) );
  XNOR U5337 ( .A(n5521), .B(n5515), .Z(n5517) );
  XOR U5338 ( .A(n5523), .B(n5524), .Z(n5515) );
  AND U5339 ( .A(n472), .B(n5525), .Z(n5524) );
  XNOR U5340 ( .A(n5526), .B(n5527), .Z(n5521) );
  AND U5341 ( .A(n464), .B(n5528), .Z(n5527) );
  XOR U5342 ( .A(p_input[638]), .B(n5526), .Z(n5528) );
  XNOR U5343 ( .A(n5529), .B(n5530), .Z(n5526) );
  AND U5344 ( .A(n468), .B(n5525), .Z(n5530) );
  XNOR U5345 ( .A(n5529), .B(n5523), .Z(n5525) );
  XOR U5346 ( .A(n5531), .B(n5532), .Z(n5523) );
  AND U5347 ( .A(n483), .B(n5533), .Z(n5532) );
  XNOR U5348 ( .A(n5534), .B(n5535), .Z(n5529) );
  AND U5349 ( .A(n475), .B(n5536), .Z(n5535) );
  XOR U5350 ( .A(p_input[654]), .B(n5534), .Z(n5536) );
  XNOR U5351 ( .A(n5537), .B(n5538), .Z(n5534) );
  AND U5352 ( .A(n479), .B(n5533), .Z(n5538) );
  XNOR U5353 ( .A(n5537), .B(n5531), .Z(n5533) );
  XOR U5354 ( .A(n5539), .B(n5540), .Z(n5531) );
  AND U5355 ( .A(n494), .B(n5541), .Z(n5540) );
  XNOR U5356 ( .A(n5542), .B(n5543), .Z(n5537) );
  AND U5357 ( .A(n486), .B(n5544), .Z(n5543) );
  XOR U5358 ( .A(p_input[670]), .B(n5542), .Z(n5544) );
  XNOR U5359 ( .A(n5545), .B(n5546), .Z(n5542) );
  AND U5360 ( .A(n490), .B(n5541), .Z(n5546) );
  XNOR U5361 ( .A(n5545), .B(n5539), .Z(n5541) );
  XOR U5362 ( .A(n5547), .B(n5548), .Z(n5539) );
  AND U5363 ( .A(n505), .B(n5549), .Z(n5548) );
  XNOR U5364 ( .A(n5550), .B(n5551), .Z(n5545) );
  AND U5365 ( .A(n497), .B(n5552), .Z(n5551) );
  XOR U5366 ( .A(p_input[686]), .B(n5550), .Z(n5552) );
  XNOR U5367 ( .A(n5553), .B(n5554), .Z(n5550) );
  AND U5368 ( .A(n501), .B(n5549), .Z(n5554) );
  XNOR U5369 ( .A(n5553), .B(n5547), .Z(n5549) );
  XOR U5370 ( .A(n5555), .B(n5556), .Z(n5547) );
  AND U5371 ( .A(n516), .B(n5557), .Z(n5556) );
  XNOR U5372 ( .A(n5558), .B(n5559), .Z(n5553) );
  AND U5373 ( .A(n508), .B(n5560), .Z(n5559) );
  XOR U5374 ( .A(p_input[702]), .B(n5558), .Z(n5560) );
  XNOR U5375 ( .A(n5561), .B(n5562), .Z(n5558) );
  AND U5376 ( .A(n512), .B(n5557), .Z(n5562) );
  XNOR U5377 ( .A(n5561), .B(n5555), .Z(n5557) );
  XOR U5378 ( .A(n5563), .B(n5564), .Z(n5555) );
  AND U5379 ( .A(n527), .B(n5565), .Z(n5564) );
  XNOR U5380 ( .A(n5566), .B(n5567), .Z(n5561) );
  AND U5381 ( .A(n519), .B(n5568), .Z(n5567) );
  XOR U5382 ( .A(p_input[718]), .B(n5566), .Z(n5568) );
  XNOR U5383 ( .A(n5569), .B(n5570), .Z(n5566) );
  AND U5384 ( .A(n523), .B(n5565), .Z(n5570) );
  XNOR U5385 ( .A(n5569), .B(n5563), .Z(n5565) );
  XOR U5386 ( .A(n5571), .B(n5572), .Z(n5563) );
  AND U5387 ( .A(n538), .B(n5573), .Z(n5572) );
  XNOR U5388 ( .A(n5574), .B(n5575), .Z(n5569) );
  AND U5389 ( .A(n530), .B(n5576), .Z(n5575) );
  XOR U5390 ( .A(p_input[734]), .B(n5574), .Z(n5576) );
  XNOR U5391 ( .A(n5577), .B(n5578), .Z(n5574) );
  AND U5392 ( .A(n534), .B(n5573), .Z(n5578) );
  XNOR U5393 ( .A(n5577), .B(n5571), .Z(n5573) );
  XOR U5394 ( .A(n5579), .B(n5580), .Z(n5571) );
  AND U5395 ( .A(n549), .B(n5581), .Z(n5580) );
  XNOR U5396 ( .A(n5582), .B(n5583), .Z(n5577) );
  AND U5397 ( .A(n541), .B(n5584), .Z(n5583) );
  XOR U5398 ( .A(p_input[750]), .B(n5582), .Z(n5584) );
  XNOR U5399 ( .A(n5585), .B(n5586), .Z(n5582) );
  AND U5400 ( .A(n545), .B(n5581), .Z(n5586) );
  XNOR U5401 ( .A(n5585), .B(n5579), .Z(n5581) );
  XOR U5402 ( .A(n5587), .B(n5588), .Z(n5579) );
  AND U5403 ( .A(n560), .B(n5589), .Z(n5588) );
  XNOR U5404 ( .A(n5590), .B(n5591), .Z(n5585) );
  AND U5405 ( .A(n552), .B(n5592), .Z(n5591) );
  XOR U5406 ( .A(p_input[766]), .B(n5590), .Z(n5592) );
  XNOR U5407 ( .A(n5593), .B(n5594), .Z(n5590) );
  AND U5408 ( .A(n556), .B(n5589), .Z(n5594) );
  XNOR U5409 ( .A(n5593), .B(n5587), .Z(n5589) );
  XOR U5410 ( .A(n5595), .B(n5596), .Z(n5587) );
  AND U5411 ( .A(n571), .B(n5597), .Z(n5596) );
  XNOR U5412 ( .A(n5598), .B(n5599), .Z(n5593) );
  AND U5413 ( .A(n563), .B(n5600), .Z(n5599) );
  XOR U5414 ( .A(p_input[782]), .B(n5598), .Z(n5600) );
  XNOR U5415 ( .A(n5601), .B(n5602), .Z(n5598) );
  AND U5416 ( .A(n567), .B(n5597), .Z(n5602) );
  XNOR U5417 ( .A(n5601), .B(n5595), .Z(n5597) );
  XOR U5418 ( .A(n5603), .B(n5604), .Z(n5595) );
  AND U5419 ( .A(n582), .B(n5605), .Z(n5604) );
  XNOR U5420 ( .A(n5606), .B(n5607), .Z(n5601) );
  AND U5421 ( .A(n574), .B(n5608), .Z(n5607) );
  XOR U5422 ( .A(p_input[798]), .B(n5606), .Z(n5608) );
  XNOR U5423 ( .A(n5609), .B(n5610), .Z(n5606) );
  AND U5424 ( .A(n578), .B(n5605), .Z(n5610) );
  XNOR U5425 ( .A(n5609), .B(n5603), .Z(n5605) );
  XOR U5426 ( .A(n5611), .B(n5612), .Z(n5603) );
  AND U5427 ( .A(n593), .B(n5613), .Z(n5612) );
  XNOR U5428 ( .A(n5614), .B(n5615), .Z(n5609) );
  AND U5429 ( .A(n585), .B(n5616), .Z(n5615) );
  XOR U5430 ( .A(p_input[814]), .B(n5614), .Z(n5616) );
  XNOR U5431 ( .A(n5617), .B(n5618), .Z(n5614) );
  AND U5432 ( .A(n589), .B(n5613), .Z(n5618) );
  XNOR U5433 ( .A(n5617), .B(n5611), .Z(n5613) );
  XOR U5434 ( .A(n5619), .B(n5620), .Z(n5611) );
  AND U5435 ( .A(n604), .B(n5621), .Z(n5620) );
  XNOR U5436 ( .A(n5622), .B(n5623), .Z(n5617) );
  AND U5437 ( .A(n596), .B(n5624), .Z(n5623) );
  XOR U5438 ( .A(p_input[830]), .B(n5622), .Z(n5624) );
  XNOR U5439 ( .A(n5625), .B(n5626), .Z(n5622) );
  AND U5440 ( .A(n600), .B(n5621), .Z(n5626) );
  XNOR U5441 ( .A(n5625), .B(n5619), .Z(n5621) );
  XOR U5442 ( .A(n5627), .B(n5628), .Z(n5619) );
  AND U5443 ( .A(n615), .B(n5629), .Z(n5628) );
  XNOR U5444 ( .A(n5630), .B(n5631), .Z(n5625) );
  AND U5445 ( .A(n607), .B(n5632), .Z(n5631) );
  XOR U5446 ( .A(p_input[846]), .B(n5630), .Z(n5632) );
  XNOR U5447 ( .A(n5633), .B(n5634), .Z(n5630) );
  AND U5448 ( .A(n611), .B(n5629), .Z(n5634) );
  XNOR U5449 ( .A(n5633), .B(n5627), .Z(n5629) );
  XOR U5450 ( .A(n5635), .B(n5636), .Z(n5627) );
  AND U5451 ( .A(n626), .B(n5637), .Z(n5636) );
  XNOR U5452 ( .A(n5638), .B(n5639), .Z(n5633) );
  AND U5453 ( .A(n618), .B(n5640), .Z(n5639) );
  XOR U5454 ( .A(p_input[862]), .B(n5638), .Z(n5640) );
  XNOR U5455 ( .A(n5641), .B(n5642), .Z(n5638) );
  AND U5456 ( .A(n622), .B(n5637), .Z(n5642) );
  XNOR U5457 ( .A(n5641), .B(n5635), .Z(n5637) );
  XOR U5458 ( .A(n5643), .B(n5644), .Z(n5635) );
  AND U5459 ( .A(n637), .B(n5645), .Z(n5644) );
  XNOR U5460 ( .A(n5646), .B(n5647), .Z(n5641) );
  AND U5461 ( .A(n629), .B(n5648), .Z(n5647) );
  XOR U5462 ( .A(p_input[878]), .B(n5646), .Z(n5648) );
  XNOR U5463 ( .A(n5649), .B(n5650), .Z(n5646) );
  AND U5464 ( .A(n633), .B(n5645), .Z(n5650) );
  XNOR U5465 ( .A(n5649), .B(n5643), .Z(n5645) );
  XOR U5466 ( .A(n5651), .B(n5652), .Z(n5643) );
  AND U5467 ( .A(n648), .B(n5653), .Z(n5652) );
  XNOR U5468 ( .A(n5654), .B(n5655), .Z(n5649) );
  AND U5469 ( .A(n640), .B(n5656), .Z(n5655) );
  XOR U5470 ( .A(p_input[894]), .B(n5654), .Z(n5656) );
  XNOR U5471 ( .A(n5657), .B(n5658), .Z(n5654) );
  AND U5472 ( .A(n644), .B(n5653), .Z(n5658) );
  XNOR U5473 ( .A(n5657), .B(n5651), .Z(n5653) );
  XOR U5474 ( .A(n5659), .B(n5660), .Z(n5651) );
  AND U5475 ( .A(n659), .B(n5661), .Z(n5660) );
  XNOR U5476 ( .A(n5662), .B(n5663), .Z(n5657) );
  AND U5477 ( .A(n651), .B(n5664), .Z(n5663) );
  XOR U5478 ( .A(p_input[910]), .B(n5662), .Z(n5664) );
  XNOR U5479 ( .A(n5665), .B(n5666), .Z(n5662) );
  AND U5480 ( .A(n655), .B(n5661), .Z(n5666) );
  XNOR U5481 ( .A(n5665), .B(n5659), .Z(n5661) );
  XOR U5482 ( .A(n5667), .B(n5668), .Z(n5659) );
  AND U5483 ( .A(n670), .B(n5669), .Z(n5668) );
  XNOR U5484 ( .A(n5670), .B(n5671), .Z(n5665) );
  AND U5485 ( .A(n662), .B(n5672), .Z(n5671) );
  XOR U5486 ( .A(p_input[926]), .B(n5670), .Z(n5672) );
  XNOR U5487 ( .A(n5673), .B(n5674), .Z(n5670) );
  AND U5488 ( .A(n666), .B(n5669), .Z(n5674) );
  XNOR U5489 ( .A(n5673), .B(n5667), .Z(n5669) );
  XOR U5490 ( .A(n5675), .B(n5676), .Z(n5667) );
  AND U5491 ( .A(n681), .B(n5677), .Z(n5676) );
  XNOR U5492 ( .A(n5678), .B(n5679), .Z(n5673) );
  AND U5493 ( .A(n673), .B(n5680), .Z(n5679) );
  XOR U5494 ( .A(p_input[942]), .B(n5678), .Z(n5680) );
  XNOR U5495 ( .A(n5681), .B(n5682), .Z(n5678) );
  AND U5496 ( .A(n677), .B(n5677), .Z(n5682) );
  XNOR U5497 ( .A(n5681), .B(n5675), .Z(n5677) );
  XOR U5498 ( .A(n5683), .B(n5684), .Z(n5675) );
  AND U5499 ( .A(n692), .B(n5685), .Z(n5684) );
  XNOR U5500 ( .A(n5686), .B(n5687), .Z(n5681) );
  AND U5501 ( .A(n684), .B(n5688), .Z(n5687) );
  XOR U5502 ( .A(p_input[958]), .B(n5686), .Z(n5688) );
  XNOR U5503 ( .A(n5689), .B(n5690), .Z(n5686) );
  AND U5504 ( .A(n688), .B(n5685), .Z(n5690) );
  XNOR U5505 ( .A(n5689), .B(n5683), .Z(n5685) );
  XOR U5506 ( .A(n5691), .B(n5692), .Z(n5683) );
  AND U5507 ( .A(n703), .B(n5693), .Z(n5692) );
  XNOR U5508 ( .A(n5694), .B(n5695), .Z(n5689) );
  AND U5509 ( .A(n695), .B(n5696), .Z(n5695) );
  XOR U5510 ( .A(p_input[974]), .B(n5694), .Z(n5696) );
  XNOR U5511 ( .A(n5697), .B(n5698), .Z(n5694) );
  AND U5512 ( .A(n699), .B(n5693), .Z(n5698) );
  XNOR U5513 ( .A(n5697), .B(n5691), .Z(n5693) );
  XOR U5514 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n5699), .Z(n5691) );
  AND U5515 ( .A(n713), .B(n5700), .Z(n5699) );
  XNOR U5516 ( .A(n5701), .B(n5702), .Z(n5697) );
  AND U5517 ( .A(n706), .B(n5703), .Z(n5702) );
  XOR U5518 ( .A(p_input[990]), .B(n5701), .Z(n5703) );
  XNOR U5519 ( .A(n5704), .B(n5705), .Z(n5701) );
  AND U5520 ( .A(n710), .B(n5700), .Z(n5705) );
  XOR U5521 ( .A(n5706), .B(n5704), .Z(n5700) );
  IV U5522 ( .A(\knn_comb_/min_val_out[0][14] ), .Z(n5706) );
  IV U5523 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n5704) );
  XOR U5524 ( .A(n21), .B(n5707), .Z(o[13]) );
  AND U5525 ( .A(n30), .B(n5708), .Z(n21) );
  XOR U5526 ( .A(n22), .B(n5707), .Z(n5708) );
  XOR U5527 ( .A(n5709), .B(n5710), .Z(n5707) );
  AND U5528 ( .A(n42), .B(n5711), .Z(n5710) );
  XOR U5529 ( .A(n5712), .B(n5713), .Z(n22) );
  AND U5530 ( .A(n34), .B(n5714), .Z(n5713) );
  XOR U5531 ( .A(p_input[13]), .B(n5712), .Z(n5714) );
  XNOR U5532 ( .A(n5715), .B(n5716), .Z(n5712) );
  AND U5533 ( .A(n38), .B(n5711), .Z(n5716) );
  XNOR U5534 ( .A(n5715), .B(n5709), .Z(n5711) );
  XOR U5535 ( .A(n5717), .B(n5718), .Z(n5709) );
  AND U5536 ( .A(n54), .B(n5719), .Z(n5718) );
  XNOR U5537 ( .A(n5720), .B(n5721), .Z(n5715) );
  AND U5538 ( .A(n46), .B(n5722), .Z(n5721) );
  XOR U5539 ( .A(p_input[29]), .B(n5720), .Z(n5722) );
  XNOR U5540 ( .A(n5723), .B(n5724), .Z(n5720) );
  AND U5541 ( .A(n50), .B(n5719), .Z(n5724) );
  XNOR U5542 ( .A(n5723), .B(n5717), .Z(n5719) );
  XOR U5543 ( .A(n5725), .B(n5726), .Z(n5717) );
  AND U5544 ( .A(n65), .B(n5727), .Z(n5726) );
  XNOR U5545 ( .A(n5728), .B(n5729), .Z(n5723) );
  AND U5546 ( .A(n57), .B(n5730), .Z(n5729) );
  XOR U5547 ( .A(p_input[45]), .B(n5728), .Z(n5730) );
  XNOR U5548 ( .A(n5731), .B(n5732), .Z(n5728) );
  AND U5549 ( .A(n61), .B(n5727), .Z(n5732) );
  XNOR U5550 ( .A(n5731), .B(n5725), .Z(n5727) );
  XOR U5551 ( .A(n5733), .B(n5734), .Z(n5725) );
  AND U5552 ( .A(n76), .B(n5735), .Z(n5734) );
  XNOR U5553 ( .A(n5736), .B(n5737), .Z(n5731) );
  AND U5554 ( .A(n68), .B(n5738), .Z(n5737) );
  XOR U5555 ( .A(p_input[61]), .B(n5736), .Z(n5738) );
  XNOR U5556 ( .A(n5739), .B(n5740), .Z(n5736) );
  AND U5557 ( .A(n72), .B(n5735), .Z(n5740) );
  XNOR U5558 ( .A(n5739), .B(n5733), .Z(n5735) );
  XOR U5559 ( .A(n5741), .B(n5742), .Z(n5733) );
  AND U5560 ( .A(n87), .B(n5743), .Z(n5742) );
  XNOR U5561 ( .A(n5744), .B(n5745), .Z(n5739) );
  AND U5562 ( .A(n79), .B(n5746), .Z(n5745) );
  XOR U5563 ( .A(p_input[77]), .B(n5744), .Z(n5746) );
  XNOR U5564 ( .A(n5747), .B(n5748), .Z(n5744) );
  AND U5565 ( .A(n83), .B(n5743), .Z(n5748) );
  XNOR U5566 ( .A(n5747), .B(n5741), .Z(n5743) );
  XOR U5567 ( .A(n5749), .B(n5750), .Z(n5741) );
  AND U5568 ( .A(n98), .B(n5751), .Z(n5750) );
  XNOR U5569 ( .A(n5752), .B(n5753), .Z(n5747) );
  AND U5570 ( .A(n90), .B(n5754), .Z(n5753) );
  XOR U5571 ( .A(p_input[93]), .B(n5752), .Z(n5754) );
  XNOR U5572 ( .A(n5755), .B(n5756), .Z(n5752) );
  AND U5573 ( .A(n94), .B(n5751), .Z(n5756) );
  XNOR U5574 ( .A(n5755), .B(n5749), .Z(n5751) );
  XOR U5575 ( .A(n5757), .B(n5758), .Z(n5749) );
  AND U5576 ( .A(n109), .B(n5759), .Z(n5758) );
  XNOR U5577 ( .A(n5760), .B(n5761), .Z(n5755) );
  AND U5578 ( .A(n101), .B(n5762), .Z(n5761) );
  XOR U5579 ( .A(p_input[109]), .B(n5760), .Z(n5762) );
  XNOR U5580 ( .A(n5763), .B(n5764), .Z(n5760) );
  AND U5581 ( .A(n105), .B(n5759), .Z(n5764) );
  XNOR U5582 ( .A(n5763), .B(n5757), .Z(n5759) );
  XOR U5583 ( .A(n5765), .B(n5766), .Z(n5757) );
  AND U5584 ( .A(n120), .B(n5767), .Z(n5766) );
  XNOR U5585 ( .A(n5768), .B(n5769), .Z(n5763) );
  AND U5586 ( .A(n112), .B(n5770), .Z(n5769) );
  XOR U5587 ( .A(p_input[125]), .B(n5768), .Z(n5770) );
  XNOR U5588 ( .A(n5771), .B(n5772), .Z(n5768) );
  AND U5589 ( .A(n116), .B(n5767), .Z(n5772) );
  XNOR U5590 ( .A(n5771), .B(n5765), .Z(n5767) );
  XOR U5591 ( .A(n5773), .B(n5774), .Z(n5765) );
  AND U5592 ( .A(n131), .B(n5775), .Z(n5774) );
  XNOR U5593 ( .A(n5776), .B(n5777), .Z(n5771) );
  AND U5594 ( .A(n123), .B(n5778), .Z(n5777) );
  XOR U5595 ( .A(p_input[141]), .B(n5776), .Z(n5778) );
  XNOR U5596 ( .A(n5779), .B(n5780), .Z(n5776) );
  AND U5597 ( .A(n127), .B(n5775), .Z(n5780) );
  XNOR U5598 ( .A(n5779), .B(n5773), .Z(n5775) );
  XOR U5599 ( .A(n5781), .B(n5782), .Z(n5773) );
  AND U5600 ( .A(n142), .B(n5783), .Z(n5782) );
  XNOR U5601 ( .A(n5784), .B(n5785), .Z(n5779) );
  AND U5602 ( .A(n134), .B(n5786), .Z(n5785) );
  XOR U5603 ( .A(p_input[157]), .B(n5784), .Z(n5786) );
  XNOR U5604 ( .A(n5787), .B(n5788), .Z(n5784) );
  AND U5605 ( .A(n138), .B(n5783), .Z(n5788) );
  XNOR U5606 ( .A(n5787), .B(n5781), .Z(n5783) );
  XOR U5607 ( .A(n5789), .B(n5790), .Z(n5781) );
  AND U5608 ( .A(n153), .B(n5791), .Z(n5790) );
  XNOR U5609 ( .A(n5792), .B(n5793), .Z(n5787) );
  AND U5610 ( .A(n145), .B(n5794), .Z(n5793) );
  XOR U5611 ( .A(p_input[173]), .B(n5792), .Z(n5794) );
  XNOR U5612 ( .A(n5795), .B(n5796), .Z(n5792) );
  AND U5613 ( .A(n149), .B(n5791), .Z(n5796) );
  XNOR U5614 ( .A(n5795), .B(n5789), .Z(n5791) );
  XOR U5615 ( .A(n5797), .B(n5798), .Z(n5789) );
  AND U5616 ( .A(n164), .B(n5799), .Z(n5798) );
  XNOR U5617 ( .A(n5800), .B(n5801), .Z(n5795) );
  AND U5618 ( .A(n156), .B(n5802), .Z(n5801) );
  XOR U5619 ( .A(p_input[189]), .B(n5800), .Z(n5802) );
  XNOR U5620 ( .A(n5803), .B(n5804), .Z(n5800) );
  AND U5621 ( .A(n160), .B(n5799), .Z(n5804) );
  XNOR U5622 ( .A(n5803), .B(n5797), .Z(n5799) );
  XOR U5623 ( .A(n5805), .B(n5806), .Z(n5797) );
  AND U5624 ( .A(n175), .B(n5807), .Z(n5806) );
  XNOR U5625 ( .A(n5808), .B(n5809), .Z(n5803) );
  AND U5626 ( .A(n167), .B(n5810), .Z(n5809) );
  XOR U5627 ( .A(p_input[205]), .B(n5808), .Z(n5810) );
  XNOR U5628 ( .A(n5811), .B(n5812), .Z(n5808) );
  AND U5629 ( .A(n171), .B(n5807), .Z(n5812) );
  XNOR U5630 ( .A(n5811), .B(n5805), .Z(n5807) );
  XOR U5631 ( .A(n5813), .B(n5814), .Z(n5805) );
  AND U5632 ( .A(n186), .B(n5815), .Z(n5814) );
  XNOR U5633 ( .A(n5816), .B(n5817), .Z(n5811) );
  AND U5634 ( .A(n178), .B(n5818), .Z(n5817) );
  XOR U5635 ( .A(p_input[221]), .B(n5816), .Z(n5818) );
  XNOR U5636 ( .A(n5819), .B(n5820), .Z(n5816) );
  AND U5637 ( .A(n182), .B(n5815), .Z(n5820) );
  XNOR U5638 ( .A(n5819), .B(n5813), .Z(n5815) );
  XOR U5639 ( .A(n5821), .B(n5822), .Z(n5813) );
  AND U5640 ( .A(n197), .B(n5823), .Z(n5822) );
  XNOR U5641 ( .A(n5824), .B(n5825), .Z(n5819) );
  AND U5642 ( .A(n189), .B(n5826), .Z(n5825) );
  XOR U5643 ( .A(p_input[237]), .B(n5824), .Z(n5826) );
  XNOR U5644 ( .A(n5827), .B(n5828), .Z(n5824) );
  AND U5645 ( .A(n193), .B(n5823), .Z(n5828) );
  XNOR U5646 ( .A(n5827), .B(n5821), .Z(n5823) );
  XOR U5647 ( .A(n5829), .B(n5830), .Z(n5821) );
  AND U5648 ( .A(n208), .B(n5831), .Z(n5830) );
  XNOR U5649 ( .A(n5832), .B(n5833), .Z(n5827) );
  AND U5650 ( .A(n200), .B(n5834), .Z(n5833) );
  XOR U5651 ( .A(p_input[253]), .B(n5832), .Z(n5834) );
  XNOR U5652 ( .A(n5835), .B(n5836), .Z(n5832) );
  AND U5653 ( .A(n204), .B(n5831), .Z(n5836) );
  XNOR U5654 ( .A(n5835), .B(n5829), .Z(n5831) );
  XOR U5655 ( .A(n5837), .B(n5838), .Z(n5829) );
  AND U5656 ( .A(n219), .B(n5839), .Z(n5838) );
  XNOR U5657 ( .A(n5840), .B(n5841), .Z(n5835) );
  AND U5658 ( .A(n211), .B(n5842), .Z(n5841) );
  XOR U5659 ( .A(p_input[269]), .B(n5840), .Z(n5842) );
  XNOR U5660 ( .A(n5843), .B(n5844), .Z(n5840) );
  AND U5661 ( .A(n215), .B(n5839), .Z(n5844) );
  XNOR U5662 ( .A(n5843), .B(n5837), .Z(n5839) );
  XOR U5663 ( .A(n5845), .B(n5846), .Z(n5837) );
  AND U5664 ( .A(n230), .B(n5847), .Z(n5846) );
  XNOR U5665 ( .A(n5848), .B(n5849), .Z(n5843) );
  AND U5666 ( .A(n222), .B(n5850), .Z(n5849) );
  XOR U5667 ( .A(p_input[285]), .B(n5848), .Z(n5850) );
  XNOR U5668 ( .A(n5851), .B(n5852), .Z(n5848) );
  AND U5669 ( .A(n226), .B(n5847), .Z(n5852) );
  XNOR U5670 ( .A(n5851), .B(n5845), .Z(n5847) );
  XOR U5671 ( .A(n5853), .B(n5854), .Z(n5845) );
  AND U5672 ( .A(n241), .B(n5855), .Z(n5854) );
  XNOR U5673 ( .A(n5856), .B(n5857), .Z(n5851) );
  AND U5674 ( .A(n233), .B(n5858), .Z(n5857) );
  XOR U5675 ( .A(p_input[301]), .B(n5856), .Z(n5858) );
  XNOR U5676 ( .A(n5859), .B(n5860), .Z(n5856) );
  AND U5677 ( .A(n237), .B(n5855), .Z(n5860) );
  XNOR U5678 ( .A(n5859), .B(n5853), .Z(n5855) );
  XOR U5679 ( .A(n5861), .B(n5862), .Z(n5853) );
  AND U5680 ( .A(n252), .B(n5863), .Z(n5862) );
  XNOR U5681 ( .A(n5864), .B(n5865), .Z(n5859) );
  AND U5682 ( .A(n244), .B(n5866), .Z(n5865) );
  XOR U5683 ( .A(p_input[317]), .B(n5864), .Z(n5866) );
  XNOR U5684 ( .A(n5867), .B(n5868), .Z(n5864) );
  AND U5685 ( .A(n248), .B(n5863), .Z(n5868) );
  XNOR U5686 ( .A(n5867), .B(n5861), .Z(n5863) );
  XOR U5687 ( .A(n5869), .B(n5870), .Z(n5861) );
  AND U5688 ( .A(n263), .B(n5871), .Z(n5870) );
  XNOR U5689 ( .A(n5872), .B(n5873), .Z(n5867) );
  AND U5690 ( .A(n255), .B(n5874), .Z(n5873) );
  XOR U5691 ( .A(p_input[333]), .B(n5872), .Z(n5874) );
  XNOR U5692 ( .A(n5875), .B(n5876), .Z(n5872) );
  AND U5693 ( .A(n259), .B(n5871), .Z(n5876) );
  XNOR U5694 ( .A(n5875), .B(n5869), .Z(n5871) );
  XOR U5695 ( .A(n5877), .B(n5878), .Z(n5869) );
  AND U5696 ( .A(n274), .B(n5879), .Z(n5878) );
  XNOR U5697 ( .A(n5880), .B(n5881), .Z(n5875) );
  AND U5698 ( .A(n266), .B(n5882), .Z(n5881) );
  XOR U5699 ( .A(p_input[349]), .B(n5880), .Z(n5882) );
  XNOR U5700 ( .A(n5883), .B(n5884), .Z(n5880) );
  AND U5701 ( .A(n270), .B(n5879), .Z(n5884) );
  XNOR U5702 ( .A(n5883), .B(n5877), .Z(n5879) );
  XOR U5703 ( .A(n5885), .B(n5886), .Z(n5877) );
  AND U5704 ( .A(n285), .B(n5887), .Z(n5886) );
  XNOR U5705 ( .A(n5888), .B(n5889), .Z(n5883) );
  AND U5706 ( .A(n277), .B(n5890), .Z(n5889) );
  XOR U5707 ( .A(p_input[365]), .B(n5888), .Z(n5890) );
  XNOR U5708 ( .A(n5891), .B(n5892), .Z(n5888) );
  AND U5709 ( .A(n281), .B(n5887), .Z(n5892) );
  XNOR U5710 ( .A(n5891), .B(n5885), .Z(n5887) );
  XOR U5711 ( .A(n5893), .B(n5894), .Z(n5885) );
  AND U5712 ( .A(n296), .B(n5895), .Z(n5894) );
  XNOR U5713 ( .A(n5896), .B(n5897), .Z(n5891) );
  AND U5714 ( .A(n288), .B(n5898), .Z(n5897) );
  XOR U5715 ( .A(p_input[381]), .B(n5896), .Z(n5898) );
  XNOR U5716 ( .A(n5899), .B(n5900), .Z(n5896) );
  AND U5717 ( .A(n292), .B(n5895), .Z(n5900) );
  XNOR U5718 ( .A(n5899), .B(n5893), .Z(n5895) );
  XOR U5719 ( .A(n5901), .B(n5902), .Z(n5893) );
  AND U5720 ( .A(n307), .B(n5903), .Z(n5902) );
  XNOR U5721 ( .A(n5904), .B(n5905), .Z(n5899) );
  AND U5722 ( .A(n299), .B(n5906), .Z(n5905) );
  XOR U5723 ( .A(p_input[397]), .B(n5904), .Z(n5906) );
  XNOR U5724 ( .A(n5907), .B(n5908), .Z(n5904) );
  AND U5725 ( .A(n303), .B(n5903), .Z(n5908) );
  XNOR U5726 ( .A(n5907), .B(n5901), .Z(n5903) );
  XOR U5727 ( .A(n5909), .B(n5910), .Z(n5901) );
  AND U5728 ( .A(n318), .B(n5911), .Z(n5910) );
  XNOR U5729 ( .A(n5912), .B(n5913), .Z(n5907) );
  AND U5730 ( .A(n310), .B(n5914), .Z(n5913) );
  XOR U5731 ( .A(p_input[413]), .B(n5912), .Z(n5914) );
  XNOR U5732 ( .A(n5915), .B(n5916), .Z(n5912) );
  AND U5733 ( .A(n314), .B(n5911), .Z(n5916) );
  XNOR U5734 ( .A(n5915), .B(n5909), .Z(n5911) );
  XOR U5735 ( .A(n5917), .B(n5918), .Z(n5909) );
  AND U5736 ( .A(n329), .B(n5919), .Z(n5918) );
  XNOR U5737 ( .A(n5920), .B(n5921), .Z(n5915) );
  AND U5738 ( .A(n321), .B(n5922), .Z(n5921) );
  XOR U5739 ( .A(p_input[429]), .B(n5920), .Z(n5922) );
  XNOR U5740 ( .A(n5923), .B(n5924), .Z(n5920) );
  AND U5741 ( .A(n325), .B(n5919), .Z(n5924) );
  XNOR U5742 ( .A(n5923), .B(n5917), .Z(n5919) );
  XOR U5743 ( .A(n5925), .B(n5926), .Z(n5917) );
  AND U5744 ( .A(n340), .B(n5927), .Z(n5926) );
  XNOR U5745 ( .A(n5928), .B(n5929), .Z(n5923) );
  AND U5746 ( .A(n332), .B(n5930), .Z(n5929) );
  XOR U5747 ( .A(p_input[445]), .B(n5928), .Z(n5930) );
  XNOR U5748 ( .A(n5931), .B(n5932), .Z(n5928) );
  AND U5749 ( .A(n336), .B(n5927), .Z(n5932) );
  XNOR U5750 ( .A(n5931), .B(n5925), .Z(n5927) );
  XOR U5751 ( .A(n5933), .B(n5934), .Z(n5925) );
  AND U5752 ( .A(n351), .B(n5935), .Z(n5934) );
  XNOR U5753 ( .A(n5936), .B(n5937), .Z(n5931) );
  AND U5754 ( .A(n343), .B(n5938), .Z(n5937) );
  XOR U5755 ( .A(p_input[461]), .B(n5936), .Z(n5938) );
  XNOR U5756 ( .A(n5939), .B(n5940), .Z(n5936) );
  AND U5757 ( .A(n347), .B(n5935), .Z(n5940) );
  XNOR U5758 ( .A(n5939), .B(n5933), .Z(n5935) );
  XOR U5759 ( .A(n5941), .B(n5942), .Z(n5933) );
  AND U5760 ( .A(n362), .B(n5943), .Z(n5942) );
  XNOR U5761 ( .A(n5944), .B(n5945), .Z(n5939) );
  AND U5762 ( .A(n354), .B(n5946), .Z(n5945) );
  XOR U5763 ( .A(p_input[477]), .B(n5944), .Z(n5946) );
  XNOR U5764 ( .A(n5947), .B(n5948), .Z(n5944) );
  AND U5765 ( .A(n358), .B(n5943), .Z(n5948) );
  XNOR U5766 ( .A(n5947), .B(n5941), .Z(n5943) );
  XOR U5767 ( .A(n5949), .B(n5950), .Z(n5941) );
  AND U5768 ( .A(n373), .B(n5951), .Z(n5950) );
  XNOR U5769 ( .A(n5952), .B(n5953), .Z(n5947) );
  AND U5770 ( .A(n365), .B(n5954), .Z(n5953) );
  XOR U5771 ( .A(p_input[493]), .B(n5952), .Z(n5954) );
  XNOR U5772 ( .A(n5955), .B(n5956), .Z(n5952) );
  AND U5773 ( .A(n369), .B(n5951), .Z(n5956) );
  XNOR U5774 ( .A(n5955), .B(n5949), .Z(n5951) );
  XOR U5775 ( .A(n5957), .B(n5958), .Z(n5949) );
  AND U5776 ( .A(n384), .B(n5959), .Z(n5958) );
  XNOR U5777 ( .A(n5960), .B(n5961), .Z(n5955) );
  AND U5778 ( .A(n376), .B(n5962), .Z(n5961) );
  XOR U5779 ( .A(p_input[509]), .B(n5960), .Z(n5962) );
  XNOR U5780 ( .A(n5963), .B(n5964), .Z(n5960) );
  AND U5781 ( .A(n380), .B(n5959), .Z(n5964) );
  XNOR U5782 ( .A(n5963), .B(n5957), .Z(n5959) );
  XOR U5783 ( .A(n5965), .B(n5966), .Z(n5957) );
  AND U5784 ( .A(n395), .B(n5967), .Z(n5966) );
  XNOR U5785 ( .A(n5968), .B(n5969), .Z(n5963) );
  AND U5786 ( .A(n387), .B(n5970), .Z(n5969) );
  XOR U5787 ( .A(p_input[525]), .B(n5968), .Z(n5970) );
  XNOR U5788 ( .A(n5971), .B(n5972), .Z(n5968) );
  AND U5789 ( .A(n391), .B(n5967), .Z(n5972) );
  XNOR U5790 ( .A(n5971), .B(n5965), .Z(n5967) );
  XOR U5791 ( .A(n5973), .B(n5974), .Z(n5965) );
  AND U5792 ( .A(n406), .B(n5975), .Z(n5974) );
  XNOR U5793 ( .A(n5976), .B(n5977), .Z(n5971) );
  AND U5794 ( .A(n398), .B(n5978), .Z(n5977) );
  XOR U5795 ( .A(p_input[541]), .B(n5976), .Z(n5978) );
  XNOR U5796 ( .A(n5979), .B(n5980), .Z(n5976) );
  AND U5797 ( .A(n402), .B(n5975), .Z(n5980) );
  XNOR U5798 ( .A(n5979), .B(n5973), .Z(n5975) );
  XOR U5799 ( .A(n5981), .B(n5982), .Z(n5973) );
  AND U5800 ( .A(n417), .B(n5983), .Z(n5982) );
  XNOR U5801 ( .A(n5984), .B(n5985), .Z(n5979) );
  AND U5802 ( .A(n409), .B(n5986), .Z(n5985) );
  XOR U5803 ( .A(p_input[557]), .B(n5984), .Z(n5986) );
  XNOR U5804 ( .A(n5987), .B(n5988), .Z(n5984) );
  AND U5805 ( .A(n413), .B(n5983), .Z(n5988) );
  XNOR U5806 ( .A(n5987), .B(n5981), .Z(n5983) );
  XOR U5807 ( .A(n5989), .B(n5990), .Z(n5981) );
  AND U5808 ( .A(n428), .B(n5991), .Z(n5990) );
  XNOR U5809 ( .A(n5992), .B(n5993), .Z(n5987) );
  AND U5810 ( .A(n420), .B(n5994), .Z(n5993) );
  XOR U5811 ( .A(p_input[573]), .B(n5992), .Z(n5994) );
  XNOR U5812 ( .A(n5995), .B(n5996), .Z(n5992) );
  AND U5813 ( .A(n424), .B(n5991), .Z(n5996) );
  XNOR U5814 ( .A(n5995), .B(n5989), .Z(n5991) );
  XOR U5815 ( .A(n5997), .B(n5998), .Z(n5989) );
  AND U5816 ( .A(n439), .B(n5999), .Z(n5998) );
  XNOR U5817 ( .A(n6000), .B(n6001), .Z(n5995) );
  AND U5818 ( .A(n431), .B(n6002), .Z(n6001) );
  XOR U5819 ( .A(p_input[589]), .B(n6000), .Z(n6002) );
  XNOR U5820 ( .A(n6003), .B(n6004), .Z(n6000) );
  AND U5821 ( .A(n435), .B(n5999), .Z(n6004) );
  XNOR U5822 ( .A(n6003), .B(n5997), .Z(n5999) );
  XOR U5823 ( .A(n6005), .B(n6006), .Z(n5997) );
  AND U5824 ( .A(n450), .B(n6007), .Z(n6006) );
  XNOR U5825 ( .A(n6008), .B(n6009), .Z(n6003) );
  AND U5826 ( .A(n442), .B(n6010), .Z(n6009) );
  XOR U5827 ( .A(p_input[605]), .B(n6008), .Z(n6010) );
  XNOR U5828 ( .A(n6011), .B(n6012), .Z(n6008) );
  AND U5829 ( .A(n446), .B(n6007), .Z(n6012) );
  XNOR U5830 ( .A(n6011), .B(n6005), .Z(n6007) );
  XOR U5831 ( .A(n6013), .B(n6014), .Z(n6005) );
  AND U5832 ( .A(n461), .B(n6015), .Z(n6014) );
  XNOR U5833 ( .A(n6016), .B(n6017), .Z(n6011) );
  AND U5834 ( .A(n453), .B(n6018), .Z(n6017) );
  XOR U5835 ( .A(p_input[621]), .B(n6016), .Z(n6018) );
  XNOR U5836 ( .A(n6019), .B(n6020), .Z(n6016) );
  AND U5837 ( .A(n457), .B(n6015), .Z(n6020) );
  XNOR U5838 ( .A(n6019), .B(n6013), .Z(n6015) );
  XOR U5839 ( .A(n6021), .B(n6022), .Z(n6013) );
  AND U5840 ( .A(n472), .B(n6023), .Z(n6022) );
  XNOR U5841 ( .A(n6024), .B(n6025), .Z(n6019) );
  AND U5842 ( .A(n464), .B(n6026), .Z(n6025) );
  XOR U5843 ( .A(p_input[637]), .B(n6024), .Z(n6026) );
  XNOR U5844 ( .A(n6027), .B(n6028), .Z(n6024) );
  AND U5845 ( .A(n468), .B(n6023), .Z(n6028) );
  XNOR U5846 ( .A(n6027), .B(n6021), .Z(n6023) );
  XOR U5847 ( .A(n6029), .B(n6030), .Z(n6021) );
  AND U5848 ( .A(n483), .B(n6031), .Z(n6030) );
  XNOR U5849 ( .A(n6032), .B(n6033), .Z(n6027) );
  AND U5850 ( .A(n475), .B(n6034), .Z(n6033) );
  XOR U5851 ( .A(p_input[653]), .B(n6032), .Z(n6034) );
  XNOR U5852 ( .A(n6035), .B(n6036), .Z(n6032) );
  AND U5853 ( .A(n479), .B(n6031), .Z(n6036) );
  XNOR U5854 ( .A(n6035), .B(n6029), .Z(n6031) );
  XOR U5855 ( .A(n6037), .B(n6038), .Z(n6029) );
  AND U5856 ( .A(n494), .B(n6039), .Z(n6038) );
  XNOR U5857 ( .A(n6040), .B(n6041), .Z(n6035) );
  AND U5858 ( .A(n486), .B(n6042), .Z(n6041) );
  XOR U5859 ( .A(p_input[669]), .B(n6040), .Z(n6042) );
  XNOR U5860 ( .A(n6043), .B(n6044), .Z(n6040) );
  AND U5861 ( .A(n490), .B(n6039), .Z(n6044) );
  XNOR U5862 ( .A(n6043), .B(n6037), .Z(n6039) );
  XOR U5863 ( .A(n6045), .B(n6046), .Z(n6037) );
  AND U5864 ( .A(n505), .B(n6047), .Z(n6046) );
  XNOR U5865 ( .A(n6048), .B(n6049), .Z(n6043) );
  AND U5866 ( .A(n497), .B(n6050), .Z(n6049) );
  XOR U5867 ( .A(p_input[685]), .B(n6048), .Z(n6050) );
  XNOR U5868 ( .A(n6051), .B(n6052), .Z(n6048) );
  AND U5869 ( .A(n501), .B(n6047), .Z(n6052) );
  XNOR U5870 ( .A(n6051), .B(n6045), .Z(n6047) );
  XOR U5871 ( .A(n6053), .B(n6054), .Z(n6045) );
  AND U5872 ( .A(n516), .B(n6055), .Z(n6054) );
  XNOR U5873 ( .A(n6056), .B(n6057), .Z(n6051) );
  AND U5874 ( .A(n508), .B(n6058), .Z(n6057) );
  XOR U5875 ( .A(p_input[701]), .B(n6056), .Z(n6058) );
  XNOR U5876 ( .A(n6059), .B(n6060), .Z(n6056) );
  AND U5877 ( .A(n512), .B(n6055), .Z(n6060) );
  XNOR U5878 ( .A(n6059), .B(n6053), .Z(n6055) );
  XOR U5879 ( .A(n6061), .B(n6062), .Z(n6053) );
  AND U5880 ( .A(n527), .B(n6063), .Z(n6062) );
  XNOR U5881 ( .A(n6064), .B(n6065), .Z(n6059) );
  AND U5882 ( .A(n519), .B(n6066), .Z(n6065) );
  XOR U5883 ( .A(p_input[717]), .B(n6064), .Z(n6066) );
  XNOR U5884 ( .A(n6067), .B(n6068), .Z(n6064) );
  AND U5885 ( .A(n523), .B(n6063), .Z(n6068) );
  XNOR U5886 ( .A(n6067), .B(n6061), .Z(n6063) );
  XOR U5887 ( .A(n6069), .B(n6070), .Z(n6061) );
  AND U5888 ( .A(n538), .B(n6071), .Z(n6070) );
  XNOR U5889 ( .A(n6072), .B(n6073), .Z(n6067) );
  AND U5890 ( .A(n530), .B(n6074), .Z(n6073) );
  XOR U5891 ( .A(p_input[733]), .B(n6072), .Z(n6074) );
  XNOR U5892 ( .A(n6075), .B(n6076), .Z(n6072) );
  AND U5893 ( .A(n534), .B(n6071), .Z(n6076) );
  XNOR U5894 ( .A(n6075), .B(n6069), .Z(n6071) );
  XOR U5895 ( .A(n6077), .B(n6078), .Z(n6069) );
  AND U5896 ( .A(n549), .B(n6079), .Z(n6078) );
  XNOR U5897 ( .A(n6080), .B(n6081), .Z(n6075) );
  AND U5898 ( .A(n541), .B(n6082), .Z(n6081) );
  XOR U5899 ( .A(p_input[749]), .B(n6080), .Z(n6082) );
  XNOR U5900 ( .A(n6083), .B(n6084), .Z(n6080) );
  AND U5901 ( .A(n545), .B(n6079), .Z(n6084) );
  XNOR U5902 ( .A(n6083), .B(n6077), .Z(n6079) );
  XOR U5903 ( .A(n6085), .B(n6086), .Z(n6077) );
  AND U5904 ( .A(n560), .B(n6087), .Z(n6086) );
  XNOR U5905 ( .A(n6088), .B(n6089), .Z(n6083) );
  AND U5906 ( .A(n552), .B(n6090), .Z(n6089) );
  XOR U5907 ( .A(p_input[765]), .B(n6088), .Z(n6090) );
  XNOR U5908 ( .A(n6091), .B(n6092), .Z(n6088) );
  AND U5909 ( .A(n556), .B(n6087), .Z(n6092) );
  XNOR U5910 ( .A(n6091), .B(n6085), .Z(n6087) );
  XOR U5911 ( .A(n6093), .B(n6094), .Z(n6085) );
  AND U5912 ( .A(n571), .B(n6095), .Z(n6094) );
  XNOR U5913 ( .A(n6096), .B(n6097), .Z(n6091) );
  AND U5914 ( .A(n563), .B(n6098), .Z(n6097) );
  XOR U5915 ( .A(p_input[781]), .B(n6096), .Z(n6098) );
  XNOR U5916 ( .A(n6099), .B(n6100), .Z(n6096) );
  AND U5917 ( .A(n567), .B(n6095), .Z(n6100) );
  XNOR U5918 ( .A(n6099), .B(n6093), .Z(n6095) );
  XOR U5919 ( .A(n6101), .B(n6102), .Z(n6093) );
  AND U5920 ( .A(n582), .B(n6103), .Z(n6102) );
  XNOR U5921 ( .A(n6104), .B(n6105), .Z(n6099) );
  AND U5922 ( .A(n574), .B(n6106), .Z(n6105) );
  XOR U5923 ( .A(p_input[797]), .B(n6104), .Z(n6106) );
  XNOR U5924 ( .A(n6107), .B(n6108), .Z(n6104) );
  AND U5925 ( .A(n578), .B(n6103), .Z(n6108) );
  XNOR U5926 ( .A(n6107), .B(n6101), .Z(n6103) );
  XOR U5927 ( .A(n6109), .B(n6110), .Z(n6101) );
  AND U5928 ( .A(n593), .B(n6111), .Z(n6110) );
  XNOR U5929 ( .A(n6112), .B(n6113), .Z(n6107) );
  AND U5930 ( .A(n585), .B(n6114), .Z(n6113) );
  XOR U5931 ( .A(p_input[813]), .B(n6112), .Z(n6114) );
  XNOR U5932 ( .A(n6115), .B(n6116), .Z(n6112) );
  AND U5933 ( .A(n589), .B(n6111), .Z(n6116) );
  XNOR U5934 ( .A(n6115), .B(n6109), .Z(n6111) );
  XOR U5935 ( .A(n6117), .B(n6118), .Z(n6109) );
  AND U5936 ( .A(n604), .B(n6119), .Z(n6118) );
  XNOR U5937 ( .A(n6120), .B(n6121), .Z(n6115) );
  AND U5938 ( .A(n596), .B(n6122), .Z(n6121) );
  XOR U5939 ( .A(p_input[829]), .B(n6120), .Z(n6122) );
  XNOR U5940 ( .A(n6123), .B(n6124), .Z(n6120) );
  AND U5941 ( .A(n600), .B(n6119), .Z(n6124) );
  XNOR U5942 ( .A(n6123), .B(n6117), .Z(n6119) );
  XOR U5943 ( .A(n6125), .B(n6126), .Z(n6117) );
  AND U5944 ( .A(n615), .B(n6127), .Z(n6126) );
  XNOR U5945 ( .A(n6128), .B(n6129), .Z(n6123) );
  AND U5946 ( .A(n607), .B(n6130), .Z(n6129) );
  XOR U5947 ( .A(p_input[845]), .B(n6128), .Z(n6130) );
  XNOR U5948 ( .A(n6131), .B(n6132), .Z(n6128) );
  AND U5949 ( .A(n611), .B(n6127), .Z(n6132) );
  XNOR U5950 ( .A(n6131), .B(n6125), .Z(n6127) );
  XOR U5951 ( .A(n6133), .B(n6134), .Z(n6125) );
  AND U5952 ( .A(n626), .B(n6135), .Z(n6134) );
  XNOR U5953 ( .A(n6136), .B(n6137), .Z(n6131) );
  AND U5954 ( .A(n618), .B(n6138), .Z(n6137) );
  XOR U5955 ( .A(p_input[861]), .B(n6136), .Z(n6138) );
  XNOR U5956 ( .A(n6139), .B(n6140), .Z(n6136) );
  AND U5957 ( .A(n622), .B(n6135), .Z(n6140) );
  XNOR U5958 ( .A(n6139), .B(n6133), .Z(n6135) );
  XOR U5959 ( .A(n6141), .B(n6142), .Z(n6133) );
  AND U5960 ( .A(n637), .B(n6143), .Z(n6142) );
  XNOR U5961 ( .A(n6144), .B(n6145), .Z(n6139) );
  AND U5962 ( .A(n629), .B(n6146), .Z(n6145) );
  XOR U5963 ( .A(p_input[877]), .B(n6144), .Z(n6146) );
  XNOR U5964 ( .A(n6147), .B(n6148), .Z(n6144) );
  AND U5965 ( .A(n633), .B(n6143), .Z(n6148) );
  XNOR U5966 ( .A(n6147), .B(n6141), .Z(n6143) );
  XOR U5967 ( .A(n6149), .B(n6150), .Z(n6141) );
  AND U5968 ( .A(n648), .B(n6151), .Z(n6150) );
  XNOR U5969 ( .A(n6152), .B(n6153), .Z(n6147) );
  AND U5970 ( .A(n640), .B(n6154), .Z(n6153) );
  XOR U5971 ( .A(p_input[893]), .B(n6152), .Z(n6154) );
  XNOR U5972 ( .A(n6155), .B(n6156), .Z(n6152) );
  AND U5973 ( .A(n644), .B(n6151), .Z(n6156) );
  XNOR U5974 ( .A(n6155), .B(n6149), .Z(n6151) );
  XOR U5975 ( .A(n6157), .B(n6158), .Z(n6149) );
  AND U5976 ( .A(n659), .B(n6159), .Z(n6158) );
  XNOR U5977 ( .A(n6160), .B(n6161), .Z(n6155) );
  AND U5978 ( .A(n651), .B(n6162), .Z(n6161) );
  XOR U5979 ( .A(p_input[909]), .B(n6160), .Z(n6162) );
  XNOR U5980 ( .A(n6163), .B(n6164), .Z(n6160) );
  AND U5981 ( .A(n655), .B(n6159), .Z(n6164) );
  XNOR U5982 ( .A(n6163), .B(n6157), .Z(n6159) );
  XOR U5983 ( .A(n6165), .B(n6166), .Z(n6157) );
  AND U5984 ( .A(n670), .B(n6167), .Z(n6166) );
  XNOR U5985 ( .A(n6168), .B(n6169), .Z(n6163) );
  AND U5986 ( .A(n662), .B(n6170), .Z(n6169) );
  XOR U5987 ( .A(p_input[925]), .B(n6168), .Z(n6170) );
  XNOR U5988 ( .A(n6171), .B(n6172), .Z(n6168) );
  AND U5989 ( .A(n666), .B(n6167), .Z(n6172) );
  XNOR U5990 ( .A(n6171), .B(n6165), .Z(n6167) );
  XOR U5991 ( .A(n6173), .B(n6174), .Z(n6165) );
  AND U5992 ( .A(n681), .B(n6175), .Z(n6174) );
  XNOR U5993 ( .A(n6176), .B(n6177), .Z(n6171) );
  AND U5994 ( .A(n673), .B(n6178), .Z(n6177) );
  XOR U5995 ( .A(p_input[941]), .B(n6176), .Z(n6178) );
  XNOR U5996 ( .A(n6179), .B(n6180), .Z(n6176) );
  AND U5997 ( .A(n677), .B(n6175), .Z(n6180) );
  XNOR U5998 ( .A(n6179), .B(n6173), .Z(n6175) );
  XOR U5999 ( .A(n6181), .B(n6182), .Z(n6173) );
  AND U6000 ( .A(n692), .B(n6183), .Z(n6182) );
  XNOR U6001 ( .A(n6184), .B(n6185), .Z(n6179) );
  AND U6002 ( .A(n684), .B(n6186), .Z(n6185) );
  XOR U6003 ( .A(p_input[957]), .B(n6184), .Z(n6186) );
  XNOR U6004 ( .A(n6187), .B(n6188), .Z(n6184) );
  AND U6005 ( .A(n688), .B(n6183), .Z(n6188) );
  XNOR U6006 ( .A(n6187), .B(n6181), .Z(n6183) );
  XOR U6007 ( .A(n6189), .B(n6190), .Z(n6181) );
  AND U6008 ( .A(n703), .B(n6191), .Z(n6190) );
  XNOR U6009 ( .A(n6192), .B(n6193), .Z(n6187) );
  AND U6010 ( .A(n695), .B(n6194), .Z(n6193) );
  XOR U6011 ( .A(p_input[973]), .B(n6192), .Z(n6194) );
  XNOR U6012 ( .A(n6195), .B(n6196), .Z(n6192) );
  AND U6013 ( .A(n699), .B(n6191), .Z(n6196) );
  XNOR U6014 ( .A(n6195), .B(n6189), .Z(n6191) );
  XOR U6015 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n6197), .Z(n6189) );
  AND U6016 ( .A(n713), .B(n6198), .Z(n6197) );
  XNOR U6017 ( .A(n6199), .B(n6200), .Z(n6195) );
  AND U6018 ( .A(n706), .B(n6201), .Z(n6200) );
  XOR U6019 ( .A(p_input[989]), .B(n6199), .Z(n6201) );
  XNOR U6020 ( .A(n6202), .B(n6203), .Z(n6199) );
  AND U6021 ( .A(n710), .B(n6198), .Z(n6203) );
  XOR U6022 ( .A(\knn_comb_/min_val_out[0][13] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n6198) );
  IV U6023 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n6202) );
  XOR U6024 ( .A(n23), .B(n6204), .Z(o[12]) );
  AND U6025 ( .A(n30), .B(n6205), .Z(n23) );
  XOR U6026 ( .A(n24), .B(n6204), .Z(n6205) );
  XOR U6027 ( .A(n6206), .B(n6207), .Z(n6204) );
  AND U6028 ( .A(n42), .B(n6208), .Z(n6207) );
  XOR U6029 ( .A(n6209), .B(n6210), .Z(n24) );
  AND U6030 ( .A(n34), .B(n6211), .Z(n6210) );
  XOR U6031 ( .A(p_input[12]), .B(n6209), .Z(n6211) );
  XNOR U6032 ( .A(n6212), .B(n6213), .Z(n6209) );
  AND U6033 ( .A(n38), .B(n6208), .Z(n6213) );
  XNOR U6034 ( .A(n6212), .B(n6206), .Z(n6208) );
  XOR U6035 ( .A(n6214), .B(n6215), .Z(n6206) );
  AND U6036 ( .A(n54), .B(n6216), .Z(n6215) );
  XNOR U6037 ( .A(n6217), .B(n6218), .Z(n6212) );
  AND U6038 ( .A(n46), .B(n6219), .Z(n6218) );
  XOR U6039 ( .A(p_input[28]), .B(n6217), .Z(n6219) );
  XNOR U6040 ( .A(n6220), .B(n6221), .Z(n6217) );
  AND U6041 ( .A(n50), .B(n6216), .Z(n6221) );
  XNOR U6042 ( .A(n6220), .B(n6214), .Z(n6216) );
  XOR U6043 ( .A(n6222), .B(n6223), .Z(n6214) );
  AND U6044 ( .A(n65), .B(n6224), .Z(n6223) );
  XNOR U6045 ( .A(n6225), .B(n6226), .Z(n6220) );
  AND U6046 ( .A(n57), .B(n6227), .Z(n6226) );
  XOR U6047 ( .A(p_input[44]), .B(n6225), .Z(n6227) );
  XNOR U6048 ( .A(n6228), .B(n6229), .Z(n6225) );
  AND U6049 ( .A(n61), .B(n6224), .Z(n6229) );
  XNOR U6050 ( .A(n6228), .B(n6222), .Z(n6224) );
  XOR U6051 ( .A(n6230), .B(n6231), .Z(n6222) );
  AND U6052 ( .A(n76), .B(n6232), .Z(n6231) );
  XNOR U6053 ( .A(n6233), .B(n6234), .Z(n6228) );
  AND U6054 ( .A(n68), .B(n6235), .Z(n6234) );
  XOR U6055 ( .A(p_input[60]), .B(n6233), .Z(n6235) );
  XNOR U6056 ( .A(n6236), .B(n6237), .Z(n6233) );
  AND U6057 ( .A(n72), .B(n6232), .Z(n6237) );
  XNOR U6058 ( .A(n6236), .B(n6230), .Z(n6232) );
  XOR U6059 ( .A(n6238), .B(n6239), .Z(n6230) );
  AND U6060 ( .A(n87), .B(n6240), .Z(n6239) );
  XNOR U6061 ( .A(n6241), .B(n6242), .Z(n6236) );
  AND U6062 ( .A(n79), .B(n6243), .Z(n6242) );
  XOR U6063 ( .A(p_input[76]), .B(n6241), .Z(n6243) );
  XNOR U6064 ( .A(n6244), .B(n6245), .Z(n6241) );
  AND U6065 ( .A(n83), .B(n6240), .Z(n6245) );
  XNOR U6066 ( .A(n6244), .B(n6238), .Z(n6240) );
  XOR U6067 ( .A(n6246), .B(n6247), .Z(n6238) );
  AND U6068 ( .A(n98), .B(n6248), .Z(n6247) );
  XNOR U6069 ( .A(n6249), .B(n6250), .Z(n6244) );
  AND U6070 ( .A(n90), .B(n6251), .Z(n6250) );
  XOR U6071 ( .A(p_input[92]), .B(n6249), .Z(n6251) );
  XNOR U6072 ( .A(n6252), .B(n6253), .Z(n6249) );
  AND U6073 ( .A(n94), .B(n6248), .Z(n6253) );
  XNOR U6074 ( .A(n6252), .B(n6246), .Z(n6248) );
  XOR U6075 ( .A(n6254), .B(n6255), .Z(n6246) );
  AND U6076 ( .A(n109), .B(n6256), .Z(n6255) );
  XNOR U6077 ( .A(n6257), .B(n6258), .Z(n6252) );
  AND U6078 ( .A(n101), .B(n6259), .Z(n6258) );
  XOR U6079 ( .A(p_input[108]), .B(n6257), .Z(n6259) );
  XNOR U6080 ( .A(n6260), .B(n6261), .Z(n6257) );
  AND U6081 ( .A(n105), .B(n6256), .Z(n6261) );
  XNOR U6082 ( .A(n6260), .B(n6254), .Z(n6256) );
  XOR U6083 ( .A(n6262), .B(n6263), .Z(n6254) );
  AND U6084 ( .A(n120), .B(n6264), .Z(n6263) );
  XNOR U6085 ( .A(n6265), .B(n6266), .Z(n6260) );
  AND U6086 ( .A(n112), .B(n6267), .Z(n6266) );
  XOR U6087 ( .A(p_input[124]), .B(n6265), .Z(n6267) );
  XNOR U6088 ( .A(n6268), .B(n6269), .Z(n6265) );
  AND U6089 ( .A(n116), .B(n6264), .Z(n6269) );
  XNOR U6090 ( .A(n6268), .B(n6262), .Z(n6264) );
  XOR U6091 ( .A(n6270), .B(n6271), .Z(n6262) );
  AND U6092 ( .A(n131), .B(n6272), .Z(n6271) );
  XNOR U6093 ( .A(n6273), .B(n6274), .Z(n6268) );
  AND U6094 ( .A(n123), .B(n6275), .Z(n6274) );
  XOR U6095 ( .A(p_input[140]), .B(n6273), .Z(n6275) );
  XNOR U6096 ( .A(n6276), .B(n6277), .Z(n6273) );
  AND U6097 ( .A(n127), .B(n6272), .Z(n6277) );
  XNOR U6098 ( .A(n6276), .B(n6270), .Z(n6272) );
  XOR U6099 ( .A(n6278), .B(n6279), .Z(n6270) );
  AND U6100 ( .A(n142), .B(n6280), .Z(n6279) );
  XNOR U6101 ( .A(n6281), .B(n6282), .Z(n6276) );
  AND U6102 ( .A(n134), .B(n6283), .Z(n6282) );
  XOR U6103 ( .A(p_input[156]), .B(n6281), .Z(n6283) );
  XNOR U6104 ( .A(n6284), .B(n6285), .Z(n6281) );
  AND U6105 ( .A(n138), .B(n6280), .Z(n6285) );
  XNOR U6106 ( .A(n6284), .B(n6278), .Z(n6280) );
  XOR U6107 ( .A(n6286), .B(n6287), .Z(n6278) );
  AND U6108 ( .A(n153), .B(n6288), .Z(n6287) );
  XNOR U6109 ( .A(n6289), .B(n6290), .Z(n6284) );
  AND U6110 ( .A(n145), .B(n6291), .Z(n6290) );
  XOR U6111 ( .A(p_input[172]), .B(n6289), .Z(n6291) );
  XNOR U6112 ( .A(n6292), .B(n6293), .Z(n6289) );
  AND U6113 ( .A(n149), .B(n6288), .Z(n6293) );
  XNOR U6114 ( .A(n6292), .B(n6286), .Z(n6288) );
  XOR U6115 ( .A(n6294), .B(n6295), .Z(n6286) );
  AND U6116 ( .A(n164), .B(n6296), .Z(n6295) );
  XNOR U6117 ( .A(n6297), .B(n6298), .Z(n6292) );
  AND U6118 ( .A(n156), .B(n6299), .Z(n6298) );
  XOR U6119 ( .A(p_input[188]), .B(n6297), .Z(n6299) );
  XNOR U6120 ( .A(n6300), .B(n6301), .Z(n6297) );
  AND U6121 ( .A(n160), .B(n6296), .Z(n6301) );
  XNOR U6122 ( .A(n6300), .B(n6294), .Z(n6296) );
  XOR U6123 ( .A(n6302), .B(n6303), .Z(n6294) );
  AND U6124 ( .A(n175), .B(n6304), .Z(n6303) );
  XNOR U6125 ( .A(n6305), .B(n6306), .Z(n6300) );
  AND U6126 ( .A(n167), .B(n6307), .Z(n6306) );
  XOR U6127 ( .A(p_input[204]), .B(n6305), .Z(n6307) );
  XNOR U6128 ( .A(n6308), .B(n6309), .Z(n6305) );
  AND U6129 ( .A(n171), .B(n6304), .Z(n6309) );
  XNOR U6130 ( .A(n6308), .B(n6302), .Z(n6304) );
  XOR U6131 ( .A(n6310), .B(n6311), .Z(n6302) );
  AND U6132 ( .A(n186), .B(n6312), .Z(n6311) );
  XNOR U6133 ( .A(n6313), .B(n6314), .Z(n6308) );
  AND U6134 ( .A(n178), .B(n6315), .Z(n6314) );
  XOR U6135 ( .A(p_input[220]), .B(n6313), .Z(n6315) );
  XNOR U6136 ( .A(n6316), .B(n6317), .Z(n6313) );
  AND U6137 ( .A(n182), .B(n6312), .Z(n6317) );
  XNOR U6138 ( .A(n6316), .B(n6310), .Z(n6312) );
  XOR U6139 ( .A(n6318), .B(n6319), .Z(n6310) );
  AND U6140 ( .A(n197), .B(n6320), .Z(n6319) );
  XNOR U6141 ( .A(n6321), .B(n6322), .Z(n6316) );
  AND U6142 ( .A(n189), .B(n6323), .Z(n6322) );
  XOR U6143 ( .A(p_input[236]), .B(n6321), .Z(n6323) );
  XNOR U6144 ( .A(n6324), .B(n6325), .Z(n6321) );
  AND U6145 ( .A(n193), .B(n6320), .Z(n6325) );
  XNOR U6146 ( .A(n6324), .B(n6318), .Z(n6320) );
  XOR U6147 ( .A(n6326), .B(n6327), .Z(n6318) );
  AND U6148 ( .A(n208), .B(n6328), .Z(n6327) );
  XNOR U6149 ( .A(n6329), .B(n6330), .Z(n6324) );
  AND U6150 ( .A(n200), .B(n6331), .Z(n6330) );
  XOR U6151 ( .A(p_input[252]), .B(n6329), .Z(n6331) );
  XNOR U6152 ( .A(n6332), .B(n6333), .Z(n6329) );
  AND U6153 ( .A(n204), .B(n6328), .Z(n6333) );
  XNOR U6154 ( .A(n6332), .B(n6326), .Z(n6328) );
  XOR U6155 ( .A(n6334), .B(n6335), .Z(n6326) );
  AND U6156 ( .A(n219), .B(n6336), .Z(n6335) );
  XNOR U6157 ( .A(n6337), .B(n6338), .Z(n6332) );
  AND U6158 ( .A(n211), .B(n6339), .Z(n6338) );
  XOR U6159 ( .A(p_input[268]), .B(n6337), .Z(n6339) );
  XNOR U6160 ( .A(n6340), .B(n6341), .Z(n6337) );
  AND U6161 ( .A(n215), .B(n6336), .Z(n6341) );
  XNOR U6162 ( .A(n6340), .B(n6334), .Z(n6336) );
  XOR U6163 ( .A(n6342), .B(n6343), .Z(n6334) );
  AND U6164 ( .A(n230), .B(n6344), .Z(n6343) );
  XNOR U6165 ( .A(n6345), .B(n6346), .Z(n6340) );
  AND U6166 ( .A(n222), .B(n6347), .Z(n6346) );
  XOR U6167 ( .A(p_input[284]), .B(n6345), .Z(n6347) );
  XNOR U6168 ( .A(n6348), .B(n6349), .Z(n6345) );
  AND U6169 ( .A(n226), .B(n6344), .Z(n6349) );
  XNOR U6170 ( .A(n6348), .B(n6342), .Z(n6344) );
  XOR U6171 ( .A(n6350), .B(n6351), .Z(n6342) );
  AND U6172 ( .A(n241), .B(n6352), .Z(n6351) );
  XNOR U6173 ( .A(n6353), .B(n6354), .Z(n6348) );
  AND U6174 ( .A(n233), .B(n6355), .Z(n6354) );
  XOR U6175 ( .A(p_input[300]), .B(n6353), .Z(n6355) );
  XNOR U6176 ( .A(n6356), .B(n6357), .Z(n6353) );
  AND U6177 ( .A(n237), .B(n6352), .Z(n6357) );
  XNOR U6178 ( .A(n6356), .B(n6350), .Z(n6352) );
  XOR U6179 ( .A(n6358), .B(n6359), .Z(n6350) );
  AND U6180 ( .A(n252), .B(n6360), .Z(n6359) );
  XNOR U6181 ( .A(n6361), .B(n6362), .Z(n6356) );
  AND U6182 ( .A(n244), .B(n6363), .Z(n6362) );
  XOR U6183 ( .A(p_input[316]), .B(n6361), .Z(n6363) );
  XNOR U6184 ( .A(n6364), .B(n6365), .Z(n6361) );
  AND U6185 ( .A(n248), .B(n6360), .Z(n6365) );
  XNOR U6186 ( .A(n6364), .B(n6358), .Z(n6360) );
  XOR U6187 ( .A(n6366), .B(n6367), .Z(n6358) );
  AND U6188 ( .A(n263), .B(n6368), .Z(n6367) );
  XNOR U6189 ( .A(n6369), .B(n6370), .Z(n6364) );
  AND U6190 ( .A(n255), .B(n6371), .Z(n6370) );
  XOR U6191 ( .A(p_input[332]), .B(n6369), .Z(n6371) );
  XNOR U6192 ( .A(n6372), .B(n6373), .Z(n6369) );
  AND U6193 ( .A(n259), .B(n6368), .Z(n6373) );
  XNOR U6194 ( .A(n6372), .B(n6366), .Z(n6368) );
  XOR U6195 ( .A(n6374), .B(n6375), .Z(n6366) );
  AND U6196 ( .A(n274), .B(n6376), .Z(n6375) );
  XNOR U6197 ( .A(n6377), .B(n6378), .Z(n6372) );
  AND U6198 ( .A(n266), .B(n6379), .Z(n6378) );
  XOR U6199 ( .A(p_input[348]), .B(n6377), .Z(n6379) );
  XNOR U6200 ( .A(n6380), .B(n6381), .Z(n6377) );
  AND U6201 ( .A(n270), .B(n6376), .Z(n6381) );
  XNOR U6202 ( .A(n6380), .B(n6374), .Z(n6376) );
  XOR U6203 ( .A(n6382), .B(n6383), .Z(n6374) );
  AND U6204 ( .A(n285), .B(n6384), .Z(n6383) );
  XNOR U6205 ( .A(n6385), .B(n6386), .Z(n6380) );
  AND U6206 ( .A(n277), .B(n6387), .Z(n6386) );
  XOR U6207 ( .A(p_input[364]), .B(n6385), .Z(n6387) );
  XNOR U6208 ( .A(n6388), .B(n6389), .Z(n6385) );
  AND U6209 ( .A(n281), .B(n6384), .Z(n6389) );
  XNOR U6210 ( .A(n6388), .B(n6382), .Z(n6384) );
  XOR U6211 ( .A(n6390), .B(n6391), .Z(n6382) );
  AND U6212 ( .A(n296), .B(n6392), .Z(n6391) );
  XNOR U6213 ( .A(n6393), .B(n6394), .Z(n6388) );
  AND U6214 ( .A(n288), .B(n6395), .Z(n6394) );
  XOR U6215 ( .A(p_input[380]), .B(n6393), .Z(n6395) );
  XNOR U6216 ( .A(n6396), .B(n6397), .Z(n6393) );
  AND U6217 ( .A(n292), .B(n6392), .Z(n6397) );
  XNOR U6218 ( .A(n6396), .B(n6390), .Z(n6392) );
  XOR U6219 ( .A(n6398), .B(n6399), .Z(n6390) );
  AND U6220 ( .A(n307), .B(n6400), .Z(n6399) );
  XNOR U6221 ( .A(n6401), .B(n6402), .Z(n6396) );
  AND U6222 ( .A(n299), .B(n6403), .Z(n6402) );
  XOR U6223 ( .A(p_input[396]), .B(n6401), .Z(n6403) );
  XNOR U6224 ( .A(n6404), .B(n6405), .Z(n6401) );
  AND U6225 ( .A(n303), .B(n6400), .Z(n6405) );
  XNOR U6226 ( .A(n6404), .B(n6398), .Z(n6400) );
  XOR U6227 ( .A(n6406), .B(n6407), .Z(n6398) );
  AND U6228 ( .A(n318), .B(n6408), .Z(n6407) );
  XNOR U6229 ( .A(n6409), .B(n6410), .Z(n6404) );
  AND U6230 ( .A(n310), .B(n6411), .Z(n6410) );
  XOR U6231 ( .A(p_input[412]), .B(n6409), .Z(n6411) );
  XNOR U6232 ( .A(n6412), .B(n6413), .Z(n6409) );
  AND U6233 ( .A(n314), .B(n6408), .Z(n6413) );
  XNOR U6234 ( .A(n6412), .B(n6406), .Z(n6408) );
  XOR U6235 ( .A(n6414), .B(n6415), .Z(n6406) );
  AND U6236 ( .A(n329), .B(n6416), .Z(n6415) );
  XNOR U6237 ( .A(n6417), .B(n6418), .Z(n6412) );
  AND U6238 ( .A(n321), .B(n6419), .Z(n6418) );
  XOR U6239 ( .A(p_input[428]), .B(n6417), .Z(n6419) );
  XNOR U6240 ( .A(n6420), .B(n6421), .Z(n6417) );
  AND U6241 ( .A(n325), .B(n6416), .Z(n6421) );
  XNOR U6242 ( .A(n6420), .B(n6414), .Z(n6416) );
  XOR U6243 ( .A(n6422), .B(n6423), .Z(n6414) );
  AND U6244 ( .A(n340), .B(n6424), .Z(n6423) );
  XNOR U6245 ( .A(n6425), .B(n6426), .Z(n6420) );
  AND U6246 ( .A(n332), .B(n6427), .Z(n6426) );
  XOR U6247 ( .A(p_input[444]), .B(n6425), .Z(n6427) );
  XNOR U6248 ( .A(n6428), .B(n6429), .Z(n6425) );
  AND U6249 ( .A(n336), .B(n6424), .Z(n6429) );
  XNOR U6250 ( .A(n6428), .B(n6422), .Z(n6424) );
  XOR U6251 ( .A(n6430), .B(n6431), .Z(n6422) );
  AND U6252 ( .A(n351), .B(n6432), .Z(n6431) );
  XNOR U6253 ( .A(n6433), .B(n6434), .Z(n6428) );
  AND U6254 ( .A(n343), .B(n6435), .Z(n6434) );
  XOR U6255 ( .A(p_input[460]), .B(n6433), .Z(n6435) );
  XNOR U6256 ( .A(n6436), .B(n6437), .Z(n6433) );
  AND U6257 ( .A(n347), .B(n6432), .Z(n6437) );
  XNOR U6258 ( .A(n6436), .B(n6430), .Z(n6432) );
  XOR U6259 ( .A(n6438), .B(n6439), .Z(n6430) );
  AND U6260 ( .A(n362), .B(n6440), .Z(n6439) );
  XNOR U6261 ( .A(n6441), .B(n6442), .Z(n6436) );
  AND U6262 ( .A(n354), .B(n6443), .Z(n6442) );
  XOR U6263 ( .A(p_input[476]), .B(n6441), .Z(n6443) );
  XNOR U6264 ( .A(n6444), .B(n6445), .Z(n6441) );
  AND U6265 ( .A(n358), .B(n6440), .Z(n6445) );
  XNOR U6266 ( .A(n6444), .B(n6438), .Z(n6440) );
  XOR U6267 ( .A(n6446), .B(n6447), .Z(n6438) );
  AND U6268 ( .A(n373), .B(n6448), .Z(n6447) );
  XNOR U6269 ( .A(n6449), .B(n6450), .Z(n6444) );
  AND U6270 ( .A(n365), .B(n6451), .Z(n6450) );
  XOR U6271 ( .A(p_input[492]), .B(n6449), .Z(n6451) );
  XNOR U6272 ( .A(n6452), .B(n6453), .Z(n6449) );
  AND U6273 ( .A(n369), .B(n6448), .Z(n6453) );
  XNOR U6274 ( .A(n6452), .B(n6446), .Z(n6448) );
  XOR U6275 ( .A(n6454), .B(n6455), .Z(n6446) );
  AND U6276 ( .A(n384), .B(n6456), .Z(n6455) );
  XNOR U6277 ( .A(n6457), .B(n6458), .Z(n6452) );
  AND U6278 ( .A(n376), .B(n6459), .Z(n6458) );
  XOR U6279 ( .A(p_input[508]), .B(n6457), .Z(n6459) );
  XNOR U6280 ( .A(n6460), .B(n6461), .Z(n6457) );
  AND U6281 ( .A(n380), .B(n6456), .Z(n6461) );
  XNOR U6282 ( .A(n6460), .B(n6454), .Z(n6456) );
  XOR U6283 ( .A(n6462), .B(n6463), .Z(n6454) );
  AND U6284 ( .A(n395), .B(n6464), .Z(n6463) );
  XNOR U6285 ( .A(n6465), .B(n6466), .Z(n6460) );
  AND U6286 ( .A(n387), .B(n6467), .Z(n6466) );
  XOR U6287 ( .A(p_input[524]), .B(n6465), .Z(n6467) );
  XNOR U6288 ( .A(n6468), .B(n6469), .Z(n6465) );
  AND U6289 ( .A(n391), .B(n6464), .Z(n6469) );
  XNOR U6290 ( .A(n6468), .B(n6462), .Z(n6464) );
  XOR U6291 ( .A(n6470), .B(n6471), .Z(n6462) );
  AND U6292 ( .A(n406), .B(n6472), .Z(n6471) );
  XNOR U6293 ( .A(n6473), .B(n6474), .Z(n6468) );
  AND U6294 ( .A(n398), .B(n6475), .Z(n6474) );
  XOR U6295 ( .A(p_input[540]), .B(n6473), .Z(n6475) );
  XNOR U6296 ( .A(n6476), .B(n6477), .Z(n6473) );
  AND U6297 ( .A(n402), .B(n6472), .Z(n6477) );
  XNOR U6298 ( .A(n6476), .B(n6470), .Z(n6472) );
  XOR U6299 ( .A(n6478), .B(n6479), .Z(n6470) );
  AND U6300 ( .A(n417), .B(n6480), .Z(n6479) );
  XNOR U6301 ( .A(n6481), .B(n6482), .Z(n6476) );
  AND U6302 ( .A(n409), .B(n6483), .Z(n6482) );
  XOR U6303 ( .A(p_input[556]), .B(n6481), .Z(n6483) );
  XNOR U6304 ( .A(n6484), .B(n6485), .Z(n6481) );
  AND U6305 ( .A(n413), .B(n6480), .Z(n6485) );
  XNOR U6306 ( .A(n6484), .B(n6478), .Z(n6480) );
  XOR U6307 ( .A(n6486), .B(n6487), .Z(n6478) );
  AND U6308 ( .A(n428), .B(n6488), .Z(n6487) );
  XNOR U6309 ( .A(n6489), .B(n6490), .Z(n6484) );
  AND U6310 ( .A(n420), .B(n6491), .Z(n6490) );
  XOR U6311 ( .A(p_input[572]), .B(n6489), .Z(n6491) );
  XNOR U6312 ( .A(n6492), .B(n6493), .Z(n6489) );
  AND U6313 ( .A(n424), .B(n6488), .Z(n6493) );
  XNOR U6314 ( .A(n6492), .B(n6486), .Z(n6488) );
  XOR U6315 ( .A(n6494), .B(n6495), .Z(n6486) );
  AND U6316 ( .A(n439), .B(n6496), .Z(n6495) );
  XNOR U6317 ( .A(n6497), .B(n6498), .Z(n6492) );
  AND U6318 ( .A(n431), .B(n6499), .Z(n6498) );
  XOR U6319 ( .A(p_input[588]), .B(n6497), .Z(n6499) );
  XNOR U6320 ( .A(n6500), .B(n6501), .Z(n6497) );
  AND U6321 ( .A(n435), .B(n6496), .Z(n6501) );
  XNOR U6322 ( .A(n6500), .B(n6494), .Z(n6496) );
  XOR U6323 ( .A(n6502), .B(n6503), .Z(n6494) );
  AND U6324 ( .A(n450), .B(n6504), .Z(n6503) );
  XNOR U6325 ( .A(n6505), .B(n6506), .Z(n6500) );
  AND U6326 ( .A(n442), .B(n6507), .Z(n6506) );
  XOR U6327 ( .A(p_input[604]), .B(n6505), .Z(n6507) );
  XNOR U6328 ( .A(n6508), .B(n6509), .Z(n6505) );
  AND U6329 ( .A(n446), .B(n6504), .Z(n6509) );
  XNOR U6330 ( .A(n6508), .B(n6502), .Z(n6504) );
  XOR U6331 ( .A(n6510), .B(n6511), .Z(n6502) );
  AND U6332 ( .A(n461), .B(n6512), .Z(n6511) );
  XNOR U6333 ( .A(n6513), .B(n6514), .Z(n6508) );
  AND U6334 ( .A(n453), .B(n6515), .Z(n6514) );
  XOR U6335 ( .A(p_input[620]), .B(n6513), .Z(n6515) );
  XNOR U6336 ( .A(n6516), .B(n6517), .Z(n6513) );
  AND U6337 ( .A(n457), .B(n6512), .Z(n6517) );
  XNOR U6338 ( .A(n6516), .B(n6510), .Z(n6512) );
  XOR U6339 ( .A(n6518), .B(n6519), .Z(n6510) );
  AND U6340 ( .A(n472), .B(n6520), .Z(n6519) );
  XNOR U6341 ( .A(n6521), .B(n6522), .Z(n6516) );
  AND U6342 ( .A(n464), .B(n6523), .Z(n6522) );
  XOR U6343 ( .A(p_input[636]), .B(n6521), .Z(n6523) );
  XNOR U6344 ( .A(n6524), .B(n6525), .Z(n6521) );
  AND U6345 ( .A(n468), .B(n6520), .Z(n6525) );
  XNOR U6346 ( .A(n6524), .B(n6518), .Z(n6520) );
  XOR U6347 ( .A(n6526), .B(n6527), .Z(n6518) );
  AND U6348 ( .A(n483), .B(n6528), .Z(n6527) );
  XNOR U6349 ( .A(n6529), .B(n6530), .Z(n6524) );
  AND U6350 ( .A(n475), .B(n6531), .Z(n6530) );
  XOR U6351 ( .A(p_input[652]), .B(n6529), .Z(n6531) );
  XNOR U6352 ( .A(n6532), .B(n6533), .Z(n6529) );
  AND U6353 ( .A(n479), .B(n6528), .Z(n6533) );
  XNOR U6354 ( .A(n6532), .B(n6526), .Z(n6528) );
  XOR U6355 ( .A(n6534), .B(n6535), .Z(n6526) );
  AND U6356 ( .A(n494), .B(n6536), .Z(n6535) );
  XNOR U6357 ( .A(n6537), .B(n6538), .Z(n6532) );
  AND U6358 ( .A(n486), .B(n6539), .Z(n6538) );
  XOR U6359 ( .A(p_input[668]), .B(n6537), .Z(n6539) );
  XNOR U6360 ( .A(n6540), .B(n6541), .Z(n6537) );
  AND U6361 ( .A(n490), .B(n6536), .Z(n6541) );
  XNOR U6362 ( .A(n6540), .B(n6534), .Z(n6536) );
  XOR U6363 ( .A(n6542), .B(n6543), .Z(n6534) );
  AND U6364 ( .A(n505), .B(n6544), .Z(n6543) );
  XNOR U6365 ( .A(n6545), .B(n6546), .Z(n6540) );
  AND U6366 ( .A(n497), .B(n6547), .Z(n6546) );
  XOR U6367 ( .A(p_input[684]), .B(n6545), .Z(n6547) );
  XNOR U6368 ( .A(n6548), .B(n6549), .Z(n6545) );
  AND U6369 ( .A(n501), .B(n6544), .Z(n6549) );
  XNOR U6370 ( .A(n6548), .B(n6542), .Z(n6544) );
  XOR U6371 ( .A(n6550), .B(n6551), .Z(n6542) );
  AND U6372 ( .A(n516), .B(n6552), .Z(n6551) );
  XNOR U6373 ( .A(n6553), .B(n6554), .Z(n6548) );
  AND U6374 ( .A(n508), .B(n6555), .Z(n6554) );
  XOR U6375 ( .A(p_input[700]), .B(n6553), .Z(n6555) );
  XNOR U6376 ( .A(n6556), .B(n6557), .Z(n6553) );
  AND U6377 ( .A(n512), .B(n6552), .Z(n6557) );
  XNOR U6378 ( .A(n6556), .B(n6550), .Z(n6552) );
  XOR U6379 ( .A(n6558), .B(n6559), .Z(n6550) );
  AND U6380 ( .A(n527), .B(n6560), .Z(n6559) );
  XNOR U6381 ( .A(n6561), .B(n6562), .Z(n6556) );
  AND U6382 ( .A(n519), .B(n6563), .Z(n6562) );
  XOR U6383 ( .A(p_input[716]), .B(n6561), .Z(n6563) );
  XNOR U6384 ( .A(n6564), .B(n6565), .Z(n6561) );
  AND U6385 ( .A(n523), .B(n6560), .Z(n6565) );
  XNOR U6386 ( .A(n6564), .B(n6558), .Z(n6560) );
  XOR U6387 ( .A(n6566), .B(n6567), .Z(n6558) );
  AND U6388 ( .A(n538), .B(n6568), .Z(n6567) );
  XNOR U6389 ( .A(n6569), .B(n6570), .Z(n6564) );
  AND U6390 ( .A(n530), .B(n6571), .Z(n6570) );
  XOR U6391 ( .A(p_input[732]), .B(n6569), .Z(n6571) );
  XNOR U6392 ( .A(n6572), .B(n6573), .Z(n6569) );
  AND U6393 ( .A(n534), .B(n6568), .Z(n6573) );
  XNOR U6394 ( .A(n6572), .B(n6566), .Z(n6568) );
  XOR U6395 ( .A(n6574), .B(n6575), .Z(n6566) );
  AND U6396 ( .A(n549), .B(n6576), .Z(n6575) );
  XNOR U6397 ( .A(n6577), .B(n6578), .Z(n6572) );
  AND U6398 ( .A(n541), .B(n6579), .Z(n6578) );
  XOR U6399 ( .A(p_input[748]), .B(n6577), .Z(n6579) );
  XNOR U6400 ( .A(n6580), .B(n6581), .Z(n6577) );
  AND U6401 ( .A(n545), .B(n6576), .Z(n6581) );
  XNOR U6402 ( .A(n6580), .B(n6574), .Z(n6576) );
  XOR U6403 ( .A(n6582), .B(n6583), .Z(n6574) );
  AND U6404 ( .A(n560), .B(n6584), .Z(n6583) );
  XNOR U6405 ( .A(n6585), .B(n6586), .Z(n6580) );
  AND U6406 ( .A(n552), .B(n6587), .Z(n6586) );
  XOR U6407 ( .A(p_input[764]), .B(n6585), .Z(n6587) );
  XNOR U6408 ( .A(n6588), .B(n6589), .Z(n6585) );
  AND U6409 ( .A(n556), .B(n6584), .Z(n6589) );
  XNOR U6410 ( .A(n6588), .B(n6582), .Z(n6584) );
  XOR U6411 ( .A(n6590), .B(n6591), .Z(n6582) );
  AND U6412 ( .A(n571), .B(n6592), .Z(n6591) );
  XNOR U6413 ( .A(n6593), .B(n6594), .Z(n6588) );
  AND U6414 ( .A(n563), .B(n6595), .Z(n6594) );
  XOR U6415 ( .A(p_input[780]), .B(n6593), .Z(n6595) );
  XNOR U6416 ( .A(n6596), .B(n6597), .Z(n6593) );
  AND U6417 ( .A(n567), .B(n6592), .Z(n6597) );
  XNOR U6418 ( .A(n6596), .B(n6590), .Z(n6592) );
  XOR U6419 ( .A(n6598), .B(n6599), .Z(n6590) );
  AND U6420 ( .A(n582), .B(n6600), .Z(n6599) );
  XNOR U6421 ( .A(n6601), .B(n6602), .Z(n6596) );
  AND U6422 ( .A(n574), .B(n6603), .Z(n6602) );
  XOR U6423 ( .A(p_input[796]), .B(n6601), .Z(n6603) );
  XNOR U6424 ( .A(n6604), .B(n6605), .Z(n6601) );
  AND U6425 ( .A(n578), .B(n6600), .Z(n6605) );
  XNOR U6426 ( .A(n6604), .B(n6598), .Z(n6600) );
  XOR U6427 ( .A(n6606), .B(n6607), .Z(n6598) );
  AND U6428 ( .A(n593), .B(n6608), .Z(n6607) );
  XNOR U6429 ( .A(n6609), .B(n6610), .Z(n6604) );
  AND U6430 ( .A(n585), .B(n6611), .Z(n6610) );
  XOR U6431 ( .A(p_input[812]), .B(n6609), .Z(n6611) );
  XNOR U6432 ( .A(n6612), .B(n6613), .Z(n6609) );
  AND U6433 ( .A(n589), .B(n6608), .Z(n6613) );
  XNOR U6434 ( .A(n6612), .B(n6606), .Z(n6608) );
  XOR U6435 ( .A(n6614), .B(n6615), .Z(n6606) );
  AND U6436 ( .A(n604), .B(n6616), .Z(n6615) );
  XNOR U6437 ( .A(n6617), .B(n6618), .Z(n6612) );
  AND U6438 ( .A(n596), .B(n6619), .Z(n6618) );
  XOR U6439 ( .A(p_input[828]), .B(n6617), .Z(n6619) );
  XNOR U6440 ( .A(n6620), .B(n6621), .Z(n6617) );
  AND U6441 ( .A(n600), .B(n6616), .Z(n6621) );
  XNOR U6442 ( .A(n6620), .B(n6614), .Z(n6616) );
  XOR U6443 ( .A(n6622), .B(n6623), .Z(n6614) );
  AND U6444 ( .A(n615), .B(n6624), .Z(n6623) );
  XNOR U6445 ( .A(n6625), .B(n6626), .Z(n6620) );
  AND U6446 ( .A(n607), .B(n6627), .Z(n6626) );
  XOR U6447 ( .A(p_input[844]), .B(n6625), .Z(n6627) );
  XNOR U6448 ( .A(n6628), .B(n6629), .Z(n6625) );
  AND U6449 ( .A(n611), .B(n6624), .Z(n6629) );
  XNOR U6450 ( .A(n6628), .B(n6622), .Z(n6624) );
  XOR U6451 ( .A(n6630), .B(n6631), .Z(n6622) );
  AND U6452 ( .A(n626), .B(n6632), .Z(n6631) );
  XNOR U6453 ( .A(n6633), .B(n6634), .Z(n6628) );
  AND U6454 ( .A(n618), .B(n6635), .Z(n6634) );
  XOR U6455 ( .A(p_input[860]), .B(n6633), .Z(n6635) );
  XNOR U6456 ( .A(n6636), .B(n6637), .Z(n6633) );
  AND U6457 ( .A(n622), .B(n6632), .Z(n6637) );
  XNOR U6458 ( .A(n6636), .B(n6630), .Z(n6632) );
  XOR U6459 ( .A(n6638), .B(n6639), .Z(n6630) );
  AND U6460 ( .A(n637), .B(n6640), .Z(n6639) );
  XNOR U6461 ( .A(n6641), .B(n6642), .Z(n6636) );
  AND U6462 ( .A(n629), .B(n6643), .Z(n6642) );
  XOR U6463 ( .A(p_input[876]), .B(n6641), .Z(n6643) );
  XNOR U6464 ( .A(n6644), .B(n6645), .Z(n6641) );
  AND U6465 ( .A(n633), .B(n6640), .Z(n6645) );
  XNOR U6466 ( .A(n6644), .B(n6638), .Z(n6640) );
  XOR U6467 ( .A(n6646), .B(n6647), .Z(n6638) );
  AND U6468 ( .A(n648), .B(n6648), .Z(n6647) );
  XNOR U6469 ( .A(n6649), .B(n6650), .Z(n6644) );
  AND U6470 ( .A(n640), .B(n6651), .Z(n6650) );
  XOR U6471 ( .A(p_input[892]), .B(n6649), .Z(n6651) );
  XNOR U6472 ( .A(n6652), .B(n6653), .Z(n6649) );
  AND U6473 ( .A(n644), .B(n6648), .Z(n6653) );
  XNOR U6474 ( .A(n6652), .B(n6646), .Z(n6648) );
  XOR U6475 ( .A(n6654), .B(n6655), .Z(n6646) );
  AND U6476 ( .A(n659), .B(n6656), .Z(n6655) );
  XNOR U6477 ( .A(n6657), .B(n6658), .Z(n6652) );
  AND U6478 ( .A(n651), .B(n6659), .Z(n6658) );
  XOR U6479 ( .A(p_input[908]), .B(n6657), .Z(n6659) );
  XNOR U6480 ( .A(n6660), .B(n6661), .Z(n6657) );
  AND U6481 ( .A(n655), .B(n6656), .Z(n6661) );
  XNOR U6482 ( .A(n6660), .B(n6654), .Z(n6656) );
  XOR U6483 ( .A(n6662), .B(n6663), .Z(n6654) );
  AND U6484 ( .A(n670), .B(n6664), .Z(n6663) );
  XNOR U6485 ( .A(n6665), .B(n6666), .Z(n6660) );
  AND U6486 ( .A(n662), .B(n6667), .Z(n6666) );
  XOR U6487 ( .A(p_input[924]), .B(n6665), .Z(n6667) );
  XNOR U6488 ( .A(n6668), .B(n6669), .Z(n6665) );
  AND U6489 ( .A(n666), .B(n6664), .Z(n6669) );
  XNOR U6490 ( .A(n6668), .B(n6662), .Z(n6664) );
  XOR U6491 ( .A(n6670), .B(n6671), .Z(n6662) );
  AND U6492 ( .A(n681), .B(n6672), .Z(n6671) );
  XNOR U6493 ( .A(n6673), .B(n6674), .Z(n6668) );
  AND U6494 ( .A(n673), .B(n6675), .Z(n6674) );
  XOR U6495 ( .A(p_input[940]), .B(n6673), .Z(n6675) );
  XNOR U6496 ( .A(n6676), .B(n6677), .Z(n6673) );
  AND U6497 ( .A(n677), .B(n6672), .Z(n6677) );
  XNOR U6498 ( .A(n6676), .B(n6670), .Z(n6672) );
  XOR U6499 ( .A(n6678), .B(n6679), .Z(n6670) );
  AND U6500 ( .A(n692), .B(n6680), .Z(n6679) );
  XNOR U6501 ( .A(n6681), .B(n6682), .Z(n6676) );
  AND U6502 ( .A(n684), .B(n6683), .Z(n6682) );
  XOR U6503 ( .A(p_input[956]), .B(n6681), .Z(n6683) );
  XNOR U6504 ( .A(n6684), .B(n6685), .Z(n6681) );
  AND U6505 ( .A(n688), .B(n6680), .Z(n6685) );
  XNOR U6506 ( .A(n6684), .B(n6678), .Z(n6680) );
  XOR U6507 ( .A(n6686), .B(n6687), .Z(n6678) );
  AND U6508 ( .A(n703), .B(n6688), .Z(n6687) );
  XNOR U6509 ( .A(n6689), .B(n6690), .Z(n6684) );
  AND U6510 ( .A(n695), .B(n6691), .Z(n6690) );
  XOR U6511 ( .A(p_input[972]), .B(n6689), .Z(n6691) );
  XNOR U6512 ( .A(n6692), .B(n6693), .Z(n6689) );
  AND U6513 ( .A(n699), .B(n6688), .Z(n6693) );
  XNOR U6514 ( .A(n6692), .B(n6686), .Z(n6688) );
  XOR U6515 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n6694), .Z(n6686) );
  AND U6516 ( .A(n713), .B(n6695), .Z(n6694) );
  XNOR U6517 ( .A(n6696), .B(n6697), .Z(n6692) );
  AND U6518 ( .A(n706), .B(n6698), .Z(n6697) );
  XOR U6519 ( .A(p_input[988]), .B(n6696), .Z(n6698) );
  XNOR U6520 ( .A(n6699), .B(n6700), .Z(n6696) );
  AND U6521 ( .A(n710), .B(n6695), .Z(n6700) );
  XOR U6522 ( .A(\knn_comb_/min_val_out[0][12] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n6695) );
  IV U6523 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n6699) );
  XOR U6524 ( .A(n25), .B(n6701), .Z(o[11]) );
  AND U6525 ( .A(n30), .B(n6702), .Z(n25) );
  XOR U6526 ( .A(n26), .B(n6701), .Z(n6702) );
  XOR U6527 ( .A(n6703), .B(n6704), .Z(n6701) );
  AND U6528 ( .A(n42), .B(n6705), .Z(n6704) );
  XOR U6529 ( .A(n6706), .B(n6707), .Z(n26) );
  AND U6530 ( .A(n34), .B(n6708), .Z(n6707) );
  XOR U6531 ( .A(p_input[11]), .B(n6706), .Z(n6708) );
  XNOR U6532 ( .A(n6709), .B(n6710), .Z(n6706) );
  AND U6533 ( .A(n38), .B(n6705), .Z(n6710) );
  XNOR U6534 ( .A(n6709), .B(n6703), .Z(n6705) );
  XOR U6535 ( .A(n6711), .B(n6712), .Z(n6703) );
  AND U6536 ( .A(n54), .B(n6713), .Z(n6712) );
  XNOR U6537 ( .A(n6714), .B(n6715), .Z(n6709) );
  AND U6538 ( .A(n46), .B(n6716), .Z(n6715) );
  XOR U6539 ( .A(p_input[27]), .B(n6714), .Z(n6716) );
  XNOR U6540 ( .A(n6717), .B(n6718), .Z(n6714) );
  AND U6541 ( .A(n50), .B(n6713), .Z(n6718) );
  XNOR U6542 ( .A(n6717), .B(n6711), .Z(n6713) );
  XOR U6543 ( .A(n6719), .B(n6720), .Z(n6711) );
  AND U6544 ( .A(n65), .B(n6721), .Z(n6720) );
  XNOR U6545 ( .A(n6722), .B(n6723), .Z(n6717) );
  AND U6546 ( .A(n57), .B(n6724), .Z(n6723) );
  XOR U6547 ( .A(p_input[43]), .B(n6722), .Z(n6724) );
  XNOR U6548 ( .A(n6725), .B(n6726), .Z(n6722) );
  AND U6549 ( .A(n61), .B(n6721), .Z(n6726) );
  XNOR U6550 ( .A(n6725), .B(n6719), .Z(n6721) );
  XOR U6551 ( .A(n6727), .B(n6728), .Z(n6719) );
  AND U6552 ( .A(n76), .B(n6729), .Z(n6728) );
  XNOR U6553 ( .A(n6730), .B(n6731), .Z(n6725) );
  AND U6554 ( .A(n68), .B(n6732), .Z(n6731) );
  XOR U6555 ( .A(p_input[59]), .B(n6730), .Z(n6732) );
  XNOR U6556 ( .A(n6733), .B(n6734), .Z(n6730) );
  AND U6557 ( .A(n72), .B(n6729), .Z(n6734) );
  XNOR U6558 ( .A(n6733), .B(n6727), .Z(n6729) );
  XOR U6559 ( .A(n6735), .B(n6736), .Z(n6727) );
  AND U6560 ( .A(n87), .B(n6737), .Z(n6736) );
  XNOR U6561 ( .A(n6738), .B(n6739), .Z(n6733) );
  AND U6562 ( .A(n79), .B(n6740), .Z(n6739) );
  XOR U6563 ( .A(p_input[75]), .B(n6738), .Z(n6740) );
  XNOR U6564 ( .A(n6741), .B(n6742), .Z(n6738) );
  AND U6565 ( .A(n83), .B(n6737), .Z(n6742) );
  XNOR U6566 ( .A(n6741), .B(n6735), .Z(n6737) );
  XOR U6567 ( .A(n6743), .B(n6744), .Z(n6735) );
  AND U6568 ( .A(n98), .B(n6745), .Z(n6744) );
  XNOR U6569 ( .A(n6746), .B(n6747), .Z(n6741) );
  AND U6570 ( .A(n90), .B(n6748), .Z(n6747) );
  XOR U6571 ( .A(p_input[91]), .B(n6746), .Z(n6748) );
  XNOR U6572 ( .A(n6749), .B(n6750), .Z(n6746) );
  AND U6573 ( .A(n94), .B(n6745), .Z(n6750) );
  XNOR U6574 ( .A(n6749), .B(n6743), .Z(n6745) );
  XOR U6575 ( .A(n6751), .B(n6752), .Z(n6743) );
  AND U6576 ( .A(n109), .B(n6753), .Z(n6752) );
  XNOR U6577 ( .A(n6754), .B(n6755), .Z(n6749) );
  AND U6578 ( .A(n101), .B(n6756), .Z(n6755) );
  XOR U6579 ( .A(p_input[107]), .B(n6754), .Z(n6756) );
  XNOR U6580 ( .A(n6757), .B(n6758), .Z(n6754) );
  AND U6581 ( .A(n105), .B(n6753), .Z(n6758) );
  XNOR U6582 ( .A(n6757), .B(n6751), .Z(n6753) );
  XOR U6583 ( .A(n6759), .B(n6760), .Z(n6751) );
  AND U6584 ( .A(n120), .B(n6761), .Z(n6760) );
  XNOR U6585 ( .A(n6762), .B(n6763), .Z(n6757) );
  AND U6586 ( .A(n112), .B(n6764), .Z(n6763) );
  XOR U6587 ( .A(p_input[123]), .B(n6762), .Z(n6764) );
  XNOR U6588 ( .A(n6765), .B(n6766), .Z(n6762) );
  AND U6589 ( .A(n116), .B(n6761), .Z(n6766) );
  XNOR U6590 ( .A(n6765), .B(n6759), .Z(n6761) );
  XOR U6591 ( .A(n6767), .B(n6768), .Z(n6759) );
  AND U6592 ( .A(n131), .B(n6769), .Z(n6768) );
  XNOR U6593 ( .A(n6770), .B(n6771), .Z(n6765) );
  AND U6594 ( .A(n123), .B(n6772), .Z(n6771) );
  XOR U6595 ( .A(p_input[139]), .B(n6770), .Z(n6772) );
  XNOR U6596 ( .A(n6773), .B(n6774), .Z(n6770) );
  AND U6597 ( .A(n127), .B(n6769), .Z(n6774) );
  XNOR U6598 ( .A(n6773), .B(n6767), .Z(n6769) );
  XOR U6599 ( .A(n6775), .B(n6776), .Z(n6767) );
  AND U6600 ( .A(n142), .B(n6777), .Z(n6776) );
  XNOR U6601 ( .A(n6778), .B(n6779), .Z(n6773) );
  AND U6602 ( .A(n134), .B(n6780), .Z(n6779) );
  XOR U6603 ( .A(p_input[155]), .B(n6778), .Z(n6780) );
  XNOR U6604 ( .A(n6781), .B(n6782), .Z(n6778) );
  AND U6605 ( .A(n138), .B(n6777), .Z(n6782) );
  XNOR U6606 ( .A(n6781), .B(n6775), .Z(n6777) );
  XOR U6607 ( .A(n6783), .B(n6784), .Z(n6775) );
  AND U6608 ( .A(n153), .B(n6785), .Z(n6784) );
  XNOR U6609 ( .A(n6786), .B(n6787), .Z(n6781) );
  AND U6610 ( .A(n145), .B(n6788), .Z(n6787) );
  XOR U6611 ( .A(p_input[171]), .B(n6786), .Z(n6788) );
  XNOR U6612 ( .A(n6789), .B(n6790), .Z(n6786) );
  AND U6613 ( .A(n149), .B(n6785), .Z(n6790) );
  XNOR U6614 ( .A(n6789), .B(n6783), .Z(n6785) );
  XOR U6615 ( .A(n6791), .B(n6792), .Z(n6783) );
  AND U6616 ( .A(n164), .B(n6793), .Z(n6792) );
  XNOR U6617 ( .A(n6794), .B(n6795), .Z(n6789) );
  AND U6618 ( .A(n156), .B(n6796), .Z(n6795) );
  XOR U6619 ( .A(p_input[187]), .B(n6794), .Z(n6796) );
  XNOR U6620 ( .A(n6797), .B(n6798), .Z(n6794) );
  AND U6621 ( .A(n160), .B(n6793), .Z(n6798) );
  XNOR U6622 ( .A(n6797), .B(n6791), .Z(n6793) );
  XOR U6623 ( .A(n6799), .B(n6800), .Z(n6791) );
  AND U6624 ( .A(n175), .B(n6801), .Z(n6800) );
  XNOR U6625 ( .A(n6802), .B(n6803), .Z(n6797) );
  AND U6626 ( .A(n167), .B(n6804), .Z(n6803) );
  XOR U6627 ( .A(p_input[203]), .B(n6802), .Z(n6804) );
  XNOR U6628 ( .A(n6805), .B(n6806), .Z(n6802) );
  AND U6629 ( .A(n171), .B(n6801), .Z(n6806) );
  XNOR U6630 ( .A(n6805), .B(n6799), .Z(n6801) );
  XOR U6631 ( .A(n6807), .B(n6808), .Z(n6799) );
  AND U6632 ( .A(n186), .B(n6809), .Z(n6808) );
  XNOR U6633 ( .A(n6810), .B(n6811), .Z(n6805) );
  AND U6634 ( .A(n178), .B(n6812), .Z(n6811) );
  XOR U6635 ( .A(p_input[219]), .B(n6810), .Z(n6812) );
  XNOR U6636 ( .A(n6813), .B(n6814), .Z(n6810) );
  AND U6637 ( .A(n182), .B(n6809), .Z(n6814) );
  XNOR U6638 ( .A(n6813), .B(n6807), .Z(n6809) );
  XOR U6639 ( .A(n6815), .B(n6816), .Z(n6807) );
  AND U6640 ( .A(n197), .B(n6817), .Z(n6816) );
  XNOR U6641 ( .A(n6818), .B(n6819), .Z(n6813) );
  AND U6642 ( .A(n189), .B(n6820), .Z(n6819) );
  XOR U6643 ( .A(p_input[235]), .B(n6818), .Z(n6820) );
  XNOR U6644 ( .A(n6821), .B(n6822), .Z(n6818) );
  AND U6645 ( .A(n193), .B(n6817), .Z(n6822) );
  XNOR U6646 ( .A(n6821), .B(n6815), .Z(n6817) );
  XOR U6647 ( .A(n6823), .B(n6824), .Z(n6815) );
  AND U6648 ( .A(n208), .B(n6825), .Z(n6824) );
  XNOR U6649 ( .A(n6826), .B(n6827), .Z(n6821) );
  AND U6650 ( .A(n200), .B(n6828), .Z(n6827) );
  XOR U6651 ( .A(p_input[251]), .B(n6826), .Z(n6828) );
  XNOR U6652 ( .A(n6829), .B(n6830), .Z(n6826) );
  AND U6653 ( .A(n204), .B(n6825), .Z(n6830) );
  XNOR U6654 ( .A(n6829), .B(n6823), .Z(n6825) );
  XOR U6655 ( .A(n6831), .B(n6832), .Z(n6823) );
  AND U6656 ( .A(n219), .B(n6833), .Z(n6832) );
  XNOR U6657 ( .A(n6834), .B(n6835), .Z(n6829) );
  AND U6658 ( .A(n211), .B(n6836), .Z(n6835) );
  XOR U6659 ( .A(p_input[267]), .B(n6834), .Z(n6836) );
  XNOR U6660 ( .A(n6837), .B(n6838), .Z(n6834) );
  AND U6661 ( .A(n215), .B(n6833), .Z(n6838) );
  XNOR U6662 ( .A(n6837), .B(n6831), .Z(n6833) );
  XOR U6663 ( .A(n6839), .B(n6840), .Z(n6831) );
  AND U6664 ( .A(n230), .B(n6841), .Z(n6840) );
  XNOR U6665 ( .A(n6842), .B(n6843), .Z(n6837) );
  AND U6666 ( .A(n222), .B(n6844), .Z(n6843) );
  XOR U6667 ( .A(p_input[283]), .B(n6842), .Z(n6844) );
  XNOR U6668 ( .A(n6845), .B(n6846), .Z(n6842) );
  AND U6669 ( .A(n226), .B(n6841), .Z(n6846) );
  XNOR U6670 ( .A(n6845), .B(n6839), .Z(n6841) );
  XOR U6671 ( .A(n6847), .B(n6848), .Z(n6839) );
  AND U6672 ( .A(n241), .B(n6849), .Z(n6848) );
  XNOR U6673 ( .A(n6850), .B(n6851), .Z(n6845) );
  AND U6674 ( .A(n233), .B(n6852), .Z(n6851) );
  XOR U6675 ( .A(p_input[299]), .B(n6850), .Z(n6852) );
  XNOR U6676 ( .A(n6853), .B(n6854), .Z(n6850) );
  AND U6677 ( .A(n237), .B(n6849), .Z(n6854) );
  XNOR U6678 ( .A(n6853), .B(n6847), .Z(n6849) );
  XOR U6679 ( .A(n6855), .B(n6856), .Z(n6847) );
  AND U6680 ( .A(n252), .B(n6857), .Z(n6856) );
  XNOR U6681 ( .A(n6858), .B(n6859), .Z(n6853) );
  AND U6682 ( .A(n244), .B(n6860), .Z(n6859) );
  XOR U6683 ( .A(p_input[315]), .B(n6858), .Z(n6860) );
  XNOR U6684 ( .A(n6861), .B(n6862), .Z(n6858) );
  AND U6685 ( .A(n248), .B(n6857), .Z(n6862) );
  XNOR U6686 ( .A(n6861), .B(n6855), .Z(n6857) );
  XOR U6687 ( .A(n6863), .B(n6864), .Z(n6855) );
  AND U6688 ( .A(n263), .B(n6865), .Z(n6864) );
  XNOR U6689 ( .A(n6866), .B(n6867), .Z(n6861) );
  AND U6690 ( .A(n255), .B(n6868), .Z(n6867) );
  XOR U6691 ( .A(p_input[331]), .B(n6866), .Z(n6868) );
  XNOR U6692 ( .A(n6869), .B(n6870), .Z(n6866) );
  AND U6693 ( .A(n259), .B(n6865), .Z(n6870) );
  XNOR U6694 ( .A(n6869), .B(n6863), .Z(n6865) );
  XOR U6695 ( .A(n6871), .B(n6872), .Z(n6863) );
  AND U6696 ( .A(n274), .B(n6873), .Z(n6872) );
  XNOR U6697 ( .A(n6874), .B(n6875), .Z(n6869) );
  AND U6698 ( .A(n266), .B(n6876), .Z(n6875) );
  XOR U6699 ( .A(p_input[347]), .B(n6874), .Z(n6876) );
  XNOR U6700 ( .A(n6877), .B(n6878), .Z(n6874) );
  AND U6701 ( .A(n270), .B(n6873), .Z(n6878) );
  XNOR U6702 ( .A(n6877), .B(n6871), .Z(n6873) );
  XOR U6703 ( .A(n6879), .B(n6880), .Z(n6871) );
  AND U6704 ( .A(n285), .B(n6881), .Z(n6880) );
  XNOR U6705 ( .A(n6882), .B(n6883), .Z(n6877) );
  AND U6706 ( .A(n277), .B(n6884), .Z(n6883) );
  XOR U6707 ( .A(p_input[363]), .B(n6882), .Z(n6884) );
  XNOR U6708 ( .A(n6885), .B(n6886), .Z(n6882) );
  AND U6709 ( .A(n281), .B(n6881), .Z(n6886) );
  XNOR U6710 ( .A(n6885), .B(n6879), .Z(n6881) );
  XOR U6711 ( .A(n6887), .B(n6888), .Z(n6879) );
  AND U6712 ( .A(n296), .B(n6889), .Z(n6888) );
  XNOR U6713 ( .A(n6890), .B(n6891), .Z(n6885) );
  AND U6714 ( .A(n288), .B(n6892), .Z(n6891) );
  XOR U6715 ( .A(p_input[379]), .B(n6890), .Z(n6892) );
  XNOR U6716 ( .A(n6893), .B(n6894), .Z(n6890) );
  AND U6717 ( .A(n292), .B(n6889), .Z(n6894) );
  XNOR U6718 ( .A(n6893), .B(n6887), .Z(n6889) );
  XOR U6719 ( .A(n6895), .B(n6896), .Z(n6887) );
  AND U6720 ( .A(n307), .B(n6897), .Z(n6896) );
  XNOR U6721 ( .A(n6898), .B(n6899), .Z(n6893) );
  AND U6722 ( .A(n299), .B(n6900), .Z(n6899) );
  XOR U6723 ( .A(p_input[395]), .B(n6898), .Z(n6900) );
  XNOR U6724 ( .A(n6901), .B(n6902), .Z(n6898) );
  AND U6725 ( .A(n303), .B(n6897), .Z(n6902) );
  XNOR U6726 ( .A(n6901), .B(n6895), .Z(n6897) );
  XOR U6727 ( .A(n6903), .B(n6904), .Z(n6895) );
  AND U6728 ( .A(n318), .B(n6905), .Z(n6904) );
  XNOR U6729 ( .A(n6906), .B(n6907), .Z(n6901) );
  AND U6730 ( .A(n310), .B(n6908), .Z(n6907) );
  XOR U6731 ( .A(p_input[411]), .B(n6906), .Z(n6908) );
  XNOR U6732 ( .A(n6909), .B(n6910), .Z(n6906) );
  AND U6733 ( .A(n314), .B(n6905), .Z(n6910) );
  XNOR U6734 ( .A(n6909), .B(n6903), .Z(n6905) );
  XOR U6735 ( .A(n6911), .B(n6912), .Z(n6903) );
  AND U6736 ( .A(n329), .B(n6913), .Z(n6912) );
  XNOR U6737 ( .A(n6914), .B(n6915), .Z(n6909) );
  AND U6738 ( .A(n321), .B(n6916), .Z(n6915) );
  XOR U6739 ( .A(p_input[427]), .B(n6914), .Z(n6916) );
  XNOR U6740 ( .A(n6917), .B(n6918), .Z(n6914) );
  AND U6741 ( .A(n325), .B(n6913), .Z(n6918) );
  XNOR U6742 ( .A(n6917), .B(n6911), .Z(n6913) );
  XOR U6743 ( .A(n6919), .B(n6920), .Z(n6911) );
  AND U6744 ( .A(n340), .B(n6921), .Z(n6920) );
  XNOR U6745 ( .A(n6922), .B(n6923), .Z(n6917) );
  AND U6746 ( .A(n332), .B(n6924), .Z(n6923) );
  XOR U6747 ( .A(p_input[443]), .B(n6922), .Z(n6924) );
  XNOR U6748 ( .A(n6925), .B(n6926), .Z(n6922) );
  AND U6749 ( .A(n336), .B(n6921), .Z(n6926) );
  XNOR U6750 ( .A(n6925), .B(n6919), .Z(n6921) );
  XOR U6751 ( .A(n6927), .B(n6928), .Z(n6919) );
  AND U6752 ( .A(n351), .B(n6929), .Z(n6928) );
  XNOR U6753 ( .A(n6930), .B(n6931), .Z(n6925) );
  AND U6754 ( .A(n343), .B(n6932), .Z(n6931) );
  XOR U6755 ( .A(p_input[459]), .B(n6930), .Z(n6932) );
  XNOR U6756 ( .A(n6933), .B(n6934), .Z(n6930) );
  AND U6757 ( .A(n347), .B(n6929), .Z(n6934) );
  XNOR U6758 ( .A(n6933), .B(n6927), .Z(n6929) );
  XOR U6759 ( .A(n6935), .B(n6936), .Z(n6927) );
  AND U6760 ( .A(n362), .B(n6937), .Z(n6936) );
  XNOR U6761 ( .A(n6938), .B(n6939), .Z(n6933) );
  AND U6762 ( .A(n354), .B(n6940), .Z(n6939) );
  XOR U6763 ( .A(p_input[475]), .B(n6938), .Z(n6940) );
  XNOR U6764 ( .A(n6941), .B(n6942), .Z(n6938) );
  AND U6765 ( .A(n358), .B(n6937), .Z(n6942) );
  XNOR U6766 ( .A(n6941), .B(n6935), .Z(n6937) );
  XOR U6767 ( .A(n6943), .B(n6944), .Z(n6935) );
  AND U6768 ( .A(n373), .B(n6945), .Z(n6944) );
  XNOR U6769 ( .A(n6946), .B(n6947), .Z(n6941) );
  AND U6770 ( .A(n365), .B(n6948), .Z(n6947) );
  XOR U6771 ( .A(p_input[491]), .B(n6946), .Z(n6948) );
  XNOR U6772 ( .A(n6949), .B(n6950), .Z(n6946) );
  AND U6773 ( .A(n369), .B(n6945), .Z(n6950) );
  XNOR U6774 ( .A(n6949), .B(n6943), .Z(n6945) );
  XOR U6775 ( .A(n6951), .B(n6952), .Z(n6943) );
  AND U6776 ( .A(n384), .B(n6953), .Z(n6952) );
  XNOR U6777 ( .A(n6954), .B(n6955), .Z(n6949) );
  AND U6778 ( .A(n376), .B(n6956), .Z(n6955) );
  XOR U6779 ( .A(p_input[507]), .B(n6954), .Z(n6956) );
  XNOR U6780 ( .A(n6957), .B(n6958), .Z(n6954) );
  AND U6781 ( .A(n380), .B(n6953), .Z(n6958) );
  XNOR U6782 ( .A(n6957), .B(n6951), .Z(n6953) );
  XOR U6783 ( .A(n6959), .B(n6960), .Z(n6951) );
  AND U6784 ( .A(n395), .B(n6961), .Z(n6960) );
  XNOR U6785 ( .A(n6962), .B(n6963), .Z(n6957) );
  AND U6786 ( .A(n387), .B(n6964), .Z(n6963) );
  XOR U6787 ( .A(p_input[523]), .B(n6962), .Z(n6964) );
  XNOR U6788 ( .A(n6965), .B(n6966), .Z(n6962) );
  AND U6789 ( .A(n391), .B(n6961), .Z(n6966) );
  XNOR U6790 ( .A(n6965), .B(n6959), .Z(n6961) );
  XOR U6791 ( .A(n6967), .B(n6968), .Z(n6959) );
  AND U6792 ( .A(n406), .B(n6969), .Z(n6968) );
  XNOR U6793 ( .A(n6970), .B(n6971), .Z(n6965) );
  AND U6794 ( .A(n398), .B(n6972), .Z(n6971) );
  XOR U6795 ( .A(p_input[539]), .B(n6970), .Z(n6972) );
  XNOR U6796 ( .A(n6973), .B(n6974), .Z(n6970) );
  AND U6797 ( .A(n402), .B(n6969), .Z(n6974) );
  XNOR U6798 ( .A(n6973), .B(n6967), .Z(n6969) );
  XOR U6799 ( .A(n6975), .B(n6976), .Z(n6967) );
  AND U6800 ( .A(n417), .B(n6977), .Z(n6976) );
  XNOR U6801 ( .A(n6978), .B(n6979), .Z(n6973) );
  AND U6802 ( .A(n409), .B(n6980), .Z(n6979) );
  XOR U6803 ( .A(p_input[555]), .B(n6978), .Z(n6980) );
  XNOR U6804 ( .A(n6981), .B(n6982), .Z(n6978) );
  AND U6805 ( .A(n413), .B(n6977), .Z(n6982) );
  XNOR U6806 ( .A(n6981), .B(n6975), .Z(n6977) );
  XOR U6807 ( .A(n6983), .B(n6984), .Z(n6975) );
  AND U6808 ( .A(n428), .B(n6985), .Z(n6984) );
  XNOR U6809 ( .A(n6986), .B(n6987), .Z(n6981) );
  AND U6810 ( .A(n420), .B(n6988), .Z(n6987) );
  XOR U6811 ( .A(p_input[571]), .B(n6986), .Z(n6988) );
  XNOR U6812 ( .A(n6989), .B(n6990), .Z(n6986) );
  AND U6813 ( .A(n424), .B(n6985), .Z(n6990) );
  XNOR U6814 ( .A(n6989), .B(n6983), .Z(n6985) );
  XOR U6815 ( .A(n6991), .B(n6992), .Z(n6983) );
  AND U6816 ( .A(n439), .B(n6993), .Z(n6992) );
  XNOR U6817 ( .A(n6994), .B(n6995), .Z(n6989) );
  AND U6818 ( .A(n431), .B(n6996), .Z(n6995) );
  XOR U6819 ( .A(p_input[587]), .B(n6994), .Z(n6996) );
  XNOR U6820 ( .A(n6997), .B(n6998), .Z(n6994) );
  AND U6821 ( .A(n435), .B(n6993), .Z(n6998) );
  XNOR U6822 ( .A(n6997), .B(n6991), .Z(n6993) );
  XOR U6823 ( .A(n6999), .B(n7000), .Z(n6991) );
  AND U6824 ( .A(n450), .B(n7001), .Z(n7000) );
  XNOR U6825 ( .A(n7002), .B(n7003), .Z(n6997) );
  AND U6826 ( .A(n442), .B(n7004), .Z(n7003) );
  XOR U6827 ( .A(p_input[603]), .B(n7002), .Z(n7004) );
  XNOR U6828 ( .A(n7005), .B(n7006), .Z(n7002) );
  AND U6829 ( .A(n446), .B(n7001), .Z(n7006) );
  XNOR U6830 ( .A(n7005), .B(n6999), .Z(n7001) );
  XOR U6831 ( .A(n7007), .B(n7008), .Z(n6999) );
  AND U6832 ( .A(n461), .B(n7009), .Z(n7008) );
  XNOR U6833 ( .A(n7010), .B(n7011), .Z(n7005) );
  AND U6834 ( .A(n453), .B(n7012), .Z(n7011) );
  XOR U6835 ( .A(p_input[619]), .B(n7010), .Z(n7012) );
  XNOR U6836 ( .A(n7013), .B(n7014), .Z(n7010) );
  AND U6837 ( .A(n457), .B(n7009), .Z(n7014) );
  XNOR U6838 ( .A(n7013), .B(n7007), .Z(n7009) );
  XOR U6839 ( .A(n7015), .B(n7016), .Z(n7007) );
  AND U6840 ( .A(n472), .B(n7017), .Z(n7016) );
  XNOR U6841 ( .A(n7018), .B(n7019), .Z(n7013) );
  AND U6842 ( .A(n464), .B(n7020), .Z(n7019) );
  XOR U6843 ( .A(p_input[635]), .B(n7018), .Z(n7020) );
  XNOR U6844 ( .A(n7021), .B(n7022), .Z(n7018) );
  AND U6845 ( .A(n468), .B(n7017), .Z(n7022) );
  XNOR U6846 ( .A(n7021), .B(n7015), .Z(n7017) );
  XOR U6847 ( .A(n7023), .B(n7024), .Z(n7015) );
  AND U6848 ( .A(n483), .B(n7025), .Z(n7024) );
  XNOR U6849 ( .A(n7026), .B(n7027), .Z(n7021) );
  AND U6850 ( .A(n475), .B(n7028), .Z(n7027) );
  XOR U6851 ( .A(p_input[651]), .B(n7026), .Z(n7028) );
  XNOR U6852 ( .A(n7029), .B(n7030), .Z(n7026) );
  AND U6853 ( .A(n479), .B(n7025), .Z(n7030) );
  XNOR U6854 ( .A(n7029), .B(n7023), .Z(n7025) );
  XOR U6855 ( .A(n7031), .B(n7032), .Z(n7023) );
  AND U6856 ( .A(n494), .B(n7033), .Z(n7032) );
  XNOR U6857 ( .A(n7034), .B(n7035), .Z(n7029) );
  AND U6858 ( .A(n486), .B(n7036), .Z(n7035) );
  XOR U6859 ( .A(p_input[667]), .B(n7034), .Z(n7036) );
  XNOR U6860 ( .A(n7037), .B(n7038), .Z(n7034) );
  AND U6861 ( .A(n490), .B(n7033), .Z(n7038) );
  XNOR U6862 ( .A(n7037), .B(n7031), .Z(n7033) );
  XOR U6863 ( .A(n7039), .B(n7040), .Z(n7031) );
  AND U6864 ( .A(n505), .B(n7041), .Z(n7040) );
  XNOR U6865 ( .A(n7042), .B(n7043), .Z(n7037) );
  AND U6866 ( .A(n497), .B(n7044), .Z(n7043) );
  XOR U6867 ( .A(p_input[683]), .B(n7042), .Z(n7044) );
  XNOR U6868 ( .A(n7045), .B(n7046), .Z(n7042) );
  AND U6869 ( .A(n501), .B(n7041), .Z(n7046) );
  XNOR U6870 ( .A(n7045), .B(n7039), .Z(n7041) );
  XOR U6871 ( .A(n7047), .B(n7048), .Z(n7039) );
  AND U6872 ( .A(n516), .B(n7049), .Z(n7048) );
  XNOR U6873 ( .A(n7050), .B(n7051), .Z(n7045) );
  AND U6874 ( .A(n508), .B(n7052), .Z(n7051) );
  XOR U6875 ( .A(p_input[699]), .B(n7050), .Z(n7052) );
  XNOR U6876 ( .A(n7053), .B(n7054), .Z(n7050) );
  AND U6877 ( .A(n512), .B(n7049), .Z(n7054) );
  XNOR U6878 ( .A(n7053), .B(n7047), .Z(n7049) );
  XOR U6879 ( .A(n7055), .B(n7056), .Z(n7047) );
  AND U6880 ( .A(n527), .B(n7057), .Z(n7056) );
  XNOR U6881 ( .A(n7058), .B(n7059), .Z(n7053) );
  AND U6882 ( .A(n519), .B(n7060), .Z(n7059) );
  XOR U6883 ( .A(p_input[715]), .B(n7058), .Z(n7060) );
  XNOR U6884 ( .A(n7061), .B(n7062), .Z(n7058) );
  AND U6885 ( .A(n523), .B(n7057), .Z(n7062) );
  XNOR U6886 ( .A(n7061), .B(n7055), .Z(n7057) );
  XOR U6887 ( .A(n7063), .B(n7064), .Z(n7055) );
  AND U6888 ( .A(n538), .B(n7065), .Z(n7064) );
  XNOR U6889 ( .A(n7066), .B(n7067), .Z(n7061) );
  AND U6890 ( .A(n530), .B(n7068), .Z(n7067) );
  XOR U6891 ( .A(p_input[731]), .B(n7066), .Z(n7068) );
  XNOR U6892 ( .A(n7069), .B(n7070), .Z(n7066) );
  AND U6893 ( .A(n534), .B(n7065), .Z(n7070) );
  XNOR U6894 ( .A(n7069), .B(n7063), .Z(n7065) );
  XOR U6895 ( .A(n7071), .B(n7072), .Z(n7063) );
  AND U6896 ( .A(n549), .B(n7073), .Z(n7072) );
  XNOR U6897 ( .A(n7074), .B(n7075), .Z(n7069) );
  AND U6898 ( .A(n541), .B(n7076), .Z(n7075) );
  XOR U6899 ( .A(p_input[747]), .B(n7074), .Z(n7076) );
  XNOR U6900 ( .A(n7077), .B(n7078), .Z(n7074) );
  AND U6901 ( .A(n545), .B(n7073), .Z(n7078) );
  XNOR U6902 ( .A(n7077), .B(n7071), .Z(n7073) );
  XOR U6903 ( .A(n7079), .B(n7080), .Z(n7071) );
  AND U6904 ( .A(n560), .B(n7081), .Z(n7080) );
  XNOR U6905 ( .A(n7082), .B(n7083), .Z(n7077) );
  AND U6906 ( .A(n552), .B(n7084), .Z(n7083) );
  XOR U6907 ( .A(p_input[763]), .B(n7082), .Z(n7084) );
  XNOR U6908 ( .A(n7085), .B(n7086), .Z(n7082) );
  AND U6909 ( .A(n556), .B(n7081), .Z(n7086) );
  XNOR U6910 ( .A(n7085), .B(n7079), .Z(n7081) );
  XOR U6911 ( .A(n7087), .B(n7088), .Z(n7079) );
  AND U6912 ( .A(n571), .B(n7089), .Z(n7088) );
  XNOR U6913 ( .A(n7090), .B(n7091), .Z(n7085) );
  AND U6914 ( .A(n563), .B(n7092), .Z(n7091) );
  XOR U6915 ( .A(p_input[779]), .B(n7090), .Z(n7092) );
  XNOR U6916 ( .A(n7093), .B(n7094), .Z(n7090) );
  AND U6917 ( .A(n567), .B(n7089), .Z(n7094) );
  XNOR U6918 ( .A(n7093), .B(n7087), .Z(n7089) );
  XOR U6919 ( .A(n7095), .B(n7096), .Z(n7087) );
  AND U6920 ( .A(n582), .B(n7097), .Z(n7096) );
  XNOR U6921 ( .A(n7098), .B(n7099), .Z(n7093) );
  AND U6922 ( .A(n574), .B(n7100), .Z(n7099) );
  XOR U6923 ( .A(p_input[795]), .B(n7098), .Z(n7100) );
  XNOR U6924 ( .A(n7101), .B(n7102), .Z(n7098) );
  AND U6925 ( .A(n578), .B(n7097), .Z(n7102) );
  XNOR U6926 ( .A(n7101), .B(n7095), .Z(n7097) );
  XOR U6927 ( .A(n7103), .B(n7104), .Z(n7095) );
  AND U6928 ( .A(n593), .B(n7105), .Z(n7104) );
  XNOR U6929 ( .A(n7106), .B(n7107), .Z(n7101) );
  AND U6930 ( .A(n585), .B(n7108), .Z(n7107) );
  XOR U6931 ( .A(p_input[811]), .B(n7106), .Z(n7108) );
  XNOR U6932 ( .A(n7109), .B(n7110), .Z(n7106) );
  AND U6933 ( .A(n589), .B(n7105), .Z(n7110) );
  XNOR U6934 ( .A(n7109), .B(n7103), .Z(n7105) );
  XOR U6935 ( .A(n7111), .B(n7112), .Z(n7103) );
  AND U6936 ( .A(n604), .B(n7113), .Z(n7112) );
  XNOR U6937 ( .A(n7114), .B(n7115), .Z(n7109) );
  AND U6938 ( .A(n596), .B(n7116), .Z(n7115) );
  XOR U6939 ( .A(p_input[827]), .B(n7114), .Z(n7116) );
  XNOR U6940 ( .A(n7117), .B(n7118), .Z(n7114) );
  AND U6941 ( .A(n600), .B(n7113), .Z(n7118) );
  XNOR U6942 ( .A(n7117), .B(n7111), .Z(n7113) );
  XOR U6943 ( .A(n7119), .B(n7120), .Z(n7111) );
  AND U6944 ( .A(n615), .B(n7121), .Z(n7120) );
  XNOR U6945 ( .A(n7122), .B(n7123), .Z(n7117) );
  AND U6946 ( .A(n607), .B(n7124), .Z(n7123) );
  XOR U6947 ( .A(p_input[843]), .B(n7122), .Z(n7124) );
  XNOR U6948 ( .A(n7125), .B(n7126), .Z(n7122) );
  AND U6949 ( .A(n611), .B(n7121), .Z(n7126) );
  XNOR U6950 ( .A(n7125), .B(n7119), .Z(n7121) );
  XOR U6951 ( .A(n7127), .B(n7128), .Z(n7119) );
  AND U6952 ( .A(n626), .B(n7129), .Z(n7128) );
  XNOR U6953 ( .A(n7130), .B(n7131), .Z(n7125) );
  AND U6954 ( .A(n618), .B(n7132), .Z(n7131) );
  XOR U6955 ( .A(p_input[859]), .B(n7130), .Z(n7132) );
  XNOR U6956 ( .A(n7133), .B(n7134), .Z(n7130) );
  AND U6957 ( .A(n622), .B(n7129), .Z(n7134) );
  XNOR U6958 ( .A(n7133), .B(n7127), .Z(n7129) );
  XOR U6959 ( .A(n7135), .B(n7136), .Z(n7127) );
  AND U6960 ( .A(n637), .B(n7137), .Z(n7136) );
  XNOR U6961 ( .A(n7138), .B(n7139), .Z(n7133) );
  AND U6962 ( .A(n629), .B(n7140), .Z(n7139) );
  XOR U6963 ( .A(p_input[875]), .B(n7138), .Z(n7140) );
  XNOR U6964 ( .A(n7141), .B(n7142), .Z(n7138) );
  AND U6965 ( .A(n633), .B(n7137), .Z(n7142) );
  XNOR U6966 ( .A(n7141), .B(n7135), .Z(n7137) );
  XOR U6967 ( .A(n7143), .B(n7144), .Z(n7135) );
  AND U6968 ( .A(n648), .B(n7145), .Z(n7144) );
  XNOR U6969 ( .A(n7146), .B(n7147), .Z(n7141) );
  AND U6970 ( .A(n640), .B(n7148), .Z(n7147) );
  XOR U6971 ( .A(p_input[891]), .B(n7146), .Z(n7148) );
  XNOR U6972 ( .A(n7149), .B(n7150), .Z(n7146) );
  AND U6973 ( .A(n644), .B(n7145), .Z(n7150) );
  XNOR U6974 ( .A(n7149), .B(n7143), .Z(n7145) );
  XOR U6975 ( .A(n7151), .B(n7152), .Z(n7143) );
  AND U6976 ( .A(n659), .B(n7153), .Z(n7152) );
  XNOR U6977 ( .A(n7154), .B(n7155), .Z(n7149) );
  AND U6978 ( .A(n651), .B(n7156), .Z(n7155) );
  XOR U6979 ( .A(p_input[907]), .B(n7154), .Z(n7156) );
  XNOR U6980 ( .A(n7157), .B(n7158), .Z(n7154) );
  AND U6981 ( .A(n655), .B(n7153), .Z(n7158) );
  XNOR U6982 ( .A(n7157), .B(n7151), .Z(n7153) );
  XOR U6983 ( .A(n7159), .B(n7160), .Z(n7151) );
  AND U6984 ( .A(n670), .B(n7161), .Z(n7160) );
  XNOR U6985 ( .A(n7162), .B(n7163), .Z(n7157) );
  AND U6986 ( .A(n662), .B(n7164), .Z(n7163) );
  XOR U6987 ( .A(p_input[923]), .B(n7162), .Z(n7164) );
  XNOR U6988 ( .A(n7165), .B(n7166), .Z(n7162) );
  AND U6989 ( .A(n666), .B(n7161), .Z(n7166) );
  XNOR U6990 ( .A(n7165), .B(n7159), .Z(n7161) );
  XOR U6991 ( .A(n7167), .B(n7168), .Z(n7159) );
  AND U6992 ( .A(n681), .B(n7169), .Z(n7168) );
  XNOR U6993 ( .A(n7170), .B(n7171), .Z(n7165) );
  AND U6994 ( .A(n673), .B(n7172), .Z(n7171) );
  XOR U6995 ( .A(p_input[939]), .B(n7170), .Z(n7172) );
  XNOR U6996 ( .A(n7173), .B(n7174), .Z(n7170) );
  AND U6997 ( .A(n677), .B(n7169), .Z(n7174) );
  XNOR U6998 ( .A(n7173), .B(n7167), .Z(n7169) );
  XOR U6999 ( .A(n7175), .B(n7176), .Z(n7167) );
  AND U7000 ( .A(n692), .B(n7177), .Z(n7176) );
  XNOR U7001 ( .A(n7178), .B(n7179), .Z(n7173) );
  AND U7002 ( .A(n684), .B(n7180), .Z(n7179) );
  XOR U7003 ( .A(p_input[955]), .B(n7178), .Z(n7180) );
  XNOR U7004 ( .A(n7181), .B(n7182), .Z(n7178) );
  AND U7005 ( .A(n688), .B(n7177), .Z(n7182) );
  XNOR U7006 ( .A(n7181), .B(n7175), .Z(n7177) );
  XOR U7007 ( .A(n7183), .B(n7184), .Z(n7175) );
  AND U7008 ( .A(n703), .B(n7185), .Z(n7184) );
  XNOR U7009 ( .A(n7186), .B(n7187), .Z(n7181) );
  AND U7010 ( .A(n695), .B(n7188), .Z(n7187) );
  XOR U7011 ( .A(p_input[971]), .B(n7186), .Z(n7188) );
  XNOR U7012 ( .A(n7189), .B(n7190), .Z(n7186) );
  AND U7013 ( .A(n699), .B(n7185), .Z(n7190) );
  XNOR U7014 ( .A(n7189), .B(n7183), .Z(n7185) );
  XOR U7015 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n7191), .Z(n7183) );
  AND U7016 ( .A(n713), .B(n7192), .Z(n7191) );
  XNOR U7017 ( .A(n7193), .B(n7194), .Z(n7189) );
  AND U7018 ( .A(n706), .B(n7195), .Z(n7194) );
  XOR U7019 ( .A(p_input[987]), .B(n7193), .Z(n7195) );
  XNOR U7020 ( .A(n7196), .B(n7197), .Z(n7193) );
  AND U7021 ( .A(n710), .B(n7192), .Z(n7197) );
  XOR U7022 ( .A(n7198), .B(n7196), .Z(n7192) );
  IV U7023 ( .A(\knn_comb_/min_val_out[0][11] ), .Z(n7198) );
  IV U7024 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n7196) );
  XOR U7025 ( .A(n27), .B(n7199), .Z(o[10]) );
  AND U7026 ( .A(n30), .B(n7200), .Z(n27) );
  XOR U7027 ( .A(n28), .B(n7199), .Z(n7200) );
  XOR U7028 ( .A(n7201), .B(n7202), .Z(n7199) );
  AND U7029 ( .A(n42), .B(n7203), .Z(n7202) );
  XOR U7030 ( .A(n7204), .B(n7205), .Z(n28) );
  AND U7031 ( .A(n34), .B(n7206), .Z(n7205) );
  XOR U7032 ( .A(p_input[10]), .B(n7204), .Z(n7206) );
  XNOR U7033 ( .A(n7207), .B(n7208), .Z(n7204) );
  AND U7034 ( .A(n38), .B(n7203), .Z(n7208) );
  XNOR U7035 ( .A(n7207), .B(n7201), .Z(n7203) );
  XOR U7036 ( .A(n7209), .B(n7210), .Z(n7201) );
  AND U7037 ( .A(n54), .B(n7211), .Z(n7210) );
  XNOR U7038 ( .A(n7212), .B(n7213), .Z(n7207) );
  AND U7039 ( .A(n46), .B(n7214), .Z(n7213) );
  XOR U7040 ( .A(p_input[26]), .B(n7212), .Z(n7214) );
  XNOR U7041 ( .A(n7215), .B(n7216), .Z(n7212) );
  AND U7042 ( .A(n50), .B(n7211), .Z(n7216) );
  XNOR U7043 ( .A(n7215), .B(n7209), .Z(n7211) );
  XOR U7044 ( .A(n7217), .B(n7218), .Z(n7209) );
  AND U7045 ( .A(n65), .B(n7219), .Z(n7218) );
  XNOR U7046 ( .A(n7220), .B(n7221), .Z(n7215) );
  AND U7047 ( .A(n57), .B(n7222), .Z(n7221) );
  XOR U7048 ( .A(p_input[42]), .B(n7220), .Z(n7222) );
  XNOR U7049 ( .A(n7223), .B(n7224), .Z(n7220) );
  AND U7050 ( .A(n61), .B(n7219), .Z(n7224) );
  XNOR U7051 ( .A(n7223), .B(n7217), .Z(n7219) );
  XOR U7052 ( .A(n7225), .B(n7226), .Z(n7217) );
  AND U7053 ( .A(n76), .B(n7227), .Z(n7226) );
  XNOR U7054 ( .A(n7228), .B(n7229), .Z(n7223) );
  AND U7055 ( .A(n68), .B(n7230), .Z(n7229) );
  XOR U7056 ( .A(p_input[58]), .B(n7228), .Z(n7230) );
  XNOR U7057 ( .A(n7231), .B(n7232), .Z(n7228) );
  AND U7058 ( .A(n72), .B(n7227), .Z(n7232) );
  XNOR U7059 ( .A(n7231), .B(n7225), .Z(n7227) );
  XOR U7060 ( .A(n7233), .B(n7234), .Z(n7225) );
  AND U7061 ( .A(n87), .B(n7235), .Z(n7234) );
  XNOR U7062 ( .A(n7236), .B(n7237), .Z(n7231) );
  AND U7063 ( .A(n79), .B(n7238), .Z(n7237) );
  XOR U7064 ( .A(p_input[74]), .B(n7236), .Z(n7238) );
  XNOR U7065 ( .A(n7239), .B(n7240), .Z(n7236) );
  AND U7066 ( .A(n83), .B(n7235), .Z(n7240) );
  XNOR U7067 ( .A(n7239), .B(n7233), .Z(n7235) );
  XOR U7068 ( .A(n7241), .B(n7242), .Z(n7233) );
  AND U7069 ( .A(n98), .B(n7243), .Z(n7242) );
  XNOR U7070 ( .A(n7244), .B(n7245), .Z(n7239) );
  AND U7071 ( .A(n90), .B(n7246), .Z(n7245) );
  XOR U7072 ( .A(p_input[90]), .B(n7244), .Z(n7246) );
  XNOR U7073 ( .A(n7247), .B(n7248), .Z(n7244) );
  AND U7074 ( .A(n94), .B(n7243), .Z(n7248) );
  XNOR U7075 ( .A(n7247), .B(n7241), .Z(n7243) );
  XOR U7076 ( .A(n7249), .B(n7250), .Z(n7241) );
  AND U7077 ( .A(n109), .B(n7251), .Z(n7250) );
  XNOR U7078 ( .A(n7252), .B(n7253), .Z(n7247) );
  AND U7079 ( .A(n101), .B(n7254), .Z(n7253) );
  XOR U7080 ( .A(p_input[106]), .B(n7252), .Z(n7254) );
  XNOR U7081 ( .A(n7255), .B(n7256), .Z(n7252) );
  AND U7082 ( .A(n105), .B(n7251), .Z(n7256) );
  XNOR U7083 ( .A(n7255), .B(n7249), .Z(n7251) );
  XOR U7084 ( .A(n7257), .B(n7258), .Z(n7249) );
  AND U7085 ( .A(n120), .B(n7259), .Z(n7258) );
  XNOR U7086 ( .A(n7260), .B(n7261), .Z(n7255) );
  AND U7087 ( .A(n112), .B(n7262), .Z(n7261) );
  XOR U7088 ( .A(p_input[122]), .B(n7260), .Z(n7262) );
  XNOR U7089 ( .A(n7263), .B(n7264), .Z(n7260) );
  AND U7090 ( .A(n116), .B(n7259), .Z(n7264) );
  XNOR U7091 ( .A(n7263), .B(n7257), .Z(n7259) );
  XOR U7092 ( .A(n7265), .B(n7266), .Z(n7257) );
  AND U7093 ( .A(n131), .B(n7267), .Z(n7266) );
  XNOR U7094 ( .A(n7268), .B(n7269), .Z(n7263) );
  AND U7095 ( .A(n123), .B(n7270), .Z(n7269) );
  XOR U7096 ( .A(p_input[138]), .B(n7268), .Z(n7270) );
  XNOR U7097 ( .A(n7271), .B(n7272), .Z(n7268) );
  AND U7098 ( .A(n127), .B(n7267), .Z(n7272) );
  XNOR U7099 ( .A(n7271), .B(n7265), .Z(n7267) );
  XOR U7100 ( .A(n7273), .B(n7274), .Z(n7265) );
  AND U7101 ( .A(n142), .B(n7275), .Z(n7274) );
  XNOR U7102 ( .A(n7276), .B(n7277), .Z(n7271) );
  AND U7103 ( .A(n134), .B(n7278), .Z(n7277) );
  XOR U7104 ( .A(p_input[154]), .B(n7276), .Z(n7278) );
  XNOR U7105 ( .A(n7279), .B(n7280), .Z(n7276) );
  AND U7106 ( .A(n138), .B(n7275), .Z(n7280) );
  XNOR U7107 ( .A(n7279), .B(n7273), .Z(n7275) );
  XOR U7108 ( .A(n7281), .B(n7282), .Z(n7273) );
  AND U7109 ( .A(n153), .B(n7283), .Z(n7282) );
  XNOR U7110 ( .A(n7284), .B(n7285), .Z(n7279) );
  AND U7111 ( .A(n145), .B(n7286), .Z(n7285) );
  XOR U7112 ( .A(p_input[170]), .B(n7284), .Z(n7286) );
  XNOR U7113 ( .A(n7287), .B(n7288), .Z(n7284) );
  AND U7114 ( .A(n149), .B(n7283), .Z(n7288) );
  XNOR U7115 ( .A(n7287), .B(n7281), .Z(n7283) );
  XOR U7116 ( .A(n7289), .B(n7290), .Z(n7281) );
  AND U7117 ( .A(n164), .B(n7291), .Z(n7290) );
  XNOR U7118 ( .A(n7292), .B(n7293), .Z(n7287) );
  AND U7119 ( .A(n156), .B(n7294), .Z(n7293) );
  XOR U7120 ( .A(p_input[186]), .B(n7292), .Z(n7294) );
  XNOR U7121 ( .A(n7295), .B(n7296), .Z(n7292) );
  AND U7122 ( .A(n160), .B(n7291), .Z(n7296) );
  XNOR U7123 ( .A(n7295), .B(n7289), .Z(n7291) );
  XOR U7124 ( .A(n7297), .B(n7298), .Z(n7289) );
  AND U7125 ( .A(n175), .B(n7299), .Z(n7298) );
  XNOR U7126 ( .A(n7300), .B(n7301), .Z(n7295) );
  AND U7127 ( .A(n167), .B(n7302), .Z(n7301) );
  XOR U7128 ( .A(p_input[202]), .B(n7300), .Z(n7302) );
  XNOR U7129 ( .A(n7303), .B(n7304), .Z(n7300) );
  AND U7130 ( .A(n171), .B(n7299), .Z(n7304) );
  XNOR U7131 ( .A(n7303), .B(n7297), .Z(n7299) );
  XOR U7132 ( .A(n7305), .B(n7306), .Z(n7297) );
  AND U7133 ( .A(n186), .B(n7307), .Z(n7306) );
  XNOR U7134 ( .A(n7308), .B(n7309), .Z(n7303) );
  AND U7135 ( .A(n178), .B(n7310), .Z(n7309) );
  XOR U7136 ( .A(p_input[218]), .B(n7308), .Z(n7310) );
  XNOR U7137 ( .A(n7311), .B(n7312), .Z(n7308) );
  AND U7138 ( .A(n182), .B(n7307), .Z(n7312) );
  XNOR U7139 ( .A(n7311), .B(n7305), .Z(n7307) );
  XOR U7140 ( .A(n7313), .B(n7314), .Z(n7305) );
  AND U7141 ( .A(n197), .B(n7315), .Z(n7314) );
  XNOR U7142 ( .A(n7316), .B(n7317), .Z(n7311) );
  AND U7143 ( .A(n189), .B(n7318), .Z(n7317) );
  XOR U7144 ( .A(p_input[234]), .B(n7316), .Z(n7318) );
  XNOR U7145 ( .A(n7319), .B(n7320), .Z(n7316) );
  AND U7146 ( .A(n193), .B(n7315), .Z(n7320) );
  XNOR U7147 ( .A(n7319), .B(n7313), .Z(n7315) );
  XOR U7148 ( .A(n7321), .B(n7322), .Z(n7313) );
  AND U7149 ( .A(n208), .B(n7323), .Z(n7322) );
  XNOR U7150 ( .A(n7324), .B(n7325), .Z(n7319) );
  AND U7151 ( .A(n200), .B(n7326), .Z(n7325) );
  XOR U7152 ( .A(p_input[250]), .B(n7324), .Z(n7326) );
  XNOR U7153 ( .A(n7327), .B(n7328), .Z(n7324) );
  AND U7154 ( .A(n204), .B(n7323), .Z(n7328) );
  XNOR U7155 ( .A(n7327), .B(n7321), .Z(n7323) );
  XOR U7156 ( .A(n7329), .B(n7330), .Z(n7321) );
  AND U7157 ( .A(n219), .B(n7331), .Z(n7330) );
  XNOR U7158 ( .A(n7332), .B(n7333), .Z(n7327) );
  AND U7159 ( .A(n211), .B(n7334), .Z(n7333) );
  XOR U7160 ( .A(p_input[266]), .B(n7332), .Z(n7334) );
  XNOR U7161 ( .A(n7335), .B(n7336), .Z(n7332) );
  AND U7162 ( .A(n215), .B(n7331), .Z(n7336) );
  XNOR U7163 ( .A(n7335), .B(n7329), .Z(n7331) );
  XOR U7164 ( .A(n7337), .B(n7338), .Z(n7329) );
  AND U7165 ( .A(n230), .B(n7339), .Z(n7338) );
  XNOR U7166 ( .A(n7340), .B(n7341), .Z(n7335) );
  AND U7167 ( .A(n222), .B(n7342), .Z(n7341) );
  XOR U7168 ( .A(p_input[282]), .B(n7340), .Z(n7342) );
  XNOR U7169 ( .A(n7343), .B(n7344), .Z(n7340) );
  AND U7170 ( .A(n226), .B(n7339), .Z(n7344) );
  XNOR U7171 ( .A(n7343), .B(n7337), .Z(n7339) );
  XOR U7172 ( .A(n7345), .B(n7346), .Z(n7337) );
  AND U7173 ( .A(n241), .B(n7347), .Z(n7346) );
  XNOR U7174 ( .A(n7348), .B(n7349), .Z(n7343) );
  AND U7175 ( .A(n233), .B(n7350), .Z(n7349) );
  XOR U7176 ( .A(p_input[298]), .B(n7348), .Z(n7350) );
  XNOR U7177 ( .A(n7351), .B(n7352), .Z(n7348) );
  AND U7178 ( .A(n237), .B(n7347), .Z(n7352) );
  XNOR U7179 ( .A(n7351), .B(n7345), .Z(n7347) );
  XOR U7180 ( .A(n7353), .B(n7354), .Z(n7345) );
  AND U7181 ( .A(n252), .B(n7355), .Z(n7354) );
  XNOR U7182 ( .A(n7356), .B(n7357), .Z(n7351) );
  AND U7183 ( .A(n244), .B(n7358), .Z(n7357) );
  XOR U7184 ( .A(p_input[314]), .B(n7356), .Z(n7358) );
  XNOR U7185 ( .A(n7359), .B(n7360), .Z(n7356) );
  AND U7186 ( .A(n248), .B(n7355), .Z(n7360) );
  XNOR U7187 ( .A(n7359), .B(n7353), .Z(n7355) );
  XOR U7188 ( .A(n7361), .B(n7362), .Z(n7353) );
  AND U7189 ( .A(n263), .B(n7363), .Z(n7362) );
  XNOR U7190 ( .A(n7364), .B(n7365), .Z(n7359) );
  AND U7191 ( .A(n255), .B(n7366), .Z(n7365) );
  XOR U7192 ( .A(p_input[330]), .B(n7364), .Z(n7366) );
  XNOR U7193 ( .A(n7367), .B(n7368), .Z(n7364) );
  AND U7194 ( .A(n259), .B(n7363), .Z(n7368) );
  XNOR U7195 ( .A(n7367), .B(n7361), .Z(n7363) );
  XOR U7196 ( .A(n7369), .B(n7370), .Z(n7361) );
  AND U7197 ( .A(n274), .B(n7371), .Z(n7370) );
  XNOR U7198 ( .A(n7372), .B(n7373), .Z(n7367) );
  AND U7199 ( .A(n266), .B(n7374), .Z(n7373) );
  XOR U7200 ( .A(p_input[346]), .B(n7372), .Z(n7374) );
  XNOR U7201 ( .A(n7375), .B(n7376), .Z(n7372) );
  AND U7202 ( .A(n270), .B(n7371), .Z(n7376) );
  XNOR U7203 ( .A(n7375), .B(n7369), .Z(n7371) );
  XOR U7204 ( .A(n7377), .B(n7378), .Z(n7369) );
  AND U7205 ( .A(n285), .B(n7379), .Z(n7378) );
  XNOR U7206 ( .A(n7380), .B(n7381), .Z(n7375) );
  AND U7207 ( .A(n277), .B(n7382), .Z(n7381) );
  XOR U7208 ( .A(p_input[362]), .B(n7380), .Z(n7382) );
  XNOR U7209 ( .A(n7383), .B(n7384), .Z(n7380) );
  AND U7210 ( .A(n281), .B(n7379), .Z(n7384) );
  XNOR U7211 ( .A(n7383), .B(n7377), .Z(n7379) );
  XOR U7212 ( .A(n7385), .B(n7386), .Z(n7377) );
  AND U7213 ( .A(n296), .B(n7387), .Z(n7386) );
  XNOR U7214 ( .A(n7388), .B(n7389), .Z(n7383) );
  AND U7215 ( .A(n288), .B(n7390), .Z(n7389) );
  XOR U7216 ( .A(p_input[378]), .B(n7388), .Z(n7390) );
  XNOR U7217 ( .A(n7391), .B(n7392), .Z(n7388) );
  AND U7218 ( .A(n292), .B(n7387), .Z(n7392) );
  XNOR U7219 ( .A(n7391), .B(n7385), .Z(n7387) );
  XOR U7220 ( .A(n7393), .B(n7394), .Z(n7385) );
  AND U7221 ( .A(n307), .B(n7395), .Z(n7394) );
  XNOR U7222 ( .A(n7396), .B(n7397), .Z(n7391) );
  AND U7223 ( .A(n299), .B(n7398), .Z(n7397) );
  XOR U7224 ( .A(p_input[394]), .B(n7396), .Z(n7398) );
  XNOR U7225 ( .A(n7399), .B(n7400), .Z(n7396) );
  AND U7226 ( .A(n303), .B(n7395), .Z(n7400) );
  XNOR U7227 ( .A(n7399), .B(n7393), .Z(n7395) );
  XOR U7228 ( .A(n7401), .B(n7402), .Z(n7393) );
  AND U7229 ( .A(n318), .B(n7403), .Z(n7402) );
  XNOR U7230 ( .A(n7404), .B(n7405), .Z(n7399) );
  AND U7231 ( .A(n310), .B(n7406), .Z(n7405) );
  XOR U7232 ( .A(p_input[410]), .B(n7404), .Z(n7406) );
  XNOR U7233 ( .A(n7407), .B(n7408), .Z(n7404) );
  AND U7234 ( .A(n314), .B(n7403), .Z(n7408) );
  XNOR U7235 ( .A(n7407), .B(n7401), .Z(n7403) );
  XOR U7236 ( .A(n7409), .B(n7410), .Z(n7401) );
  AND U7237 ( .A(n329), .B(n7411), .Z(n7410) );
  XNOR U7238 ( .A(n7412), .B(n7413), .Z(n7407) );
  AND U7239 ( .A(n321), .B(n7414), .Z(n7413) );
  XOR U7240 ( .A(p_input[426]), .B(n7412), .Z(n7414) );
  XNOR U7241 ( .A(n7415), .B(n7416), .Z(n7412) );
  AND U7242 ( .A(n325), .B(n7411), .Z(n7416) );
  XNOR U7243 ( .A(n7415), .B(n7409), .Z(n7411) );
  XOR U7244 ( .A(n7417), .B(n7418), .Z(n7409) );
  AND U7245 ( .A(n340), .B(n7419), .Z(n7418) );
  XNOR U7246 ( .A(n7420), .B(n7421), .Z(n7415) );
  AND U7247 ( .A(n332), .B(n7422), .Z(n7421) );
  XOR U7248 ( .A(p_input[442]), .B(n7420), .Z(n7422) );
  XNOR U7249 ( .A(n7423), .B(n7424), .Z(n7420) );
  AND U7250 ( .A(n336), .B(n7419), .Z(n7424) );
  XNOR U7251 ( .A(n7423), .B(n7417), .Z(n7419) );
  XOR U7252 ( .A(n7425), .B(n7426), .Z(n7417) );
  AND U7253 ( .A(n351), .B(n7427), .Z(n7426) );
  XNOR U7254 ( .A(n7428), .B(n7429), .Z(n7423) );
  AND U7255 ( .A(n343), .B(n7430), .Z(n7429) );
  XOR U7256 ( .A(p_input[458]), .B(n7428), .Z(n7430) );
  XNOR U7257 ( .A(n7431), .B(n7432), .Z(n7428) );
  AND U7258 ( .A(n347), .B(n7427), .Z(n7432) );
  XNOR U7259 ( .A(n7431), .B(n7425), .Z(n7427) );
  XOR U7260 ( .A(n7433), .B(n7434), .Z(n7425) );
  AND U7261 ( .A(n362), .B(n7435), .Z(n7434) );
  XNOR U7262 ( .A(n7436), .B(n7437), .Z(n7431) );
  AND U7263 ( .A(n354), .B(n7438), .Z(n7437) );
  XOR U7264 ( .A(p_input[474]), .B(n7436), .Z(n7438) );
  XNOR U7265 ( .A(n7439), .B(n7440), .Z(n7436) );
  AND U7266 ( .A(n358), .B(n7435), .Z(n7440) );
  XNOR U7267 ( .A(n7439), .B(n7433), .Z(n7435) );
  XOR U7268 ( .A(n7441), .B(n7442), .Z(n7433) );
  AND U7269 ( .A(n373), .B(n7443), .Z(n7442) );
  XNOR U7270 ( .A(n7444), .B(n7445), .Z(n7439) );
  AND U7271 ( .A(n365), .B(n7446), .Z(n7445) );
  XOR U7272 ( .A(p_input[490]), .B(n7444), .Z(n7446) );
  XNOR U7273 ( .A(n7447), .B(n7448), .Z(n7444) );
  AND U7274 ( .A(n369), .B(n7443), .Z(n7448) );
  XNOR U7275 ( .A(n7447), .B(n7441), .Z(n7443) );
  XOR U7276 ( .A(n7449), .B(n7450), .Z(n7441) );
  AND U7277 ( .A(n384), .B(n7451), .Z(n7450) );
  XNOR U7278 ( .A(n7452), .B(n7453), .Z(n7447) );
  AND U7279 ( .A(n376), .B(n7454), .Z(n7453) );
  XOR U7280 ( .A(p_input[506]), .B(n7452), .Z(n7454) );
  XNOR U7281 ( .A(n7455), .B(n7456), .Z(n7452) );
  AND U7282 ( .A(n380), .B(n7451), .Z(n7456) );
  XNOR U7283 ( .A(n7455), .B(n7449), .Z(n7451) );
  XOR U7284 ( .A(n7457), .B(n7458), .Z(n7449) );
  AND U7285 ( .A(n395), .B(n7459), .Z(n7458) );
  XNOR U7286 ( .A(n7460), .B(n7461), .Z(n7455) );
  AND U7287 ( .A(n387), .B(n7462), .Z(n7461) );
  XOR U7288 ( .A(p_input[522]), .B(n7460), .Z(n7462) );
  XNOR U7289 ( .A(n7463), .B(n7464), .Z(n7460) );
  AND U7290 ( .A(n391), .B(n7459), .Z(n7464) );
  XNOR U7291 ( .A(n7463), .B(n7457), .Z(n7459) );
  XOR U7292 ( .A(n7465), .B(n7466), .Z(n7457) );
  AND U7293 ( .A(n406), .B(n7467), .Z(n7466) );
  XNOR U7294 ( .A(n7468), .B(n7469), .Z(n7463) );
  AND U7295 ( .A(n398), .B(n7470), .Z(n7469) );
  XOR U7296 ( .A(p_input[538]), .B(n7468), .Z(n7470) );
  XNOR U7297 ( .A(n7471), .B(n7472), .Z(n7468) );
  AND U7298 ( .A(n402), .B(n7467), .Z(n7472) );
  XNOR U7299 ( .A(n7471), .B(n7465), .Z(n7467) );
  XOR U7300 ( .A(n7473), .B(n7474), .Z(n7465) );
  AND U7301 ( .A(n417), .B(n7475), .Z(n7474) );
  XNOR U7302 ( .A(n7476), .B(n7477), .Z(n7471) );
  AND U7303 ( .A(n409), .B(n7478), .Z(n7477) );
  XOR U7304 ( .A(p_input[554]), .B(n7476), .Z(n7478) );
  XNOR U7305 ( .A(n7479), .B(n7480), .Z(n7476) );
  AND U7306 ( .A(n413), .B(n7475), .Z(n7480) );
  XNOR U7307 ( .A(n7479), .B(n7473), .Z(n7475) );
  XOR U7308 ( .A(n7481), .B(n7482), .Z(n7473) );
  AND U7309 ( .A(n428), .B(n7483), .Z(n7482) );
  XNOR U7310 ( .A(n7484), .B(n7485), .Z(n7479) );
  AND U7311 ( .A(n420), .B(n7486), .Z(n7485) );
  XOR U7312 ( .A(p_input[570]), .B(n7484), .Z(n7486) );
  XNOR U7313 ( .A(n7487), .B(n7488), .Z(n7484) );
  AND U7314 ( .A(n424), .B(n7483), .Z(n7488) );
  XNOR U7315 ( .A(n7487), .B(n7481), .Z(n7483) );
  XOR U7316 ( .A(n7489), .B(n7490), .Z(n7481) );
  AND U7317 ( .A(n439), .B(n7491), .Z(n7490) );
  XNOR U7318 ( .A(n7492), .B(n7493), .Z(n7487) );
  AND U7319 ( .A(n431), .B(n7494), .Z(n7493) );
  XOR U7320 ( .A(p_input[586]), .B(n7492), .Z(n7494) );
  XNOR U7321 ( .A(n7495), .B(n7496), .Z(n7492) );
  AND U7322 ( .A(n435), .B(n7491), .Z(n7496) );
  XNOR U7323 ( .A(n7495), .B(n7489), .Z(n7491) );
  XOR U7324 ( .A(n7497), .B(n7498), .Z(n7489) );
  AND U7325 ( .A(n450), .B(n7499), .Z(n7498) );
  XNOR U7326 ( .A(n7500), .B(n7501), .Z(n7495) );
  AND U7327 ( .A(n442), .B(n7502), .Z(n7501) );
  XOR U7328 ( .A(p_input[602]), .B(n7500), .Z(n7502) );
  XNOR U7329 ( .A(n7503), .B(n7504), .Z(n7500) );
  AND U7330 ( .A(n446), .B(n7499), .Z(n7504) );
  XNOR U7331 ( .A(n7503), .B(n7497), .Z(n7499) );
  XOR U7332 ( .A(n7505), .B(n7506), .Z(n7497) );
  AND U7333 ( .A(n461), .B(n7507), .Z(n7506) );
  XNOR U7334 ( .A(n7508), .B(n7509), .Z(n7503) );
  AND U7335 ( .A(n453), .B(n7510), .Z(n7509) );
  XOR U7336 ( .A(p_input[618]), .B(n7508), .Z(n7510) );
  XNOR U7337 ( .A(n7511), .B(n7512), .Z(n7508) );
  AND U7338 ( .A(n457), .B(n7507), .Z(n7512) );
  XNOR U7339 ( .A(n7511), .B(n7505), .Z(n7507) );
  XOR U7340 ( .A(n7513), .B(n7514), .Z(n7505) );
  AND U7341 ( .A(n472), .B(n7515), .Z(n7514) );
  XNOR U7342 ( .A(n7516), .B(n7517), .Z(n7511) );
  AND U7343 ( .A(n464), .B(n7518), .Z(n7517) );
  XOR U7344 ( .A(p_input[634]), .B(n7516), .Z(n7518) );
  XNOR U7345 ( .A(n7519), .B(n7520), .Z(n7516) );
  AND U7346 ( .A(n468), .B(n7515), .Z(n7520) );
  XNOR U7347 ( .A(n7519), .B(n7513), .Z(n7515) );
  XOR U7348 ( .A(n7521), .B(n7522), .Z(n7513) );
  AND U7349 ( .A(n483), .B(n7523), .Z(n7522) );
  XNOR U7350 ( .A(n7524), .B(n7525), .Z(n7519) );
  AND U7351 ( .A(n475), .B(n7526), .Z(n7525) );
  XOR U7352 ( .A(p_input[650]), .B(n7524), .Z(n7526) );
  XNOR U7353 ( .A(n7527), .B(n7528), .Z(n7524) );
  AND U7354 ( .A(n479), .B(n7523), .Z(n7528) );
  XNOR U7355 ( .A(n7527), .B(n7521), .Z(n7523) );
  XOR U7356 ( .A(n7529), .B(n7530), .Z(n7521) );
  AND U7357 ( .A(n494), .B(n7531), .Z(n7530) );
  XNOR U7358 ( .A(n7532), .B(n7533), .Z(n7527) );
  AND U7359 ( .A(n486), .B(n7534), .Z(n7533) );
  XOR U7360 ( .A(p_input[666]), .B(n7532), .Z(n7534) );
  XNOR U7361 ( .A(n7535), .B(n7536), .Z(n7532) );
  AND U7362 ( .A(n490), .B(n7531), .Z(n7536) );
  XNOR U7363 ( .A(n7535), .B(n7529), .Z(n7531) );
  XOR U7364 ( .A(n7537), .B(n7538), .Z(n7529) );
  AND U7365 ( .A(n505), .B(n7539), .Z(n7538) );
  XNOR U7366 ( .A(n7540), .B(n7541), .Z(n7535) );
  AND U7367 ( .A(n497), .B(n7542), .Z(n7541) );
  XOR U7368 ( .A(p_input[682]), .B(n7540), .Z(n7542) );
  XNOR U7369 ( .A(n7543), .B(n7544), .Z(n7540) );
  AND U7370 ( .A(n501), .B(n7539), .Z(n7544) );
  XNOR U7371 ( .A(n7543), .B(n7537), .Z(n7539) );
  XOR U7372 ( .A(n7545), .B(n7546), .Z(n7537) );
  AND U7373 ( .A(n516), .B(n7547), .Z(n7546) );
  XNOR U7374 ( .A(n7548), .B(n7549), .Z(n7543) );
  AND U7375 ( .A(n508), .B(n7550), .Z(n7549) );
  XOR U7376 ( .A(p_input[698]), .B(n7548), .Z(n7550) );
  XNOR U7377 ( .A(n7551), .B(n7552), .Z(n7548) );
  AND U7378 ( .A(n512), .B(n7547), .Z(n7552) );
  XNOR U7379 ( .A(n7551), .B(n7545), .Z(n7547) );
  XOR U7380 ( .A(n7553), .B(n7554), .Z(n7545) );
  AND U7381 ( .A(n527), .B(n7555), .Z(n7554) );
  XNOR U7382 ( .A(n7556), .B(n7557), .Z(n7551) );
  AND U7383 ( .A(n519), .B(n7558), .Z(n7557) );
  XOR U7384 ( .A(p_input[714]), .B(n7556), .Z(n7558) );
  XNOR U7385 ( .A(n7559), .B(n7560), .Z(n7556) );
  AND U7386 ( .A(n523), .B(n7555), .Z(n7560) );
  XNOR U7387 ( .A(n7559), .B(n7553), .Z(n7555) );
  XOR U7388 ( .A(n7561), .B(n7562), .Z(n7553) );
  AND U7389 ( .A(n538), .B(n7563), .Z(n7562) );
  XNOR U7390 ( .A(n7564), .B(n7565), .Z(n7559) );
  AND U7391 ( .A(n530), .B(n7566), .Z(n7565) );
  XOR U7392 ( .A(p_input[730]), .B(n7564), .Z(n7566) );
  XNOR U7393 ( .A(n7567), .B(n7568), .Z(n7564) );
  AND U7394 ( .A(n534), .B(n7563), .Z(n7568) );
  XNOR U7395 ( .A(n7567), .B(n7561), .Z(n7563) );
  XOR U7396 ( .A(n7569), .B(n7570), .Z(n7561) );
  AND U7397 ( .A(n549), .B(n7571), .Z(n7570) );
  XNOR U7398 ( .A(n7572), .B(n7573), .Z(n7567) );
  AND U7399 ( .A(n541), .B(n7574), .Z(n7573) );
  XOR U7400 ( .A(p_input[746]), .B(n7572), .Z(n7574) );
  XNOR U7401 ( .A(n7575), .B(n7576), .Z(n7572) );
  AND U7402 ( .A(n545), .B(n7571), .Z(n7576) );
  XNOR U7403 ( .A(n7575), .B(n7569), .Z(n7571) );
  XOR U7404 ( .A(n7577), .B(n7578), .Z(n7569) );
  AND U7405 ( .A(n560), .B(n7579), .Z(n7578) );
  XNOR U7406 ( .A(n7580), .B(n7581), .Z(n7575) );
  AND U7407 ( .A(n552), .B(n7582), .Z(n7581) );
  XOR U7408 ( .A(p_input[762]), .B(n7580), .Z(n7582) );
  XNOR U7409 ( .A(n7583), .B(n7584), .Z(n7580) );
  AND U7410 ( .A(n556), .B(n7579), .Z(n7584) );
  XNOR U7411 ( .A(n7583), .B(n7577), .Z(n7579) );
  XOR U7412 ( .A(n7585), .B(n7586), .Z(n7577) );
  AND U7413 ( .A(n571), .B(n7587), .Z(n7586) );
  XNOR U7414 ( .A(n7588), .B(n7589), .Z(n7583) );
  AND U7415 ( .A(n563), .B(n7590), .Z(n7589) );
  XOR U7416 ( .A(p_input[778]), .B(n7588), .Z(n7590) );
  XNOR U7417 ( .A(n7591), .B(n7592), .Z(n7588) );
  AND U7418 ( .A(n567), .B(n7587), .Z(n7592) );
  XNOR U7419 ( .A(n7591), .B(n7585), .Z(n7587) );
  XOR U7420 ( .A(n7593), .B(n7594), .Z(n7585) );
  AND U7421 ( .A(n582), .B(n7595), .Z(n7594) );
  XNOR U7422 ( .A(n7596), .B(n7597), .Z(n7591) );
  AND U7423 ( .A(n574), .B(n7598), .Z(n7597) );
  XOR U7424 ( .A(p_input[794]), .B(n7596), .Z(n7598) );
  XNOR U7425 ( .A(n7599), .B(n7600), .Z(n7596) );
  AND U7426 ( .A(n578), .B(n7595), .Z(n7600) );
  XNOR U7427 ( .A(n7599), .B(n7593), .Z(n7595) );
  XOR U7428 ( .A(n7601), .B(n7602), .Z(n7593) );
  AND U7429 ( .A(n593), .B(n7603), .Z(n7602) );
  XNOR U7430 ( .A(n7604), .B(n7605), .Z(n7599) );
  AND U7431 ( .A(n585), .B(n7606), .Z(n7605) );
  XOR U7432 ( .A(p_input[810]), .B(n7604), .Z(n7606) );
  XNOR U7433 ( .A(n7607), .B(n7608), .Z(n7604) );
  AND U7434 ( .A(n589), .B(n7603), .Z(n7608) );
  XNOR U7435 ( .A(n7607), .B(n7601), .Z(n7603) );
  XOR U7436 ( .A(n7609), .B(n7610), .Z(n7601) );
  AND U7437 ( .A(n604), .B(n7611), .Z(n7610) );
  XNOR U7438 ( .A(n7612), .B(n7613), .Z(n7607) );
  AND U7439 ( .A(n596), .B(n7614), .Z(n7613) );
  XOR U7440 ( .A(p_input[826]), .B(n7612), .Z(n7614) );
  XNOR U7441 ( .A(n7615), .B(n7616), .Z(n7612) );
  AND U7442 ( .A(n600), .B(n7611), .Z(n7616) );
  XNOR U7443 ( .A(n7615), .B(n7609), .Z(n7611) );
  XOR U7444 ( .A(n7617), .B(n7618), .Z(n7609) );
  AND U7445 ( .A(n615), .B(n7619), .Z(n7618) );
  XNOR U7446 ( .A(n7620), .B(n7621), .Z(n7615) );
  AND U7447 ( .A(n607), .B(n7622), .Z(n7621) );
  XOR U7448 ( .A(p_input[842]), .B(n7620), .Z(n7622) );
  XNOR U7449 ( .A(n7623), .B(n7624), .Z(n7620) );
  AND U7450 ( .A(n611), .B(n7619), .Z(n7624) );
  XNOR U7451 ( .A(n7623), .B(n7617), .Z(n7619) );
  XOR U7452 ( .A(n7625), .B(n7626), .Z(n7617) );
  AND U7453 ( .A(n626), .B(n7627), .Z(n7626) );
  XNOR U7454 ( .A(n7628), .B(n7629), .Z(n7623) );
  AND U7455 ( .A(n618), .B(n7630), .Z(n7629) );
  XOR U7456 ( .A(p_input[858]), .B(n7628), .Z(n7630) );
  XNOR U7457 ( .A(n7631), .B(n7632), .Z(n7628) );
  AND U7458 ( .A(n622), .B(n7627), .Z(n7632) );
  XNOR U7459 ( .A(n7631), .B(n7625), .Z(n7627) );
  XOR U7460 ( .A(n7633), .B(n7634), .Z(n7625) );
  AND U7461 ( .A(n637), .B(n7635), .Z(n7634) );
  XNOR U7462 ( .A(n7636), .B(n7637), .Z(n7631) );
  AND U7463 ( .A(n629), .B(n7638), .Z(n7637) );
  XOR U7464 ( .A(p_input[874]), .B(n7636), .Z(n7638) );
  XNOR U7465 ( .A(n7639), .B(n7640), .Z(n7636) );
  AND U7466 ( .A(n633), .B(n7635), .Z(n7640) );
  XNOR U7467 ( .A(n7639), .B(n7633), .Z(n7635) );
  XOR U7468 ( .A(n7641), .B(n7642), .Z(n7633) );
  AND U7469 ( .A(n648), .B(n7643), .Z(n7642) );
  XNOR U7470 ( .A(n7644), .B(n7645), .Z(n7639) );
  AND U7471 ( .A(n640), .B(n7646), .Z(n7645) );
  XOR U7472 ( .A(p_input[890]), .B(n7644), .Z(n7646) );
  XNOR U7473 ( .A(n7647), .B(n7648), .Z(n7644) );
  AND U7474 ( .A(n644), .B(n7643), .Z(n7648) );
  XNOR U7475 ( .A(n7647), .B(n7641), .Z(n7643) );
  XOR U7476 ( .A(n7649), .B(n7650), .Z(n7641) );
  AND U7477 ( .A(n659), .B(n7651), .Z(n7650) );
  XNOR U7478 ( .A(n7652), .B(n7653), .Z(n7647) );
  AND U7479 ( .A(n651), .B(n7654), .Z(n7653) );
  XOR U7480 ( .A(p_input[906]), .B(n7652), .Z(n7654) );
  XNOR U7481 ( .A(n7655), .B(n7656), .Z(n7652) );
  AND U7482 ( .A(n655), .B(n7651), .Z(n7656) );
  XNOR U7483 ( .A(n7655), .B(n7649), .Z(n7651) );
  XOR U7484 ( .A(n7657), .B(n7658), .Z(n7649) );
  AND U7485 ( .A(n670), .B(n7659), .Z(n7658) );
  XNOR U7486 ( .A(n7660), .B(n7661), .Z(n7655) );
  AND U7487 ( .A(n662), .B(n7662), .Z(n7661) );
  XOR U7488 ( .A(p_input[922]), .B(n7660), .Z(n7662) );
  XNOR U7489 ( .A(n7663), .B(n7664), .Z(n7660) );
  AND U7490 ( .A(n666), .B(n7659), .Z(n7664) );
  XNOR U7491 ( .A(n7663), .B(n7657), .Z(n7659) );
  XOR U7492 ( .A(n7665), .B(n7666), .Z(n7657) );
  AND U7493 ( .A(n681), .B(n7667), .Z(n7666) );
  XNOR U7494 ( .A(n7668), .B(n7669), .Z(n7663) );
  AND U7495 ( .A(n673), .B(n7670), .Z(n7669) );
  XOR U7496 ( .A(p_input[938]), .B(n7668), .Z(n7670) );
  XNOR U7497 ( .A(n7671), .B(n7672), .Z(n7668) );
  AND U7498 ( .A(n677), .B(n7667), .Z(n7672) );
  XNOR U7499 ( .A(n7671), .B(n7665), .Z(n7667) );
  XOR U7500 ( .A(n7673), .B(n7674), .Z(n7665) );
  AND U7501 ( .A(n692), .B(n7675), .Z(n7674) );
  XNOR U7502 ( .A(n7676), .B(n7677), .Z(n7671) );
  AND U7503 ( .A(n684), .B(n7678), .Z(n7677) );
  XOR U7504 ( .A(p_input[954]), .B(n7676), .Z(n7678) );
  XNOR U7505 ( .A(n7679), .B(n7680), .Z(n7676) );
  AND U7506 ( .A(n688), .B(n7675), .Z(n7680) );
  XNOR U7507 ( .A(n7679), .B(n7673), .Z(n7675) );
  XOR U7508 ( .A(n7681), .B(n7682), .Z(n7673) );
  AND U7509 ( .A(n703), .B(n7683), .Z(n7682) );
  XNOR U7510 ( .A(n7684), .B(n7685), .Z(n7679) );
  AND U7511 ( .A(n695), .B(n7686), .Z(n7685) );
  XOR U7512 ( .A(p_input[970]), .B(n7684), .Z(n7686) );
  XNOR U7513 ( .A(n7687), .B(n7688), .Z(n7684) );
  AND U7514 ( .A(n699), .B(n7683), .Z(n7688) );
  XNOR U7515 ( .A(n7687), .B(n7681), .Z(n7683) );
  XOR U7516 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n7689), .Z(n7681) );
  AND U7517 ( .A(n713), .B(n7690), .Z(n7689) );
  XNOR U7518 ( .A(n7691), .B(n7692), .Z(n7687) );
  AND U7519 ( .A(n706), .B(n7693), .Z(n7692) );
  XOR U7520 ( .A(p_input[986]), .B(n7691), .Z(n7693) );
  XNOR U7521 ( .A(n7694), .B(n7695), .Z(n7691) );
  AND U7522 ( .A(n710), .B(n7690), .Z(n7695) );
  XOR U7523 ( .A(\knn_comb_/min_val_out[0][10] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n7690) );
  IV U7524 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n7694) );
  XOR U7525 ( .A(n4709), .B(n7696), .Z(o[0]) );
  AND U7526 ( .A(n30), .B(n7697), .Z(n4709) );
  XOR U7527 ( .A(n4710), .B(n7696), .Z(n7697) );
  XOR U7528 ( .A(n7698), .B(n7699), .Z(n7696) );
  AND U7529 ( .A(n42), .B(n7700), .Z(n7699) );
  XOR U7530 ( .A(n7701), .B(n7702), .Z(n4710) );
  AND U7531 ( .A(n34), .B(n7703), .Z(n7702) );
  XOR U7532 ( .A(p_input[0]), .B(n7701), .Z(n7703) );
  XNOR U7533 ( .A(n7704), .B(n7705), .Z(n7701) );
  AND U7534 ( .A(n38), .B(n7700), .Z(n7705) );
  XNOR U7535 ( .A(n7704), .B(n7698), .Z(n7700) );
  XOR U7536 ( .A(n7706), .B(n7707), .Z(n7698) );
  AND U7537 ( .A(n54), .B(n7708), .Z(n7707) );
  XNOR U7538 ( .A(n7709), .B(n7710), .Z(n7704) );
  AND U7539 ( .A(n46), .B(n7711), .Z(n7710) );
  XOR U7540 ( .A(p_input[16]), .B(n7709), .Z(n7711) );
  XNOR U7541 ( .A(n7712), .B(n7713), .Z(n7709) );
  AND U7542 ( .A(n50), .B(n7708), .Z(n7713) );
  XNOR U7543 ( .A(n7712), .B(n7706), .Z(n7708) );
  XOR U7544 ( .A(n7714), .B(n7715), .Z(n7706) );
  AND U7545 ( .A(n65), .B(n7716), .Z(n7715) );
  XNOR U7546 ( .A(n7717), .B(n7718), .Z(n7712) );
  AND U7547 ( .A(n57), .B(n7719), .Z(n7718) );
  XOR U7548 ( .A(p_input[32]), .B(n7717), .Z(n7719) );
  XNOR U7549 ( .A(n7720), .B(n7721), .Z(n7717) );
  AND U7550 ( .A(n61), .B(n7716), .Z(n7721) );
  XNOR U7551 ( .A(n7720), .B(n7714), .Z(n7716) );
  XOR U7552 ( .A(n7722), .B(n7723), .Z(n7714) );
  AND U7553 ( .A(n76), .B(n7724), .Z(n7723) );
  XNOR U7554 ( .A(n7725), .B(n7726), .Z(n7720) );
  AND U7555 ( .A(n68), .B(n7727), .Z(n7726) );
  XOR U7556 ( .A(p_input[48]), .B(n7725), .Z(n7727) );
  XNOR U7557 ( .A(n7728), .B(n7729), .Z(n7725) );
  AND U7558 ( .A(n72), .B(n7724), .Z(n7729) );
  XNOR U7559 ( .A(n7728), .B(n7722), .Z(n7724) );
  XOR U7560 ( .A(n7730), .B(n7731), .Z(n7722) );
  AND U7561 ( .A(n87), .B(n7732), .Z(n7731) );
  XNOR U7562 ( .A(n7733), .B(n7734), .Z(n7728) );
  AND U7563 ( .A(n79), .B(n7735), .Z(n7734) );
  XOR U7564 ( .A(p_input[64]), .B(n7733), .Z(n7735) );
  XNOR U7565 ( .A(n7736), .B(n7737), .Z(n7733) );
  AND U7566 ( .A(n83), .B(n7732), .Z(n7737) );
  XNOR U7567 ( .A(n7736), .B(n7730), .Z(n7732) );
  XOR U7568 ( .A(n7738), .B(n7739), .Z(n7730) );
  AND U7569 ( .A(n98), .B(n7740), .Z(n7739) );
  XNOR U7570 ( .A(n7741), .B(n7742), .Z(n7736) );
  AND U7571 ( .A(n90), .B(n7743), .Z(n7742) );
  XOR U7572 ( .A(p_input[80]), .B(n7741), .Z(n7743) );
  XNOR U7573 ( .A(n7744), .B(n7745), .Z(n7741) );
  AND U7574 ( .A(n94), .B(n7740), .Z(n7745) );
  XNOR U7575 ( .A(n7744), .B(n7738), .Z(n7740) );
  XOR U7576 ( .A(n7746), .B(n7747), .Z(n7738) );
  AND U7577 ( .A(n109), .B(n7748), .Z(n7747) );
  XNOR U7578 ( .A(n7749), .B(n7750), .Z(n7744) );
  AND U7579 ( .A(n101), .B(n7751), .Z(n7750) );
  XOR U7580 ( .A(p_input[96]), .B(n7749), .Z(n7751) );
  XNOR U7581 ( .A(n7752), .B(n7753), .Z(n7749) );
  AND U7582 ( .A(n105), .B(n7748), .Z(n7753) );
  XNOR U7583 ( .A(n7752), .B(n7746), .Z(n7748) );
  XOR U7584 ( .A(n7754), .B(n7755), .Z(n7746) );
  AND U7585 ( .A(n120), .B(n7756), .Z(n7755) );
  XNOR U7586 ( .A(n7757), .B(n7758), .Z(n7752) );
  AND U7587 ( .A(n112), .B(n7759), .Z(n7758) );
  XOR U7588 ( .A(p_input[112]), .B(n7757), .Z(n7759) );
  XNOR U7589 ( .A(n7760), .B(n7761), .Z(n7757) );
  AND U7590 ( .A(n116), .B(n7756), .Z(n7761) );
  XNOR U7591 ( .A(n7760), .B(n7754), .Z(n7756) );
  XOR U7592 ( .A(n7762), .B(n7763), .Z(n7754) );
  AND U7593 ( .A(n131), .B(n7764), .Z(n7763) );
  XNOR U7594 ( .A(n7765), .B(n7766), .Z(n7760) );
  AND U7595 ( .A(n123), .B(n7767), .Z(n7766) );
  XOR U7596 ( .A(p_input[128]), .B(n7765), .Z(n7767) );
  XNOR U7597 ( .A(n7768), .B(n7769), .Z(n7765) );
  AND U7598 ( .A(n127), .B(n7764), .Z(n7769) );
  XNOR U7599 ( .A(n7768), .B(n7762), .Z(n7764) );
  XOR U7600 ( .A(n7770), .B(n7771), .Z(n7762) );
  AND U7601 ( .A(n142), .B(n7772), .Z(n7771) );
  XNOR U7602 ( .A(n7773), .B(n7774), .Z(n7768) );
  AND U7603 ( .A(n134), .B(n7775), .Z(n7774) );
  XOR U7604 ( .A(p_input[144]), .B(n7773), .Z(n7775) );
  XNOR U7605 ( .A(n7776), .B(n7777), .Z(n7773) );
  AND U7606 ( .A(n138), .B(n7772), .Z(n7777) );
  XNOR U7607 ( .A(n7776), .B(n7770), .Z(n7772) );
  XOR U7608 ( .A(n7778), .B(n7779), .Z(n7770) );
  AND U7609 ( .A(n153), .B(n7780), .Z(n7779) );
  XNOR U7610 ( .A(n7781), .B(n7782), .Z(n7776) );
  AND U7611 ( .A(n145), .B(n7783), .Z(n7782) );
  XOR U7612 ( .A(p_input[160]), .B(n7781), .Z(n7783) );
  XNOR U7613 ( .A(n7784), .B(n7785), .Z(n7781) );
  AND U7614 ( .A(n149), .B(n7780), .Z(n7785) );
  XNOR U7615 ( .A(n7784), .B(n7778), .Z(n7780) );
  XOR U7616 ( .A(n7786), .B(n7787), .Z(n7778) );
  AND U7617 ( .A(n164), .B(n7788), .Z(n7787) );
  XNOR U7618 ( .A(n7789), .B(n7790), .Z(n7784) );
  AND U7619 ( .A(n156), .B(n7791), .Z(n7790) );
  XOR U7620 ( .A(p_input[176]), .B(n7789), .Z(n7791) );
  XNOR U7621 ( .A(n7792), .B(n7793), .Z(n7789) );
  AND U7622 ( .A(n160), .B(n7788), .Z(n7793) );
  XNOR U7623 ( .A(n7792), .B(n7786), .Z(n7788) );
  XOR U7624 ( .A(n7794), .B(n7795), .Z(n7786) );
  AND U7625 ( .A(n175), .B(n7796), .Z(n7795) );
  XNOR U7626 ( .A(n7797), .B(n7798), .Z(n7792) );
  AND U7627 ( .A(n167), .B(n7799), .Z(n7798) );
  XOR U7628 ( .A(p_input[192]), .B(n7797), .Z(n7799) );
  XNOR U7629 ( .A(n7800), .B(n7801), .Z(n7797) );
  AND U7630 ( .A(n171), .B(n7796), .Z(n7801) );
  XNOR U7631 ( .A(n7800), .B(n7794), .Z(n7796) );
  XOR U7632 ( .A(n7802), .B(n7803), .Z(n7794) );
  AND U7633 ( .A(n186), .B(n7804), .Z(n7803) );
  XNOR U7634 ( .A(n7805), .B(n7806), .Z(n7800) );
  AND U7635 ( .A(n178), .B(n7807), .Z(n7806) );
  XOR U7636 ( .A(p_input[208]), .B(n7805), .Z(n7807) );
  XNOR U7637 ( .A(n7808), .B(n7809), .Z(n7805) );
  AND U7638 ( .A(n182), .B(n7804), .Z(n7809) );
  XNOR U7639 ( .A(n7808), .B(n7802), .Z(n7804) );
  XOR U7640 ( .A(n7810), .B(n7811), .Z(n7802) );
  AND U7641 ( .A(n197), .B(n7812), .Z(n7811) );
  XNOR U7642 ( .A(n7813), .B(n7814), .Z(n7808) );
  AND U7643 ( .A(n189), .B(n7815), .Z(n7814) );
  XOR U7644 ( .A(p_input[224]), .B(n7813), .Z(n7815) );
  XNOR U7645 ( .A(n7816), .B(n7817), .Z(n7813) );
  AND U7646 ( .A(n193), .B(n7812), .Z(n7817) );
  XNOR U7647 ( .A(n7816), .B(n7810), .Z(n7812) );
  XOR U7648 ( .A(n7818), .B(n7819), .Z(n7810) );
  AND U7649 ( .A(n208), .B(n7820), .Z(n7819) );
  XNOR U7650 ( .A(n7821), .B(n7822), .Z(n7816) );
  AND U7651 ( .A(n200), .B(n7823), .Z(n7822) );
  XOR U7652 ( .A(p_input[240]), .B(n7821), .Z(n7823) );
  XNOR U7653 ( .A(n7824), .B(n7825), .Z(n7821) );
  AND U7654 ( .A(n204), .B(n7820), .Z(n7825) );
  XNOR U7655 ( .A(n7824), .B(n7818), .Z(n7820) );
  XOR U7656 ( .A(n7826), .B(n7827), .Z(n7818) );
  AND U7657 ( .A(n219), .B(n7828), .Z(n7827) );
  XNOR U7658 ( .A(n7829), .B(n7830), .Z(n7824) );
  AND U7659 ( .A(n211), .B(n7831), .Z(n7830) );
  XOR U7660 ( .A(p_input[256]), .B(n7829), .Z(n7831) );
  XNOR U7661 ( .A(n7832), .B(n7833), .Z(n7829) );
  AND U7662 ( .A(n215), .B(n7828), .Z(n7833) );
  XNOR U7663 ( .A(n7832), .B(n7826), .Z(n7828) );
  XOR U7664 ( .A(n7834), .B(n7835), .Z(n7826) );
  AND U7665 ( .A(n230), .B(n7836), .Z(n7835) );
  XNOR U7666 ( .A(n7837), .B(n7838), .Z(n7832) );
  AND U7667 ( .A(n222), .B(n7839), .Z(n7838) );
  XOR U7668 ( .A(p_input[272]), .B(n7837), .Z(n7839) );
  XNOR U7669 ( .A(n7840), .B(n7841), .Z(n7837) );
  AND U7670 ( .A(n226), .B(n7836), .Z(n7841) );
  XNOR U7671 ( .A(n7840), .B(n7834), .Z(n7836) );
  XOR U7672 ( .A(n7842), .B(n7843), .Z(n7834) );
  AND U7673 ( .A(n241), .B(n7844), .Z(n7843) );
  XNOR U7674 ( .A(n7845), .B(n7846), .Z(n7840) );
  AND U7675 ( .A(n233), .B(n7847), .Z(n7846) );
  XOR U7676 ( .A(p_input[288]), .B(n7845), .Z(n7847) );
  XNOR U7677 ( .A(n7848), .B(n7849), .Z(n7845) );
  AND U7678 ( .A(n237), .B(n7844), .Z(n7849) );
  XNOR U7679 ( .A(n7848), .B(n7842), .Z(n7844) );
  XOR U7680 ( .A(n7850), .B(n7851), .Z(n7842) );
  AND U7681 ( .A(n252), .B(n7852), .Z(n7851) );
  XNOR U7682 ( .A(n7853), .B(n7854), .Z(n7848) );
  AND U7683 ( .A(n244), .B(n7855), .Z(n7854) );
  XOR U7684 ( .A(p_input[304]), .B(n7853), .Z(n7855) );
  XNOR U7685 ( .A(n7856), .B(n7857), .Z(n7853) );
  AND U7686 ( .A(n248), .B(n7852), .Z(n7857) );
  XNOR U7687 ( .A(n7856), .B(n7850), .Z(n7852) );
  XOR U7688 ( .A(n7858), .B(n7859), .Z(n7850) );
  AND U7689 ( .A(n263), .B(n7860), .Z(n7859) );
  XNOR U7690 ( .A(n7861), .B(n7862), .Z(n7856) );
  AND U7691 ( .A(n255), .B(n7863), .Z(n7862) );
  XOR U7692 ( .A(p_input[320]), .B(n7861), .Z(n7863) );
  XNOR U7693 ( .A(n7864), .B(n7865), .Z(n7861) );
  AND U7694 ( .A(n259), .B(n7860), .Z(n7865) );
  XNOR U7695 ( .A(n7864), .B(n7858), .Z(n7860) );
  XOR U7696 ( .A(n7866), .B(n7867), .Z(n7858) );
  AND U7697 ( .A(n274), .B(n7868), .Z(n7867) );
  XNOR U7698 ( .A(n7869), .B(n7870), .Z(n7864) );
  AND U7699 ( .A(n266), .B(n7871), .Z(n7870) );
  XOR U7700 ( .A(p_input[336]), .B(n7869), .Z(n7871) );
  XNOR U7701 ( .A(n7872), .B(n7873), .Z(n7869) );
  AND U7702 ( .A(n270), .B(n7868), .Z(n7873) );
  XNOR U7703 ( .A(n7872), .B(n7866), .Z(n7868) );
  XOR U7704 ( .A(n7874), .B(n7875), .Z(n7866) );
  AND U7705 ( .A(n285), .B(n7876), .Z(n7875) );
  XNOR U7706 ( .A(n7877), .B(n7878), .Z(n7872) );
  AND U7707 ( .A(n277), .B(n7879), .Z(n7878) );
  XOR U7708 ( .A(p_input[352]), .B(n7877), .Z(n7879) );
  XNOR U7709 ( .A(n7880), .B(n7881), .Z(n7877) );
  AND U7710 ( .A(n281), .B(n7876), .Z(n7881) );
  XNOR U7711 ( .A(n7880), .B(n7874), .Z(n7876) );
  XOR U7712 ( .A(n7882), .B(n7883), .Z(n7874) );
  AND U7713 ( .A(n296), .B(n7884), .Z(n7883) );
  XNOR U7714 ( .A(n7885), .B(n7886), .Z(n7880) );
  AND U7715 ( .A(n288), .B(n7887), .Z(n7886) );
  XOR U7716 ( .A(p_input[368]), .B(n7885), .Z(n7887) );
  XNOR U7717 ( .A(n7888), .B(n7889), .Z(n7885) );
  AND U7718 ( .A(n292), .B(n7884), .Z(n7889) );
  XNOR U7719 ( .A(n7888), .B(n7882), .Z(n7884) );
  XOR U7720 ( .A(n7890), .B(n7891), .Z(n7882) );
  AND U7721 ( .A(n307), .B(n7892), .Z(n7891) );
  XNOR U7722 ( .A(n7893), .B(n7894), .Z(n7888) );
  AND U7723 ( .A(n299), .B(n7895), .Z(n7894) );
  XOR U7724 ( .A(p_input[384]), .B(n7893), .Z(n7895) );
  XNOR U7725 ( .A(n7896), .B(n7897), .Z(n7893) );
  AND U7726 ( .A(n303), .B(n7892), .Z(n7897) );
  XNOR U7727 ( .A(n7896), .B(n7890), .Z(n7892) );
  XOR U7728 ( .A(n7898), .B(n7899), .Z(n7890) );
  AND U7729 ( .A(n318), .B(n7900), .Z(n7899) );
  XNOR U7730 ( .A(n7901), .B(n7902), .Z(n7896) );
  AND U7731 ( .A(n310), .B(n7903), .Z(n7902) );
  XOR U7732 ( .A(p_input[400]), .B(n7901), .Z(n7903) );
  XNOR U7733 ( .A(n7904), .B(n7905), .Z(n7901) );
  AND U7734 ( .A(n314), .B(n7900), .Z(n7905) );
  XNOR U7735 ( .A(n7904), .B(n7898), .Z(n7900) );
  XOR U7736 ( .A(n7906), .B(n7907), .Z(n7898) );
  AND U7737 ( .A(n329), .B(n7908), .Z(n7907) );
  XNOR U7738 ( .A(n7909), .B(n7910), .Z(n7904) );
  AND U7739 ( .A(n321), .B(n7911), .Z(n7910) );
  XOR U7740 ( .A(p_input[416]), .B(n7909), .Z(n7911) );
  XNOR U7741 ( .A(n7912), .B(n7913), .Z(n7909) );
  AND U7742 ( .A(n325), .B(n7908), .Z(n7913) );
  XNOR U7743 ( .A(n7912), .B(n7906), .Z(n7908) );
  XOR U7744 ( .A(n7914), .B(n7915), .Z(n7906) );
  AND U7745 ( .A(n340), .B(n7916), .Z(n7915) );
  XNOR U7746 ( .A(n7917), .B(n7918), .Z(n7912) );
  AND U7747 ( .A(n332), .B(n7919), .Z(n7918) );
  XOR U7748 ( .A(p_input[432]), .B(n7917), .Z(n7919) );
  XNOR U7749 ( .A(n7920), .B(n7921), .Z(n7917) );
  AND U7750 ( .A(n336), .B(n7916), .Z(n7921) );
  XNOR U7751 ( .A(n7920), .B(n7914), .Z(n7916) );
  XOR U7752 ( .A(n7922), .B(n7923), .Z(n7914) );
  AND U7753 ( .A(n351), .B(n7924), .Z(n7923) );
  XNOR U7754 ( .A(n7925), .B(n7926), .Z(n7920) );
  AND U7755 ( .A(n343), .B(n7927), .Z(n7926) );
  XOR U7756 ( .A(p_input[448]), .B(n7925), .Z(n7927) );
  XNOR U7757 ( .A(n7928), .B(n7929), .Z(n7925) );
  AND U7758 ( .A(n347), .B(n7924), .Z(n7929) );
  XNOR U7759 ( .A(n7928), .B(n7922), .Z(n7924) );
  XOR U7760 ( .A(n7930), .B(n7931), .Z(n7922) );
  AND U7761 ( .A(n362), .B(n7932), .Z(n7931) );
  XNOR U7762 ( .A(n7933), .B(n7934), .Z(n7928) );
  AND U7763 ( .A(n354), .B(n7935), .Z(n7934) );
  XOR U7764 ( .A(p_input[464]), .B(n7933), .Z(n7935) );
  XNOR U7765 ( .A(n7936), .B(n7937), .Z(n7933) );
  AND U7766 ( .A(n358), .B(n7932), .Z(n7937) );
  XNOR U7767 ( .A(n7936), .B(n7930), .Z(n7932) );
  XOR U7768 ( .A(n7938), .B(n7939), .Z(n7930) );
  AND U7769 ( .A(n373), .B(n7940), .Z(n7939) );
  XNOR U7770 ( .A(n7941), .B(n7942), .Z(n7936) );
  AND U7771 ( .A(n365), .B(n7943), .Z(n7942) );
  XOR U7772 ( .A(p_input[480]), .B(n7941), .Z(n7943) );
  XNOR U7773 ( .A(n7944), .B(n7945), .Z(n7941) );
  AND U7774 ( .A(n369), .B(n7940), .Z(n7945) );
  XNOR U7775 ( .A(n7944), .B(n7938), .Z(n7940) );
  XOR U7776 ( .A(n7946), .B(n7947), .Z(n7938) );
  AND U7777 ( .A(n384), .B(n7948), .Z(n7947) );
  XNOR U7778 ( .A(n7949), .B(n7950), .Z(n7944) );
  AND U7779 ( .A(n376), .B(n7951), .Z(n7950) );
  XOR U7780 ( .A(p_input[496]), .B(n7949), .Z(n7951) );
  XNOR U7781 ( .A(n7952), .B(n7953), .Z(n7949) );
  AND U7782 ( .A(n380), .B(n7948), .Z(n7953) );
  XNOR U7783 ( .A(n7952), .B(n7946), .Z(n7948) );
  XOR U7784 ( .A(n7954), .B(n7955), .Z(n7946) );
  AND U7785 ( .A(n395), .B(n7956), .Z(n7955) );
  XNOR U7786 ( .A(n7957), .B(n7958), .Z(n7952) );
  AND U7787 ( .A(n387), .B(n7959), .Z(n7958) );
  XOR U7788 ( .A(p_input[512]), .B(n7957), .Z(n7959) );
  XNOR U7789 ( .A(n7960), .B(n7961), .Z(n7957) );
  AND U7790 ( .A(n391), .B(n7956), .Z(n7961) );
  XNOR U7791 ( .A(n7960), .B(n7954), .Z(n7956) );
  XOR U7792 ( .A(n7962), .B(n7963), .Z(n7954) );
  AND U7793 ( .A(n406), .B(n7964), .Z(n7963) );
  XNOR U7794 ( .A(n7965), .B(n7966), .Z(n7960) );
  AND U7795 ( .A(n398), .B(n7967), .Z(n7966) );
  XOR U7796 ( .A(p_input[528]), .B(n7965), .Z(n7967) );
  XNOR U7797 ( .A(n7968), .B(n7969), .Z(n7965) );
  AND U7798 ( .A(n402), .B(n7964), .Z(n7969) );
  XNOR U7799 ( .A(n7968), .B(n7962), .Z(n7964) );
  XOR U7800 ( .A(n7970), .B(n7971), .Z(n7962) );
  AND U7801 ( .A(n417), .B(n7972), .Z(n7971) );
  XNOR U7802 ( .A(n7973), .B(n7974), .Z(n7968) );
  AND U7803 ( .A(n409), .B(n7975), .Z(n7974) );
  XOR U7804 ( .A(p_input[544]), .B(n7973), .Z(n7975) );
  XNOR U7805 ( .A(n7976), .B(n7977), .Z(n7973) );
  AND U7806 ( .A(n413), .B(n7972), .Z(n7977) );
  XNOR U7807 ( .A(n7976), .B(n7970), .Z(n7972) );
  XOR U7808 ( .A(n7978), .B(n7979), .Z(n7970) );
  AND U7809 ( .A(n428), .B(n7980), .Z(n7979) );
  XNOR U7810 ( .A(n7981), .B(n7982), .Z(n7976) );
  AND U7811 ( .A(n420), .B(n7983), .Z(n7982) );
  XOR U7812 ( .A(p_input[560]), .B(n7981), .Z(n7983) );
  XNOR U7813 ( .A(n7984), .B(n7985), .Z(n7981) );
  AND U7814 ( .A(n424), .B(n7980), .Z(n7985) );
  XNOR U7815 ( .A(n7984), .B(n7978), .Z(n7980) );
  XOR U7816 ( .A(n7986), .B(n7987), .Z(n7978) );
  AND U7817 ( .A(n439), .B(n7988), .Z(n7987) );
  XNOR U7818 ( .A(n7989), .B(n7990), .Z(n7984) );
  AND U7819 ( .A(n431), .B(n7991), .Z(n7990) );
  XOR U7820 ( .A(p_input[576]), .B(n7989), .Z(n7991) );
  XNOR U7821 ( .A(n7992), .B(n7993), .Z(n7989) );
  AND U7822 ( .A(n435), .B(n7988), .Z(n7993) );
  XNOR U7823 ( .A(n7992), .B(n7986), .Z(n7988) );
  XOR U7824 ( .A(n7994), .B(n7995), .Z(n7986) );
  AND U7825 ( .A(n450), .B(n7996), .Z(n7995) );
  XNOR U7826 ( .A(n7997), .B(n7998), .Z(n7992) );
  AND U7827 ( .A(n442), .B(n7999), .Z(n7998) );
  XOR U7828 ( .A(p_input[592]), .B(n7997), .Z(n7999) );
  XNOR U7829 ( .A(n8000), .B(n8001), .Z(n7997) );
  AND U7830 ( .A(n446), .B(n7996), .Z(n8001) );
  XNOR U7831 ( .A(n8000), .B(n7994), .Z(n7996) );
  XOR U7832 ( .A(n8002), .B(n8003), .Z(n7994) );
  AND U7833 ( .A(n461), .B(n8004), .Z(n8003) );
  XNOR U7834 ( .A(n8005), .B(n8006), .Z(n8000) );
  AND U7835 ( .A(n453), .B(n8007), .Z(n8006) );
  XOR U7836 ( .A(p_input[608]), .B(n8005), .Z(n8007) );
  XNOR U7837 ( .A(n8008), .B(n8009), .Z(n8005) );
  AND U7838 ( .A(n457), .B(n8004), .Z(n8009) );
  XNOR U7839 ( .A(n8008), .B(n8002), .Z(n8004) );
  XOR U7840 ( .A(n8010), .B(n8011), .Z(n8002) );
  AND U7841 ( .A(n472), .B(n8012), .Z(n8011) );
  XNOR U7842 ( .A(n8013), .B(n8014), .Z(n8008) );
  AND U7843 ( .A(n464), .B(n8015), .Z(n8014) );
  XOR U7844 ( .A(p_input[624]), .B(n8013), .Z(n8015) );
  XNOR U7845 ( .A(n8016), .B(n8017), .Z(n8013) );
  AND U7846 ( .A(n468), .B(n8012), .Z(n8017) );
  XNOR U7847 ( .A(n8016), .B(n8010), .Z(n8012) );
  XOR U7848 ( .A(n8018), .B(n8019), .Z(n8010) );
  AND U7849 ( .A(n483), .B(n8020), .Z(n8019) );
  XNOR U7850 ( .A(n8021), .B(n8022), .Z(n8016) );
  AND U7851 ( .A(n475), .B(n8023), .Z(n8022) );
  XOR U7852 ( .A(p_input[640]), .B(n8021), .Z(n8023) );
  XNOR U7853 ( .A(n8024), .B(n8025), .Z(n8021) );
  AND U7854 ( .A(n479), .B(n8020), .Z(n8025) );
  XNOR U7855 ( .A(n8024), .B(n8018), .Z(n8020) );
  XOR U7856 ( .A(n8026), .B(n8027), .Z(n8018) );
  AND U7857 ( .A(n494), .B(n8028), .Z(n8027) );
  XNOR U7858 ( .A(n8029), .B(n8030), .Z(n8024) );
  AND U7859 ( .A(n486), .B(n8031), .Z(n8030) );
  XOR U7860 ( .A(p_input[656]), .B(n8029), .Z(n8031) );
  XNOR U7861 ( .A(n8032), .B(n8033), .Z(n8029) );
  AND U7862 ( .A(n490), .B(n8028), .Z(n8033) );
  XNOR U7863 ( .A(n8032), .B(n8026), .Z(n8028) );
  XOR U7864 ( .A(n8034), .B(n8035), .Z(n8026) );
  AND U7865 ( .A(n505), .B(n8036), .Z(n8035) );
  XNOR U7866 ( .A(n8037), .B(n8038), .Z(n8032) );
  AND U7867 ( .A(n497), .B(n8039), .Z(n8038) );
  XOR U7868 ( .A(p_input[672]), .B(n8037), .Z(n8039) );
  XNOR U7869 ( .A(n8040), .B(n8041), .Z(n8037) );
  AND U7870 ( .A(n501), .B(n8036), .Z(n8041) );
  XNOR U7871 ( .A(n8040), .B(n8034), .Z(n8036) );
  XOR U7872 ( .A(n8042), .B(n8043), .Z(n8034) );
  AND U7873 ( .A(n516), .B(n8044), .Z(n8043) );
  XNOR U7874 ( .A(n8045), .B(n8046), .Z(n8040) );
  AND U7875 ( .A(n508), .B(n8047), .Z(n8046) );
  XOR U7876 ( .A(p_input[688]), .B(n8045), .Z(n8047) );
  XNOR U7877 ( .A(n8048), .B(n8049), .Z(n8045) );
  AND U7878 ( .A(n512), .B(n8044), .Z(n8049) );
  XNOR U7879 ( .A(n8048), .B(n8042), .Z(n8044) );
  XOR U7880 ( .A(n8050), .B(n8051), .Z(n8042) );
  AND U7881 ( .A(n527), .B(n8052), .Z(n8051) );
  XNOR U7882 ( .A(n8053), .B(n8054), .Z(n8048) );
  AND U7883 ( .A(n519), .B(n8055), .Z(n8054) );
  XOR U7884 ( .A(p_input[704]), .B(n8053), .Z(n8055) );
  XNOR U7885 ( .A(n8056), .B(n8057), .Z(n8053) );
  AND U7886 ( .A(n523), .B(n8052), .Z(n8057) );
  XNOR U7887 ( .A(n8056), .B(n8050), .Z(n8052) );
  XOR U7888 ( .A(n8058), .B(n8059), .Z(n8050) );
  AND U7889 ( .A(n538), .B(n8060), .Z(n8059) );
  XNOR U7890 ( .A(n8061), .B(n8062), .Z(n8056) );
  AND U7891 ( .A(n530), .B(n8063), .Z(n8062) );
  XOR U7892 ( .A(p_input[720]), .B(n8061), .Z(n8063) );
  XNOR U7893 ( .A(n8064), .B(n8065), .Z(n8061) );
  AND U7894 ( .A(n534), .B(n8060), .Z(n8065) );
  XNOR U7895 ( .A(n8064), .B(n8058), .Z(n8060) );
  XOR U7896 ( .A(n8066), .B(n8067), .Z(n8058) );
  AND U7897 ( .A(n549), .B(n8068), .Z(n8067) );
  XNOR U7898 ( .A(n8069), .B(n8070), .Z(n8064) );
  AND U7899 ( .A(n541), .B(n8071), .Z(n8070) );
  XOR U7900 ( .A(p_input[736]), .B(n8069), .Z(n8071) );
  XNOR U7901 ( .A(n8072), .B(n8073), .Z(n8069) );
  AND U7902 ( .A(n545), .B(n8068), .Z(n8073) );
  XNOR U7903 ( .A(n8072), .B(n8066), .Z(n8068) );
  XOR U7904 ( .A(n8074), .B(n8075), .Z(n8066) );
  AND U7905 ( .A(n560), .B(n8076), .Z(n8075) );
  XNOR U7906 ( .A(n8077), .B(n8078), .Z(n8072) );
  AND U7907 ( .A(n552), .B(n8079), .Z(n8078) );
  XOR U7908 ( .A(p_input[752]), .B(n8077), .Z(n8079) );
  XNOR U7909 ( .A(n8080), .B(n8081), .Z(n8077) );
  AND U7910 ( .A(n556), .B(n8076), .Z(n8081) );
  XNOR U7911 ( .A(n8080), .B(n8074), .Z(n8076) );
  XOR U7912 ( .A(n8082), .B(n8083), .Z(n8074) );
  AND U7913 ( .A(n571), .B(n8084), .Z(n8083) );
  XNOR U7914 ( .A(n8085), .B(n8086), .Z(n8080) );
  AND U7915 ( .A(n563), .B(n8087), .Z(n8086) );
  XOR U7916 ( .A(p_input[768]), .B(n8085), .Z(n8087) );
  XNOR U7917 ( .A(n8088), .B(n8089), .Z(n8085) );
  AND U7918 ( .A(n567), .B(n8084), .Z(n8089) );
  XNOR U7919 ( .A(n8088), .B(n8082), .Z(n8084) );
  XOR U7920 ( .A(n8090), .B(n8091), .Z(n8082) );
  AND U7921 ( .A(n582), .B(n8092), .Z(n8091) );
  XNOR U7922 ( .A(n8093), .B(n8094), .Z(n8088) );
  AND U7923 ( .A(n574), .B(n8095), .Z(n8094) );
  XOR U7924 ( .A(p_input[784]), .B(n8093), .Z(n8095) );
  XNOR U7925 ( .A(n8096), .B(n8097), .Z(n8093) );
  AND U7926 ( .A(n578), .B(n8092), .Z(n8097) );
  XNOR U7927 ( .A(n8096), .B(n8090), .Z(n8092) );
  XOR U7928 ( .A(n8098), .B(n8099), .Z(n8090) );
  AND U7929 ( .A(n593), .B(n8100), .Z(n8099) );
  XNOR U7930 ( .A(n8101), .B(n8102), .Z(n8096) );
  AND U7931 ( .A(n585), .B(n8103), .Z(n8102) );
  XOR U7932 ( .A(p_input[800]), .B(n8101), .Z(n8103) );
  XNOR U7933 ( .A(n8104), .B(n8105), .Z(n8101) );
  AND U7934 ( .A(n589), .B(n8100), .Z(n8105) );
  XNOR U7935 ( .A(n8104), .B(n8098), .Z(n8100) );
  XOR U7936 ( .A(n8106), .B(n8107), .Z(n8098) );
  AND U7937 ( .A(n604), .B(n8108), .Z(n8107) );
  XNOR U7938 ( .A(n8109), .B(n8110), .Z(n8104) );
  AND U7939 ( .A(n596), .B(n8111), .Z(n8110) );
  XOR U7940 ( .A(p_input[816]), .B(n8109), .Z(n8111) );
  XNOR U7941 ( .A(n8112), .B(n8113), .Z(n8109) );
  AND U7942 ( .A(n600), .B(n8108), .Z(n8113) );
  XNOR U7943 ( .A(n8112), .B(n8106), .Z(n8108) );
  XOR U7944 ( .A(n8114), .B(n8115), .Z(n8106) );
  AND U7945 ( .A(n615), .B(n8116), .Z(n8115) );
  XNOR U7946 ( .A(n8117), .B(n8118), .Z(n8112) );
  AND U7947 ( .A(n607), .B(n8119), .Z(n8118) );
  XOR U7948 ( .A(p_input[832]), .B(n8117), .Z(n8119) );
  XNOR U7949 ( .A(n8120), .B(n8121), .Z(n8117) );
  AND U7950 ( .A(n611), .B(n8116), .Z(n8121) );
  XNOR U7951 ( .A(n8120), .B(n8114), .Z(n8116) );
  XOR U7952 ( .A(n8122), .B(n8123), .Z(n8114) );
  AND U7953 ( .A(n626), .B(n8124), .Z(n8123) );
  XNOR U7954 ( .A(n8125), .B(n8126), .Z(n8120) );
  AND U7955 ( .A(n618), .B(n8127), .Z(n8126) );
  XOR U7956 ( .A(p_input[848]), .B(n8125), .Z(n8127) );
  XNOR U7957 ( .A(n8128), .B(n8129), .Z(n8125) );
  AND U7958 ( .A(n622), .B(n8124), .Z(n8129) );
  XNOR U7959 ( .A(n8128), .B(n8122), .Z(n8124) );
  XOR U7960 ( .A(n8130), .B(n8131), .Z(n8122) );
  AND U7961 ( .A(n637), .B(n8132), .Z(n8131) );
  XNOR U7962 ( .A(n8133), .B(n8134), .Z(n8128) );
  AND U7963 ( .A(n629), .B(n8135), .Z(n8134) );
  XOR U7964 ( .A(p_input[864]), .B(n8133), .Z(n8135) );
  XNOR U7965 ( .A(n8136), .B(n8137), .Z(n8133) );
  AND U7966 ( .A(n633), .B(n8132), .Z(n8137) );
  XNOR U7967 ( .A(n8136), .B(n8130), .Z(n8132) );
  XOR U7968 ( .A(n8138), .B(n8139), .Z(n8130) );
  AND U7969 ( .A(n648), .B(n8140), .Z(n8139) );
  XNOR U7970 ( .A(n8141), .B(n8142), .Z(n8136) );
  AND U7971 ( .A(n640), .B(n8143), .Z(n8142) );
  XOR U7972 ( .A(p_input[880]), .B(n8141), .Z(n8143) );
  XNOR U7973 ( .A(n8144), .B(n8145), .Z(n8141) );
  AND U7974 ( .A(n644), .B(n8140), .Z(n8145) );
  XNOR U7975 ( .A(n8144), .B(n8138), .Z(n8140) );
  XOR U7976 ( .A(n8146), .B(n8147), .Z(n8138) );
  AND U7977 ( .A(n659), .B(n8148), .Z(n8147) );
  XNOR U7978 ( .A(n8149), .B(n8150), .Z(n8144) );
  AND U7979 ( .A(n651), .B(n8151), .Z(n8150) );
  XOR U7980 ( .A(p_input[896]), .B(n8149), .Z(n8151) );
  XNOR U7981 ( .A(n8152), .B(n8153), .Z(n8149) );
  AND U7982 ( .A(n655), .B(n8148), .Z(n8153) );
  XNOR U7983 ( .A(n8152), .B(n8146), .Z(n8148) );
  XOR U7984 ( .A(n8154), .B(n8155), .Z(n8146) );
  AND U7985 ( .A(n670), .B(n8156), .Z(n8155) );
  XNOR U7986 ( .A(n8157), .B(n8158), .Z(n8152) );
  AND U7987 ( .A(n662), .B(n8159), .Z(n8158) );
  XOR U7988 ( .A(p_input[912]), .B(n8157), .Z(n8159) );
  XNOR U7989 ( .A(n8160), .B(n8161), .Z(n8157) );
  AND U7990 ( .A(n666), .B(n8156), .Z(n8161) );
  XNOR U7991 ( .A(n8160), .B(n8154), .Z(n8156) );
  XOR U7992 ( .A(n8162), .B(n8163), .Z(n8154) );
  AND U7993 ( .A(n681), .B(n8164), .Z(n8163) );
  XNOR U7994 ( .A(n8165), .B(n8166), .Z(n8160) );
  AND U7995 ( .A(n673), .B(n8167), .Z(n8166) );
  XOR U7996 ( .A(p_input[928]), .B(n8165), .Z(n8167) );
  XNOR U7997 ( .A(n8168), .B(n8169), .Z(n8165) );
  AND U7998 ( .A(n677), .B(n8164), .Z(n8169) );
  XNOR U7999 ( .A(n8168), .B(n8162), .Z(n8164) );
  XOR U8000 ( .A(n8170), .B(n8171), .Z(n8162) );
  AND U8001 ( .A(n692), .B(n8172), .Z(n8171) );
  XNOR U8002 ( .A(n8173), .B(n8174), .Z(n8168) );
  AND U8003 ( .A(n684), .B(n8175), .Z(n8174) );
  XOR U8004 ( .A(p_input[944]), .B(n8173), .Z(n8175) );
  XNOR U8005 ( .A(n8176), .B(n8177), .Z(n8173) );
  AND U8006 ( .A(n688), .B(n8172), .Z(n8177) );
  XNOR U8007 ( .A(n8176), .B(n8170), .Z(n8172) );
  XOR U8008 ( .A(n8178), .B(n8179), .Z(n8170) );
  AND U8009 ( .A(n703), .B(n8180), .Z(n8179) );
  XNOR U8010 ( .A(n8181), .B(n8182), .Z(n8176) );
  AND U8011 ( .A(n695), .B(n8183), .Z(n8182) );
  XOR U8012 ( .A(p_input[960]), .B(n8181), .Z(n8183) );
  XNOR U8013 ( .A(n8184), .B(n8185), .Z(n8181) );
  AND U8014 ( .A(n699), .B(n8180), .Z(n8185) );
  XNOR U8015 ( .A(n8184), .B(n8178), .Z(n8180) );
  XOR U8016 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n8186), .Z(n8178) );
  AND U8017 ( .A(n713), .B(n8187), .Z(n8186) );
  XNOR U8018 ( .A(n8188), .B(n8189), .Z(n8184) );
  AND U8019 ( .A(n706), .B(n8190), .Z(n8189) );
  XOR U8020 ( .A(p_input[976]), .B(n8188), .Z(n8190) );
  XNOR U8021 ( .A(n8191), .B(n8192), .Z(n8188) );
  AND U8022 ( .A(n710), .B(n8187), .Z(n8192) );
  XOR U8023 ( .A(\knn_comb_/min_val_out[0][0] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n8187) );
  IV U8024 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n8191) );
  XNOR U8025 ( .A(n8193), .B(n8194), .Z(n30) );
  AND U8026 ( .A(n8195), .B(n8196), .Z(n8194) );
  XNOR U8027 ( .A(n8193), .B(n8197), .Z(n8196) );
  XOR U8028 ( .A(n8198), .B(n8199), .Z(n8197) );
  AND U8029 ( .A(n34), .B(n8200), .Z(n8199) );
  XNOR U8030 ( .A(n8198), .B(n8201), .Z(n8200) );
  XNOR U8031 ( .A(n8193), .B(n8202), .Z(n8195) );
  XOR U8032 ( .A(n8203), .B(n8204), .Z(n8202) );
  AND U8033 ( .A(n42), .B(n8205), .Z(n8204) );
  XOR U8034 ( .A(n8206), .B(n8207), .Z(n8193) );
  AND U8035 ( .A(n8208), .B(n8209), .Z(n8207) );
  XOR U8036 ( .A(n8210), .B(n8206), .Z(n8209) );
  XOR U8037 ( .A(n8211), .B(n8212), .Z(n8210) );
  AND U8038 ( .A(n34), .B(n8213), .Z(n8212) );
  XOR U8039 ( .A(n8214), .B(n8211), .Z(n8213) );
  XNOR U8040 ( .A(n8206), .B(n8215), .Z(n8208) );
  XOR U8041 ( .A(n8216), .B(n8217), .Z(n8215) );
  AND U8042 ( .A(n42), .B(n8218), .Z(n8217) );
  XOR U8043 ( .A(n8219), .B(n8220), .Z(n8206) );
  AND U8044 ( .A(n8221), .B(n8222), .Z(n8220) );
  XOR U8045 ( .A(n8223), .B(n8219), .Z(n8222) );
  XOR U8046 ( .A(n8224), .B(n8225), .Z(n8223) );
  AND U8047 ( .A(n34), .B(n8226), .Z(n8225) );
  XNOR U8048 ( .A(n8227), .B(n8224), .Z(n8226) );
  XNOR U8049 ( .A(n8219), .B(n8228), .Z(n8221) );
  XOR U8050 ( .A(n8229), .B(n8230), .Z(n8228) );
  AND U8051 ( .A(n42), .B(n8231), .Z(n8230) );
  XOR U8052 ( .A(n8232), .B(n8233), .Z(n8219) );
  AND U8053 ( .A(n8234), .B(n8235), .Z(n8233) );
  XOR U8054 ( .A(n8232), .B(n8236), .Z(n8235) );
  XOR U8055 ( .A(n8237), .B(n8238), .Z(n8236) );
  AND U8056 ( .A(n34), .B(n8239), .Z(n8238) );
  XOR U8057 ( .A(n8240), .B(n8237), .Z(n8239) );
  XNOR U8058 ( .A(n8241), .B(n8232), .Z(n8234) );
  XNOR U8059 ( .A(n8242), .B(n8243), .Z(n8241) );
  AND U8060 ( .A(n42), .B(n8244), .Z(n8243) );
  AND U8061 ( .A(n8245), .B(n8246), .Z(n8232) );
  XNOR U8062 ( .A(n8247), .B(n8248), .Z(n8246) );
  AND U8063 ( .A(n34), .B(n8249), .Z(n8248) );
  XNOR U8064 ( .A(n8250), .B(n8247), .Z(n8249) );
  XNOR U8065 ( .A(n8251), .B(n8252), .Z(n34) );
  AND U8066 ( .A(n8253), .B(n8254), .Z(n8252) );
  XOR U8067 ( .A(n8201), .B(n8251), .Z(n8254) );
  AND U8068 ( .A(n8255), .B(n8256), .Z(n8201) );
  XOR U8069 ( .A(n8251), .B(n8198), .Z(n8253) );
  XNOR U8070 ( .A(n8257), .B(n8258), .Z(n8198) );
  AND U8071 ( .A(n38), .B(n8205), .Z(n8258) );
  XOR U8072 ( .A(n8203), .B(n8257), .Z(n8205) );
  XOR U8073 ( .A(n8259), .B(n8260), .Z(n8251) );
  AND U8074 ( .A(n8261), .B(n8262), .Z(n8260) );
  XNOR U8075 ( .A(n8259), .B(n8255), .Z(n8262) );
  IV U8076 ( .A(n8214), .Z(n8255) );
  XOR U8077 ( .A(n8263), .B(n8264), .Z(n8214) );
  XOR U8078 ( .A(n8265), .B(n8256), .Z(n8264) );
  AND U8079 ( .A(n8227), .B(n8266), .Z(n8256) );
  AND U8080 ( .A(n8267), .B(n8268), .Z(n8265) );
  XOR U8081 ( .A(n8269), .B(n8263), .Z(n8267) );
  XNOR U8082 ( .A(n8211), .B(n8259), .Z(n8261) );
  XNOR U8083 ( .A(n8270), .B(n8271), .Z(n8211) );
  AND U8084 ( .A(n38), .B(n8218), .Z(n8271) );
  XOR U8085 ( .A(n8270), .B(n8272), .Z(n8218) );
  XOR U8086 ( .A(n8273), .B(n8274), .Z(n8259) );
  AND U8087 ( .A(n8275), .B(n8276), .Z(n8274) );
  XNOR U8088 ( .A(n8273), .B(n8227), .Z(n8276) );
  XOR U8089 ( .A(n8277), .B(n8268), .Z(n8227) );
  XNOR U8090 ( .A(n8278), .B(n8263), .Z(n8268) );
  XOR U8091 ( .A(n8279), .B(n8280), .Z(n8263) );
  AND U8092 ( .A(n8281), .B(n8282), .Z(n8280) );
  XOR U8093 ( .A(n8283), .B(n8279), .Z(n8281) );
  XNOR U8094 ( .A(n8284), .B(n8285), .Z(n8278) );
  AND U8095 ( .A(n8286), .B(n8287), .Z(n8285) );
  XOR U8096 ( .A(n8284), .B(n8288), .Z(n8286) );
  XNOR U8097 ( .A(n8269), .B(n8266), .Z(n8277) );
  AND U8098 ( .A(n8289), .B(n8290), .Z(n8266) );
  XOR U8099 ( .A(n8291), .B(n8292), .Z(n8269) );
  AND U8100 ( .A(n8293), .B(n8294), .Z(n8292) );
  XOR U8101 ( .A(n8291), .B(n8295), .Z(n8293) );
  XNOR U8102 ( .A(n8224), .B(n8273), .Z(n8275) );
  XNOR U8103 ( .A(n8296), .B(n8297), .Z(n8224) );
  AND U8104 ( .A(n38), .B(n8231), .Z(n8297) );
  XOR U8105 ( .A(n8296), .B(n8298), .Z(n8231) );
  XOR U8106 ( .A(n8299), .B(n8300), .Z(n8273) );
  AND U8107 ( .A(n8301), .B(n8302), .Z(n8300) );
  XNOR U8108 ( .A(n8299), .B(n8289), .Z(n8302) );
  IV U8109 ( .A(n8240), .Z(n8289) );
  XNOR U8110 ( .A(n8303), .B(n8282), .Z(n8240) );
  XNOR U8111 ( .A(n8304), .B(n8288), .Z(n8282) );
  XOR U8112 ( .A(n8305), .B(n8306), .Z(n8288) );
  NOR U8113 ( .A(n8307), .B(n8308), .Z(n8306) );
  XNOR U8114 ( .A(n8305), .B(n8309), .Z(n8307) );
  XNOR U8115 ( .A(n8287), .B(n8279), .Z(n8304) );
  XOR U8116 ( .A(n8310), .B(n8311), .Z(n8279) );
  AND U8117 ( .A(n8312), .B(n8313), .Z(n8311) );
  XNOR U8118 ( .A(n8310), .B(n8314), .Z(n8312) );
  XNOR U8119 ( .A(n8315), .B(n8284), .Z(n8287) );
  XOR U8120 ( .A(n8316), .B(n8317), .Z(n8284) );
  AND U8121 ( .A(n8318), .B(n8319), .Z(n8317) );
  XOR U8122 ( .A(n8316), .B(n8320), .Z(n8318) );
  XNOR U8123 ( .A(n8321), .B(n8322), .Z(n8315) );
  NOR U8124 ( .A(n8323), .B(n8324), .Z(n8322) );
  XOR U8125 ( .A(n8321), .B(n8325), .Z(n8323) );
  XNOR U8126 ( .A(n8283), .B(n8290), .Z(n8303) );
  NOR U8127 ( .A(n8250), .B(n8326), .Z(n8290) );
  XOR U8128 ( .A(n8295), .B(n8294), .Z(n8283) );
  XNOR U8129 ( .A(n8327), .B(n8291), .Z(n8294) );
  XOR U8130 ( .A(n8328), .B(n8329), .Z(n8291) );
  AND U8131 ( .A(n8330), .B(n8331), .Z(n8329) );
  XOR U8132 ( .A(n8328), .B(n8332), .Z(n8330) );
  XNOR U8133 ( .A(n8333), .B(n8334), .Z(n8327) );
  NOR U8134 ( .A(n8335), .B(n8336), .Z(n8334) );
  XNOR U8135 ( .A(n8333), .B(n8337), .Z(n8335) );
  XOR U8136 ( .A(n8338), .B(n8339), .Z(n8295) );
  NOR U8137 ( .A(n8340), .B(n8341), .Z(n8339) );
  XNOR U8138 ( .A(n8338), .B(n8342), .Z(n8340) );
  XNOR U8139 ( .A(n8237), .B(n8299), .Z(n8301) );
  XNOR U8140 ( .A(n8343), .B(n8344), .Z(n8237) );
  AND U8141 ( .A(n38), .B(n8244), .Z(n8344) );
  XOR U8142 ( .A(n8343), .B(n8242), .Z(n8244) );
  AND U8143 ( .A(n8247), .B(n8250), .Z(n8299) );
  XOR U8144 ( .A(n8345), .B(n8326), .Z(n8250) );
  XNOR U8145 ( .A(p_input[0]), .B(p_input[1024]), .Z(n8326) );
  XOR U8146 ( .A(n8314), .B(n8313), .Z(n8345) );
  XNOR U8147 ( .A(n8346), .B(n8320), .Z(n8313) );
  XNOR U8148 ( .A(n8309), .B(n8308), .Z(n8320) );
  XOR U8149 ( .A(n8347), .B(n8305), .Z(n8308) );
  XOR U8150 ( .A(p_input[1034]), .B(p_input[10]), .Z(n8305) );
  XNOR U8151 ( .A(p_input[1035]), .B(p_input[11]), .Z(n8347) );
  XOR U8152 ( .A(p_input[1036]), .B(p_input[12]), .Z(n8309) );
  XNOR U8153 ( .A(n8319), .B(n8310), .Z(n8346) );
  XOR U8154 ( .A(p_input[1025]), .B(p_input[1]), .Z(n8310) );
  XOR U8155 ( .A(n8348), .B(n8325), .Z(n8319) );
  XNOR U8156 ( .A(p_input[1039]), .B(p_input[15]), .Z(n8325) );
  XOR U8157 ( .A(n8316), .B(n8324), .Z(n8348) );
  XOR U8158 ( .A(n8349), .B(n8321), .Z(n8324) );
  XOR U8159 ( .A(p_input[1037]), .B(p_input[13]), .Z(n8321) );
  XNOR U8160 ( .A(p_input[1038]), .B(p_input[14]), .Z(n8349) );
  XOR U8161 ( .A(p_input[1033]), .B(p_input[9]), .Z(n8316) );
  XNOR U8162 ( .A(n8332), .B(n8331), .Z(n8314) );
  XNOR U8163 ( .A(n8350), .B(n8337), .Z(n8331) );
  XOR U8164 ( .A(p_input[1032]), .B(p_input[8]), .Z(n8337) );
  XOR U8165 ( .A(n8328), .B(n8336), .Z(n8350) );
  XOR U8166 ( .A(n8351), .B(n8333), .Z(n8336) );
  XOR U8167 ( .A(p_input[1030]), .B(p_input[6]), .Z(n8333) );
  XNOR U8168 ( .A(p_input[1031]), .B(p_input[7]), .Z(n8351) );
  XOR U8169 ( .A(p_input[1026]), .B(p_input[2]), .Z(n8328) );
  XNOR U8170 ( .A(n8342), .B(n8341), .Z(n8332) );
  XOR U8171 ( .A(n8352), .B(n8338), .Z(n8341) );
  XOR U8172 ( .A(p_input[1027]), .B(p_input[3]), .Z(n8338) );
  XNOR U8173 ( .A(p_input[1028]), .B(p_input[4]), .Z(n8352) );
  XOR U8174 ( .A(p_input[1029]), .B(p_input[5]), .Z(n8342) );
  XNOR U8175 ( .A(n8353), .B(n8354), .Z(n8247) );
  AND U8176 ( .A(n38), .B(n8355), .Z(n8354) );
  XNOR U8177 ( .A(n8356), .B(n8357), .Z(n38) );
  AND U8178 ( .A(n8358), .B(n8359), .Z(n8357) );
  XOR U8179 ( .A(n8356), .B(n8257), .Z(n8359) );
  XNOR U8180 ( .A(n8356), .B(n8203), .Z(n8358) );
  XOR U8181 ( .A(n8360), .B(n8361), .Z(n8356) );
  AND U8182 ( .A(n8362), .B(n8363), .Z(n8361) );
  XNOR U8183 ( .A(n8270), .B(n8360), .Z(n8363) );
  XOR U8184 ( .A(n8360), .B(n8272), .Z(n8362) );
  XOR U8185 ( .A(n8364), .B(n8365), .Z(n8360) );
  AND U8186 ( .A(n8366), .B(n8367), .Z(n8365) );
  XOR U8187 ( .A(n8364), .B(n8298), .Z(n8366) );
  IV U8188 ( .A(n8229), .Z(n8298) );
  XOR U8189 ( .A(n8368), .B(n8369), .Z(n8245) );
  AND U8190 ( .A(n42), .B(n8355), .Z(n8369) );
  XNOR U8191 ( .A(n8353), .B(n8368), .Z(n8355) );
  XNOR U8192 ( .A(n8370), .B(n8371), .Z(n42) );
  AND U8193 ( .A(n8372), .B(n8373), .Z(n8371) );
  XNOR U8194 ( .A(n8374), .B(n8370), .Z(n8373) );
  IV U8195 ( .A(n8257), .Z(n8374) );
  XNOR U8196 ( .A(n8375), .B(n8376), .Z(n8257) );
  AND U8197 ( .A(n46), .B(n8377), .Z(n8376) );
  XNOR U8198 ( .A(n8375), .B(n8378), .Z(n8377) );
  XNOR U8199 ( .A(n8203), .B(n8370), .Z(n8372) );
  XOR U8200 ( .A(n8379), .B(n8380), .Z(n8203) );
  AND U8201 ( .A(n54), .B(n8381), .Z(n8380) );
  XOR U8202 ( .A(n8382), .B(n8383), .Z(n8370) );
  AND U8203 ( .A(n8384), .B(n8385), .Z(n8383) );
  XNOR U8204 ( .A(n8382), .B(n8270), .Z(n8385) );
  XNOR U8205 ( .A(n8386), .B(n8387), .Z(n8270) );
  AND U8206 ( .A(n46), .B(n8388), .Z(n8387) );
  XOR U8207 ( .A(n8389), .B(n8386), .Z(n8388) );
  XNOR U8208 ( .A(n8216), .B(n8382), .Z(n8384) );
  IV U8209 ( .A(n8272), .Z(n8216) );
  XOR U8210 ( .A(n8390), .B(n8391), .Z(n8272) );
  AND U8211 ( .A(n54), .B(n8392), .Z(n8391) );
  XOR U8212 ( .A(n8364), .B(n8393), .Z(n8382) );
  AND U8213 ( .A(n8394), .B(n8367), .Z(n8393) );
  XNOR U8214 ( .A(n8296), .B(n8364), .Z(n8367) );
  XNOR U8215 ( .A(n8395), .B(n8396), .Z(n8296) );
  AND U8216 ( .A(n46), .B(n8397), .Z(n8396) );
  XNOR U8217 ( .A(n8398), .B(n8395), .Z(n8397) );
  XNOR U8218 ( .A(n8229), .B(n8364), .Z(n8394) );
  XNOR U8219 ( .A(n8399), .B(n8400), .Z(n8229) );
  AND U8220 ( .A(n54), .B(n8401), .Z(n8400) );
  XOR U8221 ( .A(n8402), .B(n8403), .Z(n8364) );
  AND U8222 ( .A(n8404), .B(n8405), .Z(n8403) );
  XNOR U8223 ( .A(n8402), .B(n8343), .Z(n8405) );
  XNOR U8224 ( .A(n8406), .B(n8407), .Z(n8343) );
  AND U8225 ( .A(n46), .B(n8408), .Z(n8407) );
  XOR U8226 ( .A(n8409), .B(n8406), .Z(n8408) );
  XNOR U8227 ( .A(n8410), .B(n8402), .Z(n8404) );
  IV U8228 ( .A(n8242), .Z(n8410) );
  XOR U8229 ( .A(n8411), .B(n8412), .Z(n8242) );
  AND U8230 ( .A(n54), .B(n8413), .Z(n8412) );
  AND U8231 ( .A(n8368), .B(n8353), .Z(n8402) );
  XNOR U8232 ( .A(n8414), .B(n8415), .Z(n8353) );
  AND U8233 ( .A(n46), .B(n8416), .Z(n8415) );
  XNOR U8234 ( .A(n8417), .B(n8414), .Z(n8416) );
  XNOR U8235 ( .A(n8418), .B(n8419), .Z(n46) );
  AND U8236 ( .A(n8420), .B(n8421), .Z(n8419) );
  XOR U8237 ( .A(n8378), .B(n8418), .Z(n8421) );
  AND U8238 ( .A(n8422), .B(n8423), .Z(n8378) );
  XOR U8239 ( .A(n8418), .B(n8375), .Z(n8420) );
  XNOR U8240 ( .A(n8424), .B(n8425), .Z(n8375) );
  AND U8241 ( .A(n50), .B(n8381), .Z(n8425) );
  XOR U8242 ( .A(n8379), .B(n8424), .Z(n8381) );
  XOR U8243 ( .A(n8426), .B(n8427), .Z(n8418) );
  AND U8244 ( .A(n8428), .B(n8429), .Z(n8427) );
  XNOR U8245 ( .A(n8426), .B(n8422), .Z(n8429) );
  IV U8246 ( .A(n8389), .Z(n8422) );
  XOR U8247 ( .A(n8430), .B(n8431), .Z(n8389) );
  XOR U8248 ( .A(n8432), .B(n8423), .Z(n8431) );
  AND U8249 ( .A(n8398), .B(n8433), .Z(n8423) );
  AND U8250 ( .A(n8434), .B(n8435), .Z(n8432) );
  XOR U8251 ( .A(n8436), .B(n8430), .Z(n8434) );
  XNOR U8252 ( .A(n8386), .B(n8426), .Z(n8428) );
  XNOR U8253 ( .A(n8437), .B(n8438), .Z(n8386) );
  AND U8254 ( .A(n50), .B(n8392), .Z(n8438) );
  XOR U8255 ( .A(n8437), .B(n8390), .Z(n8392) );
  XOR U8256 ( .A(n8439), .B(n8440), .Z(n8426) );
  AND U8257 ( .A(n8441), .B(n8442), .Z(n8440) );
  XNOR U8258 ( .A(n8439), .B(n8398), .Z(n8442) );
  XOR U8259 ( .A(n8443), .B(n8435), .Z(n8398) );
  XNOR U8260 ( .A(n8444), .B(n8430), .Z(n8435) );
  XOR U8261 ( .A(n8445), .B(n8446), .Z(n8430) );
  AND U8262 ( .A(n8447), .B(n8448), .Z(n8446) );
  XOR U8263 ( .A(n8449), .B(n8445), .Z(n8447) );
  XNOR U8264 ( .A(n8450), .B(n8451), .Z(n8444) );
  AND U8265 ( .A(n8452), .B(n8453), .Z(n8451) );
  XOR U8266 ( .A(n8450), .B(n8454), .Z(n8452) );
  XNOR U8267 ( .A(n8436), .B(n8433), .Z(n8443) );
  AND U8268 ( .A(n8455), .B(n8456), .Z(n8433) );
  XOR U8269 ( .A(n8457), .B(n8458), .Z(n8436) );
  AND U8270 ( .A(n8459), .B(n8460), .Z(n8458) );
  XOR U8271 ( .A(n8457), .B(n8461), .Z(n8459) );
  XNOR U8272 ( .A(n8395), .B(n8439), .Z(n8441) );
  XNOR U8273 ( .A(n8462), .B(n8463), .Z(n8395) );
  AND U8274 ( .A(n50), .B(n8401), .Z(n8463) );
  XOR U8275 ( .A(n8462), .B(n8399), .Z(n8401) );
  XOR U8276 ( .A(n8464), .B(n8465), .Z(n8439) );
  AND U8277 ( .A(n8466), .B(n8467), .Z(n8465) );
  XNOR U8278 ( .A(n8464), .B(n8455), .Z(n8467) );
  IV U8279 ( .A(n8409), .Z(n8455) );
  XNOR U8280 ( .A(n8468), .B(n8448), .Z(n8409) );
  XNOR U8281 ( .A(n8469), .B(n8454), .Z(n8448) );
  XOR U8282 ( .A(n8470), .B(n8471), .Z(n8454) );
  NOR U8283 ( .A(n8472), .B(n8473), .Z(n8471) );
  XNOR U8284 ( .A(n8470), .B(n8474), .Z(n8472) );
  XNOR U8285 ( .A(n8453), .B(n8445), .Z(n8469) );
  XOR U8286 ( .A(n8475), .B(n8476), .Z(n8445) );
  AND U8287 ( .A(n8477), .B(n8478), .Z(n8476) );
  XNOR U8288 ( .A(n8475), .B(n8479), .Z(n8477) );
  XNOR U8289 ( .A(n8480), .B(n8450), .Z(n8453) );
  XOR U8290 ( .A(n8481), .B(n8482), .Z(n8450) );
  AND U8291 ( .A(n8483), .B(n8484), .Z(n8482) );
  XOR U8292 ( .A(n8481), .B(n8485), .Z(n8483) );
  XNOR U8293 ( .A(n8486), .B(n8487), .Z(n8480) );
  NOR U8294 ( .A(n8488), .B(n8489), .Z(n8487) );
  XOR U8295 ( .A(n8486), .B(n8490), .Z(n8488) );
  XNOR U8296 ( .A(n8449), .B(n8456), .Z(n8468) );
  NOR U8297 ( .A(n8417), .B(n8491), .Z(n8456) );
  XOR U8298 ( .A(n8461), .B(n8460), .Z(n8449) );
  XNOR U8299 ( .A(n8492), .B(n8457), .Z(n8460) );
  XOR U8300 ( .A(n8493), .B(n8494), .Z(n8457) );
  AND U8301 ( .A(n8495), .B(n8496), .Z(n8494) );
  XOR U8302 ( .A(n8493), .B(n8497), .Z(n8495) );
  XNOR U8303 ( .A(n8498), .B(n8499), .Z(n8492) );
  NOR U8304 ( .A(n8500), .B(n8501), .Z(n8499) );
  XNOR U8305 ( .A(n8498), .B(n8502), .Z(n8500) );
  XOR U8306 ( .A(n8503), .B(n8504), .Z(n8461) );
  NOR U8307 ( .A(n8505), .B(n8506), .Z(n8504) );
  XNOR U8308 ( .A(n8503), .B(n8507), .Z(n8505) );
  XNOR U8309 ( .A(n8406), .B(n8464), .Z(n8466) );
  XNOR U8310 ( .A(n8508), .B(n8509), .Z(n8406) );
  AND U8311 ( .A(n50), .B(n8413), .Z(n8509) );
  XOR U8312 ( .A(n8508), .B(n8411), .Z(n8413) );
  AND U8313 ( .A(n8414), .B(n8417), .Z(n8464) );
  XOR U8314 ( .A(n8510), .B(n8491), .Z(n8417) );
  XNOR U8315 ( .A(p_input[1024]), .B(p_input[16]), .Z(n8491) );
  XOR U8316 ( .A(n8479), .B(n8478), .Z(n8510) );
  XNOR U8317 ( .A(n8511), .B(n8485), .Z(n8478) );
  XNOR U8318 ( .A(n8474), .B(n8473), .Z(n8485) );
  XOR U8319 ( .A(n8512), .B(n8470), .Z(n8473) );
  XOR U8320 ( .A(p_input[1034]), .B(p_input[26]), .Z(n8470) );
  XNOR U8321 ( .A(p_input[1035]), .B(p_input[27]), .Z(n8512) );
  XOR U8322 ( .A(p_input[1036]), .B(p_input[28]), .Z(n8474) );
  XNOR U8323 ( .A(n8484), .B(n8475), .Z(n8511) );
  XOR U8324 ( .A(p_input[1025]), .B(p_input[17]), .Z(n8475) );
  XOR U8325 ( .A(n8513), .B(n8490), .Z(n8484) );
  XNOR U8326 ( .A(p_input[1039]), .B(p_input[31]), .Z(n8490) );
  XOR U8327 ( .A(n8481), .B(n8489), .Z(n8513) );
  XOR U8328 ( .A(n8514), .B(n8486), .Z(n8489) );
  XOR U8329 ( .A(p_input[1037]), .B(p_input[29]), .Z(n8486) );
  XNOR U8330 ( .A(p_input[1038]), .B(p_input[30]), .Z(n8514) );
  XOR U8331 ( .A(p_input[1033]), .B(p_input[25]), .Z(n8481) );
  XNOR U8332 ( .A(n8497), .B(n8496), .Z(n8479) );
  XNOR U8333 ( .A(n8515), .B(n8502), .Z(n8496) );
  XOR U8334 ( .A(p_input[1032]), .B(p_input[24]), .Z(n8502) );
  XOR U8335 ( .A(n8493), .B(n8501), .Z(n8515) );
  XOR U8336 ( .A(n8516), .B(n8498), .Z(n8501) );
  XOR U8337 ( .A(p_input[1030]), .B(p_input[22]), .Z(n8498) );
  XNOR U8338 ( .A(p_input[1031]), .B(p_input[23]), .Z(n8516) );
  XOR U8339 ( .A(p_input[1026]), .B(p_input[18]), .Z(n8493) );
  XNOR U8340 ( .A(n8507), .B(n8506), .Z(n8497) );
  XOR U8341 ( .A(n8517), .B(n8503), .Z(n8506) );
  XOR U8342 ( .A(p_input[1027]), .B(p_input[19]), .Z(n8503) );
  XNOR U8343 ( .A(p_input[1028]), .B(p_input[20]), .Z(n8517) );
  XOR U8344 ( .A(p_input[1029]), .B(p_input[21]), .Z(n8507) );
  XNOR U8345 ( .A(n8518), .B(n8519), .Z(n8414) );
  AND U8346 ( .A(n50), .B(n8520), .Z(n8519) );
  XNOR U8347 ( .A(n8521), .B(n8522), .Z(n50) );
  AND U8348 ( .A(n8523), .B(n8524), .Z(n8522) );
  XOR U8349 ( .A(n8521), .B(n8424), .Z(n8524) );
  XNOR U8350 ( .A(n8521), .B(n8379), .Z(n8523) );
  XOR U8351 ( .A(n8525), .B(n8526), .Z(n8521) );
  AND U8352 ( .A(n8527), .B(n8528), .Z(n8526) );
  XOR U8353 ( .A(n8525), .B(n8390), .Z(n8527) );
  XOR U8354 ( .A(n8529), .B(n8530), .Z(n8368) );
  AND U8355 ( .A(n54), .B(n8520), .Z(n8530) );
  XNOR U8356 ( .A(n8518), .B(n8529), .Z(n8520) );
  XNOR U8357 ( .A(n8531), .B(n8532), .Z(n54) );
  AND U8358 ( .A(n8533), .B(n8534), .Z(n8532) );
  XNOR U8359 ( .A(n8535), .B(n8531), .Z(n8534) );
  IV U8360 ( .A(n8424), .Z(n8535) );
  XNOR U8361 ( .A(n8536), .B(n8537), .Z(n8424) );
  AND U8362 ( .A(n57), .B(n8538), .Z(n8537) );
  XNOR U8363 ( .A(n8536), .B(n8539), .Z(n8538) );
  XNOR U8364 ( .A(n8379), .B(n8531), .Z(n8533) );
  XOR U8365 ( .A(n8540), .B(n8541), .Z(n8379) );
  AND U8366 ( .A(n65), .B(n8542), .Z(n8541) );
  XOR U8367 ( .A(n8525), .B(n8543), .Z(n8531) );
  AND U8368 ( .A(n8544), .B(n8528), .Z(n8543) );
  XNOR U8369 ( .A(n8437), .B(n8525), .Z(n8528) );
  XNOR U8370 ( .A(n8545), .B(n8546), .Z(n8437) );
  AND U8371 ( .A(n57), .B(n8547), .Z(n8546) );
  XOR U8372 ( .A(n8548), .B(n8545), .Z(n8547) );
  XNOR U8373 ( .A(n8549), .B(n8525), .Z(n8544) );
  IV U8374 ( .A(n8390), .Z(n8549) );
  XOR U8375 ( .A(n8550), .B(n8551), .Z(n8390) );
  AND U8376 ( .A(n65), .B(n8552), .Z(n8551) );
  XOR U8377 ( .A(n8553), .B(n8554), .Z(n8525) );
  AND U8378 ( .A(n8555), .B(n8556), .Z(n8554) );
  XNOR U8379 ( .A(n8462), .B(n8553), .Z(n8556) );
  XNOR U8380 ( .A(n8557), .B(n8558), .Z(n8462) );
  AND U8381 ( .A(n57), .B(n8559), .Z(n8558) );
  XNOR U8382 ( .A(n8560), .B(n8557), .Z(n8559) );
  XOR U8383 ( .A(n8553), .B(n8399), .Z(n8555) );
  XOR U8384 ( .A(n8561), .B(n8562), .Z(n8399) );
  AND U8385 ( .A(n65), .B(n8563), .Z(n8562) );
  XOR U8386 ( .A(n8564), .B(n8565), .Z(n8553) );
  AND U8387 ( .A(n8566), .B(n8567), .Z(n8565) );
  XNOR U8388 ( .A(n8564), .B(n8508), .Z(n8567) );
  XNOR U8389 ( .A(n8568), .B(n8569), .Z(n8508) );
  AND U8390 ( .A(n57), .B(n8570), .Z(n8569) );
  XOR U8391 ( .A(n8571), .B(n8568), .Z(n8570) );
  XNOR U8392 ( .A(n8572), .B(n8564), .Z(n8566) );
  IV U8393 ( .A(n8411), .Z(n8572) );
  XOR U8394 ( .A(n8573), .B(n8574), .Z(n8411) );
  AND U8395 ( .A(n65), .B(n8575), .Z(n8574) );
  AND U8396 ( .A(n8529), .B(n8518), .Z(n8564) );
  XNOR U8397 ( .A(n8576), .B(n8577), .Z(n8518) );
  AND U8398 ( .A(n57), .B(n8578), .Z(n8577) );
  XNOR U8399 ( .A(n8579), .B(n8576), .Z(n8578) );
  XNOR U8400 ( .A(n8580), .B(n8581), .Z(n57) );
  AND U8401 ( .A(n8582), .B(n8583), .Z(n8581) );
  XOR U8402 ( .A(n8539), .B(n8580), .Z(n8583) );
  AND U8403 ( .A(n8584), .B(n8585), .Z(n8539) );
  XOR U8404 ( .A(n8580), .B(n8536), .Z(n8582) );
  XNOR U8405 ( .A(n8586), .B(n8587), .Z(n8536) );
  AND U8406 ( .A(n61), .B(n8542), .Z(n8587) );
  XOR U8407 ( .A(n8540), .B(n8586), .Z(n8542) );
  XOR U8408 ( .A(n8588), .B(n8589), .Z(n8580) );
  AND U8409 ( .A(n8590), .B(n8591), .Z(n8589) );
  XNOR U8410 ( .A(n8588), .B(n8584), .Z(n8591) );
  IV U8411 ( .A(n8548), .Z(n8584) );
  XOR U8412 ( .A(n8592), .B(n8593), .Z(n8548) );
  XOR U8413 ( .A(n8594), .B(n8585), .Z(n8593) );
  AND U8414 ( .A(n8560), .B(n8595), .Z(n8585) );
  AND U8415 ( .A(n8596), .B(n8597), .Z(n8594) );
  XOR U8416 ( .A(n8598), .B(n8592), .Z(n8596) );
  XNOR U8417 ( .A(n8545), .B(n8588), .Z(n8590) );
  XNOR U8418 ( .A(n8599), .B(n8600), .Z(n8545) );
  AND U8419 ( .A(n61), .B(n8552), .Z(n8600) );
  XOR U8420 ( .A(n8599), .B(n8550), .Z(n8552) );
  XOR U8421 ( .A(n8601), .B(n8602), .Z(n8588) );
  AND U8422 ( .A(n8603), .B(n8604), .Z(n8602) );
  XNOR U8423 ( .A(n8601), .B(n8560), .Z(n8604) );
  XOR U8424 ( .A(n8605), .B(n8597), .Z(n8560) );
  XNOR U8425 ( .A(n8606), .B(n8592), .Z(n8597) );
  XOR U8426 ( .A(n8607), .B(n8608), .Z(n8592) );
  AND U8427 ( .A(n8609), .B(n8610), .Z(n8608) );
  XOR U8428 ( .A(n8611), .B(n8607), .Z(n8609) );
  XNOR U8429 ( .A(n8612), .B(n8613), .Z(n8606) );
  AND U8430 ( .A(n8614), .B(n8615), .Z(n8613) );
  XOR U8431 ( .A(n8612), .B(n8616), .Z(n8614) );
  XNOR U8432 ( .A(n8598), .B(n8595), .Z(n8605) );
  AND U8433 ( .A(n8617), .B(n8618), .Z(n8595) );
  XOR U8434 ( .A(n8619), .B(n8620), .Z(n8598) );
  AND U8435 ( .A(n8621), .B(n8622), .Z(n8620) );
  XOR U8436 ( .A(n8619), .B(n8623), .Z(n8621) );
  XNOR U8437 ( .A(n8557), .B(n8601), .Z(n8603) );
  XNOR U8438 ( .A(n8624), .B(n8625), .Z(n8557) );
  AND U8439 ( .A(n61), .B(n8563), .Z(n8625) );
  XOR U8440 ( .A(n8624), .B(n8561), .Z(n8563) );
  XOR U8441 ( .A(n8626), .B(n8627), .Z(n8601) );
  AND U8442 ( .A(n8628), .B(n8629), .Z(n8627) );
  XNOR U8443 ( .A(n8626), .B(n8617), .Z(n8629) );
  IV U8444 ( .A(n8571), .Z(n8617) );
  XNOR U8445 ( .A(n8630), .B(n8610), .Z(n8571) );
  XNOR U8446 ( .A(n8631), .B(n8616), .Z(n8610) );
  XOR U8447 ( .A(n8632), .B(n8633), .Z(n8616) );
  NOR U8448 ( .A(n8634), .B(n8635), .Z(n8633) );
  XNOR U8449 ( .A(n8632), .B(n8636), .Z(n8634) );
  XNOR U8450 ( .A(n8615), .B(n8607), .Z(n8631) );
  XOR U8451 ( .A(n8637), .B(n8638), .Z(n8607) );
  AND U8452 ( .A(n8639), .B(n8640), .Z(n8638) );
  XNOR U8453 ( .A(n8637), .B(n8641), .Z(n8639) );
  XNOR U8454 ( .A(n8642), .B(n8612), .Z(n8615) );
  XOR U8455 ( .A(n8643), .B(n8644), .Z(n8612) );
  AND U8456 ( .A(n8645), .B(n8646), .Z(n8644) );
  XOR U8457 ( .A(n8643), .B(n8647), .Z(n8645) );
  XNOR U8458 ( .A(n8648), .B(n8649), .Z(n8642) );
  NOR U8459 ( .A(n8650), .B(n8651), .Z(n8649) );
  XOR U8460 ( .A(n8648), .B(n8652), .Z(n8650) );
  XNOR U8461 ( .A(n8611), .B(n8618), .Z(n8630) );
  NOR U8462 ( .A(n8579), .B(n8653), .Z(n8618) );
  XOR U8463 ( .A(n8623), .B(n8622), .Z(n8611) );
  XNOR U8464 ( .A(n8654), .B(n8619), .Z(n8622) );
  XOR U8465 ( .A(n8655), .B(n8656), .Z(n8619) );
  AND U8466 ( .A(n8657), .B(n8658), .Z(n8656) );
  XOR U8467 ( .A(n8655), .B(n8659), .Z(n8657) );
  XNOR U8468 ( .A(n8660), .B(n8661), .Z(n8654) );
  NOR U8469 ( .A(n8662), .B(n8663), .Z(n8661) );
  XNOR U8470 ( .A(n8660), .B(n8664), .Z(n8662) );
  XOR U8471 ( .A(n8665), .B(n8666), .Z(n8623) );
  NOR U8472 ( .A(n8667), .B(n8668), .Z(n8666) );
  XNOR U8473 ( .A(n8665), .B(n8669), .Z(n8667) );
  XNOR U8474 ( .A(n8568), .B(n8626), .Z(n8628) );
  XNOR U8475 ( .A(n8670), .B(n8671), .Z(n8568) );
  AND U8476 ( .A(n61), .B(n8575), .Z(n8671) );
  XOR U8477 ( .A(n8670), .B(n8573), .Z(n8575) );
  AND U8478 ( .A(n8576), .B(n8579), .Z(n8626) );
  XOR U8479 ( .A(n8672), .B(n8653), .Z(n8579) );
  XNOR U8480 ( .A(p_input[1024]), .B(p_input[32]), .Z(n8653) );
  XOR U8481 ( .A(n8641), .B(n8640), .Z(n8672) );
  XNOR U8482 ( .A(n8673), .B(n8647), .Z(n8640) );
  XNOR U8483 ( .A(n8636), .B(n8635), .Z(n8647) );
  XOR U8484 ( .A(n8674), .B(n8632), .Z(n8635) );
  XOR U8485 ( .A(p_input[1034]), .B(p_input[42]), .Z(n8632) );
  XNOR U8486 ( .A(p_input[1035]), .B(p_input[43]), .Z(n8674) );
  XOR U8487 ( .A(p_input[1036]), .B(p_input[44]), .Z(n8636) );
  XNOR U8488 ( .A(n8646), .B(n8637), .Z(n8673) );
  XOR U8489 ( .A(p_input[1025]), .B(p_input[33]), .Z(n8637) );
  XOR U8490 ( .A(n8675), .B(n8652), .Z(n8646) );
  XNOR U8491 ( .A(p_input[1039]), .B(p_input[47]), .Z(n8652) );
  XOR U8492 ( .A(n8643), .B(n8651), .Z(n8675) );
  XOR U8493 ( .A(n8676), .B(n8648), .Z(n8651) );
  XOR U8494 ( .A(p_input[1037]), .B(p_input[45]), .Z(n8648) );
  XNOR U8495 ( .A(p_input[1038]), .B(p_input[46]), .Z(n8676) );
  XOR U8496 ( .A(p_input[1033]), .B(p_input[41]), .Z(n8643) );
  XNOR U8497 ( .A(n8659), .B(n8658), .Z(n8641) );
  XNOR U8498 ( .A(n8677), .B(n8664), .Z(n8658) );
  XOR U8499 ( .A(p_input[1032]), .B(p_input[40]), .Z(n8664) );
  XOR U8500 ( .A(n8655), .B(n8663), .Z(n8677) );
  XOR U8501 ( .A(n8678), .B(n8660), .Z(n8663) );
  XOR U8502 ( .A(p_input[1030]), .B(p_input[38]), .Z(n8660) );
  XNOR U8503 ( .A(p_input[1031]), .B(p_input[39]), .Z(n8678) );
  XOR U8504 ( .A(p_input[1026]), .B(p_input[34]), .Z(n8655) );
  XNOR U8505 ( .A(n8669), .B(n8668), .Z(n8659) );
  XOR U8506 ( .A(n8679), .B(n8665), .Z(n8668) );
  XOR U8507 ( .A(p_input[1027]), .B(p_input[35]), .Z(n8665) );
  XNOR U8508 ( .A(p_input[1028]), .B(p_input[36]), .Z(n8679) );
  XOR U8509 ( .A(p_input[1029]), .B(p_input[37]), .Z(n8669) );
  XNOR U8510 ( .A(n8680), .B(n8681), .Z(n8576) );
  AND U8511 ( .A(n61), .B(n8682), .Z(n8681) );
  XNOR U8512 ( .A(n8683), .B(n8684), .Z(n61) );
  AND U8513 ( .A(n8685), .B(n8686), .Z(n8684) );
  XOR U8514 ( .A(n8683), .B(n8586), .Z(n8686) );
  XNOR U8515 ( .A(n8683), .B(n8540), .Z(n8685) );
  XOR U8516 ( .A(n8687), .B(n8688), .Z(n8683) );
  AND U8517 ( .A(n8689), .B(n8690), .Z(n8688) );
  XOR U8518 ( .A(n8687), .B(n8550), .Z(n8689) );
  XOR U8519 ( .A(n8691), .B(n8692), .Z(n8529) );
  AND U8520 ( .A(n65), .B(n8682), .Z(n8692) );
  XNOR U8521 ( .A(n8680), .B(n8691), .Z(n8682) );
  XNOR U8522 ( .A(n8693), .B(n8694), .Z(n65) );
  AND U8523 ( .A(n8695), .B(n8696), .Z(n8694) );
  XNOR U8524 ( .A(n8697), .B(n8693), .Z(n8696) );
  IV U8525 ( .A(n8586), .Z(n8697) );
  XNOR U8526 ( .A(n8698), .B(n8699), .Z(n8586) );
  AND U8527 ( .A(n68), .B(n8700), .Z(n8699) );
  XNOR U8528 ( .A(n8698), .B(n8701), .Z(n8700) );
  XNOR U8529 ( .A(n8540), .B(n8693), .Z(n8695) );
  XOR U8530 ( .A(n8702), .B(n8703), .Z(n8540) );
  AND U8531 ( .A(n76), .B(n8704), .Z(n8703) );
  XOR U8532 ( .A(n8687), .B(n8705), .Z(n8693) );
  AND U8533 ( .A(n8706), .B(n8690), .Z(n8705) );
  XNOR U8534 ( .A(n8599), .B(n8687), .Z(n8690) );
  XNOR U8535 ( .A(n8707), .B(n8708), .Z(n8599) );
  AND U8536 ( .A(n68), .B(n8709), .Z(n8708) );
  XOR U8537 ( .A(n8710), .B(n8707), .Z(n8709) );
  XNOR U8538 ( .A(n8711), .B(n8687), .Z(n8706) );
  IV U8539 ( .A(n8550), .Z(n8711) );
  XOR U8540 ( .A(n8712), .B(n8713), .Z(n8550) );
  AND U8541 ( .A(n76), .B(n8714), .Z(n8713) );
  XOR U8542 ( .A(n8715), .B(n8716), .Z(n8687) );
  AND U8543 ( .A(n8717), .B(n8718), .Z(n8716) );
  XNOR U8544 ( .A(n8624), .B(n8715), .Z(n8718) );
  XNOR U8545 ( .A(n8719), .B(n8720), .Z(n8624) );
  AND U8546 ( .A(n68), .B(n8721), .Z(n8720) );
  XNOR U8547 ( .A(n8722), .B(n8719), .Z(n8721) );
  XOR U8548 ( .A(n8715), .B(n8561), .Z(n8717) );
  XOR U8549 ( .A(n8723), .B(n8724), .Z(n8561) );
  AND U8550 ( .A(n76), .B(n8725), .Z(n8724) );
  XOR U8551 ( .A(n8726), .B(n8727), .Z(n8715) );
  AND U8552 ( .A(n8728), .B(n8729), .Z(n8727) );
  XNOR U8553 ( .A(n8726), .B(n8670), .Z(n8729) );
  XNOR U8554 ( .A(n8730), .B(n8731), .Z(n8670) );
  AND U8555 ( .A(n68), .B(n8732), .Z(n8731) );
  XOR U8556 ( .A(n8733), .B(n8730), .Z(n8732) );
  XNOR U8557 ( .A(n8734), .B(n8726), .Z(n8728) );
  IV U8558 ( .A(n8573), .Z(n8734) );
  XOR U8559 ( .A(n8735), .B(n8736), .Z(n8573) );
  AND U8560 ( .A(n76), .B(n8737), .Z(n8736) );
  AND U8561 ( .A(n8691), .B(n8680), .Z(n8726) );
  XNOR U8562 ( .A(n8738), .B(n8739), .Z(n8680) );
  AND U8563 ( .A(n68), .B(n8740), .Z(n8739) );
  XNOR U8564 ( .A(n8741), .B(n8738), .Z(n8740) );
  XNOR U8565 ( .A(n8742), .B(n8743), .Z(n68) );
  AND U8566 ( .A(n8744), .B(n8745), .Z(n8743) );
  XOR U8567 ( .A(n8701), .B(n8742), .Z(n8745) );
  AND U8568 ( .A(n8746), .B(n8747), .Z(n8701) );
  XOR U8569 ( .A(n8742), .B(n8698), .Z(n8744) );
  XNOR U8570 ( .A(n8748), .B(n8749), .Z(n8698) );
  AND U8571 ( .A(n72), .B(n8704), .Z(n8749) );
  XOR U8572 ( .A(n8702), .B(n8748), .Z(n8704) );
  XOR U8573 ( .A(n8750), .B(n8751), .Z(n8742) );
  AND U8574 ( .A(n8752), .B(n8753), .Z(n8751) );
  XNOR U8575 ( .A(n8750), .B(n8746), .Z(n8753) );
  IV U8576 ( .A(n8710), .Z(n8746) );
  XOR U8577 ( .A(n8754), .B(n8755), .Z(n8710) );
  XOR U8578 ( .A(n8756), .B(n8747), .Z(n8755) );
  AND U8579 ( .A(n8722), .B(n8757), .Z(n8747) );
  AND U8580 ( .A(n8758), .B(n8759), .Z(n8756) );
  XOR U8581 ( .A(n8760), .B(n8754), .Z(n8758) );
  XNOR U8582 ( .A(n8707), .B(n8750), .Z(n8752) );
  XNOR U8583 ( .A(n8761), .B(n8762), .Z(n8707) );
  AND U8584 ( .A(n72), .B(n8714), .Z(n8762) );
  XOR U8585 ( .A(n8761), .B(n8712), .Z(n8714) );
  XOR U8586 ( .A(n8763), .B(n8764), .Z(n8750) );
  AND U8587 ( .A(n8765), .B(n8766), .Z(n8764) );
  XNOR U8588 ( .A(n8763), .B(n8722), .Z(n8766) );
  XOR U8589 ( .A(n8767), .B(n8759), .Z(n8722) );
  XNOR U8590 ( .A(n8768), .B(n8754), .Z(n8759) );
  XOR U8591 ( .A(n8769), .B(n8770), .Z(n8754) );
  AND U8592 ( .A(n8771), .B(n8772), .Z(n8770) );
  XOR U8593 ( .A(n8773), .B(n8769), .Z(n8771) );
  XNOR U8594 ( .A(n8774), .B(n8775), .Z(n8768) );
  AND U8595 ( .A(n8776), .B(n8777), .Z(n8775) );
  XOR U8596 ( .A(n8774), .B(n8778), .Z(n8776) );
  XNOR U8597 ( .A(n8760), .B(n8757), .Z(n8767) );
  AND U8598 ( .A(n8779), .B(n8780), .Z(n8757) );
  XOR U8599 ( .A(n8781), .B(n8782), .Z(n8760) );
  AND U8600 ( .A(n8783), .B(n8784), .Z(n8782) );
  XOR U8601 ( .A(n8781), .B(n8785), .Z(n8783) );
  XNOR U8602 ( .A(n8719), .B(n8763), .Z(n8765) );
  XNOR U8603 ( .A(n8786), .B(n8787), .Z(n8719) );
  AND U8604 ( .A(n72), .B(n8725), .Z(n8787) );
  XOR U8605 ( .A(n8786), .B(n8723), .Z(n8725) );
  XOR U8606 ( .A(n8788), .B(n8789), .Z(n8763) );
  AND U8607 ( .A(n8790), .B(n8791), .Z(n8789) );
  XNOR U8608 ( .A(n8788), .B(n8779), .Z(n8791) );
  IV U8609 ( .A(n8733), .Z(n8779) );
  XNOR U8610 ( .A(n8792), .B(n8772), .Z(n8733) );
  XNOR U8611 ( .A(n8793), .B(n8778), .Z(n8772) );
  XOR U8612 ( .A(n8794), .B(n8795), .Z(n8778) );
  NOR U8613 ( .A(n8796), .B(n8797), .Z(n8795) );
  XNOR U8614 ( .A(n8794), .B(n8798), .Z(n8796) );
  XNOR U8615 ( .A(n8777), .B(n8769), .Z(n8793) );
  XOR U8616 ( .A(n8799), .B(n8800), .Z(n8769) );
  AND U8617 ( .A(n8801), .B(n8802), .Z(n8800) );
  XNOR U8618 ( .A(n8799), .B(n8803), .Z(n8801) );
  XNOR U8619 ( .A(n8804), .B(n8774), .Z(n8777) );
  XOR U8620 ( .A(n8805), .B(n8806), .Z(n8774) );
  AND U8621 ( .A(n8807), .B(n8808), .Z(n8806) );
  XOR U8622 ( .A(n8805), .B(n8809), .Z(n8807) );
  XNOR U8623 ( .A(n8810), .B(n8811), .Z(n8804) );
  NOR U8624 ( .A(n8812), .B(n8813), .Z(n8811) );
  XOR U8625 ( .A(n8810), .B(n8814), .Z(n8812) );
  XNOR U8626 ( .A(n8773), .B(n8780), .Z(n8792) );
  NOR U8627 ( .A(n8741), .B(n8815), .Z(n8780) );
  XOR U8628 ( .A(n8785), .B(n8784), .Z(n8773) );
  XNOR U8629 ( .A(n8816), .B(n8781), .Z(n8784) );
  XOR U8630 ( .A(n8817), .B(n8818), .Z(n8781) );
  AND U8631 ( .A(n8819), .B(n8820), .Z(n8818) );
  XOR U8632 ( .A(n8817), .B(n8821), .Z(n8819) );
  XNOR U8633 ( .A(n8822), .B(n8823), .Z(n8816) );
  NOR U8634 ( .A(n8824), .B(n8825), .Z(n8823) );
  XNOR U8635 ( .A(n8822), .B(n8826), .Z(n8824) );
  XOR U8636 ( .A(n8827), .B(n8828), .Z(n8785) );
  NOR U8637 ( .A(n8829), .B(n8830), .Z(n8828) );
  XNOR U8638 ( .A(n8827), .B(n8831), .Z(n8829) );
  XNOR U8639 ( .A(n8730), .B(n8788), .Z(n8790) );
  XNOR U8640 ( .A(n8832), .B(n8833), .Z(n8730) );
  AND U8641 ( .A(n72), .B(n8737), .Z(n8833) );
  XOR U8642 ( .A(n8832), .B(n8735), .Z(n8737) );
  AND U8643 ( .A(n8738), .B(n8741), .Z(n8788) );
  XOR U8644 ( .A(n8834), .B(n8815), .Z(n8741) );
  XNOR U8645 ( .A(p_input[1024]), .B(p_input[48]), .Z(n8815) );
  XOR U8646 ( .A(n8803), .B(n8802), .Z(n8834) );
  XNOR U8647 ( .A(n8835), .B(n8809), .Z(n8802) );
  XNOR U8648 ( .A(n8798), .B(n8797), .Z(n8809) );
  XOR U8649 ( .A(n8836), .B(n8794), .Z(n8797) );
  XOR U8650 ( .A(p_input[1034]), .B(p_input[58]), .Z(n8794) );
  XNOR U8651 ( .A(p_input[1035]), .B(p_input[59]), .Z(n8836) );
  XOR U8652 ( .A(p_input[1036]), .B(p_input[60]), .Z(n8798) );
  XNOR U8653 ( .A(n8808), .B(n8799), .Z(n8835) );
  XOR U8654 ( .A(p_input[1025]), .B(p_input[49]), .Z(n8799) );
  XOR U8655 ( .A(n8837), .B(n8814), .Z(n8808) );
  XNOR U8656 ( .A(p_input[1039]), .B(p_input[63]), .Z(n8814) );
  XOR U8657 ( .A(n8805), .B(n8813), .Z(n8837) );
  XOR U8658 ( .A(n8838), .B(n8810), .Z(n8813) );
  XOR U8659 ( .A(p_input[1037]), .B(p_input[61]), .Z(n8810) );
  XNOR U8660 ( .A(p_input[1038]), .B(p_input[62]), .Z(n8838) );
  XOR U8661 ( .A(p_input[1033]), .B(p_input[57]), .Z(n8805) );
  XNOR U8662 ( .A(n8821), .B(n8820), .Z(n8803) );
  XNOR U8663 ( .A(n8839), .B(n8826), .Z(n8820) );
  XOR U8664 ( .A(p_input[1032]), .B(p_input[56]), .Z(n8826) );
  XOR U8665 ( .A(n8817), .B(n8825), .Z(n8839) );
  XOR U8666 ( .A(n8840), .B(n8822), .Z(n8825) );
  XOR U8667 ( .A(p_input[1030]), .B(p_input[54]), .Z(n8822) );
  XNOR U8668 ( .A(p_input[1031]), .B(p_input[55]), .Z(n8840) );
  XOR U8669 ( .A(p_input[1026]), .B(p_input[50]), .Z(n8817) );
  XNOR U8670 ( .A(n8831), .B(n8830), .Z(n8821) );
  XOR U8671 ( .A(n8841), .B(n8827), .Z(n8830) );
  XOR U8672 ( .A(p_input[1027]), .B(p_input[51]), .Z(n8827) );
  XNOR U8673 ( .A(p_input[1028]), .B(p_input[52]), .Z(n8841) );
  XOR U8674 ( .A(p_input[1029]), .B(p_input[53]), .Z(n8831) );
  XNOR U8675 ( .A(n8842), .B(n8843), .Z(n8738) );
  AND U8676 ( .A(n72), .B(n8844), .Z(n8843) );
  XNOR U8677 ( .A(n8845), .B(n8846), .Z(n72) );
  AND U8678 ( .A(n8847), .B(n8848), .Z(n8846) );
  XOR U8679 ( .A(n8845), .B(n8748), .Z(n8848) );
  XNOR U8680 ( .A(n8845), .B(n8702), .Z(n8847) );
  XOR U8681 ( .A(n8849), .B(n8850), .Z(n8845) );
  AND U8682 ( .A(n8851), .B(n8852), .Z(n8850) );
  XOR U8683 ( .A(n8849), .B(n8712), .Z(n8851) );
  XOR U8684 ( .A(n8853), .B(n8854), .Z(n8691) );
  AND U8685 ( .A(n76), .B(n8844), .Z(n8854) );
  XNOR U8686 ( .A(n8842), .B(n8853), .Z(n8844) );
  XNOR U8687 ( .A(n8855), .B(n8856), .Z(n76) );
  AND U8688 ( .A(n8857), .B(n8858), .Z(n8856) );
  XNOR U8689 ( .A(n8859), .B(n8855), .Z(n8858) );
  IV U8690 ( .A(n8748), .Z(n8859) );
  XNOR U8691 ( .A(n8860), .B(n8861), .Z(n8748) );
  AND U8692 ( .A(n79), .B(n8862), .Z(n8861) );
  XNOR U8693 ( .A(n8860), .B(n8863), .Z(n8862) );
  XNOR U8694 ( .A(n8702), .B(n8855), .Z(n8857) );
  XOR U8695 ( .A(n8864), .B(n8865), .Z(n8702) );
  AND U8696 ( .A(n87), .B(n8866), .Z(n8865) );
  XOR U8697 ( .A(n8849), .B(n8867), .Z(n8855) );
  AND U8698 ( .A(n8868), .B(n8852), .Z(n8867) );
  XNOR U8699 ( .A(n8761), .B(n8849), .Z(n8852) );
  XNOR U8700 ( .A(n8869), .B(n8870), .Z(n8761) );
  AND U8701 ( .A(n79), .B(n8871), .Z(n8870) );
  XOR U8702 ( .A(n8872), .B(n8869), .Z(n8871) );
  XNOR U8703 ( .A(n8873), .B(n8849), .Z(n8868) );
  IV U8704 ( .A(n8712), .Z(n8873) );
  XOR U8705 ( .A(n8874), .B(n8875), .Z(n8712) );
  AND U8706 ( .A(n87), .B(n8876), .Z(n8875) );
  XOR U8707 ( .A(n8877), .B(n8878), .Z(n8849) );
  AND U8708 ( .A(n8879), .B(n8880), .Z(n8878) );
  XNOR U8709 ( .A(n8786), .B(n8877), .Z(n8880) );
  XNOR U8710 ( .A(n8881), .B(n8882), .Z(n8786) );
  AND U8711 ( .A(n79), .B(n8883), .Z(n8882) );
  XNOR U8712 ( .A(n8884), .B(n8881), .Z(n8883) );
  XOR U8713 ( .A(n8877), .B(n8723), .Z(n8879) );
  XOR U8714 ( .A(n8885), .B(n8886), .Z(n8723) );
  AND U8715 ( .A(n87), .B(n8887), .Z(n8886) );
  XOR U8716 ( .A(n8888), .B(n8889), .Z(n8877) );
  AND U8717 ( .A(n8890), .B(n8891), .Z(n8889) );
  XNOR U8718 ( .A(n8888), .B(n8832), .Z(n8891) );
  XNOR U8719 ( .A(n8892), .B(n8893), .Z(n8832) );
  AND U8720 ( .A(n79), .B(n8894), .Z(n8893) );
  XOR U8721 ( .A(n8895), .B(n8892), .Z(n8894) );
  XNOR U8722 ( .A(n8896), .B(n8888), .Z(n8890) );
  IV U8723 ( .A(n8735), .Z(n8896) );
  XOR U8724 ( .A(n8897), .B(n8898), .Z(n8735) );
  AND U8725 ( .A(n87), .B(n8899), .Z(n8898) );
  AND U8726 ( .A(n8853), .B(n8842), .Z(n8888) );
  XNOR U8727 ( .A(n8900), .B(n8901), .Z(n8842) );
  AND U8728 ( .A(n79), .B(n8902), .Z(n8901) );
  XNOR U8729 ( .A(n8903), .B(n8900), .Z(n8902) );
  XNOR U8730 ( .A(n8904), .B(n8905), .Z(n79) );
  AND U8731 ( .A(n8906), .B(n8907), .Z(n8905) );
  XOR U8732 ( .A(n8863), .B(n8904), .Z(n8907) );
  AND U8733 ( .A(n8908), .B(n8909), .Z(n8863) );
  XOR U8734 ( .A(n8904), .B(n8860), .Z(n8906) );
  XNOR U8735 ( .A(n8910), .B(n8911), .Z(n8860) );
  AND U8736 ( .A(n83), .B(n8866), .Z(n8911) );
  XOR U8737 ( .A(n8864), .B(n8910), .Z(n8866) );
  XOR U8738 ( .A(n8912), .B(n8913), .Z(n8904) );
  AND U8739 ( .A(n8914), .B(n8915), .Z(n8913) );
  XNOR U8740 ( .A(n8912), .B(n8908), .Z(n8915) );
  IV U8741 ( .A(n8872), .Z(n8908) );
  XOR U8742 ( .A(n8916), .B(n8917), .Z(n8872) );
  XOR U8743 ( .A(n8918), .B(n8909), .Z(n8917) );
  AND U8744 ( .A(n8884), .B(n8919), .Z(n8909) );
  AND U8745 ( .A(n8920), .B(n8921), .Z(n8918) );
  XOR U8746 ( .A(n8922), .B(n8916), .Z(n8920) );
  XNOR U8747 ( .A(n8869), .B(n8912), .Z(n8914) );
  XNOR U8748 ( .A(n8923), .B(n8924), .Z(n8869) );
  AND U8749 ( .A(n83), .B(n8876), .Z(n8924) );
  XOR U8750 ( .A(n8923), .B(n8874), .Z(n8876) );
  XOR U8751 ( .A(n8925), .B(n8926), .Z(n8912) );
  AND U8752 ( .A(n8927), .B(n8928), .Z(n8926) );
  XNOR U8753 ( .A(n8925), .B(n8884), .Z(n8928) );
  XOR U8754 ( .A(n8929), .B(n8921), .Z(n8884) );
  XNOR U8755 ( .A(n8930), .B(n8916), .Z(n8921) );
  XOR U8756 ( .A(n8931), .B(n8932), .Z(n8916) );
  AND U8757 ( .A(n8933), .B(n8934), .Z(n8932) );
  XOR U8758 ( .A(n8935), .B(n8931), .Z(n8933) );
  XNOR U8759 ( .A(n8936), .B(n8937), .Z(n8930) );
  AND U8760 ( .A(n8938), .B(n8939), .Z(n8937) );
  XOR U8761 ( .A(n8936), .B(n8940), .Z(n8938) );
  XNOR U8762 ( .A(n8922), .B(n8919), .Z(n8929) );
  AND U8763 ( .A(n8941), .B(n8942), .Z(n8919) );
  XOR U8764 ( .A(n8943), .B(n8944), .Z(n8922) );
  AND U8765 ( .A(n8945), .B(n8946), .Z(n8944) );
  XOR U8766 ( .A(n8943), .B(n8947), .Z(n8945) );
  XNOR U8767 ( .A(n8881), .B(n8925), .Z(n8927) );
  XNOR U8768 ( .A(n8948), .B(n8949), .Z(n8881) );
  AND U8769 ( .A(n83), .B(n8887), .Z(n8949) );
  XOR U8770 ( .A(n8948), .B(n8885), .Z(n8887) );
  XOR U8771 ( .A(n8950), .B(n8951), .Z(n8925) );
  AND U8772 ( .A(n8952), .B(n8953), .Z(n8951) );
  XNOR U8773 ( .A(n8950), .B(n8941), .Z(n8953) );
  IV U8774 ( .A(n8895), .Z(n8941) );
  XNOR U8775 ( .A(n8954), .B(n8934), .Z(n8895) );
  XNOR U8776 ( .A(n8955), .B(n8940), .Z(n8934) );
  XOR U8777 ( .A(n8956), .B(n8957), .Z(n8940) );
  NOR U8778 ( .A(n8958), .B(n8959), .Z(n8957) );
  XNOR U8779 ( .A(n8956), .B(n8960), .Z(n8958) );
  XNOR U8780 ( .A(n8939), .B(n8931), .Z(n8955) );
  XOR U8781 ( .A(n8961), .B(n8962), .Z(n8931) );
  AND U8782 ( .A(n8963), .B(n8964), .Z(n8962) );
  XNOR U8783 ( .A(n8961), .B(n8965), .Z(n8963) );
  XNOR U8784 ( .A(n8966), .B(n8936), .Z(n8939) );
  XOR U8785 ( .A(n8967), .B(n8968), .Z(n8936) );
  AND U8786 ( .A(n8969), .B(n8970), .Z(n8968) );
  XOR U8787 ( .A(n8967), .B(n8971), .Z(n8969) );
  XNOR U8788 ( .A(n8972), .B(n8973), .Z(n8966) );
  NOR U8789 ( .A(n8974), .B(n8975), .Z(n8973) );
  XOR U8790 ( .A(n8972), .B(n8976), .Z(n8974) );
  XNOR U8791 ( .A(n8935), .B(n8942), .Z(n8954) );
  NOR U8792 ( .A(n8903), .B(n8977), .Z(n8942) );
  XOR U8793 ( .A(n8947), .B(n8946), .Z(n8935) );
  XNOR U8794 ( .A(n8978), .B(n8943), .Z(n8946) );
  XOR U8795 ( .A(n8979), .B(n8980), .Z(n8943) );
  AND U8796 ( .A(n8981), .B(n8982), .Z(n8980) );
  XOR U8797 ( .A(n8979), .B(n8983), .Z(n8981) );
  XNOR U8798 ( .A(n8984), .B(n8985), .Z(n8978) );
  NOR U8799 ( .A(n8986), .B(n8987), .Z(n8985) );
  XNOR U8800 ( .A(n8984), .B(n8988), .Z(n8986) );
  XOR U8801 ( .A(n8989), .B(n8990), .Z(n8947) );
  NOR U8802 ( .A(n8991), .B(n8992), .Z(n8990) );
  XNOR U8803 ( .A(n8989), .B(n8993), .Z(n8991) );
  XNOR U8804 ( .A(n8892), .B(n8950), .Z(n8952) );
  XNOR U8805 ( .A(n8994), .B(n8995), .Z(n8892) );
  AND U8806 ( .A(n83), .B(n8899), .Z(n8995) );
  XOR U8807 ( .A(n8994), .B(n8897), .Z(n8899) );
  AND U8808 ( .A(n8900), .B(n8903), .Z(n8950) );
  XOR U8809 ( .A(n8996), .B(n8977), .Z(n8903) );
  XNOR U8810 ( .A(p_input[1024]), .B(p_input[64]), .Z(n8977) );
  XOR U8811 ( .A(n8965), .B(n8964), .Z(n8996) );
  XNOR U8812 ( .A(n8997), .B(n8971), .Z(n8964) );
  XNOR U8813 ( .A(n8960), .B(n8959), .Z(n8971) );
  XOR U8814 ( .A(n8998), .B(n8956), .Z(n8959) );
  XOR U8815 ( .A(p_input[1034]), .B(p_input[74]), .Z(n8956) );
  XNOR U8816 ( .A(p_input[1035]), .B(p_input[75]), .Z(n8998) );
  XOR U8817 ( .A(p_input[1036]), .B(p_input[76]), .Z(n8960) );
  XNOR U8818 ( .A(n8970), .B(n8961), .Z(n8997) );
  XOR U8819 ( .A(p_input[1025]), .B(p_input[65]), .Z(n8961) );
  XOR U8820 ( .A(n8999), .B(n8976), .Z(n8970) );
  XNOR U8821 ( .A(p_input[1039]), .B(p_input[79]), .Z(n8976) );
  XOR U8822 ( .A(n8967), .B(n8975), .Z(n8999) );
  XOR U8823 ( .A(n9000), .B(n8972), .Z(n8975) );
  XOR U8824 ( .A(p_input[1037]), .B(p_input[77]), .Z(n8972) );
  XNOR U8825 ( .A(p_input[1038]), .B(p_input[78]), .Z(n9000) );
  XOR U8826 ( .A(p_input[1033]), .B(p_input[73]), .Z(n8967) );
  XNOR U8827 ( .A(n8983), .B(n8982), .Z(n8965) );
  XNOR U8828 ( .A(n9001), .B(n8988), .Z(n8982) );
  XOR U8829 ( .A(p_input[1032]), .B(p_input[72]), .Z(n8988) );
  XOR U8830 ( .A(n8979), .B(n8987), .Z(n9001) );
  XOR U8831 ( .A(n9002), .B(n8984), .Z(n8987) );
  XOR U8832 ( .A(p_input[1030]), .B(p_input[70]), .Z(n8984) );
  XNOR U8833 ( .A(p_input[1031]), .B(p_input[71]), .Z(n9002) );
  XOR U8834 ( .A(p_input[1026]), .B(p_input[66]), .Z(n8979) );
  XNOR U8835 ( .A(n8993), .B(n8992), .Z(n8983) );
  XOR U8836 ( .A(n9003), .B(n8989), .Z(n8992) );
  XOR U8837 ( .A(p_input[1027]), .B(p_input[67]), .Z(n8989) );
  XNOR U8838 ( .A(p_input[1028]), .B(p_input[68]), .Z(n9003) );
  XOR U8839 ( .A(p_input[1029]), .B(p_input[69]), .Z(n8993) );
  XNOR U8840 ( .A(n9004), .B(n9005), .Z(n8900) );
  AND U8841 ( .A(n83), .B(n9006), .Z(n9005) );
  XNOR U8842 ( .A(n9007), .B(n9008), .Z(n83) );
  AND U8843 ( .A(n9009), .B(n9010), .Z(n9008) );
  XOR U8844 ( .A(n9007), .B(n8910), .Z(n9010) );
  XNOR U8845 ( .A(n9007), .B(n8864), .Z(n9009) );
  XOR U8846 ( .A(n9011), .B(n9012), .Z(n9007) );
  AND U8847 ( .A(n9013), .B(n9014), .Z(n9012) );
  XOR U8848 ( .A(n9011), .B(n8874), .Z(n9013) );
  XOR U8849 ( .A(n9015), .B(n9016), .Z(n8853) );
  AND U8850 ( .A(n87), .B(n9006), .Z(n9016) );
  XNOR U8851 ( .A(n9004), .B(n9015), .Z(n9006) );
  XNOR U8852 ( .A(n9017), .B(n9018), .Z(n87) );
  AND U8853 ( .A(n9019), .B(n9020), .Z(n9018) );
  XNOR U8854 ( .A(n9021), .B(n9017), .Z(n9020) );
  IV U8855 ( .A(n8910), .Z(n9021) );
  XNOR U8856 ( .A(n9022), .B(n9023), .Z(n8910) );
  AND U8857 ( .A(n90), .B(n9024), .Z(n9023) );
  XNOR U8858 ( .A(n9022), .B(n9025), .Z(n9024) );
  XNOR U8859 ( .A(n8864), .B(n9017), .Z(n9019) );
  XOR U8860 ( .A(n9026), .B(n9027), .Z(n8864) );
  AND U8861 ( .A(n98), .B(n9028), .Z(n9027) );
  XOR U8862 ( .A(n9011), .B(n9029), .Z(n9017) );
  AND U8863 ( .A(n9030), .B(n9014), .Z(n9029) );
  XNOR U8864 ( .A(n8923), .B(n9011), .Z(n9014) );
  XNOR U8865 ( .A(n9031), .B(n9032), .Z(n8923) );
  AND U8866 ( .A(n90), .B(n9033), .Z(n9032) );
  XOR U8867 ( .A(n9034), .B(n9031), .Z(n9033) );
  XNOR U8868 ( .A(n9035), .B(n9011), .Z(n9030) );
  IV U8869 ( .A(n8874), .Z(n9035) );
  XOR U8870 ( .A(n9036), .B(n9037), .Z(n8874) );
  AND U8871 ( .A(n98), .B(n9038), .Z(n9037) );
  XOR U8872 ( .A(n9039), .B(n9040), .Z(n9011) );
  AND U8873 ( .A(n9041), .B(n9042), .Z(n9040) );
  XNOR U8874 ( .A(n8948), .B(n9039), .Z(n9042) );
  XNOR U8875 ( .A(n9043), .B(n9044), .Z(n8948) );
  AND U8876 ( .A(n90), .B(n9045), .Z(n9044) );
  XNOR U8877 ( .A(n9046), .B(n9043), .Z(n9045) );
  XOR U8878 ( .A(n9039), .B(n8885), .Z(n9041) );
  XOR U8879 ( .A(n9047), .B(n9048), .Z(n8885) );
  AND U8880 ( .A(n98), .B(n9049), .Z(n9048) );
  XOR U8881 ( .A(n9050), .B(n9051), .Z(n9039) );
  AND U8882 ( .A(n9052), .B(n9053), .Z(n9051) );
  XNOR U8883 ( .A(n9050), .B(n8994), .Z(n9053) );
  XNOR U8884 ( .A(n9054), .B(n9055), .Z(n8994) );
  AND U8885 ( .A(n90), .B(n9056), .Z(n9055) );
  XOR U8886 ( .A(n9057), .B(n9054), .Z(n9056) );
  XNOR U8887 ( .A(n9058), .B(n9050), .Z(n9052) );
  IV U8888 ( .A(n8897), .Z(n9058) );
  XOR U8889 ( .A(n9059), .B(n9060), .Z(n8897) );
  AND U8890 ( .A(n98), .B(n9061), .Z(n9060) );
  AND U8891 ( .A(n9015), .B(n9004), .Z(n9050) );
  XNOR U8892 ( .A(n9062), .B(n9063), .Z(n9004) );
  AND U8893 ( .A(n90), .B(n9064), .Z(n9063) );
  XNOR U8894 ( .A(n9065), .B(n9062), .Z(n9064) );
  XNOR U8895 ( .A(n9066), .B(n9067), .Z(n90) );
  AND U8896 ( .A(n9068), .B(n9069), .Z(n9067) );
  XOR U8897 ( .A(n9025), .B(n9066), .Z(n9069) );
  AND U8898 ( .A(n9070), .B(n9071), .Z(n9025) );
  XOR U8899 ( .A(n9066), .B(n9022), .Z(n9068) );
  XNOR U8900 ( .A(n9072), .B(n9073), .Z(n9022) );
  AND U8901 ( .A(n94), .B(n9028), .Z(n9073) );
  XOR U8902 ( .A(n9026), .B(n9072), .Z(n9028) );
  XOR U8903 ( .A(n9074), .B(n9075), .Z(n9066) );
  AND U8904 ( .A(n9076), .B(n9077), .Z(n9075) );
  XNOR U8905 ( .A(n9074), .B(n9070), .Z(n9077) );
  IV U8906 ( .A(n9034), .Z(n9070) );
  XOR U8907 ( .A(n9078), .B(n9079), .Z(n9034) );
  XOR U8908 ( .A(n9080), .B(n9071), .Z(n9079) );
  AND U8909 ( .A(n9046), .B(n9081), .Z(n9071) );
  AND U8910 ( .A(n9082), .B(n9083), .Z(n9080) );
  XOR U8911 ( .A(n9084), .B(n9078), .Z(n9082) );
  XNOR U8912 ( .A(n9031), .B(n9074), .Z(n9076) );
  XNOR U8913 ( .A(n9085), .B(n9086), .Z(n9031) );
  AND U8914 ( .A(n94), .B(n9038), .Z(n9086) );
  XOR U8915 ( .A(n9085), .B(n9036), .Z(n9038) );
  XOR U8916 ( .A(n9087), .B(n9088), .Z(n9074) );
  AND U8917 ( .A(n9089), .B(n9090), .Z(n9088) );
  XNOR U8918 ( .A(n9087), .B(n9046), .Z(n9090) );
  XOR U8919 ( .A(n9091), .B(n9083), .Z(n9046) );
  XNOR U8920 ( .A(n9092), .B(n9078), .Z(n9083) );
  XOR U8921 ( .A(n9093), .B(n9094), .Z(n9078) );
  AND U8922 ( .A(n9095), .B(n9096), .Z(n9094) );
  XOR U8923 ( .A(n9097), .B(n9093), .Z(n9095) );
  XNOR U8924 ( .A(n9098), .B(n9099), .Z(n9092) );
  AND U8925 ( .A(n9100), .B(n9101), .Z(n9099) );
  XOR U8926 ( .A(n9098), .B(n9102), .Z(n9100) );
  XNOR U8927 ( .A(n9084), .B(n9081), .Z(n9091) );
  AND U8928 ( .A(n9103), .B(n9104), .Z(n9081) );
  XOR U8929 ( .A(n9105), .B(n9106), .Z(n9084) );
  AND U8930 ( .A(n9107), .B(n9108), .Z(n9106) );
  XOR U8931 ( .A(n9105), .B(n9109), .Z(n9107) );
  XNOR U8932 ( .A(n9043), .B(n9087), .Z(n9089) );
  XNOR U8933 ( .A(n9110), .B(n9111), .Z(n9043) );
  AND U8934 ( .A(n94), .B(n9049), .Z(n9111) );
  XOR U8935 ( .A(n9110), .B(n9047), .Z(n9049) );
  XOR U8936 ( .A(n9112), .B(n9113), .Z(n9087) );
  AND U8937 ( .A(n9114), .B(n9115), .Z(n9113) );
  XNOR U8938 ( .A(n9112), .B(n9103), .Z(n9115) );
  IV U8939 ( .A(n9057), .Z(n9103) );
  XNOR U8940 ( .A(n9116), .B(n9096), .Z(n9057) );
  XNOR U8941 ( .A(n9117), .B(n9102), .Z(n9096) );
  XOR U8942 ( .A(n9118), .B(n9119), .Z(n9102) );
  NOR U8943 ( .A(n9120), .B(n9121), .Z(n9119) );
  XNOR U8944 ( .A(n9118), .B(n9122), .Z(n9120) );
  XNOR U8945 ( .A(n9101), .B(n9093), .Z(n9117) );
  XOR U8946 ( .A(n9123), .B(n9124), .Z(n9093) );
  AND U8947 ( .A(n9125), .B(n9126), .Z(n9124) );
  XNOR U8948 ( .A(n9123), .B(n9127), .Z(n9125) );
  XNOR U8949 ( .A(n9128), .B(n9098), .Z(n9101) );
  XOR U8950 ( .A(n9129), .B(n9130), .Z(n9098) );
  AND U8951 ( .A(n9131), .B(n9132), .Z(n9130) );
  XOR U8952 ( .A(n9129), .B(n9133), .Z(n9131) );
  XNOR U8953 ( .A(n9134), .B(n9135), .Z(n9128) );
  NOR U8954 ( .A(n9136), .B(n9137), .Z(n9135) );
  XOR U8955 ( .A(n9134), .B(n9138), .Z(n9136) );
  XNOR U8956 ( .A(n9097), .B(n9104), .Z(n9116) );
  NOR U8957 ( .A(n9065), .B(n9139), .Z(n9104) );
  XOR U8958 ( .A(n9109), .B(n9108), .Z(n9097) );
  XNOR U8959 ( .A(n9140), .B(n9105), .Z(n9108) );
  XOR U8960 ( .A(n9141), .B(n9142), .Z(n9105) );
  AND U8961 ( .A(n9143), .B(n9144), .Z(n9142) );
  XOR U8962 ( .A(n9141), .B(n9145), .Z(n9143) );
  XNOR U8963 ( .A(n9146), .B(n9147), .Z(n9140) );
  NOR U8964 ( .A(n9148), .B(n9149), .Z(n9147) );
  XNOR U8965 ( .A(n9146), .B(n9150), .Z(n9148) );
  XOR U8966 ( .A(n9151), .B(n9152), .Z(n9109) );
  NOR U8967 ( .A(n9153), .B(n9154), .Z(n9152) );
  XNOR U8968 ( .A(n9151), .B(n9155), .Z(n9153) );
  XNOR U8969 ( .A(n9054), .B(n9112), .Z(n9114) );
  XNOR U8970 ( .A(n9156), .B(n9157), .Z(n9054) );
  AND U8971 ( .A(n94), .B(n9061), .Z(n9157) );
  XOR U8972 ( .A(n9156), .B(n9059), .Z(n9061) );
  AND U8973 ( .A(n9062), .B(n9065), .Z(n9112) );
  XOR U8974 ( .A(n9158), .B(n9139), .Z(n9065) );
  XNOR U8975 ( .A(p_input[1024]), .B(p_input[80]), .Z(n9139) );
  XOR U8976 ( .A(n9127), .B(n9126), .Z(n9158) );
  XNOR U8977 ( .A(n9159), .B(n9133), .Z(n9126) );
  XNOR U8978 ( .A(n9122), .B(n9121), .Z(n9133) );
  XOR U8979 ( .A(n9160), .B(n9118), .Z(n9121) );
  XOR U8980 ( .A(p_input[1034]), .B(p_input[90]), .Z(n9118) );
  XNOR U8981 ( .A(p_input[1035]), .B(p_input[91]), .Z(n9160) );
  XOR U8982 ( .A(p_input[1036]), .B(p_input[92]), .Z(n9122) );
  XNOR U8983 ( .A(n9132), .B(n9123), .Z(n9159) );
  XOR U8984 ( .A(p_input[1025]), .B(p_input[81]), .Z(n9123) );
  XOR U8985 ( .A(n9161), .B(n9138), .Z(n9132) );
  XNOR U8986 ( .A(p_input[1039]), .B(p_input[95]), .Z(n9138) );
  XOR U8987 ( .A(n9129), .B(n9137), .Z(n9161) );
  XOR U8988 ( .A(n9162), .B(n9134), .Z(n9137) );
  XOR U8989 ( .A(p_input[1037]), .B(p_input[93]), .Z(n9134) );
  XNOR U8990 ( .A(p_input[1038]), .B(p_input[94]), .Z(n9162) );
  XOR U8991 ( .A(p_input[1033]), .B(p_input[89]), .Z(n9129) );
  XNOR U8992 ( .A(n9145), .B(n9144), .Z(n9127) );
  XNOR U8993 ( .A(n9163), .B(n9150), .Z(n9144) );
  XOR U8994 ( .A(p_input[1032]), .B(p_input[88]), .Z(n9150) );
  XOR U8995 ( .A(n9141), .B(n9149), .Z(n9163) );
  XOR U8996 ( .A(n9164), .B(n9146), .Z(n9149) );
  XOR U8997 ( .A(p_input[1030]), .B(p_input[86]), .Z(n9146) );
  XNOR U8998 ( .A(p_input[1031]), .B(p_input[87]), .Z(n9164) );
  XOR U8999 ( .A(p_input[1026]), .B(p_input[82]), .Z(n9141) );
  XNOR U9000 ( .A(n9155), .B(n9154), .Z(n9145) );
  XOR U9001 ( .A(n9165), .B(n9151), .Z(n9154) );
  XOR U9002 ( .A(p_input[1027]), .B(p_input[83]), .Z(n9151) );
  XNOR U9003 ( .A(p_input[1028]), .B(p_input[84]), .Z(n9165) );
  XOR U9004 ( .A(p_input[1029]), .B(p_input[85]), .Z(n9155) );
  XNOR U9005 ( .A(n9166), .B(n9167), .Z(n9062) );
  AND U9006 ( .A(n94), .B(n9168), .Z(n9167) );
  XNOR U9007 ( .A(n9169), .B(n9170), .Z(n94) );
  AND U9008 ( .A(n9171), .B(n9172), .Z(n9170) );
  XOR U9009 ( .A(n9169), .B(n9072), .Z(n9172) );
  XNOR U9010 ( .A(n9169), .B(n9026), .Z(n9171) );
  XOR U9011 ( .A(n9173), .B(n9174), .Z(n9169) );
  AND U9012 ( .A(n9175), .B(n9176), .Z(n9174) );
  XOR U9013 ( .A(n9173), .B(n9036), .Z(n9175) );
  XOR U9014 ( .A(n9177), .B(n9178), .Z(n9015) );
  AND U9015 ( .A(n98), .B(n9168), .Z(n9178) );
  XNOR U9016 ( .A(n9166), .B(n9177), .Z(n9168) );
  XNOR U9017 ( .A(n9179), .B(n9180), .Z(n98) );
  AND U9018 ( .A(n9181), .B(n9182), .Z(n9180) );
  XNOR U9019 ( .A(n9183), .B(n9179), .Z(n9182) );
  IV U9020 ( .A(n9072), .Z(n9183) );
  XNOR U9021 ( .A(n9184), .B(n9185), .Z(n9072) );
  AND U9022 ( .A(n101), .B(n9186), .Z(n9185) );
  XNOR U9023 ( .A(n9184), .B(n9187), .Z(n9186) );
  XNOR U9024 ( .A(n9026), .B(n9179), .Z(n9181) );
  XOR U9025 ( .A(n9188), .B(n9189), .Z(n9026) );
  AND U9026 ( .A(n109), .B(n9190), .Z(n9189) );
  XOR U9027 ( .A(n9173), .B(n9191), .Z(n9179) );
  AND U9028 ( .A(n9192), .B(n9176), .Z(n9191) );
  XNOR U9029 ( .A(n9085), .B(n9173), .Z(n9176) );
  XNOR U9030 ( .A(n9193), .B(n9194), .Z(n9085) );
  AND U9031 ( .A(n101), .B(n9195), .Z(n9194) );
  XOR U9032 ( .A(n9196), .B(n9193), .Z(n9195) );
  XNOR U9033 ( .A(n9197), .B(n9173), .Z(n9192) );
  IV U9034 ( .A(n9036), .Z(n9197) );
  XOR U9035 ( .A(n9198), .B(n9199), .Z(n9036) );
  AND U9036 ( .A(n109), .B(n9200), .Z(n9199) );
  XOR U9037 ( .A(n9201), .B(n9202), .Z(n9173) );
  AND U9038 ( .A(n9203), .B(n9204), .Z(n9202) );
  XNOR U9039 ( .A(n9110), .B(n9201), .Z(n9204) );
  XNOR U9040 ( .A(n9205), .B(n9206), .Z(n9110) );
  AND U9041 ( .A(n101), .B(n9207), .Z(n9206) );
  XNOR U9042 ( .A(n9208), .B(n9205), .Z(n9207) );
  XOR U9043 ( .A(n9201), .B(n9047), .Z(n9203) );
  XOR U9044 ( .A(n9209), .B(n9210), .Z(n9047) );
  AND U9045 ( .A(n109), .B(n9211), .Z(n9210) );
  XOR U9046 ( .A(n9212), .B(n9213), .Z(n9201) );
  AND U9047 ( .A(n9214), .B(n9215), .Z(n9213) );
  XNOR U9048 ( .A(n9212), .B(n9156), .Z(n9215) );
  XNOR U9049 ( .A(n9216), .B(n9217), .Z(n9156) );
  AND U9050 ( .A(n101), .B(n9218), .Z(n9217) );
  XOR U9051 ( .A(n9219), .B(n9216), .Z(n9218) );
  XNOR U9052 ( .A(n9220), .B(n9212), .Z(n9214) );
  IV U9053 ( .A(n9059), .Z(n9220) );
  XOR U9054 ( .A(n9221), .B(n9222), .Z(n9059) );
  AND U9055 ( .A(n109), .B(n9223), .Z(n9222) );
  AND U9056 ( .A(n9177), .B(n9166), .Z(n9212) );
  XNOR U9057 ( .A(n9224), .B(n9225), .Z(n9166) );
  AND U9058 ( .A(n101), .B(n9226), .Z(n9225) );
  XNOR U9059 ( .A(n9227), .B(n9224), .Z(n9226) );
  XNOR U9060 ( .A(n9228), .B(n9229), .Z(n101) );
  AND U9061 ( .A(n9230), .B(n9231), .Z(n9229) );
  XOR U9062 ( .A(n9187), .B(n9228), .Z(n9231) );
  AND U9063 ( .A(n9232), .B(n9233), .Z(n9187) );
  XOR U9064 ( .A(n9228), .B(n9184), .Z(n9230) );
  XNOR U9065 ( .A(n9234), .B(n9235), .Z(n9184) );
  AND U9066 ( .A(n105), .B(n9190), .Z(n9235) );
  XOR U9067 ( .A(n9188), .B(n9234), .Z(n9190) );
  XOR U9068 ( .A(n9236), .B(n9237), .Z(n9228) );
  AND U9069 ( .A(n9238), .B(n9239), .Z(n9237) );
  XNOR U9070 ( .A(n9236), .B(n9232), .Z(n9239) );
  IV U9071 ( .A(n9196), .Z(n9232) );
  XOR U9072 ( .A(n9240), .B(n9241), .Z(n9196) );
  XOR U9073 ( .A(n9242), .B(n9233), .Z(n9241) );
  AND U9074 ( .A(n9208), .B(n9243), .Z(n9233) );
  AND U9075 ( .A(n9244), .B(n9245), .Z(n9242) );
  XOR U9076 ( .A(n9246), .B(n9240), .Z(n9244) );
  XNOR U9077 ( .A(n9193), .B(n9236), .Z(n9238) );
  XNOR U9078 ( .A(n9247), .B(n9248), .Z(n9193) );
  AND U9079 ( .A(n105), .B(n9200), .Z(n9248) );
  XOR U9080 ( .A(n9247), .B(n9198), .Z(n9200) );
  XOR U9081 ( .A(n9249), .B(n9250), .Z(n9236) );
  AND U9082 ( .A(n9251), .B(n9252), .Z(n9250) );
  XNOR U9083 ( .A(n9249), .B(n9208), .Z(n9252) );
  XOR U9084 ( .A(n9253), .B(n9245), .Z(n9208) );
  XNOR U9085 ( .A(n9254), .B(n9240), .Z(n9245) );
  XOR U9086 ( .A(n9255), .B(n9256), .Z(n9240) );
  AND U9087 ( .A(n9257), .B(n9258), .Z(n9256) );
  XOR U9088 ( .A(n9259), .B(n9255), .Z(n9257) );
  XNOR U9089 ( .A(n9260), .B(n9261), .Z(n9254) );
  AND U9090 ( .A(n9262), .B(n9263), .Z(n9261) );
  XOR U9091 ( .A(n9260), .B(n9264), .Z(n9262) );
  XNOR U9092 ( .A(n9246), .B(n9243), .Z(n9253) );
  AND U9093 ( .A(n9265), .B(n9266), .Z(n9243) );
  XOR U9094 ( .A(n9267), .B(n9268), .Z(n9246) );
  AND U9095 ( .A(n9269), .B(n9270), .Z(n9268) );
  XOR U9096 ( .A(n9267), .B(n9271), .Z(n9269) );
  XNOR U9097 ( .A(n9205), .B(n9249), .Z(n9251) );
  XNOR U9098 ( .A(n9272), .B(n9273), .Z(n9205) );
  AND U9099 ( .A(n105), .B(n9211), .Z(n9273) );
  XOR U9100 ( .A(n9272), .B(n9209), .Z(n9211) );
  XOR U9101 ( .A(n9274), .B(n9275), .Z(n9249) );
  AND U9102 ( .A(n9276), .B(n9277), .Z(n9275) );
  XNOR U9103 ( .A(n9274), .B(n9265), .Z(n9277) );
  IV U9104 ( .A(n9219), .Z(n9265) );
  XNOR U9105 ( .A(n9278), .B(n9258), .Z(n9219) );
  XNOR U9106 ( .A(n9279), .B(n9264), .Z(n9258) );
  XOR U9107 ( .A(n9280), .B(n9281), .Z(n9264) );
  NOR U9108 ( .A(n9282), .B(n9283), .Z(n9281) );
  XNOR U9109 ( .A(n9280), .B(n9284), .Z(n9282) );
  XNOR U9110 ( .A(n9263), .B(n9255), .Z(n9279) );
  XOR U9111 ( .A(n9285), .B(n9286), .Z(n9255) );
  AND U9112 ( .A(n9287), .B(n9288), .Z(n9286) );
  XNOR U9113 ( .A(n9285), .B(n9289), .Z(n9287) );
  XNOR U9114 ( .A(n9290), .B(n9260), .Z(n9263) );
  XOR U9115 ( .A(n9291), .B(n9292), .Z(n9260) );
  AND U9116 ( .A(n9293), .B(n9294), .Z(n9292) );
  XOR U9117 ( .A(n9291), .B(n9295), .Z(n9293) );
  XNOR U9118 ( .A(n9296), .B(n9297), .Z(n9290) );
  NOR U9119 ( .A(n9298), .B(n9299), .Z(n9297) );
  XOR U9120 ( .A(n9296), .B(n9300), .Z(n9298) );
  XNOR U9121 ( .A(n9259), .B(n9266), .Z(n9278) );
  NOR U9122 ( .A(n9227), .B(n9301), .Z(n9266) );
  XOR U9123 ( .A(n9271), .B(n9270), .Z(n9259) );
  XNOR U9124 ( .A(n9302), .B(n9267), .Z(n9270) );
  XOR U9125 ( .A(n9303), .B(n9304), .Z(n9267) );
  AND U9126 ( .A(n9305), .B(n9306), .Z(n9304) );
  XOR U9127 ( .A(n9303), .B(n9307), .Z(n9305) );
  XNOR U9128 ( .A(n9308), .B(n9309), .Z(n9302) );
  NOR U9129 ( .A(n9310), .B(n9311), .Z(n9309) );
  XNOR U9130 ( .A(n9308), .B(n9312), .Z(n9310) );
  XOR U9131 ( .A(n9313), .B(n9314), .Z(n9271) );
  NOR U9132 ( .A(n9315), .B(n9316), .Z(n9314) );
  XNOR U9133 ( .A(n9313), .B(n9317), .Z(n9315) );
  XNOR U9134 ( .A(n9216), .B(n9274), .Z(n9276) );
  XNOR U9135 ( .A(n9318), .B(n9319), .Z(n9216) );
  AND U9136 ( .A(n105), .B(n9223), .Z(n9319) );
  XOR U9137 ( .A(n9318), .B(n9221), .Z(n9223) );
  AND U9138 ( .A(n9224), .B(n9227), .Z(n9274) );
  XOR U9139 ( .A(n9320), .B(n9301), .Z(n9227) );
  XNOR U9140 ( .A(p_input[1024]), .B(p_input[96]), .Z(n9301) );
  XOR U9141 ( .A(n9289), .B(n9288), .Z(n9320) );
  XNOR U9142 ( .A(n9321), .B(n9295), .Z(n9288) );
  XNOR U9143 ( .A(n9284), .B(n9283), .Z(n9295) );
  XOR U9144 ( .A(n9322), .B(n9280), .Z(n9283) );
  XOR U9145 ( .A(p_input[1034]), .B(p_input[106]), .Z(n9280) );
  XNOR U9146 ( .A(p_input[1035]), .B(p_input[107]), .Z(n9322) );
  XOR U9147 ( .A(p_input[1036]), .B(p_input[108]), .Z(n9284) );
  XNOR U9148 ( .A(n9294), .B(n9285), .Z(n9321) );
  XOR U9149 ( .A(p_input[1025]), .B(p_input[97]), .Z(n9285) );
  XOR U9150 ( .A(n9323), .B(n9300), .Z(n9294) );
  XNOR U9151 ( .A(p_input[1039]), .B(p_input[111]), .Z(n9300) );
  XOR U9152 ( .A(n9291), .B(n9299), .Z(n9323) );
  XOR U9153 ( .A(n9324), .B(n9296), .Z(n9299) );
  XOR U9154 ( .A(p_input[1037]), .B(p_input[109]), .Z(n9296) );
  XNOR U9155 ( .A(p_input[1038]), .B(p_input[110]), .Z(n9324) );
  XOR U9156 ( .A(p_input[1033]), .B(p_input[105]), .Z(n9291) );
  XNOR U9157 ( .A(n9307), .B(n9306), .Z(n9289) );
  XNOR U9158 ( .A(n9325), .B(n9312), .Z(n9306) );
  XOR U9159 ( .A(p_input[1032]), .B(p_input[104]), .Z(n9312) );
  XOR U9160 ( .A(n9303), .B(n9311), .Z(n9325) );
  XOR U9161 ( .A(n9326), .B(n9308), .Z(n9311) );
  XOR U9162 ( .A(p_input[102]), .B(p_input[1030]), .Z(n9308) );
  XNOR U9163 ( .A(p_input[1031]), .B(p_input[103]), .Z(n9326) );
  XOR U9164 ( .A(p_input[1026]), .B(p_input[98]), .Z(n9303) );
  XNOR U9165 ( .A(n9317), .B(n9316), .Z(n9307) );
  XOR U9166 ( .A(n9327), .B(n9313), .Z(n9316) );
  XOR U9167 ( .A(p_input[1027]), .B(p_input[99]), .Z(n9313) );
  XOR U9168 ( .A(p_input[100]), .B(n9328), .Z(n9327) );
  XOR U9169 ( .A(p_input[101]), .B(p_input[1029]), .Z(n9317) );
  XNOR U9170 ( .A(n9329), .B(n9330), .Z(n9224) );
  AND U9171 ( .A(n105), .B(n9331), .Z(n9330) );
  XNOR U9172 ( .A(n9332), .B(n9333), .Z(n105) );
  AND U9173 ( .A(n9334), .B(n9335), .Z(n9333) );
  XOR U9174 ( .A(n9332), .B(n9234), .Z(n9335) );
  XNOR U9175 ( .A(n9332), .B(n9188), .Z(n9334) );
  XOR U9176 ( .A(n9336), .B(n9337), .Z(n9332) );
  AND U9177 ( .A(n9338), .B(n9339), .Z(n9337) );
  XOR U9178 ( .A(n9336), .B(n9198), .Z(n9338) );
  XOR U9179 ( .A(n9340), .B(n9341), .Z(n9177) );
  AND U9180 ( .A(n109), .B(n9331), .Z(n9341) );
  XNOR U9181 ( .A(n9329), .B(n9340), .Z(n9331) );
  XNOR U9182 ( .A(n9342), .B(n9343), .Z(n109) );
  AND U9183 ( .A(n9344), .B(n9345), .Z(n9343) );
  XNOR U9184 ( .A(n9346), .B(n9342), .Z(n9345) );
  IV U9185 ( .A(n9234), .Z(n9346) );
  XNOR U9186 ( .A(n9347), .B(n9348), .Z(n9234) );
  AND U9187 ( .A(n112), .B(n9349), .Z(n9348) );
  XNOR U9188 ( .A(n9347), .B(n9350), .Z(n9349) );
  XNOR U9189 ( .A(n9188), .B(n9342), .Z(n9344) );
  XOR U9190 ( .A(n9351), .B(n9352), .Z(n9188) );
  AND U9191 ( .A(n120), .B(n9353), .Z(n9352) );
  XOR U9192 ( .A(n9336), .B(n9354), .Z(n9342) );
  AND U9193 ( .A(n9355), .B(n9339), .Z(n9354) );
  XNOR U9194 ( .A(n9247), .B(n9336), .Z(n9339) );
  XNOR U9195 ( .A(n9356), .B(n9357), .Z(n9247) );
  AND U9196 ( .A(n112), .B(n9358), .Z(n9357) );
  XOR U9197 ( .A(n9359), .B(n9356), .Z(n9358) );
  XNOR U9198 ( .A(n9360), .B(n9336), .Z(n9355) );
  IV U9199 ( .A(n9198), .Z(n9360) );
  XOR U9200 ( .A(n9361), .B(n9362), .Z(n9198) );
  AND U9201 ( .A(n120), .B(n9363), .Z(n9362) );
  XOR U9202 ( .A(n9364), .B(n9365), .Z(n9336) );
  AND U9203 ( .A(n9366), .B(n9367), .Z(n9365) );
  XNOR U9204 ( .A(n9272), .B(n9364), .Z(n9367) );
  XNOR U9205 ( .A(n9368), .B(n9369), .Z(n9272) );
  AND U9206 ( .A(n112), .B(n9370), .Z(n9369) );
  XNOR U9207 ( .A(n9371), .B(n9368), .Z(n9370) );
  XOR U9208 ( .A(n9364), .B(n9209), .Z(n9366) );
  XOR U9209 ( .A(n9372), .B(n9373), .Z(n9209) );
  AND U9210 ( .A(n120), .B(n9374), .Z(n9373) );
  XOR U9211 ( .A(n9375), .B(n9376), .Z(n9364) );
  AND U9212 ( .A(n9377), .B(n9378), .Z(n9376) );
  XNOR U9213 ( .A(n9375), .B(n9318), .Z(n9378) );
  XNOR U9214 ( .A(n9379), .B(n9380), .Z(n9318) );
  AND U9215 ( .A(n112), .B(n9381), .Z(n9380) );
  XOR U9216 ( .A(n9382), .B(n9379), .Z(n9381) );
  XNOR U9217 ( .A(n9383), .B(n9375), .Z(n9377) );
  IV U9218 ( .A(n9221), .Z(n9383) );
  XOR U9219 ( .A(n9384), .B(n9385), .Z(n9221) );
  AND U9220 ( .A(n120), .B(n9386), .Z(n9385) );
  AND U9221 ( .A(n9340), .B(n9329), .Z(n9375) );
  XNOR U9222 ( .A(n9387), .B(n9388), .Z(n9329) );
  AND U9223 ( .A(n112), .B(n9389), .Z(n9388) );
  XNOR U9224 ( .A(n9390), .B(n9387), .Z(n9389) );
  XNOR U9225 ( .A(n9391), .B(n9392), .Z(n112) );
  AND U9226 ( .A(n9393), .B(n9394), .Z(n9392) );
  XOR U9227 ( .A(n9350), .B(n9391), .Z(n9394) );
  AND U9228 ( .A(n9395), .B(n9396), .Z(n9350) );
  XOR U9229 ( .A(n9391), .B(n9347), .Z(n9393) );
  XNOR U9230 ( .A(n9397), .B(n9398), .Z(n9347) );
  AND U9231 ( .A(n116), .B(n9353), .Z(n9398) );
  XOR U9232 ( .A(n9351), .B(n9397), .Z(n9353) );
  XOR U9233 ( .A(n9399), .B(n9400), .Z(n9391) );
  AND U9234 ( .A(n9401), .B(n9402), .Z(n9400) );
  XNOR U9235 ( .A(n9399), .B(n9395), .Z(n9402) );
  IV U9236 ( .A(n9359), .Z(n9395) );
  XOR U9237 ( .A(n9403), .B(n9404), .Z(n9359) );
  XOR U9238 ( .A(n9405), .B(n9396), .Z(n9404) );
  AND U9239 ( .A(n9371), .B(n9406), .Z(n9396) );
  AND U9240 ( .A(n9407), .B(n9408), .Z(n9405) );
  XOR U9241 ( .A(n9409), .B(n9403), .Z(n9407) );
  XNOR U9242 ( .A(n9356), .B(n9399), .Z(n9401) );
  XNOR U9243 ( .A(n9410), .B(n9411), .Z(n9356) );
  AND U9244 ( .A(n116), .B(n9363), .Z(n9411) );
  XOR U9245 ( .A(n9410), .B(n9361), .Z(n9363) );
  XOR U9246 ( .A(n9412), .B(n9413), .Z(n9399) );
  AND U9247 ( .A(n9414), .B(n9415), .Z(n9413) );
  XNOR U9248 ( .A(n9412), .B(n9371), .Z(n9415) );
  XOR U9249 ( .A(n9416), .B(n9408), .Z(n9371) );
  XNOR U9250 ( .A(n9417), .B(n9403), .Z(n9408) );
  XOR U9251 ( .A(n9418), .B(n9419), .Z(n9403) );
  AND U9252 ( .A(n9420), .B(n9421), .Z(n9419) );
  XOR U9253 ( .A(n9422), .B(n9418), .Z(n9420) );
  XNOR U9254 ( .A(n9423), .B(n9424), .Z(n9417) );
  AND U9255 ( .A(n9425), .B(n9426), .Z(n9424) );
  XOR U9256 ( .A(n9423), .B(n9427), .Z(n9425) );
  XNOR U9257 ( .A(n9409), .B(n9406), .Z(n9416) );
  AND U9258 ( .A(n9428), .B(n9429), .Z(n9406) );
  XOR U9259 ( .A(n9430), .B(n9431), .Z(n9409) );
  AND U9260 ( .A(n9432), .B(n9433), .Z(n9431) );
  XOR U9261 ( .A(n9430), .B(n9434), .Z(n9432) );
  XNOR U9262 ( .A(n9368), .B(n9412), .Z(n9414) );
  XNOR U9263 ( .A(n9435), .B(n9436), .Z(n9368) );
  AND U9264 ( .A(n116), .B(n9374), .Z(n9436) );
  XOR U9265 ( .A(n9435), .B(n9372), .Z(n9374) );
  XOR U9266 ( .A(n9437), .B(n9438), .Z(n9412) );
  AND U9267 ( .A(n9439), .B(n9440), .Z(n9438) );
  XNOR U9268 ( .A(n9437), .B(n9428), .Z(n9440) );
  IV U9269 ( .A(n9382), .Z(n9428) );
  XNOR U9270 ( .A(n9441), .B(n9421), .Z(n9382) );
  XNOR U9271 ( .A(n9442), .B(n9427), .Z(n9421) );
  XOR U9272 ( .A(n9443), .B(n9444), .Z(n9427) );
  NOR U9273 ( .A(n9445), .B(n9446), .Z(n9444) );
  XNOR U9274 ( .A(n9443), .B(n9447), .Z(n9445) );
  XNOR U9275 ( .A(n9426), .B(n9418), .Z(n9442) );
  XOR U9276 ( .A(n9448), .B(n9449), .Z(n9418) );
  AND U9277 ( .A(n9450), .B(n9451), .Z(n9449) );
  XNOR U9278 ( .A(n9448), .B(n9452), .Z(n9450) );
  XNOR U9279 ( .A(n9453), .B(n9423), .Z(n9426) );
  XOR U9280 ( .A(n9454), .B(n9455), .Z(n9423) );
  AND U9281 ( .A(n9456), .B(n9457), .Z(n9455) );
  XOR U9282 ( .A(n9454), .B(n9458), .Z(n9456) );
  XNOR U9283 ( .A(n9459), .B(n9460), .Z(n9453) );
  NOR U9284 ( .A(n9461), .B(n9462), .Z(n9460) );
  XOR U9285 ( .A(n9459), .B(n9463), .Z(n9461) );
  XNOR U9286 ( .A(n9422), .B(n9429), .Z(n9441) );
  NOR U9287 ( .A(n9390), .B(n9464), .Z(n9429) );
  XOR U9288 ( .A(n9434), .B(n9433), .Z(n9422) );
  XNOR U9289 ( .A(n9465), .B(n9430), .Z(n9433) );
  XOR U9290 ( .A(n9466), .B(n9467), .Z(n9430) );
  AND U9291 ( .A(n9468), .B(n9469), .Z(n9467) );
  XOR U9292 ( .A(n9466), .B(n9470), .Z(n9468) );
  XNOR U9293 ( .A(n9471), .B(n9472), .Z(n9465) );
  NOR U9294 ( .A(n9473), .B(n9474), .Z(n9472) );
  XNOR U9295 ( .A(n9471), .B(n9475), .Z(n9473) );
  XOR U9296 ( .A(n9476), .B(n9477), .Z(n9434) );
  NOR U9297 ( .A(n9478), .B(n9479), .Z(n9477) );
  XNOR U9298 ( .A(n9476), .B(n9480), .Z(n9478) );
  XNOR U9299 ( .A(n9379), .B(n9437), .Z(n9439) );
  XNOR U9300 ( .A(n9481), .B(n9482), .Z(n9379) );
  AND U9301 ( .A(n116), .B(n9386), .Z(n9482) );
  XOR U9302 ( .A(n9481), .B(n9384), .Z(n9386) );
  AND U9303 ( .A(n9387), .B(n9390), .Z(n9437) );
  XOR U9304 ( .A(n9483), .B(n9464), .Z(n9390) );
  XNOR U9305 ( .A(p_input[1024]), .B(p_input[112]), .Z(n9464) );
  XOR U9306 ( .A(n9452), .B(n9451), .Z(n9483) );
  XNOR U9307 ( .A(n9484), .B(n9458), .Z(n9451) );
  XNOR U9308 ( .A(n9447), .B(n9446), .Z(n9458) );
  XOR U9309 ( .A(n9485), .B(n9443), .Z(n9446) );
  XOR U9310 ( .A(p_input[1034]), .B(p_input[122]), .Z(n9443) );
  XNOR U9311 ( .A(p_input[1035]), .B(p_input[123]), .Z(n9485) );
  XOR U9312 ( .A(p_input[1036]), .B(p_input[124]), .Z(n9447) );
  XNOR U9313 ( .A(n9457), .B(n9448), .Z(n9484) );
  XOR U9314 ( .A(p_input[1025]), .B(p_input[113]), .Z(n9448) );
  XOR U9315 ( .A(n9486), .B(n9463), .Z(n9457) );
  XNOR U9316 ( .A(p_input[1039]), .B(p_input[127]), .Z(n9463) );
  XOR U9317 ( .A(n9454), .B(n9462), .Z(n9486) );
  XOR U9318 ( .A(n9487), .B(n9459), .Z(n9462) );
  XOR U9319 ( .A(p_input[1037]), .B(p_input[125]), .Z(n9459) );
  XNOR U9320 ( .A(p_input[1038]), .B(p_input[126]), .Z(n9487) );
  XOR U9321 ( .A(p_input[1033]), .B(p_input[121]), .Z(n9454) );
  XNOR U9322 ( .A(n9470), .B(n9469), .Z(n9452) );
  XNOR U9323 ( .A(n9488), .B(n9475), .Z(n9469) );
  XOR U9324 ( .A(p_input[1032]), .B(p_input[120]), .Z(n9475) );
  XOR U9325 ( .A(n9466), .B(n9474), .Z(n9488) );
  XOR U9326 ( .A(n9489), .B(n9471), .Z(n9474) );
  XOR U9327 ( .A(p_input[1030]), .B(p_input[118]), .Z(n9471) );
  XNOR U9328 ( .A(p_input[1031]), .B(p_input[119]), .Z(n9489) );
  XOR U9329 ( .A(p_input[1026]), .B(p_input[114]), .Z(n9466) );
  XNOR U9330 ( .A(n9480), .B(n9479), .Z(n9470) );
  XOR U9331 ( .A(n9490), .B(n9476), .Z(n9479) );
  XOR U9332 ( .A(p_input[1027]), .B(p_input[115]), .Z(n9476) );
  XNOR U9333 ( .A(p_input[1028]), .B(p_input[116]), .Z(n9490) );
  XOR U9334 ( .A(p_input[1029]), .B(p_input[117]), .Z(n9480) );
  XNOR U9335 ( .A(n9491), .B(n9492), .Z(n9387) );
  AND U9336 ( .A(n116), .B(n9493), .Z(n9492) );
  XNOR U9337 ( .A(n9494), .B(n9495), .Z(n116) );
  AND U9338 ( .A(n9496), .B(n9497), .Z(n9495) );
  XOR U9339 ( .A(n9494), .B(n9397), .Z(n9497) );
  XNOR U9340 ( .A(n9494), .B(n9351), .Z(n9496) );
  XOR U9341 ( .A(n9498), .B(n9499), .Z(n9494) );
  AND U9342 ( .A(n9500), .B(n9501), .Z(n9499) );
  XOR U9343 ( .A(n9498), .B(n9361), .Z(n9500) );
  XOR U9344 ( .A(n9502), .B(n9503), .Z(n9340) );
  AND U9345 ( .A(n120), .B(n9493), .Z(n9503) );
  XNOR U9346 ( .A(n9491), .B(n9502), .Z(n9493) );
  XNOR U9347 ( .A(n9504), .B(n9505), .Z(n120) );
  AND U9348 ( .A(n9506), .B(n9507), .Z(n9505) );
  XNOR U9349 ( .A(n9508), .B(n9504), .Z(n9507) );
  IV U9350 ( .A(n9397), .Z(n9508) );
  XNOR U9351 ( .A(n9509), .B(n9510), .Z(n9397) );
  AND U9352 ( .A(n123), .B(n9511), .Z(n9510) );
  XNOR U9353 ( .A(n9509), .B(n9512), .Z(n9511) );
  XNOR U9354 ( .A(n9351), .B(n9504), .Z(n9506) );
  XOR U9355 ( .A(n9513), .B(n9514), .Z(n9351) );
  AND U9356 ( .A(n131), .B(n9515), .Z(n9514) );
  XOR U9357 ( .A(n9498), .B(n9516), .Z(n9504) );
  AND U9358 ( .A(n9517), .B(n9501), .Z(n9516) );
  XNOR U9359 ( .A(n9410), .B(n9498), .Z(n9501) );
  XNOR U9360 ( .A(n9518), .B(n9519), .Z(n9410) );
  AND U9361 ( .A(n123), .B(n9520), .Z(n9519) );
  XOR U9362 ( .A(n9521), .B(n9518), .Z(n9520) );
  XNOR U9363 ( .A(n9522), .B(n9498), .Z(n9517) );
  IV U9364 ( .A(n9361), .Z(n9522) );
  XOR U9365 ( .A(n9523), .B(n9524), .Z(n9361) );
  AND U9366 ( .A(n131), .B(n9525), .Z(n9524) );
  XOR U9367 ( .A(n9526), .B(n9527), .Z(n9498) );
  AND U9368 ( .A(n9528), .B(n9529), .Z(n9527) );
  XNOR U9369 ( .A(n9435), .B(n9526), .Z(n9529) );
  XNOR U9370 ( .A(n9530), .B(n9531), .Z(n9435) );
  AND U9371 ( .A(n123), .B(n9532), .Z(n9531) );
  XNOR U9372 ( .A(n9533), .B(n9530), .Z(n9532) );
  XOR U9373 ( .A(n9526), .B(n9372), .Z(n9528) );
  XOR U9374 ( .A(n9534), .B(n9535), .Z(n9372) );
  AND U9375 ( .A(n131), .B(n9536), .Z(n9535) );
  XOR U9376 ( .A(n9537), .B(n9538), .Z(n9526) );
  AND U9377 ( .A(n9539), .B(n9540), .Z(n9538) );
  XNOR U9378 ( .A(n9537), .B(n9481), .Z(n9540) );
  XNOR U9379 ( .A(n9541), .B(n9542), .Z(n9481) );
  AND U9380 ( .A(n123), .B(n9543), .Z(n9542) );
  XOR U9381 ( .A(n9544), .B(n9541), .Z(n9543) );
  XNOR U9382 ( .A(n9545), .B(n9537), .Z(n9539) );
  IV U9383 ( .A(n9384), .Z(n9545) );
  XOR U9384 ( .A(n9546), .B(n9547), .Z(n9384) );
  AND U9385 ( .A(n131), .B(n9548), .Z(n9547) );
  AND U9386 ( .A(n9502), .B(n9491), .Z(n9537) );
  XNOR U9387 ( .A(n9549), .B(n9550), .Z(n9491) );
  AND U9388 ( .A(n123), .B(n9551), .Z(n9550) );
  XNOR U9389 ( .A(n9552), .B(n9549), .Z(n9551) );
  XNOR U9390 ( .A(n9553), .B(n9554), .Z(n123) );
  AND U9391 ( .A(n9555), .B(n9556), .Z(n9554) );
  XOR U9392 ( .A(n9512), .B(n9553), .Z(n9556) );
  AND U9393 ( .A(n9557), .B(n9558), .Z(n9512) );
  XOR U9394 ( .A(n9553), .B(n9509), .Z(n9555) );
  XNOR U9395 ( .A(n9559), .B(n9560), .Z(n9509) );
  AND U9396 ( .A(n127), .B(n9515), .Z(n9560) );
  XOR U9397 ( .A(n9513), .B(n9559), .Z(n9515) );
  XOR U9398 ( .A(n9561), .B(n9562), .Z(n9553) );
  AND U9399 ( .A(n9563), .B(n9564), .Z(n9562) );
  XNOR U9400 ( .A(n9561), .B(n9557), .Z(n9564) );
  IV U9401 ( .A(n9521), .Z(n9557) );
  XOR U9402 ( .A(n9565), .B(n9566), .Z(n9521) );
  XOR U9403 ( .A(n9567), .B(n9558), .Z(n9566) );
  AND U9404 ( .A(n9533), .B(n9568), .Z(n9558) );
  AND U9405 ( .A(n9569), .B(n9570), .Z(n9567) );
  XOR U9406 ( .A(n9571), .B(n9565), .Z(n9569) );
  XNOR U9407 ( .A(n9518), .B(n9561), .Z(n9563) );
  XNOR U9408 ( .A(n9572), .B(n9573), .Z(n9518) );
  AND U9409 ( .A(n127), .B(n9525), .Z(n9573) );
  XOR U9410 ( .A(n9572), .B(n9523), .Z(n9525) );
  XOR U9411 ( .A(n9574), .B(n9575), .Z(n9561) );
  AND U9412 ( .A(n9576), .B(n9577), .Z(n9575) );
  XNOR U9413 ( .A(n9574), .B(n9533), .Z(n9577) );
  XOR U9414 ( .A(n9578), .B(n9570), .Z(n9533) );
  XNOR U9415 ( .A(n9579), .B(n9565), .Z(n9570) );
  XOR U9416 ( .A(n9580), .B(n9581), .Z(n9565) );
  AND U9417 ( .A(n9582), .B(n9583), .Z(n9581) );
  XOR U9418 ( .A(n9584), .B(n9580), .Z(n9582) );
  XNOR U9419 ( .A(n9585), .B(n9586), .Z(n9579) );
  AND U9420 ( .A(n9587), .B(n9588), .Z(n9586) );
  XOR U9421 ( .A(n9585), .B(n9589), .Z(n9587) );
  XNOR U9422 ( .A(n9571), .B(n9568), .Z(n9578) );
  AND U9423 ( .A(n9590), .B(n9591), .Z(n9568) );
  XOR U9424 ( .A(n9592), .B(n9593), .Z(n9571) );
  AND U9425 ( .A(n9594), .B(n9595), .Z(n9593) );
  XOR U9426 ( .A(n9592), .B(n9596), .Z(n9594) );
  XNOR U9427 ( .A(n9530), .B(n9574), .Z(n9576) );
  XNOR U9428 ( .A(n9597), .B(n9598), .Z(n9530) );
  AND U9429 ( .A(n127), .B(n9536), .Z(n9598) );
  XOR U9430 ( .A(n9597), .B(n9534), .Z(n9536) );
  XOR U9431 ( .A(n9599), .B(n9600), .Z(n9574) );
  AND U9432 ( .A(n9601), .B(n9602), .Z(n9600) );
  XNOR U9433 ( .A(n9599), .B(n9590), .Z(n9602) );
  IV U9434 ( .A(n9544), .Z(n9590) );
  XNOR U9435 ( .A(n9603), .B(n9583), .Z(n9544) );
  XNOR U9436 ( .A(n9604), .B(n9589), .Z(n9583) );
  XOR U9437 ( .A(n9605), .B(n9606), .Z(n9589) );
  NOR U9438 ( .A(n9607), .B(n9608), .Z(n9606) );
  XNOR U9439 ( .A(n9605), .B(n9609), .Z(n9607) );
  XNOR U9440 ( .A(n9588), .B(n9580), .Z(n9604) );
  XOR U9441 ( .A(n9610), .B(n9611), .Z(n9580) );
  AND U9442 ( .A(n9612), .B(n9613), .Z(n9611) );
  XNOR U9443 ( .A(n9610), .B(n9614), .Z(n9612) );
  XNOR U9444 ( .A(n9615), .B(n9585), .Z(n9588) );
  XOR U9445 ( .A(n9616), .B(n9617), .Z(n9585) );
  AND U9446 ( .A(n9618), .B(n9619), .Z(n9617) );
  XOR U9447 ( .A(n9616), .B(n9620), .Z(n9618) );
  XNOR U9448 ( .A(n9621), .B(n9622), .Z(n9615) );
  NOR U9449 ( .A(n9623), .B(n9624), .Z(n9622) );
  XOR U9450 ( .A(n9621), .B(n9625), .Z(n9623) );
  XNOR U9451 ( .A(n9584), .B(n9591), .Z(n9603) );
  NOR U9452 ( .A(n9552), .B(n9626), .Z(n9591) );
  XOR U9453 ( .A(n9596), .B(n9595), .Z(n9584) );
  XNOR U9454 ( .A(n9627), .B(n9592), .Z(n9595) );
  XOR U9455 ( .A(n9628), .B(n9629), .Z(n9592) );
  AND U9456 ( .A(n9630), .B(n9631), .Z(n9629) );
  XOR U9457 ( .A(n9628), .B(n9632), .Z(n9630) );
  XNOR U9458 ( .A(n9633), .B(n9634), .Z(n9627) );
  NOR U9459 ( .A(n9635), .B(n9636), .Z(n9634) );
  XNOR U9460 ( .A(n9633), .B(n9637), .Z(n9635) );
  XOR U9461 ( .A(n9638), .B(n9639), .Z(n9596) );
  NOR U9462 ( .A(n9640), .B(n9641), .Z(n9639) );
  XNOR U9463 ( .A(n9638), .B(n9642), .Z(n9640) );
  XNOR U9464 ( .A(n9541), .B(n9599), .Z(n9601) );
  XNOR U9465 ( .A(n9643), .B(n9644), .Z(n9541) );
  AND U9466 ( .A(n127), .B(n9548), .Z(n9644) );
  XOR U9467 ( .A(n9643), .B(n9546), .Z(n9548) );
  AND U9468 ( .A(n9549), .B(n9552), .Z(n9599) );
  XOR U9469 ( .A(n9645), .B(n9626), .Z(n9552) );
  XNOR U9470 ( .A(p_input[1024]), .B(p_input[128]), .Z(n9626) );
  XOR U9471 ( .A(n9614), .B(n9613), .Z(n9645) );
  XNOR U9472 ( .A(n9646), .B(n9620), .Z(n9613) );
  XNOR U9473 ( .A(n9609), .B(n9608), .Z(n9620) );
  XOR U9474 ( .A(n9647), .B(n9605), .Z(n9608) );
  XOR U9475 ( .A(p_input[1034]), .B(p_input[138]), .Z(n9605) );
  XNOR U9476 ( .A(p_input[1035]), .B(p_input[139]), .Z(n9647) );
  XOR U9477 ( .A(p_input[1036]), .B(p_input[140]), .Z(n9609) );
  XNOR U9478 ( .A(n9619), .B(n9610), .Z(n9646) );
  XOR U9479 ( .A(p_input[1025]), .B(p_input[129]), .Z(n9610) );
  XOR U9480 ( .A(n9648), .B(n9625), .Z(n9619) );
  XNOR U9481 ( .A(p_input[1039]), .B(p_input[143]), .Z(n9625) );
  XOR U9482 ( .A(n9616), .B(n9624), .Z(n9648) );
  XOR U9483 ( .A(n9649), .B(n9621), .Z(n9624) );
  XOR U9484 ( .A(p_input[1037]), .B(p_input[141]), .Z(n9621) );
  XNOR U9485 ( .A(p_input[1038]), .B(p_input[142]), .Z(n9649) );
  XOR U9486 ( .A(p_input[1033]), .B(p_input[137]), .Z(n9616) );
  XNOR U9487 ( .A(n9632), .B(n9631), .Z(n9614) );
  XNOR U9488 ( .A(n9650), .B(n9637), .Z(n9631) );
  XOR U9489 ( .A(p_input[1032]), .B(p_input[136]), .Z(n9637) );
  XOR U9490 ( .A(n9628), .B(n9636), .Z(n9650) );
  XOR U9491 ( .A(n9651), .B(n9633), .Z(n9636) );
  XOR U9492 ( .A(p_input[1030]), .B(p_input[134]), .Z(n9633) );
  XNOR U9493 ( .A(p_input[1031]), .B(p_input[135]), .Z(n9651) );
  XOR U9494 ( .A(p_input[1026]), .B(p_input[130]), .Z(n9628) );
  XNOR U9495 ( .A(n9642), .B(n9641), .Z(n9632) );
  XOR U9496 ( .A(n9652), .B(n9638), .Z(n9641) );
  XOR U9497 ( .A(p_input[1027]), .B(p_input[131]), .Z(n9638) );
  XNOR U9498 ( .A(p_input[1028]), .B(p_input[132]), .Z(n9652) );
  XOR U9499 ( .A(p_input[1029]), .B(p_input[133]), .Z(n9642) );
  XNOR U9500 ( .A(n9653), .B(n9654), .Z(n9549) );
  AND U9501 ( .A(n127), .B(n9655), .Z(n9654) );
  XNOR U9502 ( .A(n9656), .B(n9657), .Z(n127) );
  AND U9503 ( .A(n9658), .B(n9659), .Z(n9657) );
  XOR U9504 ( .A(n9656), .B(n9559), .Z(n9659) );
  XNOR U9505 ( .A(n9656), .B(n9513), .Z(n9658) );
  XOR U9506 ( .A(n9660), .B(n9661), .Z(n9656) );
  AND U9507 ( .A(n9662), .B(n9663), .Z(n9661) );
  XOR U9508 ( .A(n9660), .B(n9523), .Z(n9662) );
  XOR U9509 ( .A(n9664), .B(n9665), .Z(n9502) );
  AND U9510 ( .A(n131), .B(n9655), .Z(n9665) );
  XNOR U9511 ( .A(n9653), .B(n9664), .Z(n9655) );
  XNOR U9512 ( .A(n9666), .B(n9667), .Z(n131) );
  AND U9513 ( .A(n9668), .B(n9669), .Z(n9667) );
  XNOR U9514 ( .A(n9670), .B(n9666), .Z(n9669) );
  IV U9515 ( .A(n9559), .Z(n9670) );
  XNOR U9516 ( .A(n9671), .B(n9672), .Z(n9559) );
  AND U9517 ( .A(n134), .B(n9673), .Z(n9672) );
  XNOR U9518 ( .A(n9671), .B(n9674), .Z(n9673) );
  XNOR U9519 ( .A(n9513), .B(n9666), .Z(n9668) );
  XOR U9520 ( .A(n9675), .B(n9676), .Z(n9513) );
  AND U9521 ( .A(n142), .B(n9677), .Z(n9676) );
  XOR U9522 ( .A(n9660), .B(n9678), .Z(n9666) );
  AND U9523 ( .A(n9679), .B(n9663), .Z(n9678) );
  XNOR U9524 ( .A(n9572), .B(n9660), .Z(n9663) );
  XNOR U9525 ( .A(n9680), .B(n9681), .Z(n9572) );
  AND U9526 ( .A(n134), .B(n9682), .Z(n9681) );
  XOR U9527 ( .A(n9683), .B(n9680), .Z(n9682) );
  XNOR U9528 ( .A(n9684), .B(n9660), .Z(n9679) );
  IV U9529 ( .A(n9523), .Z(n9684) );
  XOR U9530 ( .A(n9685), .B(n9686), .Z(n9523) );
  AND U9531 ( .A(n142), .B(n9687), .Z(n9686) );
  XOR U9532 ( .A(n9688), .B(n9689), .Z(n9660) );
  AND U9533 ( .A(n9690), .B(n9691), .Z(n9689) );
  XNOR U9534 ( .A(n9597), .B(n9688), .Z(n9691) );
  XNOR U9535 ( .A(n9692), .B(n9693), .Z(n9597) );
  AND U9536 ( .A(n134), .B(n9694), .Z(n9693) );
  XNOR U9537 ( .A(n9695), .B(n9692), .Z(n9694) );
  XOR U9538 ( .A(n9688), .B(n9534), .Z(n9690) );
  XOR U9539 ( .A(n9696), .B(n9697), .Z(n9534) );
  AND U9540 ( .A(n142), .B(n9698), .Z(n9697) );
  XOR U9541 ( .A(n9699), .B(n9700), .Z(n9688) );
  AND U9542 ( .A(n9701), .B(n9702), .Z(n9700) );
  XNOR U9543 ( .A(n9699), .B(n9643), .Z(n9702) );
  XNOR U9544 ( .A(n9703), .B(n9704), .Z(n9643) );
  AND U9545 ( .A(n134), .B(n9705), .Z(n9704) );
  XOR U9546 ( .A(n9706), .B(n9703), .Z(n9705) );
  XNOR U9547 ( .A(n9707), .B(n9699), .Z(n9701) );
  IV U9548 ( .A(n9546), .Z(n9707) );
  XOR U9549 ( .A(n9708), .B(n9709), .Z(n9546) );
  AND U9550 ( .A(n142), .B(n9710), .Z(n9709) );
  AND U9551 ( .A(n9664), .B(n9653), .Z(n9699) );
  XNOR U9552 ( .A(n9711), .B(n9712), .Z(n9653) );
  AND U9553 ( .A(n134), .B(n9713), .Z(n9712) );
  XNOR U9554 ( .A(n9714), .B(n9711), .Z(n9713) );
  XNOR U9555 ( .A(n9715), .B(n9716), .Z(n134) );
  AND U9556 ( .A(n9717), .B(n9718), .Z(n9716) );
  XOR U9557 ( .A(n9674), .B(n9715), .Z(n9718) );
  AND U9558 ( .A(n9719), .B(n9720), .Z(n9674) );
  XOR U9559 ( .A(n9715), .B(n9671), .Z(n9717) );
  XNOR U9560 ( .A(n9721), .B(n9722), .Z(n9671) );
  AND U9561 ( .A(n138), .B(n9677), .Z(n9722) );
  XOR U9562 ( .A(n9675), .B(n9721), .Z(n9677) );
  XOR U9563 ( .A(n9723), .B(n9724), .Z(n9715) );
  AND U9564 ( .A(n9725), .B(n9726), .Z(n9724) );
  XNOR U9565 ( .A(n9723), .B(n9719), .Z(n9726) );
  IV U9566 ( .A(n9683), .Z(n9719) );
  XOR U9567 ( .A(n9727), .B(n9728), .Z(n9683) );
  XOR U9568 ( .A(n9729), .B(n9720), .Z(n9728) );
  AND U9569 ( .A(n9695), .B(n9730), .Z(n9720) );
  AND U9570 ( .A(n9731), .B(n9732), .Z(n9729) );
  XOR U9571 ( .A(n9733), .B(n9727), .Z(n9731) );
  XNOR U9572 ( .A(n9680), .B(n9723), .Z(n9725) );
  XNOR U9573 ( .A(n9734), .B(n9735), .Z(n9680) );
  AND U9574 ( .A(n138), .B(n9687), .Z(n9735) );
  XOR U9575 ( .A(n9734), .B(n9685), .Z(n9687) );
  XOR U9576 ( .A(n9736), .B(n9737), .Z(n9723) );
  AND U9577 ( .A(n9738), .B(n9739), .Z(n9737) );
  XNOR U9578 ( .A(n9736), .B(n9695), .Z(n9739) );
  XOR U9579 ( .A(n9740), .B(n9732), .Z(n9695) );
  XNOR U9580 ( .A(n9741), .B(n9727), .Z(n9732) );
  XOR U9581 ( .A(n9742), .B(n9743), .Z(n9727) );
  AND U9582 ( .A(n9744), .B(n9745), .Z(n9743) );
  XOR U9583 ( .A(n9746), .B(n9742), .Z(n9744) );
  XNOR U9584 ( .A(n9747), .B(n9748), .Z(n9741) );
  AND U9585 ( .A(n9749), .B(n9750), .Z(n9748) );
  XOR U9586 ( .A(n9747), .B(n9751), .Z(n9749) );
  XNOR U9587 ( .A(n9733), .B(n9730), .Z(n9740) );
  AND U9588 ( .A(n9752), .B(n9753), .Z(n9730) );
  XOR U9589 ( .A(n9754), .B(n9755), .Z(n9733) );
  AND U9590 ( .A(n9756), .B(n9757), .Z(n9755) );
  XOR U9591 ( .A(n9754), .B(n9758), .Z(n9756) );
  XNOR U9592 ( .A(n9692), .B(n9736), .Z(n9738) );
  XNOR U9593 ( .A(n9759), .B(n9760), .Z(n9692) );
  AND U9594 ( .A(n138), .B(n9698), .Z(n9760) );
  XOR U9595 ( .A(n9759), .B(n9696), .Z(n9698) );
  XOR U9596 ( .A(n9761), .B(n9762), .Z(n9736) );
  AND U9597 ( .A(n9763), .B(n9764), .Z(n9762) );
  XNOR U9598 ( .A(n9761), .B(n9752), .Z(n9764) );
  IV U9599 ( .A(n9706), .Z(n9752) );
  XNOR U9600 ( .A(n9765), .B(n9745), .Z(n9706) );
  XNOR U9601 ( .A(n9766), .B(n9751), .Z(n9745) );
  XOR U9602 ( .A(n9767), .B(n9768), .Z(n9751) );
  NOR U9603 ( .A(n9769), .B(n9770), .Z(n9768) );
  XNOR U9604 ( .A(n9767), .B(n9771), .Z(n9769) );
  XNOR U9605 ( .A(n9750), .B(n9742), .Z(n9766) );
  XOR U9606 ( .A(n9772), .B(n9773), .Z(n9742) );
  AND U9607 ( .A(n9774), .B(n9775), .Z(n9773) );
  XNOR U9608 ( .A(n9772), .B(n9776), .Z(n9774) );
  XNOR U9609 ( .A(n9777), .B(n9747), .Z(n9750) );
  XOR U9610 ( .A(n9778), .B(n9779), .Z(n9747) );
  AND U9611 ( .A(n9780), .B(n9781), .Z(n9779) );
  XOR U9612 ( .A(n9778), .B(n9782), .Z(n9780) );
  XNOR U9613 ( .A(n9783), .B(n9784), .Z(n9777) );
  NOR U9614 ( .A(n9785), .B(n9786), .Z(n9784) );
  XOR U9615 ( .A(n9783), .B(n9787), .Z(n9785) );
  XNOR U9616 ( .A(n9746), .B(n9753), .Z(n9765) );
  NOR U9617 ( .A(n9714), .B(n9788), .Z(n9753) );
  XOR U9618 ( .A(n9758), .B(n9757), .Z(n9746) );
  XNOR U9619 ( .A(n9789), .B(n9754), .Z(n9757) );
  XOR U9620 ( .A(n9790), .B(n9791), .Z(n9754) );
  AND U9621 ( .A(n9792), .B(n9793), .Z(n9791) );
  XOR U9622 ( .A(n9790), .B(n9794), .Z(n9792) );
  XNOR U9623 ( .A(n9795), .B(n9796), .Z(n9789) );
  NOR U9624 ( .A(n9797), .B(n9798), .Z(n9796) );
  XNOR U9625 ( .A(n9795), .B(n9799), .Z(n9797) );
  XOR U9626 ( .A(n9800), .B(n9801), .Z(n9758) );
  NOR U9627 ( .A(n9802), .B(n9803), .Z(n9801) );
  XNOR U9628 ( .A(n9800), .B(n9804), .Z(n9802) );
  XNOR U9629 ( .A(n9703), .B(n9761), .Z(n9763) );
  XNOR U9630 ( .A(n9805), .B(n9806), .Z(n9703) );
  AND U9631 ( .A(n138), .B(n9710), .Z(n9806) );
  XOR U9632 ( .A(n9805), .B(n9708), .Z(n9710) );
  AND U9633 ( .A(n9711), .B(n9714), .Z(n9761) );
  XOR U9634 ( .A(n9807), .B(n9788), .Z(n9714) );
  XNOR U9635 ( .A(p_input[1024]), .B(p_input[144]), .Z(n9788) );
  XOR U9636 ( .A(n9776), .B(n9775), .Z(n9807) );
  XNOR U9637 ( .A(n9808), .B(n9782), .Z(n9775) );
  XNOR U9638 ( .A(n9771), .B(n9770), .Z(n9782) );
  XOR U9639 ( .A(n9809), .B(n9767), .Z(n9770) );
  XOR U9640 ( .A(p_input[1034]), .B(p_input[154]), .Z(n9767) );
  XNOR U9641 ( .A(p_input[1035]), .B(p_input[155]), .Z(n9809) );
  XOR U9642 ( .A(p_input[1036]), .B(p_input[156]), .Z(n9771) );
  XNOR U9643 ( .A(n9781), .B(n9772), .Z(n9808) );
  XOR U9644 ( .A(p_input[1025]), .B(p_input[145]), .Z(n9772) );
  XOR U9645 ( .A(n9810), .B(n9787), .Z(n9781) );
  XNOR U9646 ( .A(p_input[1039]), .B(p_input[159]), .Z(n9787) );
  XOR U9647 ( .A(n9778), .B(n9786), .Z(n9810) );
  XOR U9648 ( .A(n9811), .B(n9783), .Z(n9786) );
  XOR U9649 ( .A(p_input[1037]), .B(p_input[157]), .Z(n9783) );
  XNOR U9650 ( .A(p_input[1038]), .B(p_input[158]), .Z(n9811) );
  XOR U9651 ( .A(p_input[1033]), .B(p_input[153]), .Z(n9778) );
  XNOR U9652 ( .A(n9794), .B(n9793), .Z(n9776) );
  XNOR U9653 ( .A(n9812), .B(n9799), .Z(n9793) );
  XOR U9654 ( .A(p_input[1032]), .B(p_input[152]), .Z(n9799) );
  XOR U9655 ( .A(n9790), .B(n9798), .Z(n9812) );
  XOR U9656 ( .A(n9813), .B(n9795), .Z(n9798) );
  XOR U9657 ( .A(p_input[1030]), .B(p_input[150]), .Z(n9795) );
  XNOR U9658 ( .A(p_input[1031]), .B(p_input[151]), .Z(n9813) );
  XOR U9659 ( .A(p_input[1026]), .B(p_input[146]), .Z(n9790) );
  XNOR U9660 ( .A(n9804), .B(n9803), .Z(n9794) );
  XOR U9661 ( .A(n9814), .B(n9800), .Z(n9803) );
  XOR U9662 ( .A(p_input[1027]), .B(p_input[147]), .Z(n9800) );
  XNOR U9663 ( .A(p_input[1028]), .B(p_input[148]), .Z(n9814) );
  XOR U9664 ( .A(p_input[1029]), .B(p_input[149]), .Z(n9804) );
  XNOR U9665 ( .A(n9815), .B(n9816), .Z(n9711) );
  AND U9666 ( .A(n138), .B(n9817), .Z(n9816) );
  XNOR U9667 ( .A(n9818), .B(n9819), .Z(n138) );
  AND U9668 ( .A(n9820), .B(n9821), .Z(n9819) );
  XOR U9669 ( .A(n9818), .B(n9721), .Z(n9821) );
  XNOR U9670 ( .A(n9818), .B(n9675), .Z(n9820) );
  XOR U9671 ( .A(n9822), .B(n9823), .Z(n9818) );
  AND U9672 ( .A(n9824), .B(n9825), .Z(n9823) );
  XOR U9673 ( .A(n9822), .B(n9685), .Z(n9824) );
  XOR U9674 ( .A(n9826), .B(n9827), .Z(n9664) );
  AND U9675 ( .A(n142), .B(n9817), .Z(n9827) );
  XNOR U9676 ( .A(n9815), .B(n9826), .Z(n9817) );
  XNOR U9677 ( .A(n9828), .B(n9829), .Z(n142) );
  AND U9678 ( .A(n9830), .B(n9831), .Z(n9829) );
  XNOR U9679 ( .A(n9832), .B(n9828), .Z(n9831) );
  IV U9680 ( .A(n9721), .Z(n9832) );
  XNOR U9681 ( .A(n9833), .B(n9834), .Z(n9721) );
  AND U9682 ( .A(n145), .B(n9835), .Z(n9834) );
  XNOR U9683 ( .A(n9833), .B(n9836), .Z(n9835) );
  XNOR U9684 ( .A(n9675), .B(n9828), .Z(n9830) );
  XOR U9685 ( .A(n9837), .B(n9838), .Z(n9675) );
  AND U9686 ( .A(n153), .B(n9839), .Z(n9838) );
  XOR U9687 ( .A(n9822), .B(n9840), .Z(n9828) );
  AND U9688 ( .A(n9841), .B(n9825), .Z(n9840) );
  XNOR U9689 ( .A(n9734), .B(n9822), .Z(n9825) );
  XNOR U9690 ( .A(n9842), .B(n9843), .Z(n9734) );
  AND U9691 ( .A(n145), .B(n9844), .Z(n9843) );
  XOR U9692 ( .A(n9845), .B(n9842), .Z(n9844) );
  XNOR U9693 ( .A(n9846), .B(n9822), .Z(n9841) );
  IV U9694 ( .A(n9685), .Z(n9846) );
  XOR U9695 ( .A(n9847), .B(n9848), .Z(n9685) );
  AND U9696 ( .A(n153), .B(n9849), .Z(n9848) );
  XOR U9697 ( .A(n9850), .B(n9851), .Z(n9822) );
  AND U9698 ( .A(n9852), .B(n9853), .Z(n9851) );
  XNOR U9699 ( .A(n9759), .B(n9850), .Z(n9853) );
  XNOR U9700 ( .A(n9854), .B(n9855), .Z(n9759) );
  AND U9701 ( .A(n145), .B(n9856), .Z(n9855) );
  XNOR U9702 ( .A(n9857), .B(n9854), .Z(n9856) );
  XOR U9703 ( .A(n9850), .B(n9696), .Z(n9852) );
  XOR U9704 ( .A(n9858), .B(n9859), .Z(n9696) );
  AND U9705 ( .A(n153), .B(n9860), .Z(n9859) );
  XOR U9706 ( .A(n9861), .B(n9862), .Z(n9850) );
  AND U9707 ( .A(n9863), .B(n9864), .Z(n9862) );
  XNOR U9708 ( .A(n9861), .B(n9805), .Z(n9864) );
  XNOR U9709 ( .A(n9865), .B(n9866), .Z(n9805) );
  AND U9710 ( .A(n145), .B(n9867), .Z(n9866) );
  XOR U9711 ( .A(n9868), .B(n9865), .Z(n9867) );
  XNOR U9712 ( .A(n9869), .B(n9861), .Z(n9863) );
  IV U9713 ( .A(n9708), .Z(n9869) );
  XOR U9714 ( .A(n9870), .B(n9871), .Z(n9708) );
  AND U9715 ( .A(n153), .B(n9872), .Z(n9871) );
  AND U9716 ( .A(n9826), .B(n9815), .Z(n9861) );
  XNOR U9717 ( .A(n9873), .B(n9874), .Z(n9815) );
  AND U9718 ( .A(n145), .B(n9875), .Z(n9874) );
  XNOR U9719 ( .A(n9876), .B(n9873), .Z(n9875) );
  XNOR U9720 ( .A(n9877), .B(n9878), .Z(n145) );
  AND U9721 ( .A(n9879), .B(n9880), .Z(n9878) );
  XOR U9722 ( .A(n9836), .B(n9877), .Z(n9880) );
  AND U9723 ( .A(n9881), .B(n9882), .Z(n9836) );
  XOR U9724 ( .A(n9877), .B(n9833), .Z(n9879) );
  XNOR U9725 ( .A(n9883), .B(n9884), .Z(n9833) );
  AND U9726 ( .A(n149), .B(n9839), .Z(n9884) );
  XOR U9727 ( .A(n9837), .B(n9883), .Z(n9839) );
  XOR U9728 ( .A(n9885), .B(n9886), .Z(n9877) );
  AND U9729 ( .A(n9887), .B(n9888), .Z(n9886) );
  XNOR U9730 ( .A(n9885), .B(n9881), .Z(n9888) );
  IV U9731 ( .A(n9845), .Z(n9881) );
  XOR U9732 ( .A(n9889), .B(n9890), .Z(n9845) );
  XOR U9733 ( .A(n9891), .B(n9882), .Z(n9890) );
  AND U9734 ( .A(n9857), .B(n9892), .Z(n9882) );
  AND U9735 ( .A(n9893), .B(n9894), .Z(n9891) );
  XOR U9736 ( .A(n9895), .B(n9889), .Z(n9893) );
  XNOR U9737 ( .A(n9842), .B(n9885), .Z(n9887) );
  XNOR U9738 ( .A(n9896), .B(n9897), .Z(n9842) );
  AND U9739 ( .A(n149), .B(n9849), .Z(n9897) );
  XOR U9740 ( .A(n9896), .B(n9847), .Z(n9849) );
  XOR U9741 ( .A(n9898), .B(n9899), .Z(n9885) );
  AND U9742 ( .A(n9900), .B(n9901), .Z(n9899) );
  XNOR U9743 ( .A(n9898), .B(n9857), .Z(n9901) );
  XOR U9744 ( .A(n9902), .B(n9894), .Z(n9857) );
  XNOR U9745 ( .A(n9903), .B(n9889), .Z(n9894) );
  XOR U9746 ( .A(n9904), .B(n9905), .Z(n9889) );
  AND U9747 ( .A(n9906), .B(n9907), .Z(n9905) );
  XOR U9748 ( .A(n9908), .B(n9904), .Z(n9906) );
  XNOR U9749 ( .A(n9909), .B(n9910), .Z(n9903) );
  AND U9750 ( .A(n9911), .B(n9912), .Z(n9910) );
  XOR U9751 ( .A(n9909), .B(n9913), .Z(n9911) );
  XNOR U9752 ( .A(n9895), .B(n9892), .Z(n9902) );
  AND U9753 ( .A(n9914), .B(n9915), .Z(n9892) );
  XOR U9754 ( .A(n9916), .B(n9917), .Z(n9895) );
  AND U9755 ( .A(n9918), .B(n9919), .Z(n9917) );
  XOR U9756 ( .A(n9916), .B(n9920), .Z(n9918) );
  XNOR U9757 ( .A(n9854), .B(n9898), .Z(n9900) );
  XNOR U9758 ( .A(n9921), .B(n9922), .Z(n9854) );
  AND U9759 ( .A(n149), .B(n9860), .Z(n9922) );
  XOR U9760 ( .A(n9921), .B(n9858), .Z(n9860) );
  XOR U9761 ( .A(n9923), .B(n9924), .Z(n9898) );
  AND U9762 ( .A(n9925), .B(n9926), .Z(n9924) );
  XNOR U9763 ( .A(n9923), .B(n9914), .Z(n9926) );
  IV U9764 ( .A(n9868), .Z(n9914) );
  XNOR U9765 ( .A(n9927), .B(n9907), .Z(n9868) );
  XNOR U9766 ( .A(n9928), .B(n9913), .Z(n9907) );
  XOR U9767 ( .A(n9929), .B(n9930), .Z(n9913) );
  NOR U9768 ( .A(n9931), .B(n9932), .Z(n9930) );
  XNOR U9769 ( .A(n9929), .B(n9933), .Z(n9931) );
  XNOR U9770 ( .A(n9912), .B(n9904), .Z(n9928) );
  XOR U9771 ( .A(n9934), .B(n9935), .Z(n9904) );
  AND U9772 ( .A(n9936), .B(n9937), .Z(n9935) );
  XNOR U9773 ( .A(n9934), .B(n9938), .Z(n9936) );
  XNOR U9774 ( .A(n9939), .B(n9909), .Z(n9912) );
  XOR U9775 ( .A(n9940), .B(n9941), .Z(n9909) );
  AND U9776 ( .A(n9942), .B(n9943), .Z(n9941) );
  XOR U9777 ( .A(n9940), .B(n9944), .Z(n9942) );
  XNOR U9778 ( .A(n9945), .B(n9946), .Z(n9939) );
  NOR U9779 ( .A(n9947), .B(n9948), .Z(n9946) );
  XOR U9780 ( .A(n9945), .B(n9949), .Z(n9947) );
  XNOR U9781 ( .A(n9908), .B(n9915), .Z(n9927) );
  NOR U9782 ( .A(n9876), .B(n9950), .Z(n9915) );
  XOR U9783 ( .A(n9920), .B(n9919), .Z(n9908) );
  XNOR U9784 ( .A(n9951), .B(n9916), .Z(n9919) );
  XOR U9785 ( .A(n9952), .B(n9953), .Z(n9916) );
  AND U9786 ( .A(n9954), .B(n9955), .Z(n9953) );
  XOR U9787 ( .A(n9952), .B(n9956), .Z(n9954) );
  XNOR U9788 ( .A(n9957), .B(n9958), .Z(n9951) );
  NOR U9789 ( .A(n9959), .B(n9960), .Z(n9958) );
  XNOR U9790 ( .A(n9957), .B(n9961), .Z(n9959) );
  XOR U9791 ( .A(n9962), .B(n9963), .Z(n9920) );
  NOR U9792 ( .A(n9964), .B(n9965), .Z(n9963) );
  XNOR U9793 ( .A(n9962), .B(n9966), .Z(n9964) );
  XNOR U9794 ( .A(n9865), .B(n9923), .Z(n9925) );
  XNOR U9795 ( .A(n9967), .B(n9968), .Z(n9865) );
  AND U9796 ( .A(n149), .B(n9872), .Z(n9968) );
  XOR U9797 ( .A(n9967), .B(n9870), .Z(n9872) );
  AND U9798 ( .A(n9873), .B(n9876), .Z(n9923) );
  XOR U9799 ( .A(n9969), .B(n9950), .Z(n9876) );
  XNOR U9800 ( .A(p_input[1024]), .B(p_input[160]), .Z(n9950) );
  XOR U9801 ( .A(n9938), .B(n9937), .Z(n9969) );
  XNOR U9802 ( .A(n9970), .B(n9944), .Z(n9937) );
  XNOR U9803 ( .A(n9933), .B(n9932), .Z(n9944) );
  XOR U9804 ( .A(n9971), .B(n9929), .Z(n9932) );
  XOR U9805 ( .A(p_input[1034]), .B(p_input[170]), .Z(n9929) );
  XNOR U9806 ( .A(p_input[1035]), .B(p_input[171]), .Z(n9971) );
  XOR U9807 ( .A(p_input[1036]), .B(p_input[172]), .Z(n9933) );
  XNOR U9808 ( .A(n9943), .B(n9934), .Z(n9970) );
  XOR U9809 ( .A(p_input[1025]), .B(p_input[161]), .Z(n9934) );
  XOR U9810 ( .A(n9972), .B(n9949), .Z(n9943) );
  XNOR U9811 ( .A(p_input[1039]), .B(p_input[175]), .Z(n9949) );
  XOR U9812 ( .A(n9940), .B(n9948), .Z(n9972) );
  XOR U9813 ( .A(n9973), .B(n9945), .Z(n9948) );
  XOR U9814 ( .A(p_input[1037]), .B(p_input[173]), .Z(n9945) );
  XNOR U9815 ( .A(p_input[1038]), .B(p_input[174]), .Z(n9973) );
  XOR U9816 ( .A(p_input[1033]), .B(p_input[169]), .Z(n9940) );
  XNOR U9817 ( .A(n9956), .B(n9955), .Z(n9938) );
  XNOR U9818 ( .A(n9974), .B(n9961), .Z(n9955) );
  XOR U9819 ( .A(p_input[1032]), .B(p_input[168]), .Z(n9961) );
  XOR U9820 ( .A(n9952), .B(n9960), .Z(n9974) );
  XOR U9821 ( .A(n9975), .B(n9957), .Z(n9960) );
  XOR U9822 ( .A(p_input[1030]), .B(p_input[166]), .Z(n9957) );
  XNOR U9823 ( .A(p_input[1031]), .B(p_input[167]), .Z(n9975) );
  XOR U9824 ( .A(p_input[1026]), .B(p_input[162]), .Z(n9952) );
  XNOR U9825 ( .A(n9966), .B(n9965), .Z(n9956) );
  XOR U9826 ( .A(n9976), .B(n9962), .Z(n9965) );
  XOR U9827 ( .A(p_input[1027]), .B(p_input[163]), .Z(n9962) );
  XNOR U9828 ( .A(p_input[1028]), .B(p_input[164]), .Z(n9976) );
  XOR U9829 ( .A(p_input[1029]), .B(p_input[165]), .Z(n9966) );
  XNOR U9830 ( .A(n9977), .B(n9978), .Z(n9873) );
  AND U9831 ( .A(n149), .B(n9979), .Z(n9978) );
  XNOR U9832 ( .A(n9980), .B(n9981), .Z(n149) );
  AND U9833 ( .A(n9982), .B(n9983), .Z(n9981) );
  XOR U9834 ( .A(n9980), .B(n9883), .Z(n9983) );
  XNOR U9835 ( .A(n9980), .B(n9837), .Z(n9982) );
  XOR U9836 ( .A(n9984), .B(n9985), .Z(n9980) );
  AND U9837 ( .A(n9986), .B(n9987), .Z(n9985) );
  XOR U9838 ( .A(n9984), .B(n9847), .Z(n9986) );
  XOR U9839 ( .A(n9988), .B(n9989), .Z(n9826) );
  AND U9840 ( .A(n153), .B(n9979), .Z(n9989) );
  XNOR U9841 ( .A(n9977), .B(n9988), .Z(n9979) );
  XNOR U9842 ( .A(n9990), .B(n9991), .Z(n153) );
  AND U9843 ( .A(n9992), .B(n9993), .Z(n9991) );
  XNOR U9844 ( .A(n9994), .B(n9990), .Z(n9993) );
  IV U9845 ( .A(n9883), .Z(n9994) );
  XNOR U9846 ( .A(n9995), .B(n9996), .Z(n9883) );
  AND U9847 ( .A(n156), .B(n9997), .Z(n9996) );
  XNOR U9848 ( .A(n9995), .B(n9998), .Z(n9997) );
  XNOR U9849 ( .A(n9837), .B(n9990), .Z(n9992) );
  XOR U9850 ( .A(n9999), .B(n10000), .Z(n9837) );
  AND U9851 ( .A(n164), .B(n10001), .Z(n10000) );
  XOR U9852 ( .A(n9984), .B(n10002), .Z(n9990) );
  AND U9853 ( .A(n10003), .B(n9987), .Z(n10002) );
  XNOR U9854 ( .A(n9896), .B(n9984), .Z(n9987) );
  XNOR U9855 ( .A(n10004), .B(n10005), .Z(n9896) );
  AND U9856 ( .A(n156), .B(n10006), .Z(n10005) );
  XOR U9857 ( .A(n10007), .B(n10004), .Z(n10006) );
  XNOR U9858 ( .A(n10008), .B(n9984), .Z(n10003) );
  IV U9859 ( .A(n9847), .Z(n10008) );
  XOR U9860 ( .A(n10009), .B(n10010), .Z(n9847) );
  AND U9861 ( .A(n164), .B(n10011), .Z(n10010) );
  XOR U9862 ( .A(n10012), .B(n10013), .Z(n9984) );
  AND U9863 ( .A(n10014), .B(n10015), .Z(n10013) );
  XNOR U9864 ( .A(n9921), .B(n10012), .Z(n10015) );
  XNOR U9865 ( .A(n10016), .B(n10017), .Z(n9921) );
  AND U9866 ( .A(n156), .B(n10018), .Z(n10017) );
  XNOR U9867 ( .A(n10019), .B(n10016), .Z(n10018) );
  XOR U9868 ( .A(n10012), .B(n9858), .Z(n10014) );
  XOR U9869 ( .A(n10020), .B(n10021), .Z(n9858) );
  AND U9870 ( .A(n164), .B(n10022), .Z(n10021) );
  XOR U9871 ( .A(n10023), .B(n10024), .Z(n10012) );
  AND U9872 ( .A(n10025), .B(n10026), .Z(n10024) );
  XNOR U9873 ( .A(n10023), .B(n9967), .Z(n10026) );
  XNOR U9874 ( .A(n10027), .B(n10028), .Z(n9967) );
  AND U9875 ( .A(n156), .B(n10029), .Z(n10028) );
  XOR U9876 ( .A(n10030), .B(n10027), .Z(n10029) );
  XNOR U9877 ( .A(n10031), .B(n10023), .Z(n10025) );
  IV U9878 ( .A(n9870), .Z(n10031) );
  XOR U9879 ( .A(n10032), .B(n10033), .Z(n9870) );
  AND U9880 ( .A(n164), .B(n10034), .Z(n10033) );
  AND U9881 ( .A(n9988), .B(n9977), .Z(n10023) );
  XNOR U9882 ( .A(n10035), .B(n10036), .Z(n9977) );
  AND U9883 ( .A(n156), .B(n10037), .Z(n10036) );
  XNOR U9884 ( .A(n10038), .B(n10035), .Z(n10037) );
  XNOR U9885 ( .A(n10039), .B(n10040), .Z(n156) );
  AND U9886 ( .A(n10041), .B(n10042), .Z(n10040) );
  XOR U9887 ( .A(n9998), .B(n10039), .Z(n10042) );
  AND U9888 ( .A(n10043), .B(n10044), .Z(n9998) );
  XOR U9889 ( .A(n10039), .B(n9995), .Z(n10041) );
  XNOR U9890 ( .A(n10045), .B(n10046), .Z(n9995) );
  AND U9891 ( .A(n160), .B(n10001), .Z(n10046) );
  XOR U9892 ( .A(n9999), .B(n10045), .Z(n10001) );
  XOR U9893 ( .A(n10047), .B(n10048), .Z(n10039) );
  AND U9894 ( .A(n10049), .B(n10050), .Z(n10048) );
  XNOR U9895 ( .A(n10047), .B(n10043), .Z(n10050) );
  IV U9896 ( .A(n10007), .Z(n10043) );
  XOR U9897 ( .A(n10051), .B(n10052), .Z(n10007) );
  XOR U9898 ( .A(n10053), .B(n10044), .Z(n10052) );
  AND U9899 ( .A(n10019), .B(n10054), .Z(n10044) );
  AND U9900 ( .A(n10055), .B(n10056), .Z(n10053) );
  XOR U9901 ( .A(n10057), .B(n10051), .Z(n10055) );
  XNOR U9902 ( .A(n10004), .B(n10047), .Z(n10049) );
  XNOR U9903 ( .A(n10058), .B(n10059), .Z(n10004) );
  AND U9904 ( .A(n160), .B(n10011), .Z(n10059) );
  XOR U9905 ( .A(n10058), .B(n10009), .Z(n10011) );
  XOR U9906 ( .A(n10060), .B(n10061), .Z(n10047) );
  AND U9907 ( .A(n10062), .B(n10063), .Z(n10061) );
  XNOR U9908 ( .A(n10060), .B(n10019), .Z(n10063) );
  XOR U9909 ( .A(n10064), .B(n10056), .Z(n10019) );
  XNOR U9910 ( .A(n10065), .B(n10051), .Z(n10056) );
  XOR U9911 ( .A(n10066), .B(n10067), .Z(n10051) );
  AND U9912 ( .A(n10068), .B(n10069), .Z(n10067) );
  XOR U9913 ( .A(n10070), .B(n10066), .Z(n10068) );
  XNOR U9914 ( .A(n10071), .B(n10072), .Z(n10065) );
  AND U9915 ( .A(n10073), .B(n10074), .Z(n10072) );
  XOR U9916 ( .A(n10071), .B(n10075), .Z(n10073) );
  XNOR U9917 ( .A(n10057), .B(n10054), .Z(n10064) );
  AND U9918 ( .A(n10076), .B(n10077), .Z(n10054) );
  XOR U9919 ( .A(n10078), .B(n10079), .Z(n10057) );
  AND U9920 ( .A(n10080), .B(n10081), .Z(n10079) );
  XOR U9921 ( .A(n10078), .B(n10082), .Z(n10080) );
  XNOR U9922 ( .A(n10016), .B(n10060), .Z(n10062) );
  XNOR U9923 ( .A(n10083), .B(n10084), .Z(n10016) );
  AND U9924 ( .A(n160), .B(n10022), .Z(n10084) );
  XOR U9925 ( .A(n10083), .B(n10020), .Z(n10022) );
  XOR U9926 ( .A(n10085), .B(n10086), .Z(n10060) );
  AND U9927 ( .A(n10087), .B(n10088), .Z(n10086) );
  XNOR U9928 ( .A(n10085), .B(n10076), .Z(n10088) );
  IV U9929 ( .A(n10030), .Z(n10076) );
  XNOR U9930 ( .A(n10089), .B(n10069), .Z(n10030) );
  XNOR U9931 ( .A(n10090), .B(n10075), .Z(n10069) );
  XOR U9932 ( .A(n10091), .B(n10092), .Z(n10075) );
  NOR U9933 ( .A(n10093), .B(n10094), .Z(n10092) );
  XNOR U9934 ( .A(n10091), .B(n10095), .Z(n10093) );
  XNOR U9935 ( .A(n10074), .B(n10066), .Z(n10090) );
  XOR U9936 ( .A(n10096), .B(n10097), .Z(n10066) );
  AND U9937 ( .A(n10098), .B(n10099), .Z(n10097) );
  XNOR U9938 ( .A(n10096), .B(n10100), .Z(n10098) );
  XNOR U9939 ( .A(n10101), .B(n10071), .Z(n10074) );
  XOR U9940 ( .A(n10102), .B(n10103), .Z(n10071) );
  AND U9941 ( .A(n10104), .B(n10105), .Z(n10103) );
  XOR U9942 ( .A(n10102), .B(n10106), .Z(n10104) );
  XNOR U9943 ( .A(n10107), .B(n10108), .Z(n10101) );
  NOR U9944 ( .A(n10109), .B(n10110), .Z(n10108) );
  XOR U9945 ( .A(n10107), .B(n10111), .Z(n10109) );
  XNOR U9946 ( .A(n10070), .B(n10077), .Z(n10089) );
  NOR U9947 ( .A(n10038), .B(n10112), .Z(n10077) );
  XOR U9948 ( .A(n10082), .B(n10081), .Z(n10070) );
  XNOR U9949 ( .A(n10113), .B(n10078), .Z(n10081) );
  XOR U9950 ( .A(n10114), .B(n10115), .Z(n10078) );
  AND U9951 ( .A(n10116), .B(n10117), .Z(n10115) );
  XOR U9952 ( .A(n10114), .B(n10118), .Z(n10116) );
  XNOR U9953 ( .A(n10119), .B(n10120), .Z(n10113) );
  NOR U9954 ( .A(n10121), .B(n10122), .Z(n10120) );
  XNOR U9955 ( .A(n10119), .B(n10123), .Z(n10121) );
  XOR U9956 ( .A(n10124), .B(n10125), .Z(n10082) );
  NOR U9957 ( .A(n10126), .B(n10127), .Z(n10125) );
  XNOR U9958 ( .A(n10124), .B(n10128), .Z(n10126) );
  XNOR U9959 ( .A(n10027), .B(n10085), .Z(n10087) );
  XNOR U9960 ( .A(n10129), .B(n10130), .Z(n10027) );
  AND U9961 ( .A(n160), .B(n10034), .Z(n10130) );
  XOR U9962 ( .A(n10129), .B(n10032), .Z(n10034) );
  AND U9963 ( .A(n10035), .B(n10038), .Z(n10085) );
  XOR U9964 ( .A(n10131), .B(n10112), .Z(n10038) );
  XNOR U9965 ( .A(p_input[1024]), .B(p_input[176]), .Z(n10112) );
  XOR U9966 ( .A(n10100), .B(n10099), .Z(n10131) );
  XNOR U9967 ( .A(n10132), .B(n10106), .Z(n10099) );
  XNOR U9968 ( .A(n10095), .B(n10094), .Z(n10106) );
  XOR U9969 ( .A(n10133), .B(n10091), .Z(n10094) );
  XOR U9970 ( .A(p_input[1034]), .B(p_input[186]), .Z(n10091) );
  XNOR U9971 ( .A(p_input[1035]), .B(p_input[187]), .Z(n10133) );
  XOR U9972 ( .A(p_input[1036]), .B(p_input[188]), .Z(n10095) );
  XNOR U9973 ( .A(n10105), .B(n10096), .Z(n10132) );
  XOR U9974 ( .A(p_input[1025]), .B(p_input[177]), .Z(n10096) );
  XOR U9975 ( .A(n10134), .B(n10111), .Z(n10105) );
  XNOR U9976 ( .A(p_input[1039]), .B(p_input[191]), .Z(n10111) );
  XOR U9977 ( .A(n10102), .B(n10110), .Z(n10134) );
  XOR U9978 ( .A(n10135), .B(n10107), .Z(n10110) );
  XOR U9979 ( .A(p_input[1037]), .B(p_input[189]), .Z(n10107) );
  XNOR U9980 ( .A(p_input[1038]), .B(p_input[190]), .Z(n10135) );
  XOR U9981 ( .A(p_input[1033]), .B(p_input[185]), .Z(n10102) );
  XNOR U9982 ( .A(n10118), .B(n10117), .Z(n10100) );
  XNOR U9983 ( .A(n10136), .B(n10123), .Z(n10117) );
  XOR U9984 ( .A(p_input[1032]), .B(p_input[184]), .Z(n10123) );
  XOR U9985 ( .A(n10114), .B(n10122), .Z(n10136) );
  XOR U9986 ( .A(n10137), .B(n10119), .Z(n10122) );
  XOR U9987 ( .A(p_input[1030]), .B(p_input[182]), .Z(n10119) );
  XNOR U9988 ( .A(p_input[1031]), .B(p_input[183]), .Z(n10137) );
  XOR U9989 ( .A(p_input[1026]), .B(p_input[178]), .Z(n10114) );
  XNOR U9990 ( .A(n10128), .B(n10127), .Z(n10118) );
  XOR U9991 ( .A(n10138), .B(n10124), .Z(n10127) );
  XOR U9992 ( .A(p_input[1027]), .B(p_input[179]), .Z(n10124) );
  XNOR U9993 ( .A(p_input[1028]), .B(p_input[180]), .Z(n10138) );
  XOR U9994 ( .A(p_input[1029]), .B(p_input[181]), .Z(n10128) );
  XNOR U9995 ( .A(n10139), .B(n10140), .Z(n10035) );
  AND U9996 ( .A(n160), .B(n10141), .Z(n10140) );
  XNOR U9997 ( .A(n10142), .B(n10143), .Z(n160) );
  AND U9998 ( .A(n10144), .B(n10145), .Z(n10143) );
  XOR U9999 ( .A(n10142), .B(n10045), .Z(n10145) );
  XNOR U10000 ( .A(n10142), .B(n9999), .Z(n10144) );
  XOR U10001 ( .A(n10146), .B(n10147), .Z(n10142) );
  AND U10002 ( .A(n10148), .B(n10149), .Z(n10147) );
  XOR U10003 ( .A(n10146), .B(n10009), .Z(n10148) );
  XOR U10004 ( .A(n10150), .B(n10151), .Z(n9988) );
  AND U10005 ( .A(n164), .B(n10141), .Z(n10151) );
  XNOR U10006 ( .A(n10139), .B(n10150), .Z(n10141) );
  XNOR U10007 ( .A(n10152), .B(n10153), .Z(n164) );
  AND U10008 ( .A(n10154), .B(n10155), .Z(n10153) );
  XNOR U10009 ( .A(n10156), .B(n10152), .Z(n10155) );
  IV U10010 ( .A(n10045), .Z(n10156) );
  XNOR U10011 ( .A(n10157), .B(n10158), .Z(n10045) );
  AND U10012 ( .A(n167), .B(n10159), .Z(n10158) );
  XNOR U10013 ( .A(n10157), .B(n10160), .Z(n10159) );
  XNOR U10014 ( .A(n9999), .B(n10152), .Z(n10154) );
  XOR U10015 ( .A(n10161), .B(n10162), .Z(n9999) );
  AND U10016 ( .A(n175), .B(n10163), .Z(n10162) );
  XOR U10017 ( .A(n10146), .B(n10164), .Z(n10152) );
  AND U10018 ( .A(n10165), .B(n10149), .Z(n10164) );
  XNOR U10019 ( .A(n10058), .B(n10146), .Z(n10149) );
  XNOR U10020 ( .A(n10166), .B(n10167), .Z(n10058) );
  AND U10021 ( .A(n167), .B(n10168), .Z(n10167) );
  XOR U10022 ( .A(n10169), .B(n10166), .Z(n10168) );
  XNOR U10023 ( .A(n10170), .B(n10146), .Z(n10165) );
  IV U10024 ( .A(n10009), .Z(n10170) );
  XOR U10025 ( .A(n10171), .B(n10172), .Z(n10009) );
  AND U10026 ( .A(n175), .B(n10173), .Z(n10172) );
  XOR U10027 ( .A(n10174), .B(n10175), .Z(n10146) );
  AND U10028 ( .A(n10176), .B(n10177), .Z(n10175) );
  XNOR U10029 ( .A(n10083), .B(n10174), .Z(n10177) );
  XNOR U10030 ( .A(n10178), .B(n10179), .Z(n10083) );
  AND U10031 ( .A(n167), .B(n10180), .Z(n10179) );
  XNOR U10032 ( .A(n10181), .B(n10178), .Z(n10180) );
  XOR U10033 ( .A(n10174), .B(n10020), .Z(n10176) );
  XOR U10034 ( .A(n10182), .B(n10183), .Z(n10020) );
  AND U10035 ( .A(n175), .B(n10184), .Z(n10183) );
  XOR U10036 ( .A(n10185), .B(n10186), .Z(n10174) );
  AND U10037 ( .A(n10187), .B(n10188), .Z(n10186) );
  XNOR U10038 ( .A(n10185), .B(n10129), .Z(n10188) );
  XNOR U10039 ( .A(n10189), .B(n10190), .Z(n10129) );
  AND U10040 ( .A(n167), .B(n10191), .Z(n10190) );
  XOR U10041 ( .A(n10192), .B(n10189), .Z(n10191) );
  XNOR U10042 ( .A(n10193), .B(n10185), .Z(n10187) );
  IV U10043 ( .A(n10032), .Z(n10193) );
  XOR U10044 ( .A(n10194), .B(n10195), .Z(n10032) );
  AND U10045 ( .A(n175), .B(n10196), .Z(n10195) );
  AND U10046 ( .A(n10150), .B(n10139), .Z(n10185) );
  XNOR U10047 ( .A(n10197), .B(n10198), .Z(n10139) );
  AND U10048 ( .A(n167), .B(n10199), .Z(n10198) );
  XNOR U10049 ( .A(n10200), .B(n10197), .Z(n10199) );
  XNOR U10050 ( .A(n10201), .B(n10202), .Z(n167) );
  AND U10051 ( .A(n10203), .B(n10204), .Z(n10202) );
  XOR U10052 ( .A(n10160), .B(n10201), .Z(n10204) );
  AND U10053 ( .A(n10205), .B(n10206), .Z(n10160) );
  XOR U10054 ( .A(n10201), .B(n10157), .Z(n10203) );
  XNOR U10055 ( .A(n10207), .B(n10208), .Z(n10157) );
  AND U10056 ( .A(n171), .B(n10163), .Z(n10208) );
  XOR U10057 ( .A(n10161), .B(n10207), .Z(n10163) );
  XOR U10058 ( .A(n10209), .B(n10210), .Z(n10201) );
  AND U10059 ( .A(n10211), .B(n10212), .Z(n10210) );
  XNOR U10060 ( .A(n10209), .B(n10205), .Z(n10212) );
  IV U10061 ( .A(n10169), .Z(n10205) );
  XOR U10062 ( .A(n10213), .B(n10214), .Z(n10169) );
  XOR U10063 ( .A(n10215), .B(n10206), .Z(n10214) );
  AND U10064 ( .A(n10181), .B(n10216), .Z(n10206) );
  AND U10065 ( .A(n10217), .B(n10218), .Z(n10215) );
  XOR U10066 ( .A(n10219), .B(n10213), .Z(n10217) );
  XNOR U10067 ( .A(n10166), .B(n10209), .Z(n10211) );
  XNOR U10068 ( .A(n10220), .B(n10221), .Z(n10166) );
  AND U10069 ( .A(n171), .B(n10173), .Z(n10221) );
  XOR U10070 ( .A(n10220), .B(n10171), .Z(n10173) );
  XOR U10071 ( .A(n10222), .B(n10223), .Z(n10209) );
  AND U10072 ( .A(n10224), .B(n10225), .Z(n10223) );
  XNOR U10073 ( .A(n10222), .B(n10181), .Z(n10225) );
  XOR U10074 ( .A(n10226), .B(n10218), .Z(n10181) );
  XNOR U10075 ( .A(n10227), .B(n10213), .Z(n10218) );
  XOR U10076 ( .A(n10228), .B(n10229), .Z(n10213) );
  AND U10077 ( .A(n10230), .B(n10231), .Z(n10229) );
  XOR U10078 ( .A(n10232), .B(n10228), .Z(n10230) );
  XNOR U10079 ( .A(n10233), .B(n10234), .Z(n10227) );
  AND U10080 ( .A(n10235), .B(n10236), .Z(n10234) );
  XOR U10081 ( .A(n10233), .B(n10237), .Z(n10235) );
  XNOR U10082 ( .A(n10219), .B(n10216), .Z(n10226) );
  AND U10083 ( .A(n10238), .B(n10239), .Z(n10216) );
  XOR U10084 ( .A(n10240), .B(n10241), .Z(n10219) );
  AND U10085 ( .A(n10242), .B(n10243), .Z(n10241) );
  XOR U10086 ( .A(n10240), .B(n10244), .Z(n10242) );
  XNOR U10087 ( .A(n10178), .B(n10222), .Z(n10224) );
  XNOR U10088 ( .A(n10245), .B(n10246), .Z(n10178) );
  AND U10089 ( .A(n171), .B(n10184), .Z(n10246) );
  XOR U10090 ( .A(n10245), .B(n10182), .Z(n10184) );
  XOR U10091 ( .A(n10247), .B(n10248), .Z(n10222) );
  AND U10092 ( .A(n10249), .B(n10250), .Z(n10248) );
  XNOR U10093 ( .A(n10247), .B(n10238), .Z(n10250) );
  IV U10094 ( .A(n10192), .Z(n10238) );
  XNOR U10095 ( .A(n10251), .B(n10231), .Z(n10192) );
  XNOR U10096 ( .A(n10252), .B(n10237), .Z(n10231) );
  XOR U10097 ( .A(n10253), .B(n10254), .Z(n10237) );
  NOR U10098 ( .A(n10255), .B(n10256), .Z(n10254) );
  XNOR U10099 ( .A(n10253), .B(n10257), .Z(n10255) );
  XNOR U10100 ( .A(n10236), .B(n10228), .Z(n10252) );
  XOR U10101 ( .A(n10258), .B(n10259), .Z(n10228) );
  AND U10102 ( .A(n10260), .B(n10261), .Z(n10259) );
  XNOR U10103 ( .A(n10258), .B(n10262), .Z(n10260) );
  XNOR U10104 ( .A(n10263), .B(n10233), .Z(n10236) );
  XOR U10105 ( .A(n10264), .B(n10265), .Z(n10233) );
  AND U10106 ( .A(n10266), .B(n10267), .Z(n10265) );
  XOR U10107 ( .A(n10264), .B(n10268), .Z(n10266) );
  XNOR U10108 ( .A(n10269), .B(n10270), .Z(n10263) );
  NOR U10109 ( .A(n10271), .B(n10272), .Z(n10270) );
  XOR U10110 ( .A(n10269), .B(n10273), .Z(n10271) );
  XNOR U10111 ( .A(n10232), .B(n10239), .Z(n10251) );
  NOR U10112 ( .A(n10200), .B(n10274), .Z(n10239) );
  XOR U10113 ( .A(n10244), .B(n10243), .Z(n10232) );
  XNOR U10114 ( .A(n10275), .B(n10240), .Z(n10243) );
  XOR U10115 ( .A(n10276), .B(n10277), .Z(n10240) );
  AND U10116 ( .A(n10278), .B(n10279), .Z(n10277) );
  XOR U10117 ( .A(n10276), .B(n10280), .Z(n10278) );
  XNOR U10118 ( .A(n10281), .B(n10282), .Z(n10275) );
  NOR U10119 ( .A(n10283), .B(n10284), .Z(n10282) );
  XNOR U10120 ( .A(n10281), .B(n10285), .Z(n10283) );
  XOR U10121 ( .A(n10286), .B(n10287), .Z(n10244) );
  NOR U10122 ( .A(n10288), .B(n10289), .Z(n10287) );
  XNOR U10123 ( .A(n10286), .B(n10290), .Z(n10288) );
  XNOR U10124 ( .A(n10189), .B(n10247), .Z(n10249) );
  XNOR U10125 ( .A(n10291), .B(n10292), .Z(n10189) );
  AND U10126 ( .A(n171), .B(n10196), .Z(n10292) );
  XOR U10127 ( .A(n10291), .B(n10194), .Z(n10196) );
  AND U10128 ( .A(n10197), .B(n10200), .Z(n10247) );
  XOR U10129 ( .A(n10293), .B(n10274), .Z(n10200) );
  XNOR U10130 ( .A(p_input[1024]), .B(p_input[192]), .Z(n10274) );
  XOR U10131 ( .A(n10262), .B(n10261), .Z(n10293) );
  XNOR U10132 ( .A(n10294), .B(n10268), .Z(n10261) );
  XNOR U10133 ( .A(n10257), .B(n10256), .Z(n10268) );
  XOR U10134 ( .A(n10295), .B(n10253), .Z(n10256) );
  XOR U10135 ( .A(p_input[1034]), .B(p_input[202]), .Z(n10253) );
  XNOR U10136 ( .A(p_input[1035]), .B(p_input[203]), .Z(n10295) );
  XOR U10137 ( .A(p_input[1036]), .B(p_input[204]), .Z(n10257) );
  XNOR U10138 ( .A(n10267), .B(n10258), .Z(n10294) );
  XOR U10139 ( .A(p_input[1025]), .B(p_input[193]), .Z(n10258) );
  XOR U10140 ( .A(n10296), .B(n10273), .Z(n10267) );
  XNOR U10141 ( .A(p_input[1039]), .B(p_input[207]), .Z(n10273) );
  XOR U10142 ( .A(n10264), .B(n10272), .Z(n10296) );
  XOR U10143 ( .A(n10297), .B(n10269), .Z(n10272) );
  XOR U10144 ( .A(p_input[1037]), .B(p_input[205]), .Z(n10269) );
  XNOR U10145 ( .A(p_input[1038]), .B(p_input[206]), .Z(n10297) );
  XOR U10146 ( .A(p_input[1033]), .B(p_input[201]), .Z(n10264) );
  XNOR U10147 ( .A(n10280), .B(n10279), .Z(n10262) );
  XNOR U10148 ( .A(n10298), .B(n10285), .Z(n10279) );
  XOR U10149 ( .A(p_input[1032]), .B(p_input[200]), .Z(n10285) );
  XOR U10150 ( .A(n10276), .B(n10284), .Z(n10298) );
  XOR U10151 ( .A(n10299), .B(n10281), .Z(n10284) );
  XOR U10152 ( .A(p_input[1030]), .B(p_input[198]), .Z(n10281) );
  XNOR U10153 ( .A(p_input[1031]), .B(p_input[199]), .Z(n10299) );
  XOR U10154 ( .A(p_input[1026]), .B(p_input[194]), .Z(n10276) );
  XNOR U10155 ( .A(n10290), .B(n10289), .Z(n10280) );
  XOR U10156 ( .A(n10300), .B(n10286), .Z(n10289) );
  XOR U10157 ( .A(p_input[1027]), .B(p_input[195]), .Z(n10286) );
  XNOR U10158 ( .A(p_input[1028]), .B(p_input[196]), .Z(n10300) );
  XOR U10159 ( .A(p_input[1029]), .B(p_input[197]), .Z(n10290) );
  XNOR U10160 ( .A(n10301), .B(n10302), .Z(n10197) );
  AND U10161 ( .A(n171), .B(n10303), .Z(n10302) );
  XNOR U10162 ( .A(n10304), .B(n10305), .Z(n171) );
  AND U10163 ( .A(n10306), .B(n10307), .Z(n10305) );
  XOR U10164 ( .A(n10304), .B(n10207), .Z(n10307) );
  XNOR U10165 ( .A(n10304), .B(n10161), .Z(n10306) );
  XOR U10166 ( .A(n10308), .B(n10309), .Z(n10304) );
  AND U10167 ( .A(n10310), .B(n10311), .Z(n10309) );
  XOR U10168 ( .A(n10308), .B(n10171), .Z(n10310) );
  XOR U10169 ( .A(n10312), .B(n10313), .Z(n10150) );
  AND U10170 ( .A(n175), .B(n10303), .Z(n10313) );
  XNOR U10171 ( .A(n10301), .B(n10312), .Z(n10303) );
  XNOR U10172 ( .A(n10314), .B(n10315), .Z(n175) );
  AND U10173 ( .A(n10316), .B(n10317), .Z(n10315) );
  XNOR U10174 ( .A(n10318), .B(n10314), .Z(n10317) );
  IV U10175 ( .A(n10207), .Z(n10318) );
  XNOR U10176 ( .A(n10319), .B(n10320), .Z(n10207) );
  AND U10177 ( .A(n178), .B(n10321), .Z(n10320) );
  XNOR U10178 ( .A(n10319), .B(n10322), .Z(n10321) );
  XNOR U10179 ( .A(n10161), .B(n10314), .Z(n10316) );
  XOR U10180 ( .A(n10323), .B(n10324), .Z(n10161) );
  AND U10181 ( .A(n186), .B(n10325), .Z(n10324) );
  XOR U10182 ( .A(n10308), .B(n10326), .Z(n10314) );
  AND U10183 ( .A(n10327), .B(n10311), .Z(n10326) );
  XNOR U10184 ( .A(n10220), .B(n10308), .Z(n10311) );
  XNOR U10185 ( .A(n10328), .B(n10329), .Z(n10220) );
  AND U10186 ( .A(n178), .B(n10330), .Z(n10329) );
  XOR U10187 ( .A(n10331), .B(n10328), .Z(n10330) );
  XNOR U10188 ( .A(n10332), .B(n10308), .Z(n10327) );
  IV U10189 ( .A(n10171), .Z(n10332) );
  XOR U10190 ( .A(n10333), .B(n10334), .Z(n10171) );
  AND U10191 ( .A(n186), .B(n10335), .Z(n10334) );
  XOR U10192 ( .A(n10336), .B(n10337), .Z(n10308) );
  AND U10193 ( .A(n10338), .B(n10339), .Z(n10337) );
  XNOR U10194 ( .A(n10245), .B(n10336), .Z(n10339) );
  XNOR U10195 ( .A(n10340), .B(n10341), .Z(n10245) );
  AND U10196 ( .A(n178), .B(n10342), .Z(n10341) );
  XNOR U10197 ( .A(n10343), .B(n10340), .Z(n10342) );
  XOR U10198 ( .A(n10336), .B(n10182), .Z(n10338) );
  XOR U10199 ( .A(n10344), .B(n10345), .Z(n10182) );
  AND U10200 ( .A(n186), .B(n10346), .Z(n10345) );
  XOR U10201 ( .A(n10347), .B(n10348), .Z(n10336) );
  AND U10202 ( .A(n10349), .B(n10350), .Z(n10348) );
  XNOR U10203 ( .A(n10347), .B(n10291), .Z(n10350) );
  XNOR U10204 ( .A(n10351), .B(n10352), .Z(n10291) );
  AND U10205 ( .A(n178), .B(n10353), .Z(n10352) );
  XOR U10206 ( .A(n10354), .B(n10351), .Z(n10353) );
  XNOR U10207 ( .A(n10355), .B(n10347), .Z(n10349) );
  IV U10208 ( .A(n10194), .Z(n10355) );
  XOR U10209 ( .A(n10356), .B(n10357), .Z(n10194) );
  AND U10210 ( .A(n186), .B(n10358), .Z(n10357) );
  AND U10211 ( .A(n10312), .B(n10301), .Z(n10347) );
  XNOR U10212 ( .A(n10359), .B(n10360), .Z(n10301) );
  AND U10213 ( .A(n178), .B(n10361), .Z(n10360) );
  XNOR U10214 ( .A(n10362), .B(n10359), .Z(n10361) );
  XNOR U10215 ( .A(n10363), .B(n10364), .Z(n178) );
  AND U10216 ( .A(n10365), .B(n10366), .Z(n10364) );
  XOR U10217 ( .A(n10322), .B(n10363), .Z(n10366) );
  AND U10218 ( .A(n10367), .B(n10368), .Z(n10322) );
  XOR U10219 ( .A(n10363), .B(n10319), .Z(n10365) );
  XNOR U10220 ( .A(n10369), .B(n10370), .Z(n10319) );
  AND U10221 ( .A(n182), .B(n10325), .Z(n10370) );
  XOR U10222 ( .A(n10323), .B(n10369), .Z(n10325) );
  XOR U10223 ( .A(n10371), .B(n10372), .Z(n10363) );
  AND U10224 ( .A(n10373), .B(n10374), .Z(n10372) );
  XNOR U10225 ( .A(n10371), .B(n10367), .Z(n10374) );
  IV U10226 ( .A(n10331), .Z(n10367) );
  XOR U10227 ( .A(n10375), .B(n10376), .Z(n10331) );
  XOR U10228 ( .A(n10377), .B(n10368), .Z(n10376) );
  AND U10229 ( .A(n10343), .B(n10378), .Z(n10368) );
  AND U10230 ( .A(n10379), .B(n10380), .Z(n10377) );
  XOR U10231 ( .A(n10381), .B(n10375), .Z(n10379) );
  XNOR U10232 ( .A(n10328), .B(n10371), .Z(n10373) );
  XNOR U10233 ( .A(n10382), .B(n10383), .Z(n10328) );
  AND U10234 ( .A(n182), .B(n10335), .Z(n10383) );
  XOR U10235 ( .A(n10382), .B(n10333), .Z(n10335) );
  XOR U10236 ( .A(n10384), .B(n10385), .Z(n10371) );
  AND U10237 ( .A(n10386), .B(n10387), .Z(n10385) );
  XNOR U10238 ( .A(n10384), .B(n10343), .Z(n10387) );
  XOR U10239 ( .A(n10388), .B(n10380), .Z(n10343) );
  XNOR U10240 ( .A(n10389), .B(n10375), .Z(n10380) );
  XOR U10241 ( .A(n10390), .B(n10391), .Z(n10375) );
  AND U10242 ( .A(n10392), .B(n10393), .Z(n10391) );
  XOR U10243 ( .A(n10394), .B(n10390), .Z(n10392) );
  XNOR U10244 ( .A(n10395), .B(n10396), .Z(n10389) );
  AND U10245 ( .A(n10397), .B(n10398), .Z(n10396) );
  XOR U10246 ( .A(n10395), .B(n10399), .Z(n10397) );
  XNOR U10247 ( .A(n10381), .B(n10378), .Z(n10388) );
  AND U10248 ( .A(n10400), .B(n10401), .Z(n10378) );
  XOR U10249 ( .A(n10402), .B(n10403), .Z(n10381) );
  AND U10250 ( .A(n10404), .B(n10405), .Z(n10403) );
  XOR U10251 ( .A(n10402), .B(n10406), .Z(n10404) );
  XNOR U10252 ( .A(n10340), .B(n10384), .Z(n10386) );
  XNOR U10253 ( .A(n10407), .B(n10408), .Z(n10340) );
  AND U10254 ( .A(n182), .B(n10346), .Z(n10408) );
  XOR U10255 ( .A(n10407), .B(n10344), .Z(n10346) );
  XOR U10256 ( .A(n10409), .B(n10410), .Z(n10384) );
  AND U10257 ( .A(n10411), .B(n10412), .Z(n10410) );
  XNOR U10258 ( .A(n10409), .B(n10400), .Z(n10412) );
  IV U10259 ( .A(n10354), .Z(n10400) );
  XNOR U10260 ( .A(n10413), .B(n10393), .Z(n10354) );
  XNOR U10261 ( .A(n10414), .B(n10399), .Z(n10393) );
  XOR U10262 ( .A(n10415), .B(n10416), .Z(n10399) );
  NOR U10263 ( .A(n10417), .B(n10418), .Z(n10416) );
  XNOR U10264 ( .A(n10415), .B(n10419), .Z(n10417) );
  XNOR U10265 ( .A(n10398), .B(n10390), .Z(n10414) );
  XOR U10266 ( .A(n10420), .B(n10421), .Z(n10390) );
  AND U10267 ( .A(n10422), .B(n10423), .Z(n10421) );
  XNOR U10268 ( .A(n10420), .B(n10424), .Z(n10422) );
  XNOR U10269 ( .A(n10425), .B(n10395), .Z(n10398) );
  XOR U10270 ( .A(n10426), .B(n10427), .Z(n10395) );
  AND U10271 ( .A(n10428), .B(n10429), .Z(n10427) );
  XOR U10272 ( .A(n10426), .B(n10430), .Z(n10428) );
  XNOR U10273 ( .A(n10431), .B(n10432), .Z(n10425) );
  NOR U10274 ( .A(n10433), .B(n10434), .Z(n10432) );
  XOR U10275 ( .A(n10431), .B(n10435), .Z(n10433) );
  XNOR U10276 ( .A(n10394), .B(n10401), .Z(n10413) );
  NOR U10277 ( .A(n10362), .B(n10436), .Z(n10401) );
  XOR U10278 ( .A(n10406), .B(n10405), .Z(n10394) );
  XNOR U10279 ( .A(n10437), .B(n10402), .Z(n10405) );
  XOR U10280 ( .A(n10438), .B(n10439), .Z(n10402) );
  AND U10281 ( .A(n10440), .B(n10441), .Z(n10439) );
  XOR U10282 ( .A(n10438), .B(n10442), .Z(n10440) );
  XNOR U10283 ( .A(n10443), .B(n10444), .Z(n10437) );
  NOR U10284 ( .A(n10445), .B(n10446), .Z(n10444) );
  XNOR U10285 ( .A(n10443), .B(n10447), .Z(n10445) );
  XOR U10286 ( .A(n10448), .B(n10449), .Z(n10406) );
  NOR U10287 ( .A(n10450), .B(n10451), .Z(n10449) );
  XNOR U10288 ( .A(n10448), .B(n10452), .Z(n10450) );
  XNOR U10289 ( .A(n10351), .B(n10409), .Z(n10411) );
  XNOR U10290 ( .A(n10453), .B(n10454), .Z(n10351) );
  AND U10291 ( .A(n182), .B(n10358), .Z(n10454) );
  XOR U10292 ( .A(n10453), .B(n10356), .Z(n10358) );
  AND U10293 ( .A(n10359), .B(n10362), .Z(n10409) );
  XOR U10294 ( .A(n10455), .B(n10436), .Z(n10362) );
  XNOR U10295 ( .A(p_input[1024]), .B(p_input[208]), .Z(n10436) );
  XOR U10296 ( .A(n10424), .B(n10423), .Z(n10455) );
  XNOR U10297 ( .A(n10456), .B(n10430), .Z(n10423) );
  XNOR U10298 ( .A(n10419), .B(n10418), .Z(n10430) );
  XOR U10299 ( .A(n10457), .B(n10415), .Z(n10418) );
  XOR U10300 ( .A(p_input[1034]), .B(p_input[218]), .Z(n10415) );
  XNOR U10301 ( .A(p_input[1035]), .B(p_input[219]), .Z(n10457) );
  XOR U10302 ( .A(p_input[1036]), .B(p_input[220]), .Z(n10419) );
  XNOR U10303 ( .A(n10429), .B(n10420), .Z(n10456) );
  XOR U10304 ( .A(p_input[1025]), .B(p_input[209]), .Z(n10420) );
  XOR U10305 ( .A(n10458), .B(n10435), .Z(n10429) );
  XNOR U10306 ( .A(p_input[1039]), .B(p_input[223]), .Z(n10435) );
  XOR U10307 ( .A(n10426), .B(n10434), .Z(n10458) );
  XOR U10308 ( .A(n10459), .B(n10431), .Z(n10434) );
  XOR U10309 ( .A(p_input[1037]), .B(p_input[221]), .Z(n10431) );
  XNOR U10310 ( .A(p_input[1038]), .B(p_input[222]), .Z(n10459) );
  XOR U10311 ( .A(p_input[1033]), .B(p_input[217]), .Z(n10426) );
  XNOR U10312 ( .A(n10442), .B(n10441), .Z(n10424) );
  XNOR U10313 ( .A(n10460), .B(n10447), .Z(n10441) );
  XOR U10314 ( .A(p_input[1032]), .B(p_input[216]), .Z(n10447) );
  XOR U10315 ( .A(n10438), .B(n10446), .Z(n10460) );
  XOR U10316 ( .A(n10461), .B(n10443), .Z(n10446) );
  XOR U10317 ( .A(p_input[1030]), .B(p_input[214]), .Z(n10443) );
  XNOR U10318 ( .A(p_input[1031]), .B(p_input[215]), .Z(n10461) );
  XOR U10319 ( .A(p_input[1026]), .B(p_input[210]), .Z(n10438) );
  XNOR U10320 ( .A(n10452), .B(n10451), .Z(n10442) );
  XOR U10321 ( .A(n10462), .B(n10448), .Z(n10451) );
  XOR U10322 ( .A(p_input[1027]), .B(p_input[211]), .Z(n10448) );
  XNOR U10323 ( .A(p_input[1028]), .B(p_input[212]), .Z(n10462) );
  XOR U10324 ( .A(p_input[1029]), .B(p_input[213]), .Z(n10452) );
  XNOR U10325 ( .A(n10463), .B(n10464), .Z(n10359) );
  AND U10326 ( .A(n182), .B(n10465), .Z(n10464) );
  XNOR U10327 ( .A(n10466), .B(n10467), .Z(n182) );
  AND U10328 ( .A(n10468), .B(n10469), .Z(n10467) );
  XOR U10329 ( .A(n10466), .B(n10369), .Z(n10469) );
  XNOR U10330 ( .A(n10466), .B(n10323), .Z(n10468) );
  XOR U10331 ( .A(n10470), .B(n10471), .Z(n10466) );
  AND U10332 ( .A(n10472), .B(n10473), .Z(n10471) );
  XOR U10333 ( .A(n10470), .B(n10333), .Z(n10472) );
  XOR U10334 ( .A(n10474), .B(n10475), .Z(n10312) );
  AND U10335 ( .A(n186), .B(n10465), .Z(n10475) );
  XNOR U10336 ( .A(n10463), .B(n10474), .Z(n10465) );
  XNOR U10337 ( .A(n10476), .B(n10477), .Z(n186) );
  AND U10338 ( .A(n10478), .B(n10479), .Z(n10477) );
  XNOR U10339 ( .A(n10480), .B(n10476), .Z(n10479) );
  IV U10340 ( .A(n10369), .Z(n10480) );
  XNOR U10341 ( .A(n10481), .B(n10482), .Z(n10369) );
  AND U10342 ( .A(n189), .B(n10483), .Z(n10482) );
  XNOR U10343 ( .A(n10481), .B(n10484), .Z(n10483) );
  XNOR U10344 ( .A(n10323), .B(n10476), .Z(n10478) );
  XOR U10345 ( .A(n10485), .B(n10486), .Z(n10323) );
  AND U10346 ( .A(n197), .B(n10487), .Z(n10486) );
  XOR U10347 ( .A(n10470), .B(n10488), .Z(n10476) );
  AND U10348 ( .A(n10489), .B(n10473), .Z(n10488) );
  XNOR U10349 ( .A(n10382), .B(n10470), .Z(n10473) );
  XNOR U10350 ( .A(n10490), .B(n10491), .Z(n10382) );
  AND U10351 ( .A(n189), .B(n10492), .Z(n10491) );
  XOR U10352 ( .A(n10493), .B(n10490), .Z(n10492) );
  XNOR U10353 ( .A(n10494), .B(n10470), .Z(n10489) );
  IV U10354 ( .A(n10333), .Z(n10494) );
  XOR U10355 ( .A(n10495), .B(n10496), .Z(n10333) );
  AND U10356 ( .A(n197), .B(n10497), .Z(n10496) );
  XOR U10357 ( .A(n10498), .B(n10499), .Z(n10470) );
  AND U10358 ( .A(n10500), .B(n10501), .Z(n10499) );
  XNOR U10359 ( .A(n10407), .B(n10498), .Z(n10501) );
  XNOR U10360 ( .A(n10502), .B(n10503), .Z(n10407) );
  AND U10361 ( .A(n189), .B(n10504), .Z(n10503) );
  XNOR U10362 ( .A(n10505), .B(n10502), .Z(n10504) );
  XOR U10363 ( .A(n10498), .B(n10344), .Z(n10500) );
  XOR U10364 ( .A(n10506), .B(n10507), .Z(n10344) );
  AND U10365 ( .A(n197), .B(n10508), .Z(n10507) );
  XOR U10366 ( .A(n10509), .B(n10510), .Z(n10498) );
  AND U10367 ( .A(n10511), .B(n10512), .Z(n10510) );
  XNOR U10368 ( .A(n10509), .B(n10453), .Z(n10512) );
  XNOR U10369 ( .A(n10513), .B(n10514), .Z(n10453) );
  AND U10370 ( .A(n189), .B(n10515), .Z(n10514) );
  XOR U10371 ( .A(n10516), .B(n10513), .Z(n10515) );
  XNOR U10372 ( .A(n10517), .B(n10509), .Z(n10511) );
  IV U10373 ( .A(n10356), .Z(n10517) );
  XOR U10374 ( .A(n10518), .B(n10519), .Z(n10356) );
  AND U10375 ( .A(n197), .B(n10520), .Z(n10519) );
  AND U10376 ( .A(n10474), .B(n10463), .Z(n10509) );
  XNOR U10377 ( .A(n10521), .B(n10522), .Z(n10463) );
  AND U10378 ( .A(n189), .B(n10523), .Z(n10522) );
  XNOR U10379 ( .A(n10524), .B(n10521), .Z(n10523) );
  XNOR U10380 ( .A(n10525), .B(n10526), .Z(n189) );
  AND U10381 ( .A(n10527), .B(n10528), .Z(n10526) );
  XOR U10382 ( .A(n10484), .B(n10525), .Z(n10528) );
  AND U10383 ( .A(n10529), .B(n10530), .Z(n10484) );
  XOR U10384 ( .A(n10525), .B(n10481), .Z(n10527) );
  XNOR U10385 ( .A(n10531), .B(n10532), .Z(n10481) );
  AND U10386 ( .A(n193), .B(n10487), .Z(n10532) );
  XOR U10387 ( .A(n10485), .B(n10531), .Z(n10487) );
  XOR U10388 ( .A(n10533), .B(n10534), .Z(n10525) );
  AND U10389 ( .A(n10535), .B(n10536), .Z(n10534) );
  XNOR U10390 ( .A(n10533), .B(n10529), .Z(n10536) );
  IV U10391 ( .A(n10493), .Z(n10529) );
  XOR U10392 ( .A(n10537), .B(n10538), .Z(n10493) );
  XOR U10393 ( .A(n10539), .B(n10530), .Z(n10538) );
  AND U10394 ( .A(n10505), .B(n10540), .Z(n10530) );
  AND U10395 ( .A(n10541), .B(n10542), .Z(n10539) );
  XOR U10396 ( .A(n10543), .B(n10537), .Z(n10541) );
  XNOR U10397 ( .A(n10490), .B(n10533), .Z(n10535) );
  XNOR U10398 ( .A(n10544), .B(n10545), .Z(n10490) );
  AND U10399 ( .A(n193), .B(n10497), .Z(n10545) );
  XOR U10400 ( .A(n10544), .B(n10495), .Z(n10497) );
  XOR U10401 ( .A(n10546), .B(n10547), .Z(n10533) );
  AND U10402 ( .A(n10548), .B(n10549), .Z(n10547) );
  XNOR U10403 ( .A(n10546), .B(n10505), .Z(n10549) );
  XOR U10404 ( .A(n10550), .B(n10542), .Z(n10505) );
  XNOR U10405 ( .A(n10551), .B(n10537), .Z(n10542) );
  XOR U10406 ( .A(n10552), .B(n10553), .Z(n10537) );
  AND U10407 ( .A(n10554), .B(n10555), .Z(n10553) );
  XOR U10408 ( .A(n10556), .B(n10552), .Z(n10554) );
  XNOR U10409 ( .A(n10557), .B(n10558), .Z(n10551) );
  AND U10410 ( .A(n10559), .B(n10560), .Z(n10558) );
  XOR U10411 ( .A(n10557), .B(n10561), .Z(n10559) );
  XNOR U10412 ( .A(n10543), .B(n10540), .Z(n10550) );
  AND U10413 ( .A(n10562), .B(n10563), .Z(n10540) );
  XOR U10414 ( .A(n10564), .B(n10565), .Z(n10543) );
  AND U10415 ( .A(n10566), .B(n10567), .Z(n10565) );
  XOR U10416 ( .A(n10564), .B(n10568), .Z(n10566) );
  XNOR U10417 ( .A(n10502), .B(n10546), .Z(n10548) );
  XNOR U10418 ( .A(n10569), .B(n10570), .Z(n10502) );
  AND U10419 ( .A(n193), .B(n10508), .Z(n10570) );
  XOR U10420 ( .A(n10569), .B(n10506), .Z(n10508) );
  XOR U10421 ( .A(n10571), .B(n10572), .Z(n10546) );
  AND U10422 ( .A(n10573), .B(n10574), .Z(n10572) );
  XNOR U10423 ( .A(n10571), .B(n10562), .Z(n10574) );
  IV U10424 ( .A(n10516), .Z(n10562) );
  XNOR U10425 ( .A(n10575), .B(n10555), .Z(n10516) );
  XNOR U10426 ( .A(n10576), .B(n10561), .Z(n10555) );
  XOR U10427 ( .A(n10577), .B(n10578), .Z(n10561) );
  NOR U10428 ( .A(n10579), .B(n10580), .Z(n10578) );
  XNOR U10429 ( .A(n10577), .B(n10581), .Z(n10579) );
  XNOR U10430 ( .A(n10560), .B(n10552), .Z(n10576) );
  XOR U10431 ( .A(n10582), .B(n10583), .Z(n10552) );
  AND U10432 ( .A(n10584), .B(n10585), .Z(n10583) );
  XNOR U10433 ( .A(n10582), .B(n10586), .Z(n10584) );
  XNOR U10434 ( .A(n10587), .B(n10557), .Z(n10560) );
  XOR U10435 ( .A(n10588), .B(n10589), .Z(n10557) );
  AND U10436 ( .A(n10590), .B(n10591), .Z(n10589) );
  XOR U10437 ( .A(n10588), .B(n10592), .Z(n10590) );
  XNOR U10438 ( .A(n10593), .B(n10594), .Z(n10587) );
  NOR U10439 ( .A(n10595), .B(n10596), .Z(n10594) );
  XOR U10440 ( .A(n10593), .B(n10597), .Z(n10595) );
  XNOR U10441 ( .A(n10556), .B(n10563), .Z(n10575) );
  NOR U10442 ( .A(n10524), .B(n10598), .Z(n10563) );
  XOR U10443 ( .A(n10568), .B(n10567), .Z(n10556) );
  XNOR U10444 ( .A(n10599), .B(n10564), .Z(n10567) );
  XOR U10445 ( .A(n10600), .B(n10601), .Z(n10564) );
  AND U10446 ( .A(n10602), .B(n10603), .Z(n10601) );
  XOR U10447 ( .A(n10600), .B(n10604), .Z(n10602) );
  XNOR U10448 ( .A(n10605), .B(n10606), .Z(n10599) );
  NOR U10449 ( .A(n10607), .B(n10608), .Z(n10606) );
  XNOR U10450 ( .A(n10605), .B(n10609), .Z(n10607) );
  XOR U10451 ( .A(n10610), .B(n10611), .Z(n10568) );
  NOR U10452 ( .A(n10612), .B(n10613), .Z(n10611) );
  XNOR U10453 ( .A(n10610), .B(n10614), .Z(n10612) );
  XNOR U10454 ( .A(n10513), .B(n10571), .Z(n10573) );
  XNOR U10455 ( .A(n10615), .B(n10616), .Z(n10513) );
  AND U10456 ( .A(n193), .B(n10520), .Z(n10616) );
  XOR U10457 ( .A(n10615), .B(n10518), .Z(n10520) );
  AND U10458 ( .A(n10521), .B(n10524), .Z(n10571) );
  XOR U10459 ( .A(n10617), .B(n10598), .Z(n10524) );
  XNOR U10460 ( .A(p_input[1024]), .B(p_input[224]), .Z(n10598) );
  XOR U10461 ( .A(n10586), .B(n10585), .Z(n10617) );
  XNOR U10462 ( .A(n10618), .B(n10592), .Z(n10585) );
  XNOR U10463 ( .A(n10581), .B(n10580), .Z(n10592) );
  XOR U10464 ( .A(n10619), .B(n10577), .Z(n10580) );
  XOR U10465 ( .A(p_input[1034]), .B(p_input[234]), .Z(n10577) );
  XNOR U10466 ( .A(p_input[1035]), .B(p_input[235]), .Z(n10619) );
  XOR U10467 ( .A(p_input[1036]), .B(p_input[236]), .Z(n10581) );
  XNOR U10468 ( .A(n10591), .B(n10582), .Z(n10618) );
  XOR U10469 ( .A(p_input[1025]), .B(p_input[225]), .Z(n10582) );
  XOR U10470 ( .A(n10620), .B(n10597), .Z(n10591) );
  XNOR U10471 ( .A(p_input[1039]), .B(p_input[239]), .Z(n10597) );
  XOR U10472 ( .A(n10588), .B(n10596), .Z(n10620) );
  XOR U10473 ( .A(n10621), .B(n10593), .Z(n10596) );
  XOR U10474 ( .A(p_input[1037]), .B(p_input[237]), .Z(n10593) );
  XNOR U10475 ( .A(p_input[1038]), .B(p_input[238]), .Z(n10621) );
  XOR U10476 ( .A(p_input[1033]), .B(p_input[233]), .Z(n10588) );
  XNOR U10477 ( .A(n10604), .B(n10603), .Z(n10586) );
  XNOR U10478 ( .A(n10622), .B(n10609), .Z(n10603) );
  XOR U10479 ( .A(p_input[1032]), .B(p_input[232]), .Z(n10609) );
  XOR U10480 ( .A(n10600), .B(n10608), .Z(n10622) );
  XOR U10481 ( .A(n10623), .B(n10605), .Z(n10608) );
  XOR U10482 ( .A(p_input[1030]), .B(p_input[230]), .Z(n10605) );
  XNOR U10483 ( .A(p_input[1031]), .B(p_input[231]), .Z(n10623) );
  XOR U10484 ( .A(p_input[1026]), .B(p_input[226]), .Z(n10600) );
  XNOR U10485 ( .A(n10614), .B(n10613), .Z(n10604) );
  XOR U10486 ( .A(n10624), .B(n10610), .Z(n10613) );
  XOR U10487 ( .A(p_input[1027]), .B(p_input[227]), .Z(n10610) );
  XNOR U10488 ( .A(p_input[1028]), .B(p_input[228]), .Z(n10624) );
  XOR U10489 ( .A(p_input[1029]), .B(p_input[229]), .Z(n10614) );
  XNOR U10490 ( .A(n10625), .B(n10626), .Z(n10521) );
  AND U10491 ( .A(n193), .B(n10627), .Z(n10626) );
  XNOR U10492 ( .A(n10628), .B(n10629), .Z(n193) );
  AND U10493 ( .A(n10630), .B(n10631), .Z(n10629) );
  XOR U10494 ( .A(n10628), .B(n10531), .Z(n10631) );
  XNOR U10495 ( .A(n10628), .B(n10485), .Z(n10630) );
  XOR U10496 ( .A(n10632), .B(n10633), .Z(n10628) );
  AND U10497 ( .A(n10634), .B(n10635), .Z(n10633) );
  XOR U10498 ( .A(n10632), .B(n10495), .Z(n10634) );
  XOR U10499 ( .A(n10636), .B(n10637), .Z(n10474) );
  AND U10500 ( .A(n197), .B(n10627), .Z(n10637) );
  XNOR U10501 ( .A(n10625), .B(n10636), .Z(n10627) );
  XNOR U10502 ( .A(n10638), .B(n10639), .Z(n197) );
  AND U10503 ( .A(n10640), .B(n10641), .Z(n10639) );
  XNOR U10504 ( .A(n10642), .B(n10638), .Z(n10641) );
  IV U10505 ( .A(n10531), .Z(n10642) );
  XNOR U10506 ( .A(n10643), .B(n10644), .Z(n10531) );
  AND U10507 ( .A(n200), .B(n10645), .Z(n10644) );
  XNOR U10508 ( .A(n10643), .B(n10646), .Z(n10645) );
  XNOR U10509 ( .A(n10485), .B(n10638), .Z(n10640) );
  XOR U10510 ( .A(n10647), .B(n10648), .Z(n10485) );
  AND U10511 ( .A(n208), .B(n10649), .Z(n10648) );
  XOR U10512 ( .A(n10632), .B(n10650), .Z(n10638) );
  AND U10513 ( .A(n10651), .B(n10635), .Z(n10650) );
  XNOR U10514 ( .A(n10544), .B(n10632), .Z(n10635) );
  XNOR U10515 ( .A(n10652), .B(n10653), .Z(n10544) );
  AND U10516 ( .A(n200), .B(n10654), .Z(n10653) );
  XOR U10517 ( .A(n10655), .B(n10652), .Z(n10654) );
  XNOR U10518 ( .A(n10656), .B(n10632), .Z(n10651) );
  IV U10519 ( .A(n10495), .Z(n10656) );
  XOR U10520 ( .A(n10657), .B(n10658), .Z(n10495) );
  AND U10521 ( .A(n208), .B(n10659), .Z(n10658) );
  XOR U10522 ( .A(n10660), .B(n10661), .Z(n10632) );
  AND U10523 ( .A(n10662), .B(n10663), .Z(n10661) );
  XNOR U10524 ( .A(n10569), .B(n10660), .Z(n10663) );
  XNOR U10525 ( .A(n10664), .B(n10665), .Z(n10569) );
  AND U10526 ( .A(n200), .B(n10666), .Z(n10665) );
  XNOR U10527 ( .A(n10667), .B(n10664), .Z(n10666) );
  XOR U10528 ( .A(n10660), .B(n10506), .Z(n10662) );
  XOR U10529 ( .A(n10668), .B(n10669), .Z(n10506) );
  AND U10530 ( .A(n208), .B(n10670), .Z(n10669) );
  XOR U10531 ( .A(n10671), .B(n10672), .Z(n10660) );
  AND U10532 ( .A(n10673), .B(n10674), .Z(n10672) );
  XNOR U10533 ( .A(n10671), .B(n10615), .Z(n10674) );
  XNOR U10534 ( .A(n10675), .B(n10676), .Z(n10615) );
  AND U10535 ( .A(n200), .B(n10677), .Z(n10676) );
  XOR U10536 ( .A(n10678), .B(n10675), .Z(n10677) );
  XNOR U10537 ( .A(n10679), .B(n10671), .Z(n10673) );
  IV U10538 ( .A(n10518), .Z(n10679) );
  XOR U10539 ( .A(n10680), .B(n10681), .Z(n10518) );
  AND U10540 ( .A(n208), .B(n10682), .Z(n10681) );
  AND U10541 ( .A(n10636), .B(n10625), .Z(n10671) );
  XNOR U10542 ( .A(n10683), .B(n10684), .Z(n10625) );
  AND U10543 ( .A(n200), .B(n10685), .Z(n10684) );
  XNOR U10544 ( .A(n10686), .B(n10683), .Z(n10685) );
  XNOR U10545 ( .A(n10687), .B(n10688), .Z(n200) );
  AND U10546 ( .A(n10689), .B(n10690), .Z(n10688) );
  XOR U10547 ( .A(n10646), .B(n10687), .Z(n10690) );
  AND U10548 ( .A(n10691), .B(n10692), .Z(n10646) );
  XOR U10549 ( .A(n10687), .B(n10643), .Z(n10689) );
  XNOR U10550 ( .A(n10693), .B(n10694), .Z(n10643) );
  AND U10551 ( .A(n204), .B(n10649), .Z(n10694) );
  XOR U10552 ( .A(n10647), .B(n10693), .Z(n10649) );
  XOR U10553 ( .A(n10695), .B(n10696), .Z(n10687) );
  AND U10554 ( .A(n10697), .B(n10698), .Z(n10696) );
  XNOR U10555 ( .A(n10695), .B(n10691), .Z(n10698) );
  IV U10556 ( .A(n10655), .Z(n10691) );
  XOR U10557 ( .A(n10699), .B(n10700), .Z(n10655) );
  XOR U10558 ( .A(n10701), .B(n10692), .Z(n10700) );
  AND U10559 ( .A(n10667), .B(n10702), .Z(n10692) );
  AND U10560 ( .A(n10703), .B(n10704), .Z(n10701) );
  XOR U10561 ( .A(n10705), .B(n10699), .Z(n10703) );
  XNOR U10562 ( .A(n10652), .B(n10695), .Z(n10697) );
  XNOR U10563 ( .A(n10706), .B(n10707), .Z(n10652) );
  AND U10564 ( .A(n204), .B(n10659), .Z(n10707) );
  XOR U10565 ( .A(n10706), .B(n10657), .Z(n10659) );
  XOR U10566 ( .A(n10708), .B(n10709), .Z(n10695) );
  AND U10567 ( .A(n10710), .B(n10711), .Z(n10709) );
  XNOR U10568 ( .A(n10708), .B(n10667), .Z(n10711) );
  XOR U10569 ( .A(n10712), .B(n10704), .Z(n10667) );
  XNOR U10570 ( .A(n10713), .B(n10699), .Z(n10704) );
  XOR U10571 ( .A(n10714), .B(n10715), .Z(n10699) );
  AND U10572 ( .A(n10716), .B(n10717), .Z(n10715) );
  XOR U10573 ( .A(n10718), .B(n10714), .Z(n10716) );
  XNOR U10574 ( .A(n10719), .B(n10720), .Z(n10713) );
  AND U10575 ( .A(n10721), .B(n10722), .Z(n10720) );
  XOR U10576 ( .A(n10719), .B(n10723), .Z(n10721) );
  XNOR U10577 ( .A(n10705), .B(n10702), .Z(n10712) );
  AND U10578 ( .A(n10724), .B(n10725), .Z(n10702) );
  XOR U10579 ( .A(n10726), .B(n10727), .Z(n10705) );
  AND U10580 ( .A(n10728), .B(n10729), .Z(n10727) );
  XOR U10581 ( .A(n10726), .B(n10730), .Z(n10728) );
  XNOR U10582 ( .A(n10664), .B(n10708), .Z(n10710) );
  XNOR U10583 ( .A(n10731), .B(n10732), .Z(n10664) );
  AND U10584 ( .A(n204), .B(n10670), .Z(n10732) );
  XOR U10585 ( .A(n10731), .B(n10668), .Z(n10670) );
  XOR U10586 ( .A(n10733), .B(n10734), .Z(n10708) );
  AND U10587 ( .A(n10735), .B(n10736), .Z(n10734) );
  XNOR U10588 ( .A(n10733), .B(n10724), .Z(n10736) );
  IV U10589 ( .A(n10678), .Z(n10724) );
  XNOR U10590 ( .A(n10737), .B(n10717), .Z(n10678) );
  XNOR U10591 ( .A(n10738), .B(n10723), .Z(n10717) );
  XOR U10592 ( .A(n10739), .B(n10740), .Z(n10723) );
  NOR U10593 ( .A(n10741), .B(n10742), .Z(n10740) );
  XNOR U10594 ( .A(n10739), .B(n10743), .Z(n10741) );
  XNOR U10595 ( .A(n10722), .B(n10714), .Z(n10738) );
  XOR U10596 ( .A(n10744), .B(n10745), .Z(n10714) );
  AND U10597 ( .A(n10746), .B(n10747), .Z(n10745) );
  XNOR U10598 ( .A(n10744), .B(n10748), .Z(n10746) );
  XNOR U10599 ( .A(n10749), .B(n10719), .Z(n10722) );
  XOR U10600 ( .A(n10750), .B(n10751), .Z(n10719) );
  AND U10601 ( .A(n10752), .B(n10753), .Z(n10751) );
  XOR U10602 ( .A(n10750), .B(n10754), .Z(n10752) );
  XNOR U10603 ( .A(n10755), .B(n10756), .Z(n10749) );
  NOR U10604 ( .A(n10757), .B(n10758), .Z(n10756) );
  XOR U10605 ( .A(n10755), .B(n10759), .Z(n10757) );
  XNOR U10606 ( .A(n10718), .B(n10725), .Z(n10737) );
  NOR U10607 ( .A(n10686), .B(n10760), .Z(n10725) );
  XOR U10608 ( .A(n10730), .B(n10729), .Z(n10718) );
  XNOR U10609 ( .A(n10761), .B(n10726), .Z(n10729) );
  XOR U10610 ( .A(n10762), .B(n10763), .Z(n10726) );
  AND U10611 ( .A(n10764), .B(n10765), .Z(n10763) );
  XOR U10612 ( .A(n10762), .B(n10766), .Z(n10764) );
  XNOR U10613 ( .A(n10767), .B(n10768), .Z(n10761) );
  NOR U10614 ( .A(n10769), .B(n10770), .Z(n10768) );
  XNOR U10615 ( .A(n10767), .B(n10771), .Z(n10769) );
  XOR U10616 ( .A(n10772), .B(n10773), .Z(n10730) );
  NOR U10617 ( .A(n10774), .B(n10775), .Z(n10773) );
  XNOR U10618 ( .A(n10772), .B(n10776), .Z(n10774) );
  XNOR U10619 ( .A(n10675), .B(n10733), .Z(n10735) );
  XNOR U10620 ( .A(n10777), .B(n10778), .Z(n10675) );
  AND U10621 ( .A(n204), .B(n10682), .Z(n10778) );
  XOR U10622 ( .A(n10777), .B(n10680), .Z(n10682) );
  AND U10623 ( .A(n10683), .B(n10686), .Z(n10733) );
  XOR U10624 ( .A(n10779), .B(n10760), .Z(n10686) );
  XNOR U10625 ( .A(p_input[1024]), .B(p_input[240]), .Z(n10760) );
  XOR U10626 ( .A(n10748), .B(n10747), .Z(n10779) );
  XNOR U10627 ( .A(n10780), .B(n10754), .Z(n10747) );
  XNOR U10628 ( .A(n10743), .B(n10742), .Z(n10754) );
  XOR U10629 ( .A(n10781), .B(n10739), .Z(n10742) );
  XOR U10630 ( .A(p_input[1034]), .B(p_input[250]), .Z(n10739) );
  XNOR U10631 ( .A(p_input[1035]), .B(p_input[251]), .Z(n10781) );
  XOR U10632 ( .A(p_input[1036]), .B(p_input[252]), .Z(n10743) );
  XNOR U10633 ( .A(n10753), .B(n10744), .Z(n10780) );
  XOR U10634 ( .A(p_input[1025]), .B(p_input[241]), .Z(n10744) );
  XOR U10635 ( .A(n10782), .B(n10759), .Z(n10753) );
  XNOR U10636 ( .A(p_input[1039]), .B(p_input[255]), .Z(n10759) );
  XOR U10637 ( .A(n10750), .B(n10758), .Z(n10782) );
  XOR U10638 ( .A(n10783), .B(n10755), .Z(n10758) );
  XOR U10639 ( .A(p_input[1037]), .B(p_input[253]), .Z(n10755) );
  XNOR U10640 ( .A(p_input[1038]), .B(p_input[254]), .Z(n10783) );
  XOR U10641 ( .A(p_input[1033]), .B(p_input[249]), .Z(n10750) );
  XNOR U10642 ( .A(n10766), .B(n10765), .Z(n10748) );
  XNOR U10643 ( .A(n10784), .B(n10771), .Z(n10765) );
  XOR U10644 ( .A(p_input[1032]), .B(p_input[248]), .Z(n10771) );
  XOR U10645 ( .A(n10762), .B(n10770), .Z(n10784) );
  XOR U10646 ( .A(n10785), .B(n10767), .Z(n10770) );
  XOR U10647 ( .A(p_input[1030]), .B(p_input[246]), .Z(n10767) );
  XNOR U10648 ( .A(p_input[1031]), .B(p_input[247]), .Z(n10785) );
  XOR U10649 ( .A(p_input[1026]), .B(p_input[242]), .Z(n10762) );
  XNOR U10650 ( .A(n10776), .B(n10775), .Z(n10766) );
  XOR U10651 ( .A(n10786), .B(n10772), .Z(n10775) );
  XOR U10652 ( .A(p_input[1027]), .B(p_input[243]), .Z(n10772) );
  XNOR U10653 ( .A(p_input[1028]), .B(p_input[244]), .Z(n10786) );
  XOR U10654 ( .A(p_input[1029]), .B(p_input[245]), .Z(n10776) );
  XNOR U10655 ( .A(n10787), .B(n10788), .Z(n10683) );
  AND U10656 ( .A(n204), .B(n10789), .Z(n10788) );
  XNOR U10657 ( .A(n10790), .B(n10791), .Z(n204) );
  AND U10658 ( .A(n10792), .B(n10793), .Z(n10791) );
  XOR U10659 ( .A(n10790), .B(n10693), .Z(n10793) );
  XNOR U10660 ( .A(n10790), .B(n10647), .Z(n10792) );
  XOR U10661 ( .A(n10794), .B(n10795), .Z(n10790) );
  AND U10662 ( .A(n10796), .B(n10797), .Z(n10795) );
  XOR U10663 ( .A(n10794), .B(n10657), .Z(n10796) );
  XOR U10664 ( .A(n10798), .B(n10799), .Z(n10636) );
  AND U10665 ( .A(n208), .B(n10789), .Z(n10799) );
  XNOR U10666 ( .A(n10787), .B(n10798), .Z(n10789) );
  XNOR U10667 ( .A(n10800), .B(n10801), .Z(n208) );
  AND U10668 ( .A(n10802), .B(n10803), .Z(n10801) );
  XNOR U10669 ( .A(n10804), .B(n10800), .Z(n10803) );
  IV U10670 ( .A(n10693), .Z(n10804) );
  XNOR U10671 ( .A(n10805), .B(n10806), .Z(n10693) );
  AND U10672 ( .A(n211), .B(n10807), .Z(n10806) );
  XNOR U10673 ( .A(n10805), .B(n10808), .Z(n10807) );
  XNOR U10674 ( .A(n10647), .B(n10800), .Z(n10802) );
  XOR U10675 ( .A(n10809), .B(n10810), .Z(n10647) );
  AND U10676 ( .A(n219), .B(n10811), .Z(n10810) );
  XOR U10677 ( .A(n10794), .B(n10812), .Z(n10800) );
  AND U10678 ( .A(n10813), .B(n10797), .Z(n10812) );
  XNOR U10679 ( .A(n10706), .B(n10794), .Z(n10797) );
  XNOR U10680 ( .A(n10814), .B(n10815), .Z(n10706) );
  AND U10681 ( .A(n211), .B(n10816), .Z(n10815) );
  XOR U10682 ( .A(n10817), .B(n10814), .Z(n10816) );
  XNOR U10683 ( .A(n10818), .B(n10794), .Z(n10813) );
  IV U10684 ( .A(n10657), .Z(n10818) );
  XOR U10685 ( .A(n10819), .B(n10820), .Z(n10657) );
  AND U10686 ( .A(n219), .B(n10821), .Z(n10820) );
  XOR U10687 ( .A(n10822), .B(n10823), .Z(n10794) );
  AND U10688 ( .A(n10824), .B(n10825), .Z(n10823) );
  XNOR U10689 ( .A(n10731), .B(n10822), .Z(n10825) );
  XNOR U10690 ( .A(n10826), .B(n10827), .Z(n10731) );
  AND U10691 ( .A(n211), .B(n10828), .Z(n10827) );
  XNOR U10692 ( .A(n10829), .B(n10826), .Z(n10828) );
  XOR U10693 ( .A(n10822), .B(n10668), .Z(n10824) );
  XOR U10694 ( .A(n10830), .B(n10831), .Z(n10668) );
  AND U10695 ( .A(n219), .B(n10832), .Z(n10831) );
  XOR U10696 ( .A(n10833), .B(n10834), .Z(n10822) );
  AND U10697 ( .A(n10835), .B(n10836), .Z(n10834) );
  XNOR U10698 ( .A(n10833), .B(n10777), .Z(n10836) );
  XNOR U10699 ( .A(n10837), .B(n10838), .Z(n10777) );
  AND U10700 ( .A(n211), .B(n10839), .Z(n10838) );
  XOR U10701 ( .A(n10840), .B(n10837), .Z(n10839) );
  XNOR U10702 ( .A(n10841), .B(n10833), .Z(n10835) );
  IV U10703 ( .A(n10680), .Z(n10841) );
  XOR U10704 ( .A(n10842), .B(n10843), .Z(n10680) );
  AND U10705 ( .A(n219), .B(n10844), .Z(n10843) );
  AND U10706 ( .A(n10798), .B(n10787), .Z(n10833) );
  XNOR U10707 ( .A(n10845), .B(n10846), .Z(n10787) );
  AND U10708 ( .A(n211), .B(n10847), .Z(n10846) );
  XNOR U10709 ( .A(n10848), .B(n10845), .Z(n10847) );
  XNOR U10710 ( .A(n10849), .B(n10850), .Z(n211) );
  AND U10711 ( .A(n10851), .B(n10852), .Z(n10850) );
  XOR U10712 ( .A(n10808), .B(n10849), .Z(n10852) );
  AND U10713 ( .A(n10853), .B(n10854), .Z(n10808) );
  XOR U10714 ( .A(n10849), .B(n10805), .Z(n10851) );
  XNOR U10715 ( .A(n10855), .B(n10856), .Z(n10805) );
  AND U10716 ( .A(n215), .B(n10811), .Z(n10856) );
  XOR U10717 ( .A(n10809), .B(n10855), .Z(n10811) );
  XOR U10718 ( .A(n10857), .B(n10858), .Z(n10849) );
  AND U10719 ( .A(n10859), .B(n10860), .Z(n10858) );
  XNOR U10720 ( .A(n10857), .B(n10853), .Z(n10860) );
  IV U10721 ( .A(n10817), .Z(n10853) );
  XOR U10722 ( .A(n10861), .B(n10862), .Z(n10817) );
  XOR U10723 ( .A(n10863), .B(n10854), .Z(n10862) );
  AND U10724 ( .A(n10829), .B(n10864), .Z(n10854) );
  AND U10725 ( .A(n10865), .B(n10866), .Z(n10863) );
  XOR U10726 ( .A(n10867), .B(n10861), .Z(n10865) );
  XNOR U10727 ( .A(n10814), .B(n10857), .Z(n10859) );
  XNOR U10728 ( .A(n10868), .B(n10869), .Z(n10814) );
  AND U10729 ( .A(n215), .B(n10821), .Z(n10869) );
  XOR U10730 ( .A(n10868), .B(n10819), .Z(n10821) );
  XOR U10731 ( .A(n10870), .B(n10871), .Z(n10857) );
  AND U10732 ( .A(n10872), .B(n10873), .Z(n10871) );
  XNOR U10733 ( .A(n10870), .B(n10829), .Z(n10873) );
  XOR U10734 ( .A(n10874), .B(n10866), .Z(n10829) );
  XNOR U10735 ( .A(n10875), .B(n10861), .Z(n10866) );
  XOR U10736 ( .A(n10876), .B(n10877), .Z(n10861) );
  AND U10737 ( .A(n10878), .B(n10879), .Z(n10877) );
  XOR U10738 ( .A(n10880), .B(n10876), .Z(n10878) );
  XNOR U10739 ( .A(n10881), .B(n10882), .Z(n10875) );
  AND U10740 ( .A(n10883), .B(n10884), .Z(n10882) );
  XOR U10741 ( .A(n10881), .B(n10885), .Z(n10883) );
  XNOR U10742 ( .A(n10867), .B(n10864), .Z(n10874) );
  AND U10743 ( .A(n10886), .B(n10887), .Z(n10864) );
  XOR U10744 ( .A(n10888), .B(n10889), .Z(n10867) );
  AND U10745 ( .A(n10890), .B(n10891), .Z(n10889) );
  XOR U10746 ( .A(n10888), .B(n10892), .Z(n10890) );
  XNOR U10747 ( .A(n10826), .B(n10870), .Z(n10872) );
  XNOR U10748 ( .A(n10893), .B(n10894), .Z(n10826) );
  AND U10749 ( .A(n215), .B(n10832), .Z(n10894) );
  XOR U10750 ( .A(n10893), .B(n10830), .Z(n10832) );
  XOR U10751 ( .A(n10895), .B(n10896), .Z(n10870) );
  AND U10752 ( .A(n10897), .B(n10898), .Z(n10896) );
  XNOR U10753 ( .A(n10895), .B(n10886), .Z(n10898) );
  IV U10754 ( .A(n10840), .Z(n10886) );
  XNOR U10755 ( .A(n10899), .B(n10879), .Z(n10840) );
  XNOR U10756 ( .A(n10900), .B(n10885), .Z(n10879) );
  XOR U10757 ( .A(n10901), .B(n10902), .Z(n10885) );
  NOR U10758 ( .A(n10903), .B(n10904), .Z(n10902) );
  XNOR U10759 ( .A(n10901), .B(n10905), .Z(n10903) );
  XNOR U10760 ( .A(n10884), .B(n10876), .Z(n10900) );
  XOR U10761 ( .A(n10906), .B(n10907), .Z(n10876) );
  AND U10762 ( .A(n10908), .B(n10909), .Z(n10907) );
  XNOR U10763 ( .A(n10906), .B(n10910), .Z(n10908) );
  XNOR U10764 ( .A(n10911), .B(n10881), .Z(n10884) );
  XOR U10765 ( .A(n10912), .B(n10913), .Z(n10881) );
  AND U10766 ( .A(n10914), .B(n10915), .Z(n10913) );
  XOR U10767 ( .A(n10912), .B(n10916), .Z(n10914) );
  XNOR U10768 ( .A(n10917), .B(n10918), .Z(n10911) );
  NOR U10769 ( .A(n10919), .B(n10920), .Z(n10918) );
  XOR U10770 ( .A(n10917), .B(n10921), .Z(n10919) );
  XNOR U10771 ( .A(n10880), .B(n10887), .Z(n10899) );
  NOR U10772 ( .A(n10848), .B(n10922), .Z(n10887) );
  XOR U10773 ( .A(n10892), .B(n10891), .Z(n10880) );
  XNOR U10774 ( .A(n10923), .B(n10888), .Z(n10891) );
  XOR U10775 ( .A(n10924), .B(n10925), .Z(n10888) );
  AND U10776 ( .A(n10926), .B(n10927), .Z(n10925) );
  XOR U10777 ( .A(n10924), .B(n10928), .Z(n10926) );
  XNOR U10778 ( .A(n10929), .B(n10930), .Z(n10923) );
  NOR U10779 ( .A(n10931), .B(n10932), .Z(n10930) );
  XNOR U10780 ( .A(n10929), .B(n10933), .Z(n10931) );
  XOR U10781 ( .A(n10934), .B(n10935), .Z(n10892) );
  NOR U10782 ( .A(n10936), .B(n10937), .Z(n10935) );
  XNOR U10783 ( .A(n10934), .B(n10938), .Z(n10936) );
  XNOR U10784 ( .A(n10837), .B(n10895), .Z(n10897) );
  XNOR U10785 ( .A(n10939), .B(n10940), .Z(n10837) );
  AND U10786 ( .A(n215), .B(n10844), .Z(n10940) );
  XOR U10787 ( .A(n10939), .B(n10842), .Z(n10844) );
  AND U10788 ( .A(n10845), .B(n10848), .Z(n10895) );
  XOR U10789 ( .A(n10941), .B(n10922), .Z(n10848) );
  XNOR U10790 ( .A(p_input[1024]), .B(p_input[256]), .Z(n10922) );
  XOR U10791 ( .A(n10910), .B(n10909), .Z(n10941) );
  XNOR U10792 ( .A(n10942), .B(n10916), .Z(n10909) );
  XNOR U10793 ( .A(n10905), .B(n10904), .Z(n10916) );
  XOR U10794 ( .A(n10943), .B(n10901), .Z(n10904) );
  XOR U10795 ( .A(p_input[1034]), .B(p_input[266]), .Z(n10901) );
  XNOR U10796 ( .A(p_input[1035]), .B(p_input[267]), .Z(n10943) );
  XOR U10797 ( .A(p_input[1036]), .B(p_input[268]), .Z(n10905) );
  XNOR U10798 ( .A(n10915), .B(n10906), .Z(n10942) );
  XOR U10799 ( .A(p_input[1025]), .B(p_input[257]), .Z(n10906) );
  XOR U10800 ( .A(n10944), .B(n10921), .Z(n10915) );
  XNOR U10801 ( .A(p_input[1039]), .B(p_input[271]), .Z(n10921) );
  XOR U10802 ( .A(n10912), .B(n10920), .Z(n10944) );
  XOR U10803 ( .A(n10945), .B(n10917), .Z(n10920) );
  XOR U10804 ( .A(p_input[1037]), .B(p_input[269]), .Z(n10917) );
  XNOR U10805 ( .A(p_input[1038]), .B(p_input[270]), .Z(n10945) );
  XOR U10806 ( .A(p_input[1033]), .B(p_input[265]), .Z(n10912) );
  XNOR U10807 ( .A(n10928), .B(n10927), .Z(n10910) );
  XNOR U10808 ( .A(n10946), .B(n10933), .Z(n10927) );
  XOR U10809 ( .A(p_input[1032]), .B(p_input[264]), .Z(n10933) );
  XOR U10810 ( .A(n10924), .B(n10932), .Z(n10946) );
  XOR U10811 ( .A(n10947), .B(n10929), .Z(n10932) );
  XOR U10812 ( .A(p_input[1030]), .B(p_input[262]), .Z(n10929) );
  XNOR U10813 ( .A(p_input[1031]), .B(p_input[263]), .Z(n10947) );
  XOR U10814 ( .A(p_input[1026]), .B(p_input[258]), .Z(n10924) );
  XNOR U10815 ( .A(n10938), .B(n10937), .Z(n10928) );
  XOR U10816 ( .A(n10948), .B(n10934), .Z(n10937) );
  XOR U10817 ( .A(p_input[1027]), .B(p_input[259]), .Z(n10934) );
  XNOR U10818 ( .A(p_input[1028]), .B(p_input[260]), .Z(n10948) );
  XOR U10819 ( .A(p_input[1029]), .B(p_input[261]), .Z(n10938) );
  XNOR U10820 ( .A(n10949), .B(n10950), .Z(n10845) );
  AND U10821 ( .A(n215), .B(n10951), .Z(n10950) );
  XNOR U10822 ( .A(n10952), .B(n10953), .Z(n215) );
  AND U10823 ( .A(n10954), .B(n10955), .Z(n10953) );
  XOR U10824 ( .A(n10952), .B(n10855), .Z(n10955) );
  XNOR U10825 ( .A(n10952), .B(n10809), .Z(n10954) );
  XOR U10826 ( .A(n10956), .B(n10957), .Z(n10952) );
  AND U10827 ( .A(n10958), .B(n10959), .Z(n10957) );
  XOR U10828 ( .A(n10956), .B(n10819), .Z(n10958) );
  XOR U10829 ( .A(n10960), .B(n10961), .Z(n10798) );
  AND U10830 ( .A(n219), .B(n10951), .Z(n10961) );
  XNOR U10831 ( .A(n10949), .B(n10960), .Z(n10951) );
  XNOR U10832 ( .A(n10962), .B(n10963), .Z(n219) );
  AND U10833 ( .A(n10964), .B(n10965), .Z(n10963) );
  XNOR U10834 ( .A(n10966), .B(n10962), .Z(n10965) );
  IV U10835 ( .A(n10855), .Z(n10966) );
  XNOR U10836 ( .A(n10967), .B(n10968), .Z(n10855) );
  AND U10837 ( .A(n222), .B(n10969), .Z(n10968) );
  XNOR U10838 ( .A(n10967), .B(n10970), .Z(n10969) );
  XNOR U10839 ( .A(n10809), .B(n10962), .Z(n10964) );
  XOR U10840 ( .A(n10971), .B(n10972), .Z(n10809) );
  AND U10841 ( .A(n230), .B(n10973), .Z(n10972) );
  XOR U10842 ( .A(n10956), .B(n10974), .Z(n10962) );
  AND U10843 ( .A(n10975), .B(n10959), .Z(n10974) );
  XNOR U10844 ( .A(n10868), .B(n10956), .Z(n10959) );
  XNOR U10845 ( .A(n10976), .B(n10977), .Z(n10868) );
  AND U10846 ( .A(n222), .B(n10978), .Z(n10977) );
  XOR U10847 ( .A(n10979), .B(n10976), .Z(n10978) );
  XNOR U10848 ( .A(n10980), .B(n10956), .Z(n10975) );
  IV U10849 ( .A(n10819), .Z(n10980) );
  XOR U10850 ( .A(n10981), .B(n10982), .Z(n10819) );
  AND U10851 ( .A(n230), .B(n10983), .Z(n10982) );
  XOR U10852 ( .A(n10984), .B(n10985), .Z(n10956) );
  AND U10853 ( .A(n10986), .B(n10987), .Z(n10985) );
  XNOR U10854 ( .A(n10893), .B(n10984), .Z(n10987) );
  XNOR U10855 ( .A(n10988), .B(n10989), .Z(n10893) );
  AND U10856 ( .A(n222), .B(n10990), .Z(n10989) );
  XNOR U10857 ( .A(n10991), .B(n10988), .Z(n10990) );
  XOR U10858 ( .A(n10984), .B(n10830), .Z(n10986) );
  XOR U10859 ( .A(n10992), .B(n10993), .Z(n10830) );
  AND U10860 ( .A(n230), .B(n10994), .Z(n10993) );
  XOR U10861 ( .A(n10995), .B(n10996), .Z(n10984) );
  AND U10862 ( .A(n10997), .B(n10998), .Z(n10996) );
  XNOR U10863 ( .A(n10995), .B(n10939), .Z(n10998) );
  XNOR U10864 ( .A(n10999), .B(n11000), .Z(n10939) );
  AND U10865 ( .A(n222), .B(n11001), .Z(n11000) );
  XOR U10866 ( .A(n11002), .B(n10999), .Z(n11001) );
  XNOR U10867 ( .A(n11003), .B(n10995), .Z(n10997) );
  IV U10868 ( .A(n10842), .Z(n11003) );
  XOR U10869 ( .A(n11004), .B(n11005), .Z(n10842) );
  AND U10870 ( .A(n230), .B(n11006), .Z(n11005) );
  AND U10871 ( .A(n10960), .B(n10949), .Z(n10995) );
  XNOR U10872 ( .A(n11007), .B(n11008), .Z(n10949) );
  AND U10873 ( .A(n222), .B(n11009), .Z(n11008) );
  XNOR U10874 ( .A(n11010), .B(n11007), .Z(n11009) );
  XNOR U10875 ( .A(n11011), .B(n11012), .Z(n222) );
  AND U10876 ( .A(n11013), .B(n11014), .Z(n11012) );
  XOR U10877 ( .A(n10970), .B(n11011), .Z(n11014) );
  AND U10878 ( .A(n11015), .B(n11016), .Z(n10970) );
  XOR U10879 ( .A(n11011), .B(n10967), .Z(n11013) );
  XNOR U10880 ( .A(n11017), .B(n11018), .Z(n10967) );
  AND U10881 ( .A(n226), .B(n10973), .Z(n11018) );
  XOR U10882 ( .A(n10971), .B(n11017), .Z(n10973) );
  XOR U10883 ( .A(n11019), .B(n11020), .Z(n11011) );
  AND U10884 ( .A(n11021), .B(n11022), .Z(n11020) );
  XNOR U10885 ( .A(n11019), .B(n11015), .Z(n11022) );
  IV U10886 ( .A(n10979), .Z(n11015) );
  XOR U10887 ( .A(n11023), .B(n11024), .Z(n10979) );
  XOR U10888 ( .A(n11025), .B(n11016), .Z(n11024) );
  AND U10889 ( .A(n10991), .B(n11026), .Z(n11016) );
  AND U10890 ( .A(n11027), .B(n11028), .Z(n11025) );
  XOR U10891 ( .A(n11029), .B(n11023), .Z(n11027) );
  XNOR U10892 ( .A(n10976), .B(n11019), .Z(n11021) );
  XNOR U10893 ( .A(n11030), .B(n11031), .Z(n10976) );
  AND U10894 ( .A(n226), .B(n10983), .Z(n11031) );
  XOR U10895 ( .A(n11030), .B(n10981), .Z(n10983) );
  XOR U10896 ( .A(n11032), .B(n11033), .Z(n11019) );
  AND U10897 ( .A(n11034), .B(n11035), .Z(n11033) );
  XNOR U10898 ( .A(n11032), .B(n10991), .Z(n11035) );
  XOR U10899 ( .A(n11036), .B(n11028), .Z(n10991) );
  XNOR U10900 ( .A(n11037), .B(n11023), .Z(n11028) );
  XOR U10901 ( .A(n11038), .B(n11039), .Z(n11023) );
  AND U10902 ( .A(n11040), .B(n11041), .Z(n11039) );
  XOR U10903 ( .A(n11042), .B(n11038), .Z(n11040) );
  XNOR U10904 ( .A(n11043), .B(n11044), .Z(n11037) );
  AND U10905 ( .A(n11045), .B(n11046), .Z(n11044) );
  XOR U10906 ( .A(n11043), .B(n11047), .Z(n11045) );
  XNOR U10907 ( .A(n11029), .B(n11026), .Z(n11036) );
  AND U10908 ( .A(n11048), .B(n11049), .Z(n11026) );
  XOR U10909 ( .A(n11050), .B(n11051), .Z(n11029) );
  AND U10910 ( .A(n11052), .B(n11053), .Z(n11051) );
  XOR U10911 ( .A(n11050), .B(n11054), .Z(n11052) );
  XNOR U10912 ( .A(n10988), .B(n11032), .Z(n11034) );
  XNOR U10913 ( .A(n11055), .B(n11056), .Z(n10988) );
  AND U10914 ( .A(n226), .B(n10994), .Z(n11056) );
  XOR U10915 ( .A(n11055), .B(n10992), .Z(n10994) );
  XOR U10916 ( .A(n11057), .B(n11058), .Z(n11032) );
  AND U10917 ( .A(n11059), .B(n11060), .Z(n11058) );
  XNOR U10918 ( .A(n11057), .B(n11048), .Z(n11060) );
  IV U10919 ( .A(n11002), .Z(n11048) );
  XNOR U10920 ( .A(n11061), .B(n11041), .Z(n11002) );
  XNOR U10921 ( .A(n11062), .B(n11047), .Z(n11041) );
  XOR U10922 ( .A(n11063), .B(n11064), .Z(n11047) );
  NOR U10923 ( .A(n11065), .B(n11066), .Z(n11064) );
  XNOR U10924 ( .A(n11063), .B(n11067), .Z(n11065) );
  XNOR U10925 ( .A(n11046), .B(n11038), .Z(n11062) );
  XOR U10926 ( .A(n11068), .B(n11069), .Z(n11038) );
  AND U10927 ( .A(n11070), .B(n11071), .Z(n11069) );
  XNOR U10928 ( .A(n11068), .B(n11072), .Z(n11070) );
  XNOR U10929 ( .A(n11073), .B(n11043), .Z(n11046) );
  XOR U10930 ( .A(n11074), .B(n11075), .Z(n11043) );
  AND U10931 ( .A(n11076), .B(n11077), .Z(n11075) );
  XOR U10932 ( .A(n11074), .B(n11078), .Z(n11076) );
  XNOR U10933 ( .A(n11079), .B(n11080), .Z(n11073) );
  NOR U10934 ( .A(n11081), .B(n11082), .Z(n11080) );
  XOR U10935 ( .A(n11079), .B(n11083), .Z(n11081) );
  XNOR U10936 ( .A(n11042), .B(n11049), .Z(n11061) );
  NOR U10937 ( .A(n11010), .B(n11084), .Z(n11049) );
  XOR U10938 ( .A(n11054), .B(n11053), .Z(n11042) );
  XNOR U10939 ( .A(n11085), .B(n11050), .Z(n11053) );
  XOR U10940 ( .A(n11086), .B(n11087), .Z(n11050) );
  AND U10941 ( .A(n11088), .B(n11089), .Z(n11087) );
  XOR U10942 ( .A(n11086), .B(n11090), .Z(n11088) );
  XNOR U10943 ( .A(n11091), .B(n11092), .Z(n11085) );
  NOR U10944 ( .A(n11093), .B(n11094), .Z(n11092) );
  XNOR U10945 ( .A(n11091), .B(n11095), .Z(n11093) );
  XOR U10946 ( .A(n11096), .B(n11097), .Z(n11054) );
  NOR U10947 ( .A(n11098), .B(n11099), .Z(n11097) );
  XNOR U10948 ( .A(n11096), .B(n11100), .Z(n11098) );
  XNOR U10949 ( .A(n10999), .B(n11057), .Z(n11059) );
  XNOR U10950 ( .A(n11101), .B(n11102), .Z(n10999) );
  AND U10951 ( .A(n226), .B(n11006), .Z(n11102) );
  XOR U10952 ( .A(n11101), .B(n11004), .Z(n11006) );
  AND U10953 ( .A(n11007), .B(n11010), .Z(n11057) );
  XOR U10954 ( .A(n11103), .B(n11084), .Z(n11010) );
  XNOR U10955 ( .A(p_input[1024]), .B(p_input[272]), .Z(n11084) );
  XOR U10956 ( .A(n11072), .B(n11071), .Z(n11103) );
  XNOR U10957 ( .A(n11104), .B(n11078), .Z(n11071) );
  XNOR U10958 ( .A(n11067), .B(n11066), .Z(n11078) );
  XOR U10959 ( .A(n11105), .B(n11063), .Z(n11066) );
  XOR U10960 ( .A(p_input[1034]), .B(p_input[282]), .Z(n11063) );
  XNOR U10961 ( .A(p_input[1035]), .B(p_input[283]), .Z(n11105) );
  XOR U10962 ( .A(p_input[1036]), .B(p_input[284]), .Z(n11067) );
  XNOR U10963 ( .A(n11077), .B(n11068), .Z(n11104) );
  XOR U10964 ( .A(p_input[1025]), .B(p_input[273]), .Z(n11068) );
  XOR U10965 ( .A(n11106), .B(n11083), .Z(n11077) );
  XNOR U10966 ( .A(p_input[1039]), .B(p_input[287]), .Z(n11083) );
  XOR U10967 ( .A(n11074), .B(n11082), .Z(n11106) );
  XOR U10968 ( .A(n11107), .B(n11079), .Z(n11082) );
  XOR U10969 ( .A(p_input[1037]), .B(p_input[285]), .Z(n11079) );
  XNOR U10970 ( .A(p_input[1038]), .B(p_input[286]), .Z(n11107) );
  XOR U10971 ( .A(p_input[1033]), .B(p_input[281]), .Z(n11074) );
  XNOR U10972 ( .A(n11090), .B(n11089), .Z(n11072) );
  XNOR U10973 ( .A(n11108), .B(n11095), .Z(n11089) );
  XOR U10974 ( .A(p_input[1032]), .B(p_input[280]), .Z(n11095) );
  XOR U10975 ( .A(n11086), .B(n11094), .Z(n11108) );
  XOR U10976 ( .A(n11109), .B(n11091), .Z(n11094) );
  XOR U10977 ( .A(p_input[1030]), .B(p_input[278]), .Z(n11091) );
  XNOR U10978 ( .A(p_input[1031]), .B(p_input[279]), .Z(n11109) );
  XOR U10979 ( .A(p_input[1026]), .B(p_input[274]), .Z(n11086) );
  XNOR U10980 ( .A(n11100), .B(n11099), .Z(n11090) );
  XOR U10981 ( .A(n11110), .B(n11096), .Z(n11099) );
  XOR U10982 ( .A(p_input[1027]), .B(p_input[275]), .Z(n11096) );
  XNOR U10983 ( .A(p_input[1028]), .B(p_input[276]), .Z(n11110) );
  XOR U10984 ( .A(p_input[1029]), .B(p_input[277]), .Z(n11100) );
  XNOR U10985 ( .A(n11111), .B(n11112), .Z(n11007) );
  AND U10986 ( .A(n226), .B(n11113), .Z(n11112) );
  XNOR U10987 ( .A(n11114), .B(n11115), .Z(n226) );
  AND U10988 ( .A(n11116), .B(n11117), .Z(n11115) );
  XOR U10989 ( .A(n11114), .B(n11017), .Z(n11117) );
  XNOR U10990 ( .A(n11114), .B(n10971), .Z(n11116) );
  XOR U10991 ( .A(n11118), .B(n11119), .Z(n11114) );
  AND U10992 ( .A(n11120), .B(n11121), .Z(n11119) );
  XOR U10993 ( .A(n11118), .B(n10981), .Z(n11120) );
  XOR U10994 ( .A(n11122), .B(n11123), .Z(n10960) );
  AND U10995 ( .A(n230), .B(n11113), .Z(n11123) );
  XNOR U10996 ( .A(n11111), .B(n11122), .Z(n11113) );
  XNOR U10997 ( .A(n11124), .B(n11125), .Z(n230) );
  AND U10998 ( .A(n11126), .B(n11127), .Z(n11125) );
  XNOR U10999 ( .A(n11128), .B(n11124), .Z(n11127) );
  IV U11000 ( .A(n11017), .Z(n11128) );
  XNOR U11001 ( .A(n11129), .B(n11130), .Z(n11017) );
  AND U11002 ( .A(n233), .B(n11131), .Z(n11130) );
  XNOR U11003 ( .A(n11129), .B(n11132), .Z(n11131) );
  XNOR U11004 ( .A(n10971), .B(n11124), .Z(n11126) );
  XOR U11005 ( .A(n11133), .B(n11134), .Z(n10971) );
  AND U11006 ( .A(n241), .B(n11135), .Z(n11134) );
  XOR U11007 ( .A(n11118), .B(n11136), .Z(n11124) );
  AND U11008 ( .A(n11137), .B(n11121), .Z(n11136) );
  XNOR U11009 ( .A(n11030), .B(n11118), .Z(n11121) );
  XNOR U11010 ( .A(n11138), .B(n11139), .Z(n11030) );
  AND U11011 ( .A(n233), .B(n11140), .Z(n11139) );
  XOR U11012 ( .A(n11141), .B(n11138), .Z(n11140) );
  XNOR U11013 ( .A(n11142), .B(n11118), .Z(n11137) );
  IV U11014 ( .A(n10981), .Z(n11142) );
  XOR U11015 ( .A(n11143), .B(n11144), .Z(n10981) );
  AND U11016 ( .A(n241), .B(n11145), .Z(n11144) );
  XOR U11017 ( .A(n11146), .B(n11147), .Z(n11118) );
  AND U11018 ( .A(n11148), .B(n11149), .Z(n11147) );
  XNOR U11019 ( .A(n11055), .B(n11146), .Z(n11149) );
  XNOR U11020 ( .A(n11150), .B(n11151), .Z(n11055) );
  AND U11021 ( .A(n233), .B(n11152), .Z(n11151) );
  XNOR U11022 ( .A(n11153), .B(n11150), .Z(n11152) );
  XOR U11023 ( .A(n11146), .B(n10992), .Z(n11148) );
  XOR U11024 ( .A(n11154), .B(n11155), .Z(n10992) );
  AND U11025 ( .A(n241), .B(n11156), .Z(n11155) );
  XOR U11026 ( .A(n11157), .B(n11158), .Z(n11146) );
  AND U11027 ( .A(n11159), .B(n11160), .Z(n11158) );
  XNOR U11028 ( .A(n11157), .B(n11101), .Z(n11160) );
  XNOR U11029 ( .A(n11161), .B(n11162), .Z(n11101) );
  AND U11030 ( .A(n233), .B(n11163), .Z(n11162) );
  XOR U11031 ( .A(n11164), .B(n11161), .Z(n11163) );
  XNOR U11032 ( .A(n11165), .B(n11157), .Z(n11159) );
  IV U11033 ( .A(n11004), .Z(n11165) );
  XOR U11034 ( .A(n11166), .B(n11167), .Z(n11004) );
  AND U11035 ( .A(n241), .B(n11168), .Z(n11167) );
  AND U11036 ( .A(n11122), .B(n11111), .Z(n11157) );
  XNOR U11037 ( .A(n11169), .B(n11170), .Z(n11111) );
  AND U11038 ( .A(n233), .B(n11171), .Z(n11170) );
  XNOR U11039 ( .A(n11172), .B(n11169), .Z(n11171) );
  XNOR U11040 ( .A(n11173), .B(n11174), .Z(n233) );
  AND U11041 ( .A(n11175), .B(n11176), .Z(n11174) );
  XOR U11042 ( .A(n11132), .B(n11173), .Z(n11176) );
  AND U11043 ( .A(n11177), .B(n11178), .Z(n11132) );
  XOR U11044 ( .A(n11173), .B(n11129), .Z(n11175) );
  XNOR U11045 ( .A(n11179), .B(n11180), .Z(n11129) );
  AND U11046 ( .A(n237), .B(n11135), .Z(n11180) );
  XOR U11047 ( .A(n11133), .B(n11179), .Z(n11135) );
  XOR U11048 ( .A(n11181), .B(n11182), .Z(n11173) );
  AND U11049 ( .A(n11183), .B(n11184), .Z(n11182) );
  XNOR U11050 ( .A(n11181), .B(n11177), .Z(n11184) );
  IV U11051 ( .A(n11141), .Z(n11177) );
  XOR U11052 ( .A(n11185), .B(n11186), .Z(n11141) );
  XOR U11053 ( .A(n11187), .B(n11178), .Z(n11186) );
  AND U11054 ( .A(n11153), .B(n11188), .Z(n11178) );
  AND U11055 ( .A(n11189), .B(n11190), .Z(n11187) );
  XOR U11056 ( .A(n11191), .B(n11185), .Z(n11189) );
  XNOR U11057 ( .A(n11138), .B(n11181), .Z(n11183) );
  XNOR U11058 ( .A(n11192), .B(n11193), .Z(n11138) );
  AND U11059 ( .A(n237), .B(n11145), .Z(n11193) );
  XOR U11060 ( .A(n11192), .B(n11143), .Z(n11145) );
  XOR U11061 ( .A(n11194), .B(n11195), .Z(n11181) );
  AND U11062 ( .A(n11196), .B(n11197), .Z(n11195) );
  XNOR U11063 ( .A(n11194), .B(n11153), .Z(n11197) );
  XOR U11064 ( .A(n11198), .B(n11190), .Z(n11153) );
  XNOR U11065 ( .A(n11199), .B(n11185), .Z(n11190) );
  XOR U11066 ( .A(n11200), .B(n11201), .Z(n11185) );
  AND U11067 ( .A(n11202), .B(n11203), .Z(n11201) );
  XOR U11068 ( .A(n11204), .B(n11200), .Z(n11202) );
  XNOR U11069 ( .A(n11205), .B(n11206), .Z(n11199) );
  AND U11070 ( .A(n11207), .B(n11208), .Z(n11206) );
  XOR U11071 ( .A(n11205), .B(n11209), .Z(n11207) );
  XNOR U11072 ( .A(n11191), .B(n11188), .Z(n11198) );
  AND U11073 ( .A(n11210), .B(n11211), .Z(n11188) );
  XOR U11074 ( .A(n11212), .B(n11213), .Z(n11191) );
  AND U11075 ( .A(n11214), .B(n11215), .Z(n11213) );
  XOR U11076 ( .A(n11212), .B(n11216), .Z(n11214) );
  XNOR U11077 ( .A(n11150), .B(n11194), .Z(n11196) );
  XNOR U11078 ( .A(n11217), .B(n11218), .Z(n11150) );
  AND U11079 ( .A(n237), .B(n11156), .Z(n11218) );
  XOR U11080 ( .A(n11217), .B(n11154), .Z(n11156) );
  XOR U11081 ( .A(n11219), .B(n11220), .Z(n11194) );
  AND U11082 ( .A(n11221), .B(n11222), .Z(n11220) );
  XNOR U11083 ( .A(n11219), .B(n11210), .Z(n11222) );
  IV U11084 ( .A(n11164), .Z(n11210) );
  XNOR U11085 ( .A(n11223), .B(n11203), .Z(n11164) );
  XNOR U11086 ( .A(n11224), .B(n11209), .Z(n11203) );
  XOR U11087 ( .A(n11225), .B(n11226), .Z(n11209) );
  NOR U11088 ( .A(n11227), .B(n11228), .Z(n11226) );
  XNOR U11089 ( .A(n11225), .B(n11229), .Z(n11227) );
  XNOR U11090 ( .A(n11208), .B(n11200), .Z(n11224) );
  XOR U11091 ( .A(n11230), .B(n11231), .Z(n11200) );
  AND U11092 ( .A(n11232), .B(n11233), .Z(n11231) );
  XNOR U11093 ( .A(n11230), .B(n11234), .Z(n11232) );
  XNOR U11094 ( .A(n11235), .B(n11205), .Z(n11208) );
  XOR U11095 ( .A(n11236), .B(n11237), .Z(n11205) );
  AND U11096 ( .A(n11238), .B(n11239), .Z(n11237) );
  XOR U11097 ( .A(n11236), .B(n11240), .Z(n11238) );
  XNOR U11098 ( .A(n11241), .B(n11242), .Z(n11235) );
  NOR U11099 ( .A(n11243), .B(n11244), .Z(n11242) );
  XOR U11100 ( .A(n11241), .B(n11245), .Z(n11243) );
  XNOR U11101 ( .A(n11204), .B(n11211), .Z(n11223) );
  NOR U11102 ( .A(n11172), .B(n11246), .Z(n11211) );
  XOR U11103 ( .A(n11216), .B(n11215), .Z(n11204) );
  XNOR U11104 ( .A(n11247), .B(n11212), .Z(n11215) );
  XOR U11105 ( .A(n11248), .B(n11249), .Z(n11212) );
  AND U11106 ( .A(n11250), .B(n11251), .Z(n11249) );
  XOR U11107 ( .A(n11248), .B(n11252), .Z(n11250) );
  XNOR U11108 ( .A(n11253), .B(n11254), .Z(n11247) );
  NOR U11109 ( .A(n11255), .B(n11256), .Z(n11254) );
  XNOR U11110 ( .A(n11253), .B(n11257), .Z(n11255) );
  XOR U11111 ( .A(n11258), .B(n11259), .Z(n11216) );
  NOR U11112 ( .A(n11260), .B(n11261), .Z(n11259) );
  XNOR U11113 ( .A(n11258), .B(n11262), .Z(n11260) );
  XNOR U11114 ( .A(n11161), .B(n11219), .Z(n11221) );
  XNOR U11115 ( .A(n11263), .B(n11264), .Z(n11161) );
  AND U11116 ( .A(n237), .B(n11168), .Z(n11264) );
  XOR U11117 ( .A(n11263), .B(n11166), .Z(n11168) );
  AND U11118 ( .A(n11169), .B(n11172), .Z(n11219) );
  XOR U11119 ( .A(n11265), .B(n11246), .Z(n11172) );
  XNOR U11120 ( .A(p_input[1024]), .B(p_input[288]), .Z(n11246) );
  XOR U11121 ( .A(n11234), .B(n11233), .Z(n11265) );
  XNOR U11122 ( .A(n11266), .B(n11240), .Z(n11233) );
  XNOR U11123 ( .A(n11229), .B(n11228), .Z(n11240) );
  XOR U11124 ( .A(n11267), .B(n11225), .Z(n11228) );
  XOR U11125 ( .A(p_input[1034]), .B(p_input[298]), .Z(n11225) );
  XNOR U11126 ( .A(p_input[1035]), .B(p_input[299]), .Z(n11267) );
  XOR U11127 ( .A(p_input[1036]), .B(p_input[300]), .Z(n11229) );
  XNOR U11128 ( .A(n11239), .B(n11230), .Z(n11266) );
  XOR U11129 ( .A(p_input[1025]), .B(p_input[289]), .Z(n11230) );
  XOR U11130 ( .A(n11268), .B(n11245), .Z(n11239) );
  XNOR U11131 ( .A(p_input[1039]), .B(p_input[303]), .Z(n11245) );
  XOR U11132 ( .A(n11236), .B(n11244), .Z(n11268) );
  XOR U11133 ( .A(n11269), .B(n11241), .Z(n11244) );
  XOR U11134 ( .A(p_input[1037]), .B(p_input[301]), .Z(n11241) );
  XNOR U11135 ( .A(p_input[1038]), .B(p_input[302]), .Z(n11269) );
  XOR U11136 ( .A(p_input[1033]), .B(p_input[297]), .Z(n11236) );
  XNOR U11137 ( .A(n11252), .B(n11251), .Z(n11234) );
  XNOR U11138 ( .A(n11270), .B(n11257), .Z(n11251) );
  XOR U11139 ( .A(p_input[1032]), .B(p_input[296]), .Z(n11257) );
  XOR U11140 ( .A(n11248), .B(n11256), .Z(n11270) );
  XOR U11141 ( .A(n11271), .B(n11253), .Z(n11256) );
  XOR U11142 ( .A(p_input[1030]), .B(p_input[294]), .Z(n11253) );
  XNOR U11143 ( .A(p_input[1031]), .B(p_input[295]), .Z(n11271) );
  XOR U11144 ( .A(p_input[1026]), .B(p_input[290]), .Z(n11248) );
  XNOR U11145 ( .A(n11262), .B(n11261), .Z(n11252) );
  XOR U11146 ( .A(n11272), .B(n11258), .Z(n11261) );
  XOR U11147 ( .A(p_input[1027]), .B(p_input[291]), .Z(n11258) );
  XNOR U11148 ( .A(p_input[1028]), .B(p_input[292]), .Z(n11272) );
  XOR U11149 ( .A(p_input[1029]), .B(p_input[293]), .Z(n11262) );
  XNOR U11150 ( .A(n11273), .B(n11274), .Z(n11169) );
  AND U11151 ( .A(n237), .B(n11275), .Z(n11274) );
  XNOR U11152 ( .A(n11276), .B(n11277), .Z(n237) );
  AND U11153 ( .A(n11278), .B(n11279), .Z(n11277) );
  XOR U11154 ( .A(n11276), .B(n11179), .Z(n11279) );
  XNOR U11155 ( .A(n11276), .B(n11133), .Z(n11278) );
  XOR U11156 ( .A(n11280), .B(n11281), .Z(n11276) );
  AND U11157 ( .A(n11282), .B(n11283), .Z(n11281) );
  XOR U11158 ( .A(n11280), .B(n11143), .Z(n11282) );
  XOR U11159 ( .A(n11284), .B(n11285), .Z(n11122) );
  AND U11160 ( .A(n241), .B(n11275), .Z(n11285) );
  XNOR U11161 ( .A(n11273), .B(n11284), .Z(n11275) );
  XNOR U11162 ( .A(n11286), .B(n11287), .Z(n241) );
  AND U11163 ( .A(n11288), .B(n11289), .Z(n11287) );
  XNOR U11164 ( .A(n11290), .B(n11286), .Z(n11289) );
  IV U11165 ( .A(n11179), .Z(n11290) );
  XNOR U11166 ( .A(n11291), .B(n11292), .Z(n11179) );
  AND U11167 ( .A(n244), .B(n11293), .Z(n11292) );
  XNOR U11168 ( .A(n11291), .B(n11294), .Z(n11293) );
  XNOR U11169 ( .A(n11133), .B(n11286), .Z(n11288) );
  XOR U11170 ( .A(n11295), .B(n11296), .Z(n11133) );
  AND U11171 ( .A(n252), .B(n11297), .Z(n11296) );
  XOR U11172 ( .A(n11280), .B(n11298), .Z(n11286) );
  AND U11173 ( .A(n11299), .B(n11283), .Z(n11298) );
  XNOR U11174 ( .A(n11192), .B(n11280), .Z(n11283) );
  XNOR U11175 ( .A(n11300), .B(n11301), .Z(n11192) );
  AND U11176 ( .A(n244), .B(n11302), .Z(n11301) );
  XOR U11177 ( .A(n11303), .B(n11300), .Z(n11302) );
  XNOR U11178 ( .A(n11304), .B(n11280), .Z(n11299) );
  IV U11179 ( .A(n11143), .Z(n11304) );
  XOR U11180 ( .A(n11305), .B(n11306), .Z(n11143) );
  AND U11181 ( .A(n252), .B(n11307), .Z(n11306) );
  XOR U11182 ( .A(n11308), .B(n11309), .Z(n11280) );
  AND U11183 ( .A(n11310), .B(n11311), .Z(n11309) );
  XNOR U11184 ( .A(n11217), .B(n11308), .Z(n11311) );
  XNOR U11185 ( .A(n11312), .B(n11313), .Z(n11217) );
  AND U11186 ( .A(n244), .B(n11314), .Z(n11313) );
  XNOR U11187 ( .A(n11315), .B(n11312), .Z(n11314) );
  XOR U11188 ( .A(n11308), .B(n11154), .Z(n11310) );
  XOR U11189 ( .A(n11316), .B(n11317), .Z(n11154) );
  AND U11190 ( .A(n252), .B(n11318), .Z(n11317) );
  XOR U11191 ( .A(n11319), .B(n11320), .Z(n11308) );
  AND U11192 ( .A(n11321), .B(n11322), .Z(n11320) );
  XNOR U11193 ( .A(n11319), .B(n11263), .Z(n11322) );
  XNOR U11194 ( .A(n11323), .B(n11324), .Z(n11263) );
  AND U11195 ( .A(n244), .B(n11325), .Z(n11324) );
  XOR U11196 ( .A(n11326), .B(n11323), .Z(n11325) );
  XNOR U11197 ( .A(n11327), .B(n11319), .Z(n11321) );
  IV U11198 ( .A(n11166), .Z(n11327) );
  XOR U11199 ( .A(n11328), .B(n11329), .Z(n11166) );
  AND U11200 ( .A(n252), .B(n11330), .Z(n11329) );
  AND U11201 ( .A(n11284), .B(n11273), .Z(n11319) );
  XNOR U11202 ( .A(n11331), .B(n11332), .Z(n11273) );
  AND U11203 ( .A(n244), .B(n11333), .Z(n11332) );
  XNOR U11204 ( .A(n11334), .B(n11331), .Z(n11333) );
  XNOR U11205 ( .A(n11335), .B(n11336), .Z(n244) );
  AND U11206 ( .A(n11337), .B(n11338), .Z(n11336) );
  XOR U11207 ( .A(n11294), .B(n11335), .Z(n11338) );
  AND U11208 ( .A(n11339), .B(n11340), .Z(n11294) );
  XOR U11209 ( .A(n11335), .B(n11291), .Z(n11337) );
  XNOR U11210 ( .A(n11341), .B(n11342), .Z(n11291) );
  AND U11211 ( .A(n248), .B(n11297), .Z(n11342) );
  XOR U11212 ( .A(n11295), .B(n11341), .Z(n11297) );
  XOR U11213 ( .A(n11343), .B(n11344), .Z(n11335) );
  AND U11214 ( .A(n11345), .B(n11346), .Z(n11344) );
  XNOR U11215 ( .A(n11343), .B(n11339), .Z(n11346) );
  IV U11216 ( .A(n11303), .Z(n11339) );
  XOR U11217 ( .A(n11347), .B(n11348), .Z(n11303) );
  XOR U11218 ( .A(n11349), .B(n11340), .Z(n11348) );
  AND U11219 ( .A(n11315), .B(n11350), .Z(n11340) );
  AND U11220 ( .A(n11351), .B(n11352), .Z(n11349) );
  XOR U11221 ( .A(n11353), .B(n11347), .Z(n11351) );
  XNOR U11222 ( .A(n11300), .B(n11343), .Z(n11345) );
  XNOR U11223 ( .A(n11354), .B(n11355), .Z(n11300) );
  AND U11224 ( .A(n248), .B(n11307), .Z(n11355) );
  XOR U11225 ( .A(n11354), .B(n11305), .Z(n11307) );
  XOR U11226 ( .A(n11356), .B(n11357), .Z(n11343) );
  AND U11227 ( .A(n11358), .B(n11359), .Z(n11357) );
  XNOR U11228 ( .A(n11356), .B(n11315), .Z(n11359) );
  XOR U11229 ( .A(n11360), .B(n11352), .Z(n11315) );
  XNOR U11230 ( .A(n11361), .B(n11347), .Z(n11352) );
  XOR U11231 ( .A(n11362), .B(n11363), .Z(n11347) );
  AND U11232 ( .A(n11364), .B(n11365), .Z(n11363) );
  XOR U11233 ( .A(n11366), .B(n11362), .Z(n11364) );
  XNOR U11234 ( .A(n11367), .B(n11368), .Z(n11361) );
  AND U11235 ( .A(n11369), .B(n11370), .Z(n11368) );
  XOR U11236 ( .A(n11367), .B(n11371), .Z(n11369) );
  XNOR U11237 ( .A(n11353), .B(n11350), .Z(n11360) );
  AND U11238 ( .A(n11372), .B(n11373), .Z(n11350) );
  XOR U11239 ( .A(n11374), .B(n11375), .Z(n11353) );
  AND U11240 ( .A(n11376), .B(n11377), .Z(n11375) );
  XOR U11241 ( .A(n11374), .B(n11378), .Z(n11376) );
  XNOR U11242 ( .A(n11312), .B(n11356), .Z(n11358) );
  XNOR U11243 ( .A(n11379), .B(n11380), .Z(n11312) );
  AND U11244 ( .A(n248), .B(n11318), .Z(n11380) );
  XOR U11245 ( .A(n11379), .B(n11316), .Z(n11318) );
  XOR U11246 ( .A(n11381), .B(n11382), .Z(n11356) );
  AND U11247 ( .A(n11383), .B(n11384), .Z(n11382) );
  XNOR U11248 ( .A(n11381), .B(n11372), .Z(n11384) );
  IV U11249 ( .A(n11326), .Z(n11372) );
  XNOR U11250 ( .A(n11385), .B(n11365), .Z(n11326) );
  XNOR U11251 ( .A(n11386), .B(n11371), .Z(n11365) );
  XOR U11252 ( .A(n11387), .B(n11388), .Z(n11371) );
  NOR U11253 ( .A(n11389), .B(n11390), .Z(n11388) );
  XNOR U11254 ( .A(n11387), .B(n11391), .Z(n11389) );
  XNOR U11255 ( .A(n11370), .B(n11362), .Z(n11386) );
  XOR U11256 ( .A(n11392), .B(n11393), .Z(n11362) );
  AND U11257 ( .A(n11394), .B(n11395), .Z(n11393) );
  XNOR U11258 ( .A(n11392), .B(n11396), .Z(n11394) );
  XNOR U11259 ( .A(n11397), .B(n11367), .Z(n11370) );
  XOR U11260 ( .A(n11398), .B(n11399), .Z(n11367) );
  AND U11261 ( .A(n11400), .B(n11401), .Z(n11399) );
  XOR U11262 ( .A(n11398), .B(n11402), .Z(n11400) );
  XNOR U11263 ( .A(n11403), .B(n11404), .Z(n11397) );
  NOR U11264 ( .A(n11405), .B(n11406), .Z(n11404) );
  XOR U11265 ( .A(n11403), .B(n11407), .Z(n11405) );
  XNOR U11266 ( .A(n11366), .B(n11373), .Z(n11385) );
  NOR U11267 ( .A(n11334), .B(n11408), .Z(n11373) );
  XOR U11268 ( .A(n11378), .B(n11377), .Z(n11366) );
  XNOR U11269 ( .A(n11409), .B(n11374), .Z(n11377) );
  XOR U11270 ( .A(n11410), .B(n11411), .Z(n11374) );
  AND U11271 ( .A(n11412), .B(n11413), .Z(n11411) );
  XOR U11272 ( .A(n11410), .B(n11414), .Z(n11412) );
  XNOR U11273 ( .A(n11415), .B(n11416), .Z(n11409) );
  NOR U11274 ( .A(n11417), .B(n11418), .Z(n11416) );
  XNOR U11275 ( .A(n11415), .B(n11419), .Z(n11417) );
  XOR U11276 ( .A(n11420), .B(n11421), .Z(n11378) );
  NOR U11277 ( .A(n11422), .B(n11423), .Z(n11421) );
  XNOR U11278 ( .A(n11420), .B(n11424), .Z(n11422) );
  XNOR U11279 ( .A(n11323), .B(n11381), .Z(n11383) );
  XNOR U11280 ( .A(n11425), .B(n11426), .Z(n11323) );
  AND U11281 ( .A(n248), .B(n11330), .Z(n11426) );
  XOR U11282 ( .A(n11425), .B(n11328), .Z(n11330) );
  AND U11283 ( .A(n11331), .B(n11334), .Z(n11381) );
  XOR U11284 ( .A(n11427), .B(n11408), .Z(n11334) );
  XNOR U11285 ( .A(p_input[1024]), .B(p_input[304]), .Z(n11408) );
  XOR U11286 ( .A(n11396), .B(n11395), .Z(n11427) );
  XNOR U11287 ( .A(n11428), .B(n11402), .Z(n11395) );
  XNOR U11288 ( .A(n11391), .B(n11390), .Z(n11402) );
  XOR U11289 ( .A(n11429), .B(n11387), .Z(n11390) );
  XOR U11290 ( .A(p_input[1034]), .B(p_input[314]), .Z(n11387) );
  XNOR U11291 ( .A(p_input[1035]), .B(p_input[315]), .Z(n11429) );
  XOR U11292 ( .A(p_input[1036]), .B(p_input[316]), .Z(n11391) );
  XNOR U11293 ( .A(n11401), .B(n11392), .Z(n11428) );
  XOR U11294 ( .A(p_input[1025]), .B(p_input[305]), .Z(n11392) );
  XOR U11295 ( .A(n11430), .B(n11407), .Z(n11401) );
  XNOR U11296 ( .A(p_input[1039]), .B(p_input[319]), .Z(n11407) );
  XOR U11297 ( .A(n11398), .B(n11406), .Z(n11430) );
  XOR U11298 ( .A(n11431), .B(n11403), .Z(n11406) );
  XOR U11299 ( .A(p_input[1037]), .B(p_input[317]), .Z(n11403) );
  XNOR U11300 ( .A(p_input[1038]), .B(p_input[318]), .Z(n11431) );
  XOR U11301 ( .A(p_input[1033]), .B(p_input[313]), .Z(n11398) );
  XNOR U11302 ( .A(n11414), .B(n11413), .Z(n11396) );
  XNOR U11303 ( .A(n11432), .B(n11419), .Z(n11413) );
  XOR U11304 ( .A(p_input[1032]), .B(p_input[312]), .Z(n11419) );
  XOR U11305 ( .A(n11410), .B(n11418), .Z(n11432) );
  XOR U11306 ( .A(n11433), .B(n11415), .Z(n11418) );
  XOR U11307 ( .A(p_input[1030]), .B(p_input[310]), .Z(n11415) );
  XNOR U11308 ( .A(p_input[1031]), .B(p_input[311]), .Z(n11433) );
  XOR U11309 ( .A(p_input[1026]), .B(p_input[306]), .Z(n11410) );
  XNOR U11310 ( .A(n11424), .B(n11423), .Z(n11414) );
  XOR U11311 ( .A(n11434), .B(n11420), .Z(n11423) );
  XOR U11312 ( .A(p_input[1027]), .B(p_input[307]), .Z(n11420) );
  XNOR U11313 ( .A(p_input[1028]), .B(p_input[308]), .Z(n11434) );
  XOR U11314 ( .A(p_input[1029]), .B(p_input[309]), .Z(n11424) );
  XNOR U11315 ( .A(n11435), .B(n11436), .Z(n11331) );
  AND U11316 ( .A(n248), .B(n11437), .Z(n11436) );
  XNOR U11317 ( .A(n11438), .B(n11439), .Z(n248) );
  AND U11318 ( .A(n11440), .B(n11441), .Z(n11439) );
  XOR U11319 ( .A(n11438), .B(n11341), .Z(n11441) );
  XNOR U11320 ( .A(n11438), .B(n11295), .Z(n11440) );
  XOR U11321 ( .A(n11442), .B(n11443), .Z(n11438) );
  AND U11322 ( .A(n11444), .B(n11445), .Z(n11443) );
  XOR U11323 ( .A(n11442), .B(n11305), .Z(n11444) );
  XOR U11324 ( .A(n11446), .B(n11447), .Z(n11284) );
  AND U11325 ( .A(n252), .B(n11437), .Z(n11447) );
  XNOR U11326 ( .A(n11435), .B(n11446), .Z(n11437) );
  XNOR U11327 ( .A(n11448), .B(n11449), .Z(n252) );
  AND U11328 ( .A(n11450), .B(n11451), .Z(n11449) );
  XNOR U11329 ( .A(n11452), .B(n11448), .Z(n11451) );
  IV U11330 ( .A(n11341), .Z(n11452) );
  XNOR U11331 ( .A(n11453), .B(n11454), .Z(n11341) );
  AND U11332 ( .A(n255), .B(n11455), .Z(n11454) );
  XNOR U11333 ( .A(n11453), .B(n11456), .Z(n11455) );
  XNOR U11334 ( .A(n11295), .B(n11448), .Z(n11450) );
  XOR U11335 ( .A(n11457), .B(n11458), .Z(n11295) );
  AND U11336 ( .A(n263), .B(n11459), .Z(n11458) );
  XOR U11337 ( .A(n11442), .B(n11460), .Z(n11448) );
  AND U11338 ( .A(n11461), .B(n11445), .Z(n11460) );
  XNOR U11339 ( .A(n11354), .B(n11442), .Z(n11445) );
  XNOR U11340 ( .A(n11462), .B(n11463), .Z(n11354) );
  AND U11341 ( .A(n255), .B(n11464), .Z(n11463) );
  XOR U11342 ( .A(n11465), .B(n11462), .Z(n11464) );
  XNOR U11343 ( .A(n11466), .B(n11442), .Z(n11461) );
  IV U11344 ( .A(n11305), .Z(n11466) );
  XOR U11345 ( .A(n11467), .B(n11468), .Z(n11305) );
  AND U11346 ( .A(n263), .B(n11469), .Z(n11468) );
  XOR U11347 ( .A(n11470), .B(n11471), .Z(n11442) );
  AND U11348 ( .A(n11472), .B(n11473), .Z(n11471) );
  XNOR U11349 ( .A(n11379), .B(n11470), .Z(n11473) );
  XNOR U11350 ( .A(n11474), .B(n11475), .Z(n11379) );
  AND U11351 ( .A(n255), .B(n11476), .Z(n11475) );
  XNOR U11352 ( .A(n11477), .B(n11474), .Z(n11476) );
  XOR U11353 ( .A(n11470), .B(n11316), .Z(n11472) );
  XOR U11354 ( .A(n11478), .B(n11479), .Z(n11316) );
  AND U11355 ( .A(n263), .B(n11480), .Z(n11479) );
  XOR U11356 ( .A(n11481), .B(n11482), .Z(n11470) );
  AND U11357 ( .A(n11483), .B(n11484), .Z(n11482) );
  XNOR U11358 ( .A(n11481), .B(n11425), .Z(n11484) );
  XNOR U11359 ( .A(n11485), .B(n11486), .Z(n11425) );
  AND U11360 ( .A(n255), .B(n11487), .Z(n11486) );
  XOR U11361 ( .A(n11488), .B(n11485), .Z(n11487) );
  XNOR U11362 ( .A(n11489), .B(n11481), .Z(n11483) );
  IV U11363 ( .A(n11328), .Z(n11489) );
  XOR U11364 ( .A(n11490), .B(n11491), .Z(n11328) );
  AND U11365 ( .A(n263), .B(n11492), .Z(n11491) );
  AND U11366 ( .A(n11446), .B(n11435), .Z(n11481) );
  XNOR U11367 ( .A(n11493), .B(n11494), .Z(n11435) );
  AND U11368 ( .A(n255), .B(n11495), .Z(n11494) );
  XNOR U11369 ( .A(n11496), .B(n11493), .Z(n11495) );
  XNOR U11370 ( .A(n11497), .B(n11498), .Z(n255) );
  AND U11371 ( .A(n11499), .B(n11500), .Z(n11498) );
  XOR U11372 ( .A(n11456), .B(n11497), .Z(n11500) );
  AND U11373 ( .A(n11501), .B(n11502), .Z(n11456) );
  XOR U11374 ( .A(n11497), .B(n11453), .Z(n11499) );
  XNOR U11375 ( .A(n11503), .B(n11504), .Z(n11453) );
  AND U11376 ( .A(n259), .B(n11459), .Z(n11504) );
  XOR U11377 ( .A(n11457), .B(n11503), .Z(n11459) );
  XOR U11378 ( .A(n11505), .B(n11506), .Z(n11497) );
  AND U11379 ( .A(n11507), .B(n11508), .Z(n11506) );
  XNOR U11380 ( .A(n11505), .B(n11501), .Z(n11508) );
  IV U11381 ( .A(n11465), .Z(n11501) );
  XOR U11382 ( .A(n11509), .B(n11510), .Z(n11465) );
  XOR U11383 ( .A(n11511), .B(n11502), .Z(n11510) );
  AND U11384 ( .A(n11477), .B(n11512), .Z(n11502) );
  AND U11385 ( .A(n11513), .B(n11514), .Z(n11511) );
  XOR U11386 ( .A(n11515), .B(n11509), .Z(n11513) );
  XNOR U11387 ( .A(n11462), .B(n11505), .Z(n11507) );
  XNOR U11388 ( .A(n11516), .B(n11517), .Z(n11462) );
  AND U11389 ( .A(n259), .B(n11469), .Z(n11517) );
  XOR U11390 ( .A(n11516), .B(n11467), .Z(n11469) );
  XOR U11391 ( .A(n11518), .B(n11519), .Z(n11505) );
  AND U11392 ( .A(n11520), .B(n11521), .Z(n11519) );
  XNOR U11393 ( .A(n11518), .B(n11477), .Z(n11521) );
  XOR U11394 ( .A(n11522), .B(n11514), .Z(n11477) );
  XNOR U11395 ( .A(n11523), .B(n11509), .Z(n11514) );
  XOR U11396 ( .A(n11524), .B(n11525), .Z(n11509) );
  AND U11397 ( .A(n11526), .B(n11527), .Z(n11525) );
  XOR U11398 ( .A(n11528), .B(n11524), .Z(n11526) );
  XNOR U11399 ( .A(n11529), .B(n11530), .Z(n11523) );
  AND U11400 ( .A(n11531), .B(n11532), .Z(n11530) );
  XOR U11401 ( .A(n11529), .B(n11533), .Z(n11531) );
  XNOR U11402 ( .A(n11515), .B(n11512), .Z(n11522) );
  AND U11403 ( .A(n11534), .B(n11535), .Z(n11512) );
  XOR U11404 ( .A(n11536), .B(n11537), .Z(n11515) );
  AND U11405 ( .A(n11538), .B(n11539), .Z(n11537) );
  XOR U11406 ( .A(n11536), .B(n11540), .Z(n11538) );
  XNOR U11407 ( .A(n11474), .B(n11518), .Z(n11520) );
  XNOR U11408 ( .A(n11541), .B(n11542), .Z(n11474) );
  AND U11409 ( .A(n259), .B(n11480), .Z(n11542) );
  XOR U11410 ( .A(n11541), .B(n11478), .Z(n11480) );
  XOR U11411 ( .A(n11543), .B(n11544), .Z(n11518) );
  AND U11412 ( .A(n11545), .B(n11546), .Z(n11544) );
  XNOR U11413 ( .A(n11543), .B(n11534), .Z(n11546) );
  IV U11414 ( .A(n11488), .Z(n11534) );
  XNOR U11415 ( .A(n11547), .B(n11527), .Z(n11488) );
  XNOR U11416 ( .A(n11548), .B(n11533), .Z(n11527) );
  XOR U11417 ( .A(n11549), .B(n11550), .Z(n11533) );
  NOR U11418 ( .A(n11551), .B(n11552), .Z(n11550) );
  XNOR U11419 ( .A(n11549), .B(n11553), .Z(n11551) );
  XNOR U11420 ( .A(n11532), .B(n11524), .Z(n11548) );
  XOR U11421 ( .A(n11554), .B(n11555), .Z(n11524) );
  AND U11422 ( .A(n11556), .B(n11557), .Z(n11555) );
  XNOR U11423 ( .A(n11554), .B(n11558), .Z(n11556) );
  XNOR U11424 ( .A(n11559), .B(n11529), .Z(n11532) );
  XOR U11425 ( .A(n11560), .B(n11561), .Z(n11529) );
  AND U11426 ( .A(n11562), .B(n11563), .Z(n11561) );
  XOR U11427 ( .A(n11560), .B(n11564), .Z(n11562) );
  XNOR U11428 ( .A(n11565), .B(n11566), .Z(n11559) );
  NOR U11429 ( .A(n11567), .B(n11568), .Z(n11566) );
  XOR U11430 ( .A(n11565), .B(n11569), .Z(n11567) );
  XNOR U11431 ( .A(n11528), .B(n11535), .Z(n11547) );
  NOR U11432 ( .A(n11496), .B(n11570), .Z(n11535) );
  XOR U11433 ( .A(n11540), .B(n11539), .Z(n11528) );
  XNOR U11434 ( .A(n11571), .B(n11536), .Z(n11539) );
  XOR U11435 ( .A(n11572), .B(n11573), .Z(n11536) );
  AND U11436 ( .A(n11574), .B(n11575), .Z(n11573) );
  XOR U11437 ( .A(n11572), .B(n11576), .Z(n11574) );
  XNOR U11438 ( .A(n11577), .B(n11578), .Z(n11571) );
  NOR U11439 ( .A(n11579), .B(n11580), .Z(n11578) );
  XNOR U11440 ( .A(n11577), .B(n11581), .Z(n11579) );
  XOR U11441 ( .A(n11582), .B(n11583), .Z(n11540) );
  NOR U11442 ( .A(n11584), .B(n11585), .Z(n11583) );
  XNOR U11443 ( .A(n11582), .B(n11586), .Z(n11584) );
  XNOR U11444 ( .A(n11485), .B(n11543), .Z(n11545) );
  XNOR U11445 ( .A(n11587), .B(n11588), .Z(n11485) );
  AND U11446 ( .A(n259), .B(n11492), .Z(n11588) );
  XOR U11447 ( .A(n11587), .B(n11490), .Z(n11492) );
  AND U11448 ( .A(n11493), .B(n11496), .Z(n11543) );
  XOR U11449 ( .A(n11589), .B(n11570), .Z(n11496) );
  XNOR U11450 ( .A(p_input[1024]), .B(p_input[320]), .Z(n11570) );
  XOR U11451 ( .A(n11558), .B(n11557), .Z(n11589) );
  XNOR U11452 ( .A(n11590), .B(n11564), .Z(n11557) );
  XNOR U11453 ( .A(n11553), .B(n11552), .Z(n11564) );
  XOR U11454 ( .A(n11591), .B(n11549), .Z(n11552) );
  XOR U11455 ( .A(p_input[1034]), .B(p_input[330]), .Z(n11549) );
  XNOR U11456 ( .A(p_input[1035]), .B(p_input[331]), .Z(n11591) );
  XOR U11457 ( .A(p_input[1036]), .B(p_input[332]), .Z(n11553) );
  XNOR U11458 ( .A(n11563), .B(n11554), .Z(n11590) );
  XOR U11459 ( .A(p_input[1025]), .B(p_input[321]), .Z(n11554) );
  XOR U11460 ( .A(n11592), .B(n11569), .Z(n11563) );
  XNOR U11461 ( .A(p_input[1039]), .B(p_input[335]), .Z(n11569) );
  XOR U11462 ( .A(n11560), .B(n11568), .Z(n11592) );
  XOR U11463 ( .A(n11593), .B(n11565), .Z(n11568) );
  XOR U11464 ( .A(p_input[1037]), .B(p_input[333]), .Z(n11565) );
  XNOR U11465 ( .A(p_input[1038]), .B(p_input[334]), .Z(n11593) );
  XOR U11466 ( .A(p_input[1033]), .B(p_input[329]), .Z(n11560) );
  XNOR U11467 ( .A(n11576), .B(n11575), .Z(n11558) );
  XNOR U11468 ( .A(n11594), .B(n11581), .Z(n11575) );
  XOR U11469 ( .A(p_input[1032]), .B(p_input[328]), .Z(n11581) );
  XOR U11470 ( .A(n11572), .B(n11580), .Z(n11594) );
  XOR U11471 ( .A(n11595), .B(n11577), .Z(n11580) );
  XOR U11472 ( .A(p_input[1030]), .B(p_input[326]), .Z(n11577) );
  XNOR U11473 ( .A(p_input[1031]), .B(p_input[327]), .Z(n11595) );
  XOR U11474 ( .A(p_input[1026]), .B(p_input[322]), .Z(n11572) );
  XNOR U11475 ( .A(n11586), .B(n11585), .Z(n11576) );
  XOR U11476 ( .A(n11596), .B(n11582), .Z(n11585) );
  XOR U11477 ( .A(p_input[1027]), .B(p_input[323]), .Z(n11582) );
  XNOR U11478 ( .A(p_input[1028]), .B(p_input[324]), .Z(n11596) );
  XOR U11479 ( .A(p_input[1029]), .B(p_input[325]), .Z(n11586) );
  XNOR U11480 ( .A(n11597), .B(n11598), .Z(n11493) );
  AND U11481 ( .A(n259), .B(n11599), .Z(n11598) );
  XNOR U11482 ( .A(n11600), .B(n11601), .Z(n259) );
  AND U11483 ( .A(n11602), .B(n11603), .Z(n11601) );
  XOR U11484 ( .A(n11600), .B(n11503), .Z(n11603) );
  XNOR U11485 ( .A(n11600), .B(n11457), .Z(n11602) );
  XOR U11486 ( .A(n11604), .B(n11605), .Z(n11600) );
  AND U11487 ( .A(n11606), .B(n11607), .Z(n11605) );
  XOR U11488 ( .A(n11604), .B(n11467), .Z(n11606) );
  XOR U11489 ( .A(n11608), .B(n11609), .Z(n11446) );
  AND U11490 ( .A(n263), .B(n11599), .Z(n11609) );
  XNOR U11491 ( .A(n11597), .B(n11608), .Z(n11599) );
  XNOR U11492 ( .A(n11610), .B(n11611), .Z(n263) );
  AND U11493 ( .A(n11612), .B(n11613), .Z(n11611) );
  XNOR U11494 ( .A(n11614), .B(n11610), .Z(n11613) );
  IV U11495 ( .A(n11503), .Z(n11614) );
  XNOR U11496 ( .A(n11615), .B(n11616), .Z(n11503) );
  AND U11497 ( .A(n266), .B(n11617), .Z(n11616) );
  XNOR U11498 ( .A(n11615), .B(n11618), .Z(n11617) );
  XNOR U11499 ( .A(n11457), .B(n11610), .Z(n11612) );
  XOR U11500 ( .A(n11619), .B(n11620), .Z(n11457) );
  AND U11501 ( .A(n274), .B(n11621), .Z(n11620) );
  XOR U11502 ( .A(n11604), .B(n11622), .Z(n11610) );
  AND U11503 ( .A(n11623), .B(n11607), .Z(n11622) );
  XNOR U11504 ( .A(n11516), .B(n11604), .Z(n11607) );
  XNOR U11505 ( .A(n11624), .B(n11625), .Z(n11516) );
  AND U11506 ( .A(n266), .B(n11626), .Z(n11625) );
  XOR U11507 ( .A(n11627), .B(n11624), .Z(n11626) );
  XNOR U11508 ( .A(n11628), .B(n11604), .Z(n11623) );
  IV U11509 ( .A(n11467), .Z(n11628) );
  XOR U11510 ( .A(n11629), .B(n11630), .Z(n11467) );
  AND U11511 ( .A(n274), .B(n11631), .Z(n11630) );
  XOR U11512 ( .A(n11632), .B(n11633), .Z(n11604) );
  AND U11513 ( .A(n11634), .B(n11635), .Z(n11633) );
  XNOR U11514 ( .A(n11541), .B(n11632), .Z(n11635) );
  XNOR U11515 ( .A(n11636), .B(n11637), .Z(n11541) );
  AND U11516 ( .A(n266), .B(n11638), .Z(n11637) );
  XNOR U11517 ( .A(n11639), .B(n11636), .Z(n11638) );
  XOR U11518 ( .A(n11632), .B(n11478), .Z(n11634) );
  XOR U11519 ( .A(n11640), .B(n11641), .Z(n11478) );
  AND U11520 ( .A(n274), .B(n11642), .Z(n11641) );
  XOR U11521 ( .A(n11643), .B(n11644), .Z(n11632) );
  AND U11522 ( .A(n11645), .B(n11646), .Z(n11644) );
  XNOR U11523 ( .A(n11643), .B(n11587), .Z(n11646) );
  XNOR U11524 ( .A(n11647), .B(n11648), .Z(n11587) );
  AND U11525 ( .A(n266), .B(n11649), .Z(n11648) );
  XOR U11526 ( .A(n11650), .B(n11647), .Z(n11649) );
  XNOR U11527 ( .A(n11651), .B(n11643), .Z(n11645) );
  IV U11528 ( .A(n11490), .Z(n11651) );
  XOR U11529 ( .A(n11652), .B(n11653), .Z(n11490) );
  AND U11530 ( .A(n274), .B(n11654), .Z(n11653) );
  AND U11531 ( .A(n11608), .B(n11597), .Z(n11643) );
  XNOR U11532 ( .A(n11655), .B(n11656), .Z(n11597) );
  AND U11533 ( .A(n266), .B(n11657), .Z(n11656) );
  XNOR U11534 ( .A(n11658), .B(n11655), .Z(n11657) );
  XNOR U11535 ( .A(n11659), .B(n11660), .Z(n266) );
  AND U11536 ( .A(n11661), .B(n11662), .Z(n11660) );
  XOR U11537 ( .A(n11618), .B(n11659), .Z(n11662) );
  AND U11538 ( .A(n11663), .B(n11664), .Z(n11618) );
  XOR U11539 ( .A(n11659), .B(n11615), .Z(n11661) );
  XNOR U11540 ( .A(n11665), .B(n11666), .Z(n11615) );
  AND U11541 ( .A(n270), .B(n11621), .Z(n11666) );
  XOR U11542 ( .A(n11619), .B(n11665), .Z(n11621) );
  XOR U11543 ( .A(n11667), .B(n11668), .Z(n11659) );
  AND U11544 ( .A(n11669), .B(n11670), .Z(n11668) );
  XNOR U11545 ( .A(n11667), .B(n11663), .Z(n11670) );
  IV U11546 ( .A(n11627), .Z(n11663) );
  XOR U11547 ( .A(n11671), .B(n11672), .Z(n11627) );
  XOR U11548 ( .A(n11673), .B(n11664), .Z(n11672) );
  AND U11549 ( .A(n11639), .B(n11674), .Z(n11664) );
  AND U11550 ( .A(n11675), .B(n11676), .Z(n11673) );
  XOR U11551 ( .A(n11677), .B(n11671), .Z(n11675) );
  XNOR U11552 ( .A(n11624), .B(n11667), .Z(n11669) );
  XNOR U11553 ( .A(n11678), .B(n11679), .Z(n11624) );
  AND U11554 ( .A(n270), .B(n11631), .Z(n11679) );
  XOR U11555 ( .A(n11678), .B(n11629), .Z(n11631) );
  XOR U11556 ( .A(n11680), .B(n11681), .Z(n11667) );
  AND U11557 ( .A(n11682), .B(n11683), .Z(n11681) );
  XNOR U11558 ( .A(n11680), .B(n11639), .Z(n11683) );
  XOR U11559 ( .A(n11684), .B(n11676), .Z(n11639) );
  XNOR U11560 ( .A(n11685), .B(n11671), .Z(n11676) );
  XOR U11561 ( .A(n11686), .B(n11687), .Z(n11671) );
  AND U11562 ( .A(n11688), .B(n11689), .Z(n11687) );
  XOR U11563 ( .A(n11690), .B(n11686), .Z(n11688) );
  XNOR U11564 ( .A(n11691), .B(n11692), .Z(n11685) );
  AND U11565 ( .A(n11693), .B(n11694), .Z(n11692) );
  XOR U11566 ( .A(n11691), .B(n11695), .Z(n11693) );
  XNOR U11567 ( .A(n11677), .B(n11674), .Z(n11684) );
  AND U11568 ( .A(n11696), .B(n11697), .Z(n11674) );
  XOR U11569 ( .A(n11698), .B(n11699), .Z(n11677) );
  AND U11570 ( .A(n11700), .B(n11701), .Z(n11699) );
  XOR U11571 ( .A(n11698), .B(n11702), .Z(n11700) );
  XNOR U11572 ( .A(n11636), .B(n11680), .Z(n11682) );
  XNOR U11573 ( .A(n11703), .B(n11704), .Z(n11636) );
  AND U11574 ( .A(n270), .B(n11642), .Z(n11704) );
  XOR U11575 ( .A(n11703), .B(n11640), .Z(n11642) );
  XOR U11576 ( .A(n11705), .B(n11706), .Z(n11680) );
  AND U11577 ( .A(n11707), .B(n11708), .Z(n11706) );
  XNOR U11578 ( .A(n11705), .B(n11696), .Z(n11708) );
  IV U11579 ( .A(n11650), .Z(n11696) );
  XNOR U11580 ( .A(n11709), .B(n11689), .Z(n11650) );
  XNOR U11581 ( .A(n11710), .B(n11695), .Z(n11689) );
  XOR U11582 ( .A(n11711), .B(n11712), .Z(n11695) );
  NOR U11583 ( .A(n11713), .B(n11714), .Z(n11712) );
  XNOR U11584 ( .A(n11711), .B(n11715), .Z(n11713) );
  XNOR U11585 ( .A(n11694), .B(n11686), .Z(n11710) );
  XOR U11586 ( .A(n11716), .B(n11717), .Z(n11686) );
  AND U11587 ( .A(n11718), .B(n11719), .Z(n11717) );
  XNOR U11588 ( .A(n11716), .B(n11720), .Z(n11718) );
  XNOR U11589 ( .A(n11721), .B(n11691), .Z(n11694) );
  XOR U11590 ( .A(n11722), .B(n11723), .Z(n11691) );
  AND U11591 ( .A(n11724), .B(n11725), .Z(n11723) );
  XOR U11592 ( .A(n11722), .B(n11726), .Z(n11724) );
  XNOR U11593 ( .A(n11727), .B(n11728), .Z(n11721) );
  NOR U11594 ( .A(n11729), .B(n11730), .Z(n11728) );
  XOR U11595 ( .A(n11727), .B(n11731), .Z(n11729) );
  XNOR U11596 ( .A(n11690), .B(n11697), .Z(n11709) );
  NOR U11597 ( .A(n11658), .B(n11732), .Z(n11697) );
  XOR U11598 ( .A(n11702), .B(n11701), .Z(n11690) );
  XNOR U11599 ( .A(n11733), .B(n11698), .Z(n11701) );
  XOR U11600 ( .A(n11734), .B(n11735), .Z(n11698) );
  AND U11601 ( .A(n11736), .B(n11737), .Z(n11735) );
  XOR U11602 ( .A(n11734), .B(n11738), .Z(n11736) );
  XNOR U11603 ( .A(n11739), .B(n11740), .Z(n11733) );
  NOR U11604 ( .A(n11741), .B(n11742), .Z(n11740) );
  XNOR U11605 ( .A(n11739), .B(n11743), .Z(n11741) );
  XOR U11606 ( .A(n11744), .B(n11745), .Z(n11702) );
  NOR U11607 ( .A(n11746), .B(n11747), .Z(n11745) );
  XNOR U11608 ( .A(n11744), .B(n11748), .Z(n11746) );
  XNOR U11609 ( .A(n11647), .B(n11705), .Z(n11707) );
  XNOR U11610 ( .A(n11749), .B(n11750), .Z(n11647) );
  AND U11611 ( .A(n270), .B(n11654), .Z(n11750) );
  XOR U11612 ( .A(n11749), .B(n11652), .Z(n11654) );
  AND U11613 ( .A(n11655), .B(n11658), .Z(n11705) );
  XOR U11614 ( .A(n11751), .B(n11732), .Z(n11658) );
  XNOR U11615 ( .A(p_input[1024]), .B(p_input[336]), .Z(n11732) );
  XOR U11616 ( .A(n11720), .B(n11719), .Z(n11751) );
  XNOR U11617 ( .A(n11752), .B(n11726), .Z(n11719) );
  XNOR U11618 ( .A(n11715), .B(n11714), .Z(n11726) );
  XOR U11619 ( .A(n11753), .B(n11711), .Z(n11714) );
  XOR U11620 ( .A(p_input[1034]), .B(p_input[346]), .Z(n11711) );
  XNOR U11621 ( .A(p_input[1035]), .B(p_input[347]), .Z(n11753) );
  XOR U11622 ( .A(p_input[1036]), .B(p_input[348]), .Z(n11715) );
  XNOR U11623 ( .A(n11725), .B(n11716), .Z(n11752) );
  XOR U11624 ( .A(p_input[1025]), .B(p_input[337]), .Z(n11716) );
  XOR U11625 ( .A(n11754), .B(n11731), .Z(n11725) );
  XNOR U11626 ( .A(p_input[1039]), .B(p_input[351]), .Z(n11731) );
  XOR U11627 ( .A(n11722), .B(n11730), .Z(n11754) );
  XOR U11628 ( .A(n11755), .B(n11727), .Z(n11730) );
  XOR U11629 ( .A(p_input[1037]), .B(p_input[349]), .Z(n11727) );
  XNOR U11630 ( .A(p_input[1038]), .B(p_input[350]), .Z(n11755) );
  XOR U11631 ( .A(p_input[1033]), .B(p_input[345]), .Z(n11722) );
  XNOR U11632 ( .A(n11738), .B(n11737), .Z(n11720) );
  XNOR U11633 ( .A(n11756), .B(n11743), .Z(n11737) );
  XOR U11634 ( .A(p_input[1032]), .B(p_input[344]), .Z(n11743) );
  XOR U11635 ( .A(n11734), .B(n11742), .Z(n11756) );
  XOR U11636 ( .A(n11757), .B(n11739), .Z(n11742) );
  XOR U11637 ( .A(p_input[1030]), .B(p_input[342]), .Z(n11739) );
  XNOR U11638 ( .A(p_input[1031]), .B(p_input[343]), .Z(n11757) );
  XOR U11639 ( .A(p_input[1026]), .B(p_input[338]), .Z(n11734) );
  XNOR U11640 ( .A(n11748), .B(n11747), .Z(n11738) );
  XOR U11641 ( .A(n11758), .B(n11744), .Z(n11747) );
  XOR U11642 ( .A(p_input[1027]), .B(p_input[339]), .Z(n11744) );
  XNOR U11643 ( .A(p_input[1028]), .B(p_input[340]), .Z(n11758) );
  XOR U11644 ( .A(p_input[1029]), .B(p_input[341]), .Z(n11748) );
  XNOR U11645 ( .A(n11759), .B(n11760), .Z(n11655) );
  AND U11646 ( .A(n270), .B(n11761), .Z(n11760) );
  XNOR U11647 ( .A(n11762), .B(n11763), .Z(n270) );
  AND U11648 ( .A(n11764), .B(n11765), .Z(n11763) );
  XOR U11649 ( .A(n11762), .B(n11665), .Z(n11765) );
  XNOR U11650 ( .A(n11762), .B(n11619), .Z(n11764) );
  XOR U11651 ( .A(n11766), .B(n11767), .Z(n11762) );
  AND U11652 ( .A(n11768), .B(n11769), .Z(n11767) );
  XOR U11653 ( .A(n11766), .B(n11629), .Z(n11768) );
  XOR U11654 ( .A(n11770), .B(n11771), .Z(n11608) );
  AND U11655 ( .A(n274), .B(n11761), .Z(n11771) );
  XNOR U11656 ( .A(n11759), .B(n11770), .Z(n11761) );
  XNOR U11657 ( .A(n11772), .B(n11773), .Z(n274) );
  AND U11658 ( .A(n11774), .B(n11775), .Z(n11773) );
  XNOR U11659 ( .A(n11776), .B(n11772), .Z(n11775) );
  IV U11660 ( .A(n11665), .Z(n11776) );
  XNOR U11661 ( .A(n11777), .B(n11778), .Z(n11665) );
  AND U11662 ( .A(n277), .B(n11779), .Z(n11778) );
  XNOR U11663 ( .A(n11777), .B(n11780), .Z(n11779) );
  XNOR U11664 ( .A(n11619), .B(n11772), .Z(n11774) );
  XOR U11665 ( .A(n11781), .B(n11782), .Z(n11619) );
  AND U11666 ( .A(n285), .B(n11783), .Z(n11782) );
  XOR U11667 ( .A(n11766), .B(n11784), .Z(n11772) );
  AND U11668 ( .A(n11785), .B(n11769), .Z(n11784) );
  XNOR U11669 ( .A(n11678), .B(n11766), .Z(n11769) );
  XNOR U11670 ( .A(n11786), .B(n11787), .Z(n11678) );
  AND U11671 ( .A(n277), .B(n11788), .Z(n11787) );
  XOR U11672 ( .A(n11789), .B(n11786), .Z(n11788) );
  XNOR U11673 ( .A(n11790), .B(n11766), .Z(n11785) );
  IV U11674 ( .A(n11629), .Z(n11790) );
  XOR U11675 ( .A(n11791), .B(n11792), .Z(n11629) );
  AND U11676 ( .A(n285), .B(n11793), .Z(n11792) );
  XOR U11677 ( .A(n11794), .B(n11795), .Z(n11766) );
  AND U11678 ( .A(n11796), .B(n11797), .Z(n11795) );
  XNOR U11679 ( .A(n11703), .B(n11794), .Z(n11797) );
  XNOR U11680 ( .A(n11798), .B(n11799), .Z(n11703) );
  AND U11681 ( .A(n277), .B(n11800), .Z(n11799) );
  XNOR U11682 ( .A(n11801), .B(n11798), .Z(n11800) );
  XOR U11683 ( .A(n11794), .B(n11640), .Z(n11796) );
  XOR U11684 ( .A(n11802), .B(n11803), .Z(n11640) );
  AND U11685 ( .A(n285), .B(n11804), .Z(n11803) );
  XOR U11686 ( .A(n11805), .B(n11806), .Z(n11794) );
  AND U11687 ( .A(n11807), .B(n11808), .Z(n11806) );
  XNOR U11688 ( .A(n11805), .B(n11749), .Z(n11808) );
  XNOR U11689 ( .A(n11809), .B(n11810), .Z(n11749) );
  AND U11690 ( .A(n277), .B(n11811), .Z(n11810) );
  XOR U11691 ( .A(n11812), .B(n11809), .Z(n11811) );
  XNOR U11692 ( .A(n11813), .B(n11805), .Z(n11807) );
  IV U11693 ( .A(n11652), .Z(n11813) );
  XOR U11694 ( .A(n11814), .B(n11815), .Z(n11652) );
  AND U11695 ( .A(n285), .B(n11816), .Z(n11815) );
  AND U11696 ( .A(n11770), .B(n11759), .Z(n11805) );
  XNOR U11697 ( .A(n11817), .B(n11818), .Z(n11759) );
  AND U11698 ( .A(n277), .B(n11819), .Z(n11818) );
  XNOR U11699 ( .A(n11820), .B(n11817), .Z(n11819) );
  XNOR U11700 ( .A(n11821), .B(n11822), .Z(n277) );
  AND U11701 ( .A(n11823), .B(n11824), .Z(n11822) );
  XOR U11702 ( .A(n11780), .B(n11821), .Z(n11824) );
  AND U11703 ( .A(n11825), .B(n11826), .Z(n11780) );
  XOR U11704 ( .A(n11821), .B(n11777), .Z(n11823) );
  XNOR U11705 ( .A(n11827), .B(n11828), .Z(n11777) );
  AND U11706 ( .A(n281), .B(n11783), .Z(n11828) );
  XOR U11707 ( .A(n11781), .B(n11827), .Z(n11783) );
  XOR U11708 ( .A(n11829), .B(n11830), .Z(n11821) );
  AND U11709 ( .A(n11831), .B(n11832), .Z(n11830) );
  XNOR U11710 ( .A(n11829), .B(n11825), .Z(n11832) );
  IV U11711 ( .A(n11789), .Z(n11825) );
  XOR U11712 ( .A(n11833), .B(n11834), .Z(n11789) );
  XOR U11713 ( .A(n11835), .B(n11826), .Z(n11834) );
  AND U11714 ( .A(n11801), .B(n11836), .Z(n11826) );
  AND U11715 ( .A(n11837), .B(n11838), .Z(n11835) );
  XOR U11716 ( .A(n11839), .B(n11833), .Z(n11837) );
  XNOR U11717 ( .A(n11786), .B(n11829), .Z(n11831) );
  XNOR U11718 ( .A(n11840), .B(n11841), .Z(n11786) );
  AND U11719 ( .A(n281), .B(n11793), .Z(n11841) );
  XOR U11720 ( .A(n11840), .B(n11791), .Z(n11793) );
  XOR U11721 ( .A(n11842), .B(n11843), .Z(n11829) );
  AND U11722 ( .A(n11844), .B(n11845), .Z(n11843) );
  XNOR U11723 ( .A(n11842), .B(n11801), .Z(n11845) );
  XOR U11724 ( .A(n11846), .B(n11838), .Z(n11801) );
  XNOR U11725 ( .A(n11847), .B(n11833), .Z(n11838) );
  XOR U11726 ( .A(n11848), .B(n11849), .Z(n11833) );
  AND U11727 ( .A(n11850), .B(n11851), .Z(n11849) );
  XOR U11728 ( .A(n11852), .B(n11848), .Z(n11850) );
  XNOR U11729 ( .A(n11853), .B(n11854), .Z(n11847) );
  AND U11730 ( .A(n11855), .B(n11856), .Z(n11854) );
  XOR U11731 ( .A(n11853), .B(n11857), .Z(n11855) );
  XNOR U11732 ( .A(n11839), .B(n11836), .Z(n11846) );
  AND U11733 ( .A(n11858), .B(n11859), .Z(n11836) );
  XOR U11734 ( .A(n11860), .B(n11861), .Z(n11839) );
  AND U11735 ( .A(n11862), .B(n11863), .Z(n11861) );
  XOR U11736 ( .A(n11860), .B(n11864), .Z(n11862) );
  XNOR U11737 ( .A(n11798), .B(n11842), .Z(n11844) );
  XNOR U11738 ( .A(n11865), .B(n11866), .Z(n11798) );
  AND U11739 ( .A(n281), .B(n11804), .Z(n11866) );
  XOR U11740 ( .A(n11865), .B(n11802), .Z(n11804) );
  XOR U11741 ( .A(n11867), .B(n11868), .Z(n11842) );
  AND U11742 ( .A(n11869), .B(n11870), .Z(n11868) );
  XNOR U11743 ( .A(n11867), .B(n11858), .Z(n11870) );
  IV U11744 ( .A(n11812), .Z(n11858) );
  XNOR U11745 ( .A(n11871), .B(n11851), .Z(n11812) );
  XNOR U11746 ( .A(n11872), .B(n11857), .Z(n11851) );
  XOR U11747 ( .A(n11873), .B(n11874), .Z(n11857) );
  NOR U11748 ( .A(n11875), .B(n11876), .Z(n11874) );
  XNOR U11749 ( .A(n11873), .B(n11877), .Z(n11875) );
  XNOR U11750 ( .A(n11856), .B(n11848), .Z(n11872) );
  XOR U11751 ( .A(n11878), .B(n11879), .Z(n11848) );
  AND U11752 ( .A(n11880), .B(n11881), .Z(n11879) );
  XNOR U11753 ( .A(n11878), .B(n11882), .Z(n11880) );
  XNOR U11754 ( .A(n11883), .B(n11853), .Z(n11856) );
  XOR U11755 ( .A(n11884), .B(n11885), .Z(n11853) );
  AND U11756 ( .A(n11886), .B(n11887), .Z(n11885) );
  XOR U11757 ( .A(n11884), .B(n11888), .Z(n11886) );
  XNOR U11758 ( .A(n11889), .B(n11890), .Z(n11883) );
  NOR U11759 ( .A(n11891), .B(n11892), .Z(n11890) );
  XOR U11760 ( .A(n11889), .B(n11893), .Z(n11891) );
  XNOR U11761 ( .A(n11852), .B(n11859), .Z(n11871) );
  NOR U11762 ( .A(n11820), .B(n11894), .Z(n11859) );
  XOR U11763 ( .A(n11864), .B(n11863), .Z(n11852) );
  XNOR U11764 ( .A(n11895), .B(n11860), .Z(n11863) );
  XOR U11765 ( .A(n11896), .B(n11897), .Z(n11860) );
  AND U11766 ( .A(n11898), .B(n11899), .Z(n11897) );
  XOR U11767 ( .A(n11896), .B(n11900), .Z(n11898) );
  XNOR U11768 ( .A(n11901), .B(n11902), .Z(n11895) );
  NOR U11769 ( .A(n11903), .B(n11904), .Z(n11902) );
  XNOR U11770 ( .A(n11901), .B(n11905), .Z(n11903) );
  XOR U11771 ( .A(n11906), .B(n11907), .Z(n11864) );
  NOR U11772 ( .A(n11908), .B(n11909), .Z(n11907) );
  XNOR U11773 ( .A(n11906), .B(n11910), .Z(n11908) );
  XNOR U11774 ( .A(n11809), .B(n11867), .Z(n11869) );
  XNOR U11775 ( .A(n11911), .B(n11912), .Z(n11809) );
  AND U11776 ( .A(n281), .B(n11816), .Z(n11912) );
  XOR U11777 ( .A(n11911), .B(n11814), .Z(n11816) );
  AND U11778 ( .A(n11817), .B(n11820), .Z(n11867) );
  XOR U11779 ( .A(n11913), .B(n11894), .Z(n11820) );
  XNOR U11780 ( .A(p_input[1024]), .B(p_input[352]), .Z(n11894) );
  XOR U11781 ( .A(n11882), .B(n11881), .Z(n11913) );
  XNOR U11782 ( .A(n11914), .B(n11888), .Z(n11881) );
  XNOR U11783 ( .A(n11877), .B(n11876), .Z(n11888) );
  XOR U11784 ( .A(n11915), .B(n11873), .Z(n11876) );
  XOR U11785 ( .A(p_input[1034]), .B(p_input[362]), .Z(n11873) );
  XNOR U11786 ( .A(p_input[1035]), .B(p_input[363]), .Z(n11915) );
  XOR U11787 ( .A(p_input[1036]), .B(p_input[364]), .Z(n11877) );
  XNOR U11788 ( .A(n11887), .B(n11878), .Z(n11914) );
  XOR U11789 ( .A(p_input[1025]), .B(p_input[353]), .Z(n11878) );
  XOR U11790 ( .A(n11916), .B(n11893), .Z(n11887) );
  XNOR U11791 ( .A(p_input[1039]), .B(p_input[367]), .Z(n11893) );
  XOR U11792 ( .A(n11884), .B(n11892), .Z(n11916) );
  XOR U11793 ( .A(n11917), .B(n11889), .Z(n11892) );
  XOR U11794 ( .A(p_input[1037]), .B(p_input[365]), .Z(n11889) );
  XNOR U11795 ( .A(p_input[1038]), .B(p_input[366]), .Z(n11917) );
  XOR U11796 ( .A(p_input[1033]), .B(p_input[361]), .Z(n11884) );
  XNOR U11797 ( .A(n11900), .B(n11899), .Z(n11882) );
  XNOR U11798 ( .A(n11918), .B(n11905), .Z(n11899) );
  XOR U11799 ( .A(p_input[1032]), .B(p_input[360]), .Z(n11905) );
  XOR U11800 ( .A(n11896), .B(n11904), .Z(n11918) );
  XOR U11801 ( .A(n11919), .B(n11901), .Z(n11904) );
  XOR U11802 ( .A(p_input[1030]), .B(p_input[358]), .Z(n11901) );
  XNOR U11803 ( .A(p_input[1031]), .B(p_input[359]), .Z(n11919) );
  XOR U11804 ( .A(p_input[1026]), .B(p_input[354]), .Z(n11896) );
  XNOR U11805 ( .A(n11910), .B(n11909), .Z(n11900) );
  XOR U11806 ( .A(n11920), .B(n11906), .Z(n11909) );
  XOR U11807 ( .A(p_input[1027]), .B(p_input[355]), .Z(n11906) );
  XNOR U11808 ( .A(p_input[1028]), .B(p_input[356]), .Z(n11920) );
  XOR U11809 ( .A(p_input[1029]), .B(p_input[357]), .Z(n11910) );
  XNOR U11810 ( .A(n11921), .B(n11922), .Z(n11817) );
  AND U11811 ( .A(n281), .B(n11923), .Z(n11922) );
  XNOR U11812 ( .A(n11924), .B(n11925), .Z(n281) );
  AND U11813 ( .A(n11926), .B(n11927), .Z(n11925) );
  XOR U11814 ( .A(n11924), .B(n11827), .Z(n11927) );
  XNOR U11815 ( .A(n11924), .B(n11781), .Z(n11926) );
  XOR U11816 ( .A(n11928), .B(n11929), .Z(n11924) );
  AND U11817 ( .A(n11930), .B(n11931), .Z(n11929) );
  XOR U11818 ( .A(n11928), .B(n11791), .Z(n11930) );
  XOR U11819 ( .A(n11932), .B(n11933), .Z(n11770) );
  AND U11820 ( .A(n285), .B(n11923), .Z(n11933) );
  XNOR U11821 ( .A(n11921), .B(n11932), .Z(n11923) );
  XNOR U11822 ( .A(n11934), .B(n11935), .Z(n285) );
  AND U11823 ( .A(n11936), .B(n11937), .Z(n11935) );
  XNOR U11824 ( .A(n11938), .B(n11934), .Z(n11937) );
  IV U11825 ( .A(n11827), .Z(n11938) );
  XNOR U11826 ( .A(n11939), .B(n11940), .Z(n11827) );
  AND U11827 ( .A(n288), .B(n11941), .Z(n11940) );
  XNOR U11828 ( .A(n11939), .B(n11942), .Z(n11941) );
  XNOR U11829 ( .A(n11781), .B(n11934), .Z(n11936) );
  XOR U11830 ( .A(n11943), .B(n11944), .Z(n11781) );
  AND U11831 ( .A(n296), .B(n11945), .Z(n11944) );
  XOR U11832 ( .A(n11928), .B(n11946), .Z(n11934) );
  AND U11833 ( .A(n11947), .B(n11931), .Z(n11946) );
  XNOR U11834 ( .A(n11840), .B(n11928), .Z(n11931) );
  XNOR U11835 ( .A(n11948), .B(n11949), .Z(n11840) );
  AND U11836 ( .A(n288), .B(n11950), .Z(n11949) );
  XOR U11837 ( .A(n11951), .B(n11948), .Z(n11950) );
  XNOR U11838 ( .A(n11952), .B(n11928), .Z(n11947) );
  IV U11839 ( .A(n11791), .Z(n11952) );
  XOR U11840 ( .A(n11953), .B(n11954), .Z(n11791) );
  AND U11841 ( .A(n296), .B(n11955), .Z(n11954) );
  XOR U11842 ( .A(n11956), .B(n11957), .Z(n11928) );
  AND U11843 ( .A(n11958), .B(n11959), .Z(n11957) );
  XNOR U11844 ( .A(n11865), .B(n11956), .Z(n11959) );
  XNOR U11845 ( .A(n11960), .B(n11961), .Z(n11865) );
  AND U11846 ( .A(n288), .B(n11962), .Z(n11961) );
  XNOR U11847 ( .A(n11963), .B(n11960), .Z(n11962) );
  XOR U11848 ( .A(n11956), .B(n11802), .Z(n11958) );
  XOR U11849 ( .A(n11964), .B(n11965), .Z(n11802) );
  AND U11850 ( .A(n296), .B(n11966), .Z(n11965) );
  XOR U11851 ( .A(n11967), .B(n11968), .Z(n11956) );
  AND U11852 ( .A(n11969), .B(n11970), .Z(n11968) );
  XNOR U11853 ( .A(n11967), .B(n11911), .Z(n11970) );
  XNOR U11854 ( .A(n11971), .B(n11972), .Z(n11911) );
  AND U11855 ( .A(n288), .B(n11973), .Z(n11972) );
  XOR U11856 ( .A(n11974), .B(n11971), .Z(n11973) );
  XNOR U11857 ( .A(n11975), .B(n11967), .Z(n11969) );
  IV U11858 ( .A(n11814), .Z(n11975) );
  XOR U11859 ( .A(n11976), .B(n11977), .Z(n11814) );
  AND U11860 ( .A(n296), .B(n11978), .Z(n11977) );
  AND U11861 ( .A(n11932), .B(n11921), .Z(n11967) );
  XNOR U11862 ( .A(n11979), .B(n11980), .Z(n11921) );
  AND U11863 ( .A(n288), .B(n11981), .Z(n11980) );
  XNOR U11864 ( .A(n11982), .B(n11979), .Z(n11981) );
  XNOR U11865 ( .A(n11983), .B(n11984), .Z(n288) );
  AND U11866 ( .A(n11985), .B(n11986), .Z(n11984) );
  XOR U11867 ( .A(n11942), .B(n11983), .Z(n11986) );
  AND U11868 ( .A(n11987), .B(n11988), .Z(n11942) );
  XOR U11869 ( .A(n11983), .B(n11939), .Z(n11985) );
  XNOR U11870 ( .A(n11989), .B(n11990), .Z(n11939) );
  AND U11871 ( .A(n292), .B(n11945), .Z(n11990) );
  XOR U11872 ( .A(n11943), .B(n11989), .Z(n11945) );
  XOR U11873 ( .A(n11991), .B(n11992), .Z(n11983) );
  AND U11874 ( .A(n11993), .B(n11994), .Z(n11992) );
  XNOR U11875 ( .A(n11991), .B(n11987), .Z(n11994) );
  IV U11876 ( .A(n11951), .Z(n11987) );
  XOR U11877 ( .A(n11995), .B(n11996), .Z(n11951) );
  XOR U11878 ( .A(n11997), .B(n11988), .Z(n11996) );
  AND U11879 ( .A(n11963), .B(n11998), .Z(n11988) );
  AND U11880 ( .A(n11999), .B(n12000), .Z(n11997) );
  XOR U11881 ( .A(n12001), .B(n11995), .Z(n11999) );
  XNOR U11882 ( .A(n11948), .B(n11991), .Z(n11993) );
  XNOR U11883 ( .A(n12002), .B(n12003), .Z(n11948) );
  AND U11884 ( .A(n292), .B(n11955), .Z(n12003) );
  XOR U11885 ( .A(n12002), .B(n11953), .Z(n11955) );
  XOR U11886 ( .A(n12004), .B(n12005), .Z(n11991) );
  AND U11887 ( .A(n12006), .B(n12007), .Z(n12005) );
  XNOR U11888 ( .A(n12004), .B(n11963), .Z(n12007) );
  XOR U11889 ( .A(n12008), .B(n12000), .Z(n11963) );
  XNOR U11890 ( .A(n12009), .B(n11995), .Z(n12000) );
  XOR U11891 ( .A(n12010), .B(n12011), .Z(n11995) );
  AND U11892 ( .A(n12012), .B(n12013), .Z(n12011) );
  XOR U11893 ( .A(n12014), .B(n12010), .Z(n12012) );
  XNOR U11894 ( .A(n12015), .B(n12016), .Z(n12009) );
  AND U11895 ( .A(n12017), .B(n12018), .Z(n12016) );
  XOR U11896 ( .A(n12015), .B(n12019), .Z(n12017) );
  XNOR U11897 ( .A(n12001), .B(n11998), .Z(n12008) );
  AND U11898 ( .A(n12020), .B(n12021), .Z(n11998) );
  XOR U11899 ( .A(n12022), .B(n12023), .Z(n12001) );
  AND U11900 ( .A(n12024), .B(n12025), .Z(n12023) );
  XOR U11901 ( .A(n12022), .B(n12026), .Z(n12024) );
  XNOR U11902 ( .A(n11960), .B(n12004), .Z(n12006) );
  XNOR U11903 ( .A(n12027), .B(n12028), .Z(n11960) );
  AND U11904 ( .A(n292), .B(n11966), .Z(n12028) );
  XOR U11905 ( .A(n12027), .B(n11964), .Z(n11966) );
  XOR U11906 ( .A(n12029), .B(n12030), .Z(n12004) );
  AND U11907 ( .A(n12031), .B(n12032), .Z(n12030) );
  XNOR U11908 ( .A(n12029), .B(n12020), .Z(n12032) );
  IV U11909 ( .A(n11974), .Z(n12020) );
  XNOR U11910 ( .A(n12033), .B(n12013), .Z(n11974) );
  XNOR U11911 ( .A(n12034), .B(n12019), .Z(n12013) );
  XOR U11912 ( .A(n12035), .B(n12036), .Z(n12019) );
  NOR U11913 ( .A(n12037), .B(n12038), .Z(n12036) );
  XNOR U11914 ( .A(n12035), .B(n12039), .Z(n12037) );
  XNOR U11915 ( .A(n12018), .B(n12010), .Z(n12034) );
  XOR U11916 ( .A(n12040), .B(n12041), .Z(n12010) );
  AND U11917 ( .A(n12042), .B(n12043), .Z(n12041) );
  XNOR U11918 ( .A(n12040), .B(n12044), .Z(n12042) );
  XNOR U11919 ( .A(n12045), .B(n12015), .Z(n12018) );
  XOR U11920 ( .A(n12046), .B(n12047), .Z(n12015) );
  AND U11921 ( .A(n12048), .B(n12049), .Z(n12047) );
  XOR U11922 ( .A(n12046), .B(n12050), .Z(n12048) );
  XNOR U11923 ( .A(n12051), .B(n12052), .Z(n12045) );
  NOR U11924 ( .A(n12053), .B(n12054), .Z(n12052) );
  XOR U11925 ( .A(n12051), .B(n12055), .Z(n12053) );
  XNOR U11926 ( .A(n12014), .B(n12021), .Z(n12033) );
  NOR U11927 ( .A(n11982), .B(n12056), .Z(n12021) );
  XOR U11928 ( .A(n12026), .B(n12025), .Z(n12014) );
  XNOR U11929 ( .A(n12057), .B(n12022), .Z(n12025) );
  XOR U11930 ( .A(n12058), .B(n12059), .Z(n12022) );
  AND U11931 ( .A(n12060), .B(n12061), .Z(n12059) );
  XOR U11932 ( .A(n12058), .B(n12062), .Z(n12060) );
  XNOR U11933 ( .A(n12063), .B(n12064), .Z(n12057) );
  NOR U11934 ( .A(n12065), .B(n12066), .Z(n12064) );
  XNOR U11935 ( .A(n12063), .B(n12067), .Z(n12065) );
  XOR U11936 ( .A(n12068), .B(n12069), .Z(n12026) );
  NOR U11937 ( .A(n12070), .B(n12071), .Z(n12069) );
  XNOR U11938 ( .A(n12068), .B(n12072), .Z(n12070) );
  XNOR U11939 ( .A(n11971), .B(n12029), .Z(n12031) );
  XNOR U11940 ( .A(n12073), .B(n12074), .Z(n11971) );
  AND U11941 ( .A(n292), .B(n11978), .Z(n12074) );
  XOR U11942 ( .A(n12073), .B(n11976), .Z(n11978) );
  AND U11943 ( .A(n11979), .B(n11982), .Z(n12029) );
  XOR U11944 ( .A(n12075), .B(n12056), .Z(n11982) );
  XNOR U11945 ( .A(p_input[1024]), .B(p_input[368]), .Z(n12056) );
  XOR U11946 ( .A(n12044), .B(n12043), .Z(n12075) );
  XNOR U11947 ( .A(n12076), .B(n12050), .Z(n12043) );
  XNOR U11948 ( .A(n12039), .B(n12038), .Z(n12050) );
  XOR U11949 ( .A(n12077), .B(n12035), .Z(n12038) );
  XOR U11950 ( .A(p_input[1034]), .B(p_input[378]), .Z(n12035) );
  XNOR U11951 ( .A(p_input[1035]), .B(p_input[379]), .Z(n12077) );
  XOR U11952 ( .A(p_input[1036]), .B(p_input[380]), .Z(n12039) );
  XNOR U11953 ( .A(n12049), .B(n12040), .Z(n12076) );
  XOR U11954 ( .A(p_input[1025]), .B(p_input[369]), .Z(n12040) );
  XOR U11955 ( .A(n12078), .B(n12055), .Z(n12049) );
  XNOR U11956 ( .A(p_input[1039]), .B(p_input[383]), .Z(n12055) );
  XOR U11957 ( .A(n12046), .B(n12054), .Z(n12078) );
  XOR U11958 ( .A(n12079), .B(n12051), .Z(n12054) );
  XOR U11959 ( .A(p_input[1037]), .B(p_input[381]), .Z(n12051) );
  XNOR U11960 ( .A(p_input[1038]), .B(p_input[382]), .Z(n12079) );
  XOR U11961 ( .A(p_input[1033]), .B(p_input[377]), .Z(n12046) );
  XNOR U11962 ( .A(n12062), .B(n12061), .Z(n12044) );
  XNOR U11963 ( .A(n12080), .B(n12067), .Z(n12061) );
  XOR U11964 ( .A(p_input[1032]), .B(p_input[376]), .Z(n12067) );
  XOR U11965 ( .A(n12058), .B(n12066), .Z(n12080) );
  XOR U11966 ( .A(n12081), .B(n12063), .Z(n12066) );
  XOR U11967 ( .A(p_input[1030]), .B(p_input[374]), .Z(n12063) );
  XNOR U11968 ( .A(p_input[1031]), .B(p_input[375]), .Z(n12081) );
  XOR U11969 ( .A(p_input[1026]), .B(p_input[370]), .Z(n12058) );
  XNOR U11970 ( .A(n12072), .B(n12071), .Z(n12062) );
  XOR U11971 ( .A(n12082), .B(n12068), .Z(n12071) );
  XOR U11972 ( .A(p_input[1027]), .B(p_input[371]), .Z(n12068) );
  XNOR U11973 ( .A(p_input[1028]), .B(p_input[372]), .Z(n12082) );
  XOR U11974 ( .A(p_input[1029]), .B(p_input[373]), .Z(n12072) );
  XNOR U11975 ( .A(n12083), .B(n12084), .Z(n11979) );
  AND U11976 ( .A(n292), .B(n12085), .Z(n12084) );
  XNOR U11977 ( .A(n12086), .B(n12087), .Z(n292) );
  AND U11978 ( .A(n12088), .B(n12089), .Z(n12087) );
  XOR U11979 ( .A(n12086), .B(n11989), .Z(n12089) );
  XNOR U11980 ( .A(n12086), .B(n11943), .Z(n12088) );
  XOR U11981 ( .A(n12090), .B(n12091), .Z(n12086) );
  AND U11982 ( .A(n12092), .B(n12093), .Z(n12091) );
  XOR U11983 ( .A(n12090), .B(n11953), .Z(n12092) );
  XOR U11984 ( .A(n12094), .B(n12095), .Z(n11932) );
  AND U11985 ( .A(n296), .B(n12085), .Z(n12095) );
  XNOR U11986 ( .A(n12083), .B(n12094), .Z(n12085) );
  XNOR U11987 ( .A(n12096), .B(n12097), .Z(n296) );
  AND U11988 ( .A(n12098), .B(n12099), .Z(n12097) );
  XNOR U11989 ( .A(n12100), .B(n12096), .Z(n12099) );
  IV U11990 ( .A(n11989), .Z(n12100) );
  XNOR U11991 ( .A(n12101), .B(n12102), .Z(n11989) );
  AND U11992 ( .A(n299), .B(n12103), .Z(n12102) );
  XNOR U11993 ( .A(n12101), .B(n12104), .Z(n12103) );
  XNOR U11994 ( .A(n11943), .B(n12096), .Z(n12098) );
  XOR U11995 ( .A(n12105), .B(n12106), .Z(n11943) );
  AND U11996 ( .A(n307), .B(n12107), .Z(n12106) );
  XOR U11997 ( .A(n12090), .B(n12108), .Z(n12096) );
  AND U11998 ( .A(n12109), .B(n12093), .Z(n12108) );
  XNOR U11999 ( .A(n12002), .B(n12090), .Z(n12093) );
  XNOR U12000 ( .A(n12110), .B(n12111), .Z(n12002) );
  AND U12001 ( .A(n299), .B(n12112), .Z(n12111) );
  XOR U12002 ( .A(n12113), .B(n12110), .Z(n12112) );
  XNOR U12003 ( .A(n12114), .B(n12090), .Z(n12109) );
  IV U12004 ( .A(n11953), .Z(n12114) );
  XOR U12005 ( .A(n12115), .B(n12116), .Z(n11953) );
  AND U12006 ( .A(n307), .B(n12117), .Z(n12116) );
  XOR U12007 ( .A(n12118), .B(n12119), .Z(n12090) );
  AND U12008 ( .A(n12120), .B(n12121), .Z(n12119) );
  XNOR U12009 ( .A(n12027), .B(n12118), .Z(n12121) );
  XNOR U12010 ( .A(n12122), .B(n12123), .Z(n12027) );
  AND U12011 ( .A(n299), .B(n12124), .Z(n12123) );
  XNOR U12012 ( .A(n12125), .B(n12122), .Z(n12124) );
  XOR U12013 ( .A(n12118), .B(n11964), .Z(n12120) );
  XOR U12014 ( .A(n12126), .B(n12127), .Z(n11964) );
  AND U12015 ( .A(n307), .B(n12128), .Z(n12127) );
  XOR U12016 ( .A(n12129), .B(n12130), .Z(n12118) );
  AND U12017 ( .A(n12131), .B(n12132), .Z(n12130) );
  XNOR U12018 ( .A(n12129), .B(n12073), .Z(n12132) );
  XNOR U12019 ( .A(n12133), .B(n12134), .Z(n12073) );
  AND U12020 ( .A(n299), .B(n12135), .Z(n12134) );
  XOR U12021 ( .A(n12136), .B(n12133), .Z(n12135) );
  XNOR U12022 ( .A(n12137), .B(n12129), .Z(n12131) );
  IV U12023 ( .A(n11976), .Z(n12137) );
  XOR U12024 ( .A(n12138), .B(n12139), .Z(n11976) );
  AND U12025 ( .A(n307), .B(n12140), .Z(n12139) );
  AND U12026 ( .A(n12094), .B(n12083), .Z(n12129) );
  XNOR U12027 ( .A(n12141), .B(n12142), .Z(n12083) );
  AND U12028 ( .A(n299), .B(n12143), .Z(n12142) );
  XNOR U12029 ( .A(n12144), .B(n12141), .Z(n12143) );
  XNOR U12030 ( .A(n12145), .B(n12146), .Z(n299) );
  AND U12031 ( .A(n12147), .B(n12148), .Z(n12146) );
  XOR U12032 ( .A(n12104), .B(n12145), .Z(n12148) );
  AND U12033 ( .A(n12149), .B(n12150), .Z(n12104) );
  XOR U12034 ( .A(n12145), .B(n12101), .Z(n12147) );
  XNOR U12035 ( .A(n12151), .B(n12152), .Z(n12101) );
  AND U12036 ( .A(n303), .B(n12107), .Z(n12152) );
  XOR U12037 ( .A(n12105), .B(n12151), .Z(n12107) );
  XOR U12038 ( .A(n12153), .B(n12154), .Z(n12145) );
  AND U12039 ( .A(n12155), .B(n12156), .Z(n12154) );
  XNOR U12040 ( .A(n12153), .B(n12149), .Z(n12156) );
  IV U12041 ( .A(n12113), .Z(n12149) );
  XOR U12042 ( .A(n12157), .B(n12158), .Z(n12113) );
  XOR U12043 ( .A(n12159), .B(n12150), .Z(n12158) );
  AND U12044 ( .A(n12125), .B(n12160), .Z(n12150) );
  AND U12045 ( .A(n12161), .B(n12162), .Z(n12159) );
  XOR U12046 ( .A(n12163), .B(n12157), .Z(n12161) );
  XNOR U12047 ( .A(n12110), .B(n12153), .Z(n12155) );
  XNOR U12048 ( .A(n12164), .B(n12165), .Z(n12110) );
  AND U12049 ( .A(n303), .B(n12117), .Z(n12165) );
  XOR U12050 ( .A(n12164), .B(n12115), .Z(n12117) );
  XOR U12051 ( .A(n12166), .B(n12167), .Z(n12153) );
  AND U12052 ( .A(n12168), .B(n12169), .Z(n12167) );
  XNOR U12053 ( .A(n12166), .B(n12125), .Z(n12169) );
  XOR U12054 ( .A(n12170), .B(n12162), .Z(n12125) );
  XNOR U12055 ( .A(n12171), .B(n12157), .Z(n12162) );
  XOR U12056 ( .A(n12172), .B(n12173), .Z(n12157) );
  AND U12057 ( .A(n12174), .B(n12175), .Z(n12173) );
  XOR U12058 ( .A(n12176), .B(n12172), .Z(n12174) );
  XNOR U12059 ( .A(n12177), .B(n12178), .Z(n12171) );
  AND U12060 ( .A(n12179), .B(n12180), .Z(n12178) );
  XOR U12061 ( .A(n12177), .B(n12181), .Z(n12179) );
  XNOR U12062 ( .A(n12163), .B(n12160), .Z(n12170) );
  AND U12063 ( .A(n12182), .B(n12183), .Z(n12160) );
  XOR U12064 ( .A(n12184), .B(n12185), .Z(n12163) );
  AND U12065 ( .A(n12186), .B(n12187), .Z(n12185) );
  XOR U12066 ( .A(n12184), .B(n12188), .Z(n12186) );
  XNOR U12067 ( .A(n12122), .B(n12166), .Z(n12168) );
  XNOR U12068 ( .A(n12189), .B(n12190), .Z(n12122) );
  AND U12069 ( .A(n303), .B(n12128), .Z(n12190) );
  XOR U12070 ( .A(n12189), .B(n12126), .Z(n12128) );
  XOR U12071 ( .A(n12191), .B(n12192), .Z(n12166) );
  AND U12072 ( .A(n12193), .B(n12194), .Z(n12192) );
  XNOR U12073 ( .A(n12191), .B(n12182), .Z(n12194) );
  IV U12074 ( .A(n12136), .Z(n12182) );
  XNOR U12075 ( .A(n12195), .B(n12175), .Z(n12136) );
  XNOR U12076 ( .A(n12196), .B(n12181), .Z(n12175) );
  XOR U12077 ( .A(n12197), .B(n12198), .Z(n12181) );
  NOR U12078 ( .A(n12199), .B(n12200), .Z(n12198) );
  XNOR U12079 ( .A(n12197), .B(n12201), .Z(n12199) );
  XNOR U12080 ( .A(n12180), .B(n12172), .Z(n12196) );
  XOR U12081 ( .A(n12202), .B(n12203), .Z(n12172) );
  AND U12082 ( .A(n12204), .B(n12205), .Z(n12203) );
  XNOR U12083 ( .A(n12202), .B(n12206), .Z(n12204) );
  XNOR U12084 ( .A(n12207), .B(n12177), .Z(n12180) );
  XOR U12085 ( .A(n12208), .B(n12209), .Z(n12177) );
  AND U12086 ( .A(n12210), .B(n12211), .Z(n12209) );
  XOR U12087 ( .A(n12208), .B(n12212), .Z(n12210) );
  XNOR U12088 ( .A(n12213), .B(n12214), .Z(n12207) );
  NOR U12089 ( .A(n12215), .B(n12216), .Z(n12214) );
  XOR U12090 ( .A(n12213), .B(n12217), .Z(n12215) );
  XNOR U12091 ( .A(n12176), .B(n12183), .Z(n12195) );
  NOR U12092 ( .A(n12144), .B(n12218), .Z(n12183) );
  XOR U12093 ( .A(n12188), .B(n12187), .Z(n12176) );
  XNOR U12094 ( .A(n12219), .B(n12184), .Z(n12187) );
  XOR U12095 ( .A(n12220), .B(n12221), .Z(n12184) );
  AND U12096 ( .A(n12222), .B(n12223), .Z(n12221) );
  XOR U12097 ( .A(n12220), .B(n12224), .Z(n12222) );
  XNOR U12098 ( .A(n12225), .B(n12226), .Z(n12219) );
  NOR U12099 ( .A(n12227), .B(n12228), .Z(n12226) );
  XNOR U12100 ( .A(n12225), .B(n12229), .Z(n12227) );
  XOR U12101 ( .A(n12230), .B(n12231), .Z(n12188) );
  NOR U12102 ( .A(n12232), .B(n12233), .Z(n12231) );
  XNOR U12103 ( .A(n12230), .B(n12234), .Z(n12232) );
  XNOR U12104 ( .A(n12133), .B(n12191), .Z(n12193) );
  XNOR U12105 ( .A(n12235), .B(n12236), .Z(n12133) );
  AND U12106 ( .A(n303), .B(n12140), .Z(n12236) );
  XOR U12107 ( .A(n12235), .B(n12138), .Z(n12140) );
  AND U12108 ( .A(n12141), .B(n12144), .Z(n12191) );
  XOR U12109 ( .A(n12237), .B(n12218), .Z(n12144) );
  XNOR U12110 ( .A(p_input[1024]), .B(p_input[384]), .Z(n12218) );
  XOR U12111 ( .A(n12206), .B(n12205), .Z(n12237) );
  XNOR U12112 ( .A(n12238), .B(n12212), .Z(n12205) );
  XNOR U12113 ( .A(n12201), .B(n12200), .Z(n12212) );
  XOR U12114 ( .A(n12239), .B(n12197), .Z(n12200) );
  XOR U12115 ( .A(p_input[1034]), .B(p_input[394]), .Z(n12197) );
  XNOR U12116 ( .A(p_input[1035]), .B(p_input[395]), .Z(n12239) );
  XOR U12117 ( .A(p_input[1036]), .B(p_input[396]), .Z(n12201) );
  XNOR U12118 ( .A(n12211), .B(n12202), .Z(n12238) );
  XOR U12119 ( .A(p_input[1025]), .B(p_input[385]), .Z(n12202) );
  XOR U12120 ( .A(n12240), .B(n12217), .Z(n12211) );
  XNOR U12121 ( .A(p_input[1039]), .B(p_input[399]), .Z(n12217) );
  XOR U12122 ( .A(n12208), .B(n12216), .Z(n12240) );
  XOR U12123 ( .A(n12241), .B(n12213), .Z(n12216) );
  XOR U12124 ( .A(p_input[1037]), .B(p_input[397]), .Z(n12213) );
  XNOR U12125 ( .A(p_input[1038]), .B(p_input[398]), .Z(n12241) );
  XOR U12126 ( .A(p_input[1033]), .B(p_input[393]), .Z(n12208) );
  XNOR U12127 ( .A(n12224), .B(n12223), .Z(n12206) );
  XNOR U12128 ( .A(n12242), .B(n12229), .Z(n12223) );
  XOR U12129 ( .A(p_input[1032]), .B(p_input[392]), .Z(n12229) );
  XOR U12130 ( .A(n12220), .B(n12228), .Z(n12242) );
  XOR U12131 ( .A(n12243), .B(n12225), .Z(n12228) );
  XOR U12132 ( .A(p_input[1030]), .B(p_input[390]), .Z(n12225) );
  XNOR U12133 ( .A(p_input[1031]), .B(p_input[391]), .Z(n12243) );
  XOR U12134 ( .A(p_input[1026]), .B(p_input[386]), .Z(n12220) );
  XNOR U12135 ( .A(n12234), .B(n12233), .Z(n12224) );
  XOR U12136 ( .A(n12244), .B(n12230), .Z(n12233) );
  XOR U12137 ( .A(p_input[1027]), .B(p_input[387]), .Z(n12230) );
  XNOR U12138 ( .A(p_input[1028]), .B(p_input[388]), .Z(n12244) );
  XOR U12139 ( .A(p_input[1029]), .B(p_input[389]), .Z(n12234) );
  XNOR U12140 ( .A(n12245), .B(n12246), .Z(n12141) );
  AND U12141 ( .A(n303), .B(n12247), .Z(n12246) );
  XNOR U12142 ( .A(n12248), .B(n12249), .Z(n303) );
  AND U12143 ( .A(n12250), .B(n12251), .Z(n12249) );
  XOR U12144 ( .A(n12248), .B(n12151), .Z(n12251) );
  XNOR U12145 ( .A(n12248), .B(n12105), .Z(n12250) );
  XOR U12146 ( .A(n12252), .B(n12253), .Z(n12248) );
  AND U12147 ( .A(n12254), .B(n12255), .Z(n12253) );
  XOR U12148 ( .A(n12252), .B(n12115), .Z(n12254) );
  XOR U12149 ( .A(n12256), .B(n12257), .Z(n12094) );
  AND U12150 ( .A(n307), .B(n12247), .Z(n12257) );
  XNOR U12151 ( .A(n12245), .B(n12256), .Z(n12247) );
  XNOR U12152 ( .A(n12258), .B(n12259), .Z(n307) );
  AND U12153 ( .A(n12260), .B(n12261), .Z(n12259) );
  XNOR U12154 ( .A(n12262), .B(n12258), .Z(n12261) );
  IV U12155 ( .A(n12151), .Z(n12262) );
  XNOR U12156 ( .A(n12263), .B(n12264), .Z(n12151) );
  AND U12157 ( .A(n310), .B(n12265), .Z(n12264) );
  XNOR U12158 ( .A(n12263), .B(n12266), .Z(n12265) );
  XNOR U12159 ( .A(n12105), .B(n12258), .Z(n12260) );
  XOR U12160 ( .A(n12267), .B(n12268), .Z(n12105) );
  AND U12161 ( .A(n318), .B(n12269), .Z(n12268) );
  XOR U12162 ( .A(n12252), .B(n12270), .Z(n12258) );
  AND U12163 ( .A(n12271), .B(n12255), .Z(n12270) );
  XNOR U12164 ( .A(n12164), .B(n12252), .Z(n12255) );
  XNOR U12165 ( .A(n12272), .B(n12273), .Z(n12164) );
  AND U12166 ( .A(n310), .B(n12274), .Z(n12273) );
  XOR U12167 ( .A(n12275), .B(n12272), .Z(n12274) );
  XNOR U12168 ( .A(n12276), .B(n12252), .Z(n12271) );
  IV U12169 ( .A(n12115), .Z(n12276) );
  XOR U12170 ( .A(n12277), .B(n12278), .Z(n12115) );
  AND U12171 ( .A(n318), .B(n12279), .Z(n12278) );
  XOR U12172 ( .A(n12280), .B(n12281), .Z(n12252) );
  AND U12173 ( .A(n12282), .B(n12283), .Z(n12281) );
  XNOR U12174 ( .A(n12189), .B(n12280), .Z(n12283) );
  XNOR U12175 ( .A(n12284), .B(n12285), .Z(n12189) );
  AND U12176 ( .A(n310), .B(n12286), .Z(n12285) );
  XNOR U12177 ( .A(n12287), .B(n12284), .Z(n12286) );
  XOR U12178 ( .A(n12280), .B(n12126), .Z(n12282) );
  XOR U12179 ( .A(n12288), .B(n12289), .Z(n12126) );
  AND U12180 ( .A(n318), .B(n12290), .Z(n12289) );
  XOR U12181 ( .A(n12291), .B(n12292), .Z(n12280) );
  AND U12182 ( .A(n12293), .B(n12294), .Z(n12292) );
  XNOR U12183 ( .A(n12291), .B(n12235), .Z(n12294) );
  XNOR U12184 ( .A(n12295), .B(n12296), .Z(n12235) );
  AND U12185 ( .A(n310), .B(n12297), .Z(n12296) );
  XOR U12186 ( .A(n12298), .B(n12295), .Z(n12297) );
  XNOR U12187 ( .A(n12299), .B(n12291), .Z(n12293) );
  IV U12188 ( .A(n12138), .Z(n12299) );
  XOR U12189 ( .A(n12300), .B(n12301), .Z(n12138) );
  AND U12190 ( .A(n318), .B(n12302), .Z(n12301) );
  AND U12191 ( .A(n12256), .B(n12245), .Z(n12291) );
  XNOR U12192 ( .A(n12303), .B(n12304), .Z(n12245) );
  AND U12193 ( .A(n310), .B(n12305), .Z(n12304) );
  XNOR U12194 ( .A(n12306), .B(n12303), .Z(n12305) );
  XNOR U12195 ( .A(n12307), .B(n12308), .Z(n310) );
  AND U12196 ( .A(n12309), .B(n12310), .Z(n12308) );
  XOR U12197 ( .A(n12266), .B(n12307), .Z(n12310) );
  AND U12198 ( .A(n12311), .B(n12312), .Z(n12266) );
  XOR U12199 ( .A(n12307), .B(n12263), .Z(n12309) );
  XNOR U12200 ( .A(n12313), .B(n12314), .Z(n12263) );
  AND U12201 ( .A(n314), .B(n12269), .Z(n12314) );
  XOR U12202 ( .A(n12267), .B(n12313), .Z(n12269) );
  XOR U12203 ( .A(n12315), .B(n12316), .Z(n12307) );
  AND U12204 ( .A(n12317), .B(n12318), .Z(n12316) );
  XNOR U12205 ( .A(n12315), .B(n12311), .Z(n12318) );
  IV U12206 ( .A(n12275), .Z(n12311) );
  XOR U12207 ( .A(n12319), .B(n12320), .Z(n12275) );
  XOR U12208 ( .A(n12321), .B(n12312), .Z(n12320) );
  AND U12209 ( .A(n12287), .B(n12322), .Z(n12312) );
  AND U12210 ( .A(n12323), .B(n12324), .Z(n12321) );
  XOR U12211 ( .A(n12325), .B(n12319), .Z(n12323) );
  XNOR U12212 ( .A(n12272), .B(n12315), .Z(n12317) );
  XNOR U12213 ( .A(n12326), .B(n12327), .Z(n12272) );
  AND U12214 ( .A(n314), .B(n12279), .Z(n12327) );
  XOR U12215 ( .A(n12326), .B(n12277), .Z(n12279) );
  XOR U12216 ( .A(n12328), .B(n12329), .Z(n12315) );
  AND U12217 ( .A(n12330), .B(n12331), .Z(n12329) );
  XNOR U12218 ( .A(n12328), .B(n12287), .Z(n12331) );
  XOR U12219 ( .A(n12332), .B(n12324), .Z(n12287) );
  XNOR U12220 ( .A(n12333), .B(n12319), .Z(n12324) );
  XOR U12221 ( .A(n12334), .B(n12335), .Z(n12319) );
  AND U12222 ( .A(n12336), .B(n12337), .Z(n12335) );
  XOR U12223 ( .A(n12338), .B(n12334), .Z(n12336) );
  XNOR U12224 ( .A(n12339), .B(n12340), .Z(n12333) );
  AND U12225 ( .A(n12341), .B(n12342), .Z(n12340) );
  XOR U12226 ( .A(n12339), .B(n12343), .Z(n12341) );
  XNOR U12227 ( .A(n12325), .B(n12322), .Z(n12332) );
  AND U12228 ( .A(n12344), .B(n12345), .Z(n12322) );
  XOR U12229 ( .A(n12346), .B(n12347), .Z(n12325) );
  AND U12230 ( .A(n12348), .B(n12349), .Z(n12347) );
  XOR U12231 ( .A(n12346), .B(n12350), .Z(n12348) );
  XNOR U12232 ( .A(n12284), .B(n12328), .Z(n12330) );
  XNOR U12233 ( .A(n12351), .B(n12352), .Z(n12284) );
  AND U12234 ( .A(n314), .B(n12290), .Z(n12352) );
  XOR U12235 ( .A(n12351), .B(n12288), .Z(n12290) );
  XOR U12236 ( .A(n12353), .B(n12354), .Z(n12328) );
  AND U12237 ( .A(n12355), .B(n12356), .Z(n12354) );
  XNOR U12238 ( .A(n12353), .B(n12344), .Z(n12356) );
  IV U12239 ( .A(n12298), .Z(n12344) );
  XNOR U12240 ( .A(n12357), .B(n12337), .Z(n12298) );
  XNOR U12241 ( .A(n12358), .B(n12343), .Z(n12337) );
  XOR U12242 ( .A(n12359), .B(n12360), .Z(n12343) );
  NOR U12243 ( .A(n12361), .B(n12362), .Z(n12360) );
  XNOR U12244 ( .A(n12359), .B(n12363), .Z(n12361) );
  XNOR U12245 ( .A(n12342), .B(n12334), .Z(n12358) );
  XOR U12246 ( .A(n12364), .B(n12365), .Z(n12334) );
  AND U12247 ( .A(n12366), .B(n12367), .Z(n12365) );
  XNOR U12248 ( .A(n12364), .B(n12368), .Z(n12366) );
  XNOR U12249 ( .A(n12369), .B(n12339), .Z(n12342) );
  XOR U12250 ( .A(n12370), .B(n12371), .Z(n12339) );
  AND U12251 ( .A(n12372), .B(n12373), .Z(n12371) );
  XOR U12252 ( .A(n12370), .B(n12374), .Z(n12372) );
  XNOR U12253 ( .A(n12375), .B(n12376), .Z(n12369) );
  NOR U12254 ( .A(n12377), .B(n12378), .Z(n12376) );
  XOR U12255 ( .A(n12375), .B(n12379), .Z(n12377) );
  XNOR U12256 ( .A(n12338), .B(n12345), .Z(n12357) );
  NOR U12257 ( .A(n12306), .B(n12380), .Z(n12345) );
  XOR U12258 ( .A(n12350), .B(n12349), .Z(n12338) );
  XNOR U12259 ( .A(n12381), .B(n12346), .Z(n12349) );
  XOR U12260 ( .A(n12382), .B(n12383), .Z(n12346) );
  AND U12261 ( .A(n12384), .B(n12385), .Z(n12383) );
  XOR U12262 ( .A(n12382), .B(n12386), .Z(n12384) );
  XNOR U12263 ( .A(n12387), .B(n12388), .Z(n12381) );
  NOR U12264 ( .A(n12389), .B(n12390), .Z(n12388) );
  XNOR U12265 ( .A(n12387), .B(n12391), .Z(n12389) );
  XOR U12266 ( .A(n12392), .B(n12393), .Z(n12350) );
  NOR U12267 ( .A(n12394), .B(n12395), .Z(n12393) );
  XNOR U12268 ( .A(n12392), .B(n12396), .Z(n12394) );
  XNOR U12269 ( .A(n12295), .B(n12353), .Z(n12355) );
  XNOR U12270 ( .A(n12397), .B(n12398), .Z(n12295) );
  AND U12271 ( .A(n314), .B(n12302), .Z(n12398) );
  XOR U12272 ( .A(n12397), .B(n12300), .Z(n12302) );
  AND U12273 ( .A(n12303), .B(n12306), .Z(n12353) );
  XOR U12274 ( .A(n12399), .B(n12380), .Z(n12306) );
  XNOR U12275 ( .A(p_input[1024]), .B(p_input[400]), .Z(n12380) );
  XOR U12276 ( .A(n12368), .B(n12367), .Z(n12399) );
  XNOR U12277 ( .A(n12400), .B(n12374), .Z(n12367) );
  XNOR U12278 ( .A(n12363), .B(n12362), .Z(n12374) );
  XOR U12279 ( .A(n12401), .B(n12359), .Z(n12362) );
  XOR U12280 ( .A(p_input[1034]), .B(p_input[410]), .Z(n12359) );
  XNOR U12281 ( .A(p_input[1035]), .B(p_input[411]), .Z(n12401) );
  XOR U12282 ( .A(p_input[1036]), .B(p_input[412]), .Z(n12363) );
  XNOR U12283 ( .A(n12373), .B(n12364), .Z(n12400) );
  XOR U12284 ( .A(p_input[1025]), .B(p_input[401]), .Z(n12364) );
  XOR U12285 ( .A(n12402), .B(n12379), .Z(n12373) );
  XNOR U12286 ( .A(p_input[1039]), .B(p_input[415]), .Z(n12379) );
  XOR U12287 ( .A(n12370), .B(n12378), .Z(n12402) );
  XOR U12288 ( .A(n12403), .B(n12375), .Z(n12378) );
  XOR U12289 ( .A(p_input[1037]), .B(p_input[413]), .Z(n12375) );
  XNOR U12290 ( .A(p_input[1038]), .B(p_input[414]), .Z(n12403) );
  XOR U12291 ( .A(p_input[1033]), .B(p_input[409]), .Z(n12370) );
  XNOR U12292 ( .A(n12386), .B(n12385), .Z(n12368) );
  XNOR U12293 ( .A(n12404), .B(n12391), .Z(n12385) );
  XOR U12294 ( .A(p_input[1032]), .B(p_input[408]), .Z(n12391) );
  XOR U12295 ( .A(n12382), .B(n12390), .Z(n12404) );
  XOR U12296 ( .A(n12405), .B(n12387), .Z(n12390) );
  XOR U12297 ( .A(p_input[1030]), .B(p_input[406]), .Z(n12387) );
  XNOR U12298 ( .A(p_input[1031]), .B(p_input[407]), .Z(n12405) );
  XOR U12299 ( .A(p_input[1026]), .B(p_input[402]), .Z(n12382) );
  XNOR U12300 ( .A(n12396), .B(n12395), .Z(n12386) );
  XOR U12301 ( .A(n12406), .B(n12392), .Z(n12395) );
  XOR U12302 ( .A(p_input[1027]), .B(p_input[403]), .Z(n12392) );
  XNOR U12303 ( .A(p_input[1028]), .B(p_input[404]), .Z(n12406) );
  XOR U12304 ( .A(p_input[1029]), .B(p_input[405]), .Z(n12396) );
  XNOR U12305 ( .A(n12407), .B(n12408), .Z(n12303) );
  AND U12306 ( .A(n314), .B(n12409), .Z(n12408) );
  XNOR U12307 ( .A(n12410), .B(n12411), .Z(n314) );
  AND U12308 ( .A(n12412), .B(n12413), .Z(n12411) );
  XOR U12309 ( .A(n12410), .B(n12313), .Z(n12413) );
  XNOR U12310 ( .A(n12410), .B(n12267), .Z(n12412) );
  XOR U12311 ( .A(n12414), .B(n12415), .Z(n12410) );
  AND U12312 ( .A(n12416), .B(n12417), .Z(n12415) );
  XOR U12313 ( .A(n12414), .B(n12277), .Z(n12416) );
  XOR U12314 ( .A(n12418), .B(n12419), .Z(n12256) );
  AND U12315 ( .A(n318), .B(n12409), .Z(n12419) );
  XNOR U12316 ( .A(n12407), .B(n12418), .Z(n12409) );
  XNOR U12317 ( .A(n12420), .B(n12421), .Z(n318) );
  AND U12318 ( .A(n12422), .B(n12423), .Z(n12421) );
  XNOR U12319 ( .A(n12424), .B(n12420), .Z(n12423) );
  IV U12320 ( .A(n12313), .Z(n12424) );
  XNOR U12321 ( .A(n12425), .B(n12426), .Z(n12313) );
  AND U12322 ( .A(n321), .B(n12427), .Z(n12426) );
  XNOR U12323 ( .A(n12425), .B(n12428), .Z(n12427) );
  XNOR U12324 ( .A(n12267), .B(n12420), .Z(n12422) );
  XOR U12325 ( .A(n12429), .B(n12430), .Z(n12267) );
  AND U12326 ( .A(n329), .B(n12431), .Z(n12430) );
  XOR U12327 ( .A(n12414), .B(n12432), .Z(n12420) );
  AND U12328 ( .A(n12433), .B(n12417), .Z(n12432) );
  XNOR U12329 ( .A(n12326), .B(n12414), .Z(n12417) );
  XNOR U12330 ( .A(n12434), .B(n12435), .Z(n12326) );
  AND U12331 ( .A(n321), .B(n12436), .Z(n12435) );
  XOR U12332 ( .A(n12437), .B(n12434), .Z(n12436) );
  XNOR U12333 ( .A(n12438), .B(n12414), .Z(n12433) );
  IV U12334 ( .A(n12277), .Z(n12438) );
  XOR U12335 ( .A(n12439), .B(n12440), .Z(n12277) );
  AND U12336 ( .A(n329), .B(n12441), .Z(n12440) );
  XOR U12337 ( .A(n12442), .B(n12443), .Z(n12414) );
  AND U12338 ( .A(n12444), .B(n12445), .Z(n12443) );
  XNOR U12339 ( .A(n12351), .B(n12442), .Z(n12445) );
  XNOR U12340 ( .A(n12446), .B(n12447), .Z(n12351) );
  AND U12341 ( .A(n321), .B(n12448), .Z(n12447) );
  XNOR U12342 ( .A(n12449), .B(n12446), .Z(n12448) );
  XOR U12343 ( .A(n12442), .B(n12288), .Z(n12444) );
  XOR U12344 ( .A(n12450), .B(n12451), .Z(n12288) );
  AND U12345 ( .A(n329), .B(n12452), .Z(n12451) );
  XOR U12346 ( .A(n12453), .B(n12454), .Z(n12442) );
  AND U12347 ( .A(n12455), .B(n12456), .Z(n12454) );
  XNOR U12348 ( .A(n12453), .B(n12397), .Z(n12456) );
  XNOR U12349 ( .A(n12457), .B(n12458), .Z(n12397) );
  AND U12350 ( .A(n321), .B(n12459), .Z(n12458) );
  XOR U12351 ( .A(n12460), .B(n12457), .Z(n12459) );
  XNOR U12352 ( .A(n12461), .B(n12453), .Z(n12455) );
  IV U12353 ( .A(n12300), .Z(n12461) );
  XOR U12354 ( .A(n12462), .B(n12463), .Z(n12300) );
  AND U12355 ( .A(n329), .B(n12464), .Z(n12463) );
  AND U12356 ( .A(n12418), .B(n12407), .Z(n12453) );
  XNOR U12357 ( .A(n12465), .B(n12466), .Z(n12407) );
  AND U12358 ( .A(n321), .B(n12467), .Z(n12466) );
  XNOR U12359 ( .A(n12468), .B(n12465), .Z(n12467) );
  XNOR U12360 ( .A(n12469), .B(n12470), .Z(n321) );
  AND U12361 ( .A(n12471), .B(n12472), .Z(n12470) );
  XOR U12362 ( .A(n12428), .B(n12469), .Z(n12472) );
  AND U12363 ( .A(n12473), .B(n12474), .Z(n12428) );
  XOR U12364 ( .A(n12469), .B(n12425), .Z(n12471) );
  XNOR U12365 ( .A(n12475), .B(n12476), .Z(n12425) );
  AND U12366 ( .A(n325), .B(n12431), .Z(n12476) );
  XOR U12367 ( .A(n12429), .B(n12475), .Z(n12431) );
  XOR U12368 ( .A(n12477), .B(n12478), .Z(n12469) );
  AND U12369 ( .A(n12479), .B(n12480), .Z(n12478) );
  XNOR U12370 ( .A(n12477), .B(n12473), .Z(n12480) );
  IV U12371 ( .A(n12437), .Z(n12473) );
  XOR U12372 ( .A(n12481), .B(n12482), .Z(n12437) );
  XOR U12373 ( .A(n12483), .B(n12474), .Z(n12482) );
  AND U12374 ( .A(n12449), .B(n12484), .Z(n12474) );
  AND U12375 ( .A(n12485), .B(n12486), .Z(n12483) );
  XOR U12376 ( .A(n12487), .B(n12481), .Z(n12485) );
  XNOR U12377 ( .A(n12434), .B(n12477), .Z(n12479) );
  XNOR U12378 ( .A(n12488), .B(n12489), .Z(n12434) );
  AND U12379 ( .A(n325), .B(n12441), .Z(n12489) );
  XOR U12380 ( .A(n12488), .B(n12439), .Z(n12441) );
  XOR U12381 ( .A(n12490), .B(n12491), .Z(n12477) );
  AND U12382 ( .A(n12492), .B(n12493), .Z(n12491) );
  XNOR U12383 ( .A(n12490), .B(n12449), .Z(n12493) );
  XOR U12384 ( .A(n12494), .B(n12486), .Z(n12449) );
  XNOR U12385 ( .A(n12495), .B(n12481), .Z(n12486) );
  XOR U12386 ( .A(n12496), .B(n12497), .Z(n12481) );
  AND U12387 ( .A(n12498), .B(n12499), .Z(n12497) );
  XOR U12388 ( .A(n12500), .B(n12496), .Z(n12498) );
  XNOR U12389 ( .A(n12501), .B(n12502), .Z(n12495) );
  AND U12390 ( .A(n12503), .B(n12504), .Z(n12502) );
  XOR U12391 ( .A(n12501), .B(n12505), .Z(n12503) );
  XNOR U12392 ( .A(n12487), .B(n12484), .Z(n12494) );
  AND U12393 ( .A(n12506), .B(n12507), .Z(n12484) );
  XOR U12394 ( .A(n12508), .B(n12509), .Z(n12487) );
  AND U12395 ( .A(n12510), .B(n12511), .Z(n12509) );
  XOR U12396 ( .A(n12508), .B(n12512), .Z(n12510) );
  XNOR U12397 ( .A(n12446), .B(n12490), .Z(n12492) );
  XNOR U12398 ( .A(n12513), .B(n12514), .Z(n12446) );
  AND U12399 ( .A(n325), .B(n12452), .Z(n12514) );
  XOR U12400 ( .A(n12513), .B(n12450), .Z(n12452) );
  XOR U12401 ( .A(n12515), .B(n12516), .Z(n12490) );
  AND U12402 ( .A(n12517), .B(n12518), .Z(n12516) );
  XNOR U12403 ( .A(n12515), .B(n12506), .Z(n12518) );
  IV U12404 ( .A(n12460), .Z(n12506) );
  XNOR U12405 ( .A(n12519), .B(n12499), .Z(n12460) );
  XNOR U12406 ( .A(n12520), .B(n12505), .Z(n12499) );
  XOR U12407 ( .A(n12521), .B(n12522), .Z(n12505) );
  NOR U12408 ( .A(n12523), .B(n12524), .Z(n12522) );
  XNOR U12409 ( .A(n12521), .B(n12525), .Z(n12523) );
  XNOR U12410 ( .A(n12504), .B(n12496), .Z(n12520) );
  XOR U12411 ( .A(n12526), .B(n12527), .Z(n12496) );
  AND U12412 ( .A(n12528), .B(n12529), .Z(n12527) );
  XNOR U12413 ( .A(n12526), .B(n12530), .Z(n12528) );
  XNOR U12414 ( .A(n12531), .B(n12501), .Z(n12504) );
  XOR U12415 ( .A(n12532), .B(n12533), .Z(n12501) );
  AND U12416 ( .A(n12534), .B(n12535), .Z(n12533) );
  XOR U12417 ( .A(n12532), .B(n12536), .Z(n12534) );
  XNOR U12418 ( .A(n12537), .B(n12538), .Z(n12531) );
  NOR U12419 ( .A(n12539), .B(n12540), .Z(n12538) );
  XOR U12420 ( .A(n12537), .B(n12541), .Z(n12539) );
  XNOR U12421 ( .A(n12500), .B(n12507), .Z(n12519) );
  NOR U12422 ( .A(n12468), .B(n12542), .Z(n12507) );
  XOR U12423 ( .A(n12512), .B(n12511), .Z(n12500) );
  XNOR U12424 ( .A(n12543), .B(n12508), .Z(n12511) );
  XOR U12425 ( .A(n12544), .B(n12545), .Z(n12508) );
  AND U12426 ( .A(n12546), .B(n12547), .Z(n12545) );
  XOR U12427 ( .A(n12544), .B(n12548), .Z(n12546) );
  XNOR U12428 ( .A(n12549), .B(n12550), .Z(n12543) );
  NOR U12429 ( .A(n12551), .B(n12552), .Z(n12550) );
  XNOR U12430 ( .A(n12549), .B(n12553), .Z(n12551) );
  XOR U12431 ( .A(n12554), .B(n12555), .Z(n12512) );
  NOR U12432 ( .A(n12556), .B(n12557), .Z(n12555) );
  XNOR U12433 ( .A(n12554), .B(n12558), .Z(n12556) );
  XNOR U12434 ( .A(n12457), .B(n12515), .Z(n12517) );
  XNOR U12435 ( .A(n12559), .B(n12560), .Z(n12457) );
  AND U12436 ( .A(n325), .B(n12464), .Z(n12560) );
  XOR U12437 ( .A(n12559), .B(n12462), .Z(n12464) );
  AND U12438 ( .A(n12465), .B(n12468), .Z(n12515) );
  XOR U12439 ( .A(n12561), .B(n12542), .Z(n12468) );
  XNOR U12440 ( .A(p_input[1024]), .B(p_input[416]), .Z(n12542) );
  XOR U12441 ( .A(n12530), .B(n12529), .Z(n12561) );
  XNOR U12442 ( .A(n12562), .B(n12536), .Z(n12529) );
  XNOR U12443 ( .A(n12525), .B(n12524), .Z(n12536) );
  XOR U12444 ( .A(n12563), .B(n12521), .Z(n12524) );
  XOR U12445 ( .A(p_input[1034]), .B(p_input[426]), .Z(n12521) );
  XNOR U12446 ( .A(p_input[1035]), .B(p_input[427]), .Z(n12563) );
  XOR U12447 ( .A(p_input[1036]), .B(p_input[428]), .Z(n12525) );
  XNOR U12448 ( .A(n12535), .B(n12526), .Z(n12562) );
  XOR U12449 ( .A(p_input[1025]), .B(p_input[417]), .Z(n12526) );
  XOR U12450 ( .A(n12564), .B(n12541), .Z(n12535) );
  XNOR U12451 ( .A(p_input[1039]), .B(p_input[431]), .Z(n12541) );
  XOR U12452 ( .A(n12532), .B(n12540), .Z(n12564) );
  XOR U12453 ( .A(n12565), .B(n12537), .Z(n12540) );
  XOR U12454 ( .A(p_input[1037]), .B(p_input[429]), .Z(n12537) );
  XNOR U12455 ( .A(p_input[1038]), .B(p_input[430]), .Z(n12565) );
  XOR U12456 ( .A(p_input[1033]), .B(p_input[425]), .Z(n12532) );
  XNOR U12457 ( .A(n12548), .B(n12547), .Z(n12530) );
  XNOR U12458 ( .A(n12566), .B(n12553), .Z(n12547) );
  XOR U12459 ( .A(p_input[1032]), .B(p_input[424]), .Z(n12553) );
  XOR U12460 ( .A(n12544), .B(n12552), .Z(n12566) );
  XOR U12461 ( .A(n12567), .B(n12549), .Z(n12552) );
  XOR U12462 ( .A(p_input[1030]), .B(p_input[422]), .Z(n12549) );
  XNOR U12463 ( .A(p_input[1031]), .B(p_input[423]), .Z(n12567) );
  XOR U12464 ( .A(p_input[1026]), .B(p_input[418]), .Z(n12544) );
  XNOR U12465 ( .A(n12558), .B(n12557), .Z(n12548) );
  XOR U12466 ( .A(n12568), .B(n12554), .Z(n12557) );
  XOR U12467 ( .A(p_input[1027]), .B(p_input[419]), .Z(n12554) );
  XNOR U12468 ( .A(p_input[1028]), .B(p_input[420]), .Z(n12568) );
  XOR U12469 ( .A(p_input[1029]), .B(p_input[421]), .Z(n12558) );
  XNOR U12470 ( .A(n12569), .B(n12570), .Z(n12465) );
  AND U12471 ( .A(n325), .B(n12571), .Z(n12570) );
  XNOR U12472 ( .A(n12572), .B(n12573), .Z(n325) );
  AND U12473 ( .A(n12574), .B(n12575), .Z(n12573) );
  XOR U12474 ( .A(n12572), .B(n12475), .Z(n12575) );
  XNOR U12475 ( .A(n12572), .B(n12429), .Z(n12574) );
  XOR U12476 ( .A(n12576), .B(n12577), .Z(n12572) );
  AND U12477 ( .A(n12578), .B(n12579), .Z(n12577) );
  XOR U12478 ( .A(n12576), .B(n12439), .Z(n12578) );
  XOR U12479 ( .A(n12580), .B(n12581), .Z(n12418) );
  AND U12480 ( .A(n329), .B(n12571), .Z(n12581) );
  XNOR U12481 ( .A(n12569), .B(n12580), .Z(n12571) );
  XNOR U12482 ( .A(n12582), .B(n12583), .Z(n329) );
  AND U12483 ( .A(n12584), .B(n12585), .Z(n12583) );
  XNOR U12484 ( .A(n12586), .B(n12582), .Z(n12585) );
  IV U12485 ( .A(n12475), .Z(n12586) );
  XNOR U12486 ( .A(n12587), .B(n12588), .Z(n12475) );
  AND U12487 ( .A(n332), .B(n12589), .Z(n12588) );
  XNOR U12488 ( .A(n12587), .B(n12590), .Z(n12589) );
  XNOR U12489 ( .A(n12429), .B(n12582), .Z(n12584) );
  XOR U12490 ( .A(n12591), .B(n12592), .Z(n12429) );
  AND U12491 ( .A(n340), .B(n12593), .Z(n12592) );
  XOR U12492 ( .A(n12576), .B(n12594), .Z(n12582) );
  AND U12493 ( .A(n12595), .B(n12579), .Z(n12594) );
  XNOR U12494 ( .A(n12488), .B(n12576), .Z(n12579) );
  XNOR U12495 ( .A(n12596), .B(n12597), .Z(n12488) );
  AND U12496 ( .A(n332), .B(n12598), .Z(n12597) );
  XOR U12497 ( .A(n12599), .B(n12596), .Z(n12598) );
  XNOR U12498 ( .A(n12600), .B(n12576), .Z(n12595) );
  IV U12499 ( .A(n12439), .Z(n12600) );
  XOR U12500 ( .A(n12601), .B(n12602), .Z(n12439) );
  AND U12501 ( .A(n340), .B(n12603), .Z(n12602) );
  XOR U12502 ( .A(n12604), .B(n12605), .Z(n12576) );
  AND U12503 ( .A(n12606), .B(n12607), .Z(n12605) );
  XNOR U12504 ( .A(n12513), .B(n12604), .Z(n12607) );
  XNOR U12505 ( .A(n12608), .B(n12609), .Z(n12513) );
  AND U12506 ( .A(n332), .B(n12610), .Z(n12609) );
  XNOR U12507 ( .A(n12611), .B(n12608), .Z(n12610) );
  XOR U12508 ( .A(n12604), .B(n12450), .Z(n12606) );
  XOR U12509 ( .A(n12612), .B(n12613), .Z(n12450) );
  AND U12510 ( .A(n340), .B(n12614), .Z(n12613) );
  XOR U12511 ( .A(n12615), .B(n12616), .Z(n12604) );
  AND U12512 ( .A(n12617), .B(n12618), .Z(n12616) );
  XNOR U12513 ( .A(n12615), .B(n12559), .Z(n12618) );
  XNOR U12514 ( .A(n12619), .B(n12620), .Z(n12559) );
  AND U12515 ( .A(n332), .B(n12621), .Z(n12620) );
  XOR U12516 ( .A(n12622), .B(n12619), .Z(n12621) );
  XNOR U12517 ( .A(n12623), .B(n12615), .Z(n12617) );
  IV U12518 ( .A(n12462), .Z(n12623) );
  XOR U12519 ( .A(n12624), .B(n12625), .Z(n12462) );
  AND U12520 ( .A(n340), .B(n12626), .Z(n12625) );
  AND U12521 ( .A(n12580), .B(n12569), .Z(n12615) );
  XNOR U12522 ( .A(n12627), .B(n12628), .Z(n12569) );
  AND U12523 ( .A(n332), .B(n12629), .Z(n12628) );
  XNOR U12524 ( .A(n12630), .B(n12627), .Z(n12629) );
  XNOR U12525 ( .A(n12631), .B(n12632), .Z(n332) );
  AND U12526 ( .A(n12633), .B(n12634), .Z(n12632) );
  XOR U12527 ( .A(n12590), .B(n12631), .Z(n12634) );
  AND U12528 ( .A(n12635), .B(n12636), .Z(n12590) );
  XOR U12529 ( .A(n12631), .B(n12587), .Z(n12633) );
  XNOR U12530 ( .A(n12637), .B(n12638), .Z(n12587) );
  AND U12531 ( .A(n336), .B(n12593), .Z(n12638) );
  XOR U12532 ( .A(n12591), .B(n12637), .Z(n12593) );
  XOR U12533 ( .A(n12639), .B(n12640), .Z(n12631) );
  AND U12534 ( .A(n12641), .B(n12642), .Z(n12640) );
  XNOR U12535 ( .A(n12639), .B(n12635), .Z(n12642) );
  IV U12536 ( .A(n12599), .Z(n12635) );
  XOR U12537 ( .A(n12643), .B(n12644), .Z(n12599) );
  XOR U12538 ( .A(n12645), .B(n12636), .Z(n12644) );
  AND U12539 ( .A(n12611), .B(n12646), .Z(n12636) );
  AND U12540 ( .A(n12647), .B(n12648), .Z(n12645) );
  XOR U12541 ( .A(n12649), .B(n12643), .Z(n12647) );
  XNOR U12542 ( .A(n12596), .B(n12639), .Z(n12641) );
  XNOR U12543 ( .A(n12650), .B(n12651), .Z(n12596) );
  AND U12544 ( .A(n336), .B(n12603), .Z(n12651) );
  XOR U12545 ( .A(n12650), .B(n12601), .Z(n12603) );
  XOR U12546 ( .A(n12652), .B(n12653), .Z(n12639) );
  AND U12547 ( .A(n12654), .B(n12655), .Z(n12653) );
  XNOR U12548 ( .A(n12652), .B(n12611), .Z(n12655) );
  XOR U12549 ( .A(n12656), .B(n12648), .Z(n12611) );
  XNOR U12550 ( .A(n12657), .B(n12643), .Z(n12648) );
  XOR U12551 ( .A(n12658), .B(n12659), .Z(n12643) );
  AND U12552 ( .A(n12660), .B(n12661), .Z(n12659) );
  XOR U12553 ( .A(n12662), .B(n12658), .Z(n12660) );
  XNOR U12554 ( .A(n12663), .B(n12664), .Z(n12657) );
  AND U12555 ( .A(n12665), .B(n12666), .Z(n12664) );
  XOR U12556 ( .A(n12663), .B(n12667), .Z(n12665) );
  XNOR U12557 ( .A(n12649), .B(n12646), .Z(n12656) );
  AND U12558 ( .A(n12668), .B(n12669), .Z(n12646) );
  XOR U12559 ( .A(n12670), .B(n12671), .Z(n12649) );
  AND U12560 ( .A(n12672), .B(n12673), .Z(n12671) );
  XOR U12561 ( .A(n12670), .B(n12674), .Z(n12672) );
  XNOR U12562 ( .A(n12608), .B(n12652), .Z(n12654) );
  XNOR U12563 ( .A(n12675), .B(n12676), .Z(n12608) );
  AND U12564 ( .A(n336), .B(n12614), .Z(n12676) );
  XOR U12565 ( .A(n12675), .B(n12612), .Z(n12614) );
  XOR U12566 ( .A(n12677), .B(n12678), .Z(n12652) );
  AND U12567 ( .A(n12679), .B(n12680), .Z(n12678) );
  XNOR U12568 ( .A(n12677), .B(n12668), .Z(n12680) );
  IV U12569 ( .A(n12622), .Z(n12668) );
  XNOR U12570 ( .A(n12681), .B(n12661), .Z(n12622) );
  XNOR U12571 ( .A(n12682), .B(n12667), .Z(n12661) );
  XOR U12572 ( .A(n12683), .B(n12684), .Z(n12667) );
  NOR U12573 ( .A(n12685), .B(n12686), .Z(n12684) );
  XNOR U12574 ( .A(n12683), .B(n12687), .Z(n12685) );
  XNOR U12575 ( .A(n12666), .B(n12658), .Z(n12682) );
  XOR U12576 ( .A(n12688), .B(n12689), .Z(n12658) );
  AND U12577 ( .A(n12690), .B(n12691), .Z(n12689) );
  XNOR U12578 ( .A(n12688), .B(n12692), .Z(n12690) );
  XNOR U12579 ( .A(n12693), .B(n12663), .Z(n12666) );
  XOR U12580 ( .A(n12694), .B(n12695), .Z(n12663) );
  AND U12581 ( .A(n12696), .B(n12697), .Z(n12695) );
  XOR U12582 ( .A(n12694), .B(n12698), .Z(n12696) );
  XNOR U12583 ( .A(n12699), .B(n12700), .Z(n12693) );
  NOR U12584 ( .A(n12701), .B(n12702), .Z(n12700) );
  XOR U12585 ( .A(n12699), .B(n12703), .Z(n12701) );
  XNOR U12586 ( .A(n12662), .B(n12669), .Z(n12681) );
  NOR U12587 ( .A(n12630), .B(n12704), .Z(n12669) );
  XOR U12588 ( .A(n12674), .B(n12673), .Z(n12662) );
  XNOR U12589 ( .A(n12705), .B(n12670), .Z(n12673) );
  XOR U12590 ( .A(n12706), .B(n12707), .Z(n12670) );
  AND U12591 ( .A(n12708), .B(n12709), .Z(n12707) );
  XOR U12592 ( .A(n12706), .B(n12710), .Z(n12708) );
  XNOR U12593 ( .A(n12711), .B(n12712), .Z(n12705) );
  NOR U12594 ( .A(n12713), .B(n12714), .Z(n12712) );
  XNOR U12595 ( .A(n12711), .B(n12715), .Z(n12713) );
  XOR U12596 ( .A(n12716), .B(n12717), .Z(n12674) );
  NOR U12597 ( .A(n12718), .B(n12719), .Z(n12717) );
  XNOR U12598 ( .A(n12716), .B(n12720), .Z(n12718) );
  XNOR U12599 ( .A(n12619), .B(n12677), .Z(n12679) );
  XNOR U12600 ( .A(n12721), .B(n12722), .Z(n12619) );
  AND U12601 ( .A(n336), .B(n12626), .Z(n12722) );
  XOR U12602 ( .A(n12721), .B(n12624), .Z(n12626) );
  AND U12603 ( .A(n12627), .B(n12630), .Z(n12677) );
  XOR U12604 ( .A(n12723), .B(n12704), .Z(n12630) );
  XNOR U12605 ( .A(p_input[1024]), .B(p_input[432]), .Z(n12704) );
  XOR U12606 ( .A(n12692), .B(n12691), .Z(n12723) );
  XNOR U12607 ( .A(n12724), .B(n12698), .Z(n12691) );
  XNOR U12608 ( .A(n12687), .B(n12686), .Z(n12698) );
  XOR U12609 ( .A(n12725), .B(n12683), .Z(n12686) );
  XOR U12610 ( .A(p_input[1034]), .B(p_input[442]), .Z(n12683) );
  XNOR U12611 ( .A(p_input[1035]), .B(p_input[443]), .Z(n12725) );
  XOR U12612 ( .A(p_input[1036]), .B(p_input[444]), .Z(n12687) );
  XNOR U12613 ( .A(n12697), .B(n12688), .Z(n12724) );
  XOR U12614 ( .A(p_input[1025]), .B(p_input[433]), .Z(n12688) );
  XOR U12615 ( .A(n12726), .B(n12703), .Z(n12697) );
  XNOR U12616 ( .A(p_input[1039]), .B(p_input[447]), .Z(n12703) );
  XOR U12617 ( .A(n12694), .B(n12702), .Z(n12726) );
  XOR U12618 ( .A(n12727), .B(n12699), .Z(n12702) );
  XOR U12619 ( .A(p_input[1037]), .B(p_input[445]), .Z(n12699) );
  XNOR U12620 ( .A(p_input[1038]), .B(p_input[446]), .Z(n12727) );
  XOR U12621 ( .A(p_input[1033]), .B(p_input[441]), .Z(n12694) );
  XNOR U12622 ( .A(n12710), .B(n12709), .Z(n12692) );
  XNOR U12623 ( .A(n12728), .B(n12715), .Z(n12709) );
  XOR U12624 ( .A(p_input[1032]), .B(p_input[440]), .Z(n12715) );
  XOR U12625 ( .A(n12706), .B(n12714), .Z(n12728) );
  XOR U12626 ( .A(n12729), .B(n12711), .Z(n12714) );
  XOR U12627 ( .A(p_input[1030]), .B(p_input[438]), .Z(n12711) );
  XNOR U12628 ( .A(p_input[1031]), .B(p_input[439]), .Z(n12729) );
  XOR U12629 ( .A(p_input[1026]), .B(p_input[434]), .Z(n12706) );
  XNOR U12630 ( .A(n12720), .B(n12719), .Z(n12710) );
  XOR U12631 ( .A(n12730), .B(n12716), .Z(n12719) );
  XOR U12632 ( .A(p_input[1027]), .B(p_input[435]), .Z(n12716) );
  XNOR U12633 ( .A(p_input[1028]), .B(p_input[436]), .Z(n12730) );
  XOR U12634 ( .A(p_input[1029]), .B(p_input[437]), .Z(n12720) );
  XNOR U12635 ( .A(n12731), .B(n12732), .Z(n12627) );
  AND U12636 ( .A(n336), .B(n12733), .Z(n12732) );
  XNOR U12637 ( .A(n12734), .B(n12735), .Z(n336) );
  AND U12638 ( .A(n12736), .B(n12737), .Z(n12735) );
  XOR U12639 ( .A(n12734), .B(n12637), .Z(n12737) );
  XNOR U12640 ( .A(n12734), .B(n12591), .Z(n12736) );
  XOR U12641 ( .A(n12738), .B(n12739), .Z(n12734) );
  AND U12642 ( .A(n12740), .B(n12741), .Z(n12739) );
  XOR U12643 ( .A(n12738), .B(n12601), .Z(n12740) );
  XOR U12644 ( .A(n12742), .B(n12743), .Z(n12580) );
  AND U12645 ( .A(n340), .B(n12733), .Z(n12743) );
  XNOR U12646 ( .A(n12731), .B(n12742), .Z(n12733) );
  XNOR U12647 ( .A(n12744), .B(n12745), .Z(n340) );
  AND U12648 ( .A(n12746), .B(n12747), .Z(n12745) );
  XNOR U12649 ( .A(n12748), .B(n12744), .Z(n12747) );
  IV U12650 ( .A(n12637), .Z(n12748) );
  XNOR U12651 ( .A(n12749), .B(n12750), .Z(n12637) );
  AND U12652 ( .A(n343), .B(n12751), .Z(n12750) );
  XNOR U12653 ( .A(n12749), .B(n12752), .Z(n12751) );
  XNOR U12654 ( .A(n12591), .B(n12744), .Z(n12746) );
  XOR U12655 ( .A(n12753), .B(n12754), .Z(n12591) );
  AND U12656 ( .A(n351), .B(n12755), .Z(n12754) );
  XOR U12657 ( .A(n12738), .B(n12756), .Z(n12744) );
  AND U12658 ( .A(n12757), .B(n12741), .Z(n12756) );
  XNOR U12659 ( .A(n12650), .B(n12738), .Z(n12741) );
  XNOR U12660 ( .A(n12758), .B(n12759), .Z(n12650) );
  AND U12661 ( .A(n343), .B(n12760), .Z(n12759) );
  XOR U12662 ( .A(n12761), .B(n12758), .Z(n12760) );
  XNOR U12663 ( .A(n12762), .B(n12738), .Z(n12757) );
  IV U12664 ( .A(n12601), .Z(n12762) );
  XOR U12665 ( .A(n12763), .B(n12764), .Z(n12601) );
  AND U12666 ( .A(n351), .B(n12765), .Z(n12764) );
  XOR U12667 ( .A(n12766), .B(n12767), .Z(n12738) );
  AND U12668 ( .A(n12768), .B(n12769), .Z(n12767) );
  XNOR U12669 ( .A(n12675), .B(n12766), .Z(n12769) );
  XNOR U12670 ( .A(n12770), .B(n12771), .Z(n12675) );
  AND U12671 ( .A(n343), .B(n12772), .Z(n12771) );
  XNOR U12672 ( .A(n12773), .B(n12770), .Z(n12772) );
  XOR U12673 ( .A(n12766), .B(n12612), .Z(n12768) );
  XOR U12674 ( .A(n12774), .B(n12775), .Z(n12612) );
  AND U12675 ( .A(n351), .B(n12776), .Z(n12775) );
  XOR U12676 ( .A(n12777), .B(n12778), .Z(n12766) );
  AND U12677 ( .A(n12779), .B(n12780), .Z(n12778) );
  XNOR U12678 ( .A(n12777), .B(n12721), .Z(n12780) );
  XNOR U12679 ( .A(n12781), .B(n12782), .Z(n12721) );
  AND U12680 ( .A(n343), .B(n12783), .Z(n12782) );
  XOR U12681 ( .A(n12784), .B(n12781), .Z(n12783) );
  XNOR U12682 ( .A(n12785), .B(n12777), .Z(n12779) );
  IV U12683 ( .A(n12624), .Z(n12785) );
  XOR U12684 ( .A(n12786), .B(n12787), .Z(n12624) );
  AND U12685 ( .A(n351), .B(n12788), .Z(n12787) );
  AND U12686 ( .A(n12742), .B(n12731), .Z(n12777) );
  XNOR U12687 ( .A(n12789), .B(n12790), .Z(n12731) );
  AND U12688 ( .A(n343), .B(n12791), .Z(n12790) );
  XNOR U12689 ( .A(n12792), .B(n12789), .Z(n12791) );
  XNOR U12690 ( .A(n12793), .B(n12794), .Z(n343) );
  AND U12691 ( .A(n12795), .B(n12796), .Z(n12794) );
  XOR U12692 ( .A(n12752), .B(n12793), .Z(n12796) );
  AND U12693 ( .A(n12797), .B(n12798), .Z(n12752) );
  XOR U12694 ( .A(n12793), .B(n12749), .Z(n12795) );
  XNOR U12695 ( .A(n12799), .B(n12800), .Z(n12749) );
  AND U12696 ( .A(n347), .B(n12755), .Z(n12800) );
  XOR U12697 ( .A(n12753), .B(n12799), .Z(n12755) );
  XOR U12698 ( .A(n12801), .B(n12802), .Z(n12793) );
  AND U12699 ( .A(n12803), .B(n12804), .Z(n12802) );
  XNOR U12700 ( .A(n12801), .B(n12797), .Z(n12804) );
  IV U12701 ( .A(n12761), .Z(n12797) );
  XOR U12702 ( .A(n12805), .B(n12806), .Z(n12761) );
  XOR U12703 ( .A(n12807), .B(n12798), .Z(n12806) );
  AND U12704 ( .A(n12773), .B(n12808), .Z(n12798) );
  AND U12705 ( .A(n12809), .B(n12810), .Z(n12807) );
  XOR U12706 ( .A(n12811), .B(n12805), .Z(n12809) );
  XNOR U12707 ( .A(n12758), .B(n12801), .Z(n12803) );
  XNOR U12708 ( .A(n12812), .B(n12813), .Z(n12758) );
  AND U12709 ( .A(n347), .B(n12765), .Z(n12813) );
  XOR U12710 ( .A(n12812), .B(n12763), .Z(n12765) );
  XOR U12711 ( .A(n12814), .B(n12815), .Z(n12801) );
  AND U12712 ( .A(n12816), .B(n12817), .Z(n12815) );
  XNOR U12713 ( .A(n12814), .B(n12773), .Z(n12817) );
  XOR U12714 ( .A(n12818), .B(n12810), .Z(n12773) );
  XNOR U12715 ( .A(n12819), .B(n12805), .Z(n12810) );
  XOR U12716 ( .A(n12820), .B(n12821), .Z(n12805) );
  AND U12717 ( .A(n12822), .B(n12823), .Z(n12821) );
  XOR U12718 ( .A(n12824), .B(n12820), .Z(n12822) );
  XNOR U12719 ( .A(n12825), .B(n12826), .Z(n12819) );
  AND U12720 ( .A(n12827), .B(n12828), .Z(n12826) );
  XOR U12721 ( .A(n12825), .B(n12829), .Z(n12827) );
  XNOR U12722 ( .A(n12811), .B(n12808), .Z(n12818) );
  AND U12723 ( .A(n12830), .B(n12831), .Z(n12808) );
  XOR U12724 ( .A(n12832), .B(n12833), .Z(n12811) );
  AND U12725 ( .A(n12834), .B(n12835), .Z(n12833) );
  XOR U12726 ( .A(n12832), .B(n12836), .Z(n12834) );
  XNOR U12727 ( .A(n12770), .B(n12814), .Z(n12816) );
  XNOR U12728 ( .A(n12837), .B(n12838), .Z(n12770) );
  AND U12729 ( .A(n347), .B(n12776), .Z(n12838) );
  XOR U12730 ( .A(n12837), .B(n12774), .Z(n12776) );
  XOR U12731 ( .A(n12839), .B(n12840), .Z(n12814) );
  AND U12732 ( .A(n12841), .B(n12842), .Z(n12840) );
  XNOR U12733 ( .A(n12839), .B(n12830), .Z(n12842) );
  IV U12734 ( .A(n12784), .Z(n12830) );
  XNOR U12735 ( .A(n12843), .B(n12823), .Z(n12784) );
  XNOR U12736 ( .A(n12844), .B(n12829), .Z(n12823) );
  XOR U12737 ( .A(n12845), .B(n12846), .Z(n12829) );
  NOR U12738 ( .A(n12847), .B(n12848), .Z(n12846) );
  XNOR U12739 ( .A(n12845), .B(n12849), .Z(n12847) );
  XNOR U12740 ( .A(n12828), .B(n12820), .Z(n12844) );
  XOR U12741 ( .A(n12850), .B(n12851), .Z(n12820) );
  AND U12742 ( .A(n12852), .B(n12853), .Z(n12851) );
  XNOR U12743 ( .A(n12850), .B(n12854), .Z(n12852) );
  XNOR U12744 ( .A(n12855), .B(n12825), .Z(n12828) );
  XOR U12745 ( .A(n12856), .B(n12857), .Z(n12825) );
  AND U12746 ( .A(n12858), .B(n12859), .Z(n12857) );
  XOR U12747 ( .A(n12856), .B(n12860), .Z(n12858) );
  XNOR U12748 ( .A(n12861), .B(n12862), .Z(n12855) );
  NOR U12749 ( .A(n12863), .B(n12864), .Z(n12862) );
  XOR U12750 ( .A(n12861), .B(n12865), .Z(n12863) );
  XNOR U12751 ( .A(n12824), .B(n12831), .Z(n12843) );
  NOR U12752 ( .A(n12792), .B(n12866), .Z(n12831) );
  XOR U12753 ( .A(n12836), .B(n12835), .Z(n12824) );
  XNOR U12754 ( .A(n12867), .B(n12832), .Z(n12835) );
  XOR U12755 ( .A(n12868), .B(n12869), .Z(n12832) );
  AND U12756 ( .A(n12870), .B(n12871), .Z(n12869) );
  XOR U12757 ( .A(n12868), .B(n12872), .Z(n12870) );
  XNOR U12758 ( .A(n12873), .B(n12874), .Z(n12867) );
  NOR U12759 ( .A(n12875), .B(n12876), .Z(n12874) );
  XNOR U12760 ( .A(n12873), .B(n12877), .Z(n12875) );
  XOR U12761 ( .A(n12878), .B(n12879), .Z(n12836) );
  NOR U12762 ( .A(n12880), .B(n12881), .Z(n12879) );
  XNOR U12763 ( .A(n12878), .B(n12882), .Z(n12880) );
  XNOR U12764 ( .A(n12781), .B(n12839), .Z(n12841) );
  XNOR U12765 ( .A(n12883), .B(n12884), .Z(n12781) );
  AND U12766 ( .A(n347), .B(n12788), .Z(n12884) );
  XOR U12767 ( .A(n12883), .B(n12786), .Z(n12788) );
  AND U12768 ( .A(n12789), .B(n12792), .Z(n12839) );
  XOR U12769 ( .A(n12885), .B(n12866), .Z(n12792) );
  XNOR U12770 ( .A(p_input[1024]), .B(p_input[448]), .Z(n12866) );
  XOR U12771 ( .A(n12854), .B(n12853), .Z(n12885) );
  XNOR U12772 ( .A(n12886), .B(n12860), .Z(n12853) );
  XNOR U12773 ( .A(n12849), .B(n12848), .Z(n12860) );
  XOR U12774 ( .A(n12887), .B(n12845), .Z(n12848) );
  XOR U12775 ( .A(p_input[1034]), .B(p_input[458]), .Z(n12845) );
  XNOR U12776 ( .A(p_input[1035]), .B(p_input[459]), .Z(n12887) );
  XOR U12777 ( .A(p_input[1036]), .B(p_input[460]), .Z(n12849) );
  XNOR U12778 ( .A(n12859), .B(n12850), .Z(n12886) );
  XOR U12779 ( .A(p_input[1025]), .B(p_input[449]), .Z(n12850) );
  XOR U12780 ( .A(n12888), .B(n12865), .Z(n12859) );
  XNOR U12781 ( .A(p_input[1039]), .B(p_input[463]), .Z(n12865) );
  XOR U12782 ( .A(n12856), .B(n12864), .Z(n12888) );
  XOR U12783 ( .A(n12889), .B(n12861), .Z(n12864) );
  XOR U12784 ( .A(p_input[1037]), .B(p_input[461]), .Z(n12861) );
  XNOR U12785 ( .A(p_input[1038]), .B(p_input[462]), .Z(n12889) );
  XOR U12786 ( .A(p_input[1033]), .B(p_input[457]), .Z(n12856) );
  XNOR U12787 ( .A(n12872), .B(n12871), .Z(n12854) );
  XNOR U12788 ( .A(n12890), .B(n12877), .Z(n12871) );
  XOR U12789 ( .A(p_input[1032]), .B(p_input[456]), .Z(n12877) );
  XOR U12790 ( .A(n12868), .B(n12876), .Z(n12890) );
  XOR U12791 ( .A(n12891), .B(n12873), .Z(n12876) );
  XOR U12792 ( .A(p_input[1030]), .B(p_input[454]), .Z(n12873) );
  XNOR U12793 ( .A(p_input[1031]), .B(p_input[455]), .Z(n12891) );
  XOR U12794 ( .A(p_input[1026]), .B(p_input[450]), .Z(n12868) );
  XNOR U12795 ( .A(n12882), .B(n12881), .Z(n12872) );
  XOR U12796 ( .A(n12892), .B(n12878), .Z(n12881) );
  XOR U12797 ( .A(p_input[1027]), .B(p_input[451]), .Z(n12878) );
  XNOR U12798 ( .A(p_input[1028]), .B(p_input[452]), .Z(n12892) );
  XOR U12799 ( .A(p_input[1029]), .B(p_input[453]), .Z(n12882) );
  XNOR U12800 ( .A(n12893), .B(n12894), .Z(n12789) );
  AND U12801 ( .A(n347), .B(n12895), .Z(n12894) );
  XNOR U12802 ( .A(n12896), .B(n12897), .Z(n347) );
  AND U12803 ( .A(n12898), .B(n12899), .Z(n12897) );
  XOR U12804 ( .A(n12896), .B(n12799), .Z(n12899) );
  XNOR U12805 ( .A(n12896), .B(n12753), .Z(n12898) );
  XOR U12806 ( .A(n12900), .B(n12901), .Z(n12896) );
  AND U12807 ( .A(n12902), .B(n12903), .Z(n12901) );
  XOR U12808 ( .A(n12900), .B(n12763), .Z(n12902) );
  XOR U12809 ( .A(n12904), .B(n12905), .Z(n12742) );
  AND U12810 ( .A(n351), .B(n12895), .Z(n12905) );
  XNOR U12811 ( .A(n12893), .B(n12904), .Z(n12895) );
  XNOR U12812 ( .A(n12906), .B(n12907), .Z(n351) );
  AND U12813 ( .A(n12908), .B(n12909), .Z(n12907) );
  XNOR U12814 ( .A(n12910), .B(n12906), .Z(n12909) );
  IV U12815 ( .A(n12799), .Z(n12910) );
  XNOR U12816 ( .A(n12911), .B(n12912), .Z(n12799) );
  AND U12817 ( .A(n354), .B(n12913), .Z(n12912) );
  XNOR U12818 ( .A(n12911), .B(n12914), .Z(n12913) );
  XNOR U12819 ( .A(n12753), .B(n12906), .Z(n12908) );
  XOR U12820 ( .A(n12915), .B(n12916), .Z(n12753) );
  AND U12821 ( .A(n362), .B(n12917), .Z(n12916) );
  XOR U12822 ( .A(n12900), .B(n12918), .Z(n12906) );
  AND U12823 ( .A(n12919), .B(n12903), .Z(n12918) );
  XNOR U12824 ( .A(n12812), .B(n12900), .Z(n12903) );
  XNOR U12825 ( .A(n12920), .B(n12921), .Z(n12812) );
  AND U12826 ( .A(n354), .B(n12922), .Z(n12921) );
  XOR U12827 ( .A(n12923), .B(n12920), .Z(n12922) );
  XNOR U12828 ( .A(n12924), .B(n12900), .Z(n12919) );
  IV U12829 ( .A(n12763), .Z(n12924) );
  XOR U12830 ( .A(n12925), .B(n12926), .Z(n12763) );
  AND U12831 ( .A(n362), .B(n12927), .Z(n12926) );
  XOR U12832 ( .A(n12928), .B(n12929), .Z(n12900) );
  AND U12833 ( .A(n12930), .B(n12931), .Z(n12929) );
  XNOR U12834 ( .A(n12837), .B(n12928), .Z(n12931) );
  XNOR U12835 ( .A(n12932), .B(n12933), .Z(n12837) );
  AND U12836 ( .A(n354), .B(n12934), .Z(n12933) );
  XNOR U12837 ( .A(n12935), .B(n12932), .Z(n12934) );
  XOR U12838 ( .A(n12928), .B(n12774), .Z(n12930) );
  XOR U12839 ( .A(n12936), .B(n12937), .Z(n12774) );
  AND U12840 ( .A(n362), .B(n12938), .Z(n12937) );
  XOR U12841 ( .A(n12939), .B(n12940), .Z(n12928) );
  AND U12842 ( .A(n12941), .B(n12942), .Z(n12940) );
  XNOR U12843 ( .A(n12939), .B(n12883), .Z(n12942) );
  XNOR U12844 ( .A(n12943), .B(n12944), .Z(n12883) );
  AND U12845 ( .A(n354), .B(n12945), .Z(n12944) );
  XOR U12846 ( .A(n12946), .B(n12943), .Z(n12945) );
  XNOR U12847 ( .A(n12947), .B(n12939), .Z(n12941) );
  IV U12848 ( .A(n12786), .Z(n12947) );
  XOR U12849 ( .A(n12948), .B(n12949), .Z(n12786) );
  AND U12850 ( .A(n362), .B(n12950), .Z(n12949) );
  AND U12851 ( .A(n12904), .B(n12893), .Z(n12939) );
  XNOR U12852 ( .A(n12951), .B(n12952), .Z(n12893) );
  AND U12853 ( .A(n354), .B(n12953), .Z(n12952) );
  XNOR U12854 ( .A(n12954), .B(n12951), .Z(n12953) );
  XNOR U12855 ( .A(n12955), .B(n12956), .Z(n354) );
  AND U12856 ( .A(n12957), .B(n12958), .Z(n12956) );
  XOR U12857 ( .A(n12914), .B(n12955), .Z(n12958) );
  AND U12858 ( .A(n12959), .B(n12960), .Z(n12914) );
  XOR U12859 ( .A(n12955), .B(n12911), .Z(n12957) );
  XNOR U12860 ( .A(n12961), .B(n12962), .Z(n12911) );
  AND U12861 ( .A(n358), .B(n12917), .Z(n12962) );
  XOR U12862 ( .A(n12915), .B(n12961), .Z(n12917) );
  XOR U12863 ( .A(n12963), .B(n12964), .Z(n12955) );
  AND U12864 ( .A(n12965), .B(n12966), .Z(n12964) );
  XNOR U12865 ( .A(n12963), .B(n12959), .Z(n12966) );
  IV U12866 ( .A(n12923), .Z(n12959) );
  XOR U12867 ( .A(n12967), .B(n12968), .Z(n12923) );
  XOR U12868 ( .A(n12969), .B(n12960), .Z(n12968) );
  AND U12869 ( .A(n12935), .B(n12970), .Z(n12960) );
  AND U12870 ( .A(n12971), .B(n12972), .Z(n12969) );
  XOR U12871 ( .A(n12973), .B(n12967), .Z(n12971) );
  XNOR U12872 ( .A(n12920), .B(n12963), .Z(n12965) );
  XNOR U12873 ( .A(n12974), .B(n12975), .Z(n12920) );
  AND U12874 ( .A(n358), .B(n12927), .Z(n12975) );
  XOR U12875 ( .A(n12974), .B(n12925), .Z(n12927) );
  XOR U12876 ( .A(n12976), .B(n12977), .Z(n12963) );
  AND U12877 ( .A(n12978), .B(n12979), .Z(n12977) );
  XNOR U12878 ( .A(n12976), .B(n12935), .Z(n12979) );
  XOR U12879 ( .A(n12980), .B(n12972), .Z(n12935) );
  XNOR U12880 ( .A(n12981), .B(n12967), .Z(n12972) );
  XOR U12881 ( .A(n12982), .B(n12983), .Z(n12967) );
  AND U12882 ( .A(n12984), .B(n12985), .Z(n12983) );
  XOR U12883 ( .A(n12986), .B(n12982), .Z(n12984) );
  XNOR U12884 ( .A(n12987), .B(n12988), .Z(n12981) );
  AND U12885 ( .A(n12989), .B(n12990), .Z(n12988) );
  XOR U12886 ( .A(n12987), .B(n12991), .Z(n12989) );
  XNOR U12887 ( .A(n12973), .B(n12970), .Z(n12980) );
  AND U12888 ( .A(n12992), .B(n12993), .Z(n12970) );
  XOR U12889 ( .A(n12994), .B(n12995), .Z(n12973) );
  AND U12890 ( .A(n12996), .B(n12997), .Z(n12995) );
  XOR U12891 ( .A(n12994), .B(n12998), .Z(n12996) );
  XNOR U12892 ( .A(n12932), .B(n12976), .Z(n12978) );
  XNOR U12893 ( .A(n12999), .B(n13000), .Z(n12932) );
  AND U12894 ( .A(n358), .B(n12938), .Z(n13000) );
  XOR U12895 ( .A(n12999), .B(n12936), .Z(n12938) );
  XOR U12896 ( .A(n13001), .B(n13002), .Z(n12976) );
  AND U12897 ( .A(n13003), .B(n13004), .Z(n13002) );
  XNOR U12898 ( .A(n13001), .B(n12992), .Z(n13004) );
  IV U12899 ( .A(n12946), .Z(n12992) );
  XNOR U12900 ( .A(n13005), .B(n12985), .Z(n12946) );
  XNOR U12901 ( .A(n13006), .B(n12991), .Z(n12985) );
  XOR U12902 ( .A(n13007), .B(n13008), .Z(n12991) );
  NOR U12903 ( .A(n13009), .B(n13010), .Z(n13008) );
  XNOR U12904 ( .A(n13007), .B(n13011), .Z(n13009) );
  XNOR U12905 ( .A(n12990), .B(n12982), .Z(n13006) );
  XOR U12906 ( .A(n13012), .B(n13013), .Z(n12982) );
  AND U12907 ( .A(n13014), .B(n13015), .Z(n13013) );
  XNOR U12908 ( .A(n13012), .B(n13016), .Z(n13014) );
  XNOR U12909 ( .A(n13017), .B(n12987), .Z(n12990) );
  XOR U12910 ( .A(n13018), .B(n13019), .Z(n12987) );
  AND U12911 ( .A(n13020), .B(n13021), .Z(n13019) );
  XOR U12912 ( .A(n13018), .B(n13022), .Z(n13020) );
  XNOR U12913 ( .A(n13023), .B(n13024), .Z(n13017) );
  NOR U12914 ( .A(n13025), .B(n13026), .Z(n13024) );
  XOR U12915 ( .A(n13023), .B(n13027), .Z(n13025) );
  XNOR U12916 ( .A(n12986), .B(n12993), .Z(n13005) );
  NOR U12917 ( .A(n12954), .B(n13028), .Z(n12993) );
  XOR U12918 ( .A(n12998), .B(n12997), .Z(n12986) );
  XNOR U12919 ( .A(n13029), .B(n12994), .Z(n12997) );
  XOR U12920 ( .A(n13030), .B(n13031), .Z(n12994) );
  AND U12921 ( .A(n13032), .B(n13033), .Z(n13031) );
  XOR U12922 ( .A(n13030), .B(n13034), .Z(n13032) );
  XNOR U12923 ( .A(n13035), .B(n13036), .Z(n13029) );
  NOR U12924 ( .A(n13037), .B(n13038), .Z(n13036) );
  XNOR U12925 ( .A(n13035), .B(n13039), .Z(n13037) );
  XOR U12926 ( .A(n13040), .B(n13041), .Z(n12998) );
  NOR U12927 ( .A(n13042), .B(n13043), .Z(n13041) );
  XNOR U12928 ( .A(n13040), .B(n13044), .Z(n13042) );
  XNOR U12929 ( .A(n12943), .B(n13001), .Z(n13003) );
  XNOR U12930 ( .A(n13045), .B(n13046), .Z(n12943) );
  AND U12931 ( .A(n358), .B(n12950), .Z(n13046) );
  XOR U12932 ( .A(n13045), .B(n12948), .Z(n12950) );
  AND U12933 ( .A(n12951), .B(n12954), .Z(n13001) );
  XOR U12934 ( .A(n13047), .B(n13028), .Z(n12954) );
  XNOR U12935 ( .A(p_input[1024]), .B(p_input[464]), .Z(n13028) );
  XOR U12936 ( .A(n13016), .B(n13015), .Z(n13047) );
  XNOR U12937 ( .A(n13048), .B(n13022), .Z(n13015) );
  XNOR U12938 ( .A(n13011), .B(n13010), .Z(n13022) );
  XOR U12939 ( .A(n13049), .B(n13007), .Z(n13010) );
  XOR U12940 ( .A(p_input[1034]), .B(p_input[474]), .Z(n13007) );
  XNOR U12941 ( .A(p_input[1035]), .B(p_input[475]), .Z(n13049) );
  XOR U12942 ( .A(p_input[1036]), .B(p_input[476]), .Z(n13011) );
  XNOR U12943 ( .A(n13021), .B(n13012), .Z(n13048) );
  XOR U12944 ( .A(p_input[1025]), .B(p_input[465]), .Z(n13012) );
  XOR U12945 ( .A(n13050), .B(n13027), .Z(n13021) );
  XNOR U12946 ( .A(p_input[1039]), .B(p_input[479]), .Z(n13027) );
  XOR U12947 ( .A(n13018), .B(n13026), .Z(n13050) );
  XOR U12948 ( .A(n13051), .B(n13023), .Z(n13026) );
  XOR U12949 ( .A(p_input[1037]), .B(p_input[477]), .Z(n13023) );
  XNOR U12950 ( .A(p_input[1038]), .B(p_input[478]), .Z(n13051) );
  XOR U12951 ( .A(p_input[1033]), .B(p_input[473]), .Z(n13018) );
  XNOR U12952 ( .A(n13034), .B(n13033), .Z(n13016) );
  XNOR U12953 ( .A(n13052), .B(n13039), .Z(n13033) );
  XOR U12954 ( .A(p_input[1032]), .B(p_input[472]), .Z(n13039) );
  XOR U12955 ( .A(n13030), .B(n13038), .Z(n13052) );
  XOR U12956 ( .A(n13053), .B(n13035), .Z(n13038) );
  XOR U12957 ( .A(p_input[1030]), .B(p_input[470]), .Z(n13035) );
  XNOR U12958 ( .A(p_input[1031]), .B(p_input[471]), .Z(n13053) );
  XOR U12959 ( .A(p_input[1026]), .B(p_input[466]), .Z(n13030) );
  XNOR U12960 ( .A(n13044), .B(n13043), .Z(n13034) );
  XOR U12961 ( .A(n13054), .B(n13040), .Z(n13043) );
  XOR U12962 ( .A(p_input[1027]), .B(p_input[467]), .Z(n13040) );
  XNOR U12963 ( .A(p_input[1028]), .B(p_input[468]), .Z(n13054) );
  XOR U12964 ( .A(p_input[1029]), .B(p_input[469]), .Z(n13044) );
  XNOR U12965 ( .A(n13055), .B(n13056), .Z(n12951) );
  AND U12966 ( .A(n358), .B(n13057), .Z(n13056) );
  XNOR U12967 ( .A(n13058), .B(n13059), .Z(n358) );
  AND U12968 ( .A(n13060), .B(n13061), .Z(n13059) );
  XOR U12969 ( .A(n13058), .B(n12961), .Z(n13061) );
  XNOR U12970 ( .A(n13058), .B(n12915), .Z(n13060) );
  XOR U12971 ( .A(n13062), .B(n13063), .Z(n13058) );
  AND U12972 ( .A(n13064), .B(n13065), .Z(n13063) );
  XOR U12973 ( .A(n13062), .B(n12925), .Z(n13064) );
  XOR U12974 ( .A(n13066), .B(n13067), .Z(n12904) );
  AND U12975 ( .A(n362), .B(n13057), .Z(n13067) );
  XNOR U12976 ( .A(n13055), .B(n13066), .Z(n13057) );
  XNOR U12977 ( .A(n13068), .B(n13069), .Z(n362) );
  AND U12978 ( .A(n13070), .B(n13071), .Z(n13069) );
  XNOR U12979 ( .A(n13072), .B(n13068), .Z(n13071) );
  IV U12980 ( .A(n12961), .Z(n13072) );
  XNOR U12981 ( .A(n13073), .B(n13074), .Z(n12961) );
  AND U12982 ( .A(n365), .B(n13075), .Z(n13074) );
  XNOR U12983 ( .A(n13073), .B(n13076), .Z(n13075) );
  XNOR U12984 ( .A(n12915), .B(n13068), .Z(n13070) );
  XOR U12985 ( .A(n13077), .B(n13078), .Z(n12915) );
  AND U12986 ( .A(n373), .B(n13079), .Z(n13078) );
  XOR U12987 ( .A(n13062), .B(n13080), .Z(n13068) );
  AND U12988 ( .A(n13081), .B(n13065), .Z(n13080) );
  XNOR U12989 ( .A(n12974), .B(n13062), .Z(n13065) );
  XNOR U12990 ( .A(n13082), .B(n13083), .Z(n12974) );
  AND U12991 ( .A(n365), .B(n13084), .Z(n13083) );
  XOR U12992 ( .A(n13085), .B(n13082), .Z(n13084) );
  XNOR U12993 ( .A(n13086), .B(n13062), .Z(n13081) );
  IV U12994 ( .A(n12925), .Z(n13086) );
  XOR U12995 ( .A(n13087), .B(n13088), .Z(n12925) );
  AND U12996 ( .A(n373), .B(n13089), .Z(n13088) );
  XOR U12997 ( .A(n13090), .B(n13091), .Z(n13062) );
  AND U12998 ( .A(n13092), .B(n13093), .Z(n13091) );
  XNOR U12999 ( .A(n12999), .B(n13090), .Z(n13093) );
  XNOR U13000 ( .A(n13094), .B(n13095), .Z(n12999) );
  AND U13001 ( .A(n365), .B(n13096), .Z(n13095) );
  XNOR U13002 ( .A(n13097), .B(n13094), .Z(n13096) );
  XOR U13003 ( .A(n13090), .B(n12936), .Z(n13092) );
  XOR U13004 ( .A(n13098), .B(n13099), .Z(n12936) );
  AND U13005 ( .A(n373), .B(n13100), .Z(n13099) );
  XOR U13006 ( .A(n13101), .B(n13102), .Z(n13090) );
  AND U13007 ( .A(n13103), .B(n13104), .Z(n13102) );
  XNOR U13008 ( .A(n13101), .B(n13045), .Z(n13104) );
  XNOR U13009 ( .A(n13105), .B(n13106), .Z(n13045) );
  AND U13010 ( .A(n365), .B(n13107), .Z(n13106) );
  XOR U13011 ( .A(n13108), .B(n13105), .Z(n13107) );
  XNOR U13012 ( .A(n13109), .B(n13101), .Z(n13103) );
  IV U13013 ( .A(n12948), .Z(n13109) );
  XOR U13014 ( .A(n13110), .B(n13111), .Z(n12948) );
  AND U13015 ( .A(n373), .B(n13112), .Z(n13111) );
  AND U13016 ( .A(n13066), .B(n13055), .Z(n13101) );
  XNOR U13017 ( .A(n13113), .B(n13114), .Z(n13055) );
  AND U13018 ( .A(n365), .B(n13115), .Z(n13114) );
  XNOR U13019 ( .A(n13116), .B(n13113), .Z(n13115) );
  XNOR U13020 ( .A(n13117), .B(n13118), .Z(n365) );
  AND U13021 ( .A(n13119), .B(n13120), .Z(n13118) );
  XOR U13022 ( .A(n13076), .B(n13117), .Z(n13120) );
  AND U13023 ( .A(n13121), .B(n13122), .Z(n13076) );
  XOR U13024 ( .A(n13117), .B(n13073), .Z(n13119) );
  XNOR U13025 ( .A(n13123), .B(n13124), .Z(n13073) );
  AND U13026 ( .A(n369), .B(n13079), .Z(n13124) );
  XOR U13027 ( .A(n13077), .B(n13123), .Z(n13079) );
  XOR U13028 ( .A(n13125), .B(n13126), .Z(n13117) );
  AND U13029 ( .A(n13127), .B(n13128), .Z(n13126) );
  XNOR U13030 ( .A(n13125), .B(n13121), .Z(n13128) );
  IV U13031 ( .A(n13085), .Z(n13121) );
  XOR U13032 ( .A(n13129), .B(n13130), .Z(n13085) );
  XOR U13033 ( .A(n13131), .B(n13122), .Z(n13130) );
  AND U13034 ( .A(n13097), .B(n13132), .Z(n13122) );
  AND U13035 ( .A(n13133), .B(n13134), .Z(n13131) );
  XOR U13036 ( .A(n13135), .B(n13129), .Z(n13133) );
  XNOR U13037 ( .A(n13082), .B(n13125), .Z(n13127) );
  XNOR U13038 ( .A(n13136), .B(n13137), .Z(n13082) );
  AND U13039 ( .A(n369), .B(n13089), .Z(n13137) );
  XOR U13040 ( .A(n13136), .B(n13087), .Z(n13089) );
  XOR U13041 ( .A(n13138), .B(n13139), .Z(n13125) );
  AND U13042 ( .A(n13140), .B(n13141), .Z(n13139) );
  XNOR U13043 ( .A(n13138), .B(n13097), .Z(n13141) );
  XOR U13044 ( .A(n13142), .B(n13134), .Z(n13097) );
  XNOR U13045 ( .A(n13143), .B(n13129), .Z(n13134) );
  XOR U13046 ( .A(n13144), .B(n13145), .Z(n13129) );
  AND U13047 ( .A(n13146), .B(n13147), .Z(n13145) );
  XOR U13048 ( .A(n13148), .B(n13144), .Z(n13146) );
  XNOR U13049 ( .A(n13149), .B(n13150), .Z(n13143) );
  AND U13050 ( .A(n13151), .B(n13152), .Z(n13150) );
  XOR U13051 ( .A(n13149), .B(n13153), .Z(n13151) );
  XNOR U13052 ( .A(n13135), .B(n13132), .Z(n13142) );
  AND U13053 ( .A(n13154), .B(n13155), .Z(n13132) );
  XOR U13054 ( .A(n13156), .B(n13157), .Z(n13135) );
  AND U13055 ( .A(n13158), .B(n13159), .Z(n13157) );
  XOR U13056 ( .A(n13156), .B(n13160), .Z(n13158) );
  XNOR U13057 ( .A(n13094), .B(n13138), .Z(n13140) );
  XNOR U13058 ( .A(n13161), .B(n13162), .Z(n13094) );
  AND U13059 ( .A(n369), .B(n13100), .Z(n13162) );
  XOR U13060 ( .A(n13161), .B(n13098), .Z(n13100) );
  XOR U13061 ( .A(n13163), .B(n13164), .Z(n13138) );
  AND U13062 ( .A(n13165), .B(n13166), .Z(n13164) );
  XNOR U13063 ( .A(n13163), .B(n13154), .Z(n13166) );
  IV U13064 ( .A(n13108), .Z(n13154) );
  XNOR U13065 ( .A(n13167), .B(n13147), .Z(n13108) );
  XNOR U13066 ( .A(n13168), .B(n13153), .Z(n13147) );
  XOR U13067 ( .A(n13169), .B(n13170), .Z(n13153) );
  NOR U13068 ( .A(n13171), .B(n13172), .Z(n13170) );
  XNOR U13069 ( .A(n13169), .B(n13173), .Z(n13171) );
  XNOR U13070 ( .A(n13152), .B(n13144), .Z(n13168) );
  XOR U13071 ( .A(n13174), .B(n13175), .Z(n13144) );
  AND U13072 ( .A(n13176), .B(n13177), .Z(n13175) );
  XNOR U13073 ( .A(n13174), .B(n13178), .Z(n13176) );
  XNOR U13074 ( .A(n13179), .B(n13149), .Z(n13152) );
  XOR U13075 ( .A(n13180), .B(n13181), .Z(n13149) );
  AND U13076 ( .A(n13182), .B(n13183), .Z(n13181) );
  XOR U13077 ( .A(n13180), .B(n13184), .Z(n13182) );
  XNOR U13078 ( .A(n13185), .B(n13186), .Z(n13179) );
  NOR U13079 ( .A(n13187), .B(n13188), .Z(n13186) );
  XOR U13080 ( .A(n13185), .B(n13189), .Z(n13187) );
  XNOR U13081 ( .A(n13148), .B(n13155), .Z(n13167) );
  NOR U13082 ( .A(n13116), .B(n13190), .Z(n13155) );
  XOR U13083 ( .A(n13160), .B(n13159), .Z(n13148) );
  XNOR U13084 ( .A(n13191), .B(n13156), .Z(n13159) );
  XOR U13085 ( .A(n13192), .B(n13193), .Z(n13156) );
  AND U13086 ( .A(n13194), .B(n13195), .Z(n13193) );
  XOR U13087 ( .A(n13192), .B(n13196), .Z(n13194) );
  XNOR U13088 ( .A(n13197), .B(n13198), .Z(n13191) );
  NOR U13089 ( .A(n13199), .B(n13200), .Z(n13198) );
  XNOR U13090 ( .A(n13197), .B(n13201), .Z(n13199) );
  XOR U13091 ( .A(n13202), .B(n13203), .Z(n13160) );
  NOR U13092 ( .A(n13204), .B(n13205), .Z(n13203) );
  XNOR U13093 ( .A(n13202), .B(n13206), .Z(n13204) );
  XNOR U13094 ( .A(n13105), .B(n13163), .Z(n13165) );
  XNOR U13095 ( .A(n13207), .B(n13208), .Z(n13105) );
  AND U13096 ( .A(n369), .B(n13112), .Z(n13208) );
  XOR U13097 ( .A(n13207), .B(n13110), .Z(n13112) );
  AND U13098 ( .A(n13113), .B(n13116), .Z(n13163) );
  XOR U13099 ( .A(n13209), .B(n13190), .Z(n13116) );
  XNOR U13100 ( .A(p_input[1024]), .B(p_input[480]), .Z(n13190) );
  XOR U13101 ( .A(n13178), .B(n13177), .Z(n13209) );
  XNOR U13102 ( .A(n13210), .B(n13184), .Z(n13177) );
  XNOR U13103 ( .A(n13173), .B(n13172), .Z(n13184) );
  XOR U13104 ( .A(n13211), .B(n13169), .Z(n13172) );
  XOR U13105 ( .A(p_input[1034]), .B(p_input[490]), .Z(n13169) );
  XNOR U13106 ( .A(p_input[1035]), .B(p_input[491]), .Z(n13211) );
  XOR U13107 ( .A(p_input[1036]), .B(p_input[492]), .Z(n13173) );
  XNOR U13108 ( .A(n13183), .B(n13174), .Z(n13210) );
  XOR U13109 ( .A(p_input[1025]), .B(p_input[481]), .Z(n13174) );
  XOR U13110 ( .A(n13212), .B(n13189), .Z(n13183) );
  XNOR U13111 ( .A(p_input[1039]), .B(p_input[495]), .Z(n13189) );
  XOR U13112 ( .A(n13180), .B(n13188), .Z(n13212) );
  XOR U13113 ( .A(n13213), .B(n13185), .Z(n13188) );
  XOR U13114 ( .A(p_input[1037]), .B(p_input[493]), .Z(n13185) );
  XNOR U13115 ( .A(p_input[1038]), .B(p_input[494]), .Z(n13213) );
  XOR U13116 ( .A(p_input[1033]), .B(p_input[489]), .Z(n13180) );
  XNOR U13117 ( .A(n13196), .B(n13195), .Z(n13178) );
  XNOR U13118 ( .A(n13214), .B(n13201), .Z(n13195) );
  XOR U13119 ( .A(p_input[1032]), .B(p_input[488]), .Z(n13201) );
  XOR U13120 ( .A(n13192), .B(n13200), .Z(n13214) );
  XOR U13121 ( .A(n13215), .B(n13197), .Z(n13200) );
  XOR U13122 ( .A(p_input[1030]), .B(p_input[486]), .Z(n13197) );
  XNOR U13123 ( .A(p_input[1031]), .B(p_input[487]), .Z(n13215) );
  XOR U13124 ( .A(p_input[1026]), .B(p_input[482]), .Z(n13192) );
  XNOR U13125 ( .A(n13206), .B(n13205), .Z(n13196) );
  XOR U13126 ( .A(n13216), .B(n13202), .Z(n13205) );
  XOR U13127 ( .A(p_input[1027]), .B(p_input[483]), .Z(n13202) );
  XNOR U13128 ( .A(p_input[1028]), .B(p_input[484]), .Z(n13216) );
  XOR U13129 ( .A(p_input[1029]), .B(p_input[485]), .Z(n13206) );
  XNOR U13130 ( .A(n13217), .B(n13218), .Z(n13113) );
  AND U13131 ( .A(n369), .B(n13219), .Z(n13218) );
  XNOR U13132 ( .A(n13220), .B(n13221), .Z(n369) );
  AND U13133 ( .A(n13222), .B(n13223), .Z(n13221) );
  XOR U13134 ( .A(n13220), .B(n13123), .Z(n13223) );
  XNOR U13135 ( .A(n13220), .B(n13077), .Z(n13222) );
  XOR U13136 ( .A(n13224), .B(n13225), .Z(n13220) );
  AND U13137 ( .A(n13226), .B(n13227), .Z(n13225) );
  XOR U13138 ( .A(n13224), .B(n13087), .Z(n13226) );
  XOR U13139 ( .A(n13228), .B(n13229), .Z(n13066) );
  AND U13140 ( .A(n373), .B(n13219), .Z(n13229) );
  XNOR U13141 ( .A(n13217), .B(n13228), .Z(n13219) );
  XNOR U13142 ( .A(n13230), .B(n13231), .Z(n373) );
  AND U13143 ( .A(n13232), .B(n13233), .Z(n13231) );
  XNOR U13144 ( .A(n13234), .B(n13230), .Z(n13233) );
  IV U13145 ( .A(n13123), .Z(n13234) );
  XNOR U13146 ( .A(n13235), .B(n13236), .Z(n13123) );
  AND U13147 ( .A(n376), .B(n13237), .Z(n13236) );
  XNOR U13148 ( .A(n13235), .B(n13238), .Z(n13237) );
  XNOR U13149 ( .A(n13077), .B(n13230), .Z(n13232) );
  XOR U13150 ( .A(n13239), .B(n13240), .Z(n13077) );
  AND U13151 ( .A(n384), .B(n13241), .Z(n13240) );
  XOR U13152 ( .A(n13224), .B(n13242), .Z(n13230) );
  AND U13153 ( .A(n13243), .B(n13227), .Z(n13242) );
  XNOR U13154 ( .A(n13136), .B(n13224), .Z(n13227) );
  XNOR U13155 ( .A(n13244), .B(n13245), .Z(n13136) );
  AND U13156 ( .A(n376), .B(n13246), .Z(n13245) );
  XOR U13157 ( .A(n13247), .B(n13244), .Z(n13246) );
  XNOR U13158 ( .A(n13248), .B(n13224), .Z(n13243) );
  IV U13159 ( .A(n13087), .Z(n13248) );
  XOR U13160 ( .A(n13249), .B(n13250), .Z(n13087) );
  AND U13161 ( .A(n384), .B(n13251), .Z(n13250) );
  XOR U13162 ( .A(n13252), .B(n13253), .Z(n13224) );
  AND U13163 ( .A(n13254), .B(n13255), .Z(n13253) );
  XNOR U13164 ( .A(n13161), .B(n13252), .Z(n13255) );
  XNOR U13165 ( .A(n13256), .B(n13257), .Z(n13161) );
  AND U13166 ( .A(n376), .B(n13258), .Z(n13257) );
  XNOR U13167 ( .A(n13259), .B(n13256), .Z(n13258) );
  XOR U13168 ( .A(n13252), .B(n13098), .Z(n13254) );
  XOR U13169 ( .A(n13260), .B(n13261), .Z(n13098) );
  AND U13170 ( .A(n384), .B(n13262), .Z(n13261) );
  XOR U13171 ( .A(n13263), .B(n13264), .Z(n13252) );
  AND U13172 ( .A(n13265), .B(n13266), .Z(n13264) );
  XNOR U13173 ( .A(n13263), .B(n13207), .Z(n13266) );
  XNOR U13174 ( .A(n13267), .B(n13268), .Z(n13207) );
  AND U13175 ( .A(n376), .B(n13269), .Z(n13268) );
  XOR U13176 ( .A(n13270), .B(n13267), .Z(n13269) );
  XNOR U13177 ( .A(n13271), .B(n13263), .Z(n13265) );
  IV U13178 ( .A(n13110), .Z(n13271) );
  XOR U13179 ( .A(n13272), .B(n13273), .Z(n13110) );
  AND U13180 ( .A(n384), .B(n13274), .Z(n13273) );
  AND U13181 ( .A(n13228), .B(n13217), .Z(n13263) );
  XNOR U13182 ( .A(n13275), .B(n13276), .Z(n13217) );
  AND U13183 ( .A(n376), .B(n13277), .Z(n13276) );
  XNOR U13184 ( .A(n13278), .B(n13275), .Z(n13277) );
  XNOR U13185 ( .A(n13279), .B(n13280), .Z(n376) );
  AND U13186 ( .A(n13281), .B(n13282), .Z(n13280) );
  XOR U13187 ( .A(n13238), .B(n13279), .Z(n13282) );
  AND U13188 ( .A(n13283), .B(n13284), .Z(n13238) );
  XOR U13189 ( .A(n13279), .B(n13235), .Z(n13281) );
  XNOR U13190 ( .A(n13285), .B(n13286), .Z(n13235) );
  AND U13191 ( .A(n380), .B(n13241), .Z(n13286) );
  XOR U13192 ( .A(n13239), .B(n13285), .Z(n13241) );
  XOR U13193 ( .A(n13287), .B(n13288), .Z(n13279) );
  AND U13194 ( .A(n13289), .B(n13290), .Z(n13288) );
  XNOR U13195 ( .A(n13287), .B(n13283), .Z(n13290) );
  IV U13196 ( .A(n13247), .Z(n13283) );
  XOR U13197 ( .A(n13291), .B(n13292), .Z(n13247) );
  XOR U13198 ( .A(n13293), .B(n13284), .Z(n13292) );
  AND U13199 ( .A(n13259), .B(n13294), .Z(n13284) );
  AND U13200 ( .A(n13295), .B(n13296), .Z(n13293) );
  XOR U13201 ( .A(n13297), .B(n13291), .Z(n13295) );
  XNOR U13202 ( .A(n13244), .B(n13287), .Z(n13289) );
  XNOR U13203 ( .A(n13298), .B(n13299), .Z(n13244) );
  AND U13204 ( .A(n380), .B(n13251), .Z(n13299) );
  XOR U13205 ( .A(n13298), .B(n13249), .Z(n13251) );
  XOR U13206 ( .A(n13300), .B(n13301), .Z(n13287) );
  AND U13207 ( .A(n13302), .B(n13303), .Z(n13301) );
  XNOR U13208 ( .A(n13300), .B(n13259), .Z(n13303) );
  XOR U13209 ( .A(n13304), .B(n13296), .Z(n13259) );
  XNOR U13210 ( .A(n13305), .B(n13291), .Z(n13296) );
  XOR U13211 ( .A(n13306), .B(n13307), .Z(n13291) );
  AND U13212 ( .A(n13308), .B(n13309), .Z(n13307) );
  XOR U13213 ( .A(n13310), .B(n13306), .Z(n13308) );
  XNOR U13214 ( .A(n13311), .B(n13312), .Z(n13305) );
  AND U13215 ( .A(n13313), .B(n13314), .Z(n13312) );
  XOR U13216 ( .A(n13311), .B(n13315), .Z(n13313) );
  XNOR U13217 ( .A(n13297), .B(n13294), .Z(n13304) );
  AND U13218 ( .A(n13316), .B(n13317), .Z(n13294) );
  XOR U13219 ( .A(n13318), .B(n13319), .Z(n13297) );
  AND U13220 ( .A(n13320), .B(n13321), .Z(n13319) );
  XOR U13221 ( .A(n13318), .B(n13322), .Z(n13320) );
  XNOR U13222 ( .A(n13256), .B(n13300), .Z(n13302) );
  XNOR U13223 ( .A(n13323), .B(n13324), .Z(n13256) );
  AND U13224 ( .A(n380), .B(n13262), .Z(n13324) );
  XOR U13225 ( .A(n13323), .B(n13260), .Z(n13262) );
  XOR U13226 ( .A(n13325), .B(n13326), .Z(n13300) );
  AND U13227 ( .A(n13327), .B(n13328), .Z(n13326) );
  XNOR U13228 ( .A(n13325), .B(n13316), .Z(n13328) );
  IV U13229 ( .A(n13270), .Z(n13316) );
  XNOR U13230 ( .A(n13329), .B(n13309), .Z(n13270) );
  XNOR U13231 ( .A(n13330), .B(n13315), .Z(n13309) );
  XOR U13232 ( .A(n13331), .B(n13332), .Z(n13315) );
  NOR U13233 ( .A(n13333), .B(n13334), .Z(n13332) );
  XNOR U13234 ( .A(n13331), .B(n13335), .Z(n13333) );
  XNOR U13235 ( .A(n13314), .B(n13306), .Z(n13330) );
  XOR U13236 ( .A(n13336), .B(n13337), .Z(n13306) );
  AND U13237 ( .A(n13338), .B(n13339), .Z(n13337) );
  XNOR U13238 ( .A(n13336), .B(n13340), .Z(n13338) );
  XNOR U13239 ( .A(n13341), .B(n13311), .Z(n13314) );
  XOR U13240 ( .A(n13342), .B(n13343), .Z(n13311) );
  AND U13241 ( .A(n13344), .B(n13345), .Z(n13343) );
  XOR U13242 ( .A(n13342), .B(n13346), .Z(n13344) );
  XNOR U13243 ( .A(n13347), .B(n13348), .Z(n13341) );
  NOR U13244 ( .A(n13349), .B(n13350), .Z(n13348) );
  XOR U13245 ( .A(n13347), .B(n13351), .Z(n13349) );
  XNOR U13246 ( .A(n13310), .B(n13317), .Z(n13329) );
  NOR U13247 ( .A(n13278), .B(n13352), .Z(n13317) );
  XOR U13248 ( .A(n13322), .B(n13321), .Z(n13310) );
  XNOR U13249 ( .A(n13353), .B(n13318), .Z(n13321) );
  XOR U13250 ( .A(n13354), .B(n13355), .Z(n13318) );
  AND U13251 ( .A(n13356), .B(n13357), .Z(n13355) );
  XOR U13252 ( .A(n13354), .B(n13358), .Z(n13356) );
  XNOR U13253 ( .A(n13359), .B(n13360), .Z(n13353) );
  NOR U13254 ( .A(n13361), .B(n13362), .Z(n13360) );
  XNOR U13255 ( .A(n13359), .B(n13363), .Z(n13361) );
  XOR U13256 ( .A(n13364), .B(n13365), .Z(n13322) );
  NOR U13257 ( .A(n13366), .B(n13367), .Z(n13365) );
  XNOR U13258 ( .A(n13364), .B(n13368), .Z(n13366) );
  XNOR U13259 ( .A(n13267), .B(n13325), .Z(n13327) );
  XNOR U13260 ( .A(n13369), .B(n13370), .Z(n13267) );
  AND U13261 ( .A(n380), .B(n13274), .Z(n13370) );
  XOR U13262 ( .A(n13369), .B(n13272), .Z(n13274) );
  AND U13263 ( .A(n13275), .B(n13278), .Z(n13325) );
  XOR U13264 ( .A(n13371), .B(n13352), .Z(n13278) );
  XNOR U13265 ( .A(p_input[1024]), .B(p_input[496]), .Z(n13352) );
  XOR U13266 ( .A(n13340), .B(n13339), .Z(n13371) );
  XNOR U13267 ( .A(n13372), .B(n13346), .Z(n13339) );
  XNOR U13268 ( .A(n13335), .B(n13334), .Z(n13346) );
  XOR U13269 ( .A(n13373), .B(n13331), .Z(n13334) );
  XOR U13270 ( .A(p_input[1034]), .B(p_input[506]), .Z(n13331) );
  XNOR U13271 ( .A(p_input[1035]), .B(p_input[507]), .Z(n13373) );
  XOR U13272 ( .A(p_input[1036]), .B(p_input[508]), .Z(n13335) );
  XNOR U13273 ( .A(n13345), .B(n13336), .Z(n13372) );
  XOR U13274 ( .A(p_input[1025]), .B(p_input[497]), .Z(n13336) );
  XOR U13275 ( .A(n13374), .B(n13351), .Z(n13345) );
  XNOR U13276 ( .A(p_input[1039]), .B(p_input[511]), .Z(n13351) );
  XOR U13277 ( .A(n13342), .B(n13350), .Z(n13374) );
  XOR U13278 ( .A(n13375), .B(n13347), .Z(n13350) );
  XOR U13279 ( .A(p_input[1037]), .B(p_input[509]), .Z(n13347) );
  XNOR U13280 ( .A(p_input[1038]), .B(p_input[510]), .Z(n13375) );
  XOR U13281 ( .A(p_input[1033]), .B(p_input[505]), .Z(n13342) );
  XNOR U13282 ( .A(n13358), .B(n13357), .Z(n13340) );
  XNOR U13283 ( .A(n13376), .B(n13363), .Z(n13357) );
  XOR U13284 ( .A(p_input[1032]), .B(p_input[504]), .Z(n13363) );
  XOR U13285 ( .A(n13354), .B(n13362), .Z(n13376) );
  XOR U13286 ( .A(n13377), .B(n13359), .Z(n13362) );
  XOR U13287 ( .A(p_input[1030]), .B(p_input[502]), .Z(n13359) );
  XNOR U13288 ( .A(p_input[1031]), .B(p_input[503]), .Z(n13377) );
  XOR U13289 ( .A(p_input[1026]), .B(p_input[498]), .Z(n13354) );
  XNOR U13290 ( .A(n13368), .B(n13367), .Z(n13358) );
  XOR U13291 ( .A(n13378), .B(n13364), .Z(n13367) );
  XOR U13292 ( .A(p_input[1027]), .B(p_input[499]), .Z(n13364) );
  XNOR U13293 ( .A(p_input[1028]), .B(p_input[500]), .Z(n13378) );
  XOR U13294 ( .A(p_input[1029]), .B(p_input[501]), .Z(n13368) );
  XNOR U13295 ( .A(n13379), .B(n13380), .Z(n13275) );
  AND U13296 ( .A(n380), .B(n13381), .Z(n13380) );
  XNOR U13297 ( .A(n13382), .B(n13383), .Z(n380) );
  AND U13298 ( .A(n13384), .B(n13385), .Z(n13383) );
  XOR U13299 ( .A(n13382), .B(n13285), .Z(n13385) );
  XNOR U13300 ( .A(n13382), .B(n13239), .Z(n13384) );
  XOR U13301 ( .A(n13386), .B(n13387), .Z(n13382) );
  AND U13302 ( .A(n13388), .B(n13389), .Z(n13387) );
  XOR U13303 ( .A(n13386), .B(n13249), .Z(n13388) );
  XOR U13304 ( .A(n13390), .B(n13391), .Z(n13228) );
  AND U13305 ( .A(n384), .B(n13381), .Z(n13391) );
  XNOR U13306 ( .A(n13379), .B(n13390), .Z(n13381) );
  XNOR U13307 ( .A(n13392), .B(n13393), .Z(n384) );
  AND U13308 ( .A(n13394), .B(n13395), .Z(n13393) );
  XNOR U13309 ( .A(n13396), .B(n13392), .Z(n13395) );
  IV U13310 ( .A(n13285), .Z(n13396) );
  XNOR U13311 ( .A(n13397), .B(n13398), .Z(n13285) );
  AND U13312 ( .A(n387), .B(n13399), .Z(n13398) );
  XNOR U13313 ( .A(n13397), .B(n13400), .Z(n13399) );
  XNOR U13314 ( .A(n13239), .B(n13392), .Z(n13394) );
  XOR U13315 ( .A(n13401), .B(n13402), .Z(n13239) );
  AND U13316 ( .A(n395), .B(n13403), .Z(n13402) );
  XOR U13317 ( .A(n13386), .B(n13404), .Z(n13392) );
  AND U13318 ( .A(n13405), .B(n13389), .Z(n13404) );
  XNOR U13319 ( .A(n13298), .B(n13386), .Z(n13389) );
  XNOR U13320 ( .A(n13406), .B(n13407), .Z(n13298) );
  AND U13321 ( .A(n387), .B(n13408), .Z(n13407) );
  XOR U13322 ( .A(n13409), .B(n13406), .Z(n13408) );
  XNOR U13323 ( .A(n13410), .B(n13386), .Z(n13405) );
  IV U13324 ( .A(n13249), .Z(n13410) );
  XOR U13325 ( .A(n13411), .B(n13412), .Z(n13249) );
  AND U13326 ( .A(n395), .B(n13413), .Z(n13412) );
  XOR U13327 ( .A(n13414), .B(n13415), .Z(n13386) );
  AND U13328 ( .A(n13416), .B(n13417), .Z(n13415) );
  XNOR U13329 ( .A(n13323), .B(n13414), .Z(n13417) );
  XNOR U13330 ( .A(n13418), .B(n13419), .Z(n13323) );
  AND U13331 ( .A(n387), .B(n13420), .Z(n13419) );
  XNOR U13332 ( .A(n13421), .B(n13418), .Z(n13420) );
  XOR U13333 ( .A(n13414), .B(n13260), .Z(n13416) );
  XOR U13334 ( .A(n13422), .B(n13423), .Z(n13260) );
  AND U13335 ( .A(n395), .B(n13424), .Z(n13423) );
  XOR U13336 ( .A(n13425), .B(n13426), .Z(n13414) );
  AND U13337 ( .A(n13427), .B(n13428), .Z(n13426) );
  XNOR U13338 ( .A(n13425), .B(n13369), .Z(n13428) );
  XNOR U13339 ( .A(n13429), .B(n13430), .Z(n13369) );
  AND U13340 ( .A(n387), .B(n13431), .Z(n13430) );
  XOR U13341 ( .A(n13432), .B(n13429), .Z(n13431) );
  XNOR U13342 ( .A(n13433), .B(n13425), .Z(n13427) );
  IV U13343 ( .A(n13272), .Z(n13433) );
  XOR U13344 ( .A(n13434), .B(n13435), .Z(n13272) );
  AND U13345 ( .A(n395), .B(n13436), .Z(n13435) );
  AND U13346 ( .A(n13390), .B(n13379), .Z(n13425) );
  XNOR U13347 ( .A(n13437), .B(n13438), .Z(n13379) );
  AND U13348 ( .A(n387), .B(n13439), .Z(n13438) );
  XNOR U13349 ( .A(n13440), .B(n13437), .Z(n13439) );
  XNOR U13350 ( .A(n13441), .B(n13442), .Z(n387) );
  AND U13351 ( .A(n13443), .B(n13444), .Z(n13442) );
  XOR U13352 ( .A(n13400), .B(n13441), .Z(n13444) );
  AND U13353 ( .A(n13445), .B(n13446), .Z(n13400) );
  XOR U13354 ( .A(n13441), .B(n13397), .Z(n13443) );
  XNOR U13355 ( .A(n13447), .B(n13448), .Z(n13397) );
  AND U13356 ( .A(n391), .B(n13403), .Z(n13448) );
  XOR U13357 ( .A(n13401), .B(n13447), .Z(n13403) );
  XOR U13358 ( .A(n13449), .B(n13450), .Z(n13441) );
  AND U13359 ( .A(n13451), .B(n13452), .Z(n13450) );
  XNOR U13360 ( .A(n13449), .B(n13445), .Z(n13452) );
  IV U13361 ( .A(n13409), .Z(n13445) );
  XOR U13362 ( .A(n13453), .B(n13454), .Z(n13409) );
  XOR U13363 ( .A(n13455), .B(n13446), .Z(n13454) );
  AND U13364 ( .A(n13421), .B(n13456), .Z(n13446) );
  AND U13365 ( .A(n13457), .B(n13458), .Z(n13455) );
  XOR U13366 ( .A(n13459), .B(n13453), .Z(n13457) );
  XNOR U13367 ( .A(n13406), .B(n13449), .Z(n13451) );
  XNOR U13368 ( .A(n13460), .B(n13461), .Z(n13406) );
  AND U13369 ( .A(n391), .B(n13413), .Z(n13461) );
  XOR U13370 ( .A(n13460), .B(n13411), .Z(n13413) );
  XOR U13371 ( .A(n13462), .B(n13463), .Z(n13449) );
  AND U13372 ( .A(n13464), .B(n13465), .Z(n13463) );
  XNOR U13373 ( .A(n13462), .B(n13421), .Z(n13465) );
  XOR U13374 ( .A(n13466), .B(n13458), .Z(n13421) );
  XNOR U13375 ( .A(n13467), .B(n13453), .Z(n13458) );
  XOR U13376 ( .A(n13468), .B(n13469), .Z(n13453) );
  AND U13377 ( .A(n13470), .B(n13471), .Z(n13469) );
  XOR U13378 ( .A(n13472), .B(n13468), .Z(n13470) );
  XNOR U13379 ( .A(n13473), .B(n13474), .Z(n13467) );
  AND U13380 ( .A(n13475), .B(n13476), .Z(n13474) );
  XOR U13381 ( .A(n13473), .B(n13477), .Z(n13475) );
  XNOR U13382 ( .A(n13459), .B(n13456), .Z(n13466) );
  AND U13383 ( .A(n13478), .B(n13479), .Z(n13456) );
  XOR U13384 ( .A(n13480), .B(n13481), .Z(n13459) );
  AND U13385 ( .A(n13482), .B(n13483), .Z(n13481) );
  XOR U13386 ( .A(n13480), .B(n13484), .Z(n13482) );
  XNOR U13387 ( .A(n13418), .B(n13462), .Z(n13464) );
  XNOR U13388 ( .A(n13485), .B(n13486), .Z(n13418) );
  AND U13389 ( .A(n391), .B(n13424), .Z(n13486) );
  XOR U13390 ( .A(n13485), .B(n13422), .Z(n13424) );
  XOR U13391 ( .A(n13487), .B(n13488), .Z(n13462) );
  AND U13392 ( .A(n13489), .B(n13490), .Z(n13488) );
  XNOR U13393 ( .A(n13487), .B(n13478), .Z(n13490) );
  IV U13394 ( .A(n13432), .Z(n13478) );
  XNOR U13395 ( .A(n13491), .B(n13471), .Z(n13432) );
  XNOR U13396 ( .A(n13492), .B(n13477), .Z(n13471) );
  XOR U13397 ( .A(n13493), .B(n13494), .Z(n13477) );
  NOR U13398 ( .A(n13495), .B(n13496), .Z(n13494) );
  XNOR U13399 ( .A(n13493), .B(n13497), .Z(n13495) );
  XNOR U13400 ( .A(n13476), .B(n13468), .Z(n13492) );
  XOR U13401 ( .A(n13498), .B(n13499), .Z(n13468) );
  AND U13402 ( .A(n13500), .B(n13501), .Z(n13499) );
  XNOR U13403 ( .A(n13498), .B(n13502), .Z(n13500) );
  XNOR U13404 ( .A(n13503), .B(n13473), .Z(n13476) );
  XOR U13405 ( .A(n13504), .B(n13505), .Z(n13473) );
  AND U13406 ( .A(n13506), .B(n13507), .Z(n13505) );
  XOR U13407 ( .A(n13504), .B(n13508), .Z(n13506) );
  XNOR U13408 ( .A(n13509), .B(n13510), .Z(n13503) );
  NOR U13409 ( .A(n13511), .B(n13512), .Z(n13510) );
  XOR U13410 ( .A(n13509), .B(n13513), .Z(n13511) );
  XNOR U13411 ( .A(n13472), .B(n13479), .Z(n13491) );
  NOR U13412 ( .A(n13440), .B(n13514), .Z(n13479) );
  XOR U13413 ( .A(n13484), .B(n13483), .Z(n13472) );
  XNOR U13414 ( .A(n13515), .B(n13480), .Z(n13483) );
  XOR U13415 ( .A(n13516), .B(n13517), .Z(n13480) );
  AND U13416 ( .A(n13518), .B(n13519), .Z(n13517) );
  XOR U13417 ( .A(n13516), .B(n13520), .Z(n13518) );
  XNOR U13418 ( .A(n13521), .B(n13522), .Z(n13515) );
  NOR U13419 ( .A(n13523), .B(n13524), .Z(n13522) );
  XNOR U13420 ( .A(n13521), .B(n13525), .Z(n13523) );
  XOR U13421 ( .A(n13526), .B(n13527), .Z(n13484) );
  NOR U13422 ( .A(n13528), .B(n13529), .Z(n13527) );
  XNOR U13423 ( .A(n13526), .B(n13530), .Z(n13528) );
  XNOR U13424 ( .A(n13429), .B(n13487), .Z(n13489) );
  XNOR U13425 ( .A(n13531), .B(n13532), .Z(n13429) );
  AND U13426 ( .A(n391), .B(n13436), .Z(n13532) );
  XOR U13427 ( .A(n13531), .B(n13434), .Z(n13436) );
  AND U13428 ( .A(n13437), .B(n13440), .Z(n13487) );
  XOR U13429 ( .A(n13533), .B(n13514), .Z(n13440) );
  XNOR U13430 ( .A(p_input[1024]), .B(p_input[512]), .Z(n13514) );
  XOR U13431 ( .A(n13502), .B(n13501), .Z(n13533) );
  XNOR U13432 ( .A(n13534), .B(n13508), .Z(n13501) );
  XNOR U13433 ( .A(n13497), .B(n13496), .Z(n13508) );
  XOR U13434 ( .A(n13535), .B(n13493), .Z(n13496) );
  XOR U13435 ( .A(p_input[1034]), .B(p_input[522]), .Z(n13493) );
  XNOR U13436 ( .A(p_input[1035]), .B(p_input[523]), .Z(n13535) );
  XOR U13437 ( .A(p_input[1036]), .B(p_input[524]), .Z(n13497) );
  XNOR U13438 ( .A(n13507), .B(n13498), .Z(n13534) );
  XOR U13439 ( .A(p_input[1025]), .B(p_input[513]), .Z(n13498) );
  XOR U13440 ( .A(n13536), .B(n13513), .Z(n13507) );
  XNOR U13441 ( .A(p_input[1039]), .B(p_input[527]), .Z(n13513) );
  XOR U13442 ( .A(n13504), .B(n13512), .Z(n13536) );
  XOR U13443 ( .A(n13537), .B(n13509), .Z(n13512) );
  XOR U13444 ( .A(p_input[1037]), .B(p_input[525]), .Z(n13509) );
  XNOR U13445 ( .A(p_input[1038]), .B(p_input[526]), .Z(n13537) );
  XOR U13446 ( .A(p_input[1033]), .B(p_input[521]), .Z(n13504) );
  XNOR U13447 ( .A(n13520), .B(n13519), .Z(n13502) );
  XNOR U13448 ( .A(n13538), .B(n13525), .Z(n13519) );
  XOR U13449 ( .A(p_input[1032]), .B(p_input[520]), .Z(n13525) );
  XOR U13450 ( .A(n13516), .B(n13524), .Z(n13538) );
  XOR U13451 ( .A(n13539), .B(n13521), .Z(n13524) );
  XOR U13452 ( .A(p_input[1030]), .B(p_input[518]), .Z(n13521) );
  XNOR U13453 ( .A(p_input[1031]), .B(p_input[519]), .Z(n13539) );
  XOR U13454 ( .A(p_input[1026]), .B(p_input[514]), .Z(n13516) );
  XNOR U13455 ( .A(n13530), .B(n13529), .Z(n13520) );
  XOR U13456 ( .A(n13540), .B(n13526), .Z(n13529) );
  XOR U13457 ( .A(p_input[1027]), .B(p_input[515]), .Z(n13526) );
  XNOR U13458 ( .A(p_input[1028]), .B(p_input[516]), .Z(n13540) );
  XOR U13459 ( .A(p_input[1029]), .B(p_input[517]), .Z(n13530) );
  XNOR U13460 ( .A(n13541), .B(n13542), .Z(n13437) );
  AND U13461 ( .A(n391), .B(n13543), .Z(n13542) );
  XNOR U13462 ( .A(n13544), .B(n13545), .Z(n391) );
  AND U13463 ( .A(n13546), .B(n13547), .Z(n13545) );
  XOR U13464 ( .A(n13544), .B(n13447), .Z(n13547) );
  XNOR U13465 ( .A(n13544), .B(n13401), .Z(n13546) );
  XOR U13466 ( .A(n13548), .B(n13549), .Z(n13544) );
  AND U13467 ( .A(n13550), .B(n13551), .Z(n13549) );
  XOR U13468 ( .A(n13548), .B(n13411), .Z(n13550) );
  XOR U13469 ( .A(n13552), .B(n13553), .Z(n13390) );
  AND U13470 ( .A(n395), .B(n13543), .Z(n13553) );
  XNOR U13471 ( .A(n13541), .B(n13552), .Z(n13543) );
  XNOR U13472 ( .A(n13554), .B(n13555), .Z(n395) );
  AND U13473 ( .A(n13556), .B(n13557), .Z(n13555) );
  XNOR U13474 ( .A(n13558), .B(n13554), .Z(n13557) );
  IV U13475 ( .A(n13447), .Z(n13558) );
  XNOR U13476 ( .A(n13559), .B(n13560), .Z(n13447) );
  AND U13477 ( .A(n398), .B(n13561), .Z(n13560) );
  XNOR U13478 ( .A(n13559), .B(n13562), .Z(n13561) );
  XNOR U13479 ( .A(n13401), .B(n13554), .Z(n13556) );
  XOR U13480 ( .A(n13563), .B(n13564), .Z(n13401) );
  AND U13481 ( .A(n406), .B(n13565), .Z(n13564) );
  XOR U13482 ( .A(n13548), .B(n13566), .Z(n13554) );
  AND U13483 ( .A(n13567), .B(n13551), .Z(n13566) );
  XNOR U13484 ( .A(n13460), .B(n13548), .Z(n13551) );
  XNOR U13485 ( .A(n13568), .B(n13569), .Z(n13460) );
  AND U13486 ( .A(n398), .B(n13570), .Z(n13569) );
  XOR U13487 ( .A(n13571), .B(n13568), .Z(n13570) );
  XNOR U13488 ( .A(n13572), .B(n13548), .Z(n13567) );
  IV U13489 ( .A(n13411), .Z(n13572) );
  XOR U13490 ( .A(n13573), .B(n13574), .Z(n13411) );
  AND U13491 ( .A(n406), .B(n13575), .Z(n13574) );
  XOR U13492 ( .A(n13576), .B(n13577), .Z(n13548) );
  AND U13493 ( .A(n13578), .B(n13579), .Z(n13577) );
  XNOR U13494 ( .A(n13485), .B(n13576), .Z(n13579) );
  XNOR U13495 ( .A(n13580), .B(n13581), .Z(n13485) );
  AND U13496 ( .A(n398), .B(n13582), .Z(n13581) );
  XNOR U13497 ( .A(n13583), .B(n13580), .Z(n13582) );
  XOR U13498 ( .A(n13576), .B(n13422), .Z(n13578) );
  XOR U13499 ( .A(n13584), .B(n13585), .Z(n13422) );
  AND U13500 ( .A(n406), .B(n13586), .Z(n13585) );
  XOR U13501 ( .A(n13587), .B(n13588), .Z(n13576) );
  AND U13502 ( .A(n13589), .B(n13590), .Z(n13588) );
  XNOR U13503 ( .A(n13587), .B(n13531), .Z(n13590) );
  XNOR U13504 ( .A(n13591), .B(n13592), .Z(n13531) );
  AND U13505 ( .A(n398), .B(n13593), .Z(n13592) );
  XOR U13506 ( .A(n13594), .B(n13591), .Z(n13593) );
  XNOR U13507 ( .A(n13595), .B(n13587), .Z(n13589) );
  IV U13508 ( .A(n13434), .Z(n13595) );
  XOR U13509 ( .A(n13596), .B(n13597), .Z(n13434) );
  AND U13510 ( .A(n406), .B(n13598), .Z(n13597) );
  AND U13511 ( .A(n13552), .B(n13541), .Z(n13587) );
  XNOR U13512 ( .A(n13599), .B(n13600), .Z(n13541) );
  AND U13513 ( .A(n398), .B(n13601), .Z(n13600) );
  XNOR U13514 ( .A(n13602), .B(n13599), .Z(n13601) );
  XNOR U13515 ( .A(n13603), .B(n13604), .Z(n398) );
  AND U13516 ( .A(n13605), .B(n13606), .Z(n13604) );
  XOR U13517 ( .A(n13562), .B(n13603), .Z(n13606) );
  AND U13518 ( .A(n13607), .B(n13608), .Z(n13562) );
  XOR U13519 ( .A(n13603), .B(n13559), .Z(n13605) );
  XNOR U13520 ( .A(n13609), .B(n13610), .Z(n13559) );
  AND U13521 ( .A(n402), .B(n13565), .Z(n13610) );
  XOR U13522 ( .A(n13563), .B(n13609), .Z(n13565) );
  XOR U13523 ( .A(n13611), .B(n13612), .Z(n13603) );
  AND U13524 ( .A(n13613), .B(n13614), .Z(n13612) );
  XNOR U13525 ( .A(n13611), .B(n13607), .Z(n13614) );
  IV U13526 ( .A(n13571), .Z(n13607) );
  XOR U13527 ( .A(n13615), .B(n13616), .Z(n13571) );
  XOR U13528 ( .A(n13617), .B(n13608), .Z(n13616) );
  AND U13529 ( .A(n13583), .B(n13618), .Z(n13608) );
  AND U13530 ( .A(n13619), .B(n13620), .Z(n13617) );
  XOR U13531 ( .A(n13621), .B(n13615), .Z(n13619) );
  XNOR U13532 ( .A(n13568), .B(n13611), .Z(n13613) );
  XNOR U13533 ( .A(n13622), .B(n13623), .Z(n13568) );
  AND U13534 ( .A(n402), .B(n13575), .Z(n13623) );
  XOR U13535 ( .A(n13622), .B(n13573), .Z(n13575) );
  XOR U13536 ( .A(n13624), .B(n13625), .Z(n13611) );
  AND U13537 ( .A(n13626), .B(n13627), .Z(n13625) );
  XNOR U13538 ( .A(n13624), .B(n13583), .Z(n13627) );
  XOR U13539 ( .A(n13628), .B(n13620), .Z(n13583) );
  XNOR U13540 ( .A(n13629), .B(n13615), .Z(n13620) );
  XOR U13541 ( .A(n13630), .B(n13631), .Z(n13615) );
  AND U13542 ( .A(n13632), .B(n13633), .Z(n13631) );
  XOR U13543 ( .A(n13634), .B(n13630), .Z(n13632) );
  XNOR U13544 ( .A(n13635), .B(n13636), .Z(n13629) );
  AND U13545 ( .A(n13637), .B(n13638), .Z(n13636) );
  XOR U13546 ( .A(n13635), .B(n13639), .Z(n13637) );
  XNOR U13547 ( .A(n13621), .B(n13618), .Z(n13628) );
  AND U13548 ( .A(n13640), .B(n13641), .Z(n13618) );
  XOR U13549 ( .A(n13642), .B(n13643), .Z(n13621) );
  AND U13550 ( .A(n13644), .B(n13645), .Z(n13643) );
  XOR U13551 ( .A(n13642), .B(n13646), .Z(n13644) );
  XNOR U13552 ( .A(n13580), .B(n13624), .Z(n13626) );
  XNOR U13553 ( .A(n13647), .B(n13648), .Z(n13580) );
  AND U13554 ( .A(n402), .B(n13586), .Z(n13648) );
  XOR U13555 ( .A(n13647), .B(n13584), .Z(n13586) );
  XOR U13556 ( .A(n13649), .B(n13650), .Z(n13624) );
  AND U13557 ( .A(n13651), .B(n13652), .Z(n13650) );
  XNOR U13558 ( .A(n13649), .B(n13640), .Z(n13652) );
  IV U13559 ( .A(n13594), .Z(n13640) );
  XNOR U13560 ( .A(n13653), .B(n13633), .Z(n13594) );
  XNOR U13561 ( .A(n13654), .B(n13639), .Z(n13633) );
  XOR U13562 ( .A(n13655), .B(n13656), .Z(n13639) );
  NOR U13563 ( .A(n13657), .B(n13658), .Z(n13656) );
  XNOR U13564 ( .A(n13655), .B(n13659), .Z(n13657) );
  XNOR U13565 ( .A(n13638), .B(n13630), .Z(n13654) );
  XOR U13566 ( .A(n13660), .B(n13661), .Z(n13630) );
  AND U13567 ( .A(n13662), .B(n13663), .Z(n13661) );
  XNOR U13568 ( .A(n13660), .B(n13664), .Z(n13662) );
  XNOR U13569 ( .A(n13665), .B(n13635), .Z(n13638) );
  XOR U13570 ( .A(n13666), .B(n13667), .Z(n13635) );
  AND U13571 ( .A(n13668), .B(n13669), .Z(n13667) );
  XOR U13572 ( .A(n13666), .B(n13670), .Z(n13668) );
  XNOR U13573 ( .A(n13671), .B(n13672), .Z(n13665) );
  NOR U13574 ( .A(n13673), .B(n13674), .Z(n13672) );
  XOR U13575 ( .A(n13671), .B(n13675), .Z(n13673) );
  XNOR U13576 ( .A(n13634), .B(n13641), .Z(n13653) );
  NOR U13577 ( .A(n13602), .B(n13676), .Z(n13641) );
  XOR U13578 ( .A(n13646), .B(n13645), .Z(n13634) );
  XNOR U13579 ( .A(n13677), .B(n13642), .Z(n13645) );
  XOR U13580 ( .A(n13678), .B(n13679), .Z(n13642) );
  AND U13581 ( .A(n13680), .B(n13681), .Z(n13679) );
  XOR U13582 ( .A(n13678), .B(n13682), .Z(n13680) );
  XNOR U13583 ( .A(n13683), .B(n13684), .Z(n13677) );
  NOR U13584 ( .A(n13685), .B(n13686), .Z(n13684) );
  XNOR U13585 ( .A(n13683), .B(n13687), .Z(n13685) );
  XOR U13586 ( .A(n13688), .B(n13689), .Z(n13646) );
  NOR U13587 ( .A(n13690), .B(n13691), .Z(n13689) );
  XNOR U13588 ( .A(n13688), .B(n13692), .Z(n13690) );
  XNOR U13589 ( .A(n13591), .B(n13649), .Z(n13651) );
  XNOR U13590 ( .A(n13693), .B(n13694), .Z(n13591) );
  AND U13591 ( .A(n402), .B(n13598), .Z(n13694) );
  XOR U13592 ( .A(n13693), .B(n13596), .Z(n13598) );
  AND U13593 ( .A(n13599), .B(n13602), .Z(n13649) );
  XOR U13594 ( .A(n13695), .B(n13676), .Z(n13602) );
  XNOR U13595 ( .A(p_input[1024]), .B(p_input[528]), .Z(n13676) );
  XOR U13596 ( .A(n13664), .B(n13663), .Z(n13695) );
  XNOR U13597 ( .A(n13696), .B(n13670), .Z(n13663) );
  XNOR U13598 ( .A(n13659), .B(n13658), .Z(n13670) );
  XOR U13599 ( .A(n13697), .B(n13655), .Z(n13658) );
  XOR U13600 ( .A(p_input[1034]), .B(p_input[538]), .Z(n13655) );
  XNOR U13601 ( .A(p_input[1035]), .B(p_input[539]), .Z(n13697) );
  XOR U13602 ( .A(p_input[1036]), .B(p_input[540]), .Z(n13659) );
  XNOR U13603 ( .A(n13669), .B(n13660), .Z(n13696) );
  XOR U13604 ( .A(p_input[1025]), .B(p_input[529]), .Z(n13660) );
  XOR U13605 ( .A(n13698), .B(n13675), .Z(n13669) );
  XNOR U13606 ( .A(p_input[1039]), .B(p_input[543]), .Z(n13675) );
  XOR U13607 ( .A(n13666), .B(n13674), .Z(n13698) );
  XOR U13608 ( .A(n13699), .B(n13671), .Z(n13674) );
  XOR U13609 ( .A(p_input[1037]), .B(p_input[541]), .Z(n13671) );
  XNOR U13610 ( .A(p_input[1038]), .B(p_input[542]), .Z(n13699) );
  XOR U13611 ( .A(p_input[1033]), .B(p_input[537]), .Z(n13666) );
  XNOR U13612 ( .A(n13682), .B(n13681), .Z(n13664) );
  XNOR U13613 ( .A(n13700), .B(n13687), .Z(n13681) );
  XOR U13614 ( .A(p_input[1032]), .B(p_input[536]), .Z(n13687) );
  XOR U13615 ( .A(n13678), .B(n13686), .Z(n13700) );
  XOR U13616 ( .A(n13701), .B(n13683), .Z(n13686) );
  XOR U13617 ( .A(p_input[1030]), .B(p_input[534]), .Z(n13683) );
  XNOR U13618 ( .A(p_input[1031]), .B(p_input[535]), .Z(n13701) );
  XOR U13619 ( .A(p_input[1026]), .B(p_input[530]), .Z(n13678) );
  XNOR U13620 ( .A(n13692), .B(n13691), .Z(n13682) );
  XOR U13621 ( .A(n13702), .B(n13688), .Z(n13691) );
  XOR U13622 ( .A(p_input[1027]), .B(p_input[531]), .Z(n13688) );
  XNOR U13623 ( .A(p_input[1028]), .B(p_input[532]), .Z(n13702) );
  XOR U13624 ( .A(p_input[1029]), .B(p_input[533]), .Z(n13692) );
  XNOR U13625 ( .A(n13703), .B(n13704), .Z(n13599) );
  AND U13626 ( .A(n402), .B(n13705), .Z(n13704) );
  XNOR U13627 ( .A(n13706), .B(n13707), .Z(n402) );
  AND U13628 ( .A(n13708), .B(n13709), .Z(n13707) );
  XOR U13629 ( .A(n13706), .B(n13609), .Z(n13709) );
  XNOR U13630 ( .A(n13706), .B(n13563), .Z(n13708) );
  XOR U13631 ( .A(n13710), .B(n13711), .Z(n13706) );
  AND U13632 ( .A(n13712), .B(n13713), .Z(n13711) );
  XOR U13633 ( .A(n13710), .B(n13573), .Z(n13712) );
  XOR U13634 ( .A(n13714), .B(n13715), .Z(n13552) );
  AND U13635 ( .A(n406), .B(n13705), .Z(n13715) );
  XNOR U13636 ( .A(n13703), .B(n13714), .Z(n13705) );
  XNOR U13637 ( .A(n13716), .B(n13717), .Z(n406) );
  AND U13638 ( .A(n13718), .B(n13719), .Z(n13717) );
  XNOR U13639 ( .A(n13720), .B(n13716), .Z(n13719) );
  IV U13640 ( .A(n13609), .Z(n13720) );
  XNOR U13641 ( .A(n13721), .B(n13722), .Z(n13609) );
  AND U13642 ( .A(n409), .B(n13723), .Z(n13722) );
  XNOR U13643 ( .A(n13721), .B(n13724), .Z(n13723) );
  XNOR U13644 ( .A(n13563), .B(n13716), .Z(n13718) );
  XOR U13645 ( .A(n13725), .B(n13726), .Z(n13563) );
  AND U13646 ( .A(n417), .B(n13727), .Z(n13726) );
  XOR U13647 ( .A(n13710), .B(n13728), .Z(n13716) );
  AND U13648 ( .A(n13729), .B(n13713), .Z(n13728) );
  XNOR U13649 ( .A(n13622), .B(n13710), .Z(n13713) );
  XNOR U13650 ( .A(n13730), .B(n13731), .Z(n13622) );
  AND U13651 ( .A(n409), .B(n13732), .Z(n13731) );
  XOR U13652 ( .A(n13733), .B(n13730), .Z(n13732) );
  XNOR U13653 ( .A(n13734), .B(n13710), .Z(n13729) );
  IV U13654 ( .A(n13573), .Z(n13734) );
  XOR U13655 ( .A(n13735), .B(n13736), .Z(n13573) );
  AND U13656 ( .A(n417), .B(n13737), .Z(n13736) );
  XOR U13657 ( .A(n13738), .B(n13739), .Z(n13710) );
  AND U13658 ( .A(n13740), .B(n13741), .Z(n13739) );
  XNOR U13659 ( .A(n13647), .B(n13738), .Z(n13741) );
  XNOR U13660 ( .A(n13742), .B(n13743), .Z(n13647) );
  AND U13661 ( .A(n409), .B(n13744), .Z(n13743) );
  XNOR U13662 ( .A(n13745), .B(n13742), .Z(n13744) );
  XOR U13663 ( .A(n13738), .B(n13584), .Z(n13740) );
  XOR U13664 ( .A(n13746), .B(n13747), .Z(n13584) );
  AND U13665 ( .A(n417), .B(n13748), .Z(n13747) );
  XOR U13666 ( .A(n13749), .B(n13750), .Z(n13738) );
  AND U13667 ( .A(n13751), .B(n13752), .Z(n13750) );
  XNOR U13668 ( .A(n13749), .B(n13693), .Z(n13752) );
  XNOR U13669 ( .A(n13753), .B(n13754), .Z(n13693) );
  AND U13670 ( .A(n409), .B(n13755), .Z(n13754) );
  XOR U13671 ( .A(n13756), .B(n13753), .Z(n13755) );
  XNOR U13672 ( .A(n13757), .B(n13749), .Z(n13751) );
  IV U13673 ( .A(n13596), .Z(n13757) );
  XOR U13674 ( .A(n13758), .B(n13759), .Z(n13596) );
  AND U13675 ( .A(n417), .B(n13760), .Z(n13759) );
  AND U13676 ( .A(n13714), .B(n13703), .Z(n13749) );
  XNOR U13677 ( .A(n13761), .B(n13762), .Z(n13703) );
  AND U13678 ( .A(n409), .B(n13763), .Z(n13762) );
  XNOR U13679 ( .A(n13764), .B(n13761), .Z(n13763) );
  XNOR U13680 ( .A(n13765), .B(n13766), .Z(n409) );
  AND U13681 ( .A(n13767), .B(n13768), .Z(n13766) );
  XOR U13682 ( .A(n13724), .B(n13765), .Z(n13768) );
  AND U13683 ( .A(n13769), .B(n13770), .Z(n13724) );
  XOR U13684 ( .A(n13765), .B(n13721), .Z(n13767) );
  XNOR U13685 ( .A(n13771), .B(n13772), .Z(n13721) );
  AND U13686 ( .A(n413), .B(n13727), .Z(n13772) );
  XOR U13687 ( .A(n13725), .B(n13771), .Z(n13727) );
  XOR U13688 ( .A(n13773), .B(n13774), .Z(n13765) );
  AND U13689 ( .A(n13775), .B(n13776), .Z(n13774) );
  XNOR U13690 ( .A(n13773), .B(n13769), .Z(n13776) );
  IV U13691 ( .A(n13733), .Z(n13769) );
  XOR U13692 ( .A(n13777), .B(n13778), .Z(n13733) );
  XOR U13693 ( .A(n13779), .B(n13770), .Z(n13778) );
  AND U13694 ( .A(n13745), .B(n13780), .Z(n13770) );
  AND U13695 ( .A(n13781), .B(n13782), .Z(n13779) );
  XOR U13696 ( .A(n13783), .B(n13777), .Z(n13781) );
  XNOR U13697 ( .A(n13730), .B(n13773), .Z(n13775) );
  XNOR U13698 ( .A(n13784), .B(n13785), .Z(n13730) );
  AND U13699 ( .A(n413), .B(n13737), .Z(n13785) );
  XOR U13700 ( .A(n13784), .B(n13735), .Z(n13737) );
  XOR U13701 ( .A(n13786), .B(n13787), .Z(n13773) );
  AND U13702 ( .A(n13788), .B(n13789), .Z(n13787) );
  XNOR U13703 ( .A(n13786), .B(n13745), .Z(n13789) );
  XOR U13704 ( .A(n13790), .B(n13782), .Z(n13745) );
  XNOR U13705 ( .A(n13791), .B(n13777), .Z(n13782) );
  XOR U13706 ( .A(n13792), .B(n13793), .Z(n13777) );
  AND U13707 ( .A(n13794), .B(n13795), .Z(n13793) );
  XOR U13708 ( .A(n13796), .B(n13792), .Z(n13794) );
  XNOR U13709 ( .A(n13797), .B(n13798), .Z(n13791) );
  AND U13710 ( .A(n13799), .B(n13800), .Z(n13798) );
  XOR U13711 ( .A(n13797), .B(n13801), .Z(n13799) );
  XNOR U13712 ( .A(n13783), .B(n13780), .Z(n13790) );
  AND U13713 ( .A(n13802), .B(n13803), .Z(n13780) );
  XOR U13714 ( .A(n13804), .B(n13805), .Z(n13783) );
  AND U13715 ( .A(n13806), .B(n13807), .Z(n13805) );
  XOR U13716 ( .A(n13804), .B(n13808), .Z(n13806) );
  XNOR U13717 ( .A(n13742), .B(n13786), .Z(n13788) );
  XNOR U13718 ( .A(n13809), .B(n13810), .Z(n13742) );
  AND U13719 ( .A(n413), .B(n13748), .Z(n13810) );
  XOR U13720 ( .A(n13809), .B(n13746), .Z(n13748) );
  XOR U13721 ( .A(n13811), .B(n13812), .Z(n13786) );
  AND U13722 ( .A(n13813), .B(n13814), .Z(n13812) );
  XNOR U13723 ( .A(n13811), .B(n13802), .Z(n13814) );
  IV U13724 ( .A(n13756), .Z(n13802) );
  XNOR U13725 ( .A(n13815), .B(n13795), .Z(n13756) );
  XNOR U13726 ( .A(n13816), .B(n13801), .Z(n13795) );
  XOR U13727 ( .A(n13817), .B(n13818), .Z(n13801) );
  NOR U13728 ( .A(n13819), .B(n13820), .Z(n13818) );
  XNOR U13729 ( .A(n13817), .B(n13821), .Z(n13819) );
  XNOR U13730 ( .A(n13800), .B(n13792), .Z(n13816) );
  XOR U13731 ( .A(n13822), .B(n13823), .Z(n13792) );
  AND U13732 ( .A(n13824), .B(n13825), .Z(n13823) );
  XNOR U13733 ( .A(n13822), .B(n13826), .Z(n13824) );
  XNOR U13734 ( .A(n13827), .B(n13797), .Z(n13800) );
  XOR U13735 ( .A(n13828), .B(n13829), .Z(n13797) );
  AND U13736 ( .A(n13830), .B(n13831), .Z(n13829) );
  XOR U13737 ( .A(n13828), .B(n13832), .Z(n13830) );
  XNOR U13738 ( .A(n13833), .B(n13834), .Z(n13827) );
  NOR U13739 ( .A(n13835), .B(n13836), .Z(n13834) );
  XOR U13740 ( .A(n13833), .B(n13837), .Z(n13835) );
  XNOR U13741 ( .A(n13796), .B(n13803), .Z(n13815) );
  NOR U13742 ( .A(n13764), .B(n13838), .Z(n13803) );
  XOR U13743 ( .A(n13808), .B(n13807), .Z(n13796) );
  XNOR U13744 ( .A(n13839), .B(n13804), .Z(n13807) );
  XOR U13745 ( .A(n13840), .B(n13841), .Z(n13804) );
  AND U13746 ( .A(n13842), .B(n13843), .Z(n13841) );
  XOR U13747 ( .A(n13840), .B(n13844), .Z(n13842) );
  XNOR U13748 ( .A(n13845), .B(n13846), .Z(n13839) );
  NOR U13749 ( .A(n13847), .B(n13848), .Z(n13846) );
  XNOR U13750 ( .A(n13845), .B(n13849), .Z(n13847) );
  XOR U13751 ( .A(n13850), .B(n13851), .Z(n13808) );
  NOR U13752 ( .A(n13852), .B(n13853), .Z(n13851) );
  XNOR U13753 ( .A(n13850), .B(n13854), .Z(n13852) );
  XNOR U13754 ( .A(n13753), .B(n13811), .Z(n13813) );
  XNOR U13755 ( .A(n13855), .B(n13856), .Z(n13753) );
  AND U13756 ( .A(n413), .B(n13760), .Z(n13856) );
  XOR U13757 ( .A(n13855), .B(n13758), .Z(n13760) );
  AND U13758 ( .A(n13761), .B(n13764), .Z(n13811) );
  XOR U13759 ( .A(n13857), .B(n13838), .Z(n13764) );
  XNOR U13760 ( .A(p_input[1024]), .B(p_input[544]), .Z(n13838) );
  XOR U13761 ( .A(n13826), .B(n13825), .Z(n13857) );
  XNOR U13762 ( .A(n13858), .B(n13832), .Z(n13825) );
  XNOR U13763 ( .A(n13821), .B(n13820), .Z(n13832) );
  XOR U13764 ( .A(n13859), .B(n13817), .Z(n13820) );
  XOR U13765 ( .A(p_input[1034]), .B(p_input[554]), .Z(n13817) );
  XNOR U13766 ( .A(p_input[1035]), .B(p_input[555]), .Z(n13859) );
  XOR U13767 ( .A(p_input[1036]), .B(p_input[556]), .Z(n13821) );
  XNOR U13768 ( .A(n13831), .B(n13822), .Z(n13858) );
  XOR U13769 ( .A(p_input[1025]), .B(p_input[545]), .Z(n13822) );
  XOR U13770 ( .A(n13860), .B(n13837), .Z(n13831) );
  XNOR U13771 ( .A(p_input[1039]), .B(p_input[559]), .Z(n13837) );
  XOR U13772 ( .A(n13828), .B(n13836), .Z(n13860) );
  XOR U13773 ( .A(n13861), .B(n13833), .Z(n13836) );
  XOR U13774 ( .A(p_input[1037]), .B(p_input[557]), .Z(n13833) );
  XNOR U13775 ( .A(p_input[1038]), .B(p_input[558]), .Z(n13861) );
  XOR U13776 ( .A(p_input[1033]), .B(p_input[553]), .Z(n13828) );
  XNOR U13777 ( .A(n13844), .B(n13843), .Z(n13826) );
  XNOR U13778 ( .A(n13862), .B(n13849), .Z(n13843) );
  XOR U13779 ( .A(p_input[1032]), .B(p_input[552]), .Z(n13849) );
  XOR U13780 ( .A(n13840), .B(n13848), .Z(n13862) );
  XOR U13781 ( .A(n13863), .B(n13845), .Z(n13848) );
  XOR U13782 ( .A(p_input[1030]), .B(p_input[550]), .Z(n13845) );
  XNOR U13783 ( .A(p_input[1031]), .B(p_input[551]), .Z(n13863) );
  XOR U13784 ( .A(p_input[1026]), .B(p_input[546]), .Z(n13840) );
  XNOR U13785 ( .A(n13854), .B(n13853), .Z(n13844) );
  XOR U13786 ( .A(n13864), .B(n13850), .Z(n13853) );
  XOR U13787 ( .A(p_input[1027]), .B(p_input[547]), .Z(n13850) );
  XNOR U13788 ( .A(p_input[1028]), .B(p_input[548]), .Z(n13864) );
  XOR U13789 ( .A(p_input[1029]), .B(p_input[549]), .Z(n13854) );
  XNOR U13790 ( .A(n13865), .B(n13866), .Z(n13761) );
  AND U13791 ( .A(n413), .B(n13867), .Z(n13866) );
  XNOR U13792 ( .A(n13868), .B(n13869), .Z(n413) );
  AND U13793 ( .A(n13870), .B(n13871), .Z(n13869) );
  XOR U13794 ( .A(n13868), .B(n13771), .Z(n13871) );
  XNOR U13795 ( .A(n13868), .B(n13725), .Z(n13870) );
  XOR U13796 ( .A(n13872), .B(n13873), .Z(n13868) );
  AND U13797 ( .A(n13874), .B(n13875), .Z(n13873) );
  XOR U13798 ( .A(n13872), .B(n13735), .Z(n13874) );
  XOR U13799 ( .A(n13876), .B(n13877), .Z(n13714) );
  AND U13800 ( .A(n417), .B(n13867), .Z(n13877) );
  XNOR U13801 ( .A(n13865), .B(n13876), .Z(n13867) );
  XNOR U13802 ( .A(n13878), .B(n13879), .Z(n417) );
  AND U13803 ( .A(n13880), .B(n13881), .Z(n13879) );
  XNOR U13804 ( .A(n13882), .B(n13878), .Z(n13881) );
  IV U13805 ( .A(n13771), .Z(n13882) );
  XNOR U13806 ( .A(n13883), .B(n13884), .Z(n13771) );
  AND U13807 ( .A(n420), .B(n13885), .Z(n13884) );
  XNOR U13808 ( .A(n13883), .B(n13886), .Z(n13885) );
  XNOR U13809 ( .A(n13725), .B(n13878), .Z(n13880) );
  XOR U13810 ( .A(n13887), .B(n13888), .Z(n13725) );
  AND U13811 ( .A(n428), .B(n13889), .Z(n13888) );
  XOR U13812 ( .A(n13872), .B(n13890), .Z(n13878) );
  AND U13813 ( .A(n13891), .B(n13875), .Z(n13890) );
  XNOR U13814 ( .A(n13784), .B(n13872), .Z(n13875) );
  XNOR U13815 ( .A(n13892), .B(n13893), .Z(n13784) );
  AND U13816 ( .A(n420), .B(n13894), .Z(n13893) );
  XOR U13817 ( .A(n13895), .B(n13892), .Z(n13894) );
  XNOR U13818 ( .A(n13896), .B(n13872), .Z(n13891) );
  IV U13819 ( .A(n13735), .Z(n13896) );
  XOR U13820 ( .A(n13897), .B(n13898), .Z(n13735) );
  AND U13821 ( .A(n428), .B(n13899), .Z(n13898) );
  XOR U13822 ( .A(n13900), .B(n13901), .Z(n13872) );
  AND U13823 ( .A(n13902), .B(n13903), .Z(n13901) );
  XNOR U13824 ( .A(n13809), .B(n13900), .Z(n13903) );
  XNOR U13825 ( .A(n13904), .B(n13905), .Z(n13809) );
  AND U13826 ( .A(n420), .B(n13906), .Z(n13905) );
  XNOR U13827 ( .A(n13907), .B(n13904), .Z(n13906) );
  XOR U13828 ( .A(n13900), .B(n13746), .Z(n13902) );
  XOR U13829 ( .A(n13908), .B(n13909), .Z(n13746) );
  AND U13830 ( .A(n428), .B(n13910), .Z(n13909) );
  XOR U13831 ( .A(n13911), .B(n13912), .Z(n13900) );
  AND U13832 ( .A(n13913), .B(n13914), .Z(n13912) );
  XNOR U13833 ( .A(n13911), .B(n13855), .Z(n13914) );
  XNOR U13834 ( .A(n13915), .B(n13916), .Z(n13855) );
  AND U13835 ( .A(n420), .B(n13917), .Z(n13916) );
  XOR U13836 ( .A(n13918), .B(n13915), .Z(n13917) );
  XNOR U13837 ( .A(n13919), .B(n13911), .Z(n13913) );
  IV U13838 ( .A(n13758), .Z(n13919) );
  XOR U13839 ( .A(n13920), .B(n13921), .Z(n13758) );
  AND U13840 ( .A(n428), .B(n13922), .Z(n13921) );
  AND U13841 ( .A(n13876), .B(n13865), .Z(n13911) );
  XNOR U13842 ( .A(n13923), .B(n13924), .Z(n13865) );
  AND U13843 ( .A(n420), .B(n13925), .Z(n13924) );
  XNOR U13844 ( .A(n13926), .B(n13923), .Z(n13925) );
  XNOR U13845 ( .A(n13927), .B(n13928), .Z(n420) );
  AND U13846 ( .A(n13929), .B(n13930), .Z(n13928) );
  XOR U13847 ( .A(n13886), .B(n13927), .Z(n13930) );
  AND U13848 ( .A(n13931), .B(n13932), .Z(n13886) );
  XOR U13849 ( .A(n13927), .B(n13883), .Z(n13929) );
  XNOR U13850 ( .A(n13933), .B(n13934), .Z(n13883) );
  AND U13851 ( .A(n424), .B(n13889), .Z(n13934) );
  XOR U13852 ( .A(n13887), .B(n13933), .Z(n13889) );
  XOR U13853 ( .A(n13935), .B(n13936), .Z(n13927) );
  AND U13854 ( .A(n13937), .B(n13938), .Z(n13936) );
  XNOR U13855 ( .A(n13935), .B(n13931), .Z(n13938) );
  IV U13856 ( .A(n13895), .Z(n13931) );
  XOR U13857 ( .A(n13939), .B(n13940), .Z(n13895) );
  XOR U13858 ( .A(n13941), .B(n13932), .Z(n13940) );
  AND U13859 ( .A(n13907), .B(n13942), .Z(n13932) );
  AND U13860 ( .A(n13943), .B(n13944), .Z(n13941) );
  XOR U13861 ( .A(n13945), .B(n13939), .Z(n13943) );
  XNOR U13862 ( .A(n13892), .B(n13935), .Z(n13937) );
  XNOR U13863 ( .A(n13946), .B(n13947), .Z(n13892) );
  AND U13864 ( .A(n424), .B(n13899), .Z(n13947) );
  XOR U13865 ( .A(n13946), .B(n13897), .Z(n13899) );
  XOR U13866 ( .A(n13948), .B(n13949), .Z(n13935) );
  AND U13867 ( .A(n13950), .B(n13951), .Z(n13949) );
  XNOR U13868 ( .A(n13948), .B(n13907), .Z(n13951) );
  XOR U13869 ( .A(n13952), .B(n13944), .Z(n13907) );
  XNOR U13870 ( .A(n13953), .B(n13939), .Z(n13944) );
  XOR U13871 ( .A(n13954), .B(n13955), .Z(n13939) );
  AND U13872 ( .A(n13956), .B(n13957), .Z(n13955) );
  XOR U13873 ( .A(n13958), .B(n13954), .Z(n13956) );
  XNOR U13874 ( .A(n13959), .B(n13960), .Z(n13953) );
  AND U13875 ( .A(n13961), .B(n13962), .Z(n13960) );
  XOR U13876 ( .A(n13959), .B(n13963), .Z(n13961) );
  XNOR U13877 ( .A(n13945), .B(n13942), .Z(n13952) );
  AND U13878 ( .A(n13964), .B(n13965), .Z(n13942) );
  XOR U13879 ( .A(n13966), .B(n13967), .Z(n13945) );
  AND U13880 ( .A(n13968), .B(n13969), .Z(n13967) );
  XOR U13881 ( .A(n13966), .B(n13970), .Z(n13968) );
  XNOR U13882 ( .A(n13904), .B(n13948), .Z(n13950) );
  XNOR U13883 ( .A(n13971), .B(n13972), .Z(n13904) );
  AND U13884 ( .A(n424), .B(n13910), .Z(n13972) );
  XOR U13885 ( .A(n13971), .B(n13908), .Z(n13910) );
  XOR U13886 ( .A(n13973), .B(n13974), .Z(n13948) );
  AND U13887 ( .A(n13975), .B(n13976), .Z(n13974) );
  XNOR U13888 ( .A(n13973), .B(n13964), .Z(n13976) );
  IV U13889 ( .A(n13918), .Z(n13964) );
  XNOR U13890 ( .A(n13977), .B(n13957), .Z(n13918) );
  XNOR U13891 ( .A(n13978), .B(n13963), .Z(n13957) );
  XOR U13892 ( .A(n13979), .B(n13980), .Z(n13963) );
  NOR U13893 ( .A(n13981), .B(n13982), .Z(n13980) );
  XNOR U13894 ( .A(n13979), .B(n13983), .Z(n13981) );
  XNOR U13895 ( .A(n13962), .B(n13954), .Z(n13978) );
  XOR U13896 ( .A(n13984), .B(n13985), .Z(n13954) );
  AND U13897 ( .A(n13986), .B(n13987), .Z(n13985) );
  XNOR U13898 ( .A(n13984), .B(n13988), .Z(n13986) );
  XNOR U13899 ( .A(n13989), .B(n13959), .Z(n13962) );
  XOR U13900 ( .A(n13990), .B(n13991), .Z(n13959) );
  AND U13901 ( .A(n13992), .B(n13993), .Z(n13991) );
  XOR U13902 ( .A(n13990), .B(n13994), .Z(n13992) );
  XNOR U13903 ( .A(n13995), .B(n13996), .Z(n13989) );
  NOR U13904 ( .A(n13997), .B(n13998), .Z(n13996) );
  XOR U13905 ( .A(n13995), .B(n13999), .Z(n13997) );
  XNOR U13906 ( .A(n13958), .B(n13965), .Z(n13977) );
  NOR U13907 ( .A(n13926), .B(n14000), .Z(n13965) );
  XOR U13908 ( .A(n13970), .B(n13969), .Z(n13958) );
  XNOR U13909 ( .A(n14001), .B(n13966), .Z(n13969) );
  XOR U13910 ( .A(n14002), .B(n14003), .Z(n13966) );
  AND U13911 ( .A(n14004), .B(n14005), .Z(n14003) );
  XOR U13912 ( .A(n14002), .B(n14006), .Z(n14004) );
  XNOR U13913 ( .A(n14007), .B(n14008), .Z(n14001) );
  NOR U13914 ( .A(n14009), .B(n14010), .Z(n14008) );
  XNOR U13915 ( .A(n14007), .B(n14011), .Z(n14009) );
  XOR U13916 ( .A(n14012), .B(n14013), .Z(n13970) );
  NOR U13917 ( .A(n14014), .B(n14015), .Z(n14013) );
  XNOR U13918 ( .A(n14012), .B(n14016), .Z(n14014) );
  XNOR U13919 ( .A(n13915), .B(n13973), .Z(n13975) );
  XNOR U13920 ( .A(n14017), .B(n14018), .Z(n13915) );
  AND U13921 ( .A(n424), .B(n13922), .Z(n14018) );
  XOR U13922 ( .A(n14017), .B(n13920), .Z(n13922) );
  AND U13923 ( .A(n13923), .B(n13926), .Z(n13973) );
  XOR U13924 ( .A(n14019), .B(n14000), .Z(n13926) );
  XNOR U13925 ( .A(p_input[1024]), .B(p_input[560]), .Z(n14000) );
  XOR U13926 ( .A(n13988), .B(n13987), .Z(n14019) );
  XNOR U13927 ( .A(n14020), .B(n13994), .Z(n13987) );
  XNOR U13928 ( .A(n13983), .B(n13982), .Z(n13994) );
  XOR U13929 ( .A(n14021), .B(n13979), .Z(n13982) );
  XOR U13930 ( .A(p_input[1034]), .B(p_input[570]), .Z(n13979) );
  XNOR U13931 ( .A(p_input[1035]), .B(p_input[571]), .Z(n14021) );
  XOR U13932 ( .A(p_input[1036]), .B(p_input[572]), .Z(n13983) );
  XNOR U13933 ( .A(n13993), .B(n13984), .Z(n14020) );
  XOR U13934 ( .A(p_input[1025]), .B(p_input[561]), .Z(n13984) );
  XOR U13935 ( .A(n14022), .B(n13999), .Z(n13993) );
  XNOR U13936 ( .A(p_input[1039]), .B(p_input[575]), .Z(n13999) );
  XOR U13937 ( .A(n13990), .B(n13998), .Z(n14022) );
  XOR U13938 ( .A(n14023), .B(n13995), .Z(n13998) );
  XOR U13939 ( .A(p_input[1037]), .B(p_input[573]), .Z(n13995) );
  XNOR U13940 ( .A(p_input[1038]), .B(p_input[574]), .Z(n14023) );
  XOR U13941 ( .A(p_input[1033]), .B(p_input[569]), .Z(n13990) );
  XNOR U13942 ( .A(n14006), .B(n14005), .Z(n13988) );
  XNOR U13943 ( .A(n14024), .B(n14011), .Z(n14005) );
  XOR U13944 ( .A(p_input[1032]), .B(p_input[568]), .Z(n14011) );
  XOR U13945 ( .A(n14002), .B(n14010), .Z(n14024) );
  XOR U13946 ( .A(n14025), .B(n14007), .Z(n14010) );
  XOR U13947 ( .A(p_input[1030]), .B(p_input[566]), .Z(n14007) );
  XNOR U13948 ( .A(p_input[1031]), .B(p_input[567]), .Z(n14025) );
  XOR U13949 ( .A(p_input[1026]), .B(p_input[562]), .Z(n14002) );
  XNOR U13950 ( .A(n14016), .B(n14015), .Z(n14006) );
  XOR U13951 ( .A(n14026), .B(n14012), .Z(n14015) );
  XOR U13952 ( .A(p_input[1027]), .B(p_input[563]), .Z(n14012) );
  XNOR U13953 ( .A(p_input[1028]), .B(p_input[564]), .Z(n14026) );
  XOR U13954 ( .A(p_input[1029]), .B(p_input[565]), .Z(n14016) );
  XNOR U13955 ( .A(n14027), .B(n14028), .Z(n13923) );
  AND U13956 ( .A(n424), .B(n14029), .Z(n14028) );
  XNOR U13957 ( .A(n14030), .B(n14031), .Z(n424) );
  AND U13958 ( .A(n14032), .B(n14033), .Z(n14031) );
  XOR U13959 ( .A(n14030), .B(n13933), .Z(n14033) );
  XNOR U13960 ( .A(n14030), .B(n13887), .Z(n14032) );
  XOR U13961 ( .A(n14034), .B(n14035), .Z(n14030) );
  AND U13962 ( .A(n14036), .B(n14037), .Z(n14035) );
  XOR U13963 ( .A(n14034), .B(n13897), .Z(n14036) );
  XOR U13964 ( .A(n14038), .B(n14039), .Z(n13876) );
  AND U13965 ( .A(n428), .B(n14029), .Z(n14039) );
  XNOR U13966 ( .A(n14027), .B(n14038), .Z(n14029) );
  XNOR U13967 ( .A(n14040), .B(n14041), .Z(n428) );
  AND U13968 ( .A(n14042), .B(n14043), .Z(n14041) );
  XNOR U13969 ( .A(n14044), .B(n14040), .Z(n14043) );
  IV U13970 ( .A(n13933), .Z(n14044) );
  XNOR U13971 ( .A(n14045), .B(n14046), .Z(n13933) );
  AND U13972 ( .A(n431), .B(n14047), .Z(n14046) );
  XNOR U13973 ( .A(n14045), .B(n14048), .Z(n14047) );
  XNOR U13974 ( .A(n13887), .B(n14040), .Z(n14042) );
  XOR U13975 ( .A(n14049), .B(n14050), .Z(n13887) );
  AND U13976 ( .A(n439), .B(n14051), .Z(n14050) );
  XOR U13977 ( .A(n14034), .B(n14052), .Z(n14040) );
  AND U13978 ( .A(n14053), .B(n14037), .Z(n14052) );
  XNOR U13979 ( .A(n13946), .B(n14034), .Z(n14037) );
  XNOR U13980 ( .A(n14054), .B(n14055), .Z(n13946) );
  AND U13981 ( .A(n431), .B(n14056), .Z(n14055) );
  XOR U13982 ( .A(n14057), .B(n14054), .Z(n14056) );
  XNOR U13983 ( .A(n14058), .B(n14034), .Z(n14053) );
  IV U13984 ( .A(n13897), .Z(n14058) );
  XOR U13985 ( .A(n14059), .B(n14060), .Z(n13897) );
  AND U13986 ( .A(n439), .B(n14061), .Z(n14060) );
  XOR U13987 ( .A(n14062), .B(n14063), .Z(n14034) );
  AND U13988 ( .A(n14064), .B(n14065), .Z(n14063) );
  XNOR U13989 ( .A(n13971), .B(n14062), .Z(n14065) );
  XNOR U13990 ( .A(n14066), .B(n14067), .Z(n13971) );
  AND U13991 ( .A(n431), .B(n14068), .Z(n14067) );
  XNOR U13992 ( .A(n14069), .B(n14066), .Z(n14068) );
  XOR U13993 ( .A(n14062), .B(n13908), .Z(n14064) );
  XOR U13994 ( .A(n14070), .B(n14071), .Z(n13908) );
  AND U13995 ( .A(n439), .B(n14072), .Z(n14071) );
  XOR U13996 ( .A(n14073), .B(n14074), .Z(n14062) );
  AND U13997 ( .A(n14075), .B(n14076), .Z(n14074) );
  XNOR U13998 ( .A(n14073), .B(n14017), .Z(n14076) );
  XNOR U13999 ( .A(n14077), .B(n14078), .Z(n14017) );
  AND U14000 ( .A(n431), .B(n14079), .Z(n14078) );
  XOR U14001 ( .A(n14080), .B(n14077), .Z(n14079) );
  XNOR U14002 ( .A(n14081), .B(n14073), .Z(n14075) );
  IV U14003 ( .A(n13920), .Z(n14081) );
  XOR U14004 ( .A(n14082), .B(n14083), .Z(n13920) );
  AND U14005 ( .A(n439), .B(n14084), .Z(n14083) );
  AND U14006 ( .A(n14038), .B(n14027), .Z(n14073) );
  XNOR U14007 ( .A(n14085), .B(n14086), .Z(n14027) );
  AND U14008 ( .A(n431), .B(n14087), .Z(n14086) );
  XNOR U14009 ( .A(n14088), .B(n14085), .Z(n14087) );
  XNOR U14010 ( .A(n14089), .B(n14090), .Z(n431) );
  AND U14011 ( .A(n14091), .B(n14092), .Z(n14090) );
  XOR U14012 ( .A(n14048), .B(n14089), .Z(n14092) );
  AND U14013 ( .A(n14093), .B(n14094), .Z(n14048) );
  XOR U14014 ( .A(n14089), .B(n14045), .Z(n14091) );
  XNOR U14015 ( .A(n14095), .B(n14096), .Z(n14045) );
  AND U14016 ( .A(n435), .B(n14051), .Z(n14096) );
  XOR U14017 ( .A(n14049), .B(n14095), .Z(n14051) );
  XOR U14018 ( .A(n14097), .B(n14098), .Z(n14089) );
  AND U14019 ( .A(n14099), .B(n14100), .Z(n14098) );
  XNOR U14020 ( .A(n14097), .B(n14093), .Z(n14100) );
  IV U14021 ( .A(n14057), .Z(n14093) );
  XOR U14022 ( .A(n14101), .B(n14102), .Z(n14057) );
  XOR U14023 ( .A(n14103), .B(n14094), .Z(n14102) );
  AND U14024 ( .A(n14069), .B(n14104), .Z(n14094) );
  AND U14025 ( .A(n14105), .B(n14106), .Z(n14103) );
  XOR U14026 ( .A(n14107), .B(n14101), .Z(n14105) );
  XNOR U14027 ( .A(n14054), .B(n14097), .Z(n14099) );
  XNOR U14028 ( .A(n14108), .B(n14109), .Z(n14054) );
  AND U14029 ( .A(n435), .B(n14061), .Z(n14109) );
  XOR U14030 ( .A(n14108), .B(n14059), .Z(n14061) );
  XOR U14031 ( .A(n14110), .B(n14111), .Z(n14097) );
  AND U14032 ( .A(n14112), .B(n14113), .Z(n14111) );
  XNOR U14033 ( .A(n14110), .B(n14069), .Z(n14113) );
  XOR U14034 ( .A(n14114), .B(n14106), .Z(n14069) );
  XNOR U14035 ( .A(n14115), .B(n14101), .Z(n14106) );
  XOR U14036 ( .A(n14116), .B(n14117), .Z(n14101) );
  AND U14037 ( .A(n14118), .B(n14119), .Z(n14117) );
  XOR U14038 ( .A(n14120), .B(n14116), .Z(n14118) );
  XNOR U14039 ( .A(n14121), .B(n14122), .Z(n14115) );
  AND U14040 ( .A(n14123), .B(n14124), .Z(n14122) );
  XOR U14041 ( .A(n14121), .B(n14125), .Z(n14123) );
  XNOR U14042 ( .A(n14107), .B(n14104), .Z(n14114) );
  AND U14043 ( .A(n14126), .B(n14127), .Z(n14104) );
  XOR U14044 ( .A(n14128), .B(n14129), .Z(n14107) );
  AND U14045 ( .A(n14130), .B(n14131), .Z(n14129) );
  XOR U14046 ( .A(n14128), .B(n14132), .Z(n14130) );
  XNOR U14047 ( .A(n14066), .B(n14110), .Z(n14112) );
  XNOR U14048 ( .A(n14133), .B(n14134), .Z(n14066) );
  AND U14049 ( .A(n435), .B(n14072), .Z(n14134) );
  XOR U14050 ( .A(n14133), .B(n14070), .Z(n14072) );
  XOR U14051 ( .A(n14135), .B(n14136), .Z(n14110) );
  AND U14052 ( .A(n14137), .B(n14138), .Z(n14136) );
  XNOR U14053 ( .A(n14135), .B(n14126), .Z(n14138) );
  IV U14054 ( .A(n14080), .Z(n14126) );
  XNOR U14055 ( .A(n14139), .B(n14119), .Z(n14080) );
  XNOR U14056 ( .A(n14140), .B(n14125), .Z(n14119) );
  XOR U14057 ( .A(n14141), .B(n14142), .Z(n14125) );
  NOR U14058 ( .A(n14143), .B(n14144), .Z(n14142) );
  XNOR U14059 ( .A(n14141), .B(n14145), .Z(n14143) );
  XNOR U14060 ( .A(n14124), .B(n14116), .Z(n14140) );
  XOR U14061 ( .A(n14146), .B(n14147), .Z(n14116) );
  AND U14062 ( .A(n14148), .B(n14149), .Z(n14147) );
  XNOR U14063 ( .A(n14146), .B(n14150), .Z(n14148) );
  XNOR U14064 ( .A(n14151), .B(n14121), .Z(n14124) );
  XOR U14065 ( .A(n14152), .B(n14153), .Z(n14121) );
  AND U14066 ( .A(n14154), .B(n14155), .Z(n14153) );
  XOR U14067 ( .A(n14152), .B(n14156), .Z(n14154) );
  XNOR U14068 ( .A(n14157), .B(n14158), .Z(n14151) );
  NOR U14069 ( .A(n14159), .B(n14160), .Z(n14158) );
  XOR U14070 ( .A(n14157), .B(n14161), .Z(n14159) );
  XNOR U14071 ( .A(n14120), .B(n14127), .Z(n14139) );
  NOR U14072 ( .A(n14088), .B(n14162), .Z(n14127) );
  XOR U14073 ( .A(n14132), .B(n14131), .Z(n14120) );
  XNOR U14074 ( .A(n14163), .B(n14128), .Z(n14131) );
  XOR U14075 ( .A(n14164), .B(n14165), .Z(n14128) );
  AND U14076 ( .A(n14166), .B(n14167), .Z(n14165) );
  XOR U14077 ( .A(n14164), .B(n14168), .Z(n14166) );
  XNOR U14078 ( .A(n14169), .B(n14170), .Z(n14163) );
  NOR U14079 ( .A(n14171), .B(n14172), .Z(n14170) );
  XNOR U14080 ( .A(n14169), .B(n14173), .Z(n14171) );
  XOR U14081 ( .A(n14174), .B(n14175), .Z(n14132) );
  NOR U14082 ( .A(n14176), .B(n14177), .Z(n14175) );
  XNOR U14083 ( .A(n14174), .B(n14178), .Z(n14176) );
  XNOR U14084 ( .A(n14077), .B(n14135), .Z(n14137) );
  XNOR U14085 ( .A(n14179), .B(n14180), .Z(n14077) );
  AND U14086 ( .A(n435), .B(n14084), .Z(n14180) );
  XOR U14087 ( .A(n14179), .B(n14082), .Z(n14084) );
  AND U14088 ( .A(n14085), .B(n14088), .Z(n14135) );
  XOR U14089 ( .A(n14181), .B(n14162), .Z(n14088) );
  XNOR U14090 ( .A(p_input[1024]), .B(p_input[576]), .Z(n14162) );
  XOR U14091 ( .A(n14150), .B(n14149), .Z(n14181) );
  XNOR U14092 ( .A(n14182), .B(n14156), .Z(n14149) );
  XNOR U14093 ( .A(n14145), .B(n14144), .Z(n14156) );
  XOR U14094 ( .A(n14183), .B(n14141), .Z(n14144) );
  XOR U14095 ( .A(p_input[1034]), .B(p_input[586]), .Z(n14141) );
  XNOR U14096 ( .A(p_input[1035]), .B(p_input[587]), .Z(n14183) );
  XOR U14097 ( .A(p_input[1036]), .B(p_input[588]), .Z(n14145) );
  XNOR U14098 ( .A(n14155), .B(n14146), .Z(n14182) );
  XOR U14099 ( .A(p_input[1025]), .B(p_input[577]), .Z(n14146) );
  XOR U14100 ( .A(n14184), .B(n14161), .Z(n14155) );
  XNOR U14101 ( .A(p_input[1039]), .B(p_input[591]), .Z(n14161) );
  XOR U14102 ( .A(n14152), .B(n14160), .Z(n14184) );
  XOR U14103 ( .A(n14185), .B(n14157), .Z(n14160) );
  XOR U14104 ( .A(p_input[1037]), .B(p_input[589]), .Z(n14157) );
  XNOR U14105 ( .A(p_input[1038]), .B(p_input[590]), .Z(n14185) );
  XOR U14106 ( .A(p_input[1033]), .B(p_input[585]), .Z(n14152) );
  XNOR U14107 ( .A(n14168), .B(n14167), .Z(n14150) );
  XNOR U14108 ( .A(n14186), .B(n14173), .Z(n14167) );
  XOR U14109 ( .A(p_input[1032]), .B(p_input[584]), .Z(n14173) );
  XOR U14110 ( .A(n14164), .B(n14172), .Z(n14186) );
  XOR U14111 ( .A(n14187), .B(n14169), .Z(n14172) );
  XOR U14112 ( .A(p_input[1030]), .B(p_input[582]), .Z(n14169) );
  XNOR U14113 ( .A(p_input[1031]), .B(p_input[583]), .Z(n14187) );
  XOR U14114 ( .A(p_input[1026]), .B(p_input[578]), .Z(n14164) );
  XNOR U14115 ( .A(n14178), .B(n14177), .Z(n14168) );
  XOR U14116 ( .A(n14188), .B(n14174), .Z(n14177) );
  XOR U14117 ( .A(p_input[1027]), .B(p_input[579]), .Z(n14174) );
  XNOR U14118 ( .A(p_input[1028]), .B(p_input[580]), .Z(n14188) );
  XOR U14119 ( .A(p_input[1029]), .B(p_input[581]), .Z(n14178) );
  XNOR U14120 ( .A(n14189), .B(n14190), .Z(n14085) );
  AND U14121 ( .A(n435), .B(n14191), .Z(n14190) );
  XNOR U14122 ( .A(n14192), .B(n14193), .Z(n435) );
  AND U14123 ( .A(n14194), .B(n14195), .Z(n14193) );
  XOR U14124 ( .A(n14192), .B(n14095), .Z(n14195) );
  XNOR U14125 ( .A(n14192), .B(n14049), .Z(n14194) );
  XOR U14126 ( .A(n14196), .B(n14197), .Z(n14192) );
  AND U14127 ( .A(n14198), .B(n14199), .Z(n14197) );
  XOR U14128 ( .A(n14196), .B(n14059), .Z(n14198) );
  XOR U14129 ( .A(n14200), .B(n14201), .Z(n14038) );
  AND U14130 ( .A(n439), .B(n14191), .Z(n14201) );
  XNOR U14131 ( .A(n14189), .B(n14200), .Z(n14191) );
  XNOR U14132 ( .A(n14202), .B(n14203), .Z(n439) );
  AND U14133 ( .A(n14204), .B(n14205), .Z(n14203) );
  XNOR U14134 ( .A(n14206), .B(n14202), .Z(n14205) );
  IV U14135 ( .A(n14095), .Z(n14206) );
  XNOR U14136 ( .A(n14207), .B(n14208), .Z(n14095) );
  AND U14137 ( .A(n442), .B(n14209), .Z(n14208) );
  XNOR U14138 ( .A(n14207), .B(n14210), .Z(n14209) );
  XNOR U14139 ( .A(n14049), .B(n14202), .Z(n14204) );
  XOR U14140 ( .A(n14211), .B(n14212), .Z(n14049) );
  AND U14141 ( .A(n450), .B(n14213), .Z(n14212) );
  XOR U14142 ( .A(n14196), .B(n14214), .Z(n14202) );
  AND U14143 ( .A(n14215), .B(n14199), .Z(n14214) );
  XNOR U14144 ( .A(n14108), .B(n14196), .Z(n14199) );
  XNOR U14145 ( .A(n14216), .B(n14217), .Z(n14108) );
  AND U14146 ( .A(n442), .B(n14218), .Z(n14217) );
  XOR U14147 ( .A(n14219), .B(n14216), .Z(n14218) );
  XNOR U14148 ( .A(n14220), .B(n14196), .Z(n14215) );
  IV U14149 ( .A(n14059), .Z(n14220) );
  XOR U14150 ( .A(n14221), .B(n14222), .Z(n14059) );
  AND U14151 ( .A(n450), .B(n14223), .Z(n14222) );
  XOR U14152 ( .A(n14224), .B(n14225), .Z(n14196) );
  AND U14153 ( .A(n14226), .B(n14227), .Z(n14225) );
  XNOR U14154 ( .A(n14133), .B(n14224), .Z(n14227) );
  XNOR U14155 ( .A(n14228), .B(n14229), .Z(n14133) );
  AND U14156 ( .A(n442), .B(n14230), .Z(n14229) );
  XNOR U14157 ( .A(n14231), .B(n14228), .Z(n14230) );
  XOR U14158 ( .A(n14224), .B(n14070), .Z(n14226) );
  XOR U14159 ( .A(n14232), .B(n14233), .Z(n14070) );
  AND U14160 ( .A(n450), .B(n14234), .Z(n14233) );
  XOR U14161 ( .A(n14235), .B(n14236), .Z(n14224) );
  AND U14162 ( .A(n14237), .B(n14238), .Z(n14236) );
  XNOR U14163 ( .A(n14235), .B(n14179), .Z(n14238) );
  XNOR U14164 ( .A(n14239), .B(n14240), .Z(n14179) );
  AND U14165 ( .A(n442), .B(n14241), .Z(n14240) );
  XOR U14166 ( .A(n14242), .B(n14239), .Z(n14241) );
  XNOR U14167 ( .A(n14243), .B(n14235), .Z(n14237) );
  IV U14168 ( .A(n14082), .Z(n14243) );
  XOR U14169 ( .A(n14244), .B(n14245), .Z(n14082) );
  AND U14170 ( .A(n450), .B(n14246), .Z(n14245) );
  AND U14171 ( .A(n14200), .B(n14189), .Z(n14235) );
  XNOR U14172 ( .A(n14247), .B(n14248), .Z(n14189) );
  AND U14173 ( .A(n442), .B(n14249), .Z(n14248) );
  XNOR U14174 ( .A(n14250), .B(n14247), .Z(n14249) );
  XNOR U14175 ( .A(n14251), .B(n14252), .Z(n442) );
  AND U14176 ( .A(n14253), .B(n14254), .Z(n14252) );
  XOR U14177 ( .A(n14210), .B(n14251), .Z(n14254) );
  AND U14178 ( .A(n14255), .B(n14256), .Z(n14210) );
  XOR U14179 ( .A(n14251), .B(n14207), .Z(n14253) );
  XNOR U14180 ( .A(n14257), .B(n14258), .Z(n14207) );
  AND U14181 ( .A(n446), .B(n14213), .Z(n14258) );
  XOR U14182 ( .A(n14211), .B(n14257), .Z(n14213) );
  XOR U14183 ( .A(n14259), .B(n14260), .Z(n14251) );
  AND U14184 ( .A(n14261), .B(n14262), .Z(n14260) );
  XNOR U14185 ( .A(n14259), .B(n14255), .Z(n14262) );
  IV U14186 ( .A(n14219), .Z(n14255) );
  XOR U14187 ( .A(n14263), .B(n14264), .Z(n14219) );
  XOR U14188 ( .A(n14265), .B(n14256), .Z(n14264) );
  AND U14189 ( .A(n14231), .B(n14266), .Z(n14256) );
  AND U14190 ( .A(n14267), .B(n14268), .Z(n14265) );
  XOR U14191 ( .A(n14269), .B(n14263), .Z(n14267) );
  XNOR U14192 ( .A(n14216), .B(n14259), .Z(n14261) );
  XNOR U14193 ( .A(n14270), .B(n14271), .Z(n14216) );
  AND U14194 ( .A(n446), .B(n14223), .Z(n14271) );
  XOR U14195 ( .A(n14270), .B(n14221), .Z(n14223) );
  XOR U14196 ( .A(n14272), .B(n14273), .Z(n14259) );
  AND U14197 ( .A(n14274), .B(n14275), .Z(n14273) );
  XNOR U14198 ( .A(n14272), .B(n14231), .Z(n14275) );
  XOR U14199 ( .A(n14276), .B(n14268), .Z(n14231) );
  XNOR U14200 ( .A(n14277), .B(n14263), .Z(n14268) );
  XOR U14201 ( .A(n14278), .B(n14279), .Z(n14263) );
  AND U14202 ( .A(n14280), .B(n14281), .Z(n14279) );
  XOR U14203 ( .A(n14282), .B(n14278), .Z(n14280) );
  XNOR U14204 ( .A(n14283), .B(n14284), .Z(n14277) );
  AND U14205 ( .A(n14285), .B(n14286), .Z(n14284) );
  XOR U14206 ( .A(n14283), .B(n14287), .Z(n14285) );
  XNOR U14207 ( .A(n14269), .B(n14266), .Z(n14276) );
  AND U14208 ( .A(n14288), .B(n14289), .Z(n14266) );
  XOR U14209 ( .A(n14290), .B(n14291), .Z(n14269) );
  AND U14210 ( .A(n14292), .B(n14293), .Z(n14291) );
  XOR U14211 ( .A(n14290), .B(n14294), .Z(n14292) );
  XNOR U14212 ( .A(n14228), .B(n14272), .Z(n14274) );
  XNOR U14213 ( .A(n14295), .B(n14296), .Z(n14228) );
  AND U14214 ( .A(n446), .B(n14234), .Z(n14296) );
  XOR U14215 ( .A(n14295), .B(n14232), .Z(n14234) );
  XOR U14216 ( .A(n14297), .B(n14298), .Z(n14272) );
  AND U14217 ( .A(n14299), .B(n14300), .Z(n14298) );
  XNOR U14218 ( .A(n14297), .B(n14288), .Z(n14300) );
  IV U14219 ( .A(n14242), .Z(n14288) );
  XNOR U14220 ( .A(n14301), .B(n14281), .Z(n14242) );
  XNOR U14221 ( .A(n14302), .B(n14287), .Z(n14281) );
  XOR U14222 ( .A(n14303), .B(n14304), .Z(n14287) );
  NOR U14223 ( .A(n14305), .B(n14306), .Z(n14304) );
  XNOR U14224 ( .A(n14303), .B(n14307), .Z(n14305) );
  XNOR U14225 ( .A(n14286), .B(n14278), .Z(n14302) );
  XOR U14226 ( .A(n14308), .B(n14309), .Z(n14278) );
  AND U14227 ( .A(n14310), .B(n14311), .Z(n14309) );
  XNOR U14228 ( .A(n14308), .B(n14312), .Z(n14310) );
  XNOR U14229 ( .A(n14313), .B(n14283), .Z(n14286) );
  XOR U14230 ( .A(n14314), .B(n14315), .Z(n14283) );
  AND U14231 ( .A(n14316), .B(n14317), .Z(n14315) );
  XOR U14232 ( .A(n14314), .B(n14318), .Z(n14316) );
  XNOR U14233 ( .A(n14319), .B(n14320), .Z(n14313) );
  NOR U14234 ( .A(n14321), .B(n14322), .Z(n14320) );
  XOR U14235 ( .A(n14319), .B(n14323), .Z(n14321) );
  XNOR U14236 ( .A(n14282), .B(n14289), .Z(n14301) );
  NOR U14237 ( .A(n14250), .B(n14324), .Z(n14289) );
  XOR U14238 ( .A(n14294), .B(n14293), .Z(n14282) );
  XNOR U14239 ( .A(n14325), .B(n14290), .Z(n14293) );
  XOR U14240 ( .A(n14326), .B(n14327), .Z(n14290) );
  AND U14241 ( .A(n14328), .B(n14329), .Z(n14327) );
  XOR U14242 ( .A(n14326), .B(n14330), .Z(n14328) );
  XNOR U14243 ( .A(n14331), .B(n14332), .Z(n14325) );
  NOR U14244 ( .A(n14333), .B(n14334), .Z(n14332) );
  XNOR U14245 ( .A(n14331), .B(n14335), .Z(n14333) );
  XOR U14246 ( .A(n14336), .B(n14337), .Z(n14294) );
  NOR U14247 ( .A(n14338), .B(n14339), .Z(n14337) );
  XNOR U14248 ( .A(n14336), .B(n14340), .Z(n14338) );
  XNOR U14249 ( .A(n14239), .B(n14297), .Z(n14299) );
  XNOR U14250 ( .A(n14341), .B(n14342), .Z(n14239) );
  AND U14251 ( .A(n446), .B(n14246), .Z(n14342) );
  XOR U14252 ( .A(n14341), .B(n14244), .Z(n14246) );
  AND U14253 ( .A(n14247), .B(n14250), .Z(n14297) );
  XOR U14254 ( .A(n14343), .B(n14324), .Z(n14250) );
  XNOR U14255 ( .A(p_input[1024]), .B(p_input[592]), .Z(n14324) );
  XOR U14256 ( .A(n14312), .B(n14311), .Z(n14343) );
  XNOR U14257 ( .A(n14344), .B(n14318), .Z(n14311) );
  XNOR U14258 ( .A(n14307), .B(n14306), .Z(n14318) );
  XOR U14259 ( .A(n14345), .B(n14303), .Z(n14306) );
  XOR U14260 ( .A(p_input[1034]), .B(p_input[602]), .Z(n14303) );
  XNOR U14261 ( .A(p_input[1035]), .B(p_input[603]), .Z(n14345) );
  XOR U14262 ( .A(p_input[1036]), .B(p_input[604]), .Z(n14307) );
  XNOR U14263 ( .A(n14317), .B(n14308), .Z(n14344) );
  XOR U14264 ( .A(p_input[1025]), .B(p_input[593]), .Z(n14308) );
  XOR U14265 ( .A(n14346), .B(n14323), .Z(n14317) );
  XNOR U14266 ( .A(p_input[1039]), .B(p_input[607]), .Z(n14323) );
  XOR U14267 ( .A(n14314), .B(n14322), .Z(n14346) );
  XOR U14268 ( .A(n14347), .B(n14319), .Z(n14322) );
  XOR U14269 ( .A(p_input[1037]), .B(p_input[605]), .Z(n14319) );
  XNOR U14270 ( .A(p_input[1038]), .B(p_input[606]), .Z(n14347) );
  XOR U14271 ( .A(p_input[1033]), .B(p_input[601]), .Z(n14314) );
  XNOR U14272 ( .A(n14330), .B(n14329), .Z(n14312) );
  XNOR U14273 ( .A(n14348), .B(n14335), .Z(n14329) );
  XOR U14274 ( .A(p_input[1032]), .B(p_input[600]), .Z(n14335) );
  XOR U14275 ( .A(n14326), .B(n14334), .Z(n14348) );
  XOR U14276 ( .A(n14349), .B(n14331), .Z(n14334) );
  XOR U14277 ( .A(p_input[1030]), .B(p_input[598]), .Z(n14331) );
  XNOR U14278 ( .A(p_input[1031]), .B(p_input[599]), .Z(n14349) );
  XOR U14279 ( .A(p_input[1026]), .B(p_input[594]), .Z(n14326) );
  XNOR U14280 ( .A(n14340), .B(n14339), .Z(n14330) );
  XOR U14281 ( .A(n14350), .B(n14336), .Z(n14339) );
  XOR U14282 ( .A(p_input[1027]), .B(p_input[595]), .Z(n14336) );
  XNOR U14283 ( .A(p_input[1028]), .B(p_input[596]), .Z(n14350) );
  XOR U14284 ( .A(p_input[1029]), .B(p_input[597]), .Z(n14340) );
  XNOR U14285 ( .A(n14351), .B(n14352), .Z(n14247) );
  AND U14286 ( .A(n446), .B(n14353), .Z(n14352) );
  XNOR U14287 ( .A(n14354), .B(n14355), .Z(n446) );
  AND U14288 ( .A(n14356), .B(n14357), .Z(n14355) );
  XOR U14289 ( .A(n14354), .B(n14257), .Z(n14357) );
  XNOR U14290 ( .A(n14354), .B(n14211), .Z(n14356) );
  XOR U14291 ( .A(n14358), .B(n14359), .Z(n14354) );
  AND U14292 ( .A(n14360), .B(n14361), .Z(n14359) );
  XOR U14293 ( .A(n14358), .B(n14221), .Z(n14360) );
  XOR U14294 ( .A(n14362), .B(n14363), .Z(n14200) );
  AND U14295 ( .A(n450), .B(n14353), .Z(n14363) );
  XNOR U14296 ( .A(n14351), .B(n14362), .Z(n14353) );
  XNOR U14297 ( .A(n14364), .B(n14365), .Z(n450) );
  AND U14298 ( .A(n14366), .B(n14367), .Z(n14365) );
  XNOR U14299 ( .A(n14368), .B(n14364), .Z(n14367) );
  IV U14300 ( .A(n14257), .Z(n14368) );
  XNOR U14301 ( .A(n14369), .B(n14370), .Z(n14257) );
  AND U14302 ( .A(n453), .B(n14371), .Z(n14370) );
  XNOR U14303 ( .A(n14369), .B(n14372), .Z(n14371) );
  XNOR U14304 ( .A(n14211), .B(n14364), .Z(n14366) );
  XOR U14305 ( .A(n14373), .B(n14374), .Z(n14211) );
  AND U14306 ( .A(n461), .B(n14375), .Z(n14374) );
  XOR U14307 ( .A(n14358), .B(n14376), .Z(n14364) );
  AND U14308 ( .A(n14377), .B(n14361), .Z(n14376) );
  XNOR U14309 ( .A(n14270), .B(n14358), .Z(n14361) );
  XNOR U14310 ( .A(n14378), .B(n14379), .Z(n14270) );
  AND U14311 ( .A(n453), .B(n14380), .Z(n14379) );
  XOR U14312 ( .A(n14381), .B(n14378), .Z(n14380) );
  XNOR U14313 ( .A(n14382), .B(n14358), .Z(n14377) );
  IV U14314 ( .A(n14221), .Z(n14382) );
  XOR U14315 ( .A(n14383), .B(n14384), .Z(n14221) );
  AND U14316 ( .A(n461), .B(n14385), .Z(n14384) );
  XOR U14317 ( .A(n14386), .B(n14387), .Z(n14358) );
  AND U14318 ( .A(n14388), .B(n14389), .Z(n14387) );
  XNOR U14319 ( .A(n14295), .B(n14386), .Z(n14389) );
  XNOR U14320 ( .A(n14390), .B(n14391), .Z(n14295) );
  AND U14321 ( .A(n453), .B(n14392), .Z(n14391) );
  XNOR U14322 ( .A(n14393), .B(n14390), .Z(n14392) );
  XOR U14323 ( .A(n14386), .B(n14232), .Z(n14388) );
  XOR U14324 ( .A(n14394), .B(n14395), .Z(n14232) );
  AND U14325 ( .A(n461), .B(n14396), .Z(n14395) );
  XOR U14326 ( .A(n14397), .B(n14398), .Z(n14386) );
  AND U14327 ( .A(n14399), .B(n14400), .Z(n14398) );
  XNOR U14328 ( .A(n14397), .B(n14341), .Z(n14400) );
  XNOR U14329 ( .A(n14401), .B(n14402), .Z(n14341) );
  AND U14330 ( .A(n453), .B(n14403), .Z(n14402) );
  XOR U14331 ( .A(n14404), .B(n14401), .Z(n14403) );
  XNOR U14332 ( .A(n14405), .B(n14397), .Z(n14399) );
  IV U14333 ( .A(n14244), .Z(n14405) );
  XOR U14334 ( .A(n14406), .B(n14407), .Z(n14244) );
  AND U14335 ( .A(n461), .B(n14408), .Z(n14407) );
  AND U14336 ( .A(n14362), .B(n14351), .Z(n14397) );
  XNOR U14337 ( .A(n14409), .B(n14410), .Z(n14351) );
  AND U14338 ( .A(n453), .B(n14411), .Z(n14410) );
  XNOR U14339 ( .A(n14412), .B(n14409), .Z(n14411) );
  XNOR U14340 ( .A(n14413), .B(n14414), .Z(n453) );
  AND U14341 ( .A(n14415), .B(n14416), .Z(n14414) );
  XOR U14342 ( .A(n14372), .B(n14413), .Z(n14416) );
  AND U14343 ( .A(n14417), .B(n14418), .Z(n14372) );
  XOR U14344 ( .A(n14413), .B(n14369), .Z(n14415) );
  XNOR U14345 ( .A(n14419), .B(n14420), .Z(n14369) );
  AND U14346 ( .A(n457), .B(n14375), .Z(n14420) );
  XOR U14347 ( .A(n14373), .B(n14419), .Z(n14375) );
  XOR U14348 ( .A(n14421), .B(n14422), .Z(n14413) );
  AND U14349 ( .A(n14423), .B(n14424), .Z(n14422) );
  XNOR U14350 ( .A(n14421), .B(n14417), .Z(n14424) );
  IV U14351 ( .A(n14381), .Z(n14417) );
  XOR U14352 ( .A(n14425), .B(n14426), .Z(n14381) );
  XOR U14353 ( .A(n14427), .B(n14418), .Z(n14426) );
  AND U14354 ( .A(n14393), .B(n14428), .Z(n14418) );
  AND U14355 ( .A(n14429), .B(n14430), .Z(n14427) );
  XOR U14356 ( .A(n14431), .B(n14425), .Z(n14429) );
  XNOR U14357 ( .A(n14378), .B(n14421), .Z(n14423) );
  XNOR U14358 ( .A(n14432), .B(n14433), .Z(n14378) );
  AND U14359 ( .A(n457), .B(n14385), .Z(n14433) );
  XOR U14360 ( .A(n14432), .B(n14383), .Z(n14385) );
  XOR U14361 ( .A(n14434), .B(n14435), .Z(n14421) );
  AND U14362 ( .A(n14436), .B(n14437), .Z(n14435) );
  XNOR U14363 ( .A(n14434), .B(n14393), .Z(n14437) );
  XOR U14364 ( .A(n14438), .B(n14430), .Z(n14393) );
  XNOR U14365 ( .A(n14439), .B(n14425), .Z(n14430) );
  XOR U14366 ( .A(n14440), .B(n14441), .Z(n14425) );
  AND U14367 ( .A(n14442), .B(n14443), .Z(n14441) );
  XOR U14368 ( .A(n14444), .B(n14440), .Z(n14442) );
  XNOR U14369 ( .A(n14445), .B(n14446), .Z(n14439) );
  AND U14370 ( .A(n14447), .B(n14448), .Z(n14446) );
  XOR U14371 ( .A(n14445), .B(n14449), .Z(n14447) );
  XNOR U14372 ( .A(n14431), .B(n14428), .Z(n14438) );
  AND U14373 ( .A(n14450), .B(n14451), .Z(n14428) );
  XOR U14374 ( .A(n14452), .B(n14453), .Z(n14431) );
  AND U14375 ( .A(n14454), .B(n14455), .Z(n14453) );
  XOR U14376 ( .A(n14452), .B(n14456), .Z(n14454) );
  XNOR U14377 ( .A(n14390), .B(n14434), .Z(n14436) );
  XNOR U14378 ( .A(n14457), .B(n14458), .Z(n14390) );
  AND U14379 ( .A(n457), .B(n14396), .Z(n14458) );
  XOR U14380 ( .A(n14457), .B(n14394), .Z(n14396) );
  XOR U14381 ( .A(n14459), .B(n14460), .Z(n14434) );
  AND U14382 ( .A(n14461), .B(n14462), .Z(n14460) );
  XNOR U14383 ( .A(n14459), .B(n14450), .Z(n14462) );
  IV U14384 ( .A(n14404), .Z(n14450) );
  XNOR U14385 ( .A(n14463), .B(n14443), .Z(n14404) );
  XNOR U14386 ( .A(n14464), .B(n14449), .Z(n14443) );
  XOR U14387 ( .A(n14465), .B(n14466), .Z(n14449) );
  NOR U14388 ( .A(n14467), .B(n14468), .Z(n14466) );
  XNOR U14389 ( .A(n14465), .B(n14469), .Z(n14467) );
  XNOR U14390 ( .A(n14448), .B(n14440), .Z(n14464) );
  XOR U14391 ( .A(n14470), .B(n14471), .Z(n14440) );
  AND U14392 ( .A(n14472), .B(n14473), .Z(n14471) );
  XNOR U14393 ( .A(n14470), .B(n14474), .Z(n14472) );
  XNOR U14394 ( .A(n14475), .B(n14445), .Z(n14448) );
  XOR U14395 ( .A(n14476), .B(n14477), .Z(n14445) );
  AND U14396 ( .A(n14478), .B(n14479), .Z(n14477) );
  XOR U14397 ( .A(n14476), .B(n14480), .Z(n14478) );
  XNOR U14398 ( .A(n14481), .B(n14482), .Z(n14475) );
  NOR U14399 ( .A(n14483), .B(n14484), .Z(n14482) );
  XOR U14400 ( .A(n14481), .B(n14485), .Z(n14483) );
  XNOR U14401 ( .A(n14444), .B(n14451), .Z(n14463) );
  NOR U14402 ( .A(n14412), .B(n14486), .Z(n14451) );
  XOR U14403 ( .A(n14456), .B(n14455), .Z(n14444) );
  XNOR U14404 ( .A(n14487), .B(n14452), .Z(n14455) );
  XOR U14405 ( .A(n14488), .B(n14489), .Z(n14452) );
  AND U14406 ( .A(n14490), .B(n14491), .Z(n14489) );
  XOR U14407 ( .A(n14488), .B(n14492), .Z(n14490) );
  XNOR U14408 ( .A(n14493), .B(n14494), .Z(n14487) );
  NOR U14409 ( .A(n14495), .B(n14496), .Z(n14494) );
  XNOR U14410 ( .A(n14493), .B(n14497), .Z(n14495) );
  XOR U14411 ( .A(n14498), .B(n14499), .Z(n14456) );
  NOR U14412 ( .A(n14500), .B(n14501), .Z(n14499) );
  XNOR U14413 ( .A(n14498), .B(n14502), .Z(n14500) );
  XNOR U14414 ( .A(n14401), .B(n14459), .Z(n14461) );
  XNOR U14415 ( .A(n14503), .B(n14504), .Z(n14401) );
  AND U14416 ( .A(n457), .B(n14408), .Z(n14504) );
  XOR U14417 ( .A(n14503), .B(n14406), .Z(n14408) );
  AND U14418 ( .A(n14409), .B(n14412), .Z(n14459) );
  XOR U14419 ( .A(n14505), .B(n14486), .Z(n14412) );
  XNOR U14420 ( .A(p_input[1024]), .B(p_input[608]), .Z(n14486) );
  XOR U14421 ( .A(n14474), .B(n14473), .Z(n14505) );
  XNOR U14422 ( .A(n14506), .B(n14480), .Z(n14473) );
  XNOR U14423 ( .A(n14469), .B(n14468), .Z(n14480) );
  XOR U14424 ( .A(n14507), .B(n14465), .Z(n14468) );
  XOR U14425 ( .A(p_input[1034]), .B(p_input[618]), .Z(n14465) );
  XNOR U14426 ( .A(p_input[1035]), .B(p_input[619]), .Z(n14507) );
  XOR U14427 ( .A(p_input[1036]), .B(p_input[620]), .Z(n14469) );
  XNOR U14428 ( .A(n14479), .B(n14470), .Z(n14506) );
  XOR U14429 ( .A(p_input[1025]), .B(p_input[609]), .Z(n14470) );
  XOR U14430 ( .A(n14508), .B(n14485), .Z(n14479) );
  XNOR U14431 ( .A(p_input[1039]), .B(p_input[623]), .Z(n14485) );
  XOR U14432 ( .A(n14476), .B(n14484), .Z(n14508) );
  XOR U14433 ( .A(n14509), .B(n14481), .Z(n14484) );
  XOR U14434 ( .A(p_input[1037]), .B(p_input[621]), .Z(n14481) );
  XNOR U14435 ( .A(p_input[1038]), .B(p_input[622]), .Z(n14509) );
  XOR U14436 ( .A(p_input[1033]), .B(p_input[617]), .Z(n14476) );
  XNOR U14437 ( .A(n14492), .B(n14491), .Z(n14474) );
  XNOR U14438 ( .A(n14510), .B(n14497), .Z(n14491) );
  XOR U14439 ( .A(p_input[1032]), .B(p_input[616]), .Z(n14497) );
  XOR U14440 ( .A(n14488), .B(n14496), .Z(n14510) );
  XOR U14441 ( .A(n14511), .B(n14493), .Z(n14496) );
  XOR U14442 ( .A(p_input[1030]), .B(p_input[614]), .Z(n14493) );
  XNOR U14443 ( .A(p_input[1031]), .B(p_input[615]), .Z(n14511) );
  XOR U14444 ( .A(p_input[1026]), .B(p_input[610]), .Z(n14488) );
  XNOR U14445 ( .A(n14502), .B(n14501), .Z(n14492) );
  XOR U14446 ( .A(n14512), .B(n14498), .Z(n14501) );
  XOR U14447 ( .A(p_input[1027]), .B(p_input[611]), .Z(n14498) );
  XNOR U14448 ( .A(p_input[1028]), .B(p_input[612]), .Z(n14512) );
  XOR U14449 ( .A(p_input[1029]), .B(p_input[613]), .Z(n14502) );
  XNOR U14450 ( .A(n14513), .B(n14514), .Z(n14409) );
  AND U14451 ( .A(n457), .B(n14515), .Z(n14514) );
  XNOR U14452 ( .A(n14516), .B(n14517), .Z(n457) );
  AND U14453 ( .A(n14518), .B(n14519), .Z(n14517) );
  XOR U14454 ( .A(n14516), .B(n14419), .Z(n14519) );
  XNOR U14455 ( .A(n14516), .B(n14373), .Z(n14518) );
  XOR U14456 ( .A(n14520), .B(n14521), .Z(n14516) );
  AND U14457 ( .A(n14522), .B(n14523), .Z(n14521) );
  XOR U14458 ( .A(n14520), .B(n14383), .Z(n14522) );
  XOR U14459 ( .A(n14524), .B(n14525), .Z(n14362) );
  AND U14460 ( .A(n461), .B(n14515), .Z(n14525) );
  XNOR U14461 ( .A(n14513), .B(n14524), .Z(n14515) );
  XNOR U14462 ( .A(n14526), .B(n14527), .Z(n461) );
  AND U14463 ( .A(n14528), .B(n14529), .Z(n14527) );
  XNOR U14464 ( .A(n14530), .B(n14526), .Z(n14529) );
  IV U14465 ( .A(n14419), .Z(n14530) );
  XNOR U14466 ( .A(n14531), .B(n14532), .Z(n14419) );
  AND U14467 ( .A(n464), .B(n14533), .Z(n14532) );
  XNOR U14468 ( .A(n14531), .B(n14534), .Z(n14533) );
  XNOR U14469 ( .A(n14373), .B(n14526), .Z(n14528) );
  XOR U14470 ( .A(n14535), .B(n14536), .Z(n14373) );
  AND U14471 ( .A(n472), .B(n14537), .Z(n14536) );
  XOR U14472 ( .A(n14520), .B(n14538), .Z(n14526) );
  AND U14473 ( .A(n14539), .B(n14523), .Z(n14538) );
  XNOR U14474 ( .A(n14432), .B(n14520), .Z(n14523) );
  XNOR U14475 ( .A(n14540), .B(n14541), .Z(n14432) );
  AND U14476 ( .A(n464), .B(n14542), .Z(n14541) );
  XOR U14477 ( .A(n14543), .B(n14540), .Z(n14542) );
  XNOR U14478 ( .A(n14544), .B(n14520), .Z(n14539) );
  IV U14479 ( .A(n14383), .Z(n14544) );
  XOR U14480 ( .A(n14545), .B(n14546), .Z(n14383) );
  AND U14481 ( .A(n472), .B(n14547), .Z(n14546) );
  XOR U14482 ( .A(n14548), .B(n14549), .Z(n14520) );
  AND U14483 ( .A(n14550), .B(n14551), .Z(n14549) );
  XNOR U14484 ( .A(n14457), .B(n14548), .Z(n14551) );
  XNOR U14485 ( .A(n14552), .B(n14553), .Z(n14457) );
  AND U14486 ( .A(n464), .B(n14554), .Z(n14553) );
  XNOR U14487 ( .A(n14555), .B(n14552), .Z(n14554) );
  XOR U14488 ( .A(n14548), .B(n14394), .Z(n14550) );
  XOR U14489 ( .A(n14556), .B(n14557), .Z(n14394) );
  AND U14490 ( .A(n472), .B(n14558), .Z(n14557) );
  XOR U14491 ( .A(n14559), .B(n14560), .Z(n14548) );
  AND U14492 ( .A(n14561), .B(n14562), .Z(n14560) );
  XNOR U14493 ( .A(n14559), .B(n14503), .Z(n14562) );
  XNOR U14494 ( .A(n14563), .B(n14564), .Z(n14503) );
  AND U14495 ( .A(n464), .B(n14565), .Z(n14564) );
  XOR U14496 ( .A(n14566), .B(n14563), .Z(n14565) );
  XNOR U14497 ( .A(n14567), .B(n14559), .Z(n14561) );
  IV U14498 ( .A(n14406), .Z(n14567) );
  XOR U14499 ( .A(n14568), .B(n14569), .Z(n14406) );
  AND U14500 ( .A(n472), .B(n14570), .Z(n14569) );
  AND U14501 ( .A(n14524), .B(n14513), .Z(n14559) );
  XNOR U14502 ( .A(n14571), .B(n14572), .Z(n14513) );
  AND U14503 ( .A(n464), .B(n14573), .Z(n14572) );
  XNOR U14504 ( .A(n14574), .B(n14571), .Z(n14573) );
  XNOR U14505 ( .A(n14575), .B(n14576), .Z(n464) );
  AND U14506 ( .A(n14577), .B(n14578), .Z(n14576) );
  XOR U14507 ( .A(n14534), .B(n14575), .Z(n14578) );
  AND U14508 ( .A(n14579), .B(n14580), .Z(n14534) );
  XOR U14509 ( .A(n14575), .B(n14531), .Z(n14577) );
  XNOR U14510 ( .A(n14581), .B(n14582), .Z(n14531) );
  AND U14511 ( .A(n468), .B(n14537), .Z(n14582) );
  XOR U14512 ( .A(n14535), .B(n14581), .Z(n14537) );
  XOR U14513 ( .A(n14583), .B(n14584), .Z(n14575) );
  AND U14514 ( .A(n14585), .B(n14586), .Z(n14584) );
  XNOR U14515 ( .A(n14583), .B(n14579), .Z(n14586) );
  IV U14516 ( .A(n14543), .Z(n14579) );
  XOR U14517 ( .A(n14587), .B(n14588), .Z(n14543) );
  XOR U14518 ( .A(n14589), .B(n14580), .Z(n14588) );
  AND U14519 ( .A(n14555), .B(n14590), .Z(n14580) );
  AND U14520 ( .A(n14591), .B(n14592), .Z(n14589) );
  XOR U14521 ( .A(n14593), .B(n14587), .Z(n14591) );
  XNOR U14522 ( .A(n14540), .B(n14583), .Z(n14585) );
  XNOR U14523 ( .A(n14594), .B(n14595), .Z(n14540) );
  AND U14524 ( .A(n468), .B(n14547), .Z(n14595) );
  XOR U14525 ( .A(n14594), .B(n14545), .Z(n14547) );
  XOR U14526 ( .A(n14596), .B(n14597), .Z(n14583) );
  AND U14527 ( .A(n14598), .B(n14599), .Z(n14597) );
  XNOR U14528 ( .A(n14596), .B(n14555), .Z(n14599) );
  XOR U14529 ( .A(n14600), .B(n14592), .Z(n14555) );
  XNOR U14530 ( .A(n14601), .B(n14587), .Z(n14592) );
  XOR U14531 ( .A(n14602), .B(n14603), .Z(n14587) );
  AND U14532 ( .A(n14604), .B(n14605), .Z(n14603) );
  XOR U14533 ( .A(n14606), .B(n14602), .Z(n14604) );
  XNOR U14534 ( .A(n14607), .B(n14608), .Z(n14601) );
  AND U14535 ( .A(n14609), .B(n14610), .Z(n14608) );
  XOR U14536 ( .A(n14607), .B(n14611), .Z(n14609) );
  XNOR U14537 ( .A(n14593), .B(n14590), .Z(n14600) );
  AND U14538 ( .A(n14612), .B(n14613), .Z(n14590) );
  XOR U14539 ( .A(n14614), .B(n14615), .Z(n14593) );
  AND U14540 ( .A(n14616), .B(n14617), .Z(n14615) );
  XOR U14541 ( .A(n14614), .B(n14618), .Z(n14616) );
  XNOR U14542 ( .A(n14552), .B(n14596), .Z(n14598) );
  XNOR U14543 ( .A(n14619), .B(n14620), .Z(n14552) );
  AND U14544 ( .A(n468), .B(n14558), .Z(n14620) );
  XOR U14545 ( .A(n14619), .B(n14556), .Z(n14558) );
  XOR U14546 ( .A(n14621), .B(n14622), .Z(n14596) );
  AND U14547 ( .A(n14623), .B(n14624), .Z(n14622) );
  XNOR U14548 ( .A(n14621), .B(n14612), .Z(n14624) );
  IV U14549 ( .A(n14566), .Z(n14612) );
  XNOR U14550 ( .A(n14625), .B(n14605), .Z(n14566) );
  XNOR U14551 ( .A(n14626), .B(n14611), .Z(n14605) );
  XOR U14552 ( .A(n14627), .B(n14628), .Z(n14611) );
  NOR U14553 ( .A(n14629), .B(n14630), .Z(n14628) );
  XNOR U14554 ( .A(n14627), .B(n14631), .Z(n14629) );
  XNOR U14555 ( .A(n14610), .B(n14602), .Z(n14626) );
  XOR U14556 ( .A(n14632), .B(n14633), .Z(n14602) );
  AND U14557 ( .A(n14634), .B(n14635), .Z(n14633) );
  XNOR U14558 ( .A(n14632), .B(n14636), .Z(n14634) );
  XNOR U14559 ( .A(n14637), .B(n14607), .Z(n14610) );
  XOR U14560 ( .A(n14638), .B(n14639), .Z(n14607) );
  AND U14561 ( .A(n14640), .B(n14641), .Z(n14639) );
  XOR U14562 ( .A(n14638), .B(n14642), .Z(n14640) );
  XNOR U14563 ( .A(n14643), .B(n14644), .Z(n14637) );
  NOR U14564 ( .A(n14645), .B(n14646), .Z(n14644) );
  XOR U14565 ( .A(n14643), .B(n14647), .Z(n14645) );
  XNOR U14566 ( .A(n14606), .B(n14613), .Z(n14625) );
  NOR U14567 ( .A(n14574), .B(n14648), .Z(n14613) );
  XOR U14568 ( .A(n14618), .B(n14617), .Z(n14606) );
  XNOR U14569 ( .A(n14649), .B(n14614), .Z(n14617) );
  XOR U14570 ( .A(n14650), .B(n14651), .Z(n14614) );
  AND U14571 ( .A(n14652), .B(n14653), .Z(n14651) );
  XOR U14572 ( .A(n14650), .B(n14654), .Z(n14652) );
  XNOR U14573 ( .A(n14655), .B(n14656), .Z(n14649) );
  NOR U14574 ( .A(n14657), .B(n14658), .Z(n14656) );
  XNOR U14575 ( .A(n14655), .B(n14659), .Z(n14657) );
  XOR U14576 ( .A(n14660), .B(n14661), .Z(n14618) );
  NOR U14577 ( .A(n14662), .B(n14663), .Z(n14661) );
  XNOR U14578 ( .A(n14660), .B(n14664), .Z(n14662) );
  XNOR U14579 ( .A(n14563), .B(n14621), .Z(n14623) );
  XNOR U14580 ( .A(n14665), .B(n14666), .Z(n14563) );
  AND U14581 ( .A(n468), .B(n14570), .Z(n14666) );
  XOR U14582 ( .A(n14665), .B(n14568), .Z(n14570) );
  AND U14583 ( .A(n14571), .B(n14574), .Z(n14621) );
  XOR U14584 ( .A(n14667), .B(n14648), .Z(n14574) );
  XNOR U14585 ( .A(p_input[1024]), .B(p_input[624]), .Z(n14648) );
  XOR U14586 ( .A(n14636), .B(n14635), .Z(n14667) );
  XNOR U14587 ( .A(n14668), .B(n14642), .Z(n14635) );
  XNOR U14588 ( .A(n14631), .B(n14630), .Z(n14642) );
  XOR U14589 ( .A(n14669), .B(n14627), .Z(n14630) );
  XOR U14590 ( .A(p_input[1034]), .B(p_input[634]), .Z(n14627) );
  XNOR U14591 ( .A(p_input[1035]), .B(p_input[635]), .Z(n14669) );
  XOR U14592 ( .A(p_input[1036]), .B(p_input[636]), .Z(n14631) );
  XNOR U14593 ( .A(n14641), .B(n14632), .Z(n14668) );
  XOR U14594 ( .A(p_input[1025]), .B(p_input[625]), .Z(n14632) );
  XOR U14595 ( .A(n14670), .B(n14647), .Z(n14641) );
  XNOR U14596 ( .A(p_input[1039]), .B(p_input[639]), .Z(n14647) );
  XOR U14597 ( .A(n14638), .B(n14646), .Z(n14670) );
  XOR U14598 ( .A(n14671), .B(n14643), .Z(n14646) );
  XOR U14599 ( .A(p_input[1037]), .B(p_input[637]), .Z(n14643) );
  XNOR U14600 ( .A(p_input[1038]), .B(p_input[638]), .Z(n14671) );
  XOR U14601 ( .A(p_input[1033]), .B(p_input[633]), .Z(n14638) );
  XNOR U14602 ( .A(n14654), .B(n14653), .Z(n14636) );
  XNOR U14603 ( .A(n14672), .B(n14659), .Z(n14653) );
  XOR U14604 ( .A(p_input[1032]), .B(p_input[632]), .Z(n14659) );
  XOR U14605 ( .A(n14650), .B(n14658), .Z(n14672) );
  XOR U14606 ( .A(n14673), .B(n14655), .Z(n14658) );
  XOR U14607 ( .A(p_input[1030]), .B(p_input[630]), .Z(n14655) );
  XNOR U14608 ( .A(p_input[1031]), .B(p_input[631]), .Z(n14673) );
  XOR U14609 ( .A(p_input[1026]), .B(p_input[626]), .Z(n14650) );
  XNOR U14610 ( .A(n14664), .B(n14663), .Z(n14654) );
  XOR U14611 ( .A(n14674), .B(n14660), .Z(n14663) );
  XOR U14612 ( .A(p_input[1027]), .B(p_input[627]), .Z(n14660) );
  XNOR U14613 ( .A(p_input[1028]), .B(p_input[628]), .Z(n14674) );
  XOR U14614 ( .A(p_input[1029]), .B(p_input[629]), .Z(n14664) );
  XNOR U14615 ( .A(n14675), .B(n14676), .Z(n14571) );
  AND U14616 ( .A(n468), .B(n14677), .Z(n14676) );
  XNOR U14617 ( .A(n14678), .B(n14679), .Z(n468) );
  AND U14618 ( .A(n14680), .B(n14681), .Z(n14679) );
  XOR U14619 ( .A(n14678), .B(n14581), .Z(n14681) );
  XNOR U14620 ( .A(n14678), .B(n14535), .Z(n14680) );
  XOR U14621 ( .A(n14682), .B(n14683), .Z(n14678) );
  AND U14622 ( .A(n14684), .B(n14685), .Z(n14683) );
  XOR U14623 ( .A(n14682), .B(n14545), .Z(n14684) );
  XOR U14624 ( .A(n14686), .B(n14687), .Z(n14524) );
  AND U14625 ( .A(n472), .B(n14677), .Z(n14687) );
  XNOR U14626 ( .A(n14675), .B(n14686), .Z(n14677) );
  XNOR U14627 ( .A(n14688), .B(n14689), .Z(n472) );
  AND U14628 ( .A(n14690), .B(n14691), .Z(n14689) );
  XNOR U14629 ( .A(n14692), .B(n14688), .Z(n14691) );
  IV U14630 ( .A(n14581), .Z(n14692) );
  XNOR U14631 ( .A(n14693), .B(n14694), .Z(n14581) );
  AND U14632 ( .A(n475), .B(n14695), .Z(n14694) );
  XNOR U14633 ( .A(n14693), .B(n14696), .Z(n14695) );
  XNOR U14634 ( .A(n14535), .B(n14688), .Z(n14690) );
  XOR U14635 ( .A(n14697), .B(n14698), .Z(n14535) );
  AND U14636 ( .A(n483), .B(n14699), .Z(n14698) );
  XOR U14637 ( .A(n14682), .B(n14700), .Z(n14688) );
  AND U14638 ( .A(n14701), .B(n14685), .Z(n14700) );
  XNOR U14639 ( .A(n14594), .B(n14682), .Z(n14685) );
  XNOR U14640 ( .A(n14702), .B(n14703), .Z(n14594) );
  AND U14641 ( .A(n475), .B(n14704), .Z(n14703) );
  XOR U14642 ( .A(n14705), .B(n14702), .Z(n14704) );
  XNOR U14643 ( .A(n14706), .B(n14682), .Z(n14701) );
  IV U14644 ( .A(n14545), .Z(n14706) );
  XOR U14645 ( .A(n14707), .B(n14708), .Z(n14545) );
  AND U14646 ( .A(n483), .B(n14709), .Z(n14708) );
  XOR U14647 ( .A(n14710), .B(n14711), .Z(n14682) );
  AND U14648 ( .A(n14712), .B(n14713), .Z(n14711) );
  XNOR U14649 ( .A(n14619), .B(n14710), .Z(n14713) );
  XNOR U14650 ( .A(n14714), .B(n14715), .Z(n14619) );
  AND U14651 ( .A(n475), .B(n14716), .Z(n14715) );
  XNOR U14652 ( .A(n14717), .B(n14714), .Z(n14716) );
  XOR U14653 ( .A(n14710), .B(n14556), .Z(n14712) );
  XOR U14654 ( .A(n14718), .B(n14719), .Z(n14556) );
  AND U14655 ( .A(n483), .B(n14720), .Z(n14719) );
  XOR U14656 ( .A(n14721), .B(n14722), .Z(n14710) );
  AND U14657 ( .A(n14723), .B(n14724), .Z(n14722) );
  XNOR U14658 ( .A(n14721), .B(n14665), .Z(n14724) );
  XNOR U14659 ( .A(n14725), .B(n14726), .Z(n14665) );
  AND U14660 ( .A(n475), .B(n14727), .Z(n14726) );
  XOR U14661 ( .A(n14728), .B(n14725), .Z(n14727) );
  XNOR U14662 ( .A(n14729), .B(n14721), .Z(n14723) );
  IV U14663 ( .A(n14568), .Z(n14729) );
  XOR U14664 ( .A(n14730), .B(n14731), .Z(n14568) );
  AND U14665 ( .A(n483), .B(n14732), .Z(n14731) );
  AND U14666 ( .A(n14686), .B(n14675), .Z(n14721) );
  XNOR U14667 ( .A(n14733), .B(n14734), .Z(n14675) );
  AND U14668 ( .A(n475), .B(n14735), .Z(n14734) );
  XNOR U14669 ( .A(n14736), .B(n14733), .Z(n14735) );
  XNOR U14670 ( .A(n14737), .B(n14738), .Z(n475) );
  AND U14671 ( .A(n14739), .B(n14740), .Z(n14738) );
  XOR U14672 ( .A(n14696), .B(n14737), .Z(n14740) );
  AND U14673 ( .A(n14741), .B(n14742), .Z(n14696) );
  XOR U14674 ( .A(n14737), .B(n14693), .Z(n14739) );
  XNOR U14675 ( .A(n14743), .B(n14744), .Z(n14693) );
  AND U14676 ( .A(n479), .B(n14699), .Z(n14744) );
  XOR U14677 ( .A(n14697), .B(n14743), .Z(n14699) );
  XOR U14678 ( .A(n14745), .B(n14746), .Z(n14737) );
  AND U14679 ( .A(n14747), .B(n14748), .Z(n14746) );
  XNOR U14680 ( .A(n14745), .B(n14741), .Z(n14748) );
  IV U14681 ( .A(n14705), .Z(n14741) );
  XOR U14682 ( .A(n14749), .B(n14750), .Z(n14705) );
  XOR U14683 ( .A(n14751), .B(n14742), .Z(n14750) );
  AND U14684 ( .A(n14717), .B(n14752), .Z(n14742) );
  AND U14685 ( .A(n14753), .B(n14754), .Z(n14751) );
  XOR U14686 ( .A(n14755), .B(n14749), .Z(n14753) );
  XNOR U14687 ( .A(n14702), .B(n14745), .Z(n14747) );
  XNOR U14688 ( .A(n14756), .B(n14757), .Z(n14702) );
  AND U14689 ( .A(n479), .B(n14709), .Z(n14757) );
  XOR U14690 ( .A(n14756), .B(n14707), .Z(n14709) );
  XOR U14691 ( .A(n14758), .B(n14759), .Z(n14745) );
  AND U14692 ( .A(n14760), .B(n14761), .Z(n14759) );
  XNOR U14693 ( .A(n14758), .B(n14717), .Z(n14761) );
  XOR U14694 ( .A(n14762), .B(n14754), .Z(n14717) );
  XNOR U14695 ( .A(n14763), .B(n14749), .Z(n14754) );
  XOR U14696 ( .A(n14764), .B(n14765), .Z(n14749) );
  AND U14697 ( .A(n14766), .B(n14767), .Z(n14765) );
  XOR U14698 ( .A(n14768), .B(n14764), .Z(n14766) );
  XNOR U14699 ( .A(n14769), .B(n14770), .Z(n14763) );
  AND U14700 ( .A(n14771), .B(n14772), .Z(n14770) );
  XOR U14701 ( .A(n14769), .B(n14773), .Z(n14771) );
  XNOR U14702 ( .A(n14755), .B(n14752), .Z(n14762) );
  AND U14703 ( .A(n14774), .B(n14775), .Z(n14752) );
  XOR U14704 ( .A(n14776), .B(n14777), .Z(n14755) );
  AND U14705 ( .A(n14778), .B(n14779), .Z(n14777) );
  XOR U14706 ( .A(n14776), .B(n14780), .Z(n14778) );
  XNOR U14707 ( .A(n14714), .B(n14758), .Z(n14760) );
  XNOR U14708 ( .A(n14781), .B(n14782), .Z(n14714) );
  AND U14709 ( .A(n479), .B(n14720), .Z(n14782) );
  XOR U14710 ( .A(n14781), .B(n14718), .Z(n14720) );
  XOR U14711 ( .A(n14783), .B(n14784), .Z(n14758) );
  AND U14712 ( .A(n14785), .B(n14786), .Z(n14784) );
  XNOR U14713 ( .A(n14783), .B(n14774), .Z(n14786) );
  IV U14714 ( .A(n14728), .Z(n14774) );
  XNOR U14715 ( .A(n14787), .B(n14767), .Z(n14728) );
  XNOR U14716 ( .A(n14788), .B(n14773), .Z(n14767) );
  XOR U14717 ( .A(n14789), .B(n14790), .Z(n14773) );
  NOR U14718 ( .A(n14791), .B(n14792), .Z(n14790) );
  XNOR U14719 ( .A(n14789), .B(n14793), .Z(n14791) );
  XNOR U14720 ( .A(n14772), .B(n14764), .Z(n14788) );
  XOR U14721 ( .A(n14794), .B(n14795), .Z(n14764) );
  AND U14722 ( .A(n14796), .B(n14797), .Z(n14795) );
  XNOR U14723 ( .A(n14794), .B(n14798), .Z(n14796) );
  XNOR U14724 ( .A(n14799), .B(n14769), .Z(n14772) );
  XOR U14725 ( .A(n14800), .B(n14801), .Z(n14769) );
  AND U14726 ( .A(n14802), .B(n14803), .Z(n14801) );
  XOR U14727 ( .A(n14800), .B(n14804), .Z(n14802) );
  XNOR U14728 ( .A(n14805), .B(n14806), .Z(n14799) );
  NOR U14729 ( .A(n14807), .B(n14808), .Z(n14806) );
  XOR U14730 ( .A(n14805), .B(n14809), .Z(n14807) );
  XNOR U14731 ( .A(n14768), .B(n14775), .Z(n14787) );
  NOR U14732 ( .A(n14736), .B(n14810), .Z(n14775) );
  XOR U14733 ( .A(n14780), .B(n14779), .Z(n14768) );
  XNOR U14734 ( .A(n14811), .B(n14776), .Z(n14779) );
  XOR U14735 ( .A(n14812), .B(n14813), .Z(n14776) );
  AND U14736 ( .A(n14814), .B(n14815), .Z(n14813) );
  XOR U14737 ( .A(n14812), .B(n14816), .Z(n14814) );
  XNOR U14738 ( .A(n14817), .B(n14818), .Z(n14811) );
  NOR U14739 ( .A(n14819), .B(n14820), .Z(n14818) );
  XNOR U14740 ( .A(n14817), .B(n14821), .Z(n14819) );
  XOR U14741 ( .A(n14822), .B(n14823), .Z(n14780) );
  NOR U14742 ( .A(n14824), .B(n14825), .Z(n14823) );
  XNOR U14743 ( .A(n14822), .B(n14826), .Z(n14824) );
  XNOR U14744 ( .A(n14725), .B(n14783), .Z(n14785) );
  XNOR U14745 ( .A(n14827), .B(n14828), .Z(n14725) );
  AND U14746 ( .A(n479), .B(n14732), .Z(n14828) );
  XOR U14747 ( .A(n14827), .B(n14730), .Z(n14732) );
  AND U14748 ( .A(n14733), .B(n14736), .Z(n14783) );
  XOR U14749 ( .A(n14829), .B(n14810), .Z(n14736) );
  XNOR U14750 ( .A(p_input[1024]), .B(p_input[640]), .Z(n14810) );
  XOR U14751 ( .A(n14798), .B(n14797), .Z(n14829) );
  XNOR U14752 ( .A(n14830), .B(n14804), .Z(n14797) );
  XNOR U14753 ( .A(n14793), .B(n14792), .Z(n14804) );
  XOR U14754 ( .A(n14831), .B(n14789), .Z(n14792) );
  XOR U14755 ( .A(p_input[1034]), .B(p_input[650]), .Z(n14789) );
  XNOR U14756 ( .A(p_input[1035]), .B(p_input[651]), .Z(n14831) );
  XOR U14757 ( .A(p_input[1036]), .B(p_input[652]), .Z(n14793) );
  XNOR U14758 ( .A(n14803), .B(n14794), .Z(n14830) );
  XOR U14759 ( .A(p_input[1025]), .B(p_input[641]), .Z(n14794) );
  XOR U14760 ( .A(n14832), .B(n14809), .Z(n14803) );
  XNOR U14761 ( .A(p_input[1039]), .B(p_input[655]), .Z(n14809) );
  XOR U14762 ( .A(n14800), .B(n14808), .Z(n14832) );
  XOR U14763 ( .A(n14833), .B(n14805), .Z(n14808) );
  XOR U14764 ( .A(p_input[1037]), .B(p_input[653]), .Z(n14805) );
  XNOR U14765 ( .A(p_input[1038]), .B(p_input[654]), .Z(n14833) );
  XOR U14766 ( .A(p_input[1033]), .B(p_input[649]), .Z(n14800) );
  XNOR U14767 ( .A(n14816), .B(n14815), .Z(n14798) );
  XNOR U14768 ( .A(n14834), .B(n14821), .Z(n14815) );
  XOR U14769 ( .A(p_input[1032]), .B(p_input[648]), .Z(n14821) );
  XOR U14770 ( .A(n14812), .B(n14820), .Z(n14834) );
  XOR U14771 ( .A(n14835), .B(n14817), .Z(n14820) );
  XOR U14772 ( .A(p_input[1030]), .B(p_input[646]), .Z(n14817) );
  XNOR U14773 ( .A(p_input[1031]), .B(p_input[647]), .Z(n14835) );
  XOR U14774 ( .A(p_input[1026]), .B(p_input[642]), .Z(n14812) );
  XNOR U14775 ( .A(n14826), .B(n14825), .Z(n14816) );
  XOR U14776 ( .A(n14836), .B(n14822), .Z(n14825) );
  XOR U14777 ( .A(p_input[1027]), .B(p_input[643]), .Z(n14822) );
  XNOR U14778 ( .A(p_input[1028]), .B(p_input[644]), .Z(n14836) );
  XOR U14779 ( .A(p_input[1029]), .B(p_input[645]), .Z(n14826) );
  XNOR U14780 ( .A(n14837), .B(n14838), .Z(n14733) );
  AND U14781 ( .A(n479), .B(n14839), .Z(n14838) );
  XNOR U14782 ( .A(n14840), .B(n14841), .Z(n479) );
  AND U14783 ( .A(n14842), .B(n14843), .Z(n14841) );
  XOR U14784 ( .A(n14840), .B(n14743), .Z(n14843) );
  XNOR U14785 ( .A(n14840), .B(n14697), .Z(n14842) );
  XOR U14786 ( .A(n14844), .B(n14845), .Z(n14840) );
  AND U14787 ( .A(n14846), .B(n14847), .Z(n14845) );
  XOR U14788 ( .A(n14844), .B(n14707), .Z(n14846) );
  XOR U14789 ( .A(n14848), .B(n14849), .Z(n14686) );
  AND U14790 ( .A(n483), .B(n14839), .Z(n14849) );
  XNOR U14791 ( .A(n14837), .B(n14848), .Z(n14839) );
  XNOR U14792 ( .A(n14850), .B(n14851), .Z(n483) );
  AND U14793 ( .A(n14852), .B(n14853), .Z(n14851) );
  XNOR U14794 ( .A(n14854), .B(n14850), .Z(n14853) );
  IV U14795 ( .A(n14743), .Z(n14854) );
  XNOR U14796 ( .A(n14855), .B(n14856), .Z(n14743) );
  AND U14797 ( .A(n486), .B(n14857), .Z(n14856) );
  XNOR U14798 ( .A(n14855), .B(n14858), .Z(n14857) );
  XNOR U14799 ( .A(n14697), .B(n14850), .Z(n14852) );
  XOR U14800 ( .A(n14859), .B(n14860), .Z(n14697) );
  AND U14801 ( .A(n494), .B(n14861), .Z(n14860) );
  XOR U14802 ( .A(n14844), .B(n14862), .Z(n14850) );
  AND U14803 ( .A(n14863), .B(n14847), .Z(n14862) );
  XNOR U14804 ( .A(n14756), .B(n14844), .Z(n14847) );
  XNOR U14805 ( .A(n14864), .B(n14865), .Z(n14756) );
  AND U14806 ( .A(n486), .B(n14866), .Z(n14865) );
  XOR U14807 ( .A(n14867), .B(n14864), .Z(n14866) );
  XNOR U14808 ( .A(n14868), .B(n14844), .Z(n14863) );
  IV U14809 ( .A(n14707), .Z(n14868) );
  XOR U14810 ( .A(n14869), .B(n14870), .Z(n14707) );
  AND U14811 ( .A(n494), .B(n14871), .Z(n14870) );
  XOR U14812 ( .A(n14872), .B(n14873), .Z(n14844) );
  AND U14813 ( .A(n14874), .B(n14875), .Z(n14873) );
  XNOR U14814 ( .A(n14781), .B(n14872), .Z(n14875) );
  XNOR U14815 ( .A(n14876), .B(n14877), .Z(n14781) );
  AND U14816 ( .A(n486), .B(n14878), .Z(n14877) );
  XNOR U14817 ( .A(n14879), .B(n14876), .Z(n14878) );
  XOR U14818 ( .A(n14872), .B(n14718), .Z(n14874) );
  XOR U14819 ( .A(n14880), .B(n14881), .Z(n14718) );
  AND U14820 ( .A(n494), .B(n14882), .Z(n14881) );
  XOR U14821 ( .A(n14883), .B(n14884), .Z(n14872) );
  AND U14822 ( .A(n14885), .B(n14886), .Z(n14884) );
  XNOR U14823 ( .A(n14883), .B(n14827), .Z(n14886) );
  XNOR U14824 ( .A(n14887), .B(n14888), .Z(n14827) );
  AND U14825 ( .A(n486), .B(n14889), .Z(n14888) );
  XOR U14826 ( .A(n14890), .B(n14887), .Z(n14889) );
  XNOR U14827 ( .A(n14891), .B(n14883), .Z(n14885) );
  IV U14828 ( .A(n14730), .Z(n14891) );
  XOR U14829 ( .A(n14892), .B(n14893), .Z(n14730) );
  AND U14830 ( .A(n494), .B(n14894), .Z(n14893) );
  AND U14831 ( .A(n14848), .B(n14837), .Z(n14883) );
  XNOR U14832 ( .A(n14895), .B(n14896), .Z(n14837) );
  AND U14833 ( .A(n486), .B(n14897), .Z(n14896) );
  XNOR U14834 ( .A(n14898), .B(n14895), .Z(n14897) );
  XNOR U14835 ( .A(n14899), .B(n14900), .Z(n486) );
  AND U14836 ( .A(n14901), .B(n14902), .Z(n14900) );
  XOR U14837 ( .A(n14858), .B(n14899), .Z(n14902) );
  AND U14838 ( .A(n14903), .B(n14904), .Z(n14858) );
  XOR U14839 ( .A(n14899), .B(n14855), .Z(n14901) );
  XNOR U14840 ( .A(n14905), .B(n14906), .Z(n14855) );
  AND U14841 ( .A(n490), .B(n14861), .Z(n14906) );
  XOR U14842 ( .A(n14859), .B(n14905), .Z(n14861) );
  XOR U14843 ( .A(n14907), .B(n14908), .Z(n14899) );
  AND U14844 ( .A(n14909), .B(n14910), .Z(n14908) );
  XNOR U14845 ( .A(n14907), .B(n14903), .Z(n14910) );
  IV U14846 ( .A(n14867), .Z(n14903) );
  XOR U14847 ( .A(n14911), .B(n14912), .Z(n14867) );
  XOR U14848 ( .A(n14913), .B(n14904), .Z(n14912) );
  AND U14849 ( .A(n14879), .B(n14914), .Z(n14904) );
  AND U14850 ( .A(n14915), .B(n14916), .Z(n14913) );
  XOR U14851 ( .A(n14917), .B(n14911), .Z(n14915) );
  XNOR U14852 ( .A(n14864), .B(n14907), .Z(n14909) );
  XNOR U14853 ( .A(n14918), .B(n14919), .Z(n14864) );
  AND U14854 ( .A(n490), .B(n14871), .Z(n14919) );
  XOR U14855 ( .A(n14918), .B(n14869), .Z(n14871) );
  XOR U14856 ( .A(n14920), .B(n14921), .Z(n14907) );
  AND U14857 ( .A(n14922), .B(n14923), .Z(n14921) );
  XNOR U14858 ( .A(n14920), .B(n14879), .Z(n14923) );
  XOR U14859 ( .A(n14924), .B(n14916), .Z(n14879) );
  XNOR U14860 ( .A(n14925), .B(n14911), .Z(n14916) );
  XOR U14861 ( .A(n14926), .B(n14927), .Z(n14911) );
  AND U14862 ( .A(n14928), .B(n14929), .Z(n14927) );
  XOR U14863 ( .A(n14930), .B(n14926), .Z(n14928) );
  XNOR U14864 ( .A(n14931), .B(n14932), .Z(n14925) );
  AND U14865 ( .A(n14933), .B(n14934), .Z(n14932) );
  XOR U14866 ( .A(n14931), .B(n14935), .Z(n14933) );
  XNOR U14867 ( .A(n14917), .B(n14914), .Z(n14924) );
  AND U14868 ( .A(n14936), .B(n14937), .Z(n14914) );
  XOR U14869 ( .A(n14938), .B(n14939), .Z(n14917) );
  AND U14870 ( .A(n14940), .B(n14941), .Z(n14939) );
  XOR U14871 ( .A(n14938), .B(n14942), .Z(n14940) );
  XNOR U14872 ( .A(n14876), .B(n14920), .Z(n14922) );
  XNOR U14873 ( .A(n14943), .B(n14944), .Z(n14876) );
  AND U14874 ( .A(n490), .B(n14882), .Z(n14944) );
  XOR U14875 ( .A(n14943), .B(n14880), .Z(n14882) );
  XOR U14876 ( .A(n14945), .B(n14946), .Z(n14920) );
  AND U14877 ( .A(n14947), .B(n14948), .Z(n14946) );
  XNOR U14878 ( .A(n14945), .B(n14936), .Z(n14948) );
  IV U14879 ( .A(n14890), .Z(n14936) );
  XNOR U14880 ( .A(n14949), .B(n14929), .Z(n14890) );
  XNOR U14881 ( .A(n14950), .B(n14935), .Z(n14929) );
  XOR U14882 ( .A(n14951), .B(n14952), .Z(n14935) );
  NOR U14883 ( .A(n14953), .B(n14954), .Z(n14952) );
  XNOR U14884 ( .A(n14951), .B(n14955), .Z(n14953) );
  XNOR U14885 ( .A(n14934), .B(n14926), .Z(n14950) );
  XOR U14886 ( .A(n14956), .B(n14957), .Z(n14926) );
  AND U14887 ( .A(n14958), .B(n14959), .Z(n14957) );
  XNOR U14888 ( .A(n14956), .B(n14960), .Z(n14958) );
  XNOR U14889 ( .A(n14961), .B(n14931), .Z(n14934) );
  XOR U14890 ( .A(n14962), .B(n14963), .Z(n14931) );
  AND U14891 ( .A(n14964), .B(n14965), .Z(n14963) );
  XOR U14892 ( .A(n14962), .B(n14966), .Z(n14964) );
  XNOR U14893 ( .A(n14967), .B(n14968), .Z(n14961) );
  NOR U14894 ( .A(n14969), .B(n14970), .Z(n14968) );
  XOR U14895 ( .A(n14967), .B(n14971), .Z(n14969) );
  XNOR U14896 ( .A(n14930), .B(n14937), .Z(n14949) );
  NOR U14897 ( .A(n14898), .B(n14972), .Z(n14937) );
  XOR U14898 ( .A(n14942), .B(n14941), .Z(n14930) );
  XNOR U14899 ( .A(n14973), .B(n14938), .Z(n14941) );
  XOR U14900 ( .A(n14974), .B(n14975), .Z(n14938) );
  AND U14901 ( .A(n14976), .B(n14977), .Z(n14975) );
  XOR U14902 ( .A(n14974), .B(n14978), .Z(n14976) );
  XNOR U14903 ( .A(n14979), .B(n14980), .Z(n14973) );
  NOR U14904 ( .A(n14981), .B(n14982), .Z(n14980) );
  XNOR U14905 ( .A(n14979), .B(n14983), .Z(n14981) );
  XOR U14906 ( .A(n14984), .B(n14985), .Z(n14942) );
  NOR U14907 ( .A(n14986), .B(n14987), .Z(n14985) );
  XNOR U14908 ( .A(n14984), .B(n14988), .Z(n14986) );
  XNOR U14909 ( .A(n14887), .B(n14945), .Z(n14947) );
  XNOR U14910 ( .A(n14989), .B(n14990), .Z(n14887) );
  AND U14911 ( .A(n490), .B(n14894), .Z(n14990) );
  XOR U14912 ( .A(n14989), .B(n14892), .Z(n14894) );
  AND U14913 ( .A(n14895), .B(n14898), .Z(n14945) );
  XOR U14914 ( .A(n14991), .B(n14972), .Z(n14898) );
  XNOR U14915 ( .A(p_input[1024]), .B(p_input[656]), .Z(n14972) );
  XOR U14916 ( .A(n14960), .B(n14959), .Z(n14991) );
  XNOR U14917 ( .A(n14992), .B(n14966), .Z(n14959) );
  XNOR U14918 ( .A(n14955), .B(n14954), .Z(n14966) );
  XOR U14919 ( .A(n14993), .B(n14951), .Z(n14954) );
  XOR U14920 ( .A(p_input[1034]), .B(p_input[666]), .Z(n14951) );
  XNOR U14921 ( .A(p_input[1035]), .B(p_input[667]), .Z(n14993) );
  XOR U14922 ( .A(p_input[1036]), .B(p_input[668]), .Z(n14955) );
  XNOR U14923 ( .A(n14965), .B(n14956), .Z(n14992) );
  XOR U14924 ( .A(p_input[1025]), .B(p_input[657]), .Z(n14956) );
  XOR U14925 ( .A(n14994), .B(n14971), .Z(n14965) );
  XNOR U14926 ( .A(p_input[1039]), .B(p_input[671]), .Z(n14971) );
  XOR U14927 ( .A(n14962), .B(n14970), .Z(n14994) );
  XOR U14928 ( .A(n14995), .B(n14967), .Z(n14970) );
  XOR U14929 ( .A(p_input[1037]), .B(p_input[669]), .Z(n14967) );
  XNOR U14930 ( .A(p_input[1038]), .B(p_input[670]), .Z(n14995) );
  XOR U14931 ( .A(p_input[1033]), .B(p_input[665]), .Z(n14962) );
  XNOR U14932 ( .A(n14978), .B(n14977), .Z(n14960) );
  XNOR U14933 ( .A(n14996), .B(n14983), .Z(n14977) );
  XOR U14934 ( .A(p_input[1032]), .B(p_input[664]), .Z(n14983) );
  XOR U14935 ( .A(n14974), .B(n14982), .Z(n14996) );
  XOR U14936 ( .A(n14997), .B(n14979), .Z(n14982) );
  XOR U14937 ( .A(p_input[1030]), .B(p_input[662]), .Z(n14979) );
  XNOR U14938 ( .A(p_input[1031]), .B(p_input[663]), .Z(n14997) );
  XOR U14939 ( .A(p_input[1026]), .B(p_input[658]), .Z(n14974) );
  XNOR U14940 ( .A(n14988), .B(n14987), .Z(n14978) );
  XOR U14941 ( .A(n14998), .B(n14984), .Z(n14987) );
  XOR U14942 ( .A(p_input[1027]), .B(p_input[659]), .Z(n14984) );
  XNOR U14943 ( .A(p_input[1028]), .B(p_input[660]), .Z(n14998) );
  XOR U14944 ( .A(p_input[1029]), .B(p_input[661]), .Z(n14988) );
  XNOR U14945 ( .A(n14999), .B(n15000), .Z(n14895) );
  AND U14946 ( .A(n490), .B(n15001), .Z(n15000) );
  XNOR U14947 ( .A(n15002), .B(n15003), .Z(n490) );
  AND U14948 ( .A(n15004), .B(n15005), .Z(n15003) );
  XOR U14949 ( .A(n15002), .B(n14905), .Z(n15005) );
  XNOR U14950 ( .A(n15002), .B(n14859), .Z(n15004) );
  XOR U14951 ( .A(n15006), .B(n15007), .Z(n15002) );
  AND U14952 ( .A(n15008), .B(n15009), .Z(n15007) );
  XOR U14953 ( .A(n15006), .B(n14869), .Z(n15008) );
  XOR U14954 ( .A(n15010), .B(n15011), .Z(n14848) );
  AND U14955 ( .A(n494), .B(n15001), .Z(n15011) );
  XNOR U14956 ( .A(n14999), .B(n15010), .Z(n15001) );
  XNOR U14957 ( .A(n15012), .B(n15013), .Z(n494) );
  AND U14958 ( .A(n15014), .B(n15015), .Z(n15013) );
  XNOR U14959 ( .A(n15016), .B(n15012), .Z(n15015) );
  IV U14960 ( .A(n14905), .Z(n15016) );
  XNOR U14961 ( .A(n15017), .B(n15018), .Z(n14905) );
  AND U14962 ( .A(n497), .B(n15019), .Z(n15018) );
  XNOR U14963 ( .A(n15017), .B(n15020), .Z(n15019) );
  XNOR U14964 ( .A(n14859), .B(n15012), .Z(n15014) );
  XOR U14965 ( .A(n15021), .B(n15022), .Z(n14859) );
  AND U14966 ( .A(n505), .B(n15023), .Z(n15022) );
  XOR U14967 ( .A(n15006), .B(n15024), .Z(n15012) );
  AND U14968 ( .A(n15025), .B(n15009), .Z(n15024) );
  XNOR U14969 ( .A(n14918), .B(n15006), .Z(n15009) );
  XNOR U14970 ( .A(n15026), .B(n15027), .Z(n14918) );
  AND U14971 ( .A(n497), .B(n15028), .Z(n15027) );
  XOR U14972 ( .A(n15029), .B(n15026), .Z(n15028) );
  XNOR U14973 ( .A(n15030), .B(n15006), .Z(n15025) );
  IV U14974 ( .A(n14869), .Z(n15030) );
  XOR U14975 ( .A(n15031), .B(n15032), .Z(n14869) );
  AND U14976 ( .A(n505), .B(n15033), .Z(n15032) );
  XOR U14977 ( .A(n15034), .B(n15035), .Z(n15006) );
  AND U14978 ( .A(n15036), .B(n15037), .Z(n15035) );
  XNOR U14979 ( .A(n14943), .B(n15034), .Z(n15037) );
  XNOR U14980 ( .A(n15038), .B(n15039), .Z(n14943) );
  AND U14981 ( .A(n497), .B(n15040), .Z(n15039) );
  XNOR U14982 ( .A(n15041), .B(n15038), .Z(n15040) );
  XOR U14983 ( .A(n15034), .B(n14880), .Z(n15036) );
  XOR U14984 ( .A(n15042), .B(n15043), .Z(n14880) );
  AND U14985 ( .A(n505), .B(n15044), .Z(n15043) );
  XOR U14986 ( .A(n15045), .B(n15046), .Z(n15034) );
  AND U14987 ( .A(n15047), .B(n15048), .Z(n15046) );
  XNOR U14988 ( .A(n15045), .B(n14989), .Z(n15048) );
  XNOR U14989 ( .A(n15049), .B(n15050), .Z(n14989) );
  AND U14990 ( .A(n497), .B(n15051), .Z(n15050) );
  XOR U14991 ( .A(n15052), .B(n15049), .Z(n15051) );
  XNOR U14992 ( .A(n15053), .B(n15045), .Z(n15047) );
  IV U14993 ( .A(n14892), .Z(n15053) );
  XOR U14994 ( .A(n15054), .B(n15055), .Z(n14892) );
  AND U14995 ( .A(n505), .B(n15056), .Z(n15055) );
  AND U14996 ( .A(n15010), .B(n14999), .Z(n15045) );
  XNOR U14997 ( .A(n15057), .B(n15058), .Z(n14999) );
  AND U14998 ( .A(n497), .B(n15059), .Z(n15058) );
  XNOR U14999 ( .A(n15060), .B(n15057), .Z(n15059) );
  XNOR U15000 ( .A(n15061), .B(n15062), .Z(n497) );
  AND U15001 ( .A(n15063), .B(n15064), .Z(n15062) );
  XOR U15002 ( .A(n15020), .B(n15061), .Z(n15064) );
  AND U15003 ( .A(n15065), .B(n15066), .Z(n15020) );
  XOR U15004 ( .A(n15061), .B(n15017), .Z(n15063) );
  XNOR U15005 ( .A(n15067), .B(n15068), .Z(n15017) );
  AND U15006 ( .A(n501), .B(n15023), .Z(n15068) );
  XOR U15007 ( .A(n15021), .B(n15067), .Z(n15023) );
  XOR U15008 ( .A(n15069), .B(n15070), .Z(n15061) );
  AND U15009 ( .A(n15071), .B(n15072), .Z(n15070) );
  XNOR U15010 ( .A(n15069), .B(n15065), .Z(n15072) );
  IV U15011 ( .A(n15029), .Z(n15065) );
  XOR U15012 ( .A(n15073), .B(n15074), .Z(n15029) );
  XOR U15013 ( .A(n15075), .B(n15066), .Z(n15074) );
  AND U15014 ( .A(n15041), .B(n15076), .Z(n15066) );
  AND U15015 ( .A(n15077), .B(n15078), .Z(n15075) );
  XOR U15016 ( .A(n15079), .B(n15073), .Z(n15077) );
  XNOR U15017 ( .A(n15026), .B(n15069), .Z(n15071) );
  XNOR U15018 ( .A(n15080), .B(n15081), .Z(n15026) );
  AND U15019 ( .A(n501), .B(n15033), .Z(n15081) );
  XOR U15020 ( .A(n15080), .B(n15031), .Z(n15033) );
  XOR U15021 ( .A(n15082), .B(n15083), .Z(n15069) );
  AND U15022 ( .A(n15084), .B(n15085), .Z(n15083) );
  XNOR U15023 ( .A(n15082), .B(n15041), .Z(n15085) );
  XOR U15024 ( .A(n15086), .B(n15078), .Z(n15041) );
  XNOR U15025 ( .A(n15087), .B(n15073), .Z(n15078) );
  XOR U15026 ( .A(n15088), .B(n15089), .Z(n15073) );
  AND U15027 ( .A(n15090), .B(n15091), .Z(n15089) );
  XOR U15028 ( .A(n15092), .B(n15088), .Z(n15090) );
  XNOR U15029 ( .A(n15093), .B(n15094), .Z(n15087) );
  AND U15030 ( .A(n15095), .B(n15096), .Z(n15094) );
  XOR U15031 ( .A(n15093), .B(n15097), .Z(n15095) );
  XNOR U15032 ( .A(n15079), .B(n15076), .Z(n15086) );
  AND U15033 ( .A(n15098), .B(n15099), .Z(n15076) );
  XOR U15034 ( .A(n15100), .B(n15101), .Z(n15079) );
  AND U15035 ( .A(n15102), .B(n15103), .Z(n15101) );
  XOR U15036 ( .A(n15100), .B(n15104), .Z(n15102) );
  XNOR U15037 ( .A(n15038), .B(n15082), .Z(n15084) );
  XNOR U15038 ( .A(n15105), .B(n15106), .Z(n15038) );
  AND U15039 ( .A(n501), .B(n15044), .Z(n15106) );
  XOR U15040 ( .A(n15105), .B(n15042), .Z(n15044) );
  XOR U15041 ( .A(n15107), .B(n15108), .Z(n15082) );
  AND U15042 ( .A(n15109), .B(n15110), .Z(n15108) );
  XNOR U15043 ( .A(n15107), .B(n15098), .Z(n15110) );
  IV U15044 ( .A(n15052), .Z(n15098) );
  XNOR U15045 ( .A(n15111), .B(n15091), .Z(n15052) );
  XNOR U15046 ( .A(n15112), .B(n15097), .Z(n15091) );
  XOR U15047 ( .A(n15113), .B(n15114), .Z(n15097) );
  NOR U15048 ( .A(n15115), .B(n15116), .Z(n15114) );
  XNOR U15049 ( .A(n15113), .B(n15117), .Z(n15115) );
  XNOR U15050 ( .A(n15096), .B(n15088), .Z(n15112) );
  XOR U15051 ( .A(n15118), .B(n15119), .Z(n15088) );
  AND U15052 ( .A(n15120), .B(n15121), .Z(n15119) );
  XNOR U15053 ( .A(n15118), .B(n15122), .Z(n15120) );
  XNOR U15054 ( .A(n15123), .B(n15093), .Z(n15096) );
  XOR U15055 ( .A(n15124), .B(n15125), .Z(n15093) );
  AND U15056 ( .A(n15126), .B(n15127), .Z(n15125) );
  XOR U15057 ( .A(n15124), .B(n15128), .Z(n15126) );
  XNOR U15058 ( .A(n15129), .B(n15130), .Z(n15123) );
  NOR U15059 ( .A(n15131), .B(n15132), .Z(n15130) );
  XOR U15060 ( .A(n15129), .B(n15133), .Z(n15131) );
  XNOR U15061 ( .A(n15092), .B(n15099), .Z(n15111) );
  NOR U15062 ( .A(n15060), .B(n15134), .Z(n15099) );
  XOR U15063 ( .A(n15104), .B(n15103), .Z(n15092) );
  XNOR U15064 ( .A(n15135), .B(n15100), .Z(n15103) );
  XOR U15065 ( .A(n15136), .B(n15137), .Z(n15100) );
  AND U15066 ( .A(n15138), .B(n15139), .Z(n15137) );
  XOR U15067 ( .A(n15136), .B(n15140), .Z(n15138) );
  XNOR U15068 ( .A(n15141), .B(n15142), .Z(n15135) );
  NOR U15069 ( .A(n15143), .B(n15144), .Z(n15142) );
  XNOR U15070 ( .A(n15141), .B(n15145), .Z(n15143) );
  XOR U15071 ( .A(n15146), .B(n15147), .Z(n15104) );
  NOR U15072 ( .A(n15148), .B(n15149), .Z(n15147) );
  XNOR U15073 ( .A(n15146), .B(n15150), .Z(n15148) );
  XNOR U15074 ( .A(n15049), .B(n15107), .Z(n15109) );
  XNOR U15075 ( .A(n15151), .B(n15152), .Z(n15049) );
  AND U15076 ( .A(n501), .B(n15056), .Z(n15152) );
  XOR U15077 ( .A(n15151), .B(n15054), .Z(n15056) );
  AND U15078 ( .A(n15057), .B(n15060), .Z(n15107) );
  XOR U15079 ( .A(n15153), .B(n15134), .Z(n15060) );
  XNOR U15080 ( .A(p_input[1024]), .B(p_input[672]), .Z(n15134) );
  XOR U15081 ( .A(n15122), .B(n15121), .Z(n15153) );
  XNOR U15082 ( .A(n15154), .B(n15128), .Z(n15121) );
  XNOR U15083 ( .A(n15117), .B(n15116), .Z(n15128) );
  XOR U15084 ( .A(n15155), .B(n15113), .Z(n15116) );
  XOR U15085 ( .A(p_input[1034]), .B(p_input[682]), .Z(n15113) );
  XNOR U15086 ( .A(p_input[1035]), .B(p_input[683]), .Z(n15155) );
  XOR U15087 ( .A(p_input[1036]), .B(p_input[684]), .Z(n15117) );
  XNOR U15088 ( .A(n15127), .B(n15118), .Z(n15154) );
  XOR U15089 ( .A(p_input[1025]), .B(p_input[673]), .Z(n15118) );
  XOR U15090 ( .A(n15156), .B(n15133), .Z(n15127) );
  XNOR U15091 ( .A(p_input[1039]), .B(p_input[687]), .Z(n15133) );
  XOR U15092 ( .A(n15124), .B(n15132), .Z(n15156) );
  XOR U15093 ( .A(n15157), .B(n15129), .Z(n15132) );
  XOR U15094 ( .A(p_input[1037]), .B(p_input[685]), .Z(n15129) );
  XNOR U15095 ( .A(p_input[1038]), .B(p_input[686]), .Z(n15157) );
  XOR U15096 ( .A(p_input[1033]), .B(p_input[681]), .Z(n15124) );
  XNOR U15097 ( .A(n15140), .B(n15139), .Z(n15122) );
  XNOR U15098 ( .A(n15158), .B(n15145), .Z(n15139) );
  XOR U15099 ( .A(p_input[1032]), .B(p_input[680]), .Z(n15145) );
  XOR U15100 ( .A(n15136), .B(n15144), .Z(n15158) );
  XOR U15101 ( .A(n15159), .B(n15141), .Z(n15144) );
  XOR U15102 ( .A(p_input[1030]), .B(p_input[678]), .Z(n15141) );
  XNOR U15103 ( .A(p_input[1031]), .B(p_input[679]), .Z(n15159) );
  XOR U15104 ( .A(p_input[1026]), .B(p_input[674]), .Z(n15136) );
  XNOR U15105 ( .A(n15150), .B(n15149), .Z(n15140) );
  XOR U15106 ( .A(n15160), .B(n15146), .Z(n15149) );
  XOR U15107 ( .A(p_input[1027]), .B(p_input[675]), .Z(n15146) );
  XNOR U15108 ( .A(p_input[1028]), .B(p_input[676]), .Z(n15160) );
  XOR U15109 ( .A(p_input[1029]), .B(p_input[677]), .Z(n15150) );
  XNOR U15110 ( .A(n15161), .B(n15162), .Z(n15057) );
  AND U15111 ( .A(n501), .B(n15163), .Z(n15162) );
  XNOR U15112 ( .A(n15164), .B(n15165), .Z(n501) );
  AND U15113 ( .A(n15166), .B(n15167), .Z(n15165) );
  XOR U15114 ( .A(n15164), .B(n15067), .Z(n15167) );
  XNOR U15115 ( .A(n15164), .B(n15021), .Z(n15166) );
  XOR U15116 ( .A(n15168), .B(n15169), .Z(n15164) );
  AND U15117 ( .A(n15170), .B(n15171), .Z(n15169) );
  XOR U15118 ( .A(n15168), .B(n15031), .Z(n15170) );
  XOR U15119 ( .A(n15172), .B(n15173), .Z(n15010) );
  AND U15120 ( .A(n505), .B(n15163), .Z(n15173) );
  XNOR U15121 ( .A(n15161), .B(n15172), .Z(n15163) );
  XNOR U15122 ( .A(n15174), .B(n15175), .Z(n505) );
  AND U15123 ( .A(n15176), .B(n15177), .Z(n15175) );
  XNOR U15124 ( .A(n15178), .B(n15174), .Z(n15177) );
  IV U15125 ( .A(n15067), .Z(n15178) );
  XNOR U15126 ( .A(n15179), .B(n15180), .Z(n15067) );
  AND U15127 ( .A(n508), .B(n15181), .Z(n15180) );
  XNOR U15128 ( .A(n15179), .B(n15182), .Z(n15181) );
  XNOR U15129 ( .A(n15021), .B(n15174), .Z(n15176) );
  XOR U15130 ( .A(n15183), .B(n15184), .Z(n15021) );
  AND U15131 ( .A(n516), .B(n15185), .Z(n15184) );
  XOR U15132 ( .A(n15168), .B(n15186), .Z(n15174) );
  AND U15133 ( .A(n15187), .B(n15171), .Z(n15186) );
  XNOR U15134 ( .A(n15080), .B(n15168), .Z(n15171) );
  XNOR U15135 ( .A(n15188), .B(n15189), .Z(n15080) );
  AND U15136 ( .A(n508), .B(n15190), .Z(n15189) );
  XOR U15137 ( .A(n15191), .B(n15188), .Z(n15190) );
  XNOR U15138 ( .A(n15192), .B(n15168), .Z(n15187) );
  IV U15139 ( .A(n15031), .Z(n15192) );
  XOR U15140 ( .A(n15193), .B(n15194), .Z(n15031) );
  AND U15141 ( .A(n516), .B(n15195), .Z(n15194) );
  XOR U15142 ( .A(n15196), .B(n15197), .Z(n15168) );
  AND U15143 ( .A(n15198), .B(n15199), .Z(n15197) );
  XNOR U15144 ( .A(n15105), .B(n15196), .Z(n15199) );
  XNOR U15145 ( .A(n15200), .B(n15201), .Z(n15105) );
  AND U15146 ( .A(n508), .B(n15202), .Z(n15201) );
  XNOR U15147 ( .A(n15203), .B(n15200), .Z(n15202) );
  XOR U15148 ( .A(n15196), .B(n15042), .Z(n15198) );
  XOR U15149 ( .A(n15204), .B(n15205), .Z(n15042) );
  AND U15150 ( .A(n516), .B(n15206), .Z(n15205) );
  XOR U15151 ( .A(n15207), .B(n15208), .Z(n15196) );
  AND U15152 ( .A(n15209), .B(n15210), .Z(n15208) );
  XNOR U15153 ( .A(n15207), .B(n15151), .Z(n15210) );
  XNOR U15154 ( .A(n15211), .B(n15212), .Z(n15151) );
  AND U15155 ( .A(n508), .B(n15213), .Z(n15212) );
  XOR U15156 ( .A(n15214), .B(n15211), .Z(n15213) );
  XNOR U15157 ( .A(n15215), .B(n15207), .Z(n15209) );
  IV U15158 ( .A(n15054), .Z(n15215) );
  XOR U15159 ( .A(n15216), .B(n15217), .Z(n15054) );
  AND U15160 ( .A(n516), .B(n15218), .Z(n15217) );
  AND U15161 ( .A(n15172), .B(n15161), .Z(n15207) );
  XNOR U15162 ( .A(n15219), .B(n15220), .Z(n15161) );
  AND U15163 ( .A(n508), .B(n15221), .Z(n15220) );
  XNOR U15164 ( .A(n15222), .B(n15219), .Z(n15221) );
  XNOR U15165 ( .A(n15223), .B(n15224), .Z(n508) );
  AND U15166 ( .A(n15225), .B(n15226), .Z(n15224) );
  XOR U15167 ( .A(n15182), .B(n15223), .Z(n15226) );
  AND U15168 ( .A(n15227), .B(n15228), .Z(n15182) );
  XOR U15169 ( .A(n15223), .B(n15179), .Z(n15225) );
  XNOR U15170 ( .A(n15229), .B(n15230), .Z(n15179) );
  AND U15171 ( .A(n512), .B(n15185), .Z(n15230) );
  XOR U15172 ( .A(n15183), .B(n15229), .Z(n15185) );
  XOR U15173 ( .A(n15231), .B(n15232), .Z(n15223) );
  AND U15174 ( .A(n15233), .B(n15234), .Z(n15232) );
  XNOR U15175 ( .A(n15231), .B(n15227), .Z(n15234) );
  IV U15176 ( .A(n15191), .Z(n15227) );
  XOR U15177 ( .A(n15235), .B(n15236), .Z(n15191) );
  XOR U15178 ( .A(n15237), .B(n15228), .Z(n15236) );
  AND U15179 ( .A(n15203), .B(n15238), .Z(n15228) );
  AND U15180 ( .A(n15239), .B(n15240), .Z(n15237) );
  XOR U15181 ( .A(n15241), .B(n15235), .Z(n15239) );
  XNOR U15182 ( .A(n15188), .B(n15231), .Z(n15233) );
  XNOR U15183 ( .A(n15242), .B(n15243), .Z(n15188) );
  AND U15184 ( .A(n512), .B(n15195), .Z(n15243) );
  XOR U15185 ( .A(n15242), .B(n15193), .Z(n15195) );
  XOR U15186 ( .A(n15244), .B(n15245), .Z(n15231) );
  AND U15187 ( .A(n15246), .B(n15247), .Z(n15245) );
  XNOR U15188 ( .A(n15244), .B(n15203), .Z(n15247) );
  XOR U15189 ( .A(n15248), .B(n15240), .Z(n15203) );
  XNOR U15190 ( .A(n15249), .B(n15235), .Z(n15240) );
  XOR U15191 ( .A(n15250), .B(n15251), .Z(n15235) );
  AND U15192 ( .A(n15252), .B(n15253), .Z(n15251) );
  XOR U15193 ( .A(n15254), .B(n15250), .Z(n15252) );
  XNOR U15194 ( .A(n15255), .B(n15256), .Z(n15249) );
  AND U15195 ( .A(n15257), .B(n15258), .Z(n15256) );
  XOR U15196 ( .A(n15255), .B(n15259), .Z(n15257) );
  XNOR U15197 ( .A(n15241), .B(n15238), .Z(n15248) );
  AND U15198 ( .A(n15260), .B(n15261), .Z(n15238) );
  XOR U15199 ( .A(n15262), .B(n15263), .Z(n15241) );
  AND U15200 ( .A(n15264), .B(n15265), .Z(n15263) );
  XOR U15201 ( .A(n15262), .B(n15266), .Z(n15264) );
  XNOR U15202 ( .A(n15200), .B(n15244), .Z(n15246) );
  XNOR U15203 ( .A(n15267), .B(n15268), .Z(n15200) );
  AND U15204 ( .A(n512), .B(n15206), .Z(n15268) );
  XOR U15205 ( .A(n15267), .B(n15204), .Z(n15206) );
  XOR U15206 ( .A(n15269), .B(n15270), .Z(n15244) );
  AND U15207 ( .A(n15271), .B(n15272), .Z(n15270) );
  XNOR U15208 ( .A(n15269), .B(n15260), .Z(n15272) );
  IV U15209 ( .A(n15214), .Z(n15260) );
  XNOR U15210 ( .A(n15273), .B(n15253), .Z(n15214) );
  XNOR U15211 ( .A(n15274), .B(n15259), .Z(n15253) );
  XOR U15212 ( .A(n15275), .B(n15276), .Z(n15259) );
  NOR U15213 ( .A(n15277), .B(n15278), .Z(n15276) );
  XNOR U15214 ( .A(n15275), .B(n15279), .Z(n15277) );
  XNOR U15215 ( .A(n15258), .B(n15250), .Z(n15274) );
  XOR U15216 ( .A(n15280), .B(n15281), .Z(n15250) );
  AND U15217 ( .A(n15282), .B(n15283), .Z(n15281) );
  XNOR U15218 ( .A(n15280), .B(n15284), .Z(n15282) );
  XNOR U15219 ( .A(n15285), .B(n15255), .Z(n15258) );
  XOR U15220 ( .A(n15286), .B(n15287), .Z(n15255) );
  AND U15221 ( .A(n15288), .B(n15289), .Z(n15287) );
  XOR U15222 ( .A(n15286), .B(n15290), .Z(n15288) );
  XNOR U15223 ( .A(n15291), .B(n15292), .Z(n15285) );
  NOR U15224 ( .A(n15293), .B(n15294), .Z(n15292) );
  XOR U15225 ( .A(n15291), .B(n15295), .Z(n15293) );
  XNOR U15226 ( .A(n15254), .B(n15261), .Z(n15273) );
  NOR U15227 ( .A(n15222), .B(n15296), .Z(n15261) );
  XOR U15228 ( .A(n15266), .B(n15265), .Z(n15254) );
  XNOR U15229 ( .A(n15297), .B(n15262), .Z(n15265) );
  XOR U15230 ( .A(n15298), .B(n15299), .Z(n15262) );
  AND U15231 ( .A(n15300), .B(n15301), .Z(n15299) );
  XOR U15232 ( .A(n15298), .B(n15302), .Z(n15300) );
  XNOR U15233 ( .A(n15303), .B(n15304), .Z(n15297) );
  NOR U15234 ( .A(n15305), .B(n15306), .Z(n15304) );
  XNOR U15235 ( .A(n15303), .B(n15307), .Z(n15305) );
  XOR U15236 ( .A(n15308), .B(n15309), .Z(n15266) );
  NOR U15237 ( .A(n15310), .B(n15311), .Z(n15309) );
  XNOR U15238 ( .A(n15308), .B(n15312), .Z(n15310) );
  XNOR U15239 ( .A(n15211), .B(n15269), .Z(n15271) );
  XNOR U15240 ( .A(n15313), .B(n15314), .Z(n15211) );
  AND U15241 ( .A(n512), .B(n15218), .Z(n15314) );
  XOR U15242 ( .A(n15313), .B(n15216), .Z(n15218) );
  AND U15243 ( .A(n15219), .B(n15222), .Z(n15269) );
  XOR U15244 ( .A(n15315), .B(n15296), .Z(n15222) );
  XNOR U15245 ( .A(p_input[1024]), .B(p_input[688]), .Z(n15296) );
  XOR U15246 ( .A(n15284), .B(n15283), .Z(n15315) );
  XNOR U15247 ( .A(n15316), .B(n15290), .Z(n15283) );
  XNOR U15248 ( .A(n15279), .B(n15278), .Z(n15290) );
  XOR U15249 ( .A(n15317), .B(n15275), .Z(n15278) );
  XOR U15250 ( .A(p_input[1034]), .B(p_input[698]), .Z(n15275) );
  XNOR U15251 ( .A(p_input[1035]), .B(p_input[699]), .Z(n15317) );
  XOR U15252 ( .A(p_input[1036]), .B(p_input[700]), .Z(n15279) );
  XNOR U15253 ( .A(n15289), .B(n15280), .Z(n15316) );
  XOR U15254 ( .A(p_input[1025]), .B(p_input[689]), .Z(n15280) );
  XOR U15255 ( .A(n15318), .B(n15295), .Z(n15289) );
  XNOR U15256 ( .A(p_input[1039]), .B(p_input[703]), .Z(n15295) );
  XOR U15257 ( .A(n15286), .B(n15294), .Z(n15318) );
  XOR U15258 ( .A(n15319), .B(n15291), .Z(n15294) );
  XOR U15259 ( .A(p_input[1037]), .B(p_input[701]), .Z(n15291) );
  XNOR U15260 ( .A(p_input[1038]), .B(p_input[702]), .Z(n15319) );
  XOR U15261 ( .A(p_input[1033]), .B(p_input[697]), .Z(n15286) );
  XNOR U15262 ( .A(n15302), .B(n15301), .Z(n15284) );
  XNOR U15263 ( .A(n15320), .B(n15307), .Z(n15301) );
  XOR U15264 ( .A(p_input[1032]), .B(p_input[696]), .Z(n15307) );
  XOR U15265 ( .A(n15298), .B(n15306), .Z(n15320) );
  XOR U15266 ( .A(n15321), .B(n15303), .Z(n15306) );
  XOR U15267 ( .A(p_input[1030]), .B(p_input[694]), .Z(n15303) );
  XNOR U15268 ( .A(p_input[1031]), .B(p_input[695]), .Z(n15321) );
  XOR U15269 ( .A(p_input[1026]), .B(p_input[690]), .Z(n15298) );
  XNOR U15270 ( .A(n15312), .B(n15311), .Z(n15302) );
  XOR U15271 ( .A(n15322), .B(n15308), .Z(n15311) );
  XOR U15272 ( .A(p_input[1027]), .B(p_input[691]), .Z(n15308) );
  XNOR U15273 ( .A(p_input[1028]), .B(p_input[692]), .Z(n15322) );
  XOR U15274 ( .A(p_input[1029]), .B(p_input[693]), .Z(n15312) );
  XNOR U15275 ( .A(n15323), .B(n15324), .Z(n15219) );
  AND U15276 ( .A(n512), .B(n15325), .Z(n15324) );
  XNOR U15277 ( .A(n15326), .B(n15327), .Z(n512) );
  AND U15278 ( .A(n15328), .B(n15329), .Z(n15327) );
  XOR U15279 ( .A(n15326), .B(n15229), .Z(n15329) );
  XNOR U15280 ( .A(n15326), .B(n15183), .Z(n15328) );
  XOR U15281 ( .A(n15330), .B(n15331), .Z(n15326) );
  AND U15282 ( .A(n15332), .B(n15333), .Z(n15331) );
  XOR U15283 ( .A(n15330), .B(n15193), .Z(n15332) );
  XOR U15284 ( .A(n15334), .B(n15335), .Z(n15172) );
  AND U15285 ( .A(n516), .B(n15325), .Z(n15335) );
  XNOR U15286 ( .A(n15323), .B(n15334), .Z(n15325) );
  XNOR U15287 ( .A(n15336), .B(n15337), .Z(n516) );
  AND U15288 ( .A(n15338), .B(n15339), .Z(n15337) );
  XNOR U15289 ( .A(n15340), .B(n15336), .Z(n15339) );
  IV U15290 ( .A(n15229), .Z(n15340) );
  XNOR U15291 ( .A(n15341), .B(n15342), .Z(n15229) );
  AND U15292 ( .A(n519), .B(n15343), .Z(n15342) );
  XNOR U15293 ( .A(n15341), .B(n15344), .Z(n15343) );
  XNOR U15294 ( .A(n15183), .B(n15336), .Z(n15338) );
  XOR U15295 ( .A(n15345), .B(n15346), .Z(n15183) );
  AND U15296 ( .A(n527), .B(n15347), .Z(n15346) );
  XOR U15297 ( .A(n15330), .B(n15348), .Z(n15336) );
  AND U15298 ( .A(n15349), .B(n15333), .Z(n15348) );
  XNOR U15299 ( .A(n15242), .B(n15330), .Z(n15333) );
  XNOR U15300 ( .A(n15350), .B(n15351), .Z(n15242) );
  AND U15301 ( .A(n519), .B(n15352), .Z(n15351) );
  XOR U15302 ( .A(n15353), .B(n15350), .Z(n15352) );
  XNOR U15303 ( .A(n15354), .B(n15330), .Z(n15349) );
  IV U15304 ( .A(n15193), .Z(n15354) );
  XOR U15305 ( .A(n15355), .B(n15356), .Z(n15193) );
  AND U15306 ( .A(n527), .B(n15357), .Z(n15356) );
  XOR U15307 ( .A(n15358), .B(n15359), .Z(n15330) );
  AND U15308 ( .A(n15360), .B(n15361), .Z(n15359) );
  XNOR U15309 ( .A(n15267), .B(n15358), .Z(n15361) );
  XNOR U15310 ( .A(n15362), .B(n15363), .Z(n15267) );
  AND U15311 ( .A(n519), .B(n15364), .Z(n15363) );
  XNOR U15312 ( .A(n15365), .B(n15362), .Z(n15364) );
  XOR U15313 ( .A(n15358), .B(n15204), .Z(n15360) );
  XOR U15314 ( .A(n15366), .B(n15367), .Z(n15204) );
  AND U15315 ( .A(n527), .B(n15368), .Z(n15367) );
  XOR U15316 ( .A(n15369), .B(n15370), .Z(n15358) );
  AND U15317 ( .A(n15371), .B(n15372), .Z(n15370) );
  XNOR U15318 ( .A(n15369), .B(n15313), .Z(n15372) );
  XNOR U15319 ( .A(n15373), .B(n15374), .Z(n15313) );
  AND U15320 ( .A(n519), .B(n15375), .Z(n15374) );
  XOR U15321 ( .A(n15376), .B(n15373), .Z(n15375) );
  XNOR U15322 ( .A(n15377), .B(n15369), .Z(n15371) );
  IV U15323 ( .A(n15216), .Z(n15377) );
  XOR U15324 ( .A(n15378), .B(n15379), .Z(n15216) );
  AND U15325 ( .A(n527), .B(n15380), .Z(n15379) );
  AND U15326 ( .A(n15334), .B(n15323), .Z(n15369) );
  XNOR U15327 ( .A(n15381), .B(n15382), .Z(n15323) );
  AND U15328 ( .A(n519), .B(n15383), .Z(n15382) );
  XNOR U15329 ( .A(n15384), .B(n15381), .Z(n15383) );
  XNOR U15330 ( .A(n15385), .B(n15386), .Z(n519) );
  AND U15331 ( .A(n15387), .B(n15388), .Z(n15386) );
  XOR U15332 ( .A(n15344), .B(n15385), .Z(n15388) );
  AND U15333 ( .A(n15389), .B(n15390), .Z(n15344) );
  XOR U15334 ( .A(n15385), .B(n15341), .Z(n15387) );
  XNOR U15335 ( .A(n15391), .B(n15392), .Z(n15341) );
  AND U15336 ( .A(n523), .B(n15347), .Z(n15392) );
  XOR U15337 ( .A(n15345), .B(n15391), .Z(n15347) );
  XOR U15338 ( .A(n15393), .B(n15394), .Z(n15385) );
  AND U15339 ( .A(n15395), .B(n15396), .Z(n15394) );
  XNOR U15340 ( .A(n15393), .B(n15389), .Z(n15396) );
  IV U15341 ( .A(n15353), .Z(n15389) );
  XOR U15342 ( .A(n15397), .B(n15398), .Z(n15353) );
  XOR U15343 ( .A(n15399), .B(n15390), .Z(n15398) );
  AND U15344 ( .A(n15365), .B(n15400), .Z(n15390) );
  AND U15345 ( .A(n15401), .B(n15402), .Z(n15399) );
  XOR U15346 ( .A(n15403), .B(n15397), .Z(n15401) );
  XNOR U15347 ( .A(n15350), .B(n15393), .Z(n15395) );
  XNOR U15348 ( .A(n15404), .B(n15405), .Z(n15350) );
  AND U15349 ( .A(n523), .B(n15357), .Z(n15405) );
  XOR U15350 ( .A(n15404), .B(n15355), .Z(n15357) );
  XOR U15351 ( .A(n15406), .B(n15407), .Z(n15393) );
  AND U15352 ( .A(n15408), .B(n15409), .Z(n15407) );
  XNOR U15353 ( .A(n15406), .B(n15365), .Z(n15409) );
  XOR U15354 ( .A(n15410), .B(n15402), .Z(n15365) );
  XNOR U15355 ( .A(n15411), .B(n15397), .Z(n15402) );
  XOR U15356 ( .A(n15412), .B(n15413), .Z(n15397) );
  AND U15357 ( .A(n15414), .B(n15415), .Z(n15413) );
  XOR U15358 ( .A(n15416), .B(n15412), .Z(n15414) );
  XNOR U15359 ( .A(n15417), .B(n15418), .Z(n15411) );
  AND U15360 ( .A(n15419), .B(n15420), .Z(n15418) );
  XOR U15361 ( .A(n15417), .B(n15421), .Z(n15419) );
  XNOR U15362 ( .A(n15403), .B(n15400), .Z(n15410) );
  AND U15363 ( .A(n15422), .B(n15423), .Z(n15400) );
  XOR U15364 ( .A(n15424), .B(n15425), .Z(n15403) );
  AND U15365 ( .A(n15426), .B(n15427), .Z(n15425) );
  XOR U15366 ( .A(n15424), .B(n15428), .Z(n15426) );
  XNOR U15367 ( .A(n15362), .B(n15406), .Z(n15408) );
  XNOR U15368 ( .A(n15429), .B(n15430), .Z(n15362) );
  AND U15369 ( .A(n523), .B(n15368), .Z(n15430) );
  XOR U15370 ( .A(n15429), .B(n15366), .Z(n15368) );
  XOR U15371 ( .A(n15431), .B(n15432), .Z(n15406) );
  AND U15372 ( .A(n15433), .B(n15434), .Z(n15432) );
  XNOR U15373 ( .A(n15431), .B(n15422), .Z(n15434) );
  IV U15374 ( .A(n15376), .Z(n15422) );
  XNOR U15375 ( .A(n15435), .B(n15415), .Z(n15376) );
  XNOR U15376 ( .A(n15436), .B(n15421), .Z(n15415) );
  XOR U15377 ( .A(n15437), .B(n15438), .Z(n15421) );
  NOR U15378 ( .A(n15439), .B(n15440), .Z(n15438) );
  XNOR U15379 ( .A(n15437), .B(n15441), .Z(n15439) );
  XNOR U15380 ( .A(n15420), .B(n15412), .Z(n15436) );
  XOR U15381 ( .A(n15442), .B(n15443), .Z(n15412) );
  AND U15382 ( .A(n15444), .B(n15445), .Z(n15443) );
  XNOR U15383 ( .A(n15442), .B(n15446), .Z(n15444) );
  XNOR U15384 ( .A(n15447), .B(n15417), .Z(n15420) );
  XOR U15385 ( .A(n15448), .B(n15449), .Z(n15417) );
  AND U15386 ( .A(n15450), .B(n15451), .Z(n15449) );
  XOR U15387 ( .A(n15448), .B(n15452), .Z(n15450) );
  XNOR U15388 ( .A(n15453), .B(n15454), .Z(n15447) );
  NOR U15389 ( .A(n15455), .B(n15456), .Z(n15454) );
  XOR U15390 ( .A(n15453), .B(n15457), .Z(n15455) );
  XNOR U15391 ( .A(n15416), .B(n15423), .Z(n15435) );
  NOR U15392 ( .A(n15384), .B(n15458), .Z(n15423) );
  XOR U15393 ( .A(n15428), .B(n15427), .Z(n15416) );
  XNOR U15394 ( .A(n15459), .B(n15424), .Z(n15427) );
  XOR U15395 ( .A(n15460), .B(n15461), .Z(n15424) );
  AND U15396 ( .A(n15462), .B(n15463), .Z(n15461) );
  XOR U15397 ( .A(n15460), .B(n15464), .Z(n15462) );
  XNOR U15398 ( .A(n15465), .B(n15466), .Z(n15459) );
  NOR U15399 ( .A(n15467), .B(n15468), .Z(n15466) );
  XNOR U15400 ( .A(n15465), .B(n15469), .Z(n15467) );
  XOR U15401 ( .A(n15470), .B(n15471), .Z(n15428) );
  NOR U15402 ( .A(n15472), .B(n15473), .Z(n15471) );
  XNOR U15403 ( .A(n15470), .B(n15474), .Z(n15472) );
  XNOR U15404 ( .A(n15373), .B(n15431), .Z(n15433) );
  XNOR U15405 ( .A(n15475), .B(n15476), .Z(n15373) );
  AND U15406 ( .A(n523), .B(n15380), .Z(n15476) );
  XOR U15407 ( .A(n15475), .B(n15378), .Z(n15380) );
  AND U15408 ( .A(n15381), .B(n15384), .Z(n15431) );
  XOR U15409 ( .A(n15477), .B(n15458), .Z(n15384) );
  XNOR U15410 ( .A(p_input[1024]), .B(p_input[704]), .Z(n15458) );
  XOR U15411 ( .A(n15446), .B(n15445), .Z(n15477) );
  XNOR U15412 ( .A(n15478), .B(n15452), .Z(n15445) );
  XNOR U15413 ( .A(n15441), .B(n15440), .Z(n15452) );
  XOR U15414 ( .A(n15479), .B(n15437), .Z(n15440) );
  XOR U15415 ( .A(p_input[1034]), .B(p_input[714]), .Z(n15437) );
  XNOR U15416 ( .A(p_input[1035]), .B(p_input[715]), .Z(n15479) );
  XOR U15417 ( .A(p_input[1036]), .B(p_input[716]), .Z(n15441) );
  XNOR U15418 ( .A(n15451), .B(n15442), .Z(n15478) );
  XOR U15419 ( .A(p_input[1025]), .B(p_input[705]), .Z(n15442) );
  XOR U15420 ( .A(n15480), .B(n15457), .Z(n15451) );
  XNOR U15421 ( .A(p_input[1039]), .B(p_input[719]), .Z(n15457) );
  XOR U15422 ( .A(n15448), .B(n15456), .Z(n15480) );
  XOR U15423 ( .A(n15481), .B(n15453), .Z(n15456) );
  XOR U15424 ( .A(p_input[1037]), .B(p_input[717]), .Z(n15453) );
  XNOR U15425 ( .A(p_input[1038]), .B(p_input[718]), .Z(n15481) );
  XOR U15426 ( .A(p_input[1033]), .B(p_input[713]), .Z(n15448) );
  XNOR U15427 ( .A(n15464), .B(n15463), .Z(n15446) );
  XNOR U15428 ( .A(n15482), .B(n15469), .Z(n15463) );
  XOR U15429 ( .A(p_input[1032]), .B(p_input[712]), .Z(n15469) );
  XOR U15430 ( .A(n15460), .B(n15468), .Z(n15482) );
  XOR U15431 ( .A(n15483), .B(n15465), .Z(n15468) );
  XOR U15432 ( .A(p_input[1030]), .B(p_input[710]), .Z(n15465) );
  XNOR U15433 ( .A(p_input[1031]), .B(p_input[711]), .Z(n15483) );
  XOR U15434 ( .A(p_input[1026]), .B(p_input[706]), .Z(n15460) );
  XNOR U15435 ( .A(n15474), .B(n15473), .Z(n15464) );
  XOR U15436 ( .A(n15484), .B(n15470), .Z(n15473) );
  XOR U15437 ( .A(p_input[1027]), .B(p_input[707]), .Z(n15470) );
  XNOR U15438 ( .A(p_input[1028]), .B(p_input[708]), .Z(n15484) );
  XOR U15439 ( .A(p_input[1029]), .B(p_input[709]), .Z(n15474) );
  XNOR U15440 ( .A(n15485), .B(n15486), .Z(n15381) );
  AND U15441 ( .A(n523), .B(n15487), .Z(n15486) );
  XNOR U15442 ( .A(n15488), .B(n15489), .Z(n523) );
  AND U15443 ( .A(n15490), .B(n15491), .Z(n15489) );
  XOR U15444 ( .A(n15488), .B(n15391), .Z(n15491) );
  XNOR U15445 ( .A(n15488), .B(n15345), .Z(n15490) );
  XOR U15446 ( .A(n15492), .B(n15493), .Z(n15488) );
  AND U15447 ( .A(n15494), .B(n15495), .Z(n15493) );
  XOR U15448 ( .A(n15492), .B(n15355), .Z(n15494) );
  XOR U15449 ( .A(n15496), .B(n15497), .Z(n15334) );
  AND U15450 ( .A(n527), .B(n15487), .Z(n15497) );
  XNOR U15451 ( .A(n15485), .B(n15496), .Z(n15487) );
  XNOR U15452 ( .A(n15498), .B(n15499), .Z(n527) );
  AND U15453 ( .A(n15500), .B(n15501), .Z(n15499) );
  XNOR U15454 ( .A(n15502), .B(n15498), .Z(n15501) );
  IV U15455 ( .A(n15391), .Z(n15502) );
  XNOR U15456 ( .A(n15503), .B(n15504), .Z(n15391) );
  AND U15457 ( .A(n530), .B(n15505), .Z(n15504) );
  XNOR U15458 ( .A(n15503), .B(n15506), .Z(n15505) );
  XNOR U15459 ( .A(n15345), .B(n15498), .Z(n15500) );
  XOR U15460 ( .A(n15507), .B(n15508), .Z(n15345) );
  AND U15461 ( .A(n538), .B(n15509), .Z(n15508) );
  XOR U15462 ( .A(n15492), .B(n15510), .Z(n15498) );
  AND U15463 ( .A(n15511), .B(n15495), .Z(n15510) );
  XNOR U15464 ( .A(n15404), .B(n15492), .Z(n15495) );
  XNOR U15465 ( .A(n15512), .B(n15513), .Z(n15404) );
  AND U15466 ( .A(n530), .B(n15514), .Z(n15513) );
  XOR U15467 ( .A(n15515), .B(n15512), .Z(n15514) );
  XNOR U15468 ( .A(n15516), .B(n15492), .Z(n15511) );
  IV U15469 ( .A(n15355), .Z(n15516) );
  XOR U15470 ( .A(n15517), .B(n15518), .Z(n15355) );
  AND U15471 ( .A(n538), .B(n15519), .Z(n15518) );
  XOR U15472 ( .A(n15520), .B(n15521), .Z(n15492) );
  AND U15473 ( .A(n15522), .B(n15523), .Z(n15521) );
  XNOR U15474 ( .A(n15429), .B(n15520), .Z(n15523) );
  XNOR U15475 ( .A(n15524), .B(n15525), .Z(n15429) );
  AND U15476 ( .A(n530), .B(n15526), .Z(n15525) );
  XNOR U15477 ( .A(n15527), .B(n15524), .Z(n15526) );
  XOR U15478 ( .A(n15520), .B(n15366), .Z(n15522) );
  XOR U15479 ( .A(n15528), .B(n15529), .Z(n15366) );
  AND U15480 ( .A(n538), .B(n15530), .Z(n15529) );
  XOR U15481 ( .A(n15531), .B(n15532), .Z(n15520) );
  AND U15482 ( .A(n15533), .B(n15534), .Z(n15532) );
  XNOR U15483 ( .A(n15531), .B(n15475), .Z(n15534) );
  XNOR U15484 ( .A(n15535), .B(n15536), .Z(n15475) );
  AND U15485 ( .A(n530), .B(n15537), .Z(n15536) );
  XOR U15486 ( .A(n15538), .B(n15535), .Z(n15537) );
  XNOR U15487 ( .A(n15539), .B(n15531), .Z(n15533) );
  IV U15488 ( .A(n15378), .Z(n15539) );
  XOR U15489 ( .A(n15540), .B(n15541), .Z(n15378) );
  AND U15490 ( .A(n538), .B(n15542), .Z(n15541) );
  AND U15491 ( .A(n15496), .B(n15485), .Z(n15531) );
  XNOR U15492 ( .A(n15543), .B(n15544), .Z(n15485) );
  AND U15493 ( .A(n530), .B(n15545), .Z(n15544) );
  XNOR U15494 ( .A(n15546), .B(n15543), .Z(n15545) );
  XNOR U15495 ( .A(n15547), .B(n15548), .Z(n530) );
  AND U15496 ( .A(n15549), .B(n15550), .Z(n15548) );
  XOR U15497 ( .A(n15506), .B(n15547), .Z(n15550) );
  AND U15498 ( .A(n15551), .B(n15552), .Z(n15506) );
  XOR U15499 ( .A(n15547), .B(n15503), .Z(n15549) );
  XNOR U15500 ( .A(n15553), .B(n15554), .Z(n15503) );
  AND U15501 ( .A(n534), .B(n15509), .Z(n15554) );
  XOR U15502 ( .A(n15507), .B(n15553), .Z(n15509) );
  XOR U15503 ( .A(n15555), .B(n15556), .Z(n15547) );
  AND U15504 ( .A(n15557), .B(n15558), .Z(n15556) );
  XNOR U15505 ( .A(n15555), .B(n15551), .Z(n15558) );
  IV U15506 ( .A(n15515), .Z(n15551) );
  XOR U15507 ( .A(n15559), .B(n15560), .Z(n15515) );
  XOR U15508 ( .A(n15561), .B(n15552), .Z(n15560) );
  AND U15509 ( .A(n15527), .B(n15562), .Z(n15552) );
  AND U15510 ( .A(n15563), .B(n15564), .Z(n15561) );
  XOR U15511 ( .A(n15565), .B(n15559), .Z(n15563) );
  XNOR U15512 ( .A(n15512), .B(n15555), .Z(n15557) );
  XNOR U15513 ( .A(n15566), .B(n15567), .Z(n15512) );
  AND U15514 ( .A(n534), .B(n15519), .Z(n15567) );
  XOR U15515 ( .A(n15566), .B(n15517), .Z(n15519) );
  XOR U15516 ( .A(n15568), .B(n15569), .Z(n15555) );
  AND U15517 ( .A(n15570), .B(n15571), .Z(n15569) );
  XNOR U15518 ( .A(n15568), .B(n15527), .Z(n15571) );
  XOR U15519 ( .A(n15572), .B(n15564), .Z(n15527) );
  XNOR U15520 ( .A(n15573), .B(n15559), .Z(n15564) );
  XOR U15521 ( .A(n15574), .B(n15575), .Z(n15559) );
  AND U15522 ( .A(n15576), .B(n15577), .Z(n15575) );
  XOR U15523 ( .A(n15578), .B(n15574), .Z(n15576) );
  XNOR U15524 ( .A(n15579), .B(n15580), .Z(n15573) );
  AND U15525 ( .A(n15581), .B(n15582), .Z(n15580) );
  XOR U15526 ( .A(n15579), .B(n15583), .Z(n15581) );
  XNOR U15527 ( .A(n15565), .B(n15562), .Z(n15572) );
  AND U15528 ( .A(n15584), .B(n15585), .Z(n15562) );
  XOR U15529 ( .A(n15586), .B(n15587), .Z(n15565) );
  AND U15530 ( .A(n15588), .B(n15589), .Z(n15587) );
  XOR U15531 ( .A(n15586), .B(n15590), .Z(n15588) );
  XNOR U15532 ( .A(n15524), .B(n15568), .Z(n15570) );
  XNOR U15533 ( .A(n15591), .B(n15592), .Z(n15524) );
  AND U15534 ( .A(n534), .B(n15530), .Z(n15592) );
  XOR U15535 ( .A(n15591), .B(n15528), .Z(n15530) );
  XOR U15536 ( .A(n15593), .B(n15594), .Z(n15568) );
  AND U15537 ( .A(n15595), .B(n15596), .Z(n15594) );
  XNOR U15538 ( .A(n15593), .B(n15584), .Z(n15596) );
  IV U15539 ( .A(n15538), .Z(n15584) );
  XNOR U15540 ( .A(n15597), .B(n15577), .Z(n15538) );
  XNOR U15541 ( .A(n15598), .B(n15583), .Z(n15577) );
  XOR U15542 ( .A(n15599), .B(n15600), .Z(n15583) );
  NOR U15543 ( .A(n15601), .B(n15602), .Z(n15600) );
  XNOR U15544 ( .A(n15599), .B(n15603), .Z(n15601) );
  XNOR U15545 ( .A(n15582), .B(n15574), .Z(n15598) );
  XOR U15546 ( .A(n15604), .B(n15605), .Z(n15574) );
  AND U15547 ( .A(n15606), .B(n15607), .Z(n15605) );
  XNOR U15548 ( .A(n15604), .B(n15608), .Z(n15606) );
  XNOR U15549 ( .A(n15609), .B(n15579), .Z(n15582) );
  XOR U15550 ( .A(n15610), .B(n15611), .Z(n15579) );
  AND U15551 ( .A(n15612), .B(n15613), .Z(n15611) );
  XOR U15552 ( .A(n15610), .B(n15614), .Z(n15612) );
  XNOR U15553 ( .A(n15615), .B(n15616), .Z(n15609) );
  NOR U15554 ( .A(n15617), .B(n15618), .Z(n15616) );
  XOR U15555 ( .A(n15615), .B(n15619), .Z(n15617) );
  XNOR U15556 ( .A(n15578), .B(n15585), .Z(n15597) );
  NOR U15557 ( .A(n15546), .B(n15620), .Z(n15585) );
  XOR U15558 ( .A(n15590), .B(n15589), .Z(n15578) );
  XNOR U15559 ( .A(n15621), .B(n15586), .Z(n15589) );
  XOR U15560 ( .A(n15622), .B(n15623), .Z(n15586) );
  AND U15561 ( .A(n15624), .B(n15625), .Z(n15623) );
  XOR U15562 ( .A(n15622), .B(n15626), .Z(n15624) );
  XNOR U15563 ( .A(n15627), .B(n15628), .Z(n15621) );
  NOR U15564 ( .A(n15629), .B(n15630), .Z(n15628) );
  XNOR U15565 ( .A(n15627), .B(n15631), .Z(n15629) );
  XOR U15566 ( .A(n15632), .B(n15633), .Z(n15590) );
  NOR U15567 ( .A(n15634), .B(n15635), .Z(n15633) );
  XNOR U15568 ( .A(n15632), .B(n15636), .Z(n15634) );
  XNOR U15569 ( .A(n15535), .B(n15593), .Z(n15595) );
  XNOR U15570 ( .A(n15637), .B(n15638), .Z(n15535) );
  AND U15571 ( .A(n534), .B(n15542), .Z(n15638) );
  XOR U15572 ( .A(n15637), .B(n15540), .Z(n15542) );
  AND U15573 ( .A(n15543), .B(n15546), .Z(n15593) );
  XOR U15574 ( .A(n15639), .B(n15620), .Z(n15546) );
  XNOR U15575 ( .A(p_input[1024]), .B(p_input[720]), .Z(n15620) );
  XOR U15576 ( .A(n15608), .B(n15607), .Z(n15639) );
  XNOR U15577 ( .A(n15640), .B(n15614), .Z(n15607) );
  XNOR U15578 ( .A(n15603), .B(n15602), .Z(n15614) );
  XOR U15579 ( .A(n15641), .B(n15599), .Z(n15602) );
  XOR U15580 ( .A(p_input[1034]), .B(p_input[730]), .Z(n15599) );
  XNOR U15581 ( .A(p_input[1035]), .B(p_input[731]), .Z(n15641) );
  XOR U15582 ( .A(p_input[1036]), .B(p_input[732]), .Z(n15603) );
  XNOR U15583 ( .A(n15613), .B(n15604), .Z(n15640) );
  XOR U15584 ( .A(p_input[1025]), .B(p_input[721]), .Z(n15604) );
  XOR U15585 ( .A(n15642), .B(n15619), .Z(n15613) );
  XNOR U15586 ( .A(p_input[1039]), .B(p_input[735]), .Z(n15619) );
  XOR U15587 ( .A(n15610), .B(n15618), .Z(n15642) );
  XOR U15588 ( .A(n15643), .B(n15615), .Z(n15618) );
  XOR U15589 ( .A(p_input[1037]), .B(p_input[733]), .Z(n15615) );
  XNOR U15590 ( .A(p_input[1038]), .B(p_input[734]), .Z(n15643) );
  XOR U15591 ( .A(p_input[1033]), .B(p_input[729]), .Z(n15610) );
  XNOR U15592 ( .A(n15626), .B(n15625), .Z(n15608) );
  XNOR U15593 ( .A(n15644), .B(n15631), .Z(n15625) );
  XOR U15594 ( .A(p_input[1032]), .B(p_input[728]), .Z(n15631) );
  XOR U15595 ( .A(n15622), .B(n15630), .Z(n15644) );
  XOR U15596 ( .A(n15645), .B(n15627), .Z(n15630) );
  XOR U15597 ( .A(p_input[1030]), .B(p_input[726]), .Z(n15627) );
  XNOR U15598 ( .A(p_input[1031]), .B(p_input[727]), .Z(n15645) );
  XOR U15599 ( .A(p_input[1026]), .B(p_input[722]), .Z(n15622) );
  XNOR U15600 ( .A(n15636), .B(n15635), .Z(n15626) );
  XOR U15601 ( .A(n15646), .B(n15632), .Z(n15635) );
  XOR U15602 ( .A(p_input[1027]), .B(p_input[723]), .Z(n15632) );
  XNOR U15603 ( .A(p_input[1028]), .B(p_input[724]), .Z(n15646) );
  XOR U15604 ( .A(p_input[1029]), .B(p_input[725]), .Z(n15636) );
  XNOR U15605 ( .A(n15647), .B(n15648), .Z(n15543) );
  AND U15606 ( .A(n534), .B(n15649), .Z(n15648) );
  XNOR U15607 ( .A(n15650), .B(n15651), .Z(n534) );
  AND U15608 ( .A(n15652), .B(n15653), .Z(n15651) );
  XOR U15609 ( .A(n15650), .B(n15553), .Z(n15653) );
  XNOR U15610 ( .A(n15650), .B(n15507), .Z(n15652) );
  XOR U15611 ( .A(n15654), .B(n15655), .Z(n15650) );
  AND U15612 ( .A(n15656), .B(n15657), .Z(n15655) );
  XOR U15613 ( .A(n15654), .B(n15517), .Z(n15656) );
  XOR U15614 ( .A(n15658), .B(n15659), .Z(n15496) );
  AND U15615 ( .A(n538), .B(n15649), .Z(n15659) );
  XNOR U15616 ( .A(n15647), .B(n15658), .Z(n15649) );
  XNOR U15617 ( .A(n15660), .B(n15661), .Z(n538) );
  AND U15618 ( .A(n15662), .B(n15663), .Z(n15661) );
  XNOR U15619 ( .A(n15664), .B(n15660), .Z(n15663) );
  IV U15620 ( .A(n15553), .Z(n15664) );
  XNOR U15621 ( .A(n15665), .B(n15666), .Z(n15553) );
  AND U15622 ( .A(n541), .B(n15667), .Z(n15666) );
  XNOR U15623 ( .A(n15665), .B(n15668), .Z(n15667) );
  XNOR U15624 ( .A(n15507), .B(n15660), .Z(n15662) );
  XOR U15625 ( .A(n15669), .B(n15670), .Z(n15507) );
  AND U15626 ( .A(n549), .B(n15671), .Z(n15670) );
  XOR U15627 ( .A(n15654), .B(n15672), .Z(n15660) );
  AND U15628 ( .A(n15673), .B(n15657), .Z(n15672) );
  XNOR U15629 ( .A(n15566), .B(n15654), .Z(n15657) );
  XNOR U15630 ( .A(n15674), .B(n15675), .Z(n15566) );
  AND U15631 ( .A(n541), .B(n15676), .Z(n15675) );
  XOR U15632 ( .A(n15677), .B(n15674), .Z(n15676) );
  XNOR U15633 ( .A(n15678), .B(n15654), .Z(n15673) );
  IV U15634 ( .A(n15517), .Z(n15678) );
  XOR U15635 ( .A(n15679), .B(n15680), .Z(n15517) );
  AND U15636 ( .A(n549), .B(n15681), .Z(n15680) );
  XOR U15637 ( .A(n15682), .B(n15683), .Z(n15654) );
  AND U15638 ( .A(n15684), .B(n15685), .Z(n15683) );
  XNOR U15639 ( .A(n15591), .B(n15682), .Z(n15685) );
  XNOR U15640 ( .A(n15686), .B(n15687), .Z(n15591) );
  AND U15641 ( .A(n541), .B(n15688), .Z(n15687) );
  XNOR U15642 ( .A(n15689), .B(n15686), .Z(n15688) );
  XOR U15643 ( .A(n15682), .B(n15528), .Z(n15684) );
  XOR U15644 ( .A(n15690), .B(n15691), .Z(n15528) );
  AND U15645 ( .A(n549), .B(n15692), .Z(n15691) );
  XOR U15646 ( .A(n15693), .B(n15694), .Z(n15682) );
  AND U15647 ( .A(n15695), .B(n15696), .Z(n15694) );
  XNOR U15648 ( .A(n15693), .B(n15637), .Z(n15696) );
  XNOR U15649 ( .A(n15697), .B(n15698), .Z(n15637) );
  AND U15650 ( .A(n541), .B(n15699), .Z(n15698) );
  XOR U15651 ( .A(n15700), .B(n15697), .Z(n15699) );
  XNOR U15652 ( .A(n15701), .B(n15693), .Z(n15695) );
  IV U15653 ( .A(n15540), .Z(n15701) );
  XOR U15654 ( .A(n15702), .B(n15703), .Z(n15540) );
  AND U15655 ( .A(n549), .B(n15704), .Z(n15703) );
  AND U15656 ( .A(n15658), .B(n15647), .Z(n15693) );
  XNOR U15657 ( .A(n15705), .B(n15706), .Z(n15647) );
  AND U15658 ( .A(n541), .B(n15707), .Z(n15706) );
  XNOR U15659 ( .A(n15708), .B(n15705), .Z(n15707) );
  XNOR U15660 ( .A(n15709), .B(n15710), .Z(n541) );
  AND U15661 ( .A(n15711), .B(n15712), .Z(n15710) );
  XOR U15662 ( .A(n15668), .B(n15709), .Z(n15712) );
  AND U15663 ( .A(n15713), .B(n15714), .Z(n15668) );
  XOR U15664 ( .A(n15709), .B(n15665), .Z(n15711) );
  XNOR U15665 ( .A(n15715), .B(n15716), .Z(n15665) );
  AND U15666 ( .A(n545), .B(n15671), .Z(n15716) );
  XOR U15667 ( .A(n15669), .B(n15715), .Z(n15671) );
  XOR U15668 ( .A(n15717), .B(n15718), .Z(n15709) );
  AND U15669 ( .A(n15719), .B(n15720), .Z(n15718) );
  XNOR U15670 ( .A(n15717), .B(n15713), .Z(n15720) );
  IV U15671 ( .A(n15677), .Z(n15713) );
  XOR U15672 ( .A(n15721), .B(n15722), .Z(n15677) );
  XOR U15673 ( .A(n15723), .B(n15714), .Z(n15722) );
  AND U15674 ( .A(n15689), .B(n15724), .Z(n15714) );
  AND U15675 ( .A(n15725), .B(n15726), .Z(n15723) );
  XOR U15676 ( .A(n15727), .B(n15721), .Z(n15725) );
  XNOR U15677 ( .A(n15674), .B(n15717), .Z(n15719) );
  XNOR U15678 ( .A(n15728), .B(n15729), .Z(n15674) );
  AND U15679 ( .A(n545), .B(n15681), .Z(n15729) );
  XOR U15680 ( .A(n15728), .B(n15679), .Z(n15681) );
  XOR U15681 ( .A(n15730), .B(n15731), .Z(n15717) );
  AND U15682 ( .A(n15732), .B(n15733), .Z(n15731) );
  XNOR U15683 ( .A(n15730), .B(n15689), .Z(n15733) );
  XOR U15684 ( .A(n15734), .B(n15726), .Z(n15689) );
  XNOR U15685 ( .A(n15735), .B(n15721), .Z(n15726) );
  XOR U15686 ( .A(n15736), .B(n15737), .Z(n15721) );
  AND U15687 ( .A(n15738), .B(n15739), .Z(n15737) );
  XOR U15688 ( .A(n15740), .B(n15736), .Z(n15738) );
  XNOR U15689 ( .A(n15741), .B(n15742), .Z(n15735) );
  AND U15690 ( .A(n15743), .B(n15744), .Z(n15742) );
  XOR U15691 ( .A(n15741), .B(n15745), .Z(n15743) );
  XNOR U15692 ( .A(n15727), .B(n15724), .Z(n15734) );
  AND U15693 ( .A(n15746), .B(n15747), .Z(n15724) );
  XOR U15694 ( .A(n15748), .B(n15749), .Z(n15727) );
  AND U15695 ( .A(n15750), .B(n15751), .Z(n15749) );
  XOR U15696 ( .A(n15748), .B(n15752), .Z(n15750) );
  XNOR U15697 ( .A(n15686), .B(n15730), .Z(n15732) );
  XNOR U15698 ( .A(n15753), .B(n15754), .Z(n15686) );
  AND U15699 ( .A(n545), .B(n15692), .Z(n15754) );
  XOR U15700 ( .A(n15753), .B(n15690), .Z(n15692) );
  XOR U15701 ( .A(n15755), .B(n15756), .Z(n15730) );
  AND U15702 ( .A(n15757), .B(n15758), .Z(n15756) );
  XNOR U15703 ( .A(n15755), .B(n15746), .Z(n15758) );
  IV U15704 ( .A(n15700), .Z(n15746) );
  XNOR U15705 ( .A(n15759), .B(n15739), .Z(n15700) );
  XNOR U15706 ( .A(n15760), .B(n15745), .Z(n15739) );
  XOR U15707 ( .A(n15761), .B(n15762), .Z(n15745) );
  NOR U15708 ( .A(n15763), .B(n15764), .Z(n15762) );
  XNOR U15709 ( .A(n15761), .B(n15765), .Z(n15763) );
  XNOR U15710 ( .A(n15744), .B(n15736), .Z(n15760) );
  XOR U15711 ( .A(n15766), .B(n15767), .Z(n15736) );
  AND U15712 ( .A(n15768), .B(n15769), .Z(n15767) );
  XNOR U15713 ( .A(n15766), .B(n15770), .Z(n15768) );
  XNOR U15714 ( .A(n15771), .B(n15741), .Z(n15744) );
  XOR U15715 ( .A(n15772), .B(n15773), .Z(n15741) );
  AND U15716 ( .A(n15774), .B(n15775), .Z(n15773) );
  XOR U15717 ( .A(n15772), .B(n15776), .Z(n15774) );
  XNOR U15718 ( .A(n15777), .B(n15778), .Z(n15771) );
  NOR U15719 ( .A(n15779), .B(n15780), .Z(n15778) );
  XOR U15720 ( .A(n15777), .B(n15781), .Z(n15779) );
  XNOR U15721 ( .A(n15740), .B(n15747), .Z(n15759) );
  NOR U15722 ( .A(n15708), .B(n15782), .Z(n15747) );
  XOR U15723 ( .A(n15752), .B(n15751), .Z(n15740) );
  XNOR U15724 ( .A(n15783), .B(n15748), .Z(n15751) );
  XOR U15725 ( .A(n15784), .B(n15785), .Z(n15748) );
  AND U15726 ( .A(n15786), .B(n15787), .Z(n15785) );
  XOR U15727 ( .A(n15784), .B(n15788), .Z(n15786) );
  XNOR U15728 ( .A(n15789), .B(n15790), .Z(n15783) );
  NOR U15729 ( .A(n15791), .B(n15792), .Z(n15790) );
  XNOR U15730 ( .A(n15789), .B(n15793), .Z(n15791) );
  XOR U15731 ( .A(n15794), .B(n15795), .Z(n15752) );
  NOR U15732 ( .A(n15796), .B(n15797), .Z(n15795) );
  XNOR U15733 ( .A(n15794), .B(n15798), .Z(n15796) );
  XNOR U15734 ( .A(n15697), .B(n15755), .Z(n15757) );
  XNOR U15735 ( .A(n15799), .B(n15800), .Z(n15697) );
  AND U15736 ( .A(n545), .B(n15704), .Z(n15800) );
  XOR U15737 ( .A(n15799), .B(n15702), .Z(n15704) );
  AND U15738 ( .A(n15705), .B(n15708), .Z(n15755) );
  XOR U15739 ( .A(n15801), .B(n15782), .Z(n15708) );
  XNOR U15740 ( .A(p_input[1024]), .B(p_input[736]), .Z(n15782) );
  XOR U15741 ( .A(n15770), .B(n15769), .Z(n15801) );
  XNOR U15742 ( .A(n15802), .B(n15776), .Z(n15769) );
  XNOR U15743 ( .A(n15765), .B(n15764), .Z(n15776) );
  XOR U15744 ( .A(n15803), .B(n15761), .Z(n15764) );
  XOR U15745 ( .A(p_input[1034]), .B(p_input[746]), .Z(n15761) );
  XNOR U15746 ( .A(p_input[1035]), .B(p_input[747]), .Z(n15803) );
  XOR U15747 ( .A(p_input[1036]), .B(p_input[748]), .Z(n15765) );
  XNOR U15748 ( .A(n15775), .B(n15766), .Z(n15802) );
  XOR U15749 ( .A(p_input[1025]), .B(p_input[737]), .Z(n15766) );
  XOR U15750 ( .A(n15804), .B(n15781), .Z(n15775) );
  XNOR U15751 ( .A(p_input[1039]), .B(p_input[751]), .Z(n15781) );
  XOR U15752 ( .A(n15772), .B(n15780), .Z(n15804) );
  XOR U15753 ( .A(n15805), .B(n15777), .Z(n15780) );
  XOR U15754 ( .A(p_input[1037]), .B(p_input[749]), .Z(n15777) );
  XNOR U15755 ( .A(p_input[1038]), .B(p_input[750]), .Z(n15805) );
  XOR U15756 ( .A(p_input[1033]), .B(p_input[745]), .Z(n15772) );
  XNOR U15757 ( .A(n15788), .B(n15787), .Z(n15770) );
  XNOR U15758 ( .A(n15806), .B(n15793), .Z(n15787) );
  XOR U15759 ( .A(p_input[1032]), .B(p_input[744]), .Z(n15793) );
  XOR U15760 ( .A(n15784), .B(n15792), .Z(n15806) );
  XOR U15761 ( .A(n15807), .B(n15789), .Z(n15792) );
  XOR U15762 ( .A(p_input[1030]), .B(p_input[742]), .Z(n15789) );
  XNOR U15763 ( .A(p_input[1031]), .B(p_input[743]), .Z(n15807) );
  XOR U15764 ( .A(p_input[1026]), .B(p_input[738]), .Z(n15784) );
  XNOR U15765 ( .A(n15798), .B(n15797), .Z(n15788) );
  XOR U15766 ( .A(n15808), .B(n15794), .Z(n15797) );
  XOR U15767 ( .A(p_input[1027]), .B(p_input[739]), .Z(n15794) );
  XNOR U15768 ( .A(p_input[1028]), .B(p_input[740]), .Z(n15808) );
  XOR U15769 ( .A(p_input[1029]), .B(p_input[741]), .Z(n15798) );
  XNOR U15770 ( .A(n15809), .B(n15810), .Z(n15705) );
  AND U15771 ( .A(n545), .B(n15811), .Z(n15810) );
  XNOR U15772 ( .A(n15812), .B(n15813), .Z(n545) );
  AND U15773 ( .A(n15814), .B(n15815), .Z(n15813) );
  XOR U15774 ( .A(n15812), .B(n15715), .Z(n15815) );
  XNOR U15775 ( .A(n15812), .B(n15669), .Z(n15814) );
  XOR U15776 ( .A(n15816), .B(n15817), .Z(n15812) );
  AND U15777 ( .A(n15818), .B(n15819), .Z(n15817) );
  XOR U15778 ( .A(n15816), .B(n15679), .Z(n15818) );
  XOR U15779 ( .A(n15820), .B(n15821), .Z(n15658) );
  AND U15780 ( .A(n549), .B(n15811), .Z(n15821) );
  XNOR U15781 ( .A(n15809), .B(n15820), .Z(n15811) );
  XNOR U15782 ( .A(n15822), .B(n15823), .Z(n549) );
  AND U15783 ( .A(n15824), .B(n15825), .Z(n15823) );
  XNOR U15784 ( .A(n15826), .B(n15822), .Z(n15825) );
  IV U15785 ( .A(n15715), .Z(n15826) );
  XNOR U15786 ( .A(n15827), .B(n15828), .Z(n15715) );
  AND U15787 ( .A(n552), .B(n15829), .Z(n15828) );
  XNOR U15788 ( .A(n15827), .B(n15830), .Z(n15829) );
  XNOR U15789 ( .A(n15669), .B(n15822), .Z(n15824) );
  XOR U15790 ( .A(n15831), .B(n15832), .Z(n15669) );
  AND U15791 ( .A(n560), .B(n15833), .Z(n15832) );
  XOR U15792 ( .A(n15816), .B(n15834), .Z(n15822) );
  AND U15793 ( .A(n15835), .B(n15819), .Z(n15834) );
  XNOR U15794 ( .A(n15728), .B(n15816), .Z(n15819) );
  XNOR U15795 ( .A(n15836), .B(n15837), .Z(n15728) );
  AND U15796 ( .A(n552), .B(n15838), .Z(n15837) );
  XOR U15797 ( .A(n15839), .B(n15836), .Z(n15838) );
  XNOR U15798 ( .A(n15840), .B(n15816), .Z(n15835) );
  IV U15799 ( .A(n15679), .Z(n15840) );
  XOR U15800 ( .A(n15841), .B(n15842), .Z(n15679) );
  AND U15801 ( .A(n560), .B(n15843), .Z(n15842) );
  XOR U15802 ( .A(n15844), .B(n15845), .Z(n15816) );
  AND U15803 ( .A(n15846), .B(n15847), .Z(n15845) );
  XNOR U15804 ( .A(n15753), .B(n15844), .Z(n15847) );
  XNOR U15805 ( .A(n15848), .B(n15849), .Z(n15753) );
  AND U15806 ( .A(n552), .B(n15850), .Z(n15849) );
  XNOR U15807 ( .A(n15851), .B(n15848), .Z(n15850) );
  XOR U15808 ( .A(n15844), .B(n15690), .Z(n15846) );
  XOR U15809 ( .A(n15852), .B(n15853), .Z(n15690) );
  AND U15810 ( .A(n560), .B(n15854), .Z(n15853) );
  XOR U15811 ( .A(n15855), .B(n15856), .Z(n15844) );
  AND U15812 ( .A(n15857), .B(n15858), .Z(n15856) );
  XNOR U15813 ( .A(n15855), .B(n15799), .Z(n15858) );
  XNOR U15814 ( .A(n15859), .B(n15860), .Z(n15799) );
  AND U15815 ( .A(n552), .B(n15861), .Z(n15860) );
  XOR U15816 ( .A(n15862), .B(n15859), .Z(n15861) );
  XNOR U15817 ( .A(n15863), .B(n15855), .Z(n15857) );
  IV U15818 ( .A(n15702), .Z(n15863) );
  XOR U15819 ( .A(n15864), .B(n15865), .Z(n15702) );
  AND U15820 ( .A(n560), .B(n15866), .Z(n15865) );
  AND U15821 ( .A(n15820), .B(n15809), .Z(n15855) );
  XNOR U15822 ( .A(n15867), .B(n15868), .Z(n15809) );
  AND U15823 ( .A(n552), .B(n15869), .Z(n15868) );
  XNOR U15824 ( .A(n15870), .B(n15867), .Z(n15869) );
  XNOR U15825 ( .A(n15871), .B(n15872), .Z(n552) );
  AND U15826 ( .A(n15873), .B(n15874), .Z(n15872) );
  XOR U15827 ( .A(n15830), .B(n15871), .Z(n15874) );
  AND U15828 ( .A(n15875), .B(n15876), .Z(n15830) );
  XOR U15829 ( .A(n15871), .B(n15827), .Z(n15873) );
  XNOR U15830 ( .A(n15877), .B(n15878), .Z(n15827) );
  AND U15831 ( .A(n556), .B(n15833), .Z(n15878) );
  XOR U15832 ( .A(n15831), .B(n15877), .Z(n15833) );
  XOR U15833 ( .A(n15879), .B(n15880), .Z(n15871) );
  AND U15834 ( .A(n15881), .B(n15882), .Z(n15880) );
  XNOR U15835 ( .A(n15879), .B(n15875), .Z(n15882) );
  IV U15836 ( .A(n15839), .Z(n15875) );
  XOR U15837 ( .A(n15883), .B(n15884), .Z(n15839) );
  XOR U15838 ( .A(n15885), .B(n15876), .Z(n15884) );
  AND U15839 ( .A(n15851), .B(n15886), .Z(n15876) );
  AND U15840 ( .A(n15887), .B(n15888), .Z(n15885) );
  XOR U15841 ( .A(n15889), .B(n15883), .Z(n15887) );
  XNOR U15842 ( .A(n15836), .B(n15879), .Z(n15881) );
  XNOR U15843 ( .A(n15890), .B(n15891), .Z(n15836) );
  AND U15844 ( .A(n556), .B(n15843), .Z(n15891) );
  XOR U15845 ( .A(n15890), .B(n15841), .Z(n15843) );
  XOR U15846 ( .A(n15892), .B(n15893), .Z(n15879) );
  AND U15847 ( .A(n15894), .B(n15895), .Z(n15893) );
  XNOR U15848 ( .A(n15892), .B(n15851), .Z(n15895) );
  XOR U15849 ( .A(n15896), .B(n15888), .Z(n15851) );
  XNOR U15850 ( .A(n15897), .B(n15883), .Z(n15888) );
  XOR U15851 ( .A(n15898), .B(n15899), .Z(n15883) );
  AND U15852 ( .A(n15900), .B(n15901), .Z(n15899) );
  XOR U15853 ( .A(n15902), .B(n15898), .Z(n15900) );
  XNOR U15854 ( .A(n15903), .B(n15904), .Z(n15897) );
  AND U15855 ( .A(n15905), .B(n15906), .Z(n15904) );
  XOR U15856 ( .A(n15903), .B(n15907), .Z(n15905) );
  XNOR U15857 ( .A(n15889), .B(n15886), .Z(n15896) );
  AND U15858 ( .A(n15908), .B(n15909), .Z(n15886) );
  XOR U15859 ( .A(n15910), .B(n15911), .Z(n15889) );
  AND U15860 ( .A(n15912), .B(n15913), .Z(n15911) );
  XOR U15861 ( .A(n15910), .B(n15914), .Z(n15912) );
  XNOR U15862 ( .A(n15848), .B(n15892), .Z(n15894) );
  XNOR U15863 ( .A(n15915), .B(n15916), .Z(n15848) );
  AND U15864 ( .A(n556), .B(n15854), .Z(n15916) );
  XOR U15865 ( .A(n15915), .B(n15852), .Z(n15854) );
  XOR U15866 ( .A(n15917), .B(n15918), .Z(n15892) );
  AND U15867 ( .A(n15919), .B(n15920), .Z(n15918) );
  XNOR U15868 ( .A(n15917), .B(n15908), .Z(n15920) );
  IV U15869 ( .A(n15862), .Z(n15908) );
  XNOR U15870 ( .A(n15921), .B(n15901), .Z(n15862) );
  XNOR U15871 ( .A(n15922), .B(n15907), .Z(n15901) );
  XOR U15872 ( .A(n15923), .B(n15924), .Z(n15907) );
  NOR U15873 ( .A(n15925), .B(n15926), .Z(n15924) );
  XNOR U15874 ( .A(n15923), .B(n15927), .Z(n15925) );
  XNOR U15875 ( .A(n15906), .B(n15898), .Z(n15922) );
  XOR U15876 ( .A(n15928), .B(n15929), .Z(n15898) );
  AND U15877 ( .A(n15930), .B(n15931), .Z(n15929) );
  XNOR U15878 ( .A(n15928), .B(n15932), .Z(n15930) );
  XNOR U15879 ( .A(n15933), .B(n15903), .Z(n15906) );
  XOR U15880 ( .A(n15934), .B(n15935), .Z(n15903) );
  AND U15881 ( .A(n15936), .B(n15937), .Z(n15935) );
  XOR U15882 ( .A(n15934), .B(n15938), .Z(n15936) );
  XNOR U15883 ( .A(n15939), .B(n15940), .Z(n15933) );
  NOR U15884 ( .A(n15941), .B(n15942), .Z(n15940) );
  XOR U15885 ( .A(n15939), .B(n15943), .Z(n15941) );
  XNOR U15886 ( .A(n15902), .B(n15909), .Z(n15921) );
  NOR U15887 ( .A(n15870), .B(n15944), .Z(n15909) );
  XOR U15888 ( .A(n15914), .B(n15913), .Z(n15902) );
  XNOR U15889 ( .A(n15945), .B(n15910), .Z(n15913) );
  XOR U15890 ( .A(n15946), .B(n15947), .Z(n15910) );
  AND U15891 ( .A(n15948), .B(n15949), .Z(n15947) );
  XOR U15892 ( .A(n15946), .B(n15950), .Z(n15948) );
  XNOR U15893 ( .A(n15951), .B(n15952), .Z(n15945) );
  NOR U15894 ( .A(n15953), .B(n15954), .Z(n15952) );
  XNOR U15895 ( .A(n15951), .B(n15955), .Z(n15953) );
  XOR U15896 ( .A(n15956), .B(n15957), .Z(n15914) );
  NOR U15897 ( .A(n15958), .B(n15959), .Z(n15957) );
  XNOR U15898 ( .A(n15956), .B(n15960), .Z(n15958) );
  XNOR U15899 ( .A(n15859), .B(n15917), .Z(n15919) );
  XNOR U15900 ( .A(n15961), .B(n15962), .Z(n15859) );
  AND U15901 ( .A(n556), .B(n15866), .Z(n15962) );
  XOR U15902 ( .A(n15961), .B(n15864), .Z(n15866) );
  AND U15903 ( .A(n15867), .B(n15870), .Z(n15917) );
  XOR U15904 ( .A(n15963), .B(n15944), .Z(n15870) );
  XNOR U15905 ( .A(p_input[1024]), .B(p_input[752]), .Z(n15944) );
  XOR U15906 ( .A(n15932), .B(n15931), .Z(n15963) );
  XNOR U15907 ( .A(n15964), .B(n15938), .Z(n15931) );
  XNOR U15908 ( .A(n15927), .B(n15926), .Z(n15938) );
  XOR U15909 ( .A(n15965), .B(n15923), .Z(n15926) );
  XOR U15910 ( .A(p_input[1034]), .B(p_input[762]), .Z(n15923) );
  XNOR U15911 ( .A(p_input[1035]), .B(p_input[763]), .Z(n15965) );
  XOR U15912 ( .A(p_input[1036]), .B(p_input[764]), .Z(n15927) );
  XNOR U15913 ( .A(n15937), .B(n15928), .Z(n15964) );
  XOR U15914 ( .A(p_input[1025]), .B(p_input[753]), .Z(n15928) );
  XOR U15915 ( .A(n15966), .B(n15943), .Z(n15937) );
  XNOR U15916 ( .A(p_input[1039]), .B(p_input[767]), .Z(n15943) );
  XOR U15917 ( .A(n15934), .B(n15942), .Z(n15966) );
  XOR U15918 ( .A(n15967), .B(n15939), .Z(n15942) );
  XOR U15919 ( .A(p_input[1037]), .B(p_input[765]), .Z(n15939) );
  XNOR U15920 ( .A(p_input[1038]), .B(p_input[766]), .Z(n15967) );
  XOR U15921 ( .A(p_input[1033]), .B(p_input[761]), .Z(n15934) );
  XNOR U15922 ( .A(n15950), .B(n15949), .Z(n15932) );
  XNOR U15923 ( .A(n15968), .B(n15955), .Z(n15949) );
  XOR U15924 ( .A(p_input[1032]), .B(p_input[760]), .Z(n15955) );
  XOR U15925 ( .A(n15946), .B(n15954), .Z(n15968) );
  XOR U15926 ( .A(n15969), .B(n15951), .Z(n15954) );
  XOR U15927 ( .A(p_input[1030]), .B(p_input[758]), .Z(n15951) );
  XNOR U15928 ( .A(p_input[1031]), .B(p_input[759]), .Z(n15969) );
  XOR U15929 ( .A(p_input[1026]), .B(p_input[754]), .Z(n15946) );
  XNOR U15930 ( .A(n15960), .B(n15959), .Z(n15950) );
  XOR U15931 ( .A(n15970), .B(n15956), .Z(n15959) );
  XOR U15932 ( .A(p_input[1027]), .B(p_input[755]), .Z(n15956) );
  XNOR U15933 ( .A(p_input[1028]), .B(p_input[756]), .Z(n15970) );
  XOR U15934 ( .A(p_input[1029]), .B(p_input[757]), .Z(n15960) );
  XNOR U15935 ( .A(n15971), .B(n15972), .Z(n15867) );
  AND U15936 ( .A(n556), .B(n15973), .Z(n15972) );
  XNOR U15937 ( .A(n15974), .B(n15975), .Z(n556) );
  AND U15938 ( .A(n15976), .B(n15977), .Z(n15975) );
  XOR U15939 ( .A(n15974), .B(n15877), .Z(n15977) );
  XNOR U15940 ( .A(n15974), .B(n15831), .Z(n15976) );
  XOR U15941 ( .A(n15978), .B(n15979), .Z(n15974) );
  AND U15942 ( .A(n15980), .B(n15981), .Z(n15979) );
  XOR U15943 ( .A(n15978), .B(n15841), .Z(n15980) );
  XOR U15944 ( .A(n15982), .B(n15983), .Z(n15820) );
  AND U15945 ( .A(n560), .B(n15973), .Z(n15983) );
  XNOR U15946 ( .A(n15971), .B(n15982), .Z(n15973) );
  XNOR U15947 ( .A(n15984), .B(n15985), .Z(n560) );
  AND U15948 ( .A(n15986), .B(n15987), .Z(n15985) );
  XNOR U15949 ( .A(n15988), .B(n15984), .Z(n15987) );
  IV U15950 ( .A(n15877), .Z(n15988) );
  XNOR U15951 ( .A(n15989), .B(n15990), .Z(n15877) );
  AND U15952 ( .A(n563), .B(n15991), .Z(n15990) );
  XNOR U15953 ( .A(n15989), .B(n15992), .Z(n15991) );
  XNOR U15954 ( .A(n15831), .B(n15984), .Z(n15986) );
  XOR U15955 ( .A(n15993), .B(n15994), .Z(n15831) );
  AND U15956 ( .A(n571), .B(n15995), .Z(n15994) );
  XOR U15957 ( .A(n15978), .B(n15996), .Z(n15984) );
  AND U15958 ( .A(n15997), .B(n15981), .Z(n15996) );
  XNOR U15959 ( .A(n15890), .B(n15978), .Z(n15981) );
  XNOR U15960 ( .A(n15998), .B(n15999), .Z(n15890) );
  AND U15961 ( .A(n563), .B(n16000), .Z(n15999) );
  XOR U15962 ( .A(n16001), .B(n15998), .Z(n16000) );
  XNOR U15963 ( .A(n16002), .B(n15978), .Z(n15997) );
  IV U15964 ( .A(n15841), .Z(n16002) );
  XOR U15965 ( .A(n16003), .B(n16004), .Z(n15841) );
  AND U15966 ( .A(n571), .B(n16005), .Z(n16004) );
  XOR U15967 ( .A(n16006), .B(n16007), .Z(n15978) );
  AND U15968 ( .A(n16008), .B(n16009), .Z(n16007) );
  XNOR U15969 ( .A(n15915), .B(n16006), .Z(n16009) );
  XNOR U15970 ( .A(n16010), .B(n16011), .Z(n15915) );
  AND U15971 ( .A(n563), .B(n16012), .Z(n16011) );
  XNOR U15972 ( .A(n16013), .B(n16010), .Z(n16012) );
  XOR U15973 ( .A(n16006), .B(n15852), .Z(n16008) );
  XOR U15974 ( .A(n16014), .B(n16015), .Z(n15852) );
  AND U15975 ( .A(n571), .B(n16016), .Z(n16015) );
  XOR U15976 ( .A(n16017), .B(n16018), .Z(n16006) );
  AND U15977 ( .A(n16019), .B(n16020), .Z(n16018) );
  XNOR U15978 ( .A(n16017), .B(n15961), .Z(n16020) );
  XNOR U15979 ( .A(n16021), .B(n16022), .Z(n15961) );
  AND U15980 ( .A(n563), .B(n16023), .Z(n16022) );
  XOR U15981 ( .A(n16024), .B(n16021), .Z(n16023) );
  XNOR U15982 ( .A(n16025), .B(n16017), .Z(n16019) );
  IV U15983 ( .A(n15864), .Z(n16025) );
  XOR U15984 ( .A(n16026), .B(n16027), .Z(n15864) );
  AND U15985 ( .A(n571), .B(n16028), .Z(n16027) );
  AND U15986 ( .A(n15982), .B(n15971), .Z(n16017) );
  XNOR U15987 ( .A(n16029), .B(n16030), .Z(n15971) );
  AND U15988 ( .A(n563), .B(n16031), .Z(n16030) );
  XNOR U15989 ( .A(n16032), .B(n16029), .Z(n16031) );
  XNOR U15990 ( .A(n16033), .B(n16034), .Z(n563) );
  AND U15991 ( .A(n16035), .B(n16036), .Z(n16034) );
  XOR U15992 ( .A(n15992), .B(n16033), .Z(n16036) );
  AND U15993 ( .A(n16037), .B(n16038), .Z(n15992) );
  XOR U15994 ( .A(n16033), .B(n15989), .Z(n16035) );
  XNOR U15995 ( .A(n16039), .B(n16040), .Z(n15989) );
  AND U15996 ( .A(n567), .B(n15995), .Z(n16040) );
  XOR U15997 ( .A(n15993), .B(n16039), .Z(n15995) );
  XOR U15998 ( .A(n16041), .B(n16042), .Z(n16033) );
  AND U15999 ( .A(n16043), .B(n16044), .Z(n16042) );
  XNOR U16000 ( .A(n16041), .B(n16037), .Z(n16044) );
  IV U16001 ( .A(n16001), .Z(n16037) );
  XOR U16002 ( .A(n16045), .B(n16046), .Z(n16001) );
  XOR U16003 ( .A(n16047), .B(n16038), .Z(n16046) );
  AND U16004 ( .A(n16013), .B(n16048), .Z(n16038) );
  AND U16005 ( .A(n16049), .B(n16050), .Z(n16047) );
  XOR U16006 ( .A(n16051), .B(n16045), .Z(n16049) );
  XNOR U16007 ( .A(n15998), .B(n16041), .Z(n16043) );
  XNOR U16008 ( .A(n16052), .B(n16053), .Z(n15998) );
  AND U16009 ( .A(n567), .B(n16005), .Z(n16053) );
  XOR U16010 ( .A(n16052), .B(n16003), .Z(n16005) );
  XOR U16011 ( .A(n16054), .B(n16055), .Z(n16041) );
  AND U16012 ( .A(n16056), .B(n16057), .Z(n16055) );
  XNOR U16013 ( .A(n16054), .B(n16013), .Z(n16057) );
  XOR U16014 ( .A(n16058), .B(n16050), .Z(n16013) );
  XNOR U16015 ( .A(n16059), .B(n16045), .Z(n16050) );
  XOR U16016 ( .A(n16060), .B(n16061), .Z(n16045) );
  AND U16017 ( .A(n16062), .B(n16063), .Z(n16061) );
  XOR U16018 ( .A(n16064), .B(n16060), .Z(n16062) );
  XNOR U16019 ( .A(n16065), .B(n16066), .Z(n16059) );
  AND U16020 ( .A(n16067), .B(n16068), .Z(n16066) );
  XOR U16021 ( .A(n16065), .B(n16069), .Z(n16067) );
  XNOR U16022 ( .A(n16051), .B(n16048), .Z(n16058) );
  AND U16023 ( .A(n16070), .B(n16071), .Z(n16048) );
  XOR U16024 ( .A(n16072), .B(n16073), .Z(n16051) );
  AND U16025 ( .A(n16074), .B(n16075), .Z(n16073) );
  XOR U16026 ( .A(n16072), .B(n16076), .Z(n16074) );
  XNOR U16027 ( .A(n16010), .B(n16054), .Z(n16056) );
  XNOR U16028 ( .A(n16077), .B(n16078), .Z(n16010) );
  AND U16029 ( .A(n567), .B(n16016), .Z(n16078) );
  XOR U16030 ( .A(n16077), .B(n16014), .Z(n16016) );
  XOR U16031 ( .A(n16079), .B(n16080), .Z(n16054) );
  AND U16032 ( .A(n16081), .B(n16082), .Z(n16080) );
  XNOR U16033 ( .A(n16079), .B(n16070), .Z(n16082) );
  IV U16034 ( .A(n16024), .Z(n16070) );
  XNOR U16035 ( .A(n16083), .B(n16063), .Z(n16024) );
  XNOR U16036 ( .A(n16084), .B(n16069), .Z(n16063) );
  XOR U16037 ( .A(n16085), .B(n16086), .Z(n16069) );
  NOR U16038 ( .A(n16087), .B(n16088), .Z(n16086) );
  XNOR U16039 ( .A(n16085), .B(n16089), .Z(n16087) );
  XNOR U16040 ( .A(n16068), .B(n16060), .Z(n16084) );
  XOR U16041 ( .A(n16090), .B(n16091), .Z(n16060) );
  AND U16042 ( .A(n16092), .B(n16093), .Z(n16091) );
  XNOR U16043 ( .A(n16090), .B(n16094), .Z(n16092) );
  XNOR U16044 ( .A(n16095), .B(n16065), .Z(n16068) );
  XOR U16045 ( .A(n16096), .B(n16097), .Z(n16065) );
  AND U16046 ( .A(n16098), .B(n16099), .Z(n16097) );
  XOR U16047 ( .A(n16096), .B(n16100), .Z(n16098) );
  XNOR U16048 ( .A(n16101), .B(n16102), .Z(n16095) );
  NOR U16049 ( .A(n16103), .B(n16104), .Z(n16102) );
  XOR U16050 ( .A(n16101), .B(n16105), .Z(n16103) );
  XNOR U16051 ( .A(n16064), .B(n16071), .Z(n16083) );
  NOR U16052 ( .A(n16032), .B(n16106), .Z(n16071) );
  XOR U16053 ( .A(n16076), .B(n16075), .Z(n16064) );
  XNOR U16054 ( .A(n16107), .B(n16072), .Z(n16075) );
  XOR U16055 ( .A(n16108), .B(n16109), .Z(n16072) );
  AND U16056 ( .A(n16110), .B(n16111), .Z(n16109) );
  XOR U16057 ( .A(n16108), .B(n16112), .Z(n16110) );
  XNOR U16058 ( .A(n16113), .B(n16114), .Z(n16107) );
  NOR U16059 ( .A(n16115), .B(n16116), .Z(n16114) );
  XNOR U16060 ( .A(n16113), .B(n16117), .Z(n16115) );
  XOR U16061 ( .A(n16118), .B(n16119), .Z(n16076) );
  NOR U16062 ( .A(n16120), .B(n16121), .Z(n16119) );
  XNOR U16063 ( .A(n16118), .B(n16122), .Z(n16120) );
  XNOR U16064 ( .A(n16021), .B(n16079), .Z(n16081) );
  XNOR U16065 ( .A(n16123), .B(n16124), .Z(n16021) );
  AND U16066 ( .A(n567), .B(n16028), .Z(n16124) );
  XOR U16067 ( .A(n16123), .B(n16026), .Z(n16028) );
  AND U16068 ( .A(n16029), .B(n16032), .Z(n16079) );
  XOR U16069 ( .A(n16125), .B(n16106), .Z(n16032) );
  XNOR U16070 ( .A(p_input[1024]), .B(p_input[768]), .Z(n16106) );
  XOR U16071 ( .A(n16094), .B(n16093), .Z(n16125) );
  XNOR U16072 ( .A(n16126), .B(n16100), .Z(n16093) );
  XNOR U16073 ( .A(n16089), .B(n16088), .Z(n16100) );
  XOR U16074 ( .A(n16127), .B(n16085), .Z(n16088) );
  XOR U16075 ( .A(p_input[1034]), .B(p_input[778]), .Z(n16085) );
  XNOR U16076 ( .A(p_input[1035]), .B(p_input[779]), .Z(n16127) );
  XOR U16077 ( .A(p_input[1036]), .B(p_input[780]), .Z(n16089) );
  XNOR U16078 ( .A(n16099), .B(n16090), .Z(n16126) );
  XOR U16079 ( .A(p_input[1025]), .B(p_input[769]), .Z(n16090) );
  XOR U16080 ( .A(n16128), .B(n16105), .Z(n16099) );
  XNOR U16081 ( .A(p_input[1039]), .B(p_input[783]), .Z(n16105) );
  XOR U16082 ( .A(n16096), .B(n16104), .Z(n16128) );
  XOR U16083 ( .A(n16129), .B(n16101), .Z(n16104) );
  XOR U16084 ( .A(p_input[1037]), .B(p_input[781]), .Z(n16101) );
  XNOR U16085 ( .A(p_input[1038]), .B(p_input[782]), .Z(n16129) );
  XOR U16086 ( .A(p_input[1033]), .B(p_input[777]), .Z(n16096) );
  XNOR U16087 ( .A(n16112), .B(n16111), .Z(n16094) );
  XNOR U16088 ( .A(n16130), .B(n16117), .Z(n16111) );
  XOR U16089 ( .A(p_input[1032]), .B(p_input[776]), .Z(n16117) );
  XOR U16090 ( .A(n16108), .B(n16116), .Z(n16130) );
  XOR U16091 ( .A(n16131), .B(n16113), .Z(n16116) );
  XOR U16092 ( .A(p_input[1030]), .B(p_input[774]), .Z(n16113) );
  XNOR U16093 ( .A(p_input[1031]), .B(p_input[775]), .Z(n16131) );
  XOR U16094 ( .A(p_input[1026]), .B(p_input[770]), .Z(n16108) );
  XNOR U16095 ( .A(n16122), .B(n16121), .Z(n16112) );
  XOR U16096 ( .A(n16132), .B(n16118), .Z(n16121) );
  XOR U16097 ( .A(p_input[1027]), .B(p_input[771]), .Z(n16118) );
  XNOR U16098 ( .A(p_input[1028]), .B(p_input[772]), .Z(n16132) );
  XOR U16099 ( .A(p_input[1029]), .B(p_input[773]), .Z(n16122) );
  XNOR U16100 ( .A(n16133), .B(n16134), .Z(n16029) );
  AND U16101 ( .A(n567), .B(n16135), .Z(n16134) );
  XNOR U16102 ( .A(n16136), .B(n16137), .Z(n567) );
  AND U16103 ( .A(n16138), .B(n16139), .Z(n16137) );
  XOR U16104 ( .A(n16136), .B(n16039), .Z(n16139) );
  XNOR U16105 ( .A(n16136), .B(n15993), .Z(n16138) );
  XOR U16106 ( .A(n16140), .B(n16141), .Z(n16136) );
  AND U16107 ( .A(n16142), .B(n16143), .Z(n16141) );
  XOR U16108 ( .A(n16140), .B(n16003), .Z(n16142) );
  XOR U16109 ( .A(n16144), .B(n16145), .Z(n15982) );
  AND U16110 ( .A(n571), .B(n16135), .Z(n16145) );
  XNOR U16111 ( .A(n16133), .B(n16144), .Z(n16135) );
  XNOR U16112 ( .A(n16146), .B(n16147), .Z(n571) );
  AND U16113 ( .A(n16148), .B(n16149), .Z(n16147) );
  XNOR U16114 ( .A(n16150), .B(n16146), .Z(n16149) );
  IV U16115 ( .A(n16039), .Z(n16150) );
  XNOR U16116 ( .A(n16151), .B(n16152), .Z(n16039) );
  AND U16117 ( .A(n574), .B(n16153), .Z(n16152) );
  XNOR U16118 ( .A(n16151), .B(n16154), .Z(n16153) );
  XNOR U16119 ( .A(n15993), .B(n16146), .Z(n16148) );
  XOR U16120 ( .A(n16155), .B(n16156), .Z(n15993) );
  AND U16121 ( .A(n582), .B(n16157), .Z(n16156) );
  XOR U16122 ( .A(n16140), .B(n16158), .Z(n16146) );
  AND U16123 ( .A(n16159), .B(n16143), .Z(n16158) );
  XNOR U16124 ( .A(n16052), .B(n16140), .Z(n16143) );
  XNOR U16125 ( .A(n16160), .B(n16161), .Z(n16052) );
  AND U16126 ( .A(n574), .B(n16162), .Z(n16161) );
  XOR U16127 ( .A(n16163), .B(n16160), .Z(n16162) );
  XNOR U16128 ( .A(n16164), .B(n16140), .Z(n16159) );
  IV U16129 ( .A(n16003), .Z(n16164) );
  XOR U16130 ( .A(n16165), .B(n16166), .Z(n16003) );
  AND U16131 ( .A(n582), .B(n16167), .Z(n16166) );
  XOR U16132 ( .A(n16168), .B(n16169), .Z(n16140) );
  AND U16133 ( .A(n16170), .B(n16171), .Z(n16169) );
  XNOR U16134 ( .A(n16077), .B(n16168), .Z(n16171) );
  XNOR U16135 ( .A(n16172), .B(n16173), .Z(n16077) );
  AND U16136 ( .A(n574), .B(n16174), .Z(n16173) );
  XNOR U16137 ( .A(n16175), .B(n16172), .Z(n16174) );
  XOR U16138 ( .A(n16168), .B(n16014), .Z(n16170) );
  XOR U16139 ( .A(n16176), .B(n16177), .Z(n16014) );
  AND U16140 ( .A(n582), .B(n16178), .Z(n16177) );
  XOR U16141 ( .A(n16179), .B(n16180), .Z(n16168) );
  AND U16142 ( .A(n16181), .B(n16182), .Z(n16180) );
  XNOR U16143 ( .A(n16179), .B(n16123), .Z(n16182) );
  XNOR U16144 ( .A(n16183), .B(n16184), .Z(n16123) );
  AND U16145 ( .A(n574), .B(n16185), .Z(n16184) );
  XOR U16146 ( .A(n16186), .B(n16183), .Z(n16185) );
  XNOR U16147 ( .A(n16187), .B(n16179), .Z(n16181) );
  IV U16148 ( .A(n16026), .Z(n16187) );
  XOR U16149 ( .A(n16188), .B(n16189), .Z(n16026) );
  AND U16150 ( .A(n582), .B(n16190), .Z(n16189) );
  AND U16151 ( .A(n16144), .B(n16133), .Z(n16179) );
  XNOR U16152 ( .A(n16191), .B(n16192), .Z(n16133) );
  AND U16153 ( .A(n574), .B(n16193), .Z(n16192) );
  XNOR U16154 ( .A(n16194), .B(n16191), .Z(n16193) );
  XNOR U16155 ( .A(n16195), .B(n16196), .Z(n574) );
  AND U16156 ( .A(n16197), .B(n16198), .Z(n16196) );
  XOR U16157 ( .A(n16154), .B(n16195), .Z(n16198) );
  AND U16158 ( .A(n16199), .B(n16200), .Z(n16154) );
  XOR U16159 ( .A(n16195), .B(n16151), .Z(n16197) );
  XNOR U16160 ( .A(n16201), .B(n16202), .Z(n16151) );
  AND U16161 ( .A(n578), .B(n16157), .Z(n16202) );
  XOR U16162 ( .A(n16155), .B(n16201), .Z(n16157) );
  XOR U16163 ( .A(n16203), .B(n16204), .Z(n16195) );
  AND U16164 ( .A(n16205), .B(n16206), .Z(n16204) );
  XNOR U16165 ( .A(n16203), .B(n16199), .Z(n16206) );
  IV U16166 ( .A(n16163), .Z(n16199) );
  XOR U16167 ( .A(n16207), .B(n16208), .Z(n16163) );
  XOR U16168 ( .A(n16209), .B(n16200), .Z(n16208) );
  AND U16169 ( .A(n16175), .B(n16210), .Z(n16200) );
  AND U16170 ( .A(n16211), .B(n16212), .Z(n16209) );
  XOR U16171 ( .A(n16213), .B(n16207), .Z(n16211) );
  XNOR U16172 ( .A(n16160), .B(n16203), .Z(n16205) );
  XNOR U16173 ( .A(n16214), .B(n16215), .Z(n16160) );
  AND U16174 ( .A(n578), .B(n16167), .Z(n16215) );
  XOR U16175 ( .A(n16214), .B(n16165), .Z(n16167) );
  XOR U16176 ( .A(n16216), .B(n16217), .Z(n16203) );
  AND U16177 ( .A(n16218), .B(n16219), .Z(n16217) );
  XNOR U16178 ( .A(n16216), .B(n16175), .Z(n16219) );
  XOR U16179 ( .A(n16220), .B(n16212), .Z(n16175) );
  XNOR U16180 ( .A(n16221), .B(n16207), .Z(n16212) );
  XOR U16181 ( .A(n16222), .B(n16223), .Z(n16207) );
  AND U16182 ( .A(n16224), .B(n16225), .Z(n16223) );
  XOR U16183 ( .A(n16226), .B(n16222), .Z(n16224) );
  XNOR U16184 ( .A(n16227), .B(n16228), .Z(n16221) );
  AND U16185 ( .A(n16229), .B(n16230), .Z(n16228) );
  XOR U16186 ( .A(n16227), .B(n16231), .Z(n16229) );
  XNOR U16187 ( .A(n16213), .B(n16210), .Z(n16220) );
  AND U16188 ( .A(n16232), .B(n16233), .Z(n16210) );
  XOR U16189 ( .A(n16234), .B(n16235), .Z(n16213) );
  AND U16190 ( .A(n16236), .B(n16237), .Z(n16235) );
  XOR U16191 ( .A(n16234), .B(n16238), .Z(n16236) );
  XNOR U16192 ( .A(n16172), .B(n16216), .Z(n16218) );
  XNOR U16193 ( .A(n16239), .B(n16240), .Z(n16172) );
  AND U16194 ( .A(n578), .B(n16178), .Z(n16240) );
  XOR U16195 ( .A(n16239), .B(n16176), .Z(n16178) );
  XOR U16196 ( .A(n16241), .B(n16242), .Z(n16216) );
  AND U16197 ( .A(n16243), .B(n16244), .Z(n16242) );
  XNOR U16198 ( .A(n16241), .B(n16232), .Z(n16244) );
  IV U16199 ( .A(n16186), .Z(n16232) );
  XNOR U16200 ( .A(n16245), .B(n16225), .Z(n16186) );
  XNOR U16201 ( .A(n16246), .B(n16231), .Z(n16225) );
  XOR U16202 ( .A(n16247), .B(n16248), .Z(n16231) );
  NOR U16203 ( .A(n16249), .B(n16250), .Z(n16248) );
  XNOR U16204 ( .A(n16247), .B(n16251), .Z(n16249) );
  XNOR U16205 ( .A(n16230), .B(n16222), .Z(n16246) );
  XOR U16206 ( .A(n16252), .B(n16253), .Z(n16222) );
  AND U16207 ( .A(n16254), .B(n16255), .Z(n16253) );
  XNOR U16208 ( .A(n16252), .B(n16256), .Z(n16254) );
  XNOR U16209 ( .A(n16257), .B(n16227), .Z(n16230) );
  XOR U16210 ( .A(n16258), .B(n16259), .Z(n16227) );
  AND U16211 ( .A(n16260), .B(n16261), .Z(n16259) );
  XOR U16212 ( .A(n16258), .B(n16262), .Z(n16260) );
  XNOR U16213 ( .A(n16263), .B(n16264), .Z(n16257) );
  NOR U16214 ( .A(n16265), .B(n16266), .Z(n16264) );
  XOR U16215 ( .A(n16263), .B(n16267), .Z(n16265) );
  XNOR U16216 ( .A(n16226), .B(n16233), .Z(n16245) );
  NOR U16217 ( .A(n16194), .B(n16268), .Z(n16233) );
  XOR U16218 ( .A(n16238), .B(n16237), .Z(n16226) );
  XNOR U16219 ( .A(n16269), .B(n16234), .Z(n16237) );
  XOR U16220 ( .A(n16270), .B(n16271), .Z(n16234) );
  AND U16221 ( .A(n16272), .B(n16273), .Z(n16271) );
  XOR U16222 ( .A(n16270), .B(n16274), .Z(n16272) );
  XNOR U16223 ( .A(n16275), .B(n16276), .Z(n16269) );
  NOR U16224 ( .A(n16277), .B(n16278), .Z(n16276) );
  XNOR U16225 ( .A(n16275), .B(n16279), .Z(n16277) );
  XOR U16226 ( .A(n16280), .B(n16281), .Z(n16238) );
  NOR U16227 ( .A(n16282), .B(n16283), .Z(n16281) );
  XNOR U16228 ( .A(n16280), .B(n16284), .Z(n16282) );
  XNOR U16229 ( .A(n16183), .B(n16241), .Z(n16243) );
  XNOR U16230 ( .A(n16285), .B(n16286), .Z(n16183) );
  AND U16231 ( .A(n578), .B(n16190), .Z(n16286) );
  XOR U16232 ( .A(n16285), .B(n16188), .Z(n16190) );
  AND U16233 ( .A(n16191), .B(n16194), .Z(n16241) );
  XOR U16234 ( .A(n16287), .B(n16268), .Z(n16194) );
  XNOR U16235 ( .A(p_input[1024]), .B(p_input[784]), .Z(n16268) );
  XOR U16236 ( .A(n16256), .B(n16255), .Z(n16287) );
  XNOR U16237 ( .A(n16288), .B(n16262), .Z(n16255) );
  XNOR U16238 ( .A(n16251), .B(n16250), .Z(n16262) );
  XOR U16239 ( .A(n16289), .B(n16247), .Z(n16250) );
  XOR U16240 ( .A(p_input[1034]), .B(p_input[794]), .Z(n16247) );
  XNOR U16241 ( .A(p_input[1035]), .B(p_input[795]), .Z(n16289) );
  XOR U16242 ( .A(p_input[1036]), .B(p_input[796]), .Z(n16251) );
  XNOR U16243 ( .A(n16261), .B(n16252), .Z(n16288) );
  XOR U16244 ( .A(p_input[1025]), .B(p_input[785]), .Z(n16252) );
  XOR U16245 ( .A(n16290), .B(n16267), .Z(n16261) );
  XNOR U16246 ( .A(p_input[1039]), .B(p_input[799]), .Z(n16267) );
  XOR U16247 ( .A(n16258), .B(n16266), .Z(n16290) );
  XOR U16248 ( .A(n16291), .B(n16263), .Z(n16266) );
  XOR U16249 ( .A(p_input[1037]), .B(p_input[797]), .Z(n16263) );
  XNOR U16250 ( .A(p_input[1038]), .B(p_input[798]), .Z(n16291) );
  XOR U16251 ( .A(p_input[1033]), .B(p_input[793]), .Z(n16258) );
  XNOR U16252 ( .A(n16274), .B(n16273), .Z(n16256) );
  XNOR U16253 ( .A(n16292), .B(n16279), .Z(n16273) );
  XOR U16254 ( .A(p_input[1032]), .B(p_input[792]), .Z(n16279) );
  XOR U16255 ( .A(n16270), .B(n16278), .Z(n16292) );
  XOR U16256 ( .A(n16293), .B(n16275), .Z(n16278) );
  XOR U16257 ( .A(p_input[1030]), .B(p_input[790]), .Z(n16275) );
  XNOR U16258 ( .A(p_input[1031]), .B(p_input[791]), .Z(n16293) );
  XOR U16259 ( .A(p_input[1026]), .B(p_input[786]), .Z(n16270) );
  XNOR U16260 ( .A(n16284), .B(n16283), .Z(n16274) );
  XOR U16261 ( .A(n16294), .B(n16280), .Z(n16283) );
  XOR U16262 ( .A(p_input[1027]), .B(p_input[787]), .Z(n16280) );
  XNOR U16263 ( .A(p_input[1028]), .B(p_input[788]), .Z(n16294) );
  XOR U16264 ( .A(p_input[1029]), .B(p_input[789]), .Z(n16284) );
  XNOR U16265 ( .A(n16295), .B(n16296), .Z(n16191) );
  AND U16266 ( .A(n578), .B(n16297), .Z(n16296) );
  XNOR U16267 ( .A(n16298), .B(n16299), .Z(n578) );
  AND U16268 ( .A(n16300), .B(n16301), .Z(n16299) );
  XOR U16269 ( .A(n16298), .B(n16201), .Z(n16301) );
  XNOR U16270 ( .A(n16298), .B(n16155), .Z(n16300) );
  XOR U16271 ( .A(n16302), .B(n16303), .Z(n16298) );
  AND U16272 ( .A(n16304), .B(n16305), .Z(n16303) );
  XOR U16273 ( .A(n16302), .B(n16165), .Z(n16304) );
  XOR U16274 ( .A(n16306), .B(n16307), .Z(n16144) );
  AND U16275 ( .A(n582), .B(n16297), .Z(n16307) );
  XNOR U16276 ( .A(n16295), .B(n16306), .Z(n16297) );
  XNOR U16277 ( .A(n16308), .B(n16309), .Z(n582) );
  AND U16278 ( .A(n16310), .B(n16311), .Z(n16309) );
  XNOR U16279 ( .A(n16312), .B(n16308), .Z(n16311) );
  IV U16280 ( .A(n16201), .Z(n16312) );
  XNOR U16281 ( .A(n16313), .B(n16314), .Z(n16201) );
  AND U16282 ( .A(n585), .B(n16315), .Z(n16314) );
  XNOR U16283 ( .A(n16313), .B(n16316), .Z(n16315) );
  XNOR U16284 ( .A(n16155), .B(n16308), .Z(n16310) );
  XOR U16285 ( .A(n16317), .B(n16318), .Z(n16155) );
  AND U16286 ( .A(n593), .B(n16319), .Z(n16318) );
  XOR U16287 ( .A(n16302), .B(n16320), .Z(n16308) );
  AND U16288 ( .A(n16321), .B(n16305), .Z(n16320) );
  XNOR U16289 ( .A(n16214), .B(n16302), .Z(n16305) );
  XNOR U16290 ( .A(n16322), .B(n16323), .Z(n16214) );
  AND U16291 ( .A(n585), .B(n16324), .Z(n16323) );
  XOR U16292 ( .A(n16325), .B(n16322), .Z(n16324) );
  XNOR U16293 ( .A(n16326), .B(n16302), .Z(n16321) );
  IV U16294 ( .A(n16165), .Z(n16326) );
  XOR U16295 ( .A(n16327), .B(n16328), .Z(n16165) );
  AND U16296 ( .A(n593), .B(n16329), .Z(n16328) );
  XOR U16297 ( .A(n16330), .B(n16331), .Z(n16302) );
  AND U16298 ( .A(n16332), .B(n16333), .Z(n16331) );
  XNOR U16299 ( .A(n16239), .B(n16330), .Z(n16333) );
  XNOR U16300 ( .A(n16334), .B(n16335), .Z(n16239) );
  AND U16301 ( .A(n585), .B(n16336), .Z(n16335) );
  XNOR U16302 ( .A(n16337), .B(n16334), .Z(n16336) );
  XOR U16303 ( .A(n16330), .B(n16176), .Z(n16332) );
  XOR U16304 ( .A(n16338), .B(n16339), .Z(n16176) );
  AND U16305 ( .A(n593), .B(n16340), .Z(n16339) );
  XOR U16306 ( .A(n16341), .B(n16342), .Z(n16330) );
  AND U16307 ( .A(n16343), .B(n16344), .Z(n16342) );
  XNOR U16308 ( .A(n16341), .B(n16285), .Z(n16344) );
  XNOR U16309 ( .A(n16345), .B(n16346), .Z(n16285) );
  AND U16310 ( .A(n585), .B(n16347), .Z(n16346) );
  XOR U16311 ( .A(n16348), .B(n16345), .Z(n16347) );
  XNOR U16312 ( .A(n16349), .B(n16341), .Z(n16343) );
  IV U16313 ( .A(n16188), .Z(n16349) );
  XOR U16314 ( .A(n16350), .B(n16351), .Z(n16188) );
  AND U16315 ( .A(n593), .B(n16352), .Z(n16351) );
  AND U16316 ( .A(n16306), .B(n16295), .Z(n16341) );
  XNOR U16317 ( .A(n16353), .B(n16354), .Z(n16295) );
  AND U16318 ( .A(n585), .B(n16355), .Z(n16354) );
  XNOR U16319 ( .A(n16356), .B(n16353), .Z(n16355) );
  XNOR U16320 ( .A(n16357), .B(n16358), .Z(n585) );
  AND U16321 ( .A(n16359), .B(n16360), .Z(n16358) );
  XOR U16322 ( .A(n16316), .B(n16357), .Z(n16360) );
  AND U16323 ( .A(n16361), .B(n16362), .Z(n16316) );
  XOR U16324 ( .A(n16357), .B(n16313), .Z(n16359) );
  XNOR U16325 ( .A(n16363), .B(n16364), .Z(n16313) );
  AND U16326 ( .A(n589), .B(n16319), .Z(n16364) );
  XOR U16327 ( .A(n16317), .B(n16363), .Z(n16319) );
  XOR U16328 ( .A(n16365), .B(n16366), .Z(n16357) );
  AND U16329 ( .A(n16367), .B(n16368), .Z(n16366) );
  XNOR U16330 ( .A(n16365), .B(n16361), .Z(n16368) );
  IV U16331 ( .A(n16325), .Z(n16361) );
  XOR U16332 ( .A(n16369), .B(n16370), .Z(n16325) );
  XOR U16333 ( .A(n16371), .B(n16362), .Z(n16370) );
  AND U16334 ( .A(n16337), .B(n16372), .Z(n16362) );
  AND U16335 ( .A(n16373), .B(n16374), .Z(n16371) );
  XOR U16336 ( .A(n16375), .B(n16369), .Z(n16373) );
  XNOR U16337 ( .A(n16322), .B(n16365), .Z(n16367) );
  XNOR U16338 ( .A(n16376), .B(n16377), .Z(n16322) );
  AND U16339 ( .A(n589), .B(n16329), .Z(n16377) );
  XOR U16340 ( .A(n16376), .B(n16327), .Z(n16329) );
  XOR U16341 ( .A(n16378), .B(n16379), .Z(n16365) );
  AND U16342 ( .A(n16380), .B(n16381), .Z(n16379) );
  XNOR U16343 ( .A(n16378), .B(n16337), .Z(n16381) );
  XOR U16344 ( .A(n16382), .B(n16374), .Z(n16337) );
  XNOR U16345 ( .A(n16383), .B(n16369), .Z(n16374) );
  XOR U16346 ( .A(n16384), .B(n16385), .Z(n16369) );
  AND U16347 ( .A(n16386), .B(n16387), .Z(n16385) );
  XOR U16348 ( .A(n16388), .B(n16384), .Z(n16386) );
  XNOR U16349 ( .A(n16389), .B(n16390), .Z(n16383) );
  AND U16350 ( .A(n16391), .B(n16392), .Z(n16390) );
  XOR U16351 ( .A(n16389), .B(n16393), .Z(n16391) );
  XNOR U16352 ( .A(n16375), .B(n16372), .Z(n16382) );
  AND U16353 ( .A(n16394), .B(n16395), .Z(n16372) );
  XOR U16354 ( .A(n16396), .B(n16397), .Z(n16375) );
  AND U16355 ( .A(n16398), .B(n16399), .Z(n16397) );
  XOR U16356 ( .A(n16396), .B(n16400), .Z(n16398) );
  XNOR U16357 ( .A(n16334), .B(n16378), .Z(n16380) );
  XNOR U16358 ( .A(n16401), .B(n16402), .Z(n16334) );
  AND U16359 ( .A(n589), .B(n16340), .Z(n16402) );
  XOR U16360 ( .A(n16401), .B(n16338), .Z(n16340) );
  XOR U16361 ( .A(n16403), .B(n16404), .Z(n16378) );
  AND U16362 ( .A(n16405), .B(n16406), .Z(n16404) );
  XNOR U16363 ( .A(n16403), .B(n16394), .Z(n16406) );
  IV U16364 ( .A(n16348), .Z(n16394) );
  XNOR U16365 ( .A(n16407), .B(n16387), .Z(n16348) );
  XNOR U16366 ( .A(n16408), .B(n16393), .Z(n16387) );
  XOR U16367 ( .A(n16409), .B(n16410), .Z(n16393) );
  NOR U16368 ( .A(n16411), .B(n16412), .Z(n16410) );
  XNOR U16369 ( .A(n16409), .B(n16413), .Z(n16411) );
  XNOR U16370 ( .A(n16392), .B(n16384), .Z(n16408) );
  XOR U16371 ( .A(n16414), .B(n16415), .Z(n16384) );
  AND U16372 ( .A(n16416), .B(n16417), .Z(n16415) );
  XNOR U16373 ( .A(n16414), .B(n16418), .Z(n16416) );
  XNOR U16374 ( .A(n16419), .B(n16389), .Z(n16392) );
  XOR U16375 ( .A(n16420), .B(n16421), .Z(n16389) );
  AND U16376 ( .A(n16422), .B(n16423), .Z(n16421) );
  XOR U16377 ( .A(n16420), .B(n16424), .Z(n16422) );
  XNOR U16378 ( .A(n16425), .B(n16426), .Z(n16419) );
  NOR U16379 ( .A(n16427), .B(n16428), .Z(n16426) );
  XOR U16380 ( .A(n16425), .B(n16429), .Z(n16427) );
  XNOR U16381 ( .A(n16388), .B(n16395), .Z(n16407) );
  NOR U16382 ( .A(n16356), .B(n16430), .Z(n16395) );
  XOR U16383 ( .A(n16400), .B(n16399), .Z(n16388) );
  XNOR U16384 ( .A(n16431), .B(n16396), .Z(n16399) );
  XOR U16385 ( .A(n16432), .B(n16433), .Z(n16396) );
  AND U16386 ( .A(n16434), .B(n16435), .Z(n16433) );
  XOR U16387 ( .A(n16432), .B(n16436), .Z(n16434) );
  XNOR U16388 ( .A(n16437), .B(n16438), .Z(n16431) );
  NOR U16389 ( .A(n16439), .B(n16440), .Z(n16438) );
  XNOR U16390 ( .A(n16437), .B(n16441), .Z(n16439) );
  XOR U16391 ( .A(n16442), .B(n16443), .Z(n16400) );
  NOR U16392 ( .A(n16444), .B(n16445), .Z(n16443) );
  XNOR U16393 ( .A(n16442), .B(n16446), .Z(n16444) );
  XNOR U16394 ( .A(n16345), .B(n16403), .Z(n16405) );
  XNOR U16395 ( .A(n16447), .B(n16448), .Z(n16345) );
  AND U16396 ( .A(n589), .B(n16352), .Z(n16448) );
  XOR U16397 ( .A(n16447), .B(n16350), .Z(n16352) );
  AND U16398 ( .A(n16353), .B(n16356), .Z(n16403) );
  XOR U16399 ( .A(n16449), .B(n16430), .Z(n16356) );
  XNOR U16400 ( .A(p_input[1024]), .B(p_input[800]), .Z(n16430) );
  XOR U16401 ( .A(n16418), .B(n16417), .Z(n16449) );
  XNOR U16402 ( .A(n16450), .B(n16424), .Z(n16417) );
  XNOR U16403 ( .A(n16413), .B(n16412), .Z(n16424) );
  XOR U16404 ( .A(n16451), .B(n16409), .Z(n16412) );
  XOR U16405 ( .A(p_input[1034]), .B(p_input[810]), .Z(n16409) );
  XNOR U16406 ( .A(p_input[1035]), .B(p_input[811]), .Z(n16451) );
  XOR U16407 ( .A(p_input[1036]), .B(p_input[812]), .Z(n16413) );
  XNOR U16408 ( .A(n16423), .B(n16414), .Z(n16450) );
  XOR U16409 ( .A(p_input[1025]), .B(p_input[801]), .Z(n16414) );
  XOR U16410 ( .A(n16452), .B(n16429), .Z(n16423) );
  XNOR U16411 ( .A(p_input[1039]), .B(p_input[815]), .Z(n16429) );
  XOR U16412 ( .A(n16420), .B(n16428), .Z(n16452) );
  XOR U16413 ( .A(n16453), .B(n16425), .Z(n16428) );
  XOR U16414 ( .A(p_input[1037]), .B(p_input[813]), .Z(n16425) );
  XNOR U16415 ( .A(p_input[1038]), .B(p_input[814]), .Z(n16453) );
  XOR U16416 ( .A(p_input[1033]), .B(p_input[809]), .Z(n16420) );
  XNOR U16417 ( .A(n16436), .B(n16435), .Z(n16418) );
  XNOR U16418 ( .A(n16454), .B(n16441), .Z(n16435) );
  XOR U16419 ( .A(p_input[1032]), .B(p_input[808]), .Z(n16441) );
  XOR U16420 ( .A(n16432), .B(n16440), .Z(n16454) );
  XOR U16421 ( .A(n16455), .B(n16437), .Z(n16440) );
  XOR U16422 ( .A(p_input[1030]), .B(p_input[806]), .Z(n16437) );
  XNOR U16423 ( .A(p_input[1031]), .B(p_input[807]), .Z(n16455) );
  XOR U16424 ( .A(p_input[1026]), .B(p_input[802]), .Z(n16432) );
  XNOR U16425 ( .A(n16446), .B(n16445), .Z(n16436) );
  XOR U16426 ( .A(n16456), .B(n16442), .Z(n16445) );
  XOR U16427 ( .A(p_input[1027]), .B(p_input[803]), .Z(n16442) );
  XNOR U16428 ( .A(p_input[1028]), .B(p_input[804]), .Z(n16456) );
  XOR U16429 ( .A(p_input[1029]), .B(p_input[805]), .Z(n16446) );
  XNOR U16430 ( .A(n16457), .B(n16458), .Z(n16353) );
  AND U16431 ( .A(n589), .B(n16459), .Z(n16458) );
  XNOR U16432 ( .A(n16460), .B(n16461), .Z(n589) );
  AND U16433 ( .A(n16462), .B(n16463), .Z(n16461) );
  XOR U16434 ( .A(n16460), .B(n16363), .Z(n16463) );
  XNOR U16435 ( .A(n16460), .B(n16317), .Z(n16462) );
  XOR U16436 ( .A(n16464), .B(n16465), .Z(n16460) );
  AND U16437 ( .A(n16466), .B(n16467), .Z(n16465) );
  XOR U16438 ( .A(n16464), .B(n16327), .Z(n16466) );
  XOR U16439 ( .A(n16468), .B(n16469), .Z(n16306) );
  AND U16440 ( .A(n593), .B(n16459), .Z(n16469) );
  XNOR U16441 ( .A(n16457), .B(n16468), .Z(n16459) );
  XNOR U16442 ( .A(n16470), .B(n16471), .Z(n593) );
  AND U16443 ( .A(n16472), .B(n16473), .Z(n16471) );
  XNOR U16444 ( .A(n16474), .B(n16470), .Z(n16473) );
  IV U16445 ( .A(n16363), .Z(n16474) );
  XNOR U16446 ( .A(n16475), .B(n16476), .Z(n16363) );
  AND U16447 ( .A(n596), .B(n16477), .Z(n16476) );
  XNOR U16448 ( .A(n16475), .B(n16478), .Z(n16477) );
  XNOR U16449 ( .A(n16317), .B(n16470), .Z(n16472) );
  XOR U16450 ( .A(n16479), .B(n16480), .Z(n16317) );
  AND U16451 ( .A(n604), .B(n16481), .Z(n16480) );
  XOR U16452 ( .A(n16464), .B(n16482), .Z(n16470) );
  AND U16453 ( .A(n16483), .B(n16467), .Z(n16482) );
  XNOR U16454 ( .A(n16376), .B(n16464), .Z(n16467) );
  XNOR U16455 ( .A(n16484), .B(n16485), .Z(n16376) );
  AND U16456 ( .A(n596), .B(n16486), .Z(n16485) );
  XOR U16457 ( .A(n16487), .B(n16484), .Z(n16486) );
  XNOR U16458 ( .A(n16488), .B(n16464), .Z(n16483) );
  IV U16459 ( .A(n16327), .Z(n16488) );
  XOR U16460 ( .A(n16489), .B(n16490), .Z(n16327) );
  AND U16461 ( .A(n604), .B(n16491), .Z(n16490) );
  XOR U16462 ( .A(n16492), .B(n16493), .Z(n16464) );
  AND U16463 ( .A(n16494), .B(n16495), .Z(n16493) );
  XNOR U16464 ( .A(n16401), .B(n16492), .Z(n16495) );
  XNOR U16465 ( .A(n16496), .B(n16497), .Z(n16401) );
  AND U16466 ( .A(n596), .B(n16498), .Z(n16497) );
  XNOR U16467 ( .A(n16499), .B(n16496), .Z(n16498) );
  XOR U16468 ( .A(n16492), .B(n16338), .Z(n16494) );
  XOR U16469 ( .A(n16500), .B(n16501), .Z(n16338) );
  AND U16470 ( .A(n604), .B(n16502), .Z(n16501) );
  XOR U16471 ( .A(n16503), .B(n16504), .Z(n16492) );
  AND U16472 ( .A(n16505), .B(n16506), .Z(n16504) );
  XNOR U16473 ( .A(n16503), .B(n16447), .Z(n16506) );
  XNOR U16474 ( .A(n16507), .B(n16508), .Z(n16447) );
  AND U16475 ( .A(n596), .B(n16509), .Z(n16508) );
  XOR U16476 ( .A(n16510), .B(n16507), .Z(n16509) );
  XNOR U16477 ( .A(n16511), .B(n16503), .Z(n16505) );
  IV U16478 ( .A(n16350), .Z(n16511) );
  XOR U16479 ( .A(n16512), .B(n16513), .Z(n16350) );
  AND U16480 ( .A(n604), .B(n16514), .Z(n16513) );
  AND U16481 ( .A(n16468), .B(n16457), .Z(n16503) );
  XNOR U16482 ( .A(n16515), .B(n16516), .Z(n16457) );
  AND U16483 ( .A(n596), .B(n16517), .Z(n16516) );
  XNOR U16484 ( .A(n16518), .B(n16515), .Z(n16517) );
  XNOR U16485 ( .A(n16519), .B(n16520), .Z(n596) );
  AND U16486 ( .A(n16521), .B(n16522), .Z(n16520) );
  XOR U16487 ( .A(n16478), .B(n16519), .Z(n16522) );
  AND U16488 ( .A(n16523), .B(n16524), .Z(n16478) );
  XOR U16489 ( .A(n16519), .B(n16475), .Z(n16521) );
  XNOR U16490 ( .A(n16525), .B(n16526), .Z(n16475) );
  AND U16491 ( .A(n600), .B(n16481), .Z(n16526) );
  XOR U16492 ( .A(n16479), .B(n16525), .Z(n16481) );
  XOR U16493 ( .A(n16527), .B(n16528), .Z(n16519) );
  AND U16494 ( .A(n16529), .B(n16530), .Z(n16528) );
  XNOR U16495 ( .A(n16527), .B(n16523), .Z(n16530) );
  IV U16496 ( .A(n16487), .Z(n16523) );
  XOR U16497 ( .A(n16531), .B(n16532), .Z(n16487) );
  XOR U16498 ( .A(n16533), .B(n16524), .Z(n16532) );
  AND U16499 ( .A(n16499), .B(n16534), .Z(n16524) );
  AND U16500 ( .A(n16535), .B(n16536), .Z(n16533) );
  XOR U16501 ( .A(n16537), .B(n16531), .Z(n16535) );
  XNOR U16502 ( .A(n16484), .B(n16527), .Z(n16529) );
  XNOR U16503 ( .A(n16538), .B(n16539), .Z(n16484) );
  AND U16504 ( .A(n600), .B(n16491), .Z(n16539) );
  XOR U16505 ( .A(n16538), .B(n16489), .Z(n16491) );
  XOR U16506 ( .A(n16540), .B(n16541), .Z(n16527) );
  AND U16507 ( .A(n16542), .B(n16543), .Z(n16541) );
  XNOR U16508 ( .A(n16540), .B(n16499), .Z(n16543) );
  XOR U16509 ( .A(n16544), .B(n16536), .Z(n16499) );
  XNOR U16510 ( .A(n16545), .B(n16531), .Z(n16536) );
  XOR U16511 ( .A(n16546), .B(n16547), .Z(n16531) );
  AND U16512 ( .A(n16548), .B(n16549), .Z(n16547) );
  XOR U16513 ( .A(n16550), .B(n16546), .Z(n16548) );
  XNOR U16514 ( .A(n16551), .B(n16552), .Z(n16545) );
  AND U16515 ( .A(n16553), .B(n16554), .Z(n16552) );
  XOR U16516 ( .A(n16551), .B(n16555), .Z(n16553) );
  XNOR U16517 ( .A(n16537), .B(n16534), .Z(n16544) );
  AND U16518 ( .A(n16556), .B(n16557), .Z(n16534) );
  XOR U16519 ( .A(n16558), .B(n16559), .Z(n16537) );
  AND U16520 ( .A(n16560), .B(n16561), .Z(n16559) );
  XOR U16521 ( .A(n16558), .B(n16562), .Z(n16560) );
  XNOR U16522 ( .A(n16496), .B(n16540), .Z(n16542) );
  XNOR U16523 ( .A(n16563), .B(n16564), .Z(n16496) );
  AND U16524 ( .A(n600), .B(n16502), .Z(n16564) );
  XOR U16525 ( .A(n16563), .B(n16500), .Z(n16502) );
  XOR U16526 ( .A(n16565), .B(n16566), .Z(n16540) );
  AND U16527 ( .A(n16567), .B(n16568), .Z(n16566) );
  XNOR U16528 ( .A(n16565), .B(n16556), .Z(n16568) );
  IV U16529 ( .A(n16510), .Z(n16556) );
  XNOR U16530 ( .A(n16569), .B(n16549), .Z(n16510) );
  XNOR U16531 ( .A(n16570), .B(n16555), .Z(n16549) );
  XOR U16532 ( .A(n16571), .B(n16572), .Z(n16555) );
  NOR U16533 ( .A(n16573), .B(n16574), .Z(n16572) );
  XNOR U16534 ( .A(n16571), .B(n16575), .Z(n16573) );
  XNOR U16535 ( .A(n16554), .B(n16546), .Z(n16570) );
  XOR U16536 ( .A(n16576), .B(n16577), .Z(n16546) );
  AND U16537 ( .A(n16578), .B(n16579), .Z(n16577) );
  XNOR U16538 ( .A(n16576), .B(n16580), .Z(n16578) );
  XNOR U16539 ( .A(n16581), .B(n16551), .Z(n16554) );
  XOR U16540 ( .A(n16582), .B(n16583), .Z(n16551) );
  AND U16541 ( .A(n16584), .B(n16585), .Z(n16583) );
  XOR U16542 ( .A(n16582), .B(n16586), .Z(n16584) );
  XNOR U16543 ( .A(n16587), .B(n16588), .Z(n16581) );
  NOR U16544 ( .A(n16589), .B(n16590), .Z(n16588) );
  XOR U16545 ( .A(n16587), .B(n16591), .Z(n16589) );
  XNOR U16546 ( .A(n16550), .B(n16557), .Z(n16569) );
  NOR U16547 ( .A(n16518), .B(n16592), .Z(n16557) );
  XOR U16548 ( .A(n16562), .B(n16561), .Z(n16550) );
  XNOR U16549 ( .A(n16593), .B(n16558), .Z(n16561) );
  XOR U16550 ( .A(n16594), .B(n16595), .Z(n16558) );
  AND U16551 ( .A(n16596), .B(n16597), .Z(n16595) );
  XOR U16552 ( .A(n16594), .B(n16598), .Z(n16596) );
  XNOR U16553 ( .A(n16599), .B(n16600), .Z(n16593) );
  NOR U16554 ( .A(n16601), .B(n16602), .Z(n16600) );
  XNOR U16555 ( .A(n16599), .B(n16603), .Z(n16601) );
  XOR U16556 ( .A(n16604), .B(n16605), .Z(n16562) );
  NOR U16557 ( .A(n16606), .B(n16607), .Z(n16605) );
  XNOR U16558 ( .A(n16604), .B(n16608), .Z(n16606) );
  XNOR U16559 ( .A(n16507), .B(n16565), .Z(n16567) );
  XNOR U16560 ( .A(n16609), .B(n16610), .Z(n16507) );
  AND U16561 ( .A(n600), .B(n16514), .Z(n16610) );
  XOR U16562 ( .A(n16609), .B(n16512), .Z(n16514) );
  AND U16563 ( .A(n16515), .B(n16518), .Z(n16565) );
  XOR U16564 ( .A(n16611), .B(n16592), .Z(n16518) );
  XNOR U16565 ( .A(p_input[1024]), .B(p_input[816]), .Z(n16592) );
  XOR U16566 ( .A(n16580), .B(n16579), .Z(n16611) );
  XNOR U16567 ( .A(n16612), .B(n16586), .Z(n16579) );
  XNOR U16568 ( .A(n16575), .B(n16574), .Z(n16586) );
  XOR U16569 ( .A(n16613), .B(n16571), .Z(n16574) );
  XOR U16570 ( .A(p_input[1034]), .B(p_input[826]), .Z(n16571) );
  XNOR U16571 ( .A(p_input[1035]), .B(p_input[827]), .Z(n16613) );
  XOR U16572 ( .A(p_input[1036]), .B(p_input[828]), .Z(n16575) );
  XNOR U16573 ( .A(n16585), .B(n16576), .Z(n16612) );
  XOR U16574 ( .A(p_input[1025]), .B(p_input[817]), .Z(n16576) );
  XOR U16575 ( .A(n16614), .B(n16591), .Z(n16585) );
  XNOR U16576 ( .A(p_input[1039]), .B(p_input[831]), .Z(n16591) );
  XOR U16577 ( .A(n16582), .B(n16590), .Z(n16614) );
  XOR U16578 ( .A(n16615), .B(n16587), .Z(n16590) );
  XOR U16579 ( .A(p_input[1037]), .B(p_input[829]), .Z(n16587) );
  XNOR U16580 ( .A(p_input[1038]), .B(p_input[830]), .Z(n16615) );
  XOR U16581 ( .A(p_input[1033]), .B(p_input[825]), .Z(n16582) );
  XNOR U16582 ( .A(n16598), .B(n16597), .Z(n16580) );
  XNOR U16583 ( .A(n16616), .B(n16603), .Z(n16597) );
  XOR U16584 ( .A(p_input[1032]), .B(p_input[824]), .Z(n16603) );
  XOR U16585 ( .A(n16594), .B(n16602), .Z(n16616) );
  XOR U16586 ( .A(n16617), .B(n16599), .Z(n16602) );
  XOR U16587 ( .A(p_input[1030]), .B(p_input[822]), .Z(n16599) );
  XNOR U16588 ( .A(p_input[1031]), .B(p_input[823]), .Z(n16617) );
  XOR U16589 ( .A(p_input[1026]), .B(p_input[818]), .Z(n16594) );
  XNOR U16590 ( .A(n16608), .B(n16607), .Z(n16598) );
  XOR U16591 ( .A(n16618), .B(n16604), .Z(n16607) );
  XOR U16592 ( .A(p_input[1027]), .B(p_input[819]), .Z(n16604) );
  XNOR U16593 ( .A(p_input[1028]), .B(p_input[820]), .Z(n16618) );
  XOR U16594 ( .A(p_input[1029]), .B(p_input[821]), .Z(n16608) );
  XNOR U16595 ( .A(n16619), .B(n16620), .Z(n16515) );
  AND U16596 ( .A(n600), .B(n16621), .Z(n16620) );
  XNOR U16597 ( .A(n16622), .B(n16623), .Z(n600) );
  AND U16598 ( .A(n16624), .B(n16625), .Z(n16623) );
  XOR U16599 ( .A(n16622), .B(n16525), .Z(n16625) );
  XNOR U16600 ( .A(n16622), .B(n16479), .Z(n16624) );
  XOR U16601 ( .A(n16626), .B(n16627), .Z(n16622) );
  AND U16602 ( .A(n16628), .B(n16629), .Z(n16627) );
  XOR U16603 ( .A(n16626), .B(n16489), .Z(n16628) );
  XOR U16604 ( .A(n16630), .B(n16631), .Z(n16468) );
  AND U16605 ( .A(n604), .B(n16621), .Z(n16631) );
  XNOR U16606 ( .A(n16619), .B(n16630), .Z(n16621) );
  XNOR U16607 ( .A(n16632), .B(n16633), .Z(n604) );
  AND U16608 ( .A(n16634), .B(n16635), .Z(n16633) );
  XNOR U16609 ( .A(n16636), .B(n16632), .Z(n16635) );
  IV U16610 ( .A(n16525), .Z(n16636) );
  XNOR U16611 ( .A(n16637), .B(n16638), .Z(n16525) );
  AND U16612 ( .A(n607), .B(n16639), .Z(n16638) );
  XNOR U16613 ( .A(n16637), .B(n16640), .Z(n16639) );
  XNOR U16614 ( .A(n16479), .B(n16632), .Z(n16634) );
  XOR U16615 ( .A(n16641), .B(n16642), .Z(n16479) );
  AND U16616 ( .A(n615), .B(n16643), .Z(n16642) );
  XOR U16617 ( .A(n16626), .B(n16644), .Z(n16632) );
  AND U16618 ( .A(n16645), .B(n16629), .Z(n16644) );
  XNOR U16619 ( .A(n16538), .B(n16626), .Z(n16629) );
  XNOR U16620 ( .A(n16646), .B(n16647), .Z(n16538) );
  AND U16621 ( .A(n607), .B(n16648), .Z(n16647) );
  XOR U16622 ( .A(n16649), .B(n16646), .Z(n16648) );
  XNOR U16623 ( .A(n16650), .B(n16626), .Z(n16645) );
  IV U16624 ( .A(n16489), .Z(n16650) );
  XOR U16625 ( .A(n16651), .B(n16652), .Z(n16489) );
  AND U16626 ( .A(n615), .B(n16653), .Z(n16652) );
  XOR U16627 ( .A(n16654), .B(n16655), .Z(n16626) );
  AND U16628 ( .A(n16656), .B(n16657), .Z(n16655) );
  XNOR U16629 ( .A(n16563), .B(n16654), .Z(n16657) );
  XNOR U16630 ( .A(n16658), .B(n16659), .Z(n16563) );
  AND U16631 ( .A(n607), .B(n16660), .Z(n16659) );
  XNOR U16632 ( .A(n16661), .B(n16658), .Z(n16660) );
  XOR U16633 ( .A(n16654), .B(n16500), .Z(n16656) );
  XOR U16634 ( .A(n16662), .B(n16663), .Z(n16500) );
  AND U16635 ( .A(n615), .B(n16664), .Z(n16663) );
  XOR U16636 ( .A(n16665), .B(n16666), .Z(n16654) );
  AND U16637 ( .A(n16667), .B(n16668), .Z(n16666) );
  XNOR U16638 ( .A(n16665), .B(n16609), .Z(n16668) );
  XNOR U16639 ( .A(n16669), .B(n16670), .Z(n16609) );
  AND U16640 ( .A(n607), .B(n16671), .Z(n16670) );
  XOR U16641 ( .A(n16672), .B(n16669), .Z(n16671) );
  XNOR U16642 ( .A(n16673), .B(n16665), .Z(n16667) );
  IV U16643 ( .A(n16512), .Z(n16673) );
  XOR U16644 ( .A(n16674), .B(n16675), .Z(n16512) );
  AND U16645 ( .A(n615), .B(n16676), .Z(n16675) );
  AND U16646 ( .A(n16630), .B(n16619), .Z(n16665) );
  XNOR U16647 ( .A(n16677), .B(n16678), .Z(n16619) );
  AND U16648 ( .A(n607), .B(n16679), .Z(n16678) );
  XNOR U16649 ( .A(n16680), .B(n16677), .Z(n16679) );
  XNOR U16650 ( .A(n16681), .B(n16682), .Z(n607) );
  AND U16651 ( .A(n16683), .B(n16684), .Z(n16682) );
  XOR U16652 ( .A(n16640), .B(n16681), .Z(n16684) );
  AND U16653 ( .A(n16685), .B(n16686), .Z(n16640) );
  XOR U16654 ( .A(n16681), .B(n16637), .Z(n16683) );
  XNOR U16655 ( .A(n16687), .B(n16688), .Z(n16637) );
  AND U16656 ( .A(n611), .B(n16643), .Z(n16688) );
  XOR U16657 ( .A(n16641), .B(n16687), .Z(n16643) );
  XOR U16658 ( .A(n16689), .B(n16690), .Z(n16681) );
  AND U16659 ( .A(n16691), .B(n16692), .Z(n16690) );
  XNOR U16660 ( .A(n16689), .B(n16685), .Z(n16692) );
  IV U16661 ( .A(n16649), .Z(n16685) );
  XOR U16662 ( .A(n16693), .B(n16694), .Z(n16649) );
  XOR U16663 ( .A(n16695), .B(n16686), .Z(n16694) );
  AND U16664 ( .A(n16661), .B(n16696), .Z(n16686) );
  AND U16665 ( .A(n16697), .B(n16698), .Z(n16695) );
  XOR U16666 ( .A(n16699), .B(n16693), .Z(n16697) );
  XNOR U16667 ( .A(n16646), .B(n16689), .Z(n16691) );
  XNOR U16668 ( .A(n16700), .B(n16701), .Z(n16646) );
  AND U16669 ( .A(n611), .B(n16653), .Z(n16701) );
  XOR U16670 ( .A(n16700), .B(n16651), .Z(n16653) );
  XOR U16671 ( .A(n16702), .B(n16703), .Z(n16689) );
  AND U16672 ( .A(n16704), .B(n16705), .Z(n16703) );
  XNOR U16673 ( .A(n16702), .B(n16661), .Z(n16705) );
  XOR U16674 ( .A(n16706), .B(n16698), .Z(n16661) );
  XNOR U16675 ( .A(n16707), .B(n16693), .Z(n16698) );
  XOR U16676 ( .A(n16708), .B(n16709), .Z(n16693) );
  AND U16677 ( .A(n16710), .B(n16711), .Z(n16709) );
  XOR U16678 ( .A(n16712), .B(n16708), .Z(n16710) );
  XNOR U16679 ( .A(n16713), .B(n16714), .Z(n16707) );
  AND U16680 ( .A(n16715), .B(n16716), .Z(n16714) );
  XOR U16681 ( .A(n16713), .B(n16717), .Z(n16715) );
  XNOR U16682 ( .A(n16699), .B(n16696), .Z(n16706) );
  AND U16683 ( .A(n16718), .B(n16719), .Z(n16696) );
  XOR U16684 ( .A(n16720), .B(n16721), .Z(n16699) );
  AND U16685 ( .A(n16722), .B(n16723), .Z(n16721) );
  XOR U16686 ( .A(n16720), .B(n16724), .Z(n16722) );
  XNOR U16687 ( .A(n16658), .B(n16702), .Z(n16704) );
  XNOR U16688 ( .A(n16725), .B(n16726), .Z(n16658) );
  AND U16689 ( .A(n611), .B(n16664), .Z(n16726) );
  XOR U16690 ( .A(n16725), .B(n16662), .Z(n16664) );
  XOR U16691 ( .A(n16727), .B(n16728), .Z(n16702) );
  AND U16692 ( .A(n16729), .B(n16730), .Z(n16728) );
  XNOR U16693 ( .A(n16727), .B(n16718), .Z(n16730) );
  IV U16694 ( .A(n16672), .Z(n16718) );
  XNOR U16695 ( .A(n16731), .B(n16711), .Z(n16672) );
  XNOR U16696 ( .A(n16732), .B(n16717), .Z(n16711) );
  XOR U16697 ( .A(n16733), .B(n16734), .Z(n16717) );
  NOR U16698 ( .A(n16735), .B(n16736), .Z(n16734) );
  XNOR U16699 ( .A(n16733), .B(n16737), .Z(n16735) );
  XNOR U16700 ( .A(n16716), .B(n16708), .Z(n16732) );
  XOR U16701 ( .A(n16738), .B(n16739), .Z(n16708) );
  AND U16702 ( .A(n16740), .B(n16741), .Z(n16739) );
  XNOR U16703 ( .A(n16738), .B(n16742), .Z(n16740) );
  XNOR U16704 ( .A(n16743), .B(n16713), .Z(n16716) );
  XOR U16705 ( .A(n16744), .B(n16745), .Z(n16713) );
  AND U16706 ( .A(n16746), .B(n16747), .Z(n16745) );
  XOR U16707 ( .A(n16744), .B(n16748), .Z(n16746) );
  XNOR U16708 ( .A(n16749), .B(n16750), .Z(n16743) );
  NOR U16709 ( .A(n16751), .B(n16752), .Z(n16750) );
  XOR U16710 ( .A(n16749), .B(n16753), .Z(n16751) );
  XNOR U16711 ( .A(n16712), .B(n16719), .Z(n16731) );
  NOR U16712 ( .A(n16680), .B(n16754), .Z(n16719) );
  XOR U16713 ( .A(n16724), .B(n16723), .Z(n16712) );
  XNOR U16714 ( .A(n16755), .B(n16720), .Z(n16723) );
  XOR U16715 ( .A(n16756), .B(n16757), .Z(n16720) );
  AND U16716 ( .A(n16758), .B(n16759), .Z(n16757) );
  XOR U16717 ( .A(n16756), .B(n16760), .Z(n16758) );
  XNOR U16718 ( .A(n16761), .B(n16762), .Z(n16755) );
  NOR U16719 ( .A(n16763), .B(n16764), .Z(n16762) );
  XNOR U16720 ( .A(n16761), .B(n16765), .Z(n16763) );
  XOR U16721 ( .A(n16766), .B(n16767), .Z(n16724) );
  NOR U16722 ( .A(n16768), .B(n16769), .Z(n16767) );
  XNOR U16723 ( .A(n16766), .B(n16770), .Z(n16768) );
  XNOR U16724 ( .A(n16669), .B(n16727), .Z(n16729) );
  XNOR U16725 ( .A(n16771), .B(n16772), .Z(n16669) );
  AND U16726 ( .A(n611), .B(n16676), .Z(n16772) );
  XOR U16727 ( .A(n16771), .B(n16674), .Z(n16676) );
  AND U16728 ( .A(n16677), .B(n16680), .Z(n16727) );
  XOR U16729 ( .A(n16773), .B(n16754), .Z(n16680) );
  XNOR U16730 ( .A(p_input[1024]), .B(p_input[832]), .Z(n16754) );
  XOR U16731 ( .A(n16742), .B(n16741), .Z(n16773) );
  XNOR U16732 ( .A(n16774), .B(n16748), .Z(n16741) );
  XNOR U16733 ( .A(n16737), .B(n16736), .Z(n16748) );
  XOR U16734 ( .A(n16775), .B(n16733), .Z(n16736) );
  XOR U16735 ( .A(p_input[1034]), .B(p_input[842]), .Z(n16733) );
  XNOR U16736 ( .A(p_input[1035]), .B(p_input[843]), .Z(n16775) );
  XOR U16737 ( .A(p_input[1036]), .B(p_input[844]), .Z(n16737) );
  XNOR U16738 ( .A(n16747), .B(n16738), .Z(n16774) );
  XOR U16739 ( .A(p_input[1025]), .B(p_input[833]), .Z(n16738) );
  XOR U16740 ( .A(n16776), .B(n16753), .Z(n16747) );
  XNOR U16741 ( .A(p_input[1039]), .B(p_input[847]), .Z(n16753) );
  XOR U16742 ( .A(n16744), .B(n16752), .Z(n16776) );
  XOR U16743 ( .A(n16777), .B(n16749), .Z(n16752) );
  XOR U16744 ( .A(p_input[1037]), .B(p_input[845]), .Z(n16749) );
  XNOR U16745 ( .A(p_input[1038]), .B(p_input[846]), .Z(n16777) );
  XOR U16746 ( .A(p_input[1033]), .B(p_input[841]), .Z(n16744) );
  XNOR U16747 ( .A(n16760), .B(n16759), .Z(n16742) );
  XNOR U16748 ( .A(n16778), .B(n16765), .Z(n16759) );
  XOR U16749 ( .A(p_input[1032]), .B(p_input[840]), .Z(n16765) );
  XOR U16750 ( .A(n16756), .B(n16764), .Z(n16778) );
  XOR U16751 ( .A(n16779), .B(n16761), .Z(n16764) );
  XOR U16752 ( .A(p_input[1030]), .B(p_input[838]), .Z(n16761) );
  XNOR U16753 ( .A(p_input[1031]), .B(p_input[839]), .Z(n16779) );
  XOR U16754 ( .A(p_input[1026]), .B(p_input[834]), .Z(n16756) );
  XNOR U16755 ( .A(n16770), .B(n16769), .Z(n16760) );
  XOR U16756 ( .A(n16780), .B(n16766), .Z(n16769) );
  XOR U16757 ( .A(p_input[1027]), .B(p_input[835]), .Z(n16766) );
  XNOR U16758 ( .A(p_input[1028]), .B(p_input[836]), .Z(n16780) );
  XOR U16759 ( .A(p_input[1029]), .B(p_input[837]), .Z(n16770) );
  XNOR U16760 ( .A(n16781), .B(n16782), .Z(n16677) );
  AND U16761 ( .A(n611), .B(n16783), .Z(n16782) );
  XNOR U16762 ( .A(n16784), .B(n16785), .Z(n611) );
  AND U16763 ( .A(n16786), .B(n16787), .Z(n16785) );
  XOR U16764 ( .A(n16784), .B(n16687), .Z(n16787) );
  XNOR U16765 ( .A(n16784), .B(n16641), .Z(n16786) );
  XOR U16766 ( .A(n16788), .B(n16789), .Z(n16784) );
  AND U16767 ( .A(n16790), .B(n16791), .Z(n16789) );
  XOR U16768 ( .A(n16788), .B(n16651), .Z(n16790) );
  XOR U16769 ( .A(n16792), .B(n16793), .Z(n16630) );
  AND U16770 ( .A(n615), .B(n16783), .Z(n16793) );
  XNOR U16771 ( .A(n16781), .B(n16792), .Z(n16783) );
  XNOR U16772 ( .A(n16794), .B(n16795), .Z(n615) );
  AND U16773 ( .A(n16796), .B(n16797), .Z(n16795) );
  XNOR U16774 ( .A(n16798), .B(n16794), .Z(n16797) );
  IV U16775 ( .A(n16687), .Z(n16798) );
  XNOR U16776 ( .A(n16799), .B(n16800), .Z(n16687) );
  AND U16777 ( .A(n618), .B(n16801), .Z(n16800) );
  XNOR U16778 ( .A(n16799), .B(n16802), .Z(n16801) );
  XNOR U16779 ( .A(n16641), .B(n16794), .Z(n16796) );
  XOR U16780 ( .A(n16803), .B(n16804), .Z(n16641) );
  AND U16781 ( .A(n626), .B(n16805), .Z(n16804) );
  XOR U16782 ( .A(n16788), .B(n16806), .Z(n16794) );
  AND U16783 ( .A(n16807), .B(n16791), .Z(n16806) );
  XNOR U16784 ( .A(n16700), .B(n16788), .Z(n16791) );
  XNOR U16785 ( .A(n16808), .B(n16809), .Z(n16700) );
  AND U16786 ( .A(n618), .B(n16810), .Z(n16809) );
  XOR U16787 ( .A(n16811), .B(n16808), .Z(n16810) );
  XNOR U16788 ( .A(n16812), .B(n16788), .Z(n16807) );
  IV U16789 ( .A(n16651), .Z(n16812) );
  XOR U16790 ( .A(n16813), .B(n16814), .Z(n16651) );
  AND U16791 ( .A(n626), .B(n16815), .Z(n16814) );
  XOR U16792 ( .A(n16816), .B(n16817), .Z(n16788) );
  AND U16793 ( .A(n16818), .B(n16819), .Z(n16817) );
  XNOR U16794 ( .A(n16725), .B(n16816), .Z(n16819) );
  XNOR U16795 ( .A(n16820), .B(n16821), .Z(n16725) );
  AND U16796 ( .A(n618), .B(n16822), .Z(n16821) );
  XNOR U16797 ( .A(n16823), .B(n16820), .Z(n16822) );
  XOR U16798 ( .A(n16816), .B(n16662), .Z(n16818) );
  XOR U16799 ( .A(n16824), .B(n16825), .Z(n16662) );
  AND U16800 ( .A(n626), .B(n16826), .Z(n16825) );
  XOR U16801 ( .A(n16827), .B(n16828), .Z(n16816) );
  AND U16802 ( .A(n16829), .B(n16830), .Z(n16828) );
  XNOR U16803 ( .A(n16827), .B(n16771), .Z(n16830) );
  XNOR U16804 ( .A(n16831), .B(n16832), .Z(n16771) );
  AND U16805 ( .A(n618), .B(n16833), .Z(n16832) );
  XOR U16806 ( .A(n16834), .B(n16831), .Z(n16833) );
  XNOR U16807 ( .A(n16835), .B(n16827), .Z(n16829) );
  IV U16808 ( .A(n16674), .Z(n16835) );
  XOR U16809 ( .A(n16836), .B(n16837), .Z(n16674) );
  AND U16810 ( .A(n626), .B(n16838), .Z(n16837) );
  AND U16811 ( .A(n16792), .B(n16781), .Z(n16827) );
  XNOR U16812 ( .A(n16839), .B(n16840), .Z(n16781) );
  AND U16813 ( .A(n618), .B(n16841), .Z(n16840) );
  XNOR U16814 ( .A(n16842), .B(n16839), .Z(n16841) );
  XNOR U16815 ( .A(n16843), .B(n16844), .Z(n618) );
  AND U16816 ( .A(n16845), .B(n16846), .Z(n16844) );
  XOR U16817 ( .A(n16802), .B(n16843), .Z(n16846) );
  AND U16818 ( .A(n16847), .B(n16848), .Z(n16802) );
  XOR U16819 ( .A(n16843), .B(n16799), .Z(n16845) );
  XNOR U16820 ( .A(n16849), .B(n16850), .Z(n16799) );
  AND U16821 ( .A(n622), .B(n16805), .Z(n16850) );
  XOR U16822 ( .A(n16803), .B(n16849), .Z(n16805) );
  XOR U16823 ( .A(n16851), .B(n16852), .Z(n16843) );
  AND U16824 ( .A(n16853), .B(n16854), .Z(n16852) );
  XNOR U16825 ( .A(n16851), .B(n16847), .Z(n16854) );
  IV U16826 ( .A(n16811), .Z(n16847) );
  XOR U16827 ( .A(n16855), .B(n16856), .Z(n16811) );
  XOR U16828 ( .A(n16857), .B(n16848), .Z(n16856) );
  AND U16829 ( .A(n16823), .B(n16858), .Z(n16848) );
  AND U16830 ( .A(n16859), .B(n16860), .Z(n16857) );
  XOR U16831 ( .A(n16861), .B(n16855), .Z(n16859) );
  XNOR U16832 ( .A(n16808), .B(n16851), .Z(n16853) );
  XNOR U16833 ( .A(n16862), .B(n16863), .Z(n16808) );
  AND U16834 ( .A(n622), .B(n16815), .Z(n16863) );
  XOR U16835 ( .A(n16862), .B(n16813), .Z(n16815) );
  XOR U16836 ( .A(n16864), .B(n16865), .Z(n16851) );
  AND U16837 ( .A(n16866), .B(n16867), .Z(n16865) );
  XNOR U16838 ( .A(n16864), .B(n16823), .Z(n16867) );
  XOR U16839 ( .A(n16868), .B(n16860), .Z(n16823) );
  XNOR U16840 ( .A(n16869), .B(n16855), .Z(n16860) );
  XOR U16841 ( .A(n16870), .B(n16871), .Z(n16855) );
  AND U16842 ( .A(n16872), .B(n16873), .Z(n16871) );
  XOR U16843 ( .A(n16874), .B(n16870), .Z(n16872) );
  XNOR U16844 ( .A(n16875), .B(n16876), .Z(n16869) );
  AND U16845 ( .A(n16877), .B(n16878), .Z(n16876) );
  XOR U16846 ( .A(n16875), .B(n16879), .Z(n16877) );
  XNOR U16847 ( .A(n16861), .B(n16858), .Z(n16868) );
  AND U16848 ( .A(n16880), .B(n16881), .Z(n16858) );
  XOR U16849 ( .A(n16882), .B(n16883), .Z(n16861) );
  AND U16850 ( .A(n16884), .B(n16885), .Z(n16883) );
  XOR U16851 ( .A(n16882), .B(n16886), .Z(n16884) );
  XNOR U16852 ( .A(n16820), .B(n16864), .Z(n16866) );
  XNOR U16853 ( .A(n16887), .B(n16888), .Z(n16820) );
  AND U16854 ( .A(n622), .B(n16826), .Z(n16888) );
  XOR U16855 ( .A(n16887), .B(n16824), .Z(n16826) );
  XOR U16856 ( .A(n16889), .B(n16890), .Z(n16864) );
  AND U16857 ( .A(n16891), .B(n16892), .Z(n16890) );
  XNOR U16858 ( .A(n16889), .B(n16880), .Z(n16892) );
  IV U16859 ( .A(n16834), .Z(n16880) );
  XNOR U16860 ( .A(n16893), .B(n16873), .Z(n16834) );
  XNOR U16861 ( .A(n16894), .B(n16879), .Z(n16873) );
  XOR U16862 ( .A(n16895), .B(n16896), .Z(n16879) );
  NOR U16863 ( .A(n16897), .B(n16898), .Z(n16896) );
  XNOR U16864 ( .A(n16895), .B(n16899), .Z(n16897) );
  XNOR U16865 ( .A(n16878), .B(n16870), .Z(n16894) );
  XOR U16866 ( .A(n16900), .B(n16901), .Z(n16870) );
  AND U16867 ( .A(n16902), .B(n16903), .Z(n16901) );
  XNOR U16868 ( .A(n16900), .B(n16904), .Z(n16902) );
  XNOR U16869 ( .A(n16905), .B(n16875), .Z(n16878) );
  XOR U16870 ( .A(n16906), .B(n16907), .Z(n16875) );
  AND U16871 ( .A(n16908), .B(n16909), .Z(n16907) );
  XOR U16872 ( .A(n16906), .B(n16910), .Z(n16908) );
  XNOR U16873 ( .A(n16911), .B(n16912), .Z(n16905) );
  NOR U16874 ( .A(n16913), .B(n16914), .Z(n16912) );
  XOR U16875 ( .A(n16911), .B(n16915), .Z(n16913) );
  XNOR U16876 ( .A(n16874), .B(n16881), .Z(n16893) );
  NOR U16877 ( .A(n16842), .B(n16916), .Z(n16881) );
  XOR U16878 ( .A(n16886), .B(n16885), .Z(n16874) );
  XNOR U16879 ( .A(n16917), .B(n16882), .Z(n16885) );
  XOR U16880 ( .A(n16918), .B(n16919), .Z(n16882) );
  AND U16881 ( .A(n16920), .B(n16921), .Z(n16919) );
  XOR U16882 ( .A(n16918), .B(n16922), .Z(n16920) );
  XNOR U16883 ( .A(n16923), .B(n16924), .Z(n16917) );
  NOR U16884 ( .A(n16925), .B(n16926), .Z(n16924) );
  XNOR U16885 ( .A(n16923), .B(n16927), .Z(n16925) );
  XOR U16886 ( .A(n16928), .B(n16929), .Z(n16886) );
  NOR U16887 ( .A(n16930), .B(n16931), .Z(n16929) );
  XNOR U16888 ( .A(n16928), .B(n16932), .Z(n16930) );
  XNOR U16889 ( .A(n16831), .B(n16889), .Z(n16891) );
  XNOR U16890 ( .A(n16933), .B(n16934), .Z(n16831) );
  AND U16891 ( .A(n622), .B(n16838), .Z(n16934) );
  XOR U16892 ( .A(n16933), .B(n16836), .Z(n16838) );
  AND U16893 ( .A(n16839), .B(n16842), .Z(n16889) );
  XOR U16894 ( .A(n16935), .B(n16916), .Z(n16842) );
  XNOR U16895 ( .A(p_input[1024]), .B(p_input[848]), .Z(n16916) );
  XOR U16896 ( .A(n16904), .B(n16903), .Z(n16935) );
  XNOR U16897 ( .A(n16936), .B(n16910), .Z(n16903) );
  XNOR U16898 ( .A(n16899), .B(n16898), .Z(n16910) );
  XOR U16899 ( .A(n16937), .B(n16895), .Z(n16898) );
  XOR U16900 ( .A(p_input[1034]), .B(p_input[858]), .Z(n16895) );
  XNOR U16901 ( .A(p_input[1035]), .B(p_input[859]), .Z(n16937) );
  XOR U16902 ( .A(p_input[1036]), .B(p_input[860]), .Z(n16899) );
  XNOR U16903 ( .A(n16909), .B(n16900), .Z(n16936) );
  XOR U16904 ( .A(p_input[1025]), .B(p_input[849]), .Z(n16900) );
  XOR U16905 ( .A(n16938), .B(n16915), .Z(n16909) );
  XNOR U16906 ( .A(p_input[1039]), .B(p_input[863]), .Z(n16915) );
  XOR U16907 ( .A(n16906), .B(n16914), .Z(n16938) );
  XOR U16908 ( .A(n16939), .B(n16911), .Z(n16914) );
  XOR U16909 ( .A(p_input[1037]), .B(p_input[861]), .Z(n16911) );
  XNOR U16910 ( .A(p_input[1038]), .B(p_input[862]), .Z(n16939) );
  XOR U16911 ( .A(p_input[1033]), .B(p_input[857]), .Z(n16906) );
  XNOR U16912 ( .A(n16922), .B(n16921), .Z(n16904) );
  XNOR U16913 ( .A(n16940), .B(n16927), .Z(n16921) );
  XOR U16914 ( .A(p_input[1032]), .B(p_input[856]), .Z(n16927) );
  XOR U16915 ( .A(n16918), .B(n16926), .Z(n16940) );
  XOR U16916 ( .A(n16941), .B(n16923), .Z(n16926) );
  XOR U16917 ( .A(p_input[1030]), .B(p_input[854]), .Z(n16923) );
  XNOR U16918 ( .A(p_input[1031]), .B(p_input[855]), .Z(n16941) );
  XOR U16919 ( .A(p_input[1026]), .B(p_input[850]), .Z(n16918) );
  XNOR U16920 ( .A(n16932), .B(n16931), .Z(n16922) );
  XOR U16921 ( .A(n16942), .B(n16928), .Z(n16931) );
  XOR U16922 ( .A(p_input[1027]), .B(p_input[851]), .Z(n16928) );
  XNOR U16923 ( .A(p_input[1028]), .B(p_input[852]), .Z(n16942) );
  XOR U16924 ( .A(p_input[1029]), .B(p_input[853]), .Z(n16932) );
  XNOR U16925 ( .A(n16943), .B(n16944), .Z(n16839) );
  AND U16926 ( .A(n622), .B(n16945), .Z(n16944) );
  XNOR U16927 ( .A(n16946), .B(n16947), .Z(n622) );
  AND U16928 ( .A(n16948), .B(n16949), .Z(n16947) );
  XOR U16929 ( .A(n16946), .B(n16849), .Z(n16949) );
  XNOR U16930 ( .A(n16946), .B(n16803), .Z(n16948) );
  XOR U16931 ( .A(n16950), .B(n16951), .Z(n16946) );
  AND U16932 ( .A(n16952), .B(n16953), .Z(n16951) );
  XOR U16933 ( .A(n16950), .B(n16813), .Z(n16952) );
  XOR U16934 ( .A(n16954), .B(n16955), .Z(n16792) );
  AND U16935 ( .A(n626), .B(n16945), .Z(n16955) );
  XNOR U16936 ( .A(n16943), .B(n16954), .Z(n16945) );
  XNOR U16937 ( .A(n16956), .B(n16957), .Z(n626) );
  AND U16938 ( .A(n16958), .B(n16959), .Z(n16957) );
  XNOR U16939 ( .A(n16960), .B(n16956), .Z(n16959) );
  IV U16940 ( .A(n16849), .Z(n16960) );
  XNOR U16941 ( .A(n16961), .B(n16962), .Z(n16849) );
  AND U16942 ( .A(n629), .B(n16963), .Z(n16962) );
  XNOR U16943 ( .A(n16961), .B(n16964), .Z(n16963) );
  XNOR U16944 ( .A(n16803), .B(n16956), .Z(n16958) );
  XOR U16945 ( .A(n16965), .B(n16966), .Z(n16803) );
  AND U16946 ( .A(n637), .B(n16967), .Z(n16966) );
  XOR U16947 ( .A(n16950), .B(n16968), .Z(n16956) );
  AND U16948 ( .A(n16969), .B(n16953), .Z(n16968) );
  XNOR U16949 ( .A(n16862), .B(n16950), .Z(n16953) );
  XNOR U16950 ( .A(n16970), .B(n16971), .Z(n16862) );
  AND U16951 ( .A(n629), .B(n16972), .Z(n16971) );
  XOR U16952 ( .A(n16973), .B(n16970), .Z(n16972) );
  XNOR U16953 ( .A(n16974), .B(n16950), .Z(n16969) );
  IV U16954 ( .A(n16813), .Z(n16974) );
  XOR U16955 ( .A(n16975), .B(n16976), .Z(n16813) );
  AND U16956 ( .A(n637), .B(n16977), .Z(n16976) );
  XOR U16957 ( .A(n16978), .B(n16979), .Z(n16950) );
  AND U16958 ( .A(n16980), .B(n16981), .Z(n16979) );
  XNOR U16959 ( .A(n16887), .B(n16978), .Z(n16981) );
  XNOR U16960 ( .A(n16982), .B(n16983), .Z(n16887) );
  AND U16961 ( .A(n629), .B(n16984), .Z(n16983) );
  XNOR U16962 ( .A(n16985), .B(n16982), .Z(n16984) );
  XOR U16963 ( .A(n16978), .B(n16824), .Z(n16980) );
  XOR U16964 ( .A(n16986), .B(n16987), .Z(n16824) );
  AND U16965 ( .A(n637), .B(n16988), .Z(n16987) );
  XOR U16966 ( .A(n16989), .B(n16990), .Z(n16978) );
  AND U16967 ( .A(n16991), .B(n16992), .Z(n16990) );
  XNOR U16968 ( .A(n16989), .B(n16933), .Z(n16992) );
  XNOR U16969 ( .A(n16993), .B(n16994), .Z(n16933) );
  AND U16970 ( .A(n629), .B(n16995), .Z(n16994) );
  XOR U16971 ( .A(n16996), .B(n16993), .Z(n16995) );
  XNOR U16972 ( .A(n16997), .B(n16989), .Z(n16991) );
  IV U16973 ( .A(n16836), .Z(n16997) );
  XOR U16974 ( .A(n16998), .B(n16999), .Z(n16836) );
  AND U16975 ( .A(n637), .B(n17000), .Z(n16999) );
  AND U16976 ( .A(n16954), .B(n16943), .Z(n16989) );
  XNOR U16977 ( .A(n17001), .B(n17002), .Z(n16943) );
  AND U16978 ( .A(n629), .B(n17003), .Z(n17002) );
  XNOR U16979 ( .A(n17004), .B(n17001), .Z(n17003) );
  XNOR U16980 ( .A(n17005), .B(n17006), .Z(n629) );
  AND U16981 ( .A(n17007), .B(n17008), .Z(n17006) );
  XOR U16982 ( .A(n16964), .B(n17005), .Z(n17008) );
  AND U16983 ( .A(n17009), .B(n17010), .Z(n16964) );
  XOR U16984 ( .A(n17005), .B(n16961), .Z(n17007) );
  XNOR U16985 ( .A(n17011), .B(n17012), .Z(n16961) );
  AND U16986 ( .A(n633), .B(n16967), .Z(n17012) );
  XOR U16987 ( .A(n16965), .B(n17011), .Z(n16967) );
  XOR U16988 ( .A(n17013), .B(n17014), .Z(n17005) );
  AND U16989 ( .A(n17015), .B(n17016), .Z(n17014) );
  XNOR U16990 ( .A(n17013), .B(n17009), .Z(n17016) );
  IV U16991 ( .A(n16973), .Z(n17009) );
  XOR U16992 ( .A(n17017), .B(n17018), .Z(n16973) );
  XOR U16993 ( .A(n17019), .B(n17010), .Z(n17018) );
  AND U16994 ( .A(n16985), .B(n17020), .Z(n17010) );
  AND U16995 ( .A(n17021), .B(n17022), .Z(n17019) );
  XOR U16996 ( .A(n17023), .B(n17017), .Z(n17021) );
  XNOR U16997 ( .A(n16970), .B(n17013), .Z(n17015) );
  XNOR U16998 ( .A(n17024), .B(n17025), .Z(n16970) );
  AND U16999 ( .A(n633), .B(n16977), .Z(n17025) );
  XOR U17000 ( .A(n17024), .B(n16975), .Z(n16977) );
  XOR U17001 ( .A(n17026), .B(n17027), .Z(n17013) );
  AND U17002 ( .A(n17028), .B(n17029), .Z(n17027) );
  XNOR U17003 ( .A(n17026), .B(n16985), .Z(n17029) );
  XOR U17004 ( .A(n17030), .B(n17022), .Z(n16985) );
  XNOR U17005 ( .A(n17031), .B(n17017), .Z(n17022) );
  XOR U17006 ( .A(n17032), .B(n17033), .Z(n17017) );
  AND U17007 ( .A(n17034), .B(n17035), .Z(n17033) );
  XOR U17008 ( .A(n17036), .B(n17032), .Z(n17034) );
  XNOR U17009 ( .A(n17037), .B(n17038), .Z(n17031) );
  AND U17010 ( .A(n17039), .B(n17040), .Z(n17038) );
  XOR U17011 ( .A(n17037), .B(n17041), .Z(n17039) );
  XNOR U17012 ( .A(n17023), .B(n17020), .Z(n17030) );
  AND U17013 ( .A(n17042), .B(n17043), .Z(n17020) );
  XOR U17014 ( .A(n17044), .B(n17045), .Z(n17023) );
  AND U17015 ( .A(n17046), .B(n17047), .Z(n17045) );
  XOR U17016 ( .A(n17044), .B(n17048), .Z(n17046) );
  XNOR U17017 ( .A(n16982), .B(n17026), .Z(n17028) );
  XNOR U17018 ( .A(n17049), .B(n17050), .Z(n16982) );
  AND U17019 ( .A(n633), .B(n16988), .Z(n17050) );
  XOR U17020 ( .A(n17049), .B(n16986), .Z(n16988) );
  XOR U17021 ( .A(n17051), .B(n17052), .Z(n17026) );
  AND U17022 ( .A(n17053), .B(n17054), .Z(n17052) );
  XNOR U17023 ( .A(n17051), .B(n17042), .Z(n17054) );
  IV U17024 ( .A(n16996), .Z(n17042) );
  XNOR U17025 ( .A(n17055), .B(n17035), .Z(n16996) );
  XNOR U17026 ( .A(n17056), .B(n17041), .Z(n17035) );
  XOR U17027 ( .A(n17057), .B(n17058), .Z(n17041) );
  NOR U17028 ( .A(n17059), .B(n17060), .Z(n17058) );
  XNOR U17029 ( .A(n17057), .B(n17061), .Z(n17059) );
  XNOR U17030 ( .A(n17040), .B(n17032), .Z(n17056) );
  XOR U17031 ( .A(n17062), .B(n17063), .Z(n17032) );
  AND U17032 ( .A(n17064), .B(n17065), .Z(n17063) );
  XNOR U17033 ( .A(n17062), .B(n17066), .Z(n17064) );
  XNOR U17034 ( .A(n17067), .B(n17037), .Z(n17040) );
  XOR U17035 ( .A(n17068), .B(n17069), .Z(n17037) );
  AND U17036 ( .A(n17070), .B(n17071), .Z(n17069) );
  XOR U17037 ( .A(n17068), .B(n17072), .Z(n17070) );
  XNOR U17038 ( .A(n17073), .B(n17074), .Z(n17067) );
  NOR U17039 ( .A(n17075), .B(n17076), .Z(n17074) );
  XOR U17040 ( .A(n17073), .B(n17077), .Z(n17075) );
  XNOR U17041 ( .A(n17036), .B(n17043), .Z(n17055) );
  NOR U17042 ( .A(n17004), .B(n17078), .Z(n17043) );
  XOR U17043 ( .A(n17048), .B(n17047), .Z(n17036) );
  XNOR U17044 ( .A(n17079), .B(n17044), .Z(n17047) );
  XOR U17045 ( .A(n17080), .B(n17081), .Z(n17044) );
  AND U17046 ( .A(n17082), .B(n17083), .Z(n17081) );
  XOR U17047 ( .A(n17080), .B(n17084), .Z(n17082) );
  XNOR U17048 ( .A(n17085), .B(n17086), .Z(n17079) );
  NOR U17049 ( .A(n17087), .B(n17088), .Z(n17086) );
  XNOR U17050 ( .A(n17085), .B(n17089), .Z(n17087) );
  XOR U17051 ( .A(n17090), .B(n17091), .Z(n17048) );
  NOR U17052 ( .A(n17092), .B(n17093), .Z(n17091) );
  XNOR U17053 ( .A(n17090), .B(n17094), .Z(n17092) );
  XNOR U17054 ( .A(n16993), .B(n17051), .Z(n17053) );
  XNOR U17055 ( .A(n17095), .B(n17096), .Z(n16993) );
  AND U17056 ( .A(n633), .B(n17000), .Z(n17096) );
  XOR U17057 ( .A(n17095), .B(n16998), .Z(n17000) );
  AND U17058 ( .A(n17001), .B(n17004), .Z(n17051) );
  XOR U17059 ( .A(n17097), .B(n17078), .Z(n17004) );
  XNOR U17060 ( .A(p_input[1024]), .B(p_input[864]), .Z(n17078) );
  XOR U17061 ( .A(n17066), .B(n17065), .Z(n17097) );
  XNOR U17062 ( .A(n17098), .B(n17072), .Z(n17065) );
  XNOR U17063 ( .A(n17061), .B(n17060), .Z(n17072) );
  XOR U17064 ( .A(n17099), .B(n17057), .Z(n17060) );
  XOR U17065 ( .A(p_input[1034]), .B(p_input[874]), .Z(n17057) );
  XNOR U17066 ( .A(p_input[1035]), .B(p_input[875]), .Z(n17099) );
  XOR U17067 ( .A(p_input[1036]), .B(p_input[876]), .Z(n17061) );
  XNOR U17068 ( .A(n17071), .B(n17062), .Z(n17098) );
  XOR U17069 ( .A(p_input[1025]), .B(p_input[865]), .Z(n17062) );
  XOR U17070 ( .A(n17100), .B(n17077), .Z(n17071) );
  XNOR U17071 ( .A(p_input[1039]), .B(p_input[879]), .Z(n17077) );
  XOR U17072 ( .A(n17068), .B(n17076), .Z(n17100) );
  XOR U17073 ( .A(n17101), .B(n17073), .Z(n17076) );
  XOR U17074 ( .A(p_input[1037]), .B(p_input[877]), .Z(n17073) );
  XNOR U17075 ( .A(p_input[1038]), .B(p_input[878]), .Z(n17101) );
  XOR U17076 ( .A(p_input[1033]), .B(p_input[873]), .Z(n17068) );
  XNOR U17077 ( .A(n17084), .B(n17083), .Z(n17066) );
  XNOR U17078 ( .A(n17102), .B(n17089), .Z(n17083) );
  XOR U17079 ( .A(p_input[1032]), .B(p_input[872]), .Z(n17089) );
  XOR U17080 ( .A(n17080), .B(n17088), .Z(n17102) );
  XOR U17081 ( .A(n17103), .B(n17085), .Z(n17088) );
  XOR U17082 ( .A(p_input[1030]), .B(p_input[870]), .Z(n17085) );
  XNOR U17083 ( .A(p_input[1031]), .B(p_input[871]), .Z(n17103) );
  XOR U17084 ( .A(p_input[1026]), .B(p_input[866]), .Z(n17080) );
  XNOR U17085 ( .A(n17094), .B(n17093), .Z(n17084) );
  XOR U17086 ( .A(n17104), .B(n17090), .Z(n17093) );
  XOR U17087 ( .A(p_input[1027]), .B(p_input[867]), .Z(n17090) );
  XNOR U17088 ( .A(p_input[1028]), .B(p_input[868]), .Z(n17104) );
  XOR U17089 ( .A(p_input[1029]), .B(p_input[869]), .Z(n17094) );
  XNOR U17090 ( .A(n17105), .B(n17106), .Z(n17001) );
  AND U17091 ( .A(n633), .B(n17107), .Z(n17106) );
  XNOR U17092 ( .A(n17108), .B(n17109), .Z(n633) );
  AND U17093 ( .A(n17110), .B(n17111), .Z(n17109) );
  XOR U17094 ( .A(n17108), .B(n17011), .Z(n17111) );
  XNOR U17095 ( .A(n17108), .B(n16965), .Z(n17110) );
  XOR U17096 ( .A(n17112), .B(n17113), .Z(n17108) );
  AND U17097 ( .A(n17114), .B(n17115), .Z(n17113) );
  XOR U17098 ( .A(n17112), .B(n16975), .Z(n17114) );
  XOR U17099 ( .A(n17116), .B(n17117), .Z(n16954) );
  AND U17100 ( .A(n637), .B(n17107), .Z(n17117) );
  XNOR U17101 ( .A(n17105), .B(n17116), .Z(n17107) );
  XNOR U17102 ( .A(n17118), .B(n17119), .Z(n637) );
  AND U17103 ( .A(n17120), .B(n17121), .Z(n17119) );
  XNOR U17104 ( .A(n17122), .B(n17118), .Z(n17121) );
  IV U17105 ( .A(n17011), .Z(n17122) );
  XNOR U17106 ( .A(n17123), .B(n17124), .Z(n17011) );
  AND U17107 ( .A(n640), .B(n17125), .Z(n17124) );
  XNOR U17108 ( .A(n17123), .B(n17126), .Z(n17125) );
  XNOR U17109 ( .A(n16965), .B(n17118), .Z(n17120) );
  XOR U17110 ( .A(n17127), .B(n17128), .Z(n16965) );
  AND U17111 ( .A(n648), .B(n17129), .Z(n17128) );
  XOR U17112 ( .A(n17112), .B(n17130), .Z(n17118) );
  AND U17113 ( .A(n17131), .B(n17115), .Z(n17130) );
  XNOR U17114 ( .A(n17024), .B(n17112), .Z(n17115) );
  XNOR U17115 ( .A(n17132), .B(n17133), .Z(n17024) );
  AND U17116 ( .A(n640), .B(n17134), .Z(n17133) );
  XOR U17117 ( .A(n17135), .B(n17132), .Z(n17134) );
  XNOR U17118 ( .A(n17136), .B(n17112), .Z(n17131) );
  IV U17119 ( .A(n16975), .Z(n17136) );
  XOR U17120 ( .A(n17137), .B(n17138), .Z(n16975) );
  AND U17121 ( .A(n648), .B(n17139), .Z(n17138) );
  XOR U17122 ( .A(n17140), .B(n17141), .Z(n17112) );
  AND U17123 ( .A(n17142), .B(n17143), .Z(n17141) );
  XNOR U17124 ( .A(n17049), .B(n17140), .Z(n17143) );
  XNOR U17125 ( .A(n17144), .B(n17145), .Z(n17049) );
  AND U17126 ( .A(n640), .B(n17146), .Z(n17145) );
  XNOR U17127 ( .A(n17147), .B(n17144), .Z(n17146) );
  XOR U17128 ( .A(n17140), .B(n16986), .Z(n17142) );
  XOR U17129 ( .A(n17148), .B(n17149), .Z(n16986) );
  AND U17130 ( .A(n648), .B(n17150), .Z(n17149) );
  XOR U17131 ( .A(n17151), .B(n17152), .Z(n17140) );
  AND U17132 ( .A(n17153), .B(n17154), .Z(n17152) );
  XNOR U17133 ( .A(n17151), .B(n17095), .Z(n17154) );
  XNOR U17134 ( .A(n17155), .B(n17156), .Z(n17095) );
  AND U17135 ( .A(n640), .B(n17157), .Z(n17156) );
  XOR U17136 ( .A(n17158), .B(n17155), .Z(n17157) );
  XNOR U17137 ( .A(n17159), .B(n17151), .Z(n17153) );
  IV U17138 ( .A(n16998), .Z(n17159) );
  XOR U17139 ( .A(n17160), .B(n17161), .Z(n16998) );
  AND U17140 ( .A(n648), .B(n17162), .Z(n17161) );
  AND U17141 ( .A(n17116), .B(n17105), .Z(n17151) );
  XNOR U17142 ( .A(n17163), .B(n17164), .Z(n17105) );
  AND U17143 ( .A(n640), .B(n17165), .Z(n17164) );
  XNOR U17144 ( .A(n17166), .B(n17163), .Z(n17165) );
  XNOR U17145 ( .A(n17167), .B(n17168), .Z(n640) );
  AND U17146 ( .A(n17169), .B(n17170), .Z(n17168) );
  XOR U17147 ( .A(n17126), .B(n17167), .Z(n17170) );
  AND U17148 ( .A(n17171), .B(n17172), .Z(n17126) );
  XOR U17149 ( .A(n17167), .B(n17123), .Z(n17169) );
  XNOR U17150 ( .A(n17173), .B(n17174), .Z(n17123) );
  AND U17151 ( .A(n644), .B(n17129), .Z(n17174) );
  XOR U17152 ( .A(n17127), .B(n17173), .Z(n17129) );
  XOR U17153 ( .A(n17175), .B(n17176), .Z(n17167) );
  AND U17154 ( .A(n17177), .B(n17178), .Z(n17176) );
  XNOR U17155 ( .A(n17175), .B(n17171), .Z(n17178) );
  IV U17156 ( .A(n17135), .Z(n17171) );
  XOR U17157 ( .A(n17179), .B(n17180), .Z(n17135) );
  XOR U17158 ( .A(n17181), .B(n17172), .Z(n17180) );
  AND U17159 ( .A(n17147), .B(n17182), .Z(n17172) );
  AND U17160 ( .A(n17183), .B(n17184), .Z(n17181) );
  XOR U17161 ( .A(n17185), .B(n17179), .Z(n17183) );
  XNOR U17162 ( .A(n17132), .B(n17175), .Z(n17177) );
  XNOR U17163 ( .A(n17186), .B(n17187), .Z(n17132) );
  AND U17164 ( .A(n644), .B(n17139), .Z(n17187) );
  XOR U17165 ( .A(n17186), .B(n17137), .Z(n17139) );
  XOR U17166 ( .A(n17188), .B(n17189), .Z(n17175) );
  AND U17167 ( .A(n17190), .B(n17191), .Z(n17189) );
  XNOR U17168 ( .A(n17188), .B(n17147), .Z(n17191) );
  XOR U17169 ( .A(n17192), .B(n17184), .Z(n17147) );
  XNOR U17170 ( .A(n17193), .B(n17179), .Z(n17184) );
  XOR U17171 ( .A(n17194), .B(n17195), .Z(n17179) );
  AND U17172 ( .A(n17196), .B(n17197), .Z(n17195) );
  XOR U17173 ( .A(n17198), .B(n17194), .Z(n17196) );
  XNOR U17174 ( .A(n17199), .B(n17200), .Z(n17193) );
  AND U17175 ( .A(n17201), .B(n17202), .Z(n17200) );
  XOR U17176 ( .A(n17199), .B(n17203), .Z(n17201) );
  XNOR U17177 ( .A(n17185), .B(n17182), .Z(n17192) );
  AND U17178 ( .A(n17204), .B(n17205), .Z(n17182) );
  XOR U17179 ( .A(n17206), .B(n17207), .Z(n17185) );
  AND U17180 ( .A(n17208), .B(n17209), .Z(n17207) );
  XOR U17181 ( .A(n17206), .B(n17210), .Z(n17208) );
  XNOR U17182 ( .A(n17144), .B(n17188), .Z(n17190) );
  XNOR U17183 ( .A(n17211), .B(n17212), .Z(n17144) );
  AND U17184 ( .A(n644), .B(n17150), .Z(n17212) );
  XOR U17185 ( .A(n17211), .B(n17148), .Z(n17150) );
  XOR U17186 ( .A(n17213), .B(n17214), .Z(n17188) );
  AND U17187 ( .A(n17215), .B(n17216), .Z(n17214) );
  XNOR U17188 ( .A(n17213), .B(n17204), .Z(n17216) );
  IV U17189 ( .A(n17158), .Z(n17204) );
  XNOR U17190 ( .A(n17217), .B(n17197), .Z(n17158) );
  XNOR U17191 ( .A(n17218), .B(n17203), .Z(n17197) );
  XOR U17192 ( .A(n17219), .B(n17220), .Z(n17203) );
  NOR U17193 ( .A(n17221), .B(n17222), .Z(n17220) );
  XNOR U17194 ( .A(n17219), .B(n17223), .Z(n17221) );
  XNOR U17195 ( .A(n17202), .B(n17194), .Z(n17218) );
  XOR U17196 ( .A(n17224), .B(n17225), .Z(n17194) );
  AND U17197 ( .A(n17226), .B(n17227), .Z(n17225) );
  XNOR U17198 ( .A(n17224), .B(n17228), .Z(n17226) );
  XNOR U17199 ( .A(n17229), .B(n17199), .Z(n17202) );
  XOR U17200 ( .A(n17230), .B(n17231), .Z(n17199) );
  AND U17201 ( .A(n17232), .B(n17233), .Z(n17231) );
  XOR U17202 ( .A(n17230), .B(n17234), .Z(n17232) );
  XNOR U17203 ( .A(n17235), .B(n17236), .Z(n17229) );
  NOR U17204 ( .A(n17237), .B(n17238), .Z(n17236) );
  XOR U17205 ( .A(n17235), .B(n17239), .Z(n17237) );
  XNOR U17206 ( .A(n17198), .B(n17205), .Z(n17217) );
  NOR U17207 ( .A(n17166), .B(n17240), .Z(n17205) );
  XOR U17208 ( .A(n17210), .B(n17209), .Z(n17198) );
  XNOR U17209 ( .A(n17241), .B(n17206), .Z(n17209) );
  XOR U17210 ( .A(n17242), .B(n17243), .Z(n17206) );
  AND U17211 ( .A(n17244), .B(n17245), .Z(n17243) );
  XOR U17212 ( .A(n17242), .B(n17246), .Z(n17244) );
  XNOR U17213 ( .A(n17247), .B(n17248), .Z(n17241) );
  NOR U17214 ( .A(n17249), .B(n17250), .Z(n17248) );
  XNOR U17215 ( .A(n17247), .B(n17251), .Z(n17249) );
  XOR U17216 ( .A(n17252), .B(n17253), .Z(n17210) );
  NOR U17217 ( .A(n17254), .B(n17255), .Z(n17253) );
  XNOR U17218 ( .A(n17252), .B(n17256), .Z(n17254) );
  XNOR U17219 ( .A(n17155), .B(n17213), .Z(n17215) );
  XNOR U17220 ( .A(n17257), .B(n17258), .Z(n17155) );
  AND U17221 ( .A(n644), .B(n17162), .Z(n17258) );
  XOR U17222 ( .A(n17257), .B(n17160), .Z(n17162) );
  AND U17223 ( .A(n17163), .B(n17166), .Z(n17213) );
  XOR U17224 ( .A(n17259), .B(n17240), .Z(n17166) );
  XNOR U17225 ( .A(p_input[1024]), .B(p_input[880]), .Z(n17240) );
  XOR U17226 ( .A(n17228), .B(n17227), .Z(n17259) );
  XNOR U17227 ( .A(n17260), .B(n17234), .Z(n17227) );
  XNOR U17228 ( .A(n17223), .B(n17222), .Z(n17234) );
  XOR U17229 ( .A(n17261), .B(n17219), .Z(n17222) );
  XOR U17230 ( .A(p_input[1034]), .B(p_input[890]), .Z(n17219) );
  XNOR U17231 ( .A(p_input[1035]), .B(p_input[891]), .Z(n17261) );
  XOR U17232 ( .A(p_input[1036]), .B(p_input[892]), .Z(n17223) );
  XNOR U17233 ( .A(n17233), .B(n17224), .Z(n17260) );
  XOR U17234 ( .A(p_input[1025]), .B(p_input[881]), .Z(n17224) );
  XOR U17235 ( .A(n17262), .B(n17239), .Z(n17233) );
  XNOR U17236 ( .A(p_input[1039]), .B(p_input[895]), .Z(n17239) );
  XOR U17237 ( .A(n17230), .B(n17238), .Z(n17262) );
  XOR U17238 ( .A(n17263), .B(n17235), .Z(n17238) );
  XOR U17239 ( .A(p_input[1037]), .B(p_input[893]), .Z(n17235) );
  XNOR U17240 ( .A(p_input[1038]), .B(p_input[894]), .Z(n17263) );
  XOR U17241 ( .A(p_input[1033]), .B(p_input[889]), .Z(n17230) );
  XNOR U17242 ( .A(n17246), .B(n17245), .Z(n17228) );
  XNOR U17243 ( .A(n17264), .B(n17251), .Z(n17245) );
  XOR U17244 ( .A(p_input[1032]), .B(p_input[888]), .Z(n17251) );
  XOR U17245 ( .A(n17242), .B(n17250), .Z(n17264) );
  XOR U17246 ( .A(n17265), .B(n17247), .Z(n17250) );
  XOR U17247 ( .A(p_input[1030]), .B(p_input[886]), .Z(n17247) );
  XNOR U17248 ( .A(p_input[1031]), .B(p_input[887]), .Z(n17265) );
  XOR U17249 ( .A(p_input[1026]), .B(p_input[882]), .Z(n17242) );
  XNOR U17250 ( .A(n17256), .B(n17255), .Z(n17246) );
  XOR U17251 ( .A(n17266), .B(n17252), .Z(n17255) );
  XOR U17252 ( .A(p_input[1027]), .B(p_input[883]), .Z(n17252) );
  XNOR U17253 ( .A(p_input[1028]), .B(p_input[884]), .Z(n17266) );
  XOR U17254 ( .A(p_input[1029]), .B(p_input[885]), .Z(n17256) );
  XNOR U17255 ( .A(n17267), .B(n17268), .Z(n17163) );
  AND U17256 ( .A(n644), .B(n17269), .Z(n17268) );
  XNOR U17257 ( .A(n17270), .B(n17271), .Z(n644) );
  AND U17258 ( .A(n17272), .B(n17273), .Z(n17271) );
  XOR U17259 ( .A(n17270), .B(n17173), .Z(n17273) );
  XNOR U17260 ( .A(n17270), .B(n17127), .Z(n17272) );
  XOR U17261 ( .A(n17274), .B(n17275), .Z(n17270) );
  AND U17262 ( .A(n17276), .B(n17277), .Z(n17275) );
  XOR U17263 ( .A(n17274), .B(n17137), .Z(n17276) );
  XOR U17264 ( .A(n17278), .B(n17279), .Z(n17116) );
  AND U17265 ( .A(n648), .B(n17269), .Z(n17279) );
  XNOR U17266 ( .A(n17267), .B(n17278), .Z(n17269) );
  XNOR U17267 ( .A(n17280), .B(n17281), .Z(n648) );
  AND U17268 ( .A(n17282), .B(n17283), .Z(n17281) );
  XNOR U17269 ( .A(n17284), .B(n17280), .Z(n17283) );
  IV U17270 ( .A(n17173), .Z(n17284) );
  XNOR U17271 ( .A(n17285), .B(n17286), .Z(n17173) );
  AND U17272 ( .A(n651), .B(n17287), .Z(n17286) );
  XNOR U17273 ( .A(n17285), .B(n17288), .Z(n17287) );
  XNOR U17274 ( .A(n17127), .B(n17280), .Z(n17282) );
  XNOR U17275 ( .A(n17289), .B(n17290), .Z(n17127) );
  AND U17276 ( .A(n659), .B(n17291), .Z(n17290) );
  XNOR U17277 ( .A(n17292), .B(n17293), .Z(n17291) );
  XOR U17278 ( .A(n17274), .B(n17294), .Z(n17280) );
  AND U17279 ( .A(n17295), .B(n17277), .Z(n17294) );
  XNOR U17280 ( .A(n17186), .B(n17274), .Z(n17277) );
  XNOR U17281 ( .A(n17296), .B(n17297), .Z(n17186) );
  AND U17282 ( .A(n651), .B(n17298), .Z(n17297) );
  XOR U17283 ( .A(n17299), .B(n17296), .Z(n17298) );
  XNOR U17284 ( .A(n17300), .B(n17274), .Z(n17295) );
  IV U17285 ( .A(n17137), .Z(n17300) );
  XOR U17286 ( .A(n17301), .B(n17302), .Z(n17137) );
  AND U17287 ( .A(n659), .B(n17303), .Z(n17302) );
  XOR U17288 ( .A(n17304), .B(n17305), .Z(n17274) );
  AND U17289 ( .A(n17306), .B(n17307), .Z(n17305) );
  XNOR U17290 ( .A(n17211), .B(n17304), .Z(n17307) );
  XNOR U17291 ( .A(n17308), .B(n17309), .Z(n17211) );
  AND U17292 ( .A(n651), .B(n17310), .Z(n17309) );
  XNOR U17293 ( .A(n17311), .B(n17308), .Z(n17310) );
  XOR U17294 ( .A(n17304), .B(n17148), .Z(n17306) );
  XOR U17295 ( .A(n17312), .B(n17313), .Z(n17148) );
  AND U17296 ( .A(n659), .B(n17314), .Z(n17313) );
  XOR U17297 ( .A(n17315), .B(n17316), .Z(n17304) );
  AND U17298 ( .A(n17317), .B(n17318), .Z(n17316) );
  XNOR U17299 ( .A(n17315), .B(n17257), .Z(n17318) );
  XNOR U17300 ( .A(n17319), .B(n17320), .Z(n17257) );
  AND U17301 ( .A(n651), .B(n17321), .Z(n17320) );
  XOR U17302 ( .A(n17322), .B(n17319), .Z(n17321) );
  XNOR U17303 ( .A(n17323), .B(n17315), .Z(n17317) );
  IV U17304 ( .A(n17160), .Z(n17323) );
  XOR U17305 ( .A(n17324), .B(n17325), .Z(n17160) );
  AND U17306 ( .A(n659), .B(n17326), .Z(n17325) );
  AND U17307 ( .A(n17278), .B(n17267), .Z(n17315) );
  XNOR U17308 ( .A(n17327), .B(n17328), .Z(n17267) );
  AND U17309 ( .A(n651), .B(n17329), .Z(n17328) );
  XNOR U17310 ( .A(n17330), .B(n17327), .Z(n17329) );
  XNOR U17311 ( .A(n17331), .B(n17332), .Z(n651) );
  AND U17312 ( .A(n17333), .B(n17334), .Z(n17332) );
  XOR U17313 ( .A(n17288), .B(n17331), .Z(n17334) );
  AND U17314 ( .A(n17335), .B(n17336), .Z(n17288) );
  XOR U17315 ( .A(n17331), .B(n17285), .Z(n17333) );
  XOR U17316 ( .A(n17292), .B(n17337), .Z(n17285) );
  AND U17317 ( .A(n655), .B(n17338), .Z(n17337) );
  XOR U17318 ( .A(n17292), .B(n17289), .Z(n17338) );
  XOR U17319 ( .A(n17339), .B(n17340), .Z(n17331) );
  AND U17320 ( .A(n17341), .B(n17342), .Z(n17340) );
  XNOR U17321 ( .A(n17339), .B(n17335), .Z(n17342) );
  IV U17322 ( .A(n17299), .Z(n17335) );
  XOR U17323 ( .A(n17343), .B(n17344), .Z(n17299) );
  XOR U17324 ( .A(n17345), .B(n17336), .Z(n17344) );
  AND U17325 ( .A(n17311), .B(n17346), .Z(n17336) );
  AND U17326 ( .A(n17347), .B(n17348), .Z(n17345) );
  XOR U17327 ( .A(n17349), .B(n17343), .Z(n17347) );
  XNOR U17328 ( .A(n17296), .B(n17339), .Z(n17341) );
  XNOR U17329 ( .A(n17350), .B(n17351), .Z(n17296) );
  AND U17330 ( .A(n655), .B(n17303), .Z(n17351) );
  XOR U17331 ( .A(n17350), .B(n17301), .Z(n17303) );
  XOR U17332 ( .A(n17352), .B(n17353), .Z(n17339) );
  AND U17333 ( .A(n17354), .B(n17355), .Z(n17353) );
  XNOR U17334 ( .A(n17352), .B(n17311), .Z(n17355) );
  XOR U17335 ( .A(n17356), .B(n17348), .Z(n17311) );
  XNOR U17336 ( .A(n17357), .B(n17343), .Z(n17348) );
  XOR U17337 ( .A(n17358), .B(n17359), .Z(n17343) );
  AND U17338 ( .A(n17360), .B(n17361), .Z(n17359) );
  XOR U17339 ( .A(n17362), .B(n17358), .Z(n17360) );
  XNOR U17340 ( .A(n17363), .B(n17364), .Z(n17357) );
  AND U17341 ( .A(n17365), .B(n17366), .Z(n17364) );
  XOR U17342 ( .A(n17363), .B(n17367), .Z(n17365) );
  XNOR U17343 ( .A(n17349), .B(n17346), .Z(n17356) );
  AND U17344 ( .A(n17368), .B(n17369), .Z(n17346) );
  XOR U17345 ( .A(n17370), .B(n17371), .Z(n17349) );
  AND U17346 ( .A(n17372), .B(n17373), .Z(n17371) );
  XOR U17347 ( .A(n17370), .B(n17374), .Z(n17372) );
  XNOR U17348 ( .A(n17308), .B(n17352), .Z(n17354) );
  XNOR U17349 ( .A(n17375), .B(n17376), .Z(n17308) );
  AND U17350 ( .A(n655), .B(n17314), .Z(n17376) );
  XOR U17351 ( .A(n17375), .B(n17312), .Z(n17314) );
  XOR U17352 ( .A(n17377), .B(n17378), .Z(n17352) );
  AND U17353 ( .A(n17379), .B(n17380), .Z(n17378) );
  XNOR U17354 ( .A(n17377), .B(n17368), .Z(n17380) );
  IV U17355 ( .A(n17322), .Z(n17368) );
  XNOR U17356 ( .A(n17381), .B(n17361), .Z(n17322) );
  XNOR U17357 ( .A(n17382), .B(n17367), .Z(n17361) );
  XOR U17358 ( .A(n17383), .B(n17384), .Z(n17367) );
  NOR U17359 ( .A(n17385), .B(n17386), .Z(n17384) );
  XNOR U17360 ( .A(n17383), .B(n17387), .Z(n17385) );
  XNOR U17361 ( .A(n17366), .B(n17358), .Z(n17382) );
  XOR U17362 ( .A(n17388), .B(n17389), .Z(n17358) );
  AND U17363 ( .A(n17390), .B(n17391), .Z(n17389) );
  XNOR U17364 ( .A(n17388), .B(n17392), .Z(n17390) );
  XNOR U17365 ( .A(n17393), .B(n17363), .Z(n17366) );
  XOR U17366 ( .A(n17394), .B(n17395), .Z(n17363) );
  AND U17367 ( .A(n17396), .B(n17397), .Z(n17395) );
  XOR U17368 ( .A(n17394), .B(n17398), .Z(n17396) );
  XNOR U17369 ( .A(n17399), .B(n17400), .Z(n17393) );
  NOR U17370 ( .A(n17401), .B(n17402), .Z(n17400) );
  XOR U17371 ( .A(n17399), .B(n17403), .Z(n17401) );
  XNOR U17372 ( .A(n17362), .B(n17369), .Z(n17381) );
  NOR U17373 ( .A(n17330), .B(n17404), .Z(n17369) );
  XOR U17374 ( .A(n17374), .B(n17373), .Z(n17362) );
  XNOR U17375 ( .A(n17405), .B(n17370), .Z(n17373) );
  XOR U17376 ( .A(n17406), .B(n17407), .Z(n17370) );
  AND U17377 ( .A(n17408), .B(n17409), .Z(n17407) );
  XOR U17378 ( .A(n17406), .B(n17410), .Z(n17408) );
  XNOR U17379 ( .A(n17411), .B(n17412), .Z(n17405) );
  NOR U17380 ( .A(n17413), .B(n17414), .Z(n17412) );
  XNOR U17381 ( .A(n17411), .B(n17415), .Z(n17413) );
  XOR U17382 ( .A(n17416), .B(n17417), .Z(n17374) );
  NOR U17383 ( .A(n17418), .B(n17419), .Z(n17417) );
  XNOR U17384 ( .A(n17416), .B(n17420), .Z(n17418) );
  XNOR U17385 ( .A(n17319), .B(n17377), .Z(n17379) );
  XNOR U17386 ( .A(n17421), .B(n17422), .Z(n17319) );
  AND U17387 ( .A(n655), .B(n17326), .Z(n17422) );
  XOR U17388 ( .A(n17421), .B(n17324), .Z(n17326) );
  AND U17389 ( .A(n17327), .B(n17330), .Z(n17377) );
  XOR U17390 ( .A(n17423), .B(n17404), .Z(n17330) );
  XNOR U17391 ( .A(p_input[1024]), .B(p_input[896]), .Z(n17404) );
  XOR U17392 ( .A(n17392), .B(n17391), .Z(n17423) );
  XNOR U17393 ( .A(n17424), .B(n17398), .Z(n17391) );
  XNOR U17394 ( .A(n17387), .B(n17386), .Z(n17398) );
  XOR U17395 ( .A(n17425), .B(n17383), .Z(n17386) );
  XOR U17396 ( .A(p_input[1034]), .B(p_input[906]), .Z(n17383) );
  XNOR U17397 ( .A(p_input[1035]), .B(p_input[907]), .Z(n17425) );
  XOR U17398 ( .A(p_input[1036]), .B(p_input[908]), .Z(n17387) );
  XNOR U17399 ( .A(n17397), .B(n17388), .Z(n17424) );
  XOR U17400 ( .A(p_input[1025]), .B(p_input[897]), .Z(n17388) );
  XOR U17401 ( .A(n17426), .B(n17403), .Z(n17397) );
  XNOR U17402 ( .A(p_input[1039]), .B(p_input[911]), .Z(n17403) );
  XOR U17403 ( .A(n17394), .B(n17402), .Z(n17426) );
  XOR U17404 ( .A(n17427), .B(n17399), .Z(n17402) );
  XOR U17405 ( .A(p_input[1037]), .B(p_input[909]), .Z(n17399) );
  XNOR U17406 ( .A(p_input[1038]), .B(p_input[910]), .Z(n17427) );
  XOR U17407 ( .A(p_input[1033]), .B(p_input[905]), .Z(n17394) );
  XNOR U17408 ( .A(n17410), .B(n17409), .Z(n17392) );
  XNOR U17409 ( .A(n17428), .B(n17415), .Z(n17409) );
  XOR U17410 ( .A(p_input[1032]), .B(p_input[904]), .Z(n17415) );
  XOR U17411 ( .A(n17406), .B(n17414), .Z(n17428) );
  XOR U17412 ( .A(n17429), .B(n17411), .Z(n17414) );
  XOR U17413 ( .A(p_input[1030]), .B(p_input[902]), .Z(n17411) );
  XNOR U17414 ( .A(p_input[1031]), .B(p_input[903]), .Z(n17429) );
  XOR U17415 ( .A(p_input[1026]), .B(p_input[898]), .Z(n17406) );
  XNOR U17416 ( .A(n17420), .B(n17419), .Z(n17410) );
  XOR U17417 ( .A(n17430), .B(n17416), .Z(n17419) );
  XOR U17418 ( .A(p_input[1027]), .B(p_input[899]), .Z(n17416) );
  XNOR U17419 ( .A(p_input[1028]), .B(p_input[900]), .Z(n17430) );
  XOR U17420 ( .A(p_input[1029]), .B(p_input[901]), .Z(n17420) );
  XNOR U17421 ( .A(n17431), .B(n17432), .Z(n17327) );
  AND U17422 ( .A(n655), .B(n17433), .Z(n17432) );
  XNOR U17423 ( .A(n17434), .B(n17435), .Z(n655) );
  AND U17424 ( .A(n17436), .B(n17437), .Z(n17435) );
  XNOR U17425 ( .A(n17434), .B(n17292), .Z(n17437) );
  XOR U17426 ( .A(n17434), .B(n17289), .Z(n17436) );
  XOR U17427 ( .A(n17438), .B(n17439), .Z(n17434) );
  AND U17428 ( .A(n17440), .B(n17441), .Z(n17439) );
  XOR U17429 ( .A(n17438), .B(n17301), .Z(n17440) );
  XOR U17430 ( .A(n17442), .B(n17443), .Z(n17278) );
  AND U17431 ( .A(n659), .B(n17433), .Z(n17443) );
  XNOR U17432 ( .A(n17431), .B(n17442), .Z(n17433) );
  XNOR U17433 ( .A(n17444), .B(n17445), .Z(n659) );
  AND U17434 ( .A(n17446), .B(n17447), .Z(n17445) );
  XNOR U17435 ( .A(n17292), .B(n17444), .Z(n17447) );
  XOR U17436 ( .A(n17448), .B(n17449), .Z(n17292) );
  AND U17437 ( .A(n17450), .B(n662), .Z(n17449) );
  NOR U17438 ( .A(n17451), .B(n17448), .Z(n17450) );
  XOR U17439 ( .A(n17444), .B(n17289), .Z(n17446) );
  IV U17440 ( .A(n17293), .Z(n17289) );
  AND U17441 ( .A(n17452), .B(n17453), .Z(n17293) );
  XOR U17442 ( .A(n17438), .B(n17454), .Z(n17444) );
  AND U17443 ( .A(n17455), .B(n17441), .Z(n17454) );
  XNOR U17444 ( .A(n17350), .B(n17438), .Z(n17441) );
  XNOR U17445 ( .A(n17456), .B(n17457), .Z(n17350) );
  AND U17446 ( .A(n662), .B(n17458), .Z(n17457) );
  XOR U17447 ( .A(n17459), .B(n17456), .Z(n17458) );
  XNOR U17448 ( .A(n17460), .B(n17438), .Z(n17455) );
  IV U17449 ( .A(n17301), .Z(n17460) );
  XOR U17450 ( .A(n17461), .B(n17462), .Z(n17301) );
  AND U17451 ( .A(n670), .B(n17463), .Z(n17462) );
  XOR U17452 ( .A(n17464), .B(n17465), .Z(n17438) );
  AND U17453 ( .A(n17466), .B(n17467), .Z(n17465) );
  XNOR U17454 ( .A(n17375), .B(n17464), .Z(n17467) );
  XNOR U17455 ( .A(n17468), .B(n17469), .Z(n17375) );
  AND U17456 ( .A(n662), .B(n17470), .Z(n17469) );
  XNOR U17457 ( .A(n17471), .B(n17468), .Z(n17470) );
  XOR U17458 ( .A(n17464), .B(n17312), .Z(n17466) );
  XOR U17459 ( .A(n17472), .B(n17473), .Z(n17312) );
  AND U17460 ( .A(n670), .B(n17474), .Z(n17473) );
  XOR U17461 ( .A(n17475), .B(n17476), .Z(n17464) );
  AND U17462 ( .A(n17477), .B(n17478), .Z(n17476) );
  XNOR U17463 ( .A(n17475), .B(n17421), .Z(n17478) );
  XNOR U17464 ( .A(n17479), .B(n17480), .Z(n17421) );
  AND U17465 ( .A(n662), .B(n17481), .Z(n17480) );
  XOR U17466 ( .A(n17482), .B(n17479), .Z(n17481) );
  XNOR U17467 ( .A(n17483), .B(n17475), .Z(n17477) );
  IV U17468 ( .A(n17324), .Z(n17483) );
  XOR U17469 ( .A(n17484), .B(n17485), .Z(n17324) );
  AND U17470 ( .A(n670), .B(n17486), .Z(n17485) );
  AND U17471 ( .A(n17442), .B(n17431), .Z(n17475) );
  XNOR U17472 ( .A(n17487), .B(n17488), .Z(n17431) );
  AND U17473 ( .A(n662), .B(n17489), .Z(n17488) );
  XNOR U17474 ( .A(n17490), .B(n17487), .Z(n17489) );
  XNOR U17475 ( .A(n17491), .B(n17492), .Z(n662) );
  AND U17476 ( .A(n17493), .B(n17494), .Z(n17492) );
  XOR U17477 ( .A(n17451), .B(n17491), .Z(n17494) );
  AND U17478 ( .A(n17495), .B(n17496), .Z(n17451) );
  XOR U17479 ( .A(n17448), .B(n17491), .Z(n17493) );
  NOR U17480 ( .A(n17452), .B(n17453), .Z(n17448) );
  XOR U17481 ( .A(n17497), .B(n17498), .Z(n17491) );
  AND U17482 ( .A(n17499), .B(n17500), .Z(n17498) );
  XNOR U17483 ( .A(n17497), .B(n17495), .Z(n17500) );
  IV U17484 ( .A(n17459), .Z(n17495) );
  XOR U17485 ( .A(n17501), .B(n17502), .Z(n17459) );
  XOR U17486 ( .A(n17503), .B(n17496), .Z(n17502) );
  AND U17487 ( .A(n17471), .B(n17504), .Z(n17496) );
  AND U17488 ( .A(n17505), .B(n17506), .Z(n17503) );
  XOR U17489 ( .A(n17507), .B(n17501), .Z(n17505) );
  XNOR U17490 ( .A(n17456), .B(n17497), .Z(n17499) );
  XNOR U17491 ( .A(n17508), .B(n17509), .Z(n17456) );
  AND U17492 ( .A(n666), .B(n17463), .Z(n17509) );
  XOR U17493 ( .A(n17508), .B(n17461), .Z(n17463) );
  XOR U17494 ( .A(n17510), .B(n17511), .Z(n17497) );
  AND U17495 ( .A(n17512), .B(n17513), .Z(n17511) );
  XNOR U17496 ( .A(n17510), .B(n17471), .Z(n17513) );
  XOR U17497 ( .A(n17514), .B(n17506), .Z(n17471) );
  XNOR U17498 ( .A(n17515), .B(n17501), .Z(n17506) );
  XOR U17499 ( .A(n17516), .B(n17517), .Z(n17501) );
  AND U17500 ( .A(n17518), .B(n17519), .Z(n17517) );
  XOR U17501 ( .A(n17520), .B(n17516), .Z(n17518) );
  XNOR U17502 ( .A(n17521), .B(n17522), .Z(n17515) );
  AND U17503 ( .A(n17523), .B(n17524), .Z(n17522) );
  XOR U17504 ( .A(n17521), .B(n17525), .Z(n17523) );
  XNOR U17505 ( .A(n17507), .B(n17504), .Z(n17514) );
  AND U17506 ( .A(n17526), .B(n17527), .Z(n17504) );
  XOR U17507 ( .A(n17528), .B(n17529), .Z(n17507) );
  AND U17508 ( .A(n17530), .B(n17531), .Z(n17529) );
  XOR U17509 ( .A(n17528), .B(n17532), .Z(n17530) );
  XNOR U17510 ( .A(n17468), .B(n17510), .Z(n17512) );
  XNOR U17511 ( .A(n17533), .B(n17534), .Z(n17468) );
  AND U17512 ( .A(n666), .B(n17474), .Z(n17534) );
  XOR U17513 ( .A(n17533), .B(n17472), .Z(n17474) );
  XOR U17514 ( .A(n17535), .B(n17536), .Z(n17510) );
  AND U17515 ( .A(n17537), .B(n17538), .Z(n17536) );
  XNOR U17516 ( .A(n17535), .B(n17526), .Z(n17538) );
  IV U17517 ( .A(n17482), .Z(n17526) );
  XNOR U17518 ( .A(n17539), .B(n17519), .Z(n17482) );
  XNOR U17519 ( .A(n17540), .B(n17525), .Z(n17519) );
  XOR U17520 ( .A(n17541), .B(n17542), .Z(n17525) );
  NOR U17521 ( .A(n17543), .B(n17544), .Z(n17542) );
  XNOR U17522 ( .A(n17541), .B(n17545), .Z(n17543) );
  XNOR U17523 ( .A(n17524), .B(n17516), .Z(n17540) );
  XOR U17524 ( .A(n17546), .B(n17547), .Z(n17516) );
  AND U17525 ( .A(n17548), .B(n17549), .Z(n17547) );
  XNOR U17526 ( .A(n17546), .B(n17550), .Z(n17548) );
  XNOR U17527 ( .A(n17551), .B(n17521), .Z(n17524) );
  XOR U17528 ( .A(n17552), .B(n17553), .Z(n17521) );
  AND U17529 ( .A(n17554), .B(n17555), .Z(n17553) );
  XOR U17530 ( .A(n17552), .B(n17556), .Z(n17554) );
  XNOR U17531 ( .A(n17557), .B(n17558), .Z(n17551) );
  NOR U17532 ( .A(n17559), .B(n17560), .Z(n17558) );
  XOR U17533 ( .A(n17557), .B(n17561), .Z(n17559) );
  XNOR U17534 ( .A(n17520), .B(n17527), .Z(n17539) );
  NOR U17535 ( .A(n17490), .B(n17562), .Z(n17527) );
  XOR U17536 ( .A(n17532), .B(n17531), .Z(n17520) );
  XNOR U17537 ( .A(n17563), .B(n17528), .Z(n17531) );
  XOR U17538 ( .A(n17564), .B(n17565), .Z(n17528) );
  AND U17539 ( .A(n17566), .B(n17567), .Z(n17565) );
  XOR U17540 ( .A(n17564), .B(n17568), .Z(n17566) );
  XNOR U17541 ( .A(n17569), .B(n17570), .Z(n17563) );
  NOR U17542 ( .A(n17571), .B(n17572), .Z(n17570) );
  XNOR U17543 ( .A(n17569), .B(n17573), .Z(n17571) );
  XOR U17544 ( .A(n17574), .B(n17575), .Z(n17532) );
  NOR U17545 ( .A(n17576), .B(n17577), .Z(n17575) );
  XNOR U17546 ( .A(n17574), .B(n17578), .Z(n17576) );
  XNOR U17547 ( .A(n17479), .B(n17535), .Z(n17537) );
  XNOR U17548 ( .A(n17579), .B(n17580), .Z(n17479) );
  AND U17549 ( .A(n666), .B(n17486), .Z(n17580) );
  XOR U17550 ( .A(n17579), .B(n17484), .Z(n17486) );
  AND U17551 ( .A(n17487), .B(n17490), .Z(n17535) );
  XOR U17552 ( .A(n17581), .B(n17562), .Z(n17490) );
  XNOR U17553 ( .A(p_input[1024]), .B(p_input[912]), .Z(n17562) );
  XOR U17554 ( .A(n17550), .B(n17549), .Z(n17581) );
  XNOR U17555 ( .A(n17582), .B(n17556), .Z(n17549) );
  XNOR U17556 ( .A(n17545), .B(n17544), .Z(n17556) );
  XOR U17557 ( .A(n17583), .B(n17541), .Z(n17544) );
  XOR U17558 ( .A(p_input[1034]), .B(p_input[922]), .Z(n17541) );
  XNOR U17559 ( .A(p_input[1035]), .B(p_input[923]), .Z(n17583) );
  XOR U17560 ( .A(p_input[1036]), .B(p_input[924]), .Z(n17545) );
  XNOR U17561 ( .A(n17555), .B(n17546), .Z(n17582) );
  XOR U17562 ( .A(p_input[1025]), .B(p_input[913]), .Z(n17546) );
  XOR U17563 ( .A(n17584), .B(n17561), .Z(n17555) );
  XNOR U17564 ( .A(p_input[1039]), .B(p_input[927]), .Z(n17561) );
  XOR U17565 ( .A(n17552), .B(n17560), .Z(n17584) );
  XOR U17566 ( .A(n17585), .B(n17557), .Z(n17560) );
  XOR U17567 ( .A(p_input[1037]), .B(p_input[925]), .Z(n17557) );
  XNOR U17568 ( .A(p_input[1038]), .B(p_input[926]), .Z(n17585) );
  XOR U17569 ( .A(p_input[1033]), .B(p_input[921]), .Z(n17552) );
  XNOR U17570 ( .A(n17568), .B(n17567), .Z(n17550) );
  XNOR U17571 ( .A(n17586), .B(n17573), .Z(n17567) );
  XOR U17572 ( .A(p_input[1032]), .B(p_input[920]), .Z(n17573) );
  XOR U17573 ( .A(n17564), .B(n17572), .Z(n17586) );
  XOR U17574 ( .A(n17587), .B(n17569), .Z(n17572) );
  XOR U17575 ( .A(p_input[1030]), .B(p_input[918]), .Z(n17569) );
  XNOR U17576 ( .A(p_input[1031]), .B(p_input[919]), .Z(n17587) );
  XOR U17577 ( .A(p_input[1026]), .B(p_input[914]), .Z(n17564) );
  XNOR U17578 ( .A(n17578), .B(n17577), .Z(n17568) );
  XOR U17579 ( .A(n17588), .B(n17574), .Z(n17577) );
  XOR U17580 ( .A(p_input[1027]), .B(p_input[915]), .Z(n17574) );
  XNOR U17581 ( .A(p_input[1028]), .B(p_input[916]), .Z(n17588) );
  XOR U17582 ( .A(p_input[1029]), .B(p_input[917]), .Z(n17578) );
  XNOR U17583 ( .A(n17589), .B(n17590), .Z(n17487) );
  AND U17584 ( .A(n666), .B(n17591), .Z(n17590) );
  XNOR U17585 ( .A(n17592), .B(n17593), .Z(n666) );
  NOR U17586 ( .A(n17594), .B(n17595), .Z(n17593) );
  XOR U17587 ( .A(n17453), .B(n17592), .Z(n17595) );
  NOR U17588 ( .A(n17592), .B(n17452), .Z(n17594) );
  XOR U17589 ( .A(n17596), .B(n17597), .Z(n17592) );
  AND U17590 ( .A(n17598), .B(n17599), .Z(n17597) );
  XOR U17591 ( .A(n17596), .B(n17461), .Z(n17598) );
  XOR U17592 ( .A(n17600), .B(n17601), .Z(n17442) );
  AND U17593 ( .A(n670), .B(n17591), .Z(n17601) );
  XNOR U17594 ( .A(n17589), .B(n17600), .Z(n17591) );
  XNOR U17595 ( .A(n17602), .B(n17603), .Z(n670) );
  NOR U17596 ( .A(n17604), .B(n17605), .Z(n17603) );
  XNOR U17597 ( .A(n17453), .B(n17606), .Z(n17605) );
  IV U17598 ( .A(n17602), .Z(n17606) );
  AND U17599 ( .A(n17607), .B(n17608), .Z(n17453) );
  NOR U17600 ( .A(n17602), .B(n17452), .Z(n17604) );
  AND U17601 ( .A(n17609), .B(n17610), .Z(n17452) );
  IV U17602 ( .A(n17611), .Z(n17609) );
  XOR U17603 ( .A(n17596), .B(n17612), .Z(n17602) );
  AND U17604 ( .A(n17613), .B(n17599), .Z(n17612) );
  XNOR U17605 ( .A(n17508), .B(n17596), .Z(n17599) );
  XNOR U17606 ( .A(n17614), .B(n17615), .Z(n17508) );
  AND U17607 ( .A(n673), .B(n17616), .Z(n17615) );
  XOR U17608 ( .A(n17617), .B(n17614), .Z(n17616) );
  XNOR U17609 ( .A(n17618), .B(n17596), .Z(n17613) );
  IV U17610 ( .A(n17461), .Z(n17618) );
  XOR U17611 ( .A(n17619), .B(n17620), .Z(n17461) );
  AND U17612 ( .A(n681), .B(n17621), .Z(n17620) );
  XOR U17613 ( .A(n17622), .B(n17623), .Z(n17596) );
  AND U17614 ( .A(n17624), .B(n17625), .Z(n17623) );
  XNOR U17615 ( .A(n17533), .B(n17622), .Z(n17625) );
  XNOR U17616 ( .A(n17626), .B(n17627), .Z(n17533) );
  AND U17617 ( .A(n673), .B(n17628), .Z(n17627) );
  XNOR U17618 ( .A(n17629), .B(n17626), .Z(n17628) );
  XOR U17619 ( .A(n17622), .B(n17472), .Z(n17624) );
  XOR U17620 ( .A(n17630), .B(n17631), .Z(n17472) );
  AND U17621 ( .A(n681), .B(n17632), .Z(n17631) );
  XOR U17622 ( .A(n17633), .B(n17634), .Z(n17622) );
  AND U17623 ( .A(n17635), .B(n17636), .Z(n17634) );
  XNOR U17624 ( .A(n17633), .B(n17579), .Z(n17636) );
  XNOR U17625 ( .A(n17637), .B(n17638), .Z(n17579) );
  AND U17626 ( .A(n673), .B(n17639), .Z(n17638) );
  XOR U17627 ( .A(n17640), .B(n17637), .Z(n17639) );
  XNOR U17628 ( .A(n17641), .B(n17633), .Z(n17635) );
  IV U17629 ( .A(n17484), .Z(n17641) );
  XOR U17630 ( .A(n17642), .B(n17643), .Z(n17484) );
  AND U17631 ( .A(n681), .B(n17644), .Z(n17643) );
  AND U17632 ( .A(n17600), .B(n17589), .Z(n17633) );
  XNOR U17633 ( .A(n17645), .B(n17646), .Z(n17589) );
  AND U17634 ( .A(n673), .B(n17647), .Z(n17646) );
  XNOR U17635 ( .A(n17648), .B(n17645), .Z(n17647) );
  XNOR U17636 ( .A(n17649), .B(n17650), .Z(n673) );
  NOR U17637 ( .A(n17651), .B(n17652), .Z(n17650) );
  XNOR U17638 ( .A(n17649), .B(n17611), .Z(n17652) );
  NOR U17639 ( .A(n17607), .B(n17608), .Z(n17611) );
  NOR U17640 ( .A(n17649), .B(n17610), .Z(n17651) );
  AND U17641 ( .A(n17653), .B(n17654), .Z(n17610) );
  XOR U17642 ( .A(n17655), .B(n17656), .Z(n17649) );
  AND U17643 ( .A(n17657), .B(n17658), .Z(n17656) );
  XNOR U17644 ( .A(n17655), .B(n17653), .Z(n17658) );
  IV U17645 ( .A(n17617), .Z(n17653) );
  XOR U17646 ( .A(n17659), .B(n17660), .Z(n17617) );
  XOR U17647 ( .A(n17661), .B(n17654), .Z(n17660) );
  AND U17648 ( .A(n17629), .B(n17662), .Z(n17654) );
  AND U17649 ( .A(n17663), .B(n17664), .Z(n17661) );
  XOR U17650 ( .A(n17665), .B(n17659), .Z(n17663) );
  XNOR U17651 ( .A(n17614), .B(n17655), .Z(n17657) );
  XNOR U17652 ( .A(n17666), .B(n17667), .Z(n17614) );
  AND U17653 ( .A(n677), .B(n17621), .Z(n17667) );
  XOR U17654 ( .A(n17666), .B(n17619), .Z(n17621) );
  XOR U17655 ( .A(n17668), .B(n17669), .Z(n17655) );
  AND U17656 ( .A(n17670), .B(n17671), .Z(n17669) );
  XNOR U17657 ( .A(n17668), .B(n17629), .Z(n17671) );
  XOR U17658 ( .A(n17672), .B(n17664), .Z(n17629) );
  XNOR U17659 ( .A(n17673), .B(n17659), .Z(n17664) );
  XOR U17660 ( .A(n17674), .B(n17675), .Z(n17659) );
  AND U17661 ( .A(n17676), .B(n17677), .Z(n17675) );
  XOR U17662 ( .A(n17678), .B(n17674), .Z(n17676) );
  XNOR U17663 ( .A(n17679), .B(n17680), .Z(n17673) );
  AND U17664 ( .A(n17681), .B(n17682), .Z(n17680) );
  XOR U17665 ( .A(n17679), .B(n17683), .Z(n17681) );
  XNOR U17666 ( .A(n17665), .B(n17662), .Z(n17672) );
  AND U17667 ( .A(n17684), .B(n17685), .Z(n17662) );
  XOR U17668 ( .A(n17686), .B(n17687), .Z(n17665) );
  AND U17669 ( .A(n17688), .B(n17689), .Z(n17687) );
  XOR U17670 ( .A(n17686), .B(n17690), .Z(n17688) );
  XNOR U17671 ( .A(n17626), .B(n17668), .Z(n17670) );
  XNOR U17672 ( .A(n17691), .B(n17692), .Z(n17626) );
  AND U17673 ( .A(n677), .B(n17632), .Z(n17692) );
  XOR U17674 ( .A(n17691), .B(n17630), .Z(n17632) );
  XOR U17675 ( .A(n17693), .B(n17694), .Z(n17668) );
  AND U17676 ( .A(n17695), .B(n17696), .Z(n17694) );
  XNOR U17677 ( .A(n17693), .B(n17684), .Z(n17696) );
  IV U17678 ( .A(n17640), .Z(n17684) );
  XNOR U17679 ( .A(n17697), .B(n17677), .Z(n17640) );
  XNOR U17680 ( .A(n17698), .B(n17683), .Z(n17677) );
  XOR U17681 ( .A(n17699), .B(n17700), .Z(n17683) );
  NOR U17682 ( .A(n17701), .B(n17702), .Z(n17700) );
  XNOR U17683 ( .A(n17699), .B(n17703), .Z(n17701) );
  XNOR U17684 ( .A(n17682), .B(n17674), .Z(n17698) );
  XOR U17685 ( .A(n17704), .B(n17705), .Z(n17674) );
  AND U17686 ( .A(n17706), .B(n17707), .Z(n17705) );
  XNOR U17687 ( .A(n17704), .B(n17708), .Z(n17706) );
  XNOR U17688 ( .A(n17709), .B(n17679), .Z(n17682) );
  XOR U17689 ( .A(n17710), .B(n17711), .Z(n17679) );
  AND U17690 ( .A(n17712), .B(n17713), .Z(n17711) );
  XOR U17691 ( .A(n17710), .B(n17714), .Z(n17712) );
  XNOR U17692 ( .A(n17715), .B(n17716), .Z(n17709) );
  NOR U17693 ( .A(n17717), .B(n17718), .Z(n17716) );
  XOR U17694 ( .A(n17715), .B(n17719), .Z(n17717) );
  XNOR U17695 ( .A(n17678), .B(n17685), .Z(n17697) );
  NOR U17696 ( .A(n17648), .B(n17720), .Z(n17685) );
  XOR U17697 ( .A(n17690), .B(n17689), .Z(n17678) );
  XNOR U17698 ( .A(n17721), .B(n17686), .Z(n17689) );
  XOR U17699 ( .A(n17722), .B(n17723), .Z(n17686) );
  AND U17700 ( .A(n17724), .B(n17725), .Z(n17723) );
  XOR U17701 ( .A(n17722), .B(n17726), .Z(n17724) );
  XNOR U17702 ( .A(n17727), .B(n17728), .Z(n17721) );
  NOR U17703 ( .A(n17729), .B(n17730), .Z(n17728) );
  XNOR U17704 ( .A(n17727), .B(n17731), .Z(n17729) );
  XOR U17705 ( .A(n17732), .B(n17733), .Z(n17690) );
  NOR U17706 ( .A(n17734), .B(n17735), .Z(n17733) );
  XNOR U17707 ( .A(n17732), .B(n17736), .Z(n17734) );
  XNOR U17708 ( .A(n17637), .B(n17693), .Z(n17695) );
  XNOR U17709 ( .A(n17737), .B(n17738), .Z(n17637) );
  AND U17710 ( .A(n677), .B(n17644), .Z(n17738) );
  XOR U17711 ( .A(n17737), .B(n17642), .Z(n17644) );
  AND U17712 ( .A(n17645), .B(n17648), .Z(n17693) );
  XOR U17713 ( .A(n17739), .B(n17720), .Z(n17648) );
  XNOR U17714 ( .A(p_input[1024]), .B(p_input[928]), .Z(n17720) );
  XOR U17715 ( .A(n17708), .B(n17707), .Z(n17739) );
  XNOR U17716 ( .A(n17740), .B(n17714), .Z(n17707) );
  XNOR U17717 ( .A(n17703), .B(n17702), .Z(n17714) );
  XOR U17718 ( .A(n17741), .B(n17699), .Z(n17702) );
  XOR U17719 ( .A(p_input[1034]), .B(p_input[938]), .Z(n17699) );
  XNOR U17720 ( .A(p_input[1035]), .B(p_input[939]), .Z(n17741) );
  XOR U17721 ( .A(p_input[1036]), .B(p_input[940]), .Z(n17703) );
  XNOR U17722 ( .A(n17713), .B(n17704), .Z(n17740) );
  XOR U17723 ( .A(p_input[1025]), .B(p_input[929]), .Z(n17704) );
  XOR U17724 ( .A(n17742), .B(n17719), .Z(n17713) );
  XNOR U17725 ( .A(p_input[1039]), .B(p_input[943]), .Z(n17719) );
  XOR U17726 ( .A(n17710), .B(n17718), .Z(n17742) );
  XOR U17727 ( .A(n17743), .B(n17715), .Z(n17718) );
  XOR U17728 ( .A(p_input[1037]), .B(p_input[941]), .Z(n17715) );
  XNOR U17729 ( .A(p_input[1038]), .B(p_input[942]), .Z(n17743) );
  XOR U17730 ( .A(p_input[1033]), .B(p_input[937]), .Z(n17710) );
  XNOR U17731 ( .A(n17726), .B(n17725), .Z(n17708) );
  XNOR U17732 ( .A(n17744), .B(n17731), .Z(n17725) );
  XOR U17733 ( .A(p_input[1032]), .B(p_input[936]), .Z(n17731) );
  XOR U17734 ( .A(n17722), .B(n17730), .Z(n17744) );
  XOR U17735 ( .A(n17745), .B(n17727), .Z(n17730) );
  XOR U17736 ( .A(p_input[1030]), .B(p_input[934]), .Z(n17727) );
  XNOR U17737 ( .A(p_input[1031]), .B(p_input[935]), .Z(n17745) );
  XOR U17738 ( .A(p_input[1026]), .B(p_input[930]), .Z(n17722) );
  XNOR U17739 ( .A(n17736), .B(n17735), .Z(n17726) );
  XOR U17740 ( .A(n17746), .B(n17732), .Z(n17735) );
  XOR U17741 ( .A(p_input[1027]), .B(p_input[931]), .Z(n17732) );
  XNOR U17742 ( .A(p_input[1028]), .B(p_input[932]), .Z(n17746) );
  XOR U17743 ( .A(p_input[1029]), .B(p_input[933]), .Z(n17736) );
  XNOR U17744 ( .A(n17747), .B(n17748), .Z(n17645) );
  AND U17745 ( .A(n677), .B(n17749), .Z(n17748) );
  XNOR U17746 ( .A(n17750), .B(n17751), .Z(n677) );
  NOR U17747 ( .A(n17752), .B(n17753), .Z(n17751) );
  XOR U17748 ( .A(n17608), .B(n17750), .Z(n17753) );
  NOR U17749 ( .A(n17750), .B(n17607), .Z(n17752) );
  XOR U17750 ( .A(n17754), .B(n17755), .Z(n17750) );
  AND U17751 ( .A(n17756), .B(n17757), .Z(n17755) );
  XOR U17752 ( .A(n17754), .B(n17619), .Z(n17756) );
  XOR U17753 ( .A(n17758), .B(n17759), .Z(n17600) );
  AND U17754 ( .A(n681), .B(n17749), .Z(n17759) );
  XNOR U17755 ( .A(n17747), .B(n17758), .Z(n17749) );
  XNOR U17756 ( .A(n17760), .B(n17761), .Z(n681) );
  NOR U17757 ( .A(n17762), .B(n17763), .Z(n17761) );
  XNOR U17758 ( .A(n17608), .B(n17764), .Z(n17763) );
  IV U17759 ( .A(n17760), .Z(n17764) );
  AND U17760 ( .A(n17765), .B(n17766), .Z(n17608) );
  NOR U17761 ( .A(n17760), .B(n17607), .Z(n17762) );
  AND U17762 ( .A(n17767), .B(n17768), .Z(n17607) );
  IV U17763 ( .A(n17769), .Z(n17767) );
  XOR U17764 ( .A(n17754), .B(n17770), .Z(n17760) );
  AND U17765 ( .A(n17771), .B(n17757), .Z(n17770) );
  XNOR U17766 ( .A(n17666), .B(n17754), .Z(n17757) );
  XNOR U17767 ( .A(n17772), .B(n17773), .Z(n17666) );
  AND U17768 ( .A(n684), .B(n17774), .Z(n17773) );
  XOR U17769 ( .A(n17775), .B(n17772), .Z(n17774) );
  XNOR U17770 ( .A(n17776), .B(n17754), .Z(n17771) );
  IV U17771 ( .A(n17619), .Z(n17776) );
  XOR U17772 ( .A(n17777), .B(n17778), .Z(n17619) );
  AND U17773 ( .A(n692), .B(n17779), .Z(n17778) );
  XOR U17774 ( .A(n17780), .B(n17781), .Z(n17754) );
  AND U17775 ( .A(n17782), .B(n17783), .Z(n17781) );
  XNOR U17776 ( .A(n17691), .B(n17780), .Z(n17783) );
  XNOR U17777 ( .A(n17784), .B(n17785), .Z(n17691) );
  AND U17778 ( .A(n684), .B(n17786), .Z(n17785) );
  XNOR U17779 ( .A(n17787), .B(n17784), .Z(n17786) );
  XOR U17780 ( .A(n17780), .B(n17630), .Z(n17782) );
  XOR U17781 ( .A(n17788), .B(n17789), .Z(n17630) );
  AND U17782 ( .A(n692), .B(n17790), .Z(n17789) );
  XOR U17783 ( .A(n17791), .B(n17792), .Z(n17780) );
  AND U17784 ( .A(n17793), .B(n17794), .Z(n17792) );
  XNOR U17785 ( .A(n17791), .B(n17737), .Z(n17794) );
  XNOR U17786 ( .A(n17795), .B(n17796), .Z(n17737) );
  AND U17787 ( .A(n684), .B(n17797), .Z(n17796) );
  XOR U17788 ( .A(n17798), .B(n17795), .Z(n17797) );
  XNOR U17789 ( .A(n17799), .B(n17791), .Z(n17793) );
  IV U17790 ( .A(n17642), .Z(n17799) );
  XOR U17791 ( .A(n17800), .B(n17801), .Z(n17642) );
  AND U17792 ( .A(n692), .B(n17802), .Z(n17801) );
  AND U17793 ( .A(n17758), .B(n17747), .Z(n17791) );
  XNOR U17794 ( .A(n17803), .B(n17804), .Z(n17747) );
  AND U17795 ( .A(n684), .B(n17805), .Z(n17804) );
  XNOR U17796 ( .A(n17806), .B(n17803), .Z(n17805) );
  XNOR U17797 ( .A(n17807), .B(n17808), .Z(n684) );
  NOR U17798 ( .A(n17809), .B(n17810), .Z(n17808) );
  XNOR U17799 ( .A(n17807), .B(n17769), .Z(n17810) );
  NOR U17800 ( .A(n17765), .B(n17766), .Z(n17769) );
  NOR U17801 ( .A(n17807), .B(n17768), .Z(n17809) );
  AND U17802 ( .A(n17811), .B(n17812), .Z(n17768) );
  XOR U17803 ( .A(n17813), .B(n17814), .Z(n17807) );
  AND U17804 ( .A(n17815), .B(n17816), .Z(n17814) );
  XNOR U17805 ( .A(n17813), .B(n17811), .Z(n17816) );
  IV U17806 ( .A(n17775), .Z(n17811) );
  XOR U17807 ( .A(n17817), .B(n17818), .Z(n17775) );
  XOR U17808 ( .A(n17819), .B(n17812), .Z(n17818) );
  AND U17809 ( .A(n17787), .B(n17820), .Z(n17812) );
  AND U17810 ( .A(n17821), .B(n17822), .Z(n17819) );
  XOR U17811 ( .A(n17823), .B(n17817), .Z(n17821) );
  XNOR U17812 ( .A(n17772), .B(n17813), .Z(n17815) );
  XNOR U17813 ( .A(n17824), .B(n17825), .Z(n17772) );
  AND U17814 ( .A(n688), .B(n17779), .Z(n17825) );
  XOR U17815 ( .A(n17824), .B(n17777), .Z(n17779) );
  XOR U17816 ( .A(n17826), .B(n17827), .Z(n17813) );
  AND U17817 ( .A(n17828), .B(n17829), .Z(n17827) );
  XNOR U17818 ( .A(n17826), .B(n17787), .Z(n17829) );
  XOR U17819 ( .A(n17830), .B(n17822), .Z(n17787) );
  XNOR U17820 ( .A(n17831), .B(n17817), .Z(n17822) );
  XOR U17821 ( .A(n17832), .B(n17833), .Z(n17817) );
  AND U17822 ( .A(n17834), .B(n17835), .Z(n17833) );
  XOR U17823 ( .A(n17836), .B(n17832), .Z(n17834) );
  XNOR U17824 ( .A(n17837), .B(n17838), .Z(n17831) );
  AND U17825 ( .A(n17839), .B(n17840), .Z(n17838) );
  XOR U17826 ( .A(n17837), .B(n17841), .Z(n17839) );
  XNOR U17827 ( .A(n17823), .B(n17820), .Z(n17830) );
  AND U17828 ( .A(n17842), .B(n17843), .Z(n17820) );
  XOR U17829 ( .A(n17844), .B(n17845), .Z(n17823) );
  AND U17830 ( .A(n17846), .B(n17847), .Z(n17845) );
  XOR U17831 ( .A(n17844), .B(n17848), .Z(n17846) );
  XNOR U17832 ( .A(n17784), .B(n17826), .Z(n17828) );
  XNOR U17833 ( .A(n17849), .B(n17850), .Z(n17784) );
  AND U17834 ( .A(n688), .B(n17790), .Z(n17850) );
  XOR U17835 ( .A(n17849), .B(n17788), .Z(n17790) );
  XOR U17836 ( .A(n17851), .B(n17852), .Z(n17826) );
  AND U17837 ( .A(n17853), .B(n17854), .Z(n17852) );
  XNOR U17838 ( .A(n17851), .B(n17842), .Z(n17854) );
  IV U17839 ( .A(n17798), .Z(n17842) );
  XNOR U17840 ( .A(n17855), .B(n17835), .Z(n17798) );
  XNOR U17841 ( .A(n17856), .B(n17841), .Z(n17835) );
  XOR U17842 ( .A(n17857), .B(n17858), .Z(n17841) );
  NOR U17843 ( .A(n17859), .B(n17860), .Z(n17858) );
  XNOR U17844 ( .A(n17857), .B(n17861), .Z(n17859) );
  XNOR U17845 ( .A(n17840), .B(n17832), .Z(n17856) );
  XOR U17846 ( .A(n17862), .B(n17863), .Z(n17832) );
  AND U17847 ( .A(n17864), .B(n17865), .Z(n17863) );
  XNOR U17848 ( .A(n17862), .B(n17866), .Z(n17864) );
  XNOR U17849 ( .A(n17867), .B(n17837), .Z(n17840) );
  XOR U17850 ( .A(n17868), .B(n17869), .Z(n17837) );
  AND U17851 ( .A(n17870), .B(n17871), .Z(n17869) );
  XOR U17852 ( .A(n17868), .B(n17872), .Z(n17870) );
  XNOR U17853 ( .A(n17873), .B(n17874), .Z(n17867) );
  NOR U17854 ( .A(n17875), .B(n17876), .Z(n17874) );
  XOR U17855 ( .A(n17873), .B(n17877), .Z(n17875) );
  XNOR U17856 ( .A(n17836), .B(n17843), .Z(n17855) );
  NOR U17857 ( .A(n17806), .B(n17878), .Z(n17843) );
  XOR U17858 ( .A(n17848), .B(n17847), .Z(n17836) );
  XNOR U17859 ( .A(n17879), .B(n17844), .Z(n17847) );
  XOR U17860 ( .A(n17880), .B(n17881), .Z(n17844) );
  AND U17861 ( .A(n17882), .B(n17883), .Z(n17881) );
  XOR U17862 ( .A(n17880), .B(n17884), .Z(n17882) );
  XNOR U17863 ( .A(n17885), .B(n17886), .Z(n17879) );
  NOR U17864 ( .A(n17887), .B(n17888), .Z(n17886) );
  XNOR U17865 ( .A(n17885), .B(n17889), .Z(n17887) );
  XOR U17866 ( .A(n17890), .B(n17891), .Z(n17848) );
  NOR U17867 ( .A(n17892), .B(n17893), .Z(n17891) );
  XNOR U17868 ( .A(n17890), .B(n17894), .Z(n17892) );
  XNOR U17869 ( .A(n17795), .B(n17851), .Z(n17853) );
  XNOR U17870 ( .A(n17895), .B(n17896), .Z(n17795) );
  AND U17871 ( .A(n688), .B(n17802), .Z(n17896) );
  XOR U17872 ( .A(n17895), .B(n17800), .Z(n17802) );
  AND U17873 ( .A(n17803), .B(n17806), .Z(n17851) );
  XOR U17874 ( .A(n17897), .B(n17878), .Z(n17806) );
  XNOR U17875 ( .A(p_input[1024]), .B(p_input[944]), .Z(n17878) );
  XOR U17876 ( .A(n17866), .B(n17865), .Z(n17897) );
  XNOR U17877 ( .A(n17898), .B(n17872), .Z(n17865) );
  XNOR U17878 ( .A(n17861), .B(n17860), .Z(n17872) );
  XOR U17879 ( .A(n17899), .B(n17857), .Z(n17860) );
  XOR U17880 ( .A(p_input[1034]), .B(p_input[954]), .Z(n17857) );
  XNOR U17881 ( .A(p_input[1035]), .B(p_input[955]), .Z(n17899) );
  XOR U17882 ( .A(p_input[1036]), .B(p_input[956]), .Z(n17861) );
  XNOR U17883 ( .A(n17871), .B(n17862), .Z(n17898) );
  XOR U17884 ( .A(p_input[1025]), .B(p_input[945]), .Z(n17862) );
  XOR U17885 ( .A(n17900), .B(n17877), .Z(n17871) );
  XNOR U17886 ( .A(p_input[1039]), .B(p_input[959]), .Z(n17877) );
  XOR U17887 ( .A(n17868), .B(n17876), .Z(n17900) );
  XOR U17888 ( .A(n17901), .B(n17873), .Z(n17876) );
  XOR U17889 ( .A(p_input[1037]), .B(p_input[957]), .Z(n17873) );
  XNOR U17890 ( .A(p_input[1038]), .B(p_input[958]), .Z(n17901) );
  XOR U17891 ( .A(p_input[1033]), .B(p_input[953]), .Z(n17868) );
  XNOR U17892 ( .A(n17884), .B(n17883), .Z(n17866) );
  XNOR U17893 ( .A(n17902), .B(n17889), .Z(n17883) );
  XOR U17894 ( .A(p_input[1032]), .B(p_input[952]), .Z(n17889) );
  XOR U17895 ( .A(n17880), .B(n17888), .Z(n17902) );
  XOR U17896 ( .A(n17903), .B(n17885), .Z(n17888) );
  XOR U17897 ( .A(p_input[1030]), .B(p_input[950]), .Z(n17885) );
  XNOR U17898 ( .A(p_input[1031]), .B(p_input[951]), .Z(n17903) );
  XOR U17899 ( .A(p_input[1026]), .B(p_input[946]), .Z(n17880) );
  XNOR U17900 ( .A(n17894), .B(n17893), .Z(n17884) );
  XOR U17901 ( .A(n17904), .B(n17890), .Z(n17893) );
  XOR U17902 ( .A(p_input[1027]), .B(p_input[947]), .Z(n17890) );
  XNOR U17903 ( .A(p_input[1028]), .B(p_input[948]), .Z(n17904) );
  XOR U17904 ( .A(p_input[1029]), .B(p_input[949]), .Z(n17894) );
  XNOR U17905 ( .A(n17905), .B(n17906), .Z(n17803) );
  AND U17906 ( .A(n688), .B(n17907), .Z(n17906) );
  XNOR U17907 ( .A(n17908), .B(n17909), .Z(n688) );
  NOR U17908 ( .A(n17910), .B(n17911), .Z(n17909) );
  XOR U17909 ( .A(n17766), .B(n17908), .Z(n17911) );
  NOR U17910 ( .A(n17908), .B(n17765), .Z(n17910) );
  XOR U17911 ( .A(n17912), .B(n17913), .Z(n17908) );
  AND U17912 ( .A(n17914), .B(n17915), .Z(n17913) );
  XOR U17913 ( .A(n17912), .B(n17777), .Z(n17914) );
  XOR U17914 ( .A(n17916), .B(n17917), .Z(n17758) );
  AND U17915 ( .A(n692), .B(n17907), .Z(n17917) );
  XNOR U17916 ( .A(n17905), .B(n17916), .Z(n17907) );
  XNOR U17917 ( .A(n17918), .B(n17919), .Z(n692) );
  NOR U17918 ( .A(n17920), .B(n17921), .Z(n17919) );
  XNOR U17919 ( .A(n17766), .B(n17922), .Z(n17921) );
  IV U17920 ( .A(n17918), .Z(n17922) );
  AND U17921 ( .A(n17923), .B(n17924), .Z(n17766) );
  NOR U17922 ( .A(n17918), .B(n17765), .Z(n17920) );
  AND U17923 ( .A(n17925), .B(n17926), .Z(n17765) );
  IV U17924 ( .A(n17927), .Z(n17925) );
  XOR U17925 ( .A(n17912), .B(n17928), .Z(n17918) );
  AND U17926 ( .A(n17929), .B(n17915), .Z(n17928) );
  XNOR U17927 ( .A(n17824), .B(n17912), .Z(n17915) );
  XNOR U17928 ( .A(n17930), .B(n17931), .Z(n17824) );
  AND U17929 ( .A(n695), .B(n17932), .Z(n17931) );
  XOR U17930 ( .A(n17933), .B(n17930), .Z(n17932) );
  XNOR U17931 ( .A(n17934), .B(n17912), .Z(n17929) );
  IV U17932 ( .A(n17777), .Z(n17934) );
  XOR U17933 ( .A(n17935), .B(n17936), .Z(n17777) );
  AND U17934 ( .A(n703), .B(n17937), .Z(n17936) );
  XOR U17935 ( .A(n17938), .B(n17939), .Z(n17912) );
  AND U17936 ( .A(n17940), .B(n17941), .Z(n17939) );
  XNOR U17937 ( .A(n17849), .B(n17938), .Z(n17941) );
  XNOR U17938 ( .A(n17942), .B(n17943), .Z(n17849) );
  AND U17939 ( .A(n695), .B(n17944), .Z(n17943) );
  XNOR U17940 ( .A(n17945), .B(n17942), .Z(n17944) );
  XOR U17941 ( .A(n17938), .B(n17788), .Z(n17940) );
  XOR U17942 ( .A(n17946), .B(n17947), .Z(n17788) );
  AND U17943 ( .A(n703), .B(n17948), .Z(n17947) );
  XOR U17944 ( .A(n17949), .B(n17950), .Z(n17938) );
  AND U17945 ( .A(n17951), .B(n17952), .Z(n17950) );
  XNOR U17946 ( .A(n17949), .B(n17895), .Z(n17952) );
  XNOR U17947 ( .A(n17953), .B(n17954), .Z(n17895) );
  AND U17948 ( .A(n695), .B(n17955), .Z(n17954) );
  XOR U17949 ( .A(n17956), .B(n17953), .Z(n17955) );
  XNOR U17950 ( .A(n17957), .B(n17949), .Z(n17951) );
  IV U17951 ( .A(n17800), .Z(n17957) );
  XOR U17952 ( .A(n17958), .B(n17959), .Z(n17800) );
  AND U17953 ( .A(n703), .B(n17960), .Z(n17959) );
  AND U17954 ( .A(n17916), .B(n17905), .Z(n17949) );
  XNOR U17955 ( .A(n17961), .B(n17962), .Z(n17905) );
  AND U17956 ( .A(n695), .B(n17963), .Z(n17962) );
  XNOR U17957 ( .A(n17964), .B(n17961), .Z(n17963) );
  XNOR U17958 ( .A(n17965), .B(n17966), .Z(n695) );
  NOR U17959 ( .A(n17967), .B(n17968), .Z(n17966) );
  XNOR U17960 ( .A(n17965), .B(n17927), .Z(n17968) );
  NOR U17961 ( .A(n17923), .B(n17924), .Z(n17927) );
  NOR U17962 ( .A(n17965), .B(n17926), .Z(n17967) );
  AND U17963 ( .A(n17969), .B(n17970), .Z(n17926) );
  XOR U17964 ( .A(n17971), .B(n17972), .Z(n17965) );
  AND U17965 ( .A(n17973), .B(n17974), .Z(n17972) );
  XNOR U17966 ( .A(n17971), .B(n17969), .Z(n17974) );
  IV U17967 ( .A(n17933), .Z(n17969) );
  XOR U17968 ( .A(n17975), .B(n17976), .Z(n17933) );
  XOR U17969 ( .A(n17977), .B(n17970), .Z(n17976) );
  AND U17970 ( .A(n17945), .B(n17978), .Z(n17970) );
  AND U17971 ( .A(n17979), .B(n17980), .Z(n17977) );
  XOR U17972 ( .A(n17981), .B(n17975), .Z(n17979) );
  XNOR U17973 ( .A(n17930), .B(n17971), .Z(n17973) );
  XNOR U17974 ( .A(n17982), .B(n17983), .Z(n17930) );
  AND U17975 ( .A(n699), .B(n17937), .Z(n17983) );
  XOR U17976 ( .A(n17982), .B(n17935), .Z(n17937) );
  XOR U17977 ( .A(n17984), .B(n17985), .Z(n17971) );
  AND U17978 ( .A(n17986), .B(n17987), .Z(n17985) );
  XNOR U17979 ( .A(n17984), .B(n17945), .Z(n17987) );
  XOR U17980 ( .A(n17988), .B(n17980), .Z(n17945) );
  XNOR U17981 ( .A(n17989), .B(n17975), .Z(n17980) );
  XOR U17982 ( .A(n17990), .B(n17991), .Z(n17975) );
  AND U17983 ( .A(n17992), .B(n17993), .Z(n17991) );
  XOR U17984 ( .A(n17994), .B(n17990), .Z(n17992) );
  XNOR U17985 ( .A(n17995), .B(n17996), .Z(n17989) );
  AND U17986 ( .A(n17997), .B(n17998), .Z(n17996) );
  XOR U17987 ( .A(n17995), .B(n17999), .Z(n17997) );
  XNOR U17988 ( .A(n17981), .B(n17978), .Z(n17988) );
  AND U17989 ( .A(n18000), .B(n18001), .Z(n17978) );
  XOR U17990 ( .A(n18002), .B(n18003), .Z(n17981) );
  AND U17991 ( .A(n18004), .B(n18005), .Z(n18003) );
  XOR U17992 ( .A(n18002), .B(n18006), .Z(n18004) );
  XNOR U17993 ( .A(n17942), .B(n17984), .Z(n17986) );
  XNOR U17994 ( .A(n18007), .B(n18008), .Z(n17942) );
  AND U17995 ( .A(n699), .B(n17948), .Z(n18008) );
  XOR U17996 ( .A(n18007), .B(n17946), .Z(n17948) );
  XOR U17997 ( .A(n18009), .B(n18010), .Z(n17984) );
  AND U17998 ( .A(n18011), .B(n18012), .Z(n18010) );
  XNOR U17999 ( .A(n18009), .B(n18000), .Z(n18012) );
  IV U18000 ( .A(n17956), .Z(n18000) );
  XNOR U18001 ( .A(n18013), .B(n17993), .Z(n17956) );
  XNOR U18002 ( .A(n18014), .B(n17999), .Z(n17993) );
  XOR U18003 ( .A(n18015), .B(n18016), .Z(n17999) );
  NOR U18004 ( .A(n18017), .B(n18018), .Z(n18016) );
  XNOR U18005 ( .A(n18015), .B(n18019), .Z(n18017) );
  XNOR U18006 ( .A(n17998), .B(n17990), .Z(n18014) );
  XOR U18007 ( .A(n18020), .B(n18021), .Z(n17990) );
  AND U18008 ( .A(n18022), .B(n18023), .Z(n18021) );
  XNOR U18009 ( .A(n18020), .B(n18024), .Z(n18022) );
  XNOR U18010 ( .A(n18025), .B(n17995), .Z(n17998) );
  XOR U18011 ( .A(n18026), .B(n18027), .Z(n17995) );
  AND U18012 ( .A(n18028), .B(n18029), .Z(n18027) );
  XOR U18013 ( .A(n18026), .B(n18030), .Z(n18028) );
  XNOR U18014 ( .A(n18031), .B(n18032), .Z(n18025) );
  NOR U18015 ( .A(n18033), .B(n18034), .Z(n18032) );
  XOR U18016 ( .A(n18031), .B(n18035), .Z(n18033) );
  XNOR U18017 ( .A(n17994), .B(n18001), .Z(n18013) );
  NOR U18018 ( .A(n17964), .B(n18036), .Z(n18001) );
  XOR U18019 ( .A(n18006), .B(n18005), .Z(n17994) );
  XNOR U18020 ( .A(n18037), .B(n18002), .Z(n18005) );
  XOR U18021 ( .A(n18038), .B(n18039), .Z(n18002) );
  AND U18022 ( .A(n18040), .B(n18041), .Z(n18039) );
  XOR U18023 ( .A(n18038), .B(n18042), .Z(n18040) );
  XNOR U18024 ( .A(n18043), .B(n18044), .Z(n18037) );
  NOR U18025 ( .A(n18045), .B(n18046), .Z(n18044) );
  XNOR U18026 ( .A(n18043), .B(n18047), .Z(n18045) );
  XOR U18027 ( .A(n18048), .B(n18049), .Z(n18006) );
  NOR U18028 ( .A(n18050), .B(n18051), .Z(n18049) );
  XNOR U18029 ( .A(n18048), .B(n18052), .Z(n18050) );
  XNOR U18030 ( .A(n17953), .B(n18009), .Z(n18011) );
  XNOR U18031 ( .A(n18053), .B(n18054), .Z(n17953) );
  AND U18032 ( .A(n699), .B(n17960), .Z(n18054) );
  XOR U18033 ( .A(n18053), .B(n17958), .Z(n17960) );
  AND U18034 ( .A(n17961), .B(n17964), .Z(n18009) );
  XOR U18035 ( .A(n18055), .B(n18036), .Z(n17964) );
  XNOR U18036 ( .A(p_input[1024]), .B(p_input[960]), .Z(n18036) );
  XOR U18037 ( .A(n18024), .B(n18023), .Z(n18055) );
  XNOR U18038 ( .A(n18056), .B(n18030), .Z(n18023) );
  XNOR U18039 ( .A(n18019), .B(n18018), .Z(n18030) );
  XOR U18040 ( .A(n18057), .B(n18015), .Z(n18018) );
  XOR U18041 ( .A(p_input[1034]), .B(p_input[970]), .Z(n18015) );
  XNOR U18042 ( .A(p_input[1035]), .B(p_input[971]), .Z(n18057) );
  XOR U18043 ( .A(p_input[1036]), .B(p_input[972]), .Z(n18019) );
  XNOR U18044 ( .A(n18029), .B(n18020), .Z(n18056) );
  XOR U18045 ( .A(p_input[1025]), .B(p_input[961]), .Z(n18020) );
  XOR U18046 ( .A(n18058), .B(n18035), .Z(n18029) );
  XNOR U18047 ( .A(p_input[1039]), .B(p_input[975]), .Z(n18035) );
  XOR U18048 ( .A(n18026), .B(n18034), .Z(n18058) );
  XOR U18049 ( .A(n18059), .B(n18031), .Z(n18034) );
  XOR U18050 ( .A(p_input[1037]), .B(p_input[973]), .Z(n18031) );
  XNOR U18051 ( .A(p_input[1038]), .B(p_input[974]), .Z(n18059) );
  XOR U18052 ( .A(p_input[1033]), .B(p_input[969]), .Z(n18026) );
  XNOR U18053 ( .A(n18042), .B(n18041), .Z(n18024) );
  XNOR U18054 ( .A(n18060), .B(n18047), .Z(n18041) );
  XOR U18055 ( .A(p_input[1032]), .B(p_input[968]), .Z(n18047) );
  XOR U18056 ( .A(n18038), .B(n18046), .Z(n18060) );
  XOR U18057 ( .A(n18061), .B(n18043), .Z(n18046) );
  XOR U18058 ( .A(p_input[1030]), .B(p_input[966]), .Z(n18043) );
  XNOR U18059 ( .A(p_input[1031]), .B(p_input[967]), .Z(n18061) );
  XOR U18060 ( .A(p_input[1026]), .B(p_input[962]), .Z(n18038) );
  XNOR U18061 ( .A(n18052), .B(n18051), .Z(n18042) );
  XOR U18062 ( .A(n18062), .B(n18048), .Z(n18051) );
  XOR U18063 ( .A(p_input[1027]), .B(p_input[963]), .Z(n18048) );
  XNOR U18064 ( .A(p_input[1028]), .B(p_input[964]), .Z(n18062) );
  XOR U18065 ( .A(p_input[1029]), .B(p_input[965]), .Z(n18052) );
  XNOR U18066 ( .A(n18063), .B(n18064), .Z(n17961) );
  AND U18067 ( .A(n699), .B(n18065), .Z(n18064) );
  XNOR U18068 ( .A(n18066), .B(n18067), .Z(n699) );
  NOR U18069 ( .A(n18068), .B(n18069), .Z(n18067) );
  XOR U18070 ( .A(n17924), .B(n18066), .Z(n18069) );
  NOR U18071 ( .A(n18066), .B(n17923), .Z(n18068) );
  XOR U18072 ( .A(n18070), .B(n18071), .Z(n18066) );
  AND U18073 ( .A(n18072), .B(n18073), .Z(n18071) );
  XOR U18074 ( .A(n18070), .B(n17935), .Z(n18072) );
  XOR U18075 ( .A(n18074), .B(n18075), .Z(n17916) );
  AND U18076 ( .A(n703), .B(n18065), .Z(n18075) );
  XNOR U18077 ( .A(n18063), .B(n18074), .Z(n18065) );
  XNOR U18078 ( .A(n18076), .B(n18077), .Z(n703) );
  NOR U18079 ( .A(n18078), .B(n18079), .Z(n18077) );
  XNOR U18080 ( .A(n17924), .B(n18080), .Z(n18079) );
  IV U18081 ( .A(n18076), .Z(n18080) );
  AND U18082 ( .A(n18081), .B(n18082), .Z(n17924) );
  NOR U18083 ( .A(n18076), .B(n17923), .Z(n18078) );
  AND U18084 ( .A(n18083), .B(n18084), .Z(n17923) );
  IV U18085 ( .A(n18085), .Z(n18083) );
  XOR U18086 ( .A(n18070), .B(n18086), .Z(n18076) );
  AND U18087 ( .A(n18087), .B(n18073), .Z(n18086) );
  XNOR U18088 ( .A(n17982), .B(n18070), .Z(n18073) );
  XNOR U18089 ( .A(n18088), .B(n18089), .Z(n17982) );
  AND U18090 ( .A(n706), .B(n18090), .Z(n18089) );
  XOR U18091 ( .A(n18091), .B(n18088), .Z(n18090) );
  XNOR U18092 ( .A(n18092), .B(n18070), .Z(n18087) );
  IV U18093 ( .A(n17935), .Z(n18092) );
  XOR U18094 ( .A(n18093), .B(n18094), .Z(n17935) );
  AND U18095 ( .A(n713), .B(n18095), .Z(n18094) );
  XOR U18096 ( .A(n18096), .B(n18097), .Z(n18070) );
  AND U18097 ( .A(n18098), .B(n18099), .Z(n18097) );
  XNOR U18098 ( .A(n18007), .B(n18096), .Z(n18099) );
  XNOR U18099 ( .A(n18100), .B(n18101), .Z(n18007) );
  AND U18100 ( .A(n706), .B(n18102), .Z(n18101) );
  XNOR U18101 ( .A(n18103), .B(n18100), .Z(n18102) );
  XOR U18102 ( .A(n18096), .B(n17946), .Z(n18098) );
  XOR U18103 ( .A(n18104), .B(n18105), .Z(n17946) );
  AND U18104 ( .A(n713), .B(n18106), .Z(n18105) );
  XOR U18105 ( .A(n18107), .B(n18108), .Z(n18096) );
  AND U18106 ( .A(n18109), .B(n18110), .Z(n18108) );
  XNOR U18107 ( .A(n18107), .B(n18053), .Z(n18110) );
  XNOR U18108 ( .A(n18111), .B(n18112), .Z(n18053) );
  AND U18109 ( .A(n706), .B(n18113), .Z(n18112) );
  XOR U18110 ( .A(n18114), .B(n18111), .Z(n18113) );
  XNOR U18111 ( .A(n18115), .B(n18107), .Z(n18109) );
  IV U18112 ( .A(n17958), .Z(n18115) );
  XOR U18113 ( .A(n18116), .B(n18117), .Z(n17958) );
  AND U18114 ( .A(n713), .B(n18118), .Z(n18117) );
  AND U18115 ( .A(n18074), .B(n18063), .Z(n18107) );
  XNOR U18116 ( .A(n18119), .B(n18120), .Z(n18063) );
  AND U18117 ( .A(n706), .B(n18121), .Z(n18120) );
  XNOR U18118 ( .A(n18122), .B(n18119), .Z(n18121) );
  XNOR U18119 ( .A(n18123), .B(n18124), .Z(n706) );
  NOR U18120 ( .A(n18125), .B(n18126), .Z(n18124) );
  XNOR U18121 ( .A(n18123), .B(n18085), .Z(n18126) );
  NOR U18122 ( .A(n18081), .B(n18082), .Z(n18085) );
  NOR U18123 ( .A(n18123), .B(n18084), .Z(n18125) );
  AND U18124 ( .A(n18127), .B(n18128), .Z(n18084) );
  XOR U18125 ( .A(n18129), .B(n18130), .Z(n18123) );
  AND U18126 ( .A(n18131), .B(n18132), .Z(n18130) );
  XNOR U18127 ( .A(n18129), .B(n18127), .Z(n18132) );
  IV U18128 ( .A(n18091), .Z(n18127) );
  XOR U18129 ( .A(n18133), .B(n18134), .Z(n18091) );
  XOR U18130 ( .A(n18135), .B(n18128), .Z(n18134) );
  AND U18131 ( .A(n18103), .B(n18136), .Z(n18128) );
  AND U18132 ( .A(n18137), .B(n18138), .Z(n18135) );
  XOR U18133 ( .A(n18139), .B(n18133), .Z(n18137) );
  XNOR U18134 ( .A(n18088), .B(n18129), .Z(n18131) );
  XNOR U18135 ( .A(n18140), .B(n18141), .Z(n18088) );
  AND U18136 ( .A(n710), .B(n18095), .Z(n18141) );
  XOR U18137 ( .A(n18140), .B(n18093), .Z(n18095) );
  XOR U18138 ( .A(n18142), .B(n18143), .Z(n18129) );
  AND U18139 ( .A(n18144), .B(n18145), .Z(n18143) );
  XNOR U18140 ( .A(n18142), .B(n18103), .Z(n18145) );
  XOR U18141 ( .A(n18146), .B(n18138), .Z(n18103) );
  XNOR U18142 ( .A(n18147), .B(n18133), .Z(n18138) );
  XOR U18143 ( .A(n18148), .B(n18149), .Z(n18133) );
  AND U18144 ( .A(n18150), .B(n18151), .Z(n18149) );
  XOR U18145 ( .A(n18152), .B(n18148), .Z(n18150) );
  XNOR U18146 ( .A(n18153), .B(n18154), .Z(n18147) );
  AND U18147 ( .A(n18155), .B(n18156), .Z(n18154) );
  XOR U18148 ( .A(n18153), .B(n18157), .Z(n18155) );
  XNOR U18149 ( .A(n18139), .B(n18136), .Z(n18146) );
  AND U18150 ( .A(n18158), .B(n18159), .Z(n18136) );
  XOR U18151 ( .A(n18160), .B(n18161), .Z(n18139) );
  AND U18152 ( .A(n18162), .B(n18163), .Z(n18161) );
  XOR U18153 ( .A(n18160), .B(n18164), .Z(n18162) );
  XNOR U18154 ( .A(n18100), .B(n18142), .Z(n18144) );
  XNOR U18155 ( .A(n18165), .B(n18166), .Z(n18100) );
  AND U18156 ( .A(n710), .B(n18106), .Z(n18166) );
  XOR U18157 ( .A(n18165), .B(n18104), .Z(n18106) );
  XOR U18158 ( .A(n18167), .B(n18168), .Z(n18142) );
  AND U18159 ( .A(n18169), .B(n18170), .Z(n18168) );
  XNOR U18160 ( .A(n18167), .B(n18158), .Z(n18170) );
  IV U18161 ( .A(n18114), .Z(n18158) );
  XNOR U18162 ( .A(n18171), .B(n18151), .Z(n18114) );
  XNOR U18163 ( .A(n18172), .B(n18157), .Z(n18151) );
  XOR U18164 ( .A(n18173), .B(n18174), .Z(n18157) );
  NOR U18165 ( .A(n18175), .B(n18176), .Z(n18174) );
  XNOR U18166 ( .A(n18173), .B(n18177), .Z(n18175) );
  XNOR U18167 ( .A(n18156), .B(n18148), .Z(n18172) );
  XOR U18168 ( .A(n18178), .B(n18179), .Z(n18148) );
  AND U18169 ( .A(n18180), .B(n18181), .Z(n18179) );
  XNOR U18170 ( .A(n18178), .B(n18182), .Z(n18180) );
  XNOR U18171 ( .A(n18183), .B(n18153), .Z(n18156) );
  XOR U18172 ( .A(n18184), .B(n18185), .Z(n18153) );
  AND U18173 ( .A(n18186), .B(n18187), .Z(n18185) );
  XOR U18174 ( .A(n18184), .B(n18188), .Z(n18186) );
  XNOR U18175 ( .A(n18189), .B(n18190), .Z(n18183) );
  NOR U18176 ( .A(n18191), .B(n18192), .Z(n18190) );
  XOR U18177 ( .A(n18189), .B(n18193), .Z(n18191) );
  XNOR U18178 ( .A(n18152), .B(n18159), .Z(n18171) );
  NOR U18179 ( .A(n18122), .B(n18194), .Z(n18159) );
  XOR U18180 ( .A(n18164), .B(n18163), .Z(n18152) );
  XNOR U18181 ( .A(n18195), .B(n18160), .Z(n18163) );
  XOR U18182 ( .A(n18196), .B(n18197), .Z(n18160) );
  AND U18183 ( .A(n18198), .B(n18199), .Z(n18197) );
  XOR U18184 ( .A(n18196), .B(n18200), .Z(n18198) );
  XNOR U18185 ( .A(n18201), .B(n18202), .Z(n18195) );
  NOR U18186 ( .A(n18203), .B(n18204), .Z(n18202) );
  XNOR U18187 ( .A(n18201), .B(n18205), .Z(n18203) );
  XOR U18188 ( .A(n18206), .B(n18207), .Z(n18164) );
  NOR U18189 ( .A(n18208), .B(n18209), .Z(n18207) );
  XNOR U18190 ( .A(n18206), .B(n18210), .Z(n18208) );
  XNOR U18191 ( .A(n18111), .B(n18167), .Z(n18169) );
  XNOR U18192 ( .A(n18211), .B(n18212), .Z(n18111) );
  AND U18193 ( .A(n710), .B(n18118), .Z(n18212) );
  XOR U18194 ( .A(n18211), .B(n18116), .Z(n18118) );
  AND U18195 ( .A(n18119), .B(n18122), .Z(n18167) );
  XOR U18196 ( .A(n18213), .B(n18194), .Z(n18122) );
  XNOR U18197 ( .A(p_input[1024]), .B(p_input[976]), .Z(n18194) );
  XOR U18198 ( .A(n18182), .B(n18181), .Z(n18213) );
  XNOR U18199 ( .A(n18214), .B(n18188), .Z(n18181) );
  XNOR U18200 ( .A(n18177), .B(n18176), .Z(n18188) );
  XOR U18201 ( .A(n18215), .B(n18173), .Z(n18176) );
  XOR U18202 ( .A(p_input[1034]), .B(p_input[986]), .Z(n18173) );
  XNOR U18203 ( .A(p_input[1035]), .B(p_input[987]), .Z(n18215) );
  XOR U18204 ( .A(p_input[1036]), .B(p_input[988]), .Z(n18177) );
  XNOR U18205 ( .A(n18187), .B(n18178), .Z(n18214) );
  XOR U18206 ( .A(p_input[1025]), .B(p_input[977]), .Z(n18178) );
  XOR U18207 ( .A(n18216), .B(n18193), .Z(n18187) );
  XNOR U18208 ( .A(p_input[1039]), .B(p_input[991]), .Z(n18193) );
  XOR U18209 ( .A(n18184), .B(n18192), .Z(n18216) );
  XOR U18210 ( .A(n18217), .B(n18189), .Z(n18192) );
  XOR U18211 ( .A(p_input[1037]), .B(p_input[989]), .Z(n18189) );
  XNOR U18212 ( .A(p_input[1038]), .B(p_input[990]), .Z(n18217) );
  XOR U18213 ( .A(p_input[1033]), .B(p_input[985]), .Z(n18184) );
  XNOR U18214 ( .A(n18200), .B(n18199), .Z(n18182) );
  XNOR U18215 ( .A(n18218), .B(n18205), .Z(n18199) );
  XOR U18216 ( .A(p_input[1032]), .B(p_input[984]), .Z(n18205) );
  XOR U18217 ( .A(n18196), .B(n18204), .Z(n18218) );
  XOR U18218 ( .A(n18219), .B(n18201), .Z(n18204) );
  XOR U18219 ( .A(p_input[1030]), .B(p_input[982]), .Z(n18201) );
  XNOR U18220 ( .A(p_input[1031]), .B(p_input[983]), .Z(n18219) );
  XOR U18221 ( .A(p_input[1026]), .B(p_input[978]), .Z(n18196) );
  XNOR U18222 ( .A(n18210), .B(n18209), .Z(n18200) );
  XOR U18223 ( .A(n18220), .B(n18206), .Z(n18209) );
  XOR U18224 ( .A(p_input[1027]), .B(p_input[979]), .Z(n18206) );
  XNOR U18225 ( .A(p_input[1028]), .B(p_input[980]), .Z(n18220) );
  XOR U18226 ( .A(p_input[1029]), .B(p_input[981]), .Z(n18210) );
  XNOR U18227 ( .A(n18221), .B(n18222), .Z(n18119) );
  AND U18228 ( .A(n710), .B(n18223), .Z(n18222) );
  XNOR U18229 ( .A(n18224), .B(n18225), .Z(n710) );
  NOR U18230 ( .A(n18226), .B(n18227), .Z(n18225) );
  XOR U18231 ( .A(n18082), .B(n18224), .Z(n18227) );
  NOR U18232 ( .A(n18224), .B(n18081), .Z(n18226) );
  XOR U18233 ( .A(n18228), .B(n18229), .Z(n18224) );
  AND U18234 ( .A(n18230), .B(n18231), .Z(n18229) );
  XOR U18235 ( .A(n18228), .B(n18093), .Z(n18230) );
  XOR U18236 ( .A(n18232), .B(n18233), .Z(n18074) );
  AND U18237 ( .A(n713), .B(n18223), .Z(n18233) );
  XOR U18238 ( .A(n18234), .B(n18232), .Z(n18223) );
  XNOR U18239 ( .A(n18235), .B(n18236), .Z(n713) );
  NOR U18240 ( .A(n18237), .B(n18238), .Z(n18236) );
  XNOR U18241 ( .A(n18082), .B(n18239), .Z(n18238) );
  IV U18242 ( .A(n18235), .Z(n18239) );
  AND U18243 ( .A(n18093), .B(n18240), .Z(n18082) );
  NOR U18244 ( .A(n18235), .B(n18081), .Z(n18237) );
  AND U18245 ( .A(n18140), .B(n18241), .Z(n18081) );
  XOR U18246 ( .A(n18228), .B(n18242), .Z(n18235) );
  AND U18247 ( .A(n18243), .B(n18231), .Z(n18242) );
  XNOR U18248 ( .A(n18140), .B(n18228), .Z(n18231) );
  XNOR U18249 ( .A(n18244), .B(n18245), .Z(n18140) );
  XOR U18250 ( .A(n18246), .B(n18241), .Z(n18245) );
  AND U18251 ( .A(n18165), .B(n18247), .Z(n18241) );
  AND U18252 ( .A(n18248), .B(n18249), .Z(n18246) );
  XOR U18253 ( .A(n18250), .B(n18244), .Z(n18248) );
  XNOR U18254 ( .A(n18251), .B(n18228), .Z(n18243) );
  IV U18255 ( .A(n18093), .Z(n18251) );
  XNOR U18256 ( .A(n18252), .B(n18253), .Z(n18093) );
  XOR U18257 ( .A(n18254), .B(n18240), .Z(n18253) );
  AND U18258 ( .A(n18104), .B(n18255), .Z(n18240) );
  AND U18259 ( .A(n18256), .B(n18257), .Z(n18254) );
  XNOR U18260 ( .A(n18252), .B(n18258), .Z(n18256) );
  XOR U18261 ( .A(n18259), .B(n18260), .Z(n18228) );
  AND U18262 ( .A(n18261), .B(n18262), .Z(n18260) );
  XNOR U18263 ( .A(n18165), .B(n18259), .Z(n18262) );
  XOR U18264 ( .A(n18263), .B(n18249), .Z(n18165) );
  XNOR U18265 ( .A(n18264), .B(n18244), .Z(n18249) );
  XOR U18266 ( .A(n18265), .B(n18266), .Z(n18244) );
  AND U18267 ( .A(n18267), .B(n18268), .Z(n18266) );
  XOR U18268 ( .A(n18269), .B(n18265), .Z(n18267) );
  XNOR U18269 ( .A(n18270), .B(n18271), .Z(n18264) );
  AND U18270 ( .A(n18272), .B(n18273), .Z(n18271) );
  XOR U18271 ( .A(n18270), .B(n18274), .Z(n18272) );
  XNOR U18272 ( .A(n18250), .B(n18247), .Z(n18263) );
  AND U18273 ( .A(n18211), .B(n18275), .Z(n18247) );
  XOR U18274 ( .A(n18276), .B(n18277), .Z(n18250) );
  AND U18275 ( .A(n18278), .B(n18279), .Z(n18277) );
  XOR U18276 ( .A(n18276), .B(n18280), .Z(n18278) );
  XOR U18277 ( .A(n18259), .B(n18104), .Z(n18261) );
  XNOR U18278 ( .A(n18281), .B(n18258), .Z(n18104) );
  XNOR U18279 ( .A(n18282), .B(n18283), .Z(n18258) );
  AND U18280 ( .A(n18284), .B(n18285), .Z(n18283) );
  XOR U18281 ( .A(n18282), .B(n18286), .Z(n18284) );
  XNOR U18282 ( .A(n18257), .B(n18255), .Z(n18281) );
  AND U18283 ( .A(n18116), .B(n18287), .Z(n18255) );
  XNOR U18284 ( .A(n18288), .B(n18252), .Z(n18257) );
  XOR U18285 ( .A(n18289), .B(n18290), .Z(n18252) );
  AND U18286 ( .A(n18291), .B(n18292), .Z(n18290) );
  XOR U18287 ( .A(n18289), .B(n18293), .Z(n18291) );
  XNOR U18288 ( .A(n18294), .B(n18295), .Z(n18288) );
  AND U18289 ( .A(n18296), .B(n18297), .Z(n18295) );
  XNOR U18290 ( .A(n18294), .B(n18298), .Z(n18296) );
  XOR U18291 ( .A(n18299), .B(n18300), .Z(n18259) );
  AND U18292 ( .A(n18301), .B(n18302), .Z(n18300) );
  XNOR U18293 ( .A(n18299), .B(n18211), .Z(n18302) );
  XOR U18294 ( .A(n18303), .B(n18268), .Z(n18211) );
  XNOR U18295 ( .A(n18304), .B(n18274), .Z(n18268) );
  XOR U18296 ( .A(n18305), .B(n18306), .Z(n18274) );
  AND U18297 ( .A(n18307), .B(n18308), .Z(n18306) );
  XOR U18298 ( .A(n18305), .B(n18309), .Z(n18307) );
  XNOR U18299 ( .A(n18273), .B(n18265), .Z(n18304) );
  XOR U18300 ( .A(n18310), .B(n18311), .Z(n18265) );
  AND U18301 ( .A(n18312), .B(n18313), .Z(n18311) );
  XNOR U18302 ( .A(n18310), .B(n18314), .Z(n18312) );
  XNOR U18303 ( .A(n18315), .B(n18270), .Z(n18273) );
  XOR U18304 ( .A(n18316), .B(n18317), .Z(n18270) );
  AND U18305 ( .A(n18318), .B(n18319), .Z(n18317) );
  XNOR U18306 ( .A(n18320), .B(n18321), .Z(n18318) );
  XNOR U18307 ( .A(n18322), .B(n18323), .Z(n18315) );
  AND U18308 ( .A(n18324), .B(n18325), .Z(n18323) );
  XNOR U18309 ( .A(n18322), .B(n18326), .Z(n18324) );
  XNOR U18310 ( .A(n18269), .B(n18275), .Z(n18303) );
  AND U18311 ( .A(n18234), .B(n18327), .Z(n18275) );
  IV U18312 ( .A(n18221), .Z(n18234) );
  XOR U18313 ( .A(n18280), .B(n18279), .Z(n18269) );
  XNOR U18314 ( .A(n18328), .B(n18276), .Z(n18279) );
  XOR U18315 ( .A(n18329), .B(n18330), .Z(n18276) );
  AND U18316 ( .A(n18331), .B(n18332), .Z(n18330) );
  XNOR U18317 ( .A(n18333), .B(n18334), .Z(n18331) );
  XNOR U18318 ( .A(n18335), .B(n18336), .Z(n18328) );
  NOR U18319 ( .A(n18337), .B(n18338), .Z(n18336) );
  XOR U18320 ( .A(n18335), .B(n18339), .Z(n18337) );
  XOR U18321 ( .A(n18340), .B(n18341), .Z(n18280) );
  AND U18322 ( .A(n18342), .B(n18343), .Z(n18341) );
  XOR U18323 ( .A(n18340), .B(n18344), .Z(n18342) );
  XNOR U18324 ( .A(n18345), .B(n18299), .Z(n18301) );
  IV U18325 ( .A(n18116), .Z(n18345) );
  XOR U18326 ( .A(n18346), .B(n18293), .Z(n18116) );
  XOR U18327 ( .A(n18286), .B(n18285), .Z(n18293) );
  XNOR U18328 ( .A(n18347), .B(n18282), .Z(n18285) );
  XOR U18329 ( .A(n18348), .B(n18349), .Z(n18282) );
  AND U18330 ( .A(n18350), .B(n18351), .Z(n18349) );
  XOR U18331 ( .A(n18348), .B(n18352), .Z(n18350) );
  XNOR U18332 ( .A(n18353), .B(n18354), .Z(n18347) );
  NOR U18333 ( .A(n18355), .B(n18356), .Z(n18354) );
  XNOR U18334 ( .A(n18353), .B(n18357), .Z(n18355) );
  XOR U18335 ( .A(n18358), .B(n18359), .Z(n18286) );
  NOR U18336 ( .A(n18360), .B(n18361), .Z(n18359) );
  XNOR U18337 ( .A(n18358), .B(n18362), .Z(n18360) );
  XNOR U18338 ( .A(n18292), .B(n18287), .Z(n18346) );
  AND U18339 ( .A(n18232), .B(n18363), .Z(n18287) );
  XOR U18340 ( .A(n18364), .B(n18298), .Z(n18292) );
  XNOR U18341 ( .A(n18365), .B(n18366), .Z(n18298) );
  NOR U18342 ( .A(n18367), .B(n18368), .Z(n18366) );
  XNOR U18343 ( .A(n18365), .B(n18369), .Z(n18367) );
  XNOR U18344 ( .A(n18297), .B(n18289), .Z(n18364) );
  XOR U18345 ( .A(n18370), .B(n18371), .Z(n18289) );
  AND U18346 ( .A(n18372), .B(n18373), .Z(n18371) );
  XOR U18347 ( .A(n18370), .B(n18374), .Z(n18372) );
  XNOR U18348 ( .A(n18375), .B(n18294), .Z(n18297) );
  XOR U18349 ( .A(n18376), .B(n18377), .Z(n18294) );
  AND U18350 ( .A(n18378), .B(n18379), .Z(n18377) );
  XOR U18351 ( .A(n18376), .B(n18380), .Z(n18378) );
  XNOR U18352 ( .A(n18381), .B(n18382), .Z(n18375) );
  NOR U18353 ( .A(n18383), .B(n18384), .Z(n18382) );
  XOR U18354 ( .A(n18381), .B(n18385), .Z(n18383) );
  AND U18355 ( .A(n18232), .B(n18221), .Z(n18299) );
  XNOR U18356 ( .A(n18386), .B(n18327), .Z(n18221) );
  XOR U18357 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(
        p_input[1024]), .Z(n18327) );
  XOR U18358 ( .A(n18314), .B(n18313), .Z(n18386) );
  XNOR U18359 ( .A(n18387), .B(n18321), .Z(n18313) );
  XOR U18360 ( .A(n18309), .B(n18308), .Z(n18321) );
  XNOR U18361 ( .A(n18388), .B(n18305), .Z(n18308) );
  XOR U18362 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(
        p_input[1034]), .Z(n18305) );
  XNOR U18363 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(
        p_input[1035]), .Z(n18388) );
  XOR U18364 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(
        p_input[1036]), .Z(n18309) );
  XNOR U18365 ( .A(n18319), .B(n18310), .Z(n18387) );
  XOR U18366 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(
        p_input[1025]), .Z(n18310) );
  XOR U18367 ( .A(n18389), .B(n18326), .Z(n18319) );
  XOR U18368 ( .A(n5206), .B(p_input[1039]), .Z(n18326) );
  IV U18369 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .Z(n5206) );
  XNOR U18370 ( .A(n18316), .B(n18325), .Z(n18389) );
  XNOR U18371 ( .A(n18390), .B(n18322), .Z(n18325) );
  XOR U18372 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(
        p_input[1037]), .Z(n18322) );
  XNOR U18373 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(
        p_input[1038]), .Z(n18390) );
  IV U18374 ( .A(n18320), .Z(n18316) );
  XOR U18375 ( .A(n708), .B(p_input[1033]), .Z(n18320) );
  IV U18376 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .Z(n708) );
  XNOR U18377 ( .A(n18334), .B(n18332), .Z(n18314) );
  XOR U18378 ( .A(n18391), .B(n18339), .Z(n18332) );
  XOR U18379 ( .A(n1209), .B(p_input[1032]), .Z(n18339) );
  IV U18380 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .Z(n1209) );
  XOR U18381 ( .A(n18329), .B(n18338), .Z(n18391) );
  XOR U18382 ( .A(n18392), .B(n18335), .Z(n18338) );
  XNOR U18383 ( .A(n2207), .B(p_input[1030]), .Z(n18335) );
  IV U18384 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .Z(n2207) );
  XNOR U18385 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(
        p_input[1031]), .Z(n18392) );
  IV U18386 ( .A(n18333), .Z(n18329) );
  XOR U18387 ( .A(n4205), .B(p_input[1026]), .Z(n18333) );
  IV U18388 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n4205) );
  XOR U18389 ( .A(n18344), .B(n18343), .Z(n18334) );
  XNOR U18390 ( .A(n18393), .B(n18340), .Z(n18343) );
  XOR U18391 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .B(
        p_input[1027]), .Z(n18340) );
  XOR U18392 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(n9328), 
        .Z(n18393) );
  XNOR U18393 ( .A(n2706), .B(p_input[1029]), .Z(n18344) );
  IV U18394 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .Z(n2706) );
  XOR U18395 ( .A(n18394), .B(n18374), .Z(n18232) );
  XOR U18396 ( .A(n18352), .B(n18351), .Z(n18374) );
  XNOR U18397 ( .A(n18395), .B(n18357), .Z(n18351) );
  XNOR U18398 ( .A(n1213), .B(p_input[1032]), .Z(n18357) );
  IV U18399 ( .A(\knn_comb_/min_val_out[0][8] ), .Z(n1213) );
  XOR U18400 ( .A(n18348), .B(n18356), .Z(n18395) );
  XOR U18401 ( .A(n18396), .B(n18353), .Z(n18356) );
  XNOR U18402 ( .A(n2211), .B(p_input[1030]), .Z(n18353) );
  IV U18403 ( .A(\knn_comb_/min_val_out[0][6] ), .Z(n2211) );
  XNOR U18404 ( .A(\knn_comb_/min_val_out[0][7] ), .B(p_input[1031]), .Z(
        n18396) );
  XNOR U18405 ( .A(n4209), .B(p_input[1026]), .Z(n18348) );
  IV U18406 ( .A(\knn_comb_/min_val_out[0][2] ), .Z(n4209) );
  XNOR U18407 ( .A(n18362), .B(n18361), .Z(n18352) );
  XOR U18408 ( .A(n18397), .B(n18358), .Z(n18361) );
  XNOR U18409 ( .A(n3710), .B(p_input[1027]), .Z(n18358) );
  IV U18410 ( .A(\knn_comb_/min_val_out[0][3] ), .Z(n3710) );
  XOR U18411 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n9328), .Z(n18397) );
  IV U18412 ( .A(p_input[1028]), .Z(n9328) );
  XNOR U18413 ( .A(n2710), .B(p_input[1029]), .Z(n18362) );
  IV U18414 ( .A(\knn_comb_/min_val_out[0][5] ), .Z(n2710) );
  XNOR U18415 ( .A(n18373), .B(n18363), .Z(n18394) );
  XOR U18416 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[1024]), .Z(n18363) );
  XNOR U18417 ( .A(n18398), .B(n18380), .Z(n18373) );
  XNOR U18418 ( .A(n18369), .B(n18368), .Z(n18380) );
  XOR U18419 ( .A(n18399), .B(n18365), .Z(n18368) );
  XOR U18420 ( .A(\knn_comb_/min_val_out[0][10] ), .B(p_input[1034]), .Z(
        n18365) );
  XNOR U18421 ( .A(\knn_comb_/min_val_out[0][11] ), .B(p_input[1035]), .Z(
        n18399) );
  XOR U18422 ( .A(\knn_comb_/min_val_out[0][12] ), .B(p_input[1036]), .Z(
        n18369) );
  XNOR U18423 ( .A(n18379), .B(n18370), .Z(n18398) );
  XNOR U18424 ( .A(n4708), .B(p_input[1025]), .Z(n18370) );
  IV U18425 ( .A(\knn_comb_/min_val_out[0][1] ), .Z(n4708) );
  XOR U18426 ( .A(n18400), .B(n18385), .Z(n18379) );
  XNOR U18427 ( .A(\knn_comb_/min_val_out[0][15] ), .B(p_input[1039]), .Z(
        n18385) );
  XOR U18428 ( .A(n18376), .B(n18384), .Z(n18400) );
  XOR U18429 ( .A(n18401), .B(n18381), .Z(n18384) );
  XOR U18430 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[1037]), .Z(
        n18381) );
  XNOR U18431 ( .A(\knn_comb_/min_val_out[0][14] ), .B(p_input[1038]), .Z(
        n18401) );
  XNOR U18432 ( .A(n714), .B(p_input[1033]), .Z(n18376) );
  IV U18433 ( .A(\knn_comb_/min_val_out[0][9] ), .Z(n714) );
endmodule

