
module auction_BMR_N4_W16 ( p_input, o );
  input [255:0] p_input;
  output [19:0] o;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704;

  XNOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  AND U2 ( .A(o[3]), .B(n3), .Z(n1) );
  XOR U3 ( .A(n2), .B(n4), .Z(n3) );
  XOR U4 ( .A(n5), .B(n6), .Z(o[8]) );
  AND U5 ( .A(o[3]), .B(n7), .Z(n5) );
  XOR U6 ( .A(n8), .B(n9), .Z(n7) );
  XOR U7 ( .A(n10), .B(n11), .Z(o[7]) );
  AND U8 ( .A(o[3]), .B(n12), .Z(n10) );
  XOR U9 ( .A(n13), .B(n14), .Z(n12) );
  XOR U10 ( .A(n15), .B(n16), .Z(o[6]) );
  AND U11 ( .A(o[3]), .B(n17), .Z(n15) );
  XOR U12 ( .A(n18), .B(n19), .Z(n17) );
  XOR U13 ( .A(n20), .B(n21), .Z(o[5]) );
  AND U14 ( .A(o[3]), .B(n22), .Z(n20) );
  XOR U15 ( .A(n23), .B(n24), .Z(n22) );
  XNOR U16 ( .A(n25), .B(n26), .Z(o[4]) );
  AND U17 ( .A(o[3]), .B(n27), .Z(n25) );
  XNOR U18 ( .A(n28), .B(n26), .Z(n27) );
  XOR U19 ( .A(n29), .B(n30), .Z(o[19]) );
  AND U20 ( .A(n31), .B(o[3]), .Z(n29) );
  AND U21 ( .A(n30), .B(n32), .Z(n31) );
  XOR U22 ( .A(n33), .B(n34), .Z(o[18]) );
  AND U23 ( .A(o[3]), .B(n35), .Z(n33) );
  XOR U24 ( .A(n36), .B(n37), .Z(n35) );
  XOR U25 ( .A(n38), .B(n39), .Z(o[17]) );
  AND U26 ( .A(o[3]), .B(n40), .Z(n38) );
  XOR U27 ( .A(n41), .B(n42), .Z(n40) );
  XOR U28 ( .A(n43), .B(n44), .Z(o[16]) );
  AND U29 ( .A(o[3]), .B(n45), .Z(n43) );
  XOR U30 ( .A(n46), .B(n47), .Z(n45) );
  XOR U31 ( .A(n48), .B(n49), .Z(o[15]) );
  AND U32 ( .A(o[3]), .B(n50), .Z(n48) );
  XOR U33 ( .A(n51), .B(n52), .Z(n50) );
  XOR U34 ( .A(n53), .B(n54), .Z(o[14]) );
  AND U35 ( .A(o[3]), .B(n55), .Z(n53) );
  XOR U36 ( .A(n56), .B(n57), .Z(n55) );
  XOR U37 ( .A(n58), .B(n59), .Z(o[13]) );
  AND U38 ( .A(o[3]), .B(n60), .Z(n58) );
  XOR U39 ( .A(n61), .B(n62), .Z(n60) );
  XOR U40 ( .A(n63), .B(n64), .Z(o[12]) );
  AND U41 ( .A(o[3]), .B(n65), .Z(n63) );
  XOR U42 ( .A(n66), .B(n67), .Z(n65) );
  XOR U43 ( .A(n68), .B(n69), .Z(o[11]) );
  AND U44 ( .A(o[3]), .B(n70), .Z(n68) );
  XOR U45 ( .A(n71), .B(n72), .Z(n70) );
  XOR U46 ( .A(n73), .B(n74), .Z(o[10]) );
  AND U47 ( .A(o[3]), .B(n75), .Z(n73) );
  XOR U48 ( .A(n76), .B(n77), .Z(n75) );
  XOR U49 ( .A(n78), .B(n79), .Z(o[0]) );
  AND U50 ( .A(o[1]), .B(n80), .Z(n79) );
  XNOR U51 ( .A(n81), .B(n82), .Z(n80) );
  XNOR U52 ( .A(n83), .B(n78), .Z(n82) );
  AND U53 ( .A(o[2]), .B(n84), .Z(n83) );
  XNOR U54 ( .A(n81), .B(n85), .Z(n84) );
  XNOR U55 ( .A(n86), .B(n87), .Z(n85) );
  AND U56 ( .A(o[3]), .B(n88), .Z(n86) );
  XOR U57 ( .A(n87), .B(n89), .Z(n88) );
  XOR U58 ( .A(n90), .B(n91), .Z(n81) );
  AND U59 ( .A(o[3]), .B(n92), .Z(n91) );
  XOR U60 ( .A(n90), .B(n93), .Z(n92) );
  XOR U61 ( .A(n94), .B(n95), .Z(o[1]) );
  AND U62 ( .A(o[2]), .B(n96), .Z(n95) );
  XNOR U63 ( .A(n94), .B(n97), .Z(n96) );
  XNOR U64 ( .A(n98), .B(n99), .Z(n97) );
  AND U65 ( .A(o[3]), .B(n100), .Z(n98) );
  XOR U66 ( .A(n99), .B(n101), .Z(n100) );
  XOR U67 ( .A(n102), .B(n103), .Z(n94) );
  AND U68 ( .A(o[3]), .B(n104), .Z(n103) );
  XOR U69 ( .A(n102), .B(n105), .Z(n104) );
  XOR U70 ( .A(n106), .B(n107), .Z(n78) );
  AND U71 ( .A(o[2]), .B(n108), .Z(n107) );
  XNOR U72 ( .A(n106), .B(n109), .Z(n108) );
  XNOR U73 ( .A(n110), .B(n111), .Z(n109) );
  AND U74 ( .A(o[3]), .B(n112), .Z(n110) );
  XOR U75 ( .A(n111), .B(n113), .Z(n112) );
  XOR U76 ( .A(n114), .B(n115), .Z(o[2]) );
  AND U77 ( .A(o[3]), .B(n116), .Z(n115) );
  XOR U78 ( .A(n114), .B(n117), .Z(n116) );
  XOR U79 ( .A(n118), .B(n119), .Z(n106) );
  AND U80 ( .A(o[3]), .B(n120), .Z(n119) );
  XOR U81 ( .A(n118), .B(n121), .Z(n120) );
  XOR U82 ( .A(n122), .B(n123), .Z(o[3]) );
  AND U83 ( .A(n124), .B(n125), .Z(n123) );
  XOR U84 ( .A(n32), .B(n122), .Z(n125) );
  IV U85 ( .A(n126), .Z(n32) );
  AND U86 ( .A(n127), .B(n128), .Z(n126) );
  XOR U87 ( .A(n122), .B(n30), .Z(n124) );
  AND U88 ( .A(n129), .B(n130), .Z(n30) );
  XOR U89 ( .A(n131), .B(n132), .Z(n122) );
  AND U90 ( .A(n133), .B(n134), .Z(n132) );
  XOR U91 ( .A(n131), .B(n36), .Z(n134) );
  XOR U92 ( .A(n135), .B(n136), .Z(n36) );
  AND U93 ( .A(n117), .B(n137), .Z(n136) );
  XOR U94 ( .A(n138), .B(n135), .Z(n137) );
  XNOR U95 ( .A(n37), .B(n131), .Z(n133) );
  IV U96 ( .A(n34), .Z(n37) );
  XNOR U97 ( .A(n139), .B(n140), .Z(n34) );
  AND U98 ( .A(n114), .B(n141), .Z(n140) );
  XOR U99 ( .A(n142), .B(n139), .Z(n141) );
  XOR U100 ( .A(n143), .B(n144), .Z(n131) );
  AND U101 ( .A(n145), .B(n146), .Z(n144) );
  XOR U102 ( .A(n143), .B(n41), .Z(n146) );
  XOR U103 ( .A(n147), .B(n148), .Z(n41) );
  AND U104 ( .A(n117), .B(n149), .Z(n148) );
  XOR U105 ( .A(n150), .B(n147), .Z(n149) );
  XNOR U106 ( .A(n42), .B(n143), .Z(n145) );
  IV U107 ( .A(n39), .Z(n42) );
  XNOR U108 ( .A(n151), .B(n152), .Z(n39) );
  AND U109 ( .A(n114), .B(n153), .Z(n152) );
  XOR U110 ( .A(n154), .B(n151), .Z(n153) );
  XOR U111 ( .A(n155), .B(n156), .Z(n143) );
  AND U112 ( .A(n157), .B(n158), .Z(n156) );
  XOR U113 ( .A(n155), .B(n46), .Z(n158) );
  XOR U114 ( .A(n159), .B(n160), .Z(n46) );
  AND U115 ( .A(n117), .B(n161), .Z(n160) );
  XOR U116 ( .A(n162), .B(n159), .Z(n161) );
  XNOR U117 ( .A(n47), .B(n155), .Z(n157) );
  IV U118 ( .A(n44), .Z(n47) );
  XNOR U119 ( .A(n163), .B(n164), .Z(n44) );
  AND U120 ( .A(n114), .B(n165), .Z(n164) );
  XOR U121 ( .A(n166), .B(n163), .Z(n165) );
  XOR U122 ( .A(n167), .B(n168), .Z(n155) );
  AND U123 ( .A(n169), .B(n170), .Z(n168) );
  XOR U124 ( .A(n167), .B(n51), .Z(n170) );
  XOR U125 ( .A(n171), .B(n172), .Z(n51) );
  AND U126 ( .A(n117), .B(n173), .Z(n172) );
  XOR U127 ( .A(n174), .B(n171), .Z(n173) );
  XNOR U128 ( .A(n52), .B(n167), .Z(n169) );
  IV U129 ( .A(n49), .Z(n52) );
  XNOR U130 ( .A(n175), .B(n176), .Z(n49) );
  AND U131 ( .A(n114), .B(n177), .Z(n176) );
  XOR U132 ( .A(n178), .B(n175), .Z(n177) );
  XOR U133 ( .A(n179), .B(n180), .Z(n167) );
  AND U134 ( .A(n181), .B(n182), .Z(n180) );
  XOR U135 ( .A(n179), .B(n56), .Z(n182) );
  XOR U136 ( .A(n183), .B(n184), .Z(n56) );
  AND U137 ( .A(n117), .B(n185), .Z(n184) );
  XOR U138 ( .A(n186), .B(n183), .Z(n185) );
  XNOR U139 ( .A(n57), .B(n179), .Z(n181) );
  IV U140 ( .A(n54), .Z(n57) );
  XNOR U141 ( .A(n187), .B(n188), .Z(n54) );
  AND U142 ( .A(n114), .B(n189), .Z(n188) );
  XOR U143 ( .A(n190), .B(n187), .Z(n189) );
  XOR U144 ( .A(n191), .B(n192), .Z(n179) );
  AND U145 ( .A(n193), .B(n194), .Z(n192) );
  XOR U146 ( .A(n191), .B(n61), .Z(n194) );
  XOR U147 ( .A(n195), .B(n196), .Z(n61) );
  AND U148 ( .A(n117), .B(n197), .Z(n196) );
  XOR U149 ( .A(n198), .B(n195), .Z(n197) );
  XNOR U150 ( .A(n62), .B(n191), .Z(n193) );
  IV U151 ( .A(n59), .Z(n62) );
  XNOR U152 ( .A(n199), .B(n200), .Z(n59) );
  AND U153 ( .A(n114), .B(n201), .Z(n200) );
  XOR U154 ( .A(n202), .B(n199), .Z(n201) );
  XOR U155 ( .A(n203), .B(n204), .Z(n191) );
  AND U156 ( .A(n205), .B(n206), .Z(n204) );
  XOR U157 ( .A(n203), .B(n66), .Z(n206) );
  XOR U158 ( .A(n207), .B(n208), .Z(n66) );
  AND U159 ( .A(n117), .B(n209), .Z(n208) );
  XOR U160 ( .A(n210), .B(n207), .Z(n209) );
  XNOR U161 ( .A(n67), .B(n203), .Z(n205) );
  IV U162 ( .A(n64), .Z(n67) );
  XNOR U163 ( .A(n211), .B(n212), .Z(n64) );
  AND U164 ( .A(n114), .B(n213), .Z(n212) );
  XOR U165 ( .A(n214), .B(n211), .Z(n213) );
  XOR U166 ( .A(n215), .B(n216), .Z(n203) );
  AND U167 ( .A(n217), .B(n218), .Z(n216) );
  XOR U168 ( .A(n215), .B(n71), .Z(n218) );
  XOR U169 ( .A(n219), .B(n220), .Z(n71) );
  AND U170 ( .A(n117), .B(n221), .Z(n220) );
  XOR U171 ( .A(n222), .B(n219), .Z(n221) );
  XNOR U172 ( .A(n72), .B(n215), .Z(n217) );
  IV U173 ( .A(n69), .Z(n72) );
  XNOR U174 ( .A(n223), .B(n224), .Z(n69) );
  AND U175 ( .A(n114), .B(n225), .Z(n224) );
  XOR U176 ( .A(n226), .B(n223), .Z(n225) );
  XOR U177 ( .A(n227), .B(n228), .Z(n215) );
  AND U178 ( .A(n229), .B(n230), .Z(n228) );
  XOR U179 ( .A(n227), .B(n76), .Z(n230) );
  XOR U180 ( .A(n231), .B(n232), .Z(n76) );
  AND U181 ( .A(n117), .B(n233), .Z(n232) );
  XOR U182 ( .A(n234), .B(n231), .Z(n233) );
  XNOR U183 ( .A(n77), .B(n227), .Z(n229) );
  IV U184 ( .A(n74), .Z(n77) );
  XNOR U185 ( .A(n235), .B(n236), .Z(n74) );
  AND U186 ( .A(n114), .B(n237), .Z(n236) );
  XOR U187 ( .A(n238), .B(n235), .Z(n237) );
  XOR U188 ( .A(n239), .B(n240), .Z(n227) );
  AND U189 ( .A(n241), .B(n242), .Z(n240) );
  XOR U190 ( .A(n4), .B(n239), .Z(n242) );
  XOR U191 ( .A(n243), .B(n244), .Z(n4) );
  AND U192 ( .A(n117), .B(n245), .Z(n244) );
  XOR U193 ( .A(n243), .B(n246), .Z(n245) );
  XNOR U194 ( .A(n239), .B(n2), .Z(n241) );
  XOR U195 ( .A(n247), .B(n248), .Z(n2) );
  AND U196 ( .A(n114), .B(n249), .Z(n248) );
  XOR U197 ( .A(n247), .B(n250), .Z(n249) );
  XOR U198 ( .A(n251), .B(n252), .Z(n239) );
  AND U199 ( .A(n253), .B(n254), .Z(n252) );
  XOR U200 ( .A(n251), .B(n8), .Z(n254) );
  XOR U201 ( .A(n255), .B(n256), .Z(n8) );
  AND U202 ( .A(n117), .B(n257), .Z(n256) );
  XOR U203 ( .A(n258), .B(n255), .Z(n257) );
  XNOR U204 ( .A(n9), .B(n251), .Z(n253) );
  IV U205 ( .A(n6), .Z(n9) );
  XNOR U206 ( .A(n259), .B(n260), .Z(n6) );
  AND U207 ( .A(n114), .B(n261), .Z(n260) );
  XOR U208 ( .A(n262), .B(n259), .Z(n261) );
  XOR U209 ( .A(n263), .B(n264), .Z(n251) );
  AND U210 ( .A(n265), .B(n266), .Z(n264) );
  XOR U211 ( .A(n263), .B(n13), .Z(n266) );
  XOR U212 ( .A(n267), .B(n268), .Z(n13) );
  AND U213 ( .A(n117), .B(n269), .Z(n268) );
  XOR U214 ( .A(n270), .B(n267), .Z(n269) );
  XNOR U215 ( .A(n14), .B(n263), .Z(n265) );
  IV U216 ( .A(n11), .Z(n14) );
  XNOR U217 ( .A(n271), .B(n272), .Z(n11) );
  AND U218 ( .A(n114), .B(n273), .Z(n272) );
  XOR U219 ( .A(n274), .B(n271), .Z(n273) );
  XOR U220 ( .A(n275), .B(n276), .Z(n263) );
  AND U221 ( .A(n277), .B(n278), .Z(n276) );
  XOR U222 ( .A(n275), .B(n18), .Z(n278) );
  XOR U223 ( .A(n279), .B(n280), .Z(n18) );
  AND U224 ( .A(n117), .B(n281), .Z(n280) );
  XOR U225 ( .A(n282), .B(n279), .Z(n281) );
  XNOR U226 ( .A(n19), .B(n275), .Z(n277) );
  IV U227 ( .A(n16), .Z(n19) );
  XNOR U228 ( .A(n283), .B(n284), .Z(n16) );
  AND U229 ( .A(n114), .B(n285), .Z(n284) );
  XOR U230 ( .A(n286), .B(n283), .Z(n285) );
  XNOR U231 ( .A(n287), .B(n288), .Z(n275) );
  AND U232 ( .A(n289), .B(n290), .Z(n288) );
  XNOR U233 ( .A(n287), .B(n23), .Z(n290) );
  XOR U234 ( .A(n291), .B(n292), .Z(n23) );
  AND U235 ( .A(n117), .B(n293), .Z(n292) );
  XOR U236 ( .A(n294), .B(n291), .Z(n293) );
  XOR U237 ( .A(n24), .B(n287), .Z(n289) );
  IV U238 ( .A(n21), .Z(n24) );
  XNOR U239 ( .A(n295), .B(n296), .Z(n21) );
  AND U240 ( .A(n114), .B(n297), .Z(n296) );
  XOR U241 ( .A(n298), .B(n295), .Z(n297) );
  AND U242 ( .A(n26), .B(n28), .Z(n287) );
  XNOR U243 ( .A(n299), .B(n300), .Z(n28) );
  AND U244 ( .A(n117), .B(n301), .Z(n300) );
  XNOR U245 ( .A(n302), .B(n299), .Z(n301) );
  XOR U246 ( .A(n303), .B(n304), .Z(n117) );
  AND U247 ( .A(n305), .B(n306), .Z(n304) );
  XNOR U248 ( .A(n127), .B(n303), .Z(n306) );
  AND U249 ( .A(n307), .B(n308), .Z(n127) );
  XOR U250 ( .A(n303), .B(n128), .Z(n305) );
  AND U251 ( .A(n309), .B(n310), .Z(n128) );
  XOR U252 ( .A(n311), .B(n312), .Z(n303) );
  AND U253 ( .A(n313), .B(n314), .Z(n312) );
  XOR U254 ( .A(n311), .B(n138), .Z(n314) );
  XOR U255 ( .A(n315), .B(n316), .Z(n138) );
  AND U256 ( .A(n101), .B(n317), .Z(n316) );
  XOR U257 ( .A(n318), .B(n315), .Z(n317) );
  XNOR U258 ( .A(n135), .B(n311), .Z(n313) );
  XOR U259 ( .A(n319), .B(n320), .Z(n135) );
  AND U260 ( .A(n99), .B(n321), .Z(n320) );
  XOR U261 ( .A(n322), .B(n319), .Z(n321) );
  XOR U262 ( .A(n323), .B(n324), .Z(n311) );
  AND U263 ( .A(n325), .B(n326), .Z(n324) );
  XOR U264 ( .A(n323), .B(n150), .Z(n326) );
  XOR U265 ( .A(n327), .B(n328), .Z(n150) );
  AND U266 ( .A(n101), .B(n329), .Z(n328) );
  XOR U267 ( .A(n330), .B(n327), .Z(n329) );
  XNOR U268 ( .A(n147), .B(n323), .Z(n325) );
  XOR U269 ( .A(n331), .B(n332), .Z(n147) );
  AND U270 ( .A(n99), .B(n333), .Z(n332) );
  XOR U271 ( .A(n334), .B(n331), .Z(n333) );
  XOR U272 ( .A(n335), .B(n336), .Z(n323) );
  AND U273 ( .A(n337), .B(n338), .Z(n336) );
  XOR U274 ( .A(n335), .B(n162), .Z(n338) );
  XOR U275 ( .A(n339), .B(n340), .Z(n162) );
  AND U276 ( .A(n101), .B(n341), .Z(n340) );
  XOR U277 ( .A(n342), .B(n339), .Z(n341) );
  XNOR U278 ( .A(n159), .B(n335), .Z(n337) );
  XOR U279 ( .A(n343), .B(n344), .Z(n159) );
  AND U280 ( .A(n99), .B(n345), .Z(n344) );
  XOR U281 ( .A(n346), .B(n343), .Z(n345) );
  XOR U282 ( .A(n347), .B(n348), .Z(n335) );
  AND U283 ( .A(n349), .B(n350), .Z(n348) );
  XOR U284 ( .A(n347), .B(n174), .Z(n350) );
  XOR U285 ( .A(n351), .B(n352), .Z(n174) );
  AND U286 ( .A(n101), .B(n353), .Z(n352) );
  XOR U287 ( .A(n354), .B(n351), .Z(n353) );
  XNOR U288 ( .A(n171), .B(n347), .Z(n349) );
  XOR U289 ( .A(n355), .B(n356), .Z(n171) );
  AND U290 ( .A(n99), .B(n357), .Z(n356) );
  XOR U291 ( .A(n358), .B(n355), .Z(n357) );
  XOR U292 ( .A(n359), .B(n360), .Z(n347) );
  AND U293 ( .A(n361), .B(n362), .Z(n360) );
  XOR U294 ( .A(n359), .B(n186), .Z(n362) );
  XOR U295 ( .A(n363), .B(n364), .Z(n186) );
  AND U296 ( .A(n101), .B(n365), .Z(n364) );
  XOR U297 ( .A(n366), .B(n363), .Z(n365) );
  XNOR U298 ( .A(n183), .B(n359), .Z(n361) );
  XOR U299 ( .A(n367), .B(n368), .Z(n183) );
  AND U300 ( .A(n99), .B(n369), .Z(n368) );
  XOR U301 ( .A(n370), .B(n367), .Z(n369) );
  XOR U302 ( .A(n371), .B(n372), .Z(n359) );
  AND U303 ( .A(n373), .B(n374), .Z(n372) );
  XOR U304 ( .A(n371), .B(n198), .Z(n374) );
  XOR U305 ( .A(n375), .B(n376), .Z(n198) );
  AND U306 ( .A(n101), .B(n377), .Z(n376) );
  XOR U307 ( .A(n378), .B(n375), .Z(n377) );
  XNOR U308 ( .A(n195), .B(n371), .Z(n373) );
  XOR U309 ( .A(n379), .B(n380), .Z(n195) );
  AND U310 ( .A(n99), .B(n381), .Z(n380) );
  XOR U311 ( .A(n382), .B(n379), .Z(n381) );
  XOR U312 ( .A(n383), .B(n384), .Z(n371) );
  AND U313 ( .A(n385), .B(n386), .Z(n384) );
  XOR U314 ( .A(n383), .B(n210), .Z(n386) );
  XOR U315 ( .A(n387), .B(n388), .Z(n210) );
  AND U316 ( .A(n101), .B(n389), .Z(n388) );
  XOR U317 ( .A(n390), .B(n387), .Z(n389) );
  XNOR U318 ( .A(n207), .B(n383), .Z(n385) );
  XOR U319 ( .A(n391), .B(n392), .Z(n207) );
  AND U320 ( .A(n99), .B(n393), .Z(n392) );
  XOR U321 ( .A(n394), .B(n391), .Z(n393) );
  XOR U322 ( .A(n395), .B(n396), .Z(n383) );
  AND U323 ( .A(n397), .B(n398), .Z(n396) );
  XOR U324 ( .A(n395), .B(n222), .Z(n398) );
  XOR U325 ( .A(n399), .B(n400), .Z(n222) );
  AND U326 ( .A(n101), .B(n401), .Z(n400) );
  XOR U327 ( .A(n402), .B(n399), .Z(n401) );
  XNOR U328 ( .A(n219), .B(n395), .Z(n397) );
  XOR U329 ( .A(n403), .B(n404), .Z(n219) );
  AND U330 ( .A(n99), .B(n405), .Z(n404) );
  XOR U331 ( .A(n406), .B(n403), .Z(n405) );
  XOR U332 ( .A(n407), .B(n408), .Z(n395) );
  AND U333 ( .A(n409), .B(n410), .Z(n408) );
  XOR U334 ( .A(n407), .B(n234), .Z(n410) );
  XOR U335 ( .A(n411), .B(n412), .Z(n234) );
  AND U336 ( .A(n101), .B(n413), .Z(n412) );
  XOR U337 ( .A(n414), .B(n411), .Z(n413) );
  XNOR U338 ( .A(n231), .B(n407), .Z(n409) );
  XOR U339 ( .A(n415), .B(n416), .Z(n231) );
  AND U340 ( .A(n99), .B(n417), .Z(n416) );
  XOR U341 ( .A(n418), .B(n415), .Z(n417) );
  XOR U342 ( .A(n419), .B(n420), .Z(n407) );
  AND U343 ( .A(n421), .B(n422), .Z(n420) );
  XOR U344 ( .A(n246), .B(n419), .Z(n422) );
  XOR U345 ( .A(n423), .B(n424), .Z(n246) );
  AND U346 ( .A(n101), .B(n425), .Z(n424) );
  XOR U347 ( .A(n423), .B(n426), .Z(n425) );
  XNOR U348 ( .A(n419), .B(n243), .Z(n421) );
  XOR U349 ( .A(n427), .B(n428), .Z(n243) );
  AND U350 ( .A(n99), .B(n429), .Z(n428) );
  XOR U351 ( .A(n427), .B(n430), .Z(n429) );
  XOR U352 ( .A(n431), .B(n432), .Z(n419) );
  AND U353 ( .A(n433), .B(n434), .Z(n432) );
  XOR U354 ( .A(n431), .B(n258), .Z(n434) );
  XOR U355 ( .A(n435), .B(n436), .Z(n258) );
  AND U356 ( .A(n101), .B(n437), .Z(n436) );
  XOR U357 ( .A(n438), .B(n435), .Z(n437) );
  XNOR U358 ( .A(n255), .B(n431), .Z(n433) );
  XOR U359 ( .A(n439), .B(n440), .Z(n255) );
  AND U360 ( .A(n99), .B(n441), .Z(n440) );
  XOR U361 ( .A(n442), .B(n439), .Z(n441) );
  XOR U362 ( .A(n443), .B(n444), .Z(n431) );
  AND U363 ( .A(n445), .B(n446), .Z(n444) );
  XOR U364 ( .A(n443), .B(n270), .Z(n446) );
  XOR U365 ( .A(n447), .B(n448), .Z(n270) );
  AND U366 ( .A(n101), .B(n449), .Z(n448) );
  XOR U367 ( .A(n450), .B(n447), .Z(n449) );
  XNOR U368 ( .A(n267), .B(n443), .Z(n445) );
  XOR U369 ( .A(n451), .B(n452), .Z(n267) );
  AND U370 ( .A(n99), .B(n453), .Z(n452) );
  XOR U371 ( .A(n454), .B(n451), .Z(n453) );
  XOR U372 ( .A(n455), .B(n456), .Z(n443) );
  AND U373 ( .A(n457), .B(n458), .Z(n456) );
  XOR U374 ( .A(n455), .B(n282), .Z(n458) );
  XOR U375 ( .A(n459), .B(n460), .Z(n282) );
  AND U376 ( .A(n101), .B(n461), .Z(n460) );
  XOR U377 ( .A(n462), .B(n459), .Z(n461) );
  XNOR U378 ( .A(n279), .B(n455), .Z(n457) );
  XOR U379 ( .A(n463), .B(n464), .Z(n279) );
  AND U380 ( .A(n99), .B(n465), .Z(n464) );
  XOR U381 ( .A(n466), .B(n463), .Z(n465) );
  XOR U382 ( .A(n467), .B(n468), .Z(n455) );
  AND U383 ( .A(n469), .B(n470), .Z(n468) );
  XNOR U384 ( .A(n471), .B(n294), .Z(n470) );
  XOR U385 ( .A(n472), .B(n473), .Z(n294) );
  AND U386 ( .A(n101), .B(n474), .Z(n473) );
  XOR U387 ( .A(n475), .B(n472), .Z(n474) );
  XNOR U388 ( .A(n291), .B(n467), .Z(n469) );
  XOR U389 ( .A(n476), .B(n477), .Z(n291) );
  AND U390 ( .A(n99), .B(n478), .Z(n477) );
  XOR U391 ( .A(n479), .B(n476), .Z(n478) );
  IV U392 ( .A(n471), .Z(n467) );
  AND U393 ( .A(n299), .B(n302), .Z(n471) );
  XNOR U394 ( .A(n480), .B(n481), .Z(n302) );
  AND U395 ( .A(n101), .B(n482), .Z(n481) );
  XNOR U396 ( .A(n483), .B(n480), .Z(n482) );
  XOR U397 ( .A(n484), .B(n485), .Z(n101) );
  AND U398 ( .A(n486), .B(n487), .Z(n485) );
  XNOR U399 ( .A(n307), .B(n484), .Z(n487) );
  AND U400 ( .A(p_input[255]), .B(p_input[239]), .Z(n307) );
  XOR U401 ( .A(n484), .B(n308), .Z(n486) );
  AND U402 ( .A(p_input[223]), .B(p_input[207]), .Z(n308) );
  XOR U403 ( .A(n488), .B(n489), .Z(n484) );
  AND U404 ( .A(n490), .B(n491), .Z(n489) );
  XOR U405 ( .A(n488), .B(n318), .Z(n491) );
  XNOR U406 ( .A(p_input[238]), .B(n492), .Z(n318) );
  AND U407 ( .A(n89), .B(n493), .Z(n492) );
  XOR U408 ( .A(p_input[254]), .B(p_input[238]), .Z(n493) );
  XNOR U409 ( .A(n315), .B(n488), .Z(n490) );
  XOR U410 ( .A(n494), .B(n495), .Z(n315) );
  AND U411 ( .A(n87), .B(n496), .Z(n495) );
  XOR U412 ( .A(p_input[222]), .B(p_input[206]), .Z(n496) );
  XOR U413 ( .A(n497), .B(n498), .Z(n488) );
  AND U414 ( .A(n499), .B(n500), .Z(n498) );
  XOR U415 ( .A(n497), .B(n330), .Z(n500) );
  XNOR U416 ( .A(p_input[237]), .B(n501), .Z(n330) );
  AND U417 ( .A(n89), .B(n502), .Z(n501) );
  XOR U418 ( .A(p_input[253]), .B(p_input[237]), .Z(n502) );
  XNOR U419 ( .A(n327), .B(n497), .Z(n499) );
  XOR U420 ( .A(n503), .B(n504), .Z(n327) );
  AND U421 ( .A(n87), .B(n505), .Z(n504) );
  XOR U422 ( .A(p_input[221]), .B(p_input[205]), .Z(n505) );
  XOR U423 ( .A(n506), .B(n507), .Z(n497) );
  AND U424 ( .A(n508), .B(n509), .Z(n507) );
  XOR U425 ( .A(n506), .B(n342), .Z(n509) );
  XNOR U426 ( .A(p_input[236]), .B(n510), .Z(n342) );
  AND U427 ( .A(n89), .B(n511), .Z(n510) );
  XOR U428 ( .A(p_input[252]), .B(p_input[236]), .Z(n511) );
  XNOR U429 ( .A(n339), .B(n506), .Z(n508) );
  XOR U430 ( .A(n512), .B(n513), .Z(n339) );
  AND U431 ( .A(n87), .B(n514), .Z(n513) );
  XOR U432 ( .A(p_input[220]), .B(p_input[204]), .Z(n514) );
  XOR U433 ( .A(n515), .B(n516), .Z(n506) );
  AND U434 ( .A(n517), .B(n518), .Z(n516) );
  XOR U435 ( .A(n515), .B(n354), .Z(n518) );
  XNOR U436 ( .A(p_input[235]), .B(n519), .Z(n354) );
  AND U437 ( .A(n89), .B(n520), .Z(n519) );
  XOR U438 ( .A(p_input[251]), .B(p_input[235]), .Z(n520) );
  XNOR U439 ( .A(n351), .B(n515), .Z(n517) );
  XOR U440 ( .A(n521), .B(n522), .Z(n351) );
  AND U441 ( .A(n87), .B(n523), .Z(n522) );
  XOR U442 ( .A(p_input[219]), .B(p_input[203]), .Z(n523) );
  XOR U443 ( .A(n524), .B(n525), .Z(n515) );
  AND U444 ( .A(n526), .B(n527), .Z(n525) );
  XOR U445 ( .A(n524), .B(n366), .Z(n527) );
  XNOR U446 ( .A(p_input[234]), .B(n528), .Z(n366) );
  AND U447 ( .A(n89), .B(n529), .Z(n528) );
  XOR U448 ( .A(p_input[250]), .B(p_input[234]), .Z(n529) );
  XNOR U449 ( .A(n363), .B(n524), .Z(n526) );
  XOR U450 ( .A(n530), .B(n531), .Z(n363) );
  AND U451 ( .A(n87), .B(n532), .Z(n531) );
  XOR U452 ( .A(p_input[218]), .B(p_input[202]), .Z(n532) );
  XOR U453 ( .A(n533), .B(n534), .Z(n524) );
  AND U454 ( .A(n535), .B(n536), .Z(n534) );
  XOR U455 ( .A(n533), .B(n378), .Z(n536) );
  XNOR U456 ( .A(p_input[233]), .B(n537), .Z(n378) );
  AND U457 ( .A(n89), .B(n538), .Z(n537) );
  XOR U458 ( .A(p_input[249]), .B(p_input[233]), .Z(n538) );
  XNOR U459 ( .A(n375), .B(n533), .Z(n535) );
  XOR U460 ( .A(n539), .B(n540), .Z(n375) );
  AND U461 ( .A(n87), .B(n541), .Z(n540) );
  XOR U462 ( .A(p_input[217]), .B(p_input[201]), .Z(n541) );
  XOR U463 ( .A(n542), .B(n543), .Z(n533) );
  AND U464 ( .A(n544), .B(n545), .Z(n543) );
  XOR U465 ( .A(n542), .B(n390), .Z(n545) );
  XNOR U466 ( .A(p_input[232]), .B(n546), .Z(n390) );
  AND U467 ( .A(n89), .B(n547), .Z(n546) );
  XOR U468 ( .A(p_input[248]), .B(p_input[232]), .Z(n547) );
  XNOR U469 ( .A(n387), .B(n542), .Z(n544) );
  XOR U470 ( .A(n548), .B(n549), .Z(n387) );
  AND U471 ( .A(n87), .B(n550), .Z(n549) );
  XOR U472 ( .A(p_input[216]), .B(p_input[200]), .Z(n550) );
  XOR U473 ( .A(n551), .B(n552), .Z(n542) );
  AND U474 ( .A(n553), .B(n554), .Z(n552) );
  XOR U475 ( .A(n551), .B(n402), .Z(n554) );
  XNOR U476 ( .A(p_input[231]), .B(n555), .Z(n402) );
  AND U477 ( .A(n89), .B(n556), .Z(n555) );
  XOR U478 ( .A(p_input[247]), .B(p_input[231]), .Z(n556) );
  XNOR U479 ( .A(n399), .B(n551), .Z(n553) );
  XOR U480 ( .A(n557), .B(n558), .Z(n399) );
  AND U481 ( .A(n87), .B(n559), .Z(n558) );
  XOR U482 ( .A(p_input[215]), .B(p_input[199]), .Z(n559) );
  XOR U483 ( .A(n560), .B(n561), .Z(n551) );
  AND U484 ( .A(n562), .B(n563), .Z(n561) );
  XOR U485 ( .A(n560), .B(n414), .Z(n563) );
  XNOR U486 ( .A(p_input[230]), .B(n564), .Z(n414) );
  AND U487 ( .A(n89), .B(n565), .Z(n564) );
  XOR U488 ( .A(p_input[246]), .B(p_input[230]), .Z(n565) );
  XNOR U489 ( .A(n411), .B(n560), .Z(n562) );
  XOR U490 ( .A(n566), .B(n567), .Z(n411) );
  AND U491 ( .A(n87), .B(n568), .Z(n567) );
  XOR U492 ( .A(p_input[214]), .B(p_input[198]), .Z(n568) );
  XOR U493 ( .A(n569), .B(n570), .Z(n560) );
  AND U494 ( .A(n571), .B(n572), .Z(n570) );
  XOR U495 ( .A(n426), .B(n569), .Z(n572) );
  XNOR U496 ( .A(p_input[229]), .B(n573), .Z(n426) );
  AND U497 ( .A(n89), .B(n574), .Z(n573) );
  XOR U498 ( .A(p_input[245]), .B(p_input[229]), .Z(n574) );
  XNOR U499 ( .A(n569), .B(n423), .Z(n571) );
  XOR U500 ( .A(n575), .B(n576), .Z(n423) );
  AND U501 ( .A(n87), .B(n577), .Z(n576) );
  XOR U502 ( .A(p_input[213]), .B(p_input[197]), .Z(n577) );
  XOR U503 ( .A(n578), .B(n579), .Z(n569) );
  AND U504 ( .A(n580), .B(n581), .Z(n579) );
  XOR U505 ( .A(n578), .B(n438), .Z(n581) );
  XNOR U506 ( .A(p_input[228]), .B(n582), .Z(n438) );
  AND U507 ( .A(n89), .B(n583), .Z(n582) );
  XOR U508 ( .A(p_input[244]), .B(p_input[228]), .Z(n583) );
  XNOR U509 ( .A(n435), .B(n578), .Z(n580) );
  XOR U510 ( .A(n584), .B(n585), .Z(n435) );
  AND U511 ( .A(n87), .B(n586), .Z(n585) );
  XOR U512 ( .A(p_input[212]), .B(p_input[196]), .Z(n586) );
  XOR U513 ( .A(n587), .B(n588), .Z(n578) );
  AND U514 ( .A(n589), .B(n590), .Z(n588) );
  XOR U515 ( .A(n587), .B(n450), .Z(n590) );
  XNOR U516 ( .A(p_input[227]), .B(n591), .Z(n450) );
  AND U517 ( .A(n89), .B(n592), .Z(n591) );
  XOR U518 ( .A(p_input[243]), .B(p_input[227]), .Z(n592) );
  XNOR U519 ( .A(n447), .B(n587), .Z(n589) );
  XOR U520 ( .A(n593), .B(n594), .Z(n447) );
  AND U521 ( .A(n87), .B(n595), .Z(n594) );
  XOR U522 ( .A(p_input[211]), .B(p_input[195]), .Z(n595) );
  XOR U523 ( .A(n596), .B(n597), .Z(n587) );
  AND U524 ( .A(n598), .B(n599), .Z(n597) );
  XOR U525 ( .A(n596), .B(n462), .Z(n599) );
  XNOR U526 ( .A(p_input[226]), .B(n600), .Z(n462) );
  AND U527 ( .A(n89), .B(n601), .Z(n600) );
  XOR U528 ( .A(p_input[242]), .B(p_input[226]), .Z(n601) );
  XNOR U529 ( .A(n459), .B(n596), .Z(n598) );
  XOR U530 ( .A(n602), .B(n603), .Z(n459) );
  AND U531 ( .A(n87), .B(n604), .Z(n603) );
  XOR U532 ( .A(p_input[210]), .B(p_input[194]), .Z(n604) );
  XOR U533 ( .A(n605), .B(n606), .Z(n596) );
  AND U534 ( .A(n607), .B(n608), .Z(n606) );
  XNOR U535 ( .A(n609), .B(n475), .Z(n608) );
  XNOR U536 ( .A(p_input[225]), .B(n610), .Z(n475) );
  AND U537 ( .A(n89), .B(n611), .Z(n610) );
  XNOR U538 ( .A(p_input[241]), .B(n612), .Z(n611) );
  IV U539 ( .A(p_input[225]), .Z(n612) );
  XNOR U540 ( .A(n472), .B(n605), .Z(n607) );
  XNOR U541 ( .A(p_input[193]), .B(n613), .Z(n472) );
  AND U542 ( .A(n87), .B(n614), .Z(n613) );
  XOR U543 ( .A(p_input[209]), .B(p_input[193]), .Z(n614) );
  IV U544 ( .A(n609), .Z(n605) );
  AND U545 ( .A(n480), .B(n483), .Z(n609) );
  XOR U546 ( .A(p_input[224]), .B(n615), .Z(n483) );
  AND U547 ( .A(n89), .B(n616), .Z(n615) );
  XOR U548 ( .A(p_input[240]), .B(p_input[224]), .Z(n616) );
  XOR U549 ( .A(n617), .B(n618), .Z(n89) );
  AND U550 ( .A(n619), .B(n620), .Z(n618) );
  XNOR U551 ( .A(p_input[255]), .B(n617), .Z(n620) );
  XOR U552 ( .A(n617), .B(p_input[239]), .Z(n619) );
  XOR U553 ( .A(n621), .B(n622), .Z(n617) );
  AND U554 ( .A(n623), .B(n624), .Z(n622) );
  XNOR U555 ( .A(p_input[254]), .B(n621), .Z(n624) );
  XOR U556 ( .A(n621), .B(p_input[238]), .Z(n623) );
  XOR U557 ( .A(n625), .B(n626), .Z(n621) );
  AND U558 ( .A(n627), .B(n628), .Z(n626) );
  XNOR U559 ( .A(p_input[253]), .B(n625), .Z(n628) );
  XOR U560 ( .A(n625), .B(p_input[237]), .Z(n627) );
  XOR U561 ( .A(n629), .B(n630), .Z(n625) );
  AND U562 ( .A(n631), .B(n632), .Z(n630) );
  XNOR U563 ( .A(p_input[252]), .B(n629), .Z(n632) );
  XOR U564 ( .A(n629), .B(p_input[236]), .Z(n631) );
  XOR U565 ( .A(n633), .B(n634), .Z(n629) );
  AND U566 ( .A(n635), .B(n636), .Z(n634) );
  XNOR U567 ( .A(p_input[251]), .B(n633), .Z(n636) );
  XOR U568 ( .A(n633), .B(p_input[235]), .Z(n635) );
  XOR U569 ( .A(n637), .B(n638), .Z(n633) );
  AND U570 ( .A(n639), .B(n640), .Z(n638) );
  XNOR U571 ( .A(p_input[250]), .B(n637), .Z(n640) );
  XOR U572 ( .A(n637), .B(p_input[234]), .Z(n639) );
  XOR U573 ( .A(n641), .B(n642), .Z(n637) );
  AND U574 ( .A(n643), .B(n644), .Z(n642) );
  XNOR U575 ( .A(p_input[249]), .B(n641), .Z(n644) );
  XOR U576 ( .A(n641), .B(p_input[233]), .Z(n643) );
  XOR U577 ( .A(n645), .B(n646), .Z(n641) );
  AND U578 ( .A(n647), .B(n648), .Z(n646) );
  XNOR U579 ( .A(p_input[248]), .B(n645), .Z(n648) );
  XOR U580 ( .A(n645), .B(p_input[232]), .Z(n647) );
  XOR U581 ( .A(n649), .B(n650), .Z(n645) );
  AND U582 ( .A(n651), .B(n652), .Z(n650) );
  XNOR U583 ( .A(p_input[247]), .B(n649), .Z(n652) );
  XOR U584 ( .A(n649), .B(p_input[231]), .Z(n651) );
  XOR U585 ( .A(n653), .B(n654), .Z(n649) );
  AND U586 ( .A(n655), .B(n656), .Z(n654) );
  XNOR U587 ( .A(p_input[246]), .B(n653), .Z(n656) );
  XOR U588 ( .A(n653), .B(p_input[230]), .Z(n655) );
  XOR U589 ( .A(n657), .B(n658), .Z(n653) );
  AND U590 ( .A(n659), .B(n660), .Z(n658) );
  XNOR U591 ( .A(p_input[245]), .B(n657), .Z(n660) );
  XOR U592 ( .A(n657), .B(p_input[229]), .Z(n659) );
  XOR U593 ( .A(n661), .B(n662), .Z(n657) );
  AND U594 ( .A(n663), .B(n664), .Z(n662) );
  XNOR U595 ( .A(p_input[244]), .B(n661), .Z(n664) );
  XOR U596 ( .A(n661), .B(p_input[228]), .Z(n663) );
  XOR U597 ( .A(n665), .B(n666), .Z(n661) );
  AND U598 ( .A(n667), .B(n668), .Z(n666) );
  XNOR U599 ( .A(p_input[243]), .B(n665), .Z(n668) );
  XOR U600 ( .A(n665), .B(p_input[227]), .Z(n667) );
  XOR U601 ( .A(n669), .B(n670), .Z(n665) );
  AND U602 ( .A(n671), .B(n672), .Z(n670) );
  XNOR U603 ( .A(p_input[242]), .B(n669), .Z(n672) );
  XOR U604 ( .A(n669), .B(p_input[226]), .Z(n671) );
  XNOR U605 ( .A(n673), .B(n674), .Z(n669) );
  AND U606 ( .A(n675), .B(n676), .Z(n674) );
  XOR U607 ( .A(p_input[241]), .B(n673), .Z(n676) );
  XNOR U608 ( .A(p_input[225]), .B(n673), .Z(n675) );
  AND U609 ( .A(p_input[240]), .B(n677), .Z(n673) );
  IV U610 ( .A(p_input[224]), .Z(n677) );
  XNOR U611 ( .A(p_input[192]), .B(n678), .Z(n480) );
  AND U612 ( .A(n87), .B(n679), .Z(n678) );
  XOR U613 ( .A(p_input[208]), .B(p_input[192]), .Z(n679) );
  XOR U614 ( .A(n680), .B(n681), .Z(n87) );
  AND U615 ( .A(n682), .B(n683), .Z(n681) );
  XNOR U616 ( .A(p_input[223]), .B(n680), .Z(n683) );
  XOR U617 ( .A(n680), .B(p_input[207]), .Z(n682) );
  XOR U618 ( .A(n684), .B(n685), .Z(n680) );
  AND U619 ( .A(n686), .B(n687), .Z(n685) );
  XNOR U620 ( .A(p_input[222]), .B(n684), .Z(n687) );
  XNOR U621 ( .A(n684), .B(n494), .Z(n686) );
  IV U622 ( .A(p_input[206]), .Z(n494) );
  XOR U623 ( .A(n688), .B(n689), .Z(n684) );
  AND U624 ( .A(n690), .B(n691), .Z(n689) );
  XNOR U625 ( .A(p_input[221]), .B(n688), .Z(n691) );
  XNOR U626 ( .A(n688), .B(n503), .Z(n690) );
  IV U627 ( .A(p_input[205]), .Z(n503) );
  XOR U628 ( .A(n692), .B(n693), .Z(n688) );
  AND U629 ( .A(n694), .B(n695), .Z(n693) );
  XNOR U630 ( .A(p_input[220]), .B(n692), .Z(n695) );
  XNOR U631 ( .A(n692), .B(n512), .Z(n694) );
  IV U632 ( .A(p_input[204]), .Z(n512) );
  XOR U633 ( .A(n696), .B(n697), .Z(n692) );
  AND U634 ( .A(n698), .B(n699), .Z(n697) );
  XNOR U635 ( .A(p_input[219]), .B(n696), .Z(n699) );
  XNOR U636 ( .A(n696), .B(n521), .Z(n698) );
  IV U637 ( .A(p_input[203]), .Z(n521) );
  XOR U638 ( .A(n700), .B(n701), .Z(n696) );
  AND U639 ( .A(n702), .B(n703), .Z(n701) );
  XNOR U640 ( .A(p_input[218]), .B(n700), .Z(n703) );
  XNOR U641 ( .A(n700), .B(n530), .Z(n702) );
  IV U642 ( .A(p_input[202]), .Z(n530) );
  XOR U643 ( .A(n704), .B(n705), .Z(n700) );
  AND U644 ( .A(n706), .B(n707), .Z(n705) );
  XNOR U645 ( .A(p_input[217]), .B(n704), .Z(n707) );
  XNOR U646 ( .A(n704), .B(n539), .Z(n706) );
  IV U647 ( .A(p_input[201]), .Z(n539) );
  XOR U648 ( .A(n708), .B(n709), .Z(n704) );
  AND U649 ( .A(n710), .B(n711), .Z(n709) );
  XNOR U650 ( .A(p_input[216]), .B(n708), .Z(n711) );
  XNOR U651 ( .A(n708), .B(n548), .Z(n710) );
  IV U652 ( .A(p_input[200]), .Z(n548) );
  XOR U653 ( .A(n712), .B(n713), .Z(n708) );
  AND U654 ( .A(n714), .B(n715), .Z(n713) );
  XNOR U655 ( .A(p_input[215]), .B(n712), .Z(n715) );
  XNOR U656 ( .A(n712), .B(n557), .Z(n714) );
  IV U657 ( .A(p_input[199]), .Z(n557) );
  XOR U658 ( .A(n716), .B(n717), .Z(n712) );
  AND U659 ( .A(n718), .B(n719), .Z(n717) );
  XNOR U660 ( .A(p_input[214]), .B(n716), .Z(n719) );
  XNOR U661 ( .A(n716), .B(n566), .Z(n718) );
  IV U662 ( .A(p_input[198]), .Z(n566) );
  XOR U663 ( .A(n720), .B(n721), .Z(n716) );
  AND U664 ( .A(n722), .B(n723), .Z(n721) );
  XNOR U665 ( .A(p_input[213]), .B(n720), .Z(n723) );
  XNOR U666 ( .A(n720), .B(n575), .Z(n722) );
  IV U667 ( .A(p_input[197]), .Z(n575) );
  XOR U668 ( .A(n724), .B(n725), .Z(n720) );
  AND U669 ( .A(n726), .B(n727), .Z(n725) );
  XNOR U670 ( .A(p_input[212]), .B(n724), .Z(n727) );
  XNOR U671 ( .A(n724), .B(n584), .Z(n726) );
  IV U672 ( .A(p_input[196]), .Z(n584) );
  XOR U673 ( .A(n728), .B(n729), .Z(n724) );
  AND U674 ( .A(n730), .B(n731), .Z(n729) );
  XNOR U675 ( .A(p_input[211]), .B(n728), .Z(n731) );
  XNOR U676 ( .A(n728), .B(n593), .Z(n730) );
  IV U677 ( .A(p_input[195]), .Z(n593) );
  XOR U678 ( .A(n732), .B(n733), .Z(n728) );
  AND U679 ( .A(n734), .B(n735), .Z(n733) );
  XNOR U680 ( .A(p_input[210]), .B(n732), .Z(n735) );
  XNOR U681 ( .A(n732), .B(n602), .Z(n734) );
  IV U682 ( .A(p_input[194]), .Z(n602) );
  XNOR U683 ( .A(n736), .B(n737), .Z(n732) );
  AND U684 ( .A(n738), .B(n739), .Z(n737) );
  XOR U685 ( .A(p_input[209]), .B(n736), .Z(n739) );
  XNOR U686 ( .A(p_input[193]), .B(n736), .Z(n738) );
  AND U687 ( .A(p_input[208]), .B(n740), .Z(n736) );
  IV U688 ( .A(p_input[192]), .Z(n740) );
  XOR U689 ( .A(n741), .B(n742), .Z(n299) );
  AND U690 ( .A(n99), .B(n743), .Z(n742) );
  XNOR U691 ( .A(n744), .B(n741), .Z(n743) );
  XOR U692 ( .A(n745), .B(n746), .Z(n99) );
  AND U693 ( .A(n747), .B(n748), .Z(n746) );
  XNOR U694 ( .A(n309), .B(n745), .Z(n748) );
  AND U695 ( .A(p_input[191]), .B(p_input[175]), .Z(n309) );
  XOR U696 ( .A(n745), .B(n310), .Z(n747) );
  AND U697 ( .A(p_input[159]), .B(p_input[143]), .Z(n310) );
  XOR U698 ( .A(n749), .B(n750), .Z(n745) );
  AND U699 ( .A(n751), .B(n752), .Z(n750) );
  XOR U700 ( .A(n749), .B(n322), .Z(n752) );
  XNOR U701 ( .A(p_input[174]), .B(n753), .Z(n322) );
  AND U702 ( .A(n93), .B(n754), .Z(n753) );
  XOR U703 ( .A(p_input[190]), .B(p_input[174]), .Z(n754) );
  XNOR U704 ( .A(n319), .B(n749), .Z(n751) );
  XOR U705 ( .A(n755), .B(n756), .Z(n319) );
  AND U706 ( .A(n90), .B(n757), .Z(n756) );
  XOR U707 ( .A(p_input[158]), .B(p_input[142]), .Z(n757) );
  XOR U708 ( .A(n758), .B(n759), .Z(n749) );
  AND U709 ( .A(n760), .B(n761), .Z(n759) );
  XOR U710 ( .A(n758), .B(n334), .Z(n761) );
  XNOR U711 ( .A(p_input[173]), .B(n762), .Z(n334) );
  AND U712 ( .A(n93), .B(n763), .Z(n762) );
  XOR U713 ( .A(p_input[189]), .B(p_input[173]), .Z(n763) );
  XNOR U714 ( .A(n331), .B(n758), .Z(n760) );
  XOR U715 ( .A(n764), .B(n765), .Z(n331) );
  AND U716 ( .A(n90), .B(n766), .Z(n765) );
  XOR U717 ( .A(p_input[157]), .B(p_input[141]), .Z(n766) );
  XOR U718 ( .A(n767), .B(n768), .Z(n758) );
  AND U719 ( .A(n769), .B(n770), .Z(n768) );
  XOR U720 ( .A(n767), .B(n346), .Z(n770) );
  XNOR U721 ( .A(p_input[172]), .B(n771), .Z(n346) );
  AND U722 ( .A(n93), .B(n772), .Z(n771) );
  XOR U723 ( .A(p_input[188]), .B(p_input[172]), .Z(n772) );
  XNOR U724 ( .A(n343), .B(n767), .Z(n769) );
  XOR U725 ( .A(n773), .B(n774), .Z(n343) );
  AND U726 ( .A(n90), .B(n775), .Z(n774) );
  XOR U727 ( .A(p_input[156]), .B(p_input[140]), .Z(n775) );
  XOR U728 ( .A(n776), .B(n777), .Z(n767) );
  AND U729 ( .A(n778), .B(n779), .Z(n777) );
  XOR U730 ( .A(n776), .B(n358), .Z(n779) );
  XNOR U731 ( .A(p_input[171]), .B(n780), .Z(n358) );
  AND U732 ( .A(n93), .B(n781), .Z(n780) );
  XOR U733 ( .A(p_input[187]), .B(p_input[171]), .Z(n781) );
  XNOR U734 ( .A(n355), .B(n776), .Z(n778) );
  XOR U735 ( .A(n782), .B(n783), .Z(n355) );
  AND U736 ( .A(n90), .B(n784), .Z(n783) );
  XOR U737 ( .A(p_input[155]), .B(p_input[139]), .Z(n784) );
  XOR U738 ( .A(n785), .B(n786), .Z(n776) );
  AND U739 ( .A(n787), .B(n788), .Z(n786) );
  XOR U740 ( .A(n785), .B(n370), .Z(n788) );
  XNOR U741 ( .A(p_input[170]), .B(n789), .Z(n370) );
  AND U742 ( .A(n93), .B(n790), .Z(n789) );
  XOR U743 ( .A(p_input[186]), .B(p_input[170]), .Z(n790) );
  XNOR U744 ( .A(n367), .B(n785), .Z(n787) );
  XOR U745 ( .A(n791), .B(n792), .Z(n367) );
  AND U746 ( .A(n90), .B(n793), .Z(n792) );
  XOR U747 ( .A(p_input[154]), .B(p_input[138]), .Z(n793) );
  XOR U748 ( .A(n794), .B(n795), .Z(n785) );
  AND U749 ( .A(n796), .B(n797), .Z(n795) );
  XOR U750 ( .A(n794), .B(n382), .Z(n797) );
  XNOR U751 ( .A(p_input[169]), .B(n798), .Z(n382) );
  AND U752 ( .A(n93), .B(n799), .Z(n798) );
  XOR U753 ( .A(p_input[185]), .B(p_input[169]), .Z(n799) );
  XNOR U754 ( .A(n379), .B(n794), .Z(n796) );
  XOR U755 ( .A(n800), .B(n801), .Z(n379) );
  AND U756 ( .A(n90), .B(n802), .Z(n801) );
  XOR U757 ( .A(p_input[153]), .B(p_input[137]), .Z(n802) );
  XOR U758 ( .A(n803), .B(n804), .Z(n794) );
  AND U759 ( .A(n805), .B(n806), .Z(n804) );
  XOR U760 ( .A(n803), .B(n394), .Z(n806) );
  XNOR U761 ( .A(p_input[168]), .B(n807), .Z(n394) );
  AND U762 ( .A(n93), .B(n808), .Z(n807) );
  XOR U763 ( .A(p_input[184]), .B(p_input[168]), .Z(n808) );
  XNOR U764 ( .A(n391), .B(n803), .Z(n805) );
  XOR U765 ( .A(n809), .B(n810), .Z(n391) );
  AND U766 ( .A(n90), .B(n811), .Z(n810) );
  XOR U767 ( .A(p_input[152]), .B(p_input[136]), .Z(n811) );
  XOR U768 ( .A(n812), .B(n813), .Z(n803) );
  AND U769 ( .A(n814), .B(n815), .Z(n813) );
  XOR U770 ( .A(n812), .B(n406), .Z(n815) );
  XNOR U771 ( .A(p_input[167]), .B(n816), .Z(n406) );
  AND U772 ( .A(n93), .B(n817), .Z(n816) );
  XOR U773 ( .A(p_input[183]), .B(p_input[167]), .Z(n817) );
  XNOR U774 ( .A(n403), .B(n812), .Z(n814) );
  XOR U775 ( .A(n818), .B(n819), .Z(n403) );
  AND U776 ( .A(n90), .B(n820), .Z(n819) );
  XOR U777 ( .A(p_input[151]), .B(p_input[135]), .Z(n820) );
  XOR U778 ( .A(n821), .B(n822), .Z(n812) );
  AND U779 ( .A(n823), .B(n824), .Z(n822) );
  XOR U780 ( .A(n821), .B(n418), .Z(n824) );
  XNOR U781 ( .A(p_input[166]), .B(n825), .Z(n418) );
  AND U782 ( .A(n93), .B(n826), .Z(n825) );
  XOR U783 ( .A(p_input[182]), .B(p_input[166]), .Z(n826) );
  XNOR U784 ( .A(n415), .B(n821), .Z(n823) );
  XOR U785 ( .A(n827), .B(n828), .Z(n415) );
  AND U786 ( .A(n90), .B(n829), .Z(n828) );
  XOR U787 ( .A(p_input[150]), .B(p_input[134]), .Z(n829) );
  XOR U788 ( .A(n830), .B(n831), .Z(n821) );
  AND U789 ( .A(n832), .B(n833), .Z(n831) );
  XOR U790 ( .A(n430), .B(n830), .Z(n833) );
  XNOR U791 ( .A(p_input[165]), .B(n834), .Z(n430) );
  AND U792 ( .A(n93), .B(n835), .Z(n834) );
  XOR U793 ( .A(p_input[181]), .B(p_input[165]), .Z(n835) );
  XNOR U794 ( .A(n830), .B(n427), .Z(n832) );
  XOR U795 ( .A(n836), .B(n837), .Z(n427) );
  AND U796 ( .A(n90), .B(n838), .Z(n837) );
  XOR U797 ( .A(p_input[149]), .B(p_input[133]), .Z(n838) );
  XOR U798 ( .A(n839), .B(n840), .Z(n830) );
  AND U799 ( .A(n841), .B(n842), .Z(n840) );
  XOR U800 ( .A(n839), .B(n442), .Z(n842) );
  XNOR U801 ( .A(p_input[164]), .B(n843), .Z(n442) );
  AND U802 ( .A(n93), .B(n844), .Z(n843) );
  XOR U803 ( .A(p_input[180]), .B(p_input[164]), .Z(n844) );
  XNOR U804 ( .A(n439), .B(n839), .Z(n841) );
  XOR U805 ( .A(n845), .B(n846), .Z(n439) );
  AND U806 ( .A(n90), .B(n847), .Z(n846) );
  XOR U807 ( .A(p_input[148]), .B(p_input[132]), .Z(n847) );
  XOR U808 ( .A(n848), .B(n849), .Z(n839) );
  AND U809 ( .A(n850), .B(n851), .Z(n849) );
  XOR U810 ( .A(n848), .B(n454), .Z(n851) );
  XNOR U811 ( .A(p_input[163]), .B(n852), .Z(n454) );
  AND U812 ( .A(n93), .B(n853), .Z(n852) );
  XOR U813 ( .A(p_input[179]), .B(p_input[163]), .Z(n853) );
  XNOR U814 ( .A(n451), .B(n848), .Z(n850) );
  XOR U815 ( .A(n854), .B(n855), .Z(n451) );
  AND U816 ( .A(n90), .B(n856), .Z(n855) );
  XOR U817 ( .A(p_input[147]), .B(p_input[131]), .Z(n856) );
  XOR U818 ( .A(n857), .B(n858), .Z(n848) );
  AND U819 ( .A(n859), .B(n860), .Z(n858) );
  XOR U820 ( .A(n857), .B(n466), .Z(n860) );
  XNOR U821 ( .A(p_input[162]), .B(n861), .Z(n466) );
  AND U822 ( .A(n93), .B(n862), .Z(n861) );
  XOR U823 ( .A(p_input[178]), .B(p_input[162]), .Z(n862) );
  XNOR U824 ( .A(n463), .B(n857), .Z(n859) );
  XOR U825 ( .A(n863), .B(n864), .Z(n463) );
  AND U826 ( .A(n90), .B(n865), .Z(n864) );
  XOR U827 ( .A(p_input[146]), .B(p_input[130]), .Z(n865) );
  XOR U828 ( .A(n866), .B(n867), .Z(n857) );
  AND U829 ( .A(n868), .B(n869), .Z(n867) );
  XNOR U830 ( .A(n870), .B(n479), .Z(n869) );
  XNOR U831 ( .A(p_input[161]), .B(n871), .Z(n479) );
  AND U832 ( .A(n93), .B(n872), .Z(n871) );
  XNOR U833 ( .A(p_input[177]), .B(n873), .Z(n872) );
  IV U834 ( .A(p_input[161]), .Z(n873) );
  XNOR U835 ( .A(n476), .B(n866), .Z(n868) );
  XNOR U836 ( .A(p_input[129]), .B(n874), .Z(n476) );
  AND U837 ( .A(n90), .B(n875), .Z(n874) );
  XOR U838 ( .A(p_input[145]), .B(p_input[129]), .Z(n875) );
  IV U839 ( .A(n870), .Z(n866) );
  AND U840 ( .A(n741), .B(n744), .Z(n870) );
  XOR U841 ( .A(p_input[160]), .B(n876), .Z(n744) );
  AND U842 ( .A(n93), .B(n877), .Z(n876) );
  XOR U843 ( .A(p_input[176]), .B(p_input[160]), .Z(n877) );
  XOR U844 ( .A(n878), .B(n879), .Z(n93) );
  AND U845 ( .A(n880), .B(n881), .Z(n879) );
  XNOR U846 ( .A(p_input[191]), .B(n878), .Z(n881) );
  XOR U847 ( .A(n878), .B(p_input[175]), .Z(n880) );
  XOR U848 ( .A(n882), .B(n883), .Z(n878) );
  AND U849 ( .A(n884), .B(n885), .Z(n883) );
  XNOR U850 ( .A(p_input[190]), .B(n882), .Z(n885) );
  XOR U851 ( .A(n882), .B(p_input[174]), .Z(n884) );
  XOR U852 ( .A(n886), .B(n887), .Z(n882) );
  AND U853 ( .A(n888), .B(n889), .Z(n887) );
  XNOR U854 ( .A(p_input[189]), .B(n886), .Z(n889) );
  XOR U855 ( .A(n886), .B(p_input[173]), .Z(n888) );
  XOR U856 ( .A(n890), .B(n891), .Z(n886) );
  AND U857 ( .A(n892), .B(n893), .Z(n891) );
  XNOR U858 ( .A(p_input[188]), .B(n890), .Z(n893) );
  XOR U859 ( .A(n890), .B(p_input[172]), .Z(n892) );
  XOR U860 ( .A(n894), .B(n895), .Z(n890) );
  AND U861 ( .A(n896), .B(n897), .Z(n895) );
  XNOR U862 ( .A(p_input[187]), .B(n894), .Z(n897) );
  XOR U863 ( .A(n894), .B(p_input[171]), .Z(n896) );
  XOR U864 ( .A(n898), .B(n899), .Z(n894) );
  AND U865 ( .A(n900), .B(n901), .Z(n899) );
  XNOR U866 ( .A(p_input[186]), .B(n898), .Z(n901) );
  XOR U867 ( .A(n898), .B(p_input[170]), .Z(n900) );
  XOR U868 ( .A(n902), .B(n903), .Z(n898) );
  AND U869 ( .A(n904), .B(n905), .Z(n903) );
  XNOR U870 ( .A(p_input[185]), .B(n902), .Z(n905) );
  XOR U871 ( .A(n902), .B(p_input[169]), .Z(n904) );
  XOR U872 ( .A(n906), .B(n907), .Z(n902) );
  AND U873 ( .A(n908), .B(n909), .Z(n907) );
  XNOR U874 ( .A(p_input[184]), .B(n906), .Z(n909) );
  XOR U875 ( .A(n906), .B(p_input[168]), .Z(n908) );
  XOR U876 ( .A(n910), .B(n911), .Z(n906) );
  AND U877 ( .A(n912), .B(n913), .Z(n911) );
  XNOR U878 ( .A(p_input[183]), .B(n910), .Z(n913) );
  XOR U879 ( .A(n910), .B(p_input[167]), .Z(n912) );
  XOR U880 ( .A(n914), .B(n915), .Z(n910) );
  AND U881 ( .A(n916), .B(n917), .Z(n915) );
  XNOR U882 ( .A(p_input[182]), .B(n914), .Z(n917) );
  XOR U883 ( .A(n914), .B(p_input[166]), .Z(n916) );
  XOR U884 ( .A(n918), .B(n919), .Z(n914) );
  AND U885 ( .A(n920), .B(n921), .Z(n919) );
  XNOR U886 ( .A(p_input[181]), .B(n918), .Z(n921) );
  XOR U887 ( .A(n918), .B(p_input[165]), .Z(n920) );
  XOR U888 ( .A(n922), .B(n923), .Z(n918) );
  AND U889 ( .A(n924), .B(n925), .Z(n923) );
  XNOR U890 ( .A(p_input[180]), .B(n922), .Z(n925) );
  XOR U891 ( .A(n922), .B(p_input[164]), .Z(n924) );
  XOR U892 ( .A(n926), .B(n927), .Z(n922) );
  AND U893 ( .A(n928), .B(n929), .Z(n927) );
  XNOR U894 ( .A(p_input[179]), .B(n926), .Z(n929) );
  XOR U895 ( .A(n926), .B(p_input[163]), .Z(n928) );
  XOR U896 ( .A(n930), .B(n931), .Z(n926) );
  AND U897 ( .A(n932), .B(n933), .Z(n931) );
  XNOR U898 ( .A(p_input[178]), .B(n930), .Z(n933) );
  XOR U899 ( .A(n930), .B(p_input[162]), .Z(n932) );
  XNOR U900 ( .A(n934), .B(n935), .Z(n930) );
  AND U901 ( .A(n936), .B(n937), .Z(n935) );
  XOR U902 ( .A(p_input[177]), .B(n934), .Z(n937) );
  XNOR U903 ( .A(p_input[161]), .B(n934), .Z(n936) );
  AND U904 ( .A(p_input[176]), .B(n938), .Z(n934) );
  IV U905 ( .A(p_input[160]), .Z(n938) );
  XNOR U906 ( .A(p_input[128]), .B(n939), .Z(n741) );
  AND U907 ( .A(n90), .B(n940), .Z(n939) );
  XOR U908 ( .A(p_input[144]), .B(p_input[128]), .Z(n940) );
  XOR U909 ( .A(n941), .B(n942), .Z(n90) );
  AND U910 ( .A(n943), .B(n944), .Z(n942) );
  XNOR U911 ( .A(p_input[159]), .B(n941), .Z(n944) );
  XOR U912 ( .A(n941), .B(p_input[143]), .Z(n943) );
  XOR U913 ( .A(n945), .B(n946), .Z(n941) );
  AND U914 ( .A(n947), .B(n948), .Z(n946) );
  XNOR U915 ( .A(p_input[158]), .B(n945), .Z(n948) );
  XNOR U916 ( .A(n945), .B(n755), .Z(n947) );
  IV U917 ( .A(p_input[142]), .Z(n755) );
  XOR U918 ( .A(n949), .B(n950), .Z(n945) );
  AND U919 ( .A(n951), .B(n952), .Z(n950) );
  XNOR U920 ( .A(p_input[157]), .B(n949), .Z(n952) );
  XNOR U921 ( .A(n949), .B(n764), .Z(n951) );
  IV U922 ( .A(p_input[141]), .Z(n764) );
  XOR U923 ( .A(n953), .B(n954), .Z(n949) );
  AND U924 ( .A(n955), .B(n956), .Z(n954) );
  XNOR U925 ( .A(p_input[156]), .B(n953), .Z(n956) );
  XNOR U926 ( .A(n953), .B(n773), .Z(n955) );
  IV U927 ( .A(p_input[140]), .Z(n773) );
  XOR U928 ( .A(n957), .B(n958), .Z(n953) );
  AND U929 ( .A(n959), .B(n960), .Z(n958) );
  XNOR U930 ( .A(p_input[155]), .B(n957), .Z(n960) );
  XNOR U931 ( .A(n957), .B(n782), .Z(n959) );
  IV U932 ( .A(p_input[139]), .Z(n782) );
  XOR U933 ( .A(n961), .B(n962), .Z(n957) );
  AND U934 ( .A(n963), .B(n964), .Z(n962) );
  XNOR U935 ( .A(p_input[154]), .B(n961), .Z(n964) );
  XNOR U936 ( .A(n961), .B(n791), .Z(n963) );
  IV U937 ( .A(p_input[138]), .Z(n791) );
  XOR U938 ( .A(n965), .B(n966), .Z(n961) );
  AND U939 ( .A(n967), .B(n968), .Z(n966) );
  XNOR U940 ( .A(p_input[153]), .B(n965), .Z(n968) );
  XNOR U941 ( .A(n965), .B(n800), .Z(n967) );
  IV U942 ( .A(p_input[137]), .Z(n800) );
  XOR U943 ( .A(n969), .B(n970), .Z(n965) );
  AND U944 ( .A(n971), .B(n972), .Z(n970) );
  XNOR U945 ( .A(p_input[152]), .B(n969), .Z(n972) );
  XNOR U946 ( .A(n969), .B(n809), .Z(n971) );
  IV U947 ( .A(p_input[136]), .Z(n809) );
  XOR U948 ( .A(n973), .B(n974), .Z(n969) );
  AND U949 ( .A(n975), .B(n976), .Z(n974) );
  XNOR U950 ( .A(p_input[151]), .B(n973), .Z(n976) );
  XNOR U951 ( .A(n973), .B(n818), .Z(n975) );
  IV U952 ( .A(p_input[135]), .Z(n818) );
  XOR U953 ( .A(n977), .B(n978), .Z(n973) );
  AND U954 ( .A(n979), .B(n980), .Z(n978) );
  XNOR U955 ( .A(p_input[150]), .B(n977), .Z(n980) );
  XNOR U956 ( .A(n977), .B(n827), .Z(n979) );
  IV U957 ( .A(p_input[134]), .Z(n827) );
  XOR U958 ( .A(n981), .B(n982), .Z(n977) );
  AND U959 ( .A(n983), .B(n984), .Z(n982) );
  XNOR U960 ( .A(p_input[149]), .B(n981), .Z(n984) );
  XNOR U961 ( .A(n981), .B(n836), .Z(n983) );
  IV U962 ( .A(p_input[133]), .Z(n836) );
  XOR U963 ( .A(n985), .B(n986), .Z(n981) );
  AND U964 ( .A(n987), .B(n988), .Z(n986) );
  XNOR U965 ( .A(p_input[148]), .B(n985), .Z(n988) );
  XNOR U966 ( .A(n985), .B(n845), .Z(n987) );
  IV U967 ( .A(p_input[132]), .Z(n845) );
  XOR U968 ( .A(n989), .B(n990), .Z(n985) );
  AND U969 ( .A(n991), .B(n992), .Z(n990) );
  XNOR U970 ( .A(p_input[147]), .B(n989), .Z(n992) );
  XNOR U971 ( .A(n989), .B(n854), .Z(n991) );
  IV U972 ( .A(p_input[131]), .Z(n854) );
  XOR U973 ( .A(n993), .B(n994), .Z(n989) );
  AND U974 ( .A(n995), .B(n996), .Z(n994) );
  XNOR U975 ( .A(p_input[146]), .B(n993), .Z(n996) );
  XNOR U976 ( .A(n993), .B(n863), .Z(n995) );
  IV U977 ( .A(p_input[130]), .Z(n863) );
  XNOR U978 ( .A(n997), .B(n998), .Z(n993) );
  AND U979 ( .A(n999), .B(n1000), .Z(n998) );
  XOR U980 ( .A(p_input[145]), .B(n997), .Z(n1000) );
  XNOR U981 ( .A(p_input[129]), .B(n997), .Z(n999) );
  AND U982 ( .A(p_input[144]), .B(n1001), .Z(n997) );
  IV U983 ( .A(p_input[128]), .Z(n1001) );
  XOR U984 ( .A(n1002), .B(n1003), .Z(n26) );
  AND U985 ( .A(n114), .B(n1004), .Z(n1003) );
  XNOR U986 ( .A(n1005), .B(n1002), .Z(n1004) );
  XOR U987 ( .A(n1006), .B(n1007), .Z(n114) );
  AND U988 ( .A(n1008), .B(n1009), .Z(n1007) );
  XNOR U989 ( .A(n130), .B(n1006), .Z(n1009) );
  AND U990 ( .A(n1010), .B(n1011), .Z(n130) );
  XOR U991 ( .A(n1006), .B(n129), .Z(n1008) );
  AND U992 ( .A(n1012), .B(n1013), .Z(n129) );
  XOR U993 ( .A(n1014), .B(n1015), .Z(n1006) );
  AND U994 ( .A(n1016), .B(n1017), .Z(n1015) );
  XOR U995 ( .A(n1014), .B(n142), .Z(n1017) );
  XOR U996 ( .A(n1018), .B(n1019), .Z(n142) );
  AND U997 ( .A(n105), .B(n1020), .Z(n1019) );
  XOR U998 ( .A(n1021), .B(n1018), .Z(n1020) );
  XNOR U999 ( .A(n139), .B(n1014), .Z(n1016) );
  XOR U1000 ( .A(n1022), .B(n1023), .Z(n139) );
  AND U1001 ( .A(n102), .B(n1024), .Z(n1023) );
  XOR U1002 ( .A(n1025), .B(n1022), .Z(n1024) );
  XOR U1003 ( .A(n1026), .B(n1027), .Z(n1014) );
  AND U1004 ( .A(n1028), .B(n1029), .Z(n1027) );
  XOR U1005 ( .A(n1026), .B(n154), .Z(n1029) );
  XOR U1006 ( .A(n1030), .B(n1031), .Z(n154) );
  AND U1007 ( .A(n105), .B(n1032), .Z(n1031) );
  XOR U1008 ( .A(n1033), .B(n1030), .Z(n1032) );
  XNOR U1009 ( .A(n151), .B(n1026), .Z(n1028) );
  XOR U1010 ( .A(n1034), .B(n1035), .Z(n151) );
  AND U1011 ( .A(n102), .B(n1036), .Z(n1035) );
  XOR U1012 ( .A(n1037), .B(n1034), .Z(n1036) );
  XOR U1013 ( .A(n1038), .B(n1039), .Z(n1026) );
  AND U1014 ( .A(n1040), .B(n1041), .Z(n1039) );
  XOR U1015 ( .A(n1038), .B(n166), .Z(n1041) );
  XOR U1016 ( .A(n1042), .B(n1043), .Z(n166) );
  AND U1017 ( .A(n105), .B(n1044), .Z(n1043) );
  XOR U1018 ( .A(n1045), .B(n1042), .Z(n1044) );
  XNOR U1019 ( .A(n163), .B(n1038), .Z(n1040) );
  XOR U1020 ( .A(n1046), .B(n1047), .Z(n163) );
  AND U1021 ( .A(n102), .B(n1048), .Z(n1047) );
  XOR U1022 ( .A(n1049), .B(n1046), .Z(n1048) );
  XOR U1023 ( .A(n1050), .B(n1051), .Z(n1038) );
  AND U1024 ( .A(n1052), .B(n1053), .Z(n1051) );
  XOR U1025 ( .A(n1050), .B(n178), .Z(n1053) );
  XOR U1026 ( .A(n1054), .B(n1055), .Z(n178) );
  AND U1027 ( .A(n105), .B(n1056), .Z(n1055) );
  XOR U1028 ( .A(n1057), .B(n1054), .Z(n1056) );
  XNOR U1029 ( .A(n175), .B(n1050), .Z(n1052) );
  XOR U1030 ( .A(n1058), .B(n1059), .Z(n175) );
  AND U1031 ( .A(n102), .B(n1060), .Z(n1059) );
  XOR U1032 ( .A(n1061), .B(n1058), .Z(n1060) );
  XOR U1033 ( .A(n1062), .B(n1063), .Z(n1050) );
  AND U1034 ( .A(n1064), .B(n1065), .Z(n1063) );
  XOR U1035 ( .A(n1062), .B(n190), .Z(n1065) );
  XOR U1036 ( .A(n1066), .B(n1067), .Z(n190) );
  AND U1037 ( .A(n105), .B(n1068), .Z(n1067) );
  XOR U1038 ( .A(n1069), .B(n1066), .Z(n1068) );
  XNOR U1039 ( .A(n187), .B(n1062), .Z(n1064) );
  XOR U1040 ( .A(n1070), .B(n1071), .Z(n187) );
  AND U1041 ( .A(n102), .B(n1072), .Z(n1071) );
  XOR U1042 ( .A(n1073), .B(n1070), .Z(n1072) );
  XOR U1043 ( .A(n1074), .B(n1075), .Z(n1062) );
  AND U1044 ( .A(n1076), .B(n1077), .Z(n1075) );
  XOR U1045 ( .A(n1074), .B(n202), .Z(n1077) );
  XOR U1046 ( .A(n1078), .B(n1079), .Z(n202) );
  AND U1047 ( .A(n105), .B(n1080), .Z(n1079) );
  XOR U1048 ( .A(n1081), .B(n1078), .Z(n1080) );
  XNOR U1049 ( .A(n199), .B(n1074), .Z(n1076) );
  XOR U1050 ( .A(n1082), .B(n1083), .Z(n199) );
  AND U1051 ( .A(n102), .B(n1084), .Z(n1083) );
  XOR U1052 ( .A(n1085), .B(n1082), .Z(n1084) );
  XOR U1053 ( .A(n1086), .B(n1087), .Z(n1074) );
  AND U1054 ( .A(n1088), .B(n1089), .Z(n1087) );
  XOR U1055 ( .A(n1086), .B(n214), .Z(n1089) );
  XOR U1056 ( .A(n1090), .B(n1091), .Z(n214) );
  AND U1057 ( .A(n105), .B(n1092), .Z(n1091) );
  XOR U1058 ( .A(n1093), .B(n1090), .Z(n1092) );
  XNOR U1059 ( .A(n211), .B(n1086), .Z(n1088) );
  XOR U1060 ( .A(n1094), .B(n1095), .Z(n211) );
  AND U1061 ( .A(n102), .B(n1096), .Z(n1095) );
  XOR U1062 ( .A(n1097), .B(n1094), .Z(n1096) );
  XOR U1063 ( .A(n1098), .B(n1099), .Z(n1086) );
  AND U1064 ( .A(n1100), .B(n1101), .Z(n1099) );
  XOR U1065 ( .A(n1098), .B(n226), .Z(n1101) );
  XOR U1066 ( .A(n1102), .B(n1103), .Z(n226) );
  AND U1067 ( .A(n105), .B(n1104), .Z(n1103) );
  XOR U1068 ( .A(n1105), .B(n1102), .Z(n1104) );
  XNOR U1069 ( .A(n223), .B(n1098), .Z(n1100) );
  XOR U1070 ( .A(n1106), .B(n1107), .Z(n223) );
  AND U1071 ( .A(n102), .B(n1108), .Z(n1107) );
  XOR U1072 ( .A(n1109), .B(n1106), .Z(n1108) );
  XOR U1073 ( .A(n1110), .B(n1111), .Z(n1098) );
  AND U1074 ( .A(n1112), .B(n1113), .Z(n1111) );
  XOR U1075 ( .A(n1110), .B(n238), .Z(n1113) );
  XOR U1076 ( .A(n1114), .B(n1115), .Z(n238) );
  AND U1077 ( .A(n105), .B(n1116), .Z(n1115) );
  XOR U1078 ( .A(n1117), .B(n1114), .Z(n1116) );
  XNOR U1079 ( .A(n235), .B(n1110), .Z(n1112) );
  XOR U1080 ( .A(n1118), .B(n1119), .Z(n235) );
  AND U1081 ( .A(n102), .B(n1120), .Z(n1119) );
  XOR U1082 ( .A(n1121), .B(n1118), .Z(n1120) );
  XOR U1083 ( .A(n1122), .B(n1123), .Z(n1110) );
  AND U1084 ( .A(n1124), .B(n1125), .Z(n1123) );
  XOR U1085 ( .A(n250), .B(n1122), .Z(n1125) );
  XOR U1086 ( .A(n1126), .B(n1127), .Z(n250) );
  AND U1087 ( .A(n105), .B(n1128), .Z(n1127) );
  XOR U1088 ( .A(n1126), .B(n1129), .Z(n1128) );
  XNOR U1089 ( .A(n1122), .B(n247), .Z(n1124) );
  XOR U1090 ( .A(n1130), .B(n1131), .Z(n247) );
  AND U1091 ( .A(n102), .B(n1132), .Z(n1131) );
  XOR U1092 ( .A(n1130), .B(n1133), .Z(n1132) );
  XOR U1093 ( .A(n1134), .B(n1135), .Z(n1122) );
  AND U1094 ( .A(n1136), .B(n1137), .Z(n1135) );
  XOR U1095 ( .A(n1134), .B(n262), .Z(n1137) );
  XOR U1096 ( .A(n1138), .B(n1139), .Z(n262) );
  AND U1097 ( .A(n105), .B(n1140), .Z(n1139) );
  XOR U1098 ( .A(n1141), .B(n1138), .Z(n1140) );
  XNOR U1099 ( .A(n259), .B(n1134), .Z(n1136) );
  XOR U1100 ( .A(n1142), .B(n1143), .Z(n259) );
  AND U1101 ( .A(n102), .B(n1144), .Z(n1143) );
  XOR U1102 ( .A(n1145), .B(n1142), .Z(n1144) );
  XOR U1103 ( .A(n1146), .B(n1147), .Z(n1134) );
  AND U1104 ( .A(n1148), .B(n1149), .Z(n1147) );
  XOR U1105 ( .A(n1146), .B(n274), .Z(n1149) );
  XOR U1106 ( .A(n1150), .B(n1151), .Z(n274) );
  AND U1107 ( .A(n105), .B(n1152), .Z(n1151) );
  XOR U1108 ( .A(n1153), .B(n1150), .Z(n1152) );
  XNOR U1109 ( .A(n271), .B(n1146), .Z(n1148) );
  XOR U1110 ( .A(n1154), .B(n1155), .Z(n271) );
  AND U1111 ( .A(n102), .B(n1156), .Z(n1155) );
  XOR U1112 ( .A(n1157), .B(n1154), .Z(n1156) );
  XOR U1113 ( .A(n1158), .B(n1159), .Z(n1146) );
  AND U1114 ( .A(n1160), .B(n1161), .Z(n1159) );
  XOR U1115 ( .A(n1158), .B(n286), .Z(n1161) );
  XOR U1116 ( .A(n1162), .B(n1163), .Z(n286) );
  AND U1117 ( .A(n105), .B(n1164), .Z(n1163) );
  XOR U1118 ( .A(n1165), .B(n1162), .Z(n1164) );
  XNOR U1119 ( .A(n283), .B(n1158), .Z(n1160) );
  XOR U1120 ( .A(n1166), .B(n1167), .Z(n283) );
  AND U1121 ( .A(n102), .B(n1168), .Z(n1167) );
  XOR U1122 ( .A(n1169), .B(n1166), .Z(n1168) );
  XOR U1123 ( .A(n1170), .B(n1171), .Z(n1158) );
  AND U1124 ( .A(n1172), .B(n1173), .Z(n1171) );
  XNOR U1125 ( .A(n1174), .B(n298), .Z(n1173) );
  XOR U1126 ( .A(n1175), .B(n1176), .Z(n298) );
  AND U1127 ( .A(n105), .B(n1177), .Z(n1176) );
  XOR U1128 ( .A(n1178), .B(n1175), .Z(n1177) );
  XNOR U1129 ( .A(n295), .B(n1170), .Z(n1172) );
  XOR U1130 ( .A(n1179), .B(n1180), .Z(n295) );
  AND U1131 ( .A(n102), .B(n1181), .Z(n1180) );
  XOR U1132 ( .A(n1182), .B(n1179), .Z(n1181) );
  IV U1133 ( .A(n1174), .Z(n1170) );
  AND U1134 ( .A(n1002), .B(n1005), .Z(n1174) );
  XNOR U1135 ( .A(n1183), .B(n1184), .Z(n1005) );
  AND U1136 ( .A(n105), .B(n1185), .Z(n1184) );
  XNOR U1137 ( .A(n1186), .B(n1183), .Z(n1185) );
  XOR U1138 ( .A(n1187), .B(n1188), .Z(n105) );
  AND U1139 ( .A(n1189), .B(n1190), .Z(n1188) );
  XNOR U1140 ( .A(n1010), .B(n1187), .Z(n1190) );
  AND U1141 ( .A(p_input[127]), .B(p_input[111]), .Z(n1010) );
  XOR U1142 ( .A(n1187), .B(n1011), .Z(n1189) );
  AND U1143 ( .A(p_input[95]), .B(p_input[79]), .Z(n1011) );
  XOR U1144 ( .A(n1191), .B(n1192), .Z(n1187) );
  AND U1145 ( .A(n1193), .B(n1194), .Z(n1192) );
  XOR U1146 ( .A(n1191), .B(n1021), .Z(n1194) );
  XNOR U1147 ( .A(p_input[110]), .B(n1195), .Z(n1021) );
  AND U1148 ( .A(n113), .B(n1196), .Z(n1195) );
  XOR U1149 ( .A(p_input[126]), .B(p_input[110]), .Z(n1196) );
  XNOR U1150 ( .A(n1018), .B(n1191), .Z(n1193) );
  XOR U1151 ( .A(n1197), .B(n1198), .Z(n1018) );
  AND U1152 ( .A(n111), .B(n1199), .Z(n1198) );
  XOR U1153 ( .A(p_input[94]), .B(p_input[78]), .Z(n1199) );
  XOR U1154 ( .A(n1200), .B(n1201), .Z(n1191) );
  AND U1155 ( .A(n1202), .B(n1203), .Z(n1201) );
  XOR U1156 ( .A(n1200), .B(n1033), .Z(n1203) );
  XNOR U1157 ( .A(p_input[109]), .B(n1204), .Z(n1033) );
  AND U1158 ( .A(n113), .B(n1205), .Z(n1204) );
  XOR U1159 ( .A(p_input[125]), .B(p_input[109]), .Z(n1205) );
  XNOR U1160 ( .A(n1030), .B(n1200), .Z(n1202) );
  XOR U1161 ( .A(n1206), .B(n1207), .Z(n1030) );
  AND U1162 ( .A(n111), .B(n1208), .Z(n1207) );
  XOR U1163 ( .A(p_input[93]), .B(p_input[77]), .Z(n1208) );
  XOR U1164 ( .A(n1209), .B(n1210), .Z(n1200) );
  AND U1165 ( .A(n1211), .B(n1212), .Z(n1210) );
  XOR U1166 ( .A(n1209), .B(n1045), .Z(n1212) );
  XNOR U1167 ( .A(p_input[108]), .B(n1213), .Z(n1045) );
  AND U1168 ( .A(n113), .B(n1214), .Z(n1213) );
  XOR U1169 ( .A(p_input[124]), .B(p_input[108]), .Z(n1214) );
  XNOR U1170 ( .A(n1042), .B(n1209), .Z(n1211) );
  XOR U1171 ( .A(n1215), .B(n1216), .Z(n1042) );
  AND U1172 ( .A(n111), .B(n1217), .Z(n1216) );
  XOR U1173 ( .A(p_input[92]), .B(p_input[76]), .Z(n1217) );
  XOR U1174 ( .A(n1218), .B(n1219), .Z(n1209) );
  AND U1175 ( .A(n1220), .B(n1221), .Z(n1219) );
  XOR U1176 ( .A(n1218), .B(n1057), .Z(n1221) );
  XNOR U1177 ( .A(p_input[107]), .B(n1222), .Z(n1057) );
  AND U1178 ( .A(n113), .B(n1223), .Z(n1222) );
  XOR U1179 ( .A(p_input[123]), .B(p_input[107]), .Z(n1223) );
  XNOR U1180 ( .A(n1054), .B(n1218), .Z(n1220) );
  XOR U1181 ( .A(n1224), .B(n1225), .Z(n1054) );
  AND U1182 ( .A(n111), .B(n1226), .Z(n1225) );
  XOR U1183 ( .A(p_input[91]), .B(p_input[75]), .Z(n1226) );
  XOR U1184 ( .A(n1227), .B(n1228), .Z(n1218) );
  AND U1185 ( .A(n1229), .B(n1230), .Z(n1228) );
  XOR U1186 ( .A(n1227), .B(n1069), .Z(n1230) );
  XNOR U1187 ( .A(p_input[106]), .B(n1231), .Z(n1069) );
  AND U1188 ( .A(n113), .B(n1232), .Z(n1231) );
  XOR U1189 ( .A(p_input[122]), .B(p_input[106]), .Z(n1232) );
  XNOR U1190 ( .A(n1066), .B(n1227), .Z(n1229) );
  XOR U1191 ( .A(n1233), .B(n1234), .Z(n1066) );
  AND U1192 ( .A(n111), .B(n1235), .Z(n1234) );
  XOR U1193 ( .A(p_input[90]), .B(p_input[74]), .Z(n1235) );
  XOR U1194 ( .A(n1236), .B(n1237), .Z(n1227) );
  AND U1195 ( .A(n1238), .B(n1239), .Z(n1237) );
  XOR U1196 ( .A(n1236), .B(n1081), .Z(n1239) );
  XNOR U1197 ( .A(p_input[105]), .B(n1240), .Z(n1081) );
  AND U1198 ( .A(n113), .B(n1241), .Z(n1240) );
  XOR U1199 ( .A(p_input[121]), .B(p_input[105]), .Z(n1241) );
  XNOR U1200 ( .A(n1078), .B(n1236), .Z(n1238) );
  XOR U1201 ( .A(n1242), .B(n1243), .Z(n1078) );
  AND U1202 ( .A(n111), .B(n1244), .Z(n1243) );
  XOR U1203 ( .A(p_input[89]), .B(p_input[73]), .Z(n1244) );
  XOR U1204 ( .A(n1245), .B(n1246), .Z(n1236) );
  AND U1205 ( .A(n1247), .B(n1248), .Z(n1246) );
  XOR U1206 ( .A(n1245), .B(n1093), .Z(n1248) );
  XNOR U1207 ( .A(p_input[104]), .B(n1249), .Z(n1093) );
  AND U1208 ( .A(n113), .B(n1250), .Z(n1249) );
  XOR U1209 ( .A(p_input[120]), .B(p_input[104]), .Z(n1250) );
  XNOR U1210 ( .A(n1090), .B(n1245), .Z(n1247) );
  XOR U1211 ( .A(n1251), .B(n1252), .Z(n1090) );
  AND U1212 ( .A(n111), .B(n1253), .Z(n1252) );
  XOR U1213 ( .A(p_input[88]), .B(p_input[72]), .Z(n1253) );
  XOR U1214 ( .A(n1254), .B(n1255), .Z(n1245) );
  AND U1215 ( .A(n1256), .B(n1257), .Z(n1255) );
  XOR U1216 ( .A(n1254), .B(n1105), .Z(n1257) );
  XNOR U1217 ( .A(p_input[103]), .B(n1258), .Z(n1105) );
  AND U1218 ( .A(n113), .B(n1259), .Z(n1258) );
  XOR U1219 ( .A(p_input[119]), .B(p_input[103]), .Z(n1259) );
  XNOR U1220 ( .A(n1102), .B(n1254), .Z(n1256) );
  XOR U1221 ( .A(n1260), .B(n1261), .Z(n1102) );
  AND U1222 ( .A(n111), .B(n1262), .Z(n1261) );
  XOR U1223 ( .A(p_input[87]), .B(p_input[71]), .Z(n1262) );
  XOR U1224 ( .A(n1263), .B(n1264), .Z(n1254) );
  AND U1225 ( .A(n1265), .B(n1266), .Z(n1264) );
  XOR U1226 ( .A(n1263), .B(n1117), .Z(n1266) );
  XNOR U1227 ( .A(p_input[102]), .B(n1267), .Z(n1117) );
  AND U1228 ( .A(n113), .B(n1268), .Z(n1267) );
  XOR U1229 ( .A(p_input[118]), .B(p_input[102]), .Z(n1268) );
  XNOR U1230 ( .A(n1114), .B(n1263), .Z(n1265) );
  XOR U1231 ( .A(n1269), .B(n1270), .Z(n1114) );
  AND U1232 ( .A(n111), .B(n1271), .Z(n1270) );
  XOR U1233 ( .A(p_input[86]), .B(p_input[70]), .Z(n1271) );
  XOR U1234 ( .A(n1272), .B(n1273), .Z(n1263) );
  AND U1235 ( .A(n1274), .B(n1275), .Z(n1273) );
  XOR U1236 ( .A(n1129), .B(n1272), .Z(n1275) );
  XNOR U1237 ( .A(p_input[101]), .B(n1276), .Z(n1129) );
  AND U1238 ( .A(n113), .B(n1277), .Z(n1276) );
  XOR U1239 ( .A(p_input[117]), .B(p_input[101]), .Z(n1277) );
  XNOR U1240 ( .A(n1272), .B(n1126), .Z(n1274) );
  XOR U1241 ( .A(n1278), .B(n1279), .Z(n1126) );
  AND U1242 ( .A(n111), .B(n1280), .Z(n1279) );
  XOR U1243 ( .A(p_input[85]), .B(p_input[69]), .Z(n1280) );
  XOR U1244 ( .A(n1281), .B(n1282), .Z(n1272) );
  AND U1245 ( .A(n1283), .B(n1284), .Z(n1282) );
  XOR U1246 ( .A(n1281), .B(n1141), .Z(n1284) );
  XNOR U1247 ( .A(p_input[100]), .B(n1285), .Z(n1141) );
  AND U1248 ( .A(n113), .B(n1286), .Z(n1285) );
  XOR U1249 ( .A(p_input[116]), .B(p_input[100]), .Z(n1286) );
  XNOR U1250 ( .A(n1138), .B(n1281), .Z(n1283) );
  XOR U1251 ( .A(n1287), .B(n1288), .Z(n1138) );
  AND U1252 ( .A(n111), .B(n1289), .Z(n1288) );
  XOR U1253 ( .A(p_input[84]), .B(p_input[68]), .Z(n1289) );
  XOR U1254 ( .A(n1290), .B(n1291), .Z(n1281) );
  AND U1255 ( .A(n1292), .B(n1293), .Z(n1291) );
  XOR U1256 ( .A(n1290), .B(n1153), .Z(n1293) );
  XNOR U1257 ( .A(p_input[99]), .B(n1294), .Z(n1153) );
  AND U1258 ( .A(n113), .B(n1295), .Z(n1294) );
  XOR U1259 ( .A(p_input[99]), .B(p_input[115]), .Z(n1295) );
  XNOR U1260 ( .A(n1150), .B(n1290), .Z(n1292) );
  XOR U1261 ( .A(n1296), .B(n1297), .Z(n1150) );
  AND U1262 ( .A(n111), .B(n1298), .Z(n1297) );
  XOR U1263 ( .A(p_input[83]), .B(p_input[67]), .Z(n1298) );
  XOR U1264 ( .A(n1299), .B(n1300), .Z(n1290) );
  AND U1265 ( .A(n1301), .B(n1302), .Z(n1300) );
  XOR U1266 ( .A(n1299), .B(n1165), .Z(n1302) );
  XNOR U1267 ( .A(p_input[98]), .B(n1303), .Z(n1165) );
  AND U1268 ( .A(n113), .B(n1304), .Z(n1303) );
  XOR U1269 ( .A(p_input[98]), .B(p_input[114]), .Z(n1304) );
  XNOR U1270 ( .A(n1162), .B(n1299), .Z(n1301) );
  XOR U1271 ( .A(n1305), .B(n1306), .Z(n1162) );
  AND U1272 ( .A(n111), .B(n1307), .Z(n1306) );
  XOR U1273 ( .A(p_input[82]), .B(p_input[66]), .Z(n1307) );
  XOR U1274 ( .A(n1308), .B(n1309), .Z(n1299) );
  AND U1275 ( .A(n1310), .B(n1311), .Z(n1309) );
  XNOR U1276 ( .A(n1312), .B(n1178), .Z(n1311) );
  XNOR U1277 ( .A(p_input[97]), .B(n1313), .Z(n1178) );
  AND U1278 ( .A(n113), .B(n1314), .Z(n1313) );
  XNOR U1279 ( .A(n1315), .B(p_input[113]), .Z(n1314) );
  IV U1280 ( .A(p_input[97]), .Z(n1315) );
  XNOR U1281 ( .A(n1175), .B(n1308), .Z(n1310) );
  XNOR U1282 ( .A(p_input[65]), .B(n1316), .Z(n1175) );
  AND U1283 ( .A(n111), .B(n1317), .Z(n1316) );
  XOR U1284 ( .A(p_input[81]), .B(p_input[65]), .Z(n1317) );
  IV U1285 ( .A(n1312), .Z(n1308) );
  AND U1286 ( .A(n1183), .B(n1186), .Z(n1312) );
  XOR U1287 ( .A(p_input[96]), .B(n1318), .Z(n1186) );
  AND U1288 ( .A(n113), .B(n1319), .Z(n1318) );
  XOR U1289 ( .A(p_input[96]), .B(p_input[112]), .Z(n1319) );
  XOR U1290 ( .A(n1320), .B(n1321), .Z(n113) );
  AND U1291 ( .A(n1322), .B(n1323), .Z(n1321) );
  XNOR U1292 ( .A(p_input[127]), .B(n1320), .Z(n1323) );
  XOR U1293 ( .A(n1320), .B(p_input[111]), .Z(n1322) );
  XOR U1294 ( .A(n1324), .B(n1325), .Z(n1320) );
  AND U1295 ( .A(n1326), .B(n1327), .Z(n1325) );
  XNOR U1296 ( .A(p_input[126]), .B(n1324), .Z(n1327) );
  XOR U1297 ( .A(n1324), .B(p_input[110]), .Z(n1326) );
  XOR U1298 ( .A(n1328), .B(n1329), .Z(n1324) );
  AND U1299 ( .A(n1330), .B(n1331), .Z(n1329) );
  XNOR U1300 ( .A(p_input[125]), .B(n1328), .Z(n1331) );
  XOR U1301 ( .A(n1328), .B(p_input[109]), .Z(n1330) );
  XOR U1302 ( .A(n1332), .B(n1333), .Z(n1328) );
  AND U1303 ( .A(n1334), .B(n1335), .Z(n1333) );
  XNOR U1304 ( .A(p_input[124]), .B(n1332), .Z(n1335) );
  XOR U1305 ( .A(n1332), .B(p_input[108]), .Z(n1334) );
  XOR U1306 ( .A(n1336), .B(n1337), .Z(n1332) );
  AND U1307 ( .A(n1338), .B(n1339), .Z(n1337) );
  XNOR U1308 ( .A(p_input[123]), .B(n1336), .Z(n1339) );
  XOR U1309 ( .A(n1336), .B(p_input[107]), .Z(n1338) );
  XOR U1310 ( .A(n1340), .B(n1341), .Z(n1336) );
  AND U1311 ( .A(n1342), .B(n1343), .Z(n1341) );
  XNOR U1312 ( .A(p_input[122]), .B(n1340), .Z(n1343) );
  XOR U1313 ( .A(n1340), .B(p_input[106]), .Z(n1342) );
  XOR U1314 ( .A(n1344), .B(n1345), .Z(n1340) );
  AND U1315 ( .A(n1346), .B(n1347), .Z(n1345) );
  XNOR U1316 ( .A(p_input[121]), .B(n1344), .Z(n1347) );
  XOR U1317 ( .A(n1344), .B(p_input[105]), .Z(n1346) );
  XOR U1318 ( .A(n1348), .B(n1349), .Z(n1344) );
  AND U1319 ( .A(n1350), .B(n1351), .Z(n1349) );
  XNOR U1320 ( .A(p_input[120]), .B(n1348), .Z(n1351) );
  XOR U1321 ( .A(n1348), .B(p_input[104]), .Z(n1350) );
  XOR U1322 ( .A(n1352), .B(n1353), .Z(n1348) );
  AND U1323 ( .A(n1354), .B(n1355), .Z(n1353) );
  XNOR U1324 ( .A(p_input[119]), .B(n1352), .Z(n1355) );
  XOR U1325 ( .A(n1352), .B(p_input[103]), .Z(n1354) );
  XOR U1326 ( .A(n1356), .B(n1357), .Z(n1352) );
  AND U1327 ( .A(n1358), .B(n1359), .Z(n1357) );
  XNOR U1328 ( .A(p_input[118]), .B(n1356), .Z(n1359) );
  XOR U1329 ( .A(n1356), .B(p_input[102]), .Z(n1358) );
  XOR U1330 ( .A(n1360), .B(n1361), .Z(n1356) );
  AND U1331 ( .A(n1362), .B(n1363), .Z(n1361) );
  XNOR U1332 ( .A(p_input[117]), .B(n1360), .Z(n1363) );
  XOR U1333 ( .A(n1360), .B(p_input[101]), .Z(n1362) );
  XOR U1334 ( .A(n1364), .B(n1365), .Z(n1360) );
  AND U1335 ( .A(n1366), .B(n1367), .Z(n1365) );
  XNOR U1336 ( .A(p_input[116]), .B(n1364), .Z(n1367) );
  XOR U1337 ( .A(n1364), .B(p_input[100]), .Z(n1366) );
  XOR U1338 ( .A(n1368), .B(n1369), .Z(n1364) );
  AND U1339 ( .A(n1370), .B(n1371), .Z(n1369) );
  XNOR U1340 ( .A(p_input[115]), .B(n1368), .Z(n1371) );
  XOR U1341 ( .A(n1368), .B(p_input[99]), .Z(n1370) );
  XOR U1342 ( .A(n1372), .B(n1373), .Z(n1368) );
  AND U1343 ( .A(n1374), .B(n1375), .Z(n1373) );
  XNOR U1344 ( .A(p_input[114]), .B(n1372), .Z(n1375) );
  XOR U1345 ( .A(n1372), .B(p_input[98]), .Z(n1374) );
  XNOR U1346 ( .A(n1376), .B(n1377), .Z(n1372) );
  AND U1347 ( .A(n1378), .B(n1379), .Z(n1377) );
  XOR U1348 ( .A(p_input[113]), .B(n1376), .Z(n1379) );
  XNOR U1349 ( .A(p_input[97]), .B(n1376), .Z(n1378) );
  AND U1350 ( .A(p_input[112]), .B(n1380), .Z(n1376) );
  IV U1351 ( .A(p_input[96]), .Z(n1380) );
  XNOR U1352 ( .A(p_input[64]), .B(n1381), .Z(n1183) );
  AND U1353 ( .A(n111), .B(n1382), .Z(n1381) );
  XOR U1354 ( .A(p_input[80]), .B(p_input[64]), .Z(n1382) );
  XOR U1355 ( .A(n1383), .B(n1384), .Z(n111) );
  AND U1356 ( .A(n1385), .B(n1386), .Z(n1384) );
  XNOR U1357 ( .A(p_input[95]), .B(n1383), .Z(n1386) );
  XOR U1358 ( .A(n1383), .B(p_input[79]), .Z(n1385) );
  XOR U1359 ( .A(n1387), .B(n1388), .Z(n1383) );
  AND U1360 ( .A(n1389), .B(n1390), .Z(n1388) );
  XNOR U1361 ( .A(p_input[94]), .B(n1387), .Z(n1390) );
  XNOR U1362 ( .A(n1387), .B(n1197), .Z(n1389) );
  IV U1363 ( .A(p_input[78]), .Z(n1197) );
  XOR U1364 ( .A(n1391), .B(n1392), .Z(n1387) );
  AND U1365 ( .A(n1393), .B(n1394), .Z(n1392) );
  XNOR U1366 ( .A(p_input[93]), .B(n1391), .Z(n1394) );
  XNOR U1367 ( .A(n1391), .B(n1206), .Z(n1393) );
  IV U1368 ( .A(p_input[77]), .Z(n1206) );
  XOR U1369 ( .A(n1395), .B(n1396), .Z(n1391) );
  AND U1370 ( .A(n1397), .B(n1398), .Z(n1396) );
  XNOR U1371 ( .A(p_input[92]), .B(n1395), .Z(n1398) );
  XNOR U1372 ( .A(n1395), .B(n1215), .Z(n1397) );
  IV U1373 ( .A(p_input[76]), .Z(n1215) );
  XOR U1374 ( .A(n1399), .B(n1400), .Z(n1395) );
  AND U1375 ( .A(n1401), .B(n1402), .Z(n1400) );
  XNOR U1376 ( .A(p_input[91]), .B(n1399), .Z(n1402) );
  XNOR U1377 ( .A(n1399), .B(n1224), .Z(n1401) );
  IV U1378 ( .A(p_input[75]), .Z(n1224) );
  XOR U1379 ( .A(n1403), .B(n1404), .Z(n1399) );
  AND U1380 ( .A(n1405), .B(n1406), .Z(n1404) );
  XNOR U1381 ( .A(p_input[90]), .B(n1403), .Z(n1406) );
  XNOR U1382 ( .A(n1403), .B(n1233), .Z(n1405) );
  IV U1383 ( .A(p_input[74]), .Z(n1233) );
  XOR U1384 ( .A(n1407), .B(n1408), .Z(n1403) );
  AND U1385 ( .A(n1409), .B(n1410), .Z(n1408) );
  XNOR U1386 ( .A(p_input[89]), .B(n1407), .Z(n1410) );
  XNOR U1387 ( .A(n1407), .B(n1242), .Z(n1409) );
  IV U1388 ( .A(p_input[73]), .Z(n1242) );
  XOR U1389 ( .A(n1411), .B(n1412), .Z(n1407) );
  AND U1390 ( .A(n1413), .B(n1414), .Z(n1412) );
  XNOR U1391 ( .A(p_input[88]), .B(n1411), .Z(n1414) );
  XNOR U1392 ( .A(n1411), .B(n1251), .Z(n1413) );
  IV U1393 ( .A(p_input[72]), .Z(n1251) );
  XOR U1394 ( .A(n1415), .B(n1416), .Z(n1411) );
  AND U1395 ( .A(n1417), .B(n1418), .Z(n1416) );
  XNOR U1396 ( .A(p_input[87]), .B(n1415), .Z(n1418) );
  XNOR U1397 ( .A(n1415), .B(n1260), .Z(n1417) );
  IV U1398 ( .A(p_input[71]), .Z(n1260) );
  XOR U1399 ( .A(n1419), .B(n1420), .Z(n1415) );
  AND U1400 ( .A(n1421), .B(n1422), .Z(n1420) );
  XNOR U1401 ( .A(p_input[86]), .B(n1419), .Z(n1422) );
  XNOR U1402 ( .A(n1419), .B(n1269), .Z(n1421) );
  IV U1403 ( .A(p_input[70]), .Z(n1269) );
  XOR U1404 ( .A(n1423), .B(n1424), .Z(n1419) );
  AND U1405 ( .A(n1425), .B(n1426), .Z(n1424) );
  XNOR U1406 ( .A(p_input[85]), .B(n1423), .Z(n1426) );
  XNOR U1407 ( .A(n1423), .B(n1278), .Z(n1425) );
  IV U1408 ( .A(p_input[69]), .Z(n1278) );
  XOR U1409 ( .A(n1427), .B(n1428), .Z(n1423) );
  AND U1410 ( .A(n1429), .B(n1430), .Z(n1428) );
  XNOR U1411 ( .A(p_input[84]), .B(n1427), .Z(n1430) );
  XNOR U1412 ( .A(n1427), .B(n1287), .Z(n1429) );
  IV U1413 ( .A(p_input[68]), .Z(n1287) );
  XOR U1414 ( .A(n1431), .B(n1432), .Z(n1427) );
  AND U1415 ( .A(n1433), .B(n1434), .Z(n1432) );
  XNOR U1416 ( .A(p_input[83]), .B(n1431), .Z(n1434) );
  XNOR U1417 ( .A(n1431), .B(n1296), .Z(n1433) );
  IV U1418 ( .A(p_input[67]), .Z(n1296) );
  XOR U1419 ( .A(n1435), .B(n1436), .Z(n1431) );
  AND U1420 ( .A(n1437), .B(n1438), .Z(n1436) );
  XNOR U1421 ( .A(p_input[82]), .B(n1435), .Z(n1438) );
  XNOR U1422 ( .A(n1435), .B(n1305), .Z(n1437) );
  IV U1423 ( .A(p_input[66]), .Z(n1305) );
  XNOR U1424 ( .A(n1439), .B(n1440), .Z(n1435) );
  AND U1425 ( .A(n1441), .B(n1442), .Z(n1440) );
  XOR U1426 ( .A(p_input[81]), .B(n1439), .Z(n1442) );
  XNOR U1427 ( .A(p_input[65]), .B(n1439), .Z(n1441) );
  AND U1428 ( .A(p_input[80]), .B(n1443), .Z(n1439) );
  IV U1429 ( .A(p_input[64]), .Z(n1443) );
  XOR U1430 ( .A(n1444), .B(n1445), .Z(n1002) );
  AND U1431 ( .A(n102), .B(n1446), .Z(n1445) );
  XNOR U1432 ( .A(n1447), .B(n1444), .Z(n1446) );
  XOR U1433 ( .A(n1448), .B(n1449), .Z(n102) );
  AND U1434 ( .A(n1450), .B(n1451), .Z(n1449) );
  XNOR U1435 ( .A(n1013), .B(n1448), .Z(n1451) );
  AND U1436 ( .A(p_input[63]), .B(p_input[47]), .Z(n1013) );
  XOR U1437 ( .A(n1448), .B(n1012), .Z(n1450) );
  AND U1438 ( .A(p_input[15]), .B(p_input[31]), .Z(n1012) );
  XOR U1439 ( .A(n1452), .B(n1453), .Z(n1448) );
  AND U1440 ( .A(n1454), .B(n1455), .Z(n1453) );
  XOR U1441 ( .A(n1452), .B(n1025), .Z(n1455) );
  XNOR U1442 ( .A(p_input[46]), .B(n1456), .Z(n1025) );
  AND U1443 ( .A(n121), .B(n1457), .Z(n1456) );
  XOR U1444 ( .A(p_input[62]), .B(p_input[46]), .Z(n1457) );
  XNOR U1445 ( .A(n1022), .B(n1452), .Z(n1454) );
  XOR U1446 ( .A(n1458), .B(n1459), .Z(n1022) );
  AND U1447 ( .A(n118), .B(n1460), .Z(n1459) );
  XOR U1448 ( .A(p_input[30]), .B(p_input[14]), .Z(n1460) );
  XOR U1449 ( .A(n1461), .B(n1462), .Z(n1452) );
  AND U1450 ( .A(n1463), .B(n1464), .Z(n1462) );
  XOR U1451 ( .A(n1461), .B(n1037), .Z(n1464) );
  XNOR U1452 ( .A(p_input[45]), .B(n1465), .Z(n1037) );
  AND U1453 ( .A(n121), .B(n1466), .Z(n1465) );
  XOR U1454 ( .A(p_input[61]), .B(p_input[45]), .Z(n1466) );
  XNOR U1455 ( .A(n1034), .B(n1461), .Z(n1463) );
  XOR U1456 ( .A(n1467), .B(n1468), .Z(n1034) );
  AND U1457 ( .A(n118), .B(n1469), .Z(n1468) );
  XOR U1458 ( .A(p_input[29]), .B(p_input[13]), .Z(n1469) );
  XOR U1459 ( .A(n1470), .B(n1471), .Z(n1461) );
  AND U1460 ( .A(n1472), .B(n1473), .Z(n1471) );
  XOR U1461 ( .A(n1470), .B(n1049), .Z(n1473) );
  XNOR U1462 ( .A(p_input[44]), .B(n1474), .Z(n1049) );
  AND U1463 ( .A(n121), .B(n1475), .Z(n1474) );
  XOR U1464 ( .A(p_input[60]), .B(p_input[44]), .Z(n1475) );
  XNOR U1465 ( .A(n1046), .B(n1470), .Z(n1472) );
  XOR U1466 ( .A(n1476), .B(n1477), .Z(n1046) );
  AND U1467 ( .A(n118), .B(n1478), .Z(n1477) );
  XOR U1468 ( .A(p_input[28]), .B(p_input[12]), .Z(n1478) );
  XOR U1469 ( .A(n1479), .B(n1480), .Z(n1470) );
  AND U1470 ( .A(n1481), .B(n1482), .Z(n1480) );
  XOR U1471 ( .A(n1479), .B(n1061), .Z(n1482) );
  XNOR U1472 ( .A(p_input[43]), .B(n1483), .Z(n1061) );
  AND U1473 ( .A(n121), .B(n1484), .Z(n1483) );
  XOR U1474 ( .A(p_input[59]), .B(p_input[43]), .Z(n1484) );
  XNOR U1475 ( .A(n1058), .B(n1479), .Z(n1481) );
  XOR U1476 ( .A(n1485), .B(n1486), .Z(n1058) );
  AND U1477 ( .A(n118), .B(n1487), .Z(n1486) );
  XOR U1478 ( .A(p_input[27]), .B(p_input[11]), .Z(n1487) );
  XOR U1479 ( .A(n1488), .B(n1489), .Z(n1479) );
  AND U1480 ( .A(n1490), .B(n1491), .Z(n1489) );
  XOR U1481 ( .A(n1488), .B(n1073), .Z(n1491) );
  XNOR U1482 ( .A(p_input[42]), .B(n1492), .Z(n1073) );
  AND U1483 ( .A(n121), .B(n1493), .Z(n1492) );
  XOR U1484 ( .A(p_input[58]), .B(p_input[42]), .Z(n1493) );
  XNOR U1485 ( .A(n1070), .B(n1488), .Z(n1490) );
  XOR U1486 ( .A(n1494), .B(n1495), .Z(n1070) );
  AND U1487 ( .A(n118), .B(n1496), .Z(n1495) );
  XOR U1488 ( .A(p_input[26]), .B(p_input[10]), .Z(n1496) );
  XOR U1489 ( .A(n1497), .B(n1498), .Z(n1488) );
  AND U1490 ( .A(n1499), .B(n1500), .Z(n1498) );
  XOR U1491 ( .A(n1497), .B(n1085), .Z(n1500) );
  XNOR U1492 ( .A(p_input[41]), .B(n1501), .Z(n1085) );
  AND U1493 ( .A(n121), .B(n1502), .Z(n1501) );
  XOR U1494 ( .A(p_input[57]), .B(p_input[41]), .Z(n1502) );
  XNOR U1495 ( .A(n1082), .B(n1497), .Z(n1499) );
  XOR U1496 ( .A(n1503), .B(n1504), .Z(n1082) );
  AND U1497 ( .A(n118), .B(n1505), .Z(n1504) );
  XOR U1498 ( .A(p_input[9]), .B(p_input[25]), .Z(n1505) );
  XOR U1499 ( .A(n1506), .B(n1507), .Z(n1497) );
  AND U1500 ( .A(n1508), .B(n1509), .Z(n1507) );
  XOR U1501 ( .A(n1506), .B(n1097), .Z(n1509) );
  XNOR U1502 ( .A(p_input[40]), .B(n1510), .Z(n1097) );
  AND U1503 ( .A(n121), .B(n1511), .Z(n1510) );
  XOR U1504 ( .A(p_input[56]), .B(p_input[40]), .Z(n1511) );
  XNOR U1505 ( .A(n1094), .B(n1506), .Z(n1508) );
  XOR U1506 ( .A(n1512), .B(n1513), .Z(n1094) );
  AND U1507 ( .A(n118), .B(n1514), .Z(n1513) );
  XOR U1508 ( .A(p_input[8]), .B(p_input[24]), .Z(n1514) );
  XOR U1509 ( .A(n1515), .B(n1516), .Z(n1506) );
  AND U1510 ( .A(n1517), .B(n1518), .Z(n1516) );
  XOR U1511 ( .A(n1515), .B(n1109), .Z(n1518) );
  XNOR U1512 ( .A(p_input[39]), .B(n1519), .Z(n1109) );
  AND U1513 ( .A(n121), .B(n1520), .Z(n1519) );
  XOR U1514 ( .A(p_input[55]), .B(p_input[39]), .Z(n1520) );
  XNOR U1515 ( .A(n1106), .B(n1515), .Z(n1517) );
  XOR U1516 ( .A(n1521), .B(n1522), .Z(n1106) );
  AND U1517 ( .A(n118), .B(n1523), .Z(n1522) );
  XOR U1518 ( .A(p_input[7]), .B(p_input[23]), .Z(n1523) );
  XOR U1519 ( .A(n1524), .B(n1525), .Z(n1515) );
  AND U1520 ( .A(n1526), .B(n1527), .Z(n1525) );
  XOR U1521 ( .A(n1524), .B(n1121), .Z(n1527) );
  XNOR U1522 ( .A(p_input[38]), .B(n1528), .Z(n1121) );
  AND U1523 ( .A(n121), .B(n1529), .Z(n1528) );
  XOR U1524 ( .A(p_input[54]), .B(p_input[38]), .Z(n1529) );
  XNOR U1525 ( .A(n1118), .B(n1524), .Z(n1526) );
  XOR U1526 ( .A(n1530), .B(n1531), .Z(n1118) );
  AND U1527 ( .A(n118), .B(n1532), .Z(n1531) );
  XOR U1528 ( .A(p_input[6]), .B(p_input[22]), .Z(n1532) );
  XOR U1529 ( .A(n1533), .B(n1534), .Z(n1524) );
  AND U1530 ( .A(n1535), .B(n1536), .Z(n1534) );
  XOR U1531 ( .A(n1133), .B(n1533), .Z(n1536) );
  XNOR U1532 ( .A(p_input[37]), .B(n1537), .Z(n1133) );
  AND U1533 ( .A(n121), .B(n1538), .Z(n1537) );
  XOR U1534 ( .A(p_input[53]), .B(p_input[37]), .Z(n1538) );
  XNOR U1535 ( .A(n1533), .B(n1130), .Z(n1535) );
  XOR U1536 ( .A(n1539), .B(n1540), .Z(n1130) );
  AND U1537 ( .A(n118), .B(n1541), .Z(n1540) );
  XOR U1538 ( .A(p_input[5]), .B(p_input[21]), .Z(n1541) );
  XOR U1539 ( .A(n1542), .B(n1543), .Z(n1533) );
  AND U1540 ( .A(n1544), .B(n1545), .Z(n1543) );
  XOR U1541 ( .A(n1542), .B(n1145), .Z(n1545) );
  XNOR U1542 ( .A(p_input[36]), .B(n1546), .Z(n1145) );
  AND U1543 ( .A(n121), .B(n1547), .Z(n1546) );
  XOR U1544 ( .A(p_input[52]), .B(p_input[36]), .Z(n1547) );
  XNOR U1545 ( .A(n1142), .B(n1542), .Z(n1544) );
  XOR U1546 ( .A(n1548), .B(n1549), .Z(n1142) );
  AND U1547 ( .A(n118), .B(n1550), .Z(n1549) );
  XOR U1548 ( .A(p_input[4]), .B(p_input[20]), .Z(n1550) );
  XOR U1549 ( .A(n1551), .B(n1552), .Z(n1542) );
  AND U1550 ( .A(n1553), .B(n1554), .Z(n1552) );
  XOR U1551 ( .A(n1551), .B(n1157), .Z(n1554) );
  XNOR U1552 ( .A(p_input[35]), .B(n1555), .Z(n1157) );
  AND U1553 ( .A(n121), .B(n1556), .Z(n1555) );
  XOR U1554 ( .A(p_input[51]), .B(p_input[35]), .Z(n1556) );
  XNOR U1555 ( .A(n1154), .B(n1551), .Z(n1553) );
  XOR U1556 ( .A(n1557), .B(n1558), .Z(n1154) );
  AND U1557 ( .A(n118), .B(n1559), .Z(n1558) );
  XOR U1558 ( .A(p_input[3]), .B(p_input[19]), .Z(n1559) );
  XOR U1559 ( .A(n1560), .B(n1561), .Z(n1551) );
  AND U1560 ( .A(n1562), .B(n1563), .Z(n1561) );
  XOR U1561 ( .A(n1560), .B(n1169), .Z(n1563) );
  XNOR U1562 ( .A(p_input[34]), .B(n1564), .Z(n1169) );
  AND U1563 ( .A(n121), .B(n1565), .Z(n1564) );
  XOR U1564 ( .A(p_input[50]), .B(p_input[34]), .Z(n1565) );
  XNOR U1565 ( .A(n1166), .B(n1560), .Z(n1562) );
  XOR U1566 ( .A(n1566), .B(n1567), .Z(n1166) );
  AND U1567 ( .A(n118), .B(n1568), .Z(n1567) );
  XOR U1568 ( .A(p_input[2]), .B(p_input[18]), .Z(n1568) );
  XOR U1569 ( .A(n1569), .B(n1570), .Z(n1560) );
  AND U1570 ( .A(n1571), .B(n1572), .Z(n1570) );
  XNOR U1571 ( .A(n1573), .B(n1182), .Z(n1572) );
  XNOR U1572 ( .A(p_input[33]), .B(n1574), .Z(n1182) );
  AND U1573 ( .A(n121), .B(n1575), .Z(n1574) );
  XNOR U1574 ( .A(p_input[49]), .B(n1576), .Z(n1575) );
  IV U1575 ( .A(p_input[33]), .Z(n1576) );
  XNOR U1576 ( .A(n1179), .B(n1569), .Z(n1571) );
  XNOR U1577 ( .A(p_input[1]), .B(n1577), .Z(n1179) );
  AND U1578 ( .A(n118), .B(n1578), .Z(n1577) );
  XOR U1579 ( .A(p_input[1]), .B(p_input[17]), .Z(n1578) );
  IV U1580 ( .A(n1573), .Z(n1569) );
  AND U1581 ( .A(n1444), .B(n1447), .Z(n1573) );
  XOR U1582 ( .A(p_input[32]), .B(n1579), .Z(n1447) );
  AND U1583 ( .A(n121), .B(n1580), .Z(n1579) );
  XOR U1584 ( .A(p_input[48]), .B(p_input[32]), .Z(n1580) );
  XOR U1585 ( .A(n1581), .B(n1582), .Z(n121) );
  AND U1586 ( .A(n1583), .B(n1584), .Z(n1582) );
  XNOR U1587 ( .A(p_input[63]), .B(n1581), .Z(n1584) );
  XOR U1588 ( .A(n1581), .B(p_input[47]), .Z(n1583) );
  XOR U1589 ( .A(n1585), .B(n1586), .Z(n1581) );
  AND U1590 ( .A(n1587), .B(n1588), .Z(n1586) );
  XNOR U1591 ( .A(p_input[62]), .B(n1585), .Z(n1588) );
  XOR U1592 ( .A(n1585), .B(p_input[46]), .Z(n1587) );
  XOR U1593 ( .A(n1589), .B(n1590), .Z(n1585) );
  AND U1594 ( .A(n1591), .B(n1592), .Z(n1590) );
  XNOR U1595 ( .A(p_input[61]), .B(n1589), .Z(n1592) );
  XOR U1596 ( .A(n1589), .B(p_input[45]), .Z(n1591) );
  XOR U1597 ( .A(n1593), .B(n1594), .Z(n1589) );
  AND U1598 ( .A(n1595), .B(n1596), .Z(n1594) );
  XNOR U1599 ( .A(p_input[60]), .B(n1593), .Z(n1596) );
  XOR U1600 ( .A(n1593), .B(p_input[44]), .Z(n1595) );
  XOR U1601 ( .A(n1597), .B(n1598), .Z(n1593) );
  AND U1602 ( .A(n1599), .B(n1600), .Z(n1598) );
  XNOR U1603 ( .A(p_input[59]), .B(n1597), .Z(n1600) );
  XOR U1604 ( .A(n1597), .B(p_input[43]), .Z(n1599) );
  XOR U1605 ( .A(n1601), .B(n1602), .Z(n1597) );
  AND U1606 ( .A(n1603), .B(n1604), .Z(n1602) );
  XNOR U1607 ( .A(p_input[58]), .B(n1601), .Z(n1604) );
  XOR U1608 ( .A(n1601), .B(p_input[42]), .Z(n1603) );
  XOR U1609 ( .A(n1605), .B(n1606), .Z(n1601) );
  AND U1610 ( .A(n1607), .B(n1608), .Z(n1606) );
  XNOR U1611 ( .A(p_input[57]), .B(n1605), .Z(n1608) );
  XOR U1612 ( .A(n1605), .B(p_input[41]), .Z(n1607) );
  XOR U1613 ( .A(n1609), .B(n1610), .Z(n1605) );
  AND U1614 ( .A(n1611), .B(n1612), .Z(n1610) );
  XNOR U1615 ( .A(p_input[56]), .B(n1609), .Z(n1612) );
  XOR U1616 ( .A(n1609), .B(p_input[40]), .Z(n1611) );
  XOR U1617 ( .A(n1613), .B(n1614), .Z(n1609) );
  AND U1618 ( .A(n1615), .B(n1616), .Z(n1614) );
  XNOR U1619 ( .A(p_input[55]), .B(n1613), .Z(n1616) );
  XOR U1620 ( .A(n1613), .B(p_input[39]), .Z(n1615) );
  XOR U1621 ( .A(n1617), .B(n1618), .Z(n1613) );
  AND U1622 ( .A(n1619), .B(n1620), .Z(n1618) );
  XNOR U1623 ( .A(p_input[54]), .B(n1617), .Z(n1620) );
  XOR U1624 ( .A(n1617), .B(p_input[38]), .Z(n1619) );
  XOR U1625 ( .A(n1621), .B(n1622), .Z(n1617) );
  AND U1626 ( .A(n1623), .B(n1624), .Z(n1622) );
  XNOR U1627 ( .A(p_input[53]), .B(n1621), .Z(n1624) );
  XOR U1628 ( .A(n1621), .B(p_input[37]), .Z(n1623) );
  XOR U1629 ( .A(n1625), .B(n1626), .Z(n1621) );
  AND U1630 ( .A(n1627), .B(n1628), .Z(n1626) );
  XNOR U1631 ( .A(p_input[52]), .B(n1625), .Z(n1628) );
  XOR U1632 ( .A(n1625), .B(p_input[36]), .Z(n1627) );
  XOR U1633 ( .A(n1629), .B(n1630), .Z(n1625) );
  AND U1634 ( .A(n1631), .B(n1632), .Z(n1630) );
  XNOR U1635 ( .A(p_input[51]), .B(n1629), .Z(n1632) );
  XOR U1636 ( .A(n1629), .B(p_input[35]), .Z(n1631) );
  XOR U1637 ( .A(n1633), .B(n1634), .Z(n1629) );
  AND U1638 ( .A(n1635), .B(n1636), .Z(n1634) );
  XNOR U1639 ( .A(p_input[50]), .B(n1633), .Z(n1636) );
  XOR U1640 ( .A(n1633), .B(p_input[34]), .Z(n1635) );
  XNOR U1641 ( .A(n1637), .B(n1638), .Z(n1633) );
  AND U1642 ( .A(n1639), .B(n1640), .Z(n1638) );
  XOR U1643 ( .A(p_input[49]), .B(n1637), .Z(n1640) );
  XNOR U1644 ( .A(p_input[33]), .B(n1637), .Z(n1639) );
  AND U1645 ( .A(p_input[48]), .B(n1641), .Z(n1637) );
  IV U1646 ( .A(p_input[32]), .Z(n1641) );
  XNOR U1647 ( .A(p_input[0]), .B(n1642), .Z(n1444) );
  AND U1648 ( .A(n118), .B(n1643), .Z(n1642) );
  XOR U1649 ( .A(p_input[16]), .B(p_input[0]), .Z(n1643) );
  XOR U1650 ( .A(n1644), .B(n1645), .Z(n118) );
  AND U1651 ( .A(n1646), .B(n1647), .Z(n1645) );
  XNOR U1652 ( .A(p_input[31]), .B(n1644), .Z(n1647) );
  XOR U1653 ( .A(n1644), .B(p_input[15]), .Z(n1646) );
  XOR U1654 ( .A(n1648), .B(n1649), .Z(n1644) );
  AND U1655 ( .A(n1650), .B(n1651), .Z(n1649) );
  XNOR U1656 ( .A(p_input[30]), .B(n1648), .Z(n1651) );
  XNOR U1657 ( .A(n1648), .B(n1458), .Z(n1650) );
  IV U1658 ( .A(p_input[14]), .Z(n1458) );
  XOR U1659 ( .A(n1652), .B(n1653), .Z(n1648) );
  AND U1660 ( .A(n1654), .B(n1655), .Z(n1653) );
  XNOR U1661 ( .A(p_input[29]), .B(n1652), .Z(n1655) );
  XNOR U1662 ( .A(n1652), .B(n1467), .Z(n1654) );
  IV U1663 ( .A(p_input[13]), .Z(n1467) );
  XOR U1664 ( .A(n1656), .B(n1657), .Z(n1652) );
  AND U1665 ( .A(n1658), .B(n1659), .Z(n1657) );
  XNOR U1666 ( .A(p_input[28]), .B(n1656), .Z(n1659) );
  XNOR U1667 ( .A(n1656), .B(n1476), .Z(n1658) );
  IV U1668 ( .A(p_input[12]), .Z(n1476) );
  XOR U1669 ( .A(n1660), .B(n1661), .Z(n1656) );
  AND U1670 ( .A(n1662), .B(n1663), .Z(n1661) );
  XNOR U1671 ( .A(p_input[27]), .B(n1660), .Z(n1663) );
  XNOR U1672 ( .A(n1660), .B(n1485), .Z(n1662) );
  IV U1673 ( .A(p_input[11]), .Z(n1485) );
  XOR U1674 ( .A(n1664), .B(n1665), .Z(n1660) );
  AND U1675 ( .A(n1666), .B(n1667), .Z(n1665) );
  XNOR U1676 ( .A(p_input[26]), .B(n1664), .Z(n1667) );
  XNOR U1677 ( .A(n1664), .B(n1494), .Z(n1666) );
  IV U1678 ( .A(p_input[10]), .Z(n1494) );
  XOR U1679 ( .A(n1668), .B(n1669), .Z(n1664) );
  AND U1680 ( .A(n1670), .B(n1671), .Z(n1669) );
  XNOR U1681 ( .A(p_input[25]), .B(n1668), .Z(n1671) );
  XNOR U1682 ( .A(n1668), .B(n1503), .Z(n1670) );
  IV U1683 ( .A(p_input[9]), .Z(n1503) );
  XOR U1684 ( .A(n1672), .B(n1673), .Z(n1668) );
  AND U1685 ( .A(n1674), .B(n1675), .Z(n1673) );
  XNOR U1686 ( .A(p_input[24]), .B(n1672), .Z(n1675) );
  XNOR U1687 ( .A(n1672), .B(n1512), .Z(n1674) );
  IV U1688 ( .A(p_input[8]), .Z(n1512) );
  XOR U1689 ( .A(n1676), .B(n1677), .Z(n1672) );
  AND U1690 ( .A(n1678), .B(n1679), .Z(n1677) );
  XNOR U1691 ( .A(p_input[23]), .B(n1676), .Z(n1679) );
  XNOR U1692 ( .A(n1676), .B(n1521), .Z(n1678) );
  IV U1693 ( .A(p_input[7]), .Z(n1521) );
  XOR U1694 ( .A(n1680), .B(n1681), .Z(n1676) );
  AND U1695 ( .A(n1682), .B(n1683), .Z(n1681) );
  XNOR U1696 ( .A(p_input[22]), .B(n1680), .Z(n1683) );
  XNOR U1697 ( .A(n1680), .B(n1530), .Z(n1682) );
  IV U1698 ( .A(p_input[6]), .Z(n1530) );
  XOR U1699 ( .A(n1684), .B(n1685), .Z(n1680) );
  AND U1700 ( .A(n1686), .B(n1687), .Z(n1685) );
  XNOR U1701 ( .A(p_input[21]), .B(n1684), .Z(n1687) );
  XNOR U1702 ( .A(n1684), .B(n1539), .Z(n1686) );
  IV U1703 ( .A(p_input[5]), .Z(n1539) );
  XOR U1704 ( .A(n1688), .B(n1689), .Z(n1684) );
  AND U1705 ( .A(n1690), .B(n1691), .Z(n1689) );
  XNOR U1706 ( .A(p_input[20]), .B(n1688), .Z(n1691) );
  XNOR U1707 ( .A(n1688), .B(n1548), .Z(n1690) );
  IV U1708 ( .A(p_input[4]), .Z(n1548) );
  XOR U1709 ( .A(n1692), .B(n1693), .Z(n1688) );
  AND U1710 ( .A(n1694), .B(n1695), .Z(n1693) );
  XNOR U1711 ( .A(p_input[19]), .B(n1692), .Z(n1695) );
  XNOR U1712 ( .A(n1692), .B(n1557), .Z(n1694) );
  IV U1713 ( .A(p_input[3]), .Z(n1557) );
  XOR U1714 ( .A(n1696), .B(n1697), .Z(n1692) );
  AND U1715 ( .A(n1698), .B(n1699), .Z(n1697) );
  XNOR U1716 ( .A(p_input[18]), .B(n1696), .Z(n1699) );
  XNOR U1717 ( .A(n1696), .B(n1566), .Z(n1698) );
  IV U1718 ( .A(p_input[2]), .Z(n1566) );
  XNOR U1719 ( .A(n1700), .B(n1701), .Z(n1696) );
  AND U1720 ( .A(n1702), .B(n1703), .Z(n1701) );
  XOR U1721 ( .A(p_input[17]), .B(n1700), .Z(n1703) );
  XNOR U1722 ( .A(p_input[1]), .B(n1700), .Z(n1702) );
  AND U1723 ( .A(p_input[16]), .B(n1704), .Z(n1700) );
  IV U1724 ( .A(p_input[0]), .Z(n1704) );
endmodule

