
module knn_comb_BMR_W16_K2_N8 ( p_input, o );
  input [143:0] p_input;
  output [31:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][15] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992;
  assign \knn_comb_/min_val_out[0][0]  = p_input[112];
  assign \knn_comb_/min_val_out[0][1]  = p_input[113];
  assign \knn_comb_/min_val_out[0][2]  = p_input[114];
  assign \knn_comb_/min_val_out[0][3]  = p_input[115];
  assign \knn_comb_/min_val_out[0][4]  = p_input[116];
  assign \knn_comb_/min_val_out[0][5]  = p_input[117];
  assign \knn_comb_/min_val_out[0][6]  = p_input[118];
  assign \knn_comb_/min_val_out[0][7]  = p_input[119];
  assign \knn_comb_/min_val_out[0][8]  = p_input[120];
  assign \knn_comb_/min_val_out[0][9]  = p_input[121];
  assign \knn_comb_/min_val_out[0][10]  = p_input[122];
  assign \knn_comb_/min_val_out[0][11]  = p_input[123];
  assign \knn_comb_/min_val_out[0][12]  = p_input[124];
  assign \knn_comb_/min_val_out[0][13]  = p_input[125];
  assign \knn_comb_/min_val_out[0][14]  = p_input[126];
  assign \knn_comb_/min_val_out[0][15]  = p_input[127];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][0]  = p_input[96];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][1]  = p_input[97];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][2]  = p_input[98];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][3]  = p_input[99];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][4]  = p_input[100];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][5]  = p_input[101];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][6]  = p_input[102];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][7]  = p_input[103];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][8]  = p_input[104];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][9]  = p_input[105];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][10]  = p_input[106];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][11]  = p_input[107];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][12]  = p_input[108];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][13]  = p_input[109];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][14]  = p_input[110];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][15]  = p_input[111];

  XOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  XOR U2 ( .A(n3), .B(n4), .Z(o[8]) );
  XOR U3 ( .A(n5), .B(n6), .Z(o[7]) );
  XOR U4 ( .A(n7), .B(n8), .Z(o[6]) );
  XOR U5 ( .A(n9), .B(n10), .Z(o[5]) );
  XOR U6 ( .A(n11), .B(n12), .Z(o[4]) );
  XOR U7 ( .A(n13), .B(n14), .Z(o[3]) );
  XOR U8 ( .A(n15), .B(n16), .Z(o[31]) );
  XOR U9 ( .A(n17), .B(n18), .Z(o[30]) );
  XOR U10 ( .A(n19), .B(n20), .Z(o[2]) );
  XOR U11 ( .A(n21), .B(n22), .Z(o[29]) );
  XOR U12 ( .A(n23), .B(n24), .Z(o[28]) );
  XOR U13 ( .A(n25), .B(n26), .Z(o[27]) );
  XOR U14 ( .A(n27), .B(n28), .Z(o[26]) );
  XOR U15 ( .A(n1), .B(n29), .Z(o[25]) );
  AND U16 ( .A(n30), .B(n31), .Z(n1) );
  XOR U17 ( .A(n2), .B(n29), .Z(n31) );
  XOR U18 ( .A(n32), .B(n33), .Z(n29) );
  AND U19 ( .A(n34), .B(n35), .Z(n33) );
  XOR U20 ( .A(p_input[9]), .B(n32), .Z(n35) );
  XOR U21 ( .A(n36), .B(n37), .Z(n32) );
  AND U22 ( .A(n38), .B(n39), .Z(n37) );
  XOR U23 ( .A(n40), .B(n41), .Z(n2) );
  AND U24 ( .A(n42), .B(n39), .Z(n41) );
  XNOR U25 ( .A(n43), .B(n36), .Z(n39) );
  XOR U26 ( .A(n44), .B(n45), .Z(n36) );
  AND U27 ( .A(n46), .B(n47), .Z(n45) );
  XOR U28 ( .A(p_input[25]), .B(n44), .Z(n47) );
  XOR U29 ( .A(n48), .B(n49), .Z(n44) );
  AND U30 ( .A(n50), .B(n51), .Z(n49) );
  IV U31 ( .A(n40), .Z(n43) );
  XNOR U32 ( .A(n52), .B(n53), .Z(n40) );
  AND U33 ( .A(n54), .B(n51), .Z(n53) );
  XNOR U34 ( .A(n52), .B(n48), .Z(n51) );
  XOR U35 ( .A(n55), .B(n56), .Z(n48) );
  AND U36 ( .A(n57), .B(n58), .Z(n56) );
  XOR U37 ( .A(p_input[41]), .B(n55), .Z(n58) );
  XOR U38 ( .A(n59), .B(n60), .Z(n55) );
  AND U39 ( .A(n61), .B(n62), .Z(n60) );
  XOR U40 ( .A(n63), .B(n64), .Z(n52) );
  AND U41 ( .A(n65), .B(n62), .Z(n64) );
  XNOR U42 ( .A(n63), .B(n59), .Z(n62) );
  XOR U43 ( .A(n66), .B(n67), .Z(n59) );
  AND U44 ( .A(n68), .B(n69), .Z(n67) );
  XOR U45 ( .A(p_input[57]), .B(n66), .Z(n69) );
  XOR U46 ( .A(n70), .B(n71), .Z(n66) );
  AND U47 ( .A(n72), .B(n73), .Z(n71) );
  XOR U48 ( .A(n74), .B(n75), .Z(n63) );
  AND U49 ( .A(n76), .B(n73), .Z(n75) );
  XNOR U50 ( .A(n74), .B(n70), .Z(n73) );
  XOR U51 ( .A(n77), .B(n78), .Z(n70) );
  AND U52 ( .A(n79), .B(n80), .Z(n78) );
  XOR U53 ( .A(p_input[73]), .B(n77), .Z(n80) );
  XOR U54 ( .A(n81), .B(n82), .Z(n77) );
  AND U55 ( .A(n83), .B(n84), .Z(n82) );
  XOR U56 ( .A(n85), .B(n86), .Z(n74) );
  AND U57 ( .A(n87), .B(n84), .Z(n86) );
  XNOR U58 ( .A(n85), .B(n81), .Z(n84) );
  XOR U59 ( .A(n88), .B(n89), .Z(n81) );
  AND U60 ( .A(n90), .B(n91), .Z(n89) );
  XOR U61 ( .A(p_input[89]), .B(n88), .Z(n91) );
  XNOR U62 ( .A(n92), .B(n93), .Z(n88) );
  AND U63 ( .A(n94), .B(n95), .Z(n93) );
  XNOR U64 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n96), .Z(n85) );
  AND U65 ( .A(n97), .B(n95), .Z(n96) );
  XOR U66 ( .A(n98), .B(n92), .Z(n95) );
  XOR U67 ( .A(n3), .B(n99), .Z(o[24]) );
  AND U68 ( .A(n30), .B(n100), .Z(n3) );
  XOR U69 ( .A(n4), .B(n99), .Z(n100) );
  XOR U70 ( .A(n101), .B(n102), .Z(n99) );
  AND U71 ( .A(n34), .B(n103), .Z(n102) );
  XOR U72 ( .A(p_input[8]), .B(n101), .Z(n103) );
  XOR U73 ( .A(n104), .B(n105), .Z(n101) );
  AND U74 ( .A(n38), .B(n106), .Z(n105) );
  XOR U75 ( .A(n107), .B(n108), .Z(n4) );
  AND U76 ( .A(n42), .B(n106), .Z(n108) );
  XNOR U77 ( .A(n109), .B(n104), .Z(n106) );
  XOR U78 ( .A(n110), .B(n111), .Z(n104) );
  AND U79 ( .A(n46), .B(n112), .Z(n111) );
  XOR U80 ( .A(p_input[24]), .B(n110), .Z(n112) );
  XOR U81 ( .A(n113), .B(n114), .Z(n110) );
  AND U82 ( .A(n50), .B(n115), .Z(n114) );
  IV U83 ( .A(n107), .Z(n109) );
  XNOR U84 ( .A(n116), .B(n117), .Z(n107) );
  AND U85 ( .A(n54), .B(n115), .Z(n117) );
  XNOR U86 ( .A(n116), .B(n113), .Z(n115) );
  XOR U87 ( .A(n118), .B(n119), .Z(n113) );
  AND U88 ( .A(n57), .B(n120), .Z(n119) );
  XOR U89 ( .A(p_input[40]), .B(n118), .Z(n120) );
  XOR U90 ( .A(n121), .B(n122), .Z(n118) );
  AND U91 ( .A(n61), .B(n123), .Z(n122) );
  XOR U92 ( .A(n124), .B(n125), .Z(n116) );
  AND U93 ( .A(n65), .B(n123), .Z(n125) );
  XNOR U94 ( .A(n124), .B(n121), .Z(n123) );
  XOR U95 ( .A(n126), .B(n127), .Z(n121) );
  AND U96 ( .A(n68), .B(n128), .Z(n127) );
  XOR U97 ( .A(p_input[56]), .B(n126), .Z(n128) );
  XOR U98 ( .A(n129), .B(n130), .Z(n126) );
  AND U99 ( .A(n72), .B(n131), .Z(n130) );
  XOR U100 ( .A(n132), .B(n133), .Z(n124) );
  AND U101 ( .A(n76), .B(n131), .Z(n133) );
  XNOR U102 ( .A(n132), .B(n129), .Z(n131) );
  XOR U103 ( .A(n134), .B(n135), .Z(n129) );
  AND U104 ( .A(n79), .B(n136), .Z(n135) );
  XOR U105 ( .A(p_input[72]), .B(n134), .Z(n136) );
  XOR U106 ( .A(n137), .B(n138), .Z(n134) );
  AND U107 ( .A(n83), .B(n139), .Z(n138) );
  XOR U108 ( .A(n140), .B(n141), .Z(n132) );
  AND U109 ( .A(n87), .B(n139), .Z(n141) );
  XNOR U110 ( .A(n140), .B(n137), .Z(n139) );
  XOR U111 ( .A(n142), .B(n143), .Z(n137) );
  AND U112 ( .A(n90), .B(n144), .Z(n143) );
  XOR U113 ( .A(p_input[88]), .B(n142), .Z(n144) );
  XNOR U114 ( .A(n145), .B(n146), .Z(n142) );
  AND U115 ( .A(n94), .B(n147), .Z(n146) );
  XNOR U116 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n148), .Z(n140) );
  AND U117 ( .A(n97), .B(n147), .Z(n148) );
  XOR U118 ( .A(n149), .B(n145), .Z(n147) );
  XOR U119 ( .A(n5), .B(n150), .Z(o[23]) );
  AND U120 ( .A(n30), .B(n151), .Z(n5) );
  XOR U121 ( .A(n6), .B(n150), .Z(n151) );
  XOR U122 ( .A(n152), .B(n153), .Z(n150) );
  AND U123 ( .A(n34), .B(n154), .Z(n153) );
  XOR U124 ( .A(p_input[7]), .B(n152), .Z(n154) );
  XOR U125 ( .A(n155), .B(n156), .Z(n152) );
  AND U126 ( .A(n38), .B(n157), .Z(n156) );
  XOR U127 ( .A(n158), .B(n159), .Z(n6) );
  AND U128 ( .A(n42), .B(n157), .Z(n159) );
  XNOR U129 ( .A(n160), .B(n155), .Z(n157) );
  XOR U130 ( .A(n161), .B(n162), .Z(n155) );
  AND U131 ( .A(n46), .B(n163), .Z(n162) );
  XOR U132 ( .A(p_input[23]), .B(n161), .Z(n163) );
  XOR U133 ( .A(n164), .B(n165), .Z(n161) );
  AND U134 ( .A(n50), .B(n166), .Z(n165) );
  IV U135 ( .A(n158), .Z(n160) );
  XNOR U136 ( .A(n167), .B(n168), .Z(n158) );
  AND U137 ( .A(n54), .B(n166), .Z(n168) );
  XNOR U138 ( .A(n167), .B(n164), .Z(n166) );
  XOR U139 ( .A(n169), .B(n170), .Z(n164) );
  AND U140 ( .A(n57), .B(n171), .Z(n170) );
  XOR U141 ( .A(p_input[39]), .B(n169), .Z(n171) );
  XOR U142 ( .A(n172), .B(n173), .Z(n169) );
  AND U143 ( .A(n61), .B(n174), .Z(n173) );
  XOR U144 ( .A(n175), .B(n176), .Z(n167) );
  AND U145 ( .A(n65), .B(n174), .Z(n176) );
  XNOR U146 ( .A(n175), .B(n172), .Z(n174) );
  XOR U147 ( .A(n177), .B(n178), .Z(n172) );
  AND U148 ( .A(n68), .B(n179), .Z(n178) );
  XOR U149 ( .A(p_input[55]), .B(n177), .Z(n179) );
  XOR U150 ( .A(n180), .B(n181), .Z(n177) );
  AND U151 ( .A(n72), .B(n182), .Z(n181) );
  XOR U152 ( .A(n183), .B(n184), .Z(n175) );
  AND U153 ( .A(n76), .B(n182), .Z(n184) );
  XNOR U154 ( .A(n183), .B(n180), .Z(n182) );
  XOR U155 ( .A(n185), .B(n186), .Z(n180) );
  AND U156 ( .A(n79), .B(n187), .Z(n186) );
  XOR U157 ( .A(p_input[71]), .B(n185), .Z(n187) );
  XOR U158 ( .A(n188), .B(n189), .Z(n185) );
  AND U159 ( .A(n83), .B(n190), .Z(n189) );
  XOR U160 ( .A(n191), .B(n192), .Z(n183) );
  AND U161 ( .A(n87), .B(n190), .Z(n192) );
  XNOR U162 ( .A(n191), .B(n188), .Z(n190) );
  XOR U163 ( .A(n193), .B(n194), .Z(n188) );
  AND U164 ( .A(n90), .B(n195), .Z(n194) );
  XOR U165 ( .A(p_input[87]), .B(n193), .Z(n195) );
  XNOR U166 ( .A(n196), .B(n197), .Z(n193) );
  AND U167 ( .A(n94), .B(n198), .Z(n197) );
  XNOR U168 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n199), .Z(n191) );
  AND U169 ( .A(n97), .B(n198), .Z(n199) );
  XOR U170 ( .A(n200), .B(n196), .Z(n198) );
  IV U171 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .Z(n196) );
  IV U172 ( .A(\knn_comb_/min_val_out[0][7] ), .Z(n200) );
  XOR U173 ( .A(n7), .B(n201), .Z(o[22]) );
  AND U174 ( .A(n30), .B(n202), .Z(n7) );
  XOR U175 ( .A(n8), .B(n201), .Z(n202) );
  XOR U176 ( .A(n203), .B(n204), .Z(n201) );
  AND U177 ( .A(n34), .B(n205), .Z(n204) );
  XOR U178 ( .A(p_input[6]), .B(n203), .Z(n205) );
  XOR U179 ( .A(n206), .B(n207), .Z(n203) );
  AND U180 ( .A(n38), .B(n208), .Z(n207) );
  XOR U181 ( .A(n209), .B(n210), .Z(n8) );
  AND U182 ( .A(n42), .B(n208), .Z(n210) );
  XNOR U183 ( .A(n211), .B(n206), .Z(n208) );
  XOR U184 ( .A(n212), .B(n213), .Z(n206) );
  AND U185 ( .A(n46), .B(n214), .Z(n213) );
  XOR U186 ( .A(p_input[22]), .B(n212), .Z(n214) );
  XOR U187 ( .A(n215), .B(n216), .Z(n212) );
  AND U188 ( .A(n50), .B(n217), .Z(n216) );
  IV U189 ( .A(n209), .Z(n211) );
  XNOR U190 ( .A(n218), .B(n219), .Z(n209) );
  AND U191 ( .A(n54), .B(n217), .Z(n219) );
  XNOR U192 ( .A(n218), .B(n215), .Z(n217) );
  XOR U193 ( .A(n220), .B(n221), .Z(n215) );
  AND U194 ( .A(n57), .B(n222), .Z(n221) );
  XOR U195 ( .A(p_input[38]), .B(n220), .Z(n222) );
  XOR U196 ( .A(n223), .B(n224), .Z(n220) );
  AND U197 ( .A(n61), .B(n225), .Z(n224) );
  XOR U198 ( .A(n226), .B(n227), .Z(n218) );
  AND U199 ( .A(n65), .B(n225), .Z(n227) );
  XNOR U200 ( .A(n226), .B(n223), .Z(n225) );
  XOR U201 ( .A(n228), .B(n229), .Z(n223) );
  AND U202 ( .A(n68), .B(n230), .Z(n229) );
  XOR U203 ( .A(p_input[54]), .B(n228), .Z(n230) );
  XOR U204 ( .A(n231), .B(n232), .Z(n228) );
  AND U205 ( .A(n72), .B(n233), .Z(n232) );
  XOR U206 ( .A(n234), .B(n235), .Z(n226) );
  AND U207 ( .A(n76), .B(n233), .Z(n235) );
  XNOR U208 ( .A(n234), .B(n231), .Z(n233) );
  XOR U209 ( .A(n236), .B(n237), .Z(n231) );
  AND U210 ( .A(n79), .B(n238), .Z(n237) );
  XOR U211 ( .A(p_input[70]), .B(n236), .Z(n238) );
  XOR U212 ( .A(n239), .B(n240), .Z(n236) );
  AND U213 ( .A(n83), .B(n241), .Z(n240) );
  XOR U214 ( .A(n242), .B(n243), .Z(n234) );
  AND U215 ( .A(n87), .B(n241), .Z(n243) );
  XNOR U216 ( .A(n242), .B(n239), .Z(n241) );
  XOR U217 ( .A(n244), .B(n245), .Z(n239) );
  AND U218 ( .A(n90), .B(n246), .Z(n245) );
  XOR U219 ( .A(p_input[86]), .B(n244), .Z(n246) );
  XNOR U220 ( .A(n247), .B(n248), .Z(n244) );
  AND U221 ( .A(n94), .B(n249), .Z(n248) );
  XNOR U222 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n250), .Z(n242) );
  AND U223 ( .A(n97), .B(n249), .Z(n250) );
  XOR U224 ( .A(n251), .B(n247), .Z(n249) );
  IV U225 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .Z(n247) );
  XOR U226 ( .A(n9), .B(n252), .Z(o[21]) );
  AND U227 ( .A(n30), .B(n253), .Z(n9) );
  XOR U228 ( .A(n10), .B(n252), .Z(n253) );
  XOR U229 ( .A(n254), .B(n255), .Z(n252) );
  AND U230 ( .A(n34), .B(n256), .Z(n255) );
  XOR U231 ( .A(p_input[5]), .B(n254), .Z(n256) );
  XOR U232 ( .A(n257), .B(n258), .Z(n254) );
  AND U233 ( .A(n38), .B(n259), .Z(n258) );
  XOR U234 ( .A(n260), .B(n261), .Z(n10) );
  AND U235 ( .A(n42), .B(n259), .Z(n261) );
  XNOR U236 ( .A(n262), .B(n257), .Z(n259) );
  XOR U237 ( .A(n263), .B(n264), .Z(n257) );
  AND U238 ( .A(n46), .B(n265), .Z(n264) );
  XOR U239 ( .A(p_input[21]), .B(n263), .Z(n265) );
  XOR U240 ( .A(n266), .B(n267), .Z(n263) );
  AND U241 ( .A(n50), .B(n268), .Z(n267) );
  IV U242 ( .A(n260), .Z(n262) );
  XNOR U243 ( .A(n269), .B(n270), .Z(n260) );
  AND U244 ( .A(n54), .B(n268), .Z(n270) );
  XNOR U245 ( .A(n269), .B(n266), .Z(n268) );
  XOR U246 ( .A(n271), .B(n272), .Z(n266) );
  AND U247 ( .A(n57), .B(n273), .Z(n272) );
  XOR U248 ( .A(p_input[37]), .B(n271), .Z(n273) );
  XOR U249 ( .A(n274), .B(n275), .Z(n271) );
  AND U250 ( .A(n61), .B(n276), .Z(n275) );
  XOR U251 ( .A(n277), .B(n278), .Z(n269) );
  AND U252 ( .A(n65), .B(n276), .Z(n278) );
  XNOR U253 ( .A(n277), .B(n274), .Z(n276) );
  XOR U254 ( .A(n279), .B(n280), .Z(n274) );
  AND U255 ( .A(n68), .B(n281), .Z(n280) );
  XOR U256 ( .A(p_input[53]), .B(n279), .Z(n281) );
  XOR U257 ( .A(n282), .B(n283), .Z(n279) );
  AND U258 ( .A(n72), .B(n284), .Z(n283) );
  XOR U259 ( .A(n285), .B(n286), .Z(n277) );
  AND U260 ( .A(n76), .B(n284), .Z(n286) );
  XNOR U261 ( .A(n285), .B(n282), .Z(n284) );
  XOR U262 ( .A(n287), .B(n288), .Z(n282) );
  AND U263 ( .A(n79), .B(n289), .Z(n288) );
  XOR U264 ( .A(p_input[69]), .B(n287), .Z(n289) );
  XOR U265 ( .A(n290), .B(n291), .Z(n287) );
  AND U266 ( .A(n83), .B(n292), .Z(n291) );
  XOR U267 ( .A(n293), .B(n294), .Z(n285) );
  AND U268 ( .A(n87), .B(n292), .Z(n294) );
  XNOR U269 ( .A(n293), .B(n290), .Z(n292) );
  XOR U270 ( .A(n295), .B(n296), .Z(n290) );
  AND U271 ( .A(n90), .B(n297), .Z(n296) );
  XOR U272 ( .A(p_input[85]), .B(n295), .Z(n297) );
  XNOR U273 ( .A(n298), .B(n299), .Z(n295) );
  AND U274 ( .A(n94), .B(n300), .Z(n299) );
  XNOR U275 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n301), .Z(n293) );
  AND U276 ( .A(n97), .B(n300), .Z(n301) );
  XOR U277 ( .A(n302), .B(n298), .Z(n300) );
  IV U278 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .Z(n298) );
  XOR U279 ( .A(n11), .B(n303), .Z(o[20]) );
  AND U280 ( .A(n30), .B(n304), .Z(n11) );
  XOR U281 ( .A(n12), .B(n303), .Z(n304) );
  XOR U282 ( .A(n305), .B(n306), .Z(n303) );
  AND U283 ( .A(n34), .B(n307), .Z(n306) );
  XOR U284 ( .A(p_input[4]), .B(n305), .Z(n307) );
  XOR U285 ( .A(n308), .B(n309), .Z(n305) );
  AND U286 ( .A(n38), .B(n310), .Z(n309) );
  XOR U287 ( .A(n311), .B(n312), .Z(n12) );
  AND U288 ( .A(n42), .B(n310), .Z(n312) );
  XNOR U289 ( .A(n313), .B(n308), .Z(n310) );
  XOR U290 ( .A(n314), .B(n315), .Z(n308) );
  AND U291 ( .A(n46), .B(n316), .Z(n315) );
  XOR U292 ( .A(p_input[20]), .B(n314), .Z(n316) );
  XOR U293 ( .A(n317), .B(n318), .Z(n314) );
  AND U294 ( .A(n50), .B(n319), .Z(n318) );
  IV U295 ( .A(n311), .Z(n313) );
  XNOR U296 ( .A(n320), .B(n321), .Z(n311) );
  AND U297 ( .A(n54), .B(n319), .Z(n321) );
  XNOR U298 ( .A(n320), .B(n317), .Z(n319) );
  XOR U299 ( .A(n322), .B(n323), .Z(n317) );
  AND U300 ( .A(n57), .B(n324), .Z(n323) );
  XOR U301 ( .A(p_input[36]), .B(n322), .Z(n324) );
  XOR U302 ( .A(n325), .B(n326), .Z(n322) );
  AND U303 ( .A(n61), .B(n327), .Z(n326) );
  XOR U304 ( .A(n328), .B(n329), .Z(n320) );
  AND U305 ( .A(n65), .B(n327), .Z(n329) );
  XNOR U306 ( .A(n328), .B(n325), .Z(n327) );
  XOR U307 ( .A(n330), .B(n331), .Z(n325) );
  AND U308 ( .A(n68), .B(n332), .Z(n331) );
  XOR U309 ( .A(p_input[52]), .B(n330), .Z(n332) );
  XOR U310 ( .A(n333), .B(n334), .Z(n330) );
  AND U311 ( .A(n72), .B(n335), .Z(n334) );
  XOR U312 ( .A(n336), .B(n337), .Z(n328) );
  AND U313 ( .A(n76), .B(n335), .Z(n337) );
  XNOR U314 ( .A(n336), .B(n333), .Z(n335) );
  XOR U315 ( .A(n338), .B(n339), .Z(n333) );
  AND U316 ( .A(n79), .B(n340), .Z(n339) );
  XOR U317 ( .A(p_input[68]), .B(n338), .Z(n340) );
  XOR U318 ( .A(n341), .B(n342), .Z(n338) );
  AND U319 ( .A(n83), .B(n343), .Z(n342) );
  XOR U320 ( .A(n344), .B(n345), .Z(n336) );
  AND U321 ( .A(n87), .B(n343), .Z(n345) );
  XNOR U322 ( .A(n344), .B(n341), .Z(n343) );
  XOR U323 ( .A(n346), .B(n347), .Z(n341) );
  AND U324 ( .A(n90), .B(n348), .Z(n347) );
  XOR U325 ( .A(p_input[84]), .B(n346), .Z(n348) );
  XNOR U326 ( .A(n349), .B(n350), .Z(n346) );
  AND U327 ( .A(n94), .B(n351), .Z(n350) );
  XNOR U328 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n352), .Z(n344) );
  AND U329 ( .A(n97), .B(n351), .Z(n352) );
  XOR U330 ( .A(n353), .B(n349), .Z(n351) );
  IV U331 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .Z(n349) );
  IV U332 ( .A(\knn_comb_/min_val_out[0][4] ), .Z(n353) );
  XOR U333 ( .A(n354), .B(n355), .Z(o[1]) );
  XOR U334 ( .A(n13), .B(n356), .Z(o[19]) );
  AND U335 ( .A(n30), .B(n357), .Z(n13) );
  XOR U336 ( .A(n14), .B(n356), .Z(n357) );
  XOR U337 ( .A(n358), .B(n359), .Z(n356) );
  AND U338 ( .A(n34), .B(n360), .Z(n359) );
  XOR U339 ( .A(p_input[3]), .B(n358), .Z(n360) );
  XOR U340 ( .A(n361), .B(n362), .Z(n358) );
  AND U341 ( .A(n38), .B(n363), .Z(n362) );
  XOR U342 ( .A(n364), .B(n365), .Z(n14) );
  AND U343 ( .A(n42), .B(n363), .Z(n365) );
  XNOR U344 ( .A(n366), .B(n361), .Z(n363) );
  XOR U345 ( .A(n367), .B(n368), .Z(n361) );
  AND U346 ( .A(n46), .B(n369), .Z(n368) );
  XOR U347 ( .A(p_input[19]), .B(n367), .Z(n369) );
  XOR U348 ( .A(n370), .B(n371), .Z(n367) );
  AND U349 ( .A(n50), .B(n372), .Z(n371) );
  IV U350 ( .A(n364), .Z(n366) );
  XNOR U351 ( .A(n373), .B(n374), .Z(n364) );
  AND U352 ( .A(n54), .B(n372), .Z(n374) );
  XNOR U353 ( .A(n373), .B(n370), .Z(n372) );
  XOR U354 ( .A(n375), .B(n376), .Z(n370) );
  AND U355 ( .A(n57), .B(n377), .Z(n376) );
  XOR U356 ( .A(p_input[35]), .B(n375), .Z(n377) );
  XOR U357 ( .A(n378), .B(n379), .Z(n375) );
  AND U358 ( .A(n61), .B(n380), .Z(n379) );
  XOR U359 ( .A(n381), .B(n382), .Z(n373) );
  AND U360 ( .A(n65), .B(n380), .Z(n382) );
  XNOR U361 ( .A(n381), .B(n378), .Z(n380) );
  XOR U362 ( .A(n383), .B(n384), .Z(n378) );
  AND U363 ( .A(n68), .B(n385), .Z(n384) );
  XOR U364 ( .A(p_input[51]), .B(n383), .Z(n385) );
  XOR U365 ( .A(n386), .B(n387), .Z(n383) );
  AND U366 ( .A(n72), .B(n388), .Z(n387) );
  XOR U367 ( .A(n389), .B(n390), .Z(n381) );
  AND U368 ( .A(n76), .B(n388), .Z(n390) );
  XNOR U369 ( .A(n389), .B(n386), .Z(n388) );
  XOR U370 ( .A(n391), .B(n392), .Z(n386) );
  AND U371 ( .A(n79), .B(n393), .Z(n392) );
  XOR U372 ( .A(p_input[67]), .B(n391), .Z(n393) );
  XOR U373 ( .A(n394), .B(n395), .Z(n391) );
  AND U374 ( .A(n83), .B(n396), .Z(n395) );
  XOR U375 ( .A(n397), .B(n398), .Z(n389) );
  AND U376 ( .A(n87), .B(n396), .Z(n398) );
  XNOR U377 ( .A(n397), .B(n394), .Z(n396) );
  XOR U378 ( .A(n399), .B(n400), .Z(n394) );
  AND U379 ( .A(n90), .B(n401), .Z(n400) );
  XOR U380 ( .A(p_input[83]), .B(n399), .Z(n401) );
  XNOR U381 ( .A(n402), .B(n403), .Z(n399) );
  AND U382 ( .A(n94), .B(n404), .Z(n403) );
  XNOR U383 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n405), .Z(n397) );
  AND U384 ( .A(n97), .B(n404), .Z(n405) );
  XOR U385 ( .A(n406), .B(n402), .Z(n404) );
  IV U386 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .Z(n402) );
  XOR U387 ( .A(n19), .B(n407), .Z(o[18]) );
  AND U388 ( .A(n30), .B(n408), .Z(n19) );
  XOR U389 ( .A(n20), .B(n407), .Z(n408) );
  XOR U390 ( .A(n409), .B(n410), .Z(n407) );
  AND U391 ( .A(n34), .B(n411), .Z(n410) );
  XOR U392 ( .A(p_input[2]), .B(n409), .Z(n411) );
  XOR U393 ( .A(n412), .B(n413), .Z(n409) );
  AND U394 ( .A(n38), .B(n414), .Z(n413) );
  XOR U395 ( .A(n415), .B(n416), .Z(n20) );
  AND U396 ( .A(n42), .B(n414), .Z(n416) );
  XNOR U397 ( .A(n417), .B(n412), .Z(n414) );
  XOR U398 ( .A(n418), .B(n419), .Z(n412) );
  AND U399 ( .A(n46), .B(n420), .Z(n419) );
  XOR U400 ( .A(p_input[18]), .B(n418), .Z(n420) );
  XOR U401 ( .A(n421), .B(n422), .Z(n418) );
  AND U402 ( .A(n50), .B(n423), .Z(n422) );
  IV U403 ( .A(n415), .Z(n417) );
  XNOR U404 ( .A(n424), .B(n425), .Z(n415) );
  AND U405 ( .A(n54), .B(n423), .Z(n425) );
  XNOR U406 ( .A(n424), .B(n421), .Z(n423) );
  XOR U407 ( .A(n426), .B(n427), .Z(n421) );
  AND U408 ( .A(n57), .B(n428), .Z(n427) );
  XOR U409 ( .A(p_input[34]), .B(n426), .Z(n428) );
  XOR U410 ( .A(n429), .B(n430), .Z(n426) );
  AND U411 ( .A(n61), .B(n431), .Z(n430) );
  XOR U412 ( .A(n432), .B(n433), .Z(n424) );
  AND U413 ( .A(n65), .B(n431), .Z(n433) );
  XNOR U414 ( .A(n432), .B(n429), .Z(n431) );
  XOR U415 ( .A(n434), .B(n435), .Z(n429) );
  AND U416 ( .A(n68), .B(n436), .Z(n435) );
  XOR U417 ( .A(p_input[50]), .B(n434), .Z(n436) );
  XOR U418 ( .A(n437), .B(n438), .Z(n434) );
  AND U419 ( .A(n72), .B(n439), .Z(n438) );
  XOR U420 ( .A(n440), .B(n441), .Z(n432) );
  AND U421 ( .A(n76), .B(n439), .Z(n441) );
  XNOR U422 ( .A(n440), .B(n437), .Z(n439) );
  XOR U423 ( .A(n442), .B(n443), .Z(n437) );
  AND U424 ( .A(n79), .B(n444), .Z(n443) );
  XOR U425 ( .A(p_input[66]), .B(n442), .Z(n444) );
  XOR U426 ( .A(n445), .B(n446), .Z(n442) );
  AND U427 ( .A(n83), .B(n447), .Z(n446) );
  XOR U428 ( .A(n448), .B(n449), .Z(n440) );
  AND U429 ( .A(n87), .B(n447), .Z(n449) );
  XNOR U430 ( .A(n448), .B(n445), .Z(n447) );
  XOR U431 ( .A(n450), .B(n451), .Z(n445) );
  AND U432 ( .A(n90), .B(n452), .Z(n451) );
  XOR U433 ( .A(p_input[82]), .B(n450), .Z(n452) );
  XNOR U434 ( .A(n453), .B(n454), .Z(n450) );
  AND U435 ( .A(n94), .B(n455), .Z(n454) );
  XNOR U436 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n456), .Z(n448) );
  AND U437 ( .A(n97), .B(n455), .Z(n456) );
  XOR U438 ( .A(n457), .B(n453), .Z(n455) );
  XOR U439 ( .A(n354), .B(n458), .Z(o[17]) );
  AND U440 ( .A(n30), .B(n459), .Z(n354) );
  XOR U441 ( .A(n355), .B(n458), .Z(n459) );
  XOR U442 ( .A(n460), .B(n461), .Z(n458) );
  AND U443 ( .A(n34), .B(n462), .Z(n461) );
  XOR U444 ( .A(p_input[1]), .B(n460), .Z(n462) );
  XOR U445 ( .A(n463), .B(n464), .Z(n460) );
  AND U446 ( .A(n38), .B(n465), .Z(n464) );
  XOR U447 ( .A(n466), .B(n467), .Z(n355) );
  AND U448 ( .A(n42), .B(n465), .Z(n467) );
  XNOR U449 ( .A(n468), .B(n463), .Z(n465) );
  XOR U450 ( .A(n469), .B(n470), .Z(n463) );
  AND U451 ( .A(n46), .B(n471), .Z(n470) );
  XOR U452 ( .A(p_input[17]), .B(n469), .Z(n471) );
  XOR U453 ( .A(n472), .B(n473), .Z(n469) );
  AND U454 ( .A(n50), .B(n474), .Z(n473) );
  IV U455 ( .A(n466), .Z(n468) );
  XNOR U456 ( .A(n475), .B(n476), .Z(n466) );
  AND U457 ( .A(n54), .B(n474), .Z(n476) );
  XNOR U458 ( .A(n475), .B(n472), .Z(n474) );
  XOR U459 ( .A(n477), .B(n478), .Z(n472) );
  AND U460 ( .A(n57), .B(n479), .Z(n478) );
  XOR U461 ( .A(p_input[33]), .B(n477), .Z(n479) );
  XOR U462 ( .A(n480), .B(n481), .Z(n477) );
  AND U463 ( .A(n61), .B(n482), .Z(n481) );
  XOR U464 ( .A(n483), .B(n484), .Z(n475) );
  AND U465 ( .A(n65), .B(n482), .Z(n484) );
  XNOR U466 ( .A(n483), .B(n480), .Z(n482) );
  XOR U467 ( .A(n485), .B(n486), .Z(n480) );
  AND U468 ( .A(n68), .B(n487), .Z(n486) );
  XOR U469 ( .A(p_input[49]), .B(n485), .Z(n487) );
  XOR U470 ( .A(n488), .B(n489), .Z(n485) );
  AND U471 ( .A(n72), .B(n490), .Z(n489) );
  XOR U472 ( .A(n491), .B(n492), .Z(n483) );
  AND U473 ( .A(n76), .B(n490), .Z(n492) );
  XNOR U474 ( .A(n491), .B(n488), .Z(n490) );
  XOR U475 ( .A(n493), .B(n494), .Z(n488) );
  AND U476 ( .A(n79), .B(n495), .Z(n494) );
  XOR U477 ( .A(p_input[65]), .B(n493), .Z(n495) );
  XOR U478 ( .A(n496), .B(n497), .Z(n493) );
  AND U479 ( .A(n83), .B(n498), .Z(n497) );
  XOR U480 ( .A(n499), .B(n500), .Z(n491) );
  AND U481 ( .A(n87), .B(n498), .Z(n500) );
  XNOR U482 ( .A(n499), .B(n496), .Z(n498) );
  XOR U483 ( .A(n501), .B(n502), .Z(n496) );
  AND U484 ( .A(n90), .B(n503), .Z(n502) );
  XOR U485 ( .A(p_input[81]), .B(n501), .Z(n503) );
  XNOR U486 ( .A(n504), .B(n505), .Z(n501) );
  AND U487 ( .A(n94), .B(n506), .Z(n505) );
  XNOR U488 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n507), .Z(n499) );
  AND U489 ( .A(n97), .B(n506), .Z(n507) );
  XOR U490 ( .A(n508), .B(n504), .Z(n506) );
  IV U491 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n504) );
  XOR U492 ( .A(n509), .B(n510), .Z(o[16]) );
  XOR U493 ( .A(n15), .B(n511), .Z(o[15]) );
  AND U494 ( .A(n30), .B(n512), .Z(n15) );
  XOR U495 ( .A(n16), .B(n511), .Z(n512) );
  XOR U496 ( .A(n513), .B(n514), .Z(n511) );
  AND U497 ( .A(n42), .B(n515), .Z(n514) );
  XOR U498 ( .A(n516), .B(n517), .Z(n16) );
  AND U499 ( .A(n34), .B(n518), .Z(n517) );
  XOR U500 ( .A(p_input[15]), .B(n516), .Z(n518) );
  XNOR U501 ( .A(n519), .B(n520), .Z(n516) );
  AND U502 ( .A(n38), .B(n515), .Z(n520) );
  XNOR U503 ( .A(n519), .B(n513), .Z(n515) );
  XOR U504 ( .A(n521), .B(n522), .Z(n513) );
  AND U505 ( .A(n54), .B(n523), .Z(n522) );
  XNOR U506 ( .A(n524), .B(n525), .Z(n519) );
  AND U507 ( .A(n46), .B(n526), .Z(n525) );
  XOR U508 ( .A(p_input[31]), .B(n524), .Z(n526) );
  XNOR U509 ( .A(n527), .B(n528), .Z(n524) );
  AND U510 ( .A(n50), .B(n523), .Z(n528) );
  XNOR U511 ( .A(n527), .B(n521), .Z(n523) );
  XOR U512 ( .A(n529), .B(n530), .Z(n521) );
  AND U513 ( .A(n65), .B(n531), .Z(n530) );
  XNOR U514 ( .A(n532), .B(n533), .Z(n527) );
  AND U515 ( .A(n57), .B(n534), .Z(n533) );
  XOR U516 ( .A(p_input[47]), .B(n532), .Z(n534) );
  XNOR U517 ( .A(n535), .B(n536), .Z(n532) );
  AND U518 ( .A(n61), .B(n531), .Z(n536) );
  XNOR U519 ( .A(n535), .B(n529), .Z(n531) );
  XOR U520 ( .A(n537), .B(n538), .Z(n529) );
  AND U521 ( .A(n76), .B(n539), .Z(n538) );
  XNOR U522 ( .A(n540), .B(n541), .Z(n535) );
  AND U523 ( .A(n68), .B(n542), .Z(n541) );
  XOR U524 ( .A(p_input[63]), .B(n540), .Z(n542) );
  XNOR U525 ( .A(n543), .B(n544), .Z(n540) );
  AND U526 ( .A(n72), .B(n539), .Z(n544) );
  XNOR U527 ( .A(n543), .B(n537), .Z(n539) );
  XOR U528 ( .A(n545), .B(n546), .Z(n537) );
  AND U529 ( .A(n87), .B(n547), .Z(n546) );
  XNOR U530 ( .A(n548), .B(n549), .Z(n543) );
  AND U531 ( .A(n79), .B(n550), .Z(n549) );
  XOR U532 ( .A(p_input[79]), .B(n548), .Z(n550) );
  XNOR U533 ( .A(n551), .B(n552), .Z(n548) );
  AND U534 ( .A(n83), .B(n547), .Z(n552) );
  XNOR U535 ( .A(n551), .B(n545), .Z(n547) );
  XOR U536 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n553), .Z(n545) );
  AND U537 ( .A(n97), .B(n554), .Z(n553) );
  XNOR U538 ( .A(n555), .B(n556), .Z(n551) );
  AND U539 ( .A(n90), .B(n557), .Z(n556) );
  XOR U540 ( .A(p_input[95]), .B(n555), .Z(n557) );
  XNOR U541 ( .A(n558), .B(n559), .Z(n555) );
  AND U542 ( .A(n94), .B(n554), .Z(n559) );
  XOR U543 ( .A(n560), .B(n558), .Z(n554) );
  IV U544 ( .A(\knn_comb_/min_val_out[0][15] ), .Z(n560) );
  XOR U545 ( .A(n17), .B(n561), .Z(o[14]) );
  AND U546 ( .A(n30), .B(n562), .Z(n17) );
  XOR U547 ( .A(n18), .B(n561), .Z(n562) );
  XOR U548 ( .A(n563), .B(n564), .Z(n561) );
  AND U549 ( .A(n42), .B(n565), .Z(n564) );
  XOR U550 ( .A(n566), .B(n567), .Z(n18) );
  AND U551 ( .A(n34), .B(n568), .Z(n567) );
  XOR U552 ( .A(p_input[14]), .B(n566), .Z(n568) );
  XNOR U553 ( .A(n569), .B(n570), .Z(n566) );
  AND U554 ( .A(n38), .B(n565), .Z(n570) );
  XNOR U555 ( .A(n569), .B(n563), .Z(n565) );
  XOR U556 ( .A(n571), .B(n572), .Z(n563) );
  AND U557 ( .A(n54), .B(n573), .Z(n572) );
  XNOR U558 ( .A(n574), .B(n575), .Z(n569) );
  AND U559 ( .A(n46), .B(n576), .Z(n575) );
  XOR U560 ( .A(p_input[30]), .B(n574), .Z(n576) );
  XNOR U561 ( .A(n577), .B(n578), .Z(n574) );
  AND U562 ( .A(n50), .B(n573), .Z(n578) );
  XNOR U563 ( .A(n577), .B(n571), .Z(n573) );
  XOR U564 ( .A(n579), .B(n580), .Z(n571) );
  AND U565 ( .A(n65), .B(n581), .Z(n580) );
  XNOR U566 ( .A(n582), .B(n583), .Z(n577) );
  AND U567 ( .A(n57), .B(n584), .Z(n583) );
  XOR U568 ( .A(p_input[46]), .B(n582), .Z(n584) );
  XNOR U569 ( .A(n585), .B(n586), .Z(n582) );
  AND U570 ( .A(n61), .B(n581), .Z(n586) );
  XNOR U571 ( .A(n585), .B(n579), .Z(n581) );
  XOR U572 ( .A(n587), .B(n588), .Z(n579) );
  AND U573 ( .A(n76), .B(n589), .Z(n588) );
  XNOR U574 ( .A(n590), .B(n591), .Z(n585) );
  AND U575 ( .A(n68), .B(n592), .Z(n591) );
  XOR U576 ( .A(p_input[62]), .B(n590), .Z(n592) );
  XNOR U577 ( .A(n593), .B(n594), .Z(n590) );
  AND U578 ( .A(n72), .B(n589), .Z(n594) );
  XNOR U579 ( .A(n593), .B(n587), .Z(n589) );
  XOR U580 ( .A(n595), .B(n596), .Z(n587) );
  AND U581 ( .A(n87), .B(n597), .Z(n596) );
  XNOR U582 ( .A(n598), .B(n599), .Z(n593) );
  AND U583 ( .A(n79), .B(n600), .Z(n599) );
  XOR U584 ( .A(p_input[78]), .B(n598), .Z(n600) );
  XNOR U585 ( .A(n601), .B(n602), .Z(n598) );
  AND U586 ( .A(n83), .B(n597), .Z(n602) );
  XNOR U587 ( .A(n601), .B(n595), .Z(n597) );
  XOR U588 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n603), .Z(n595) );
  AND U589 ( .A(n97), .B(n604), .Z(n603) );
  XNOR U590 ( .A(n605), .B(n606), .Z(n601) );
  AND U591 ( .A(n90), .B(n607), .Z(n606) );
  XOR U592 ( .A(p_input[94]), .B(n605), .Z(n607) );
  XNOR U593 ( .A(n608), .B(n609), .Z(n605) );
  AND U594 ( .A(n94), .B(n604), .Z(n609) );
  XOR U595 ( .A(n610), .B(n608), .Z(n604) );
  IV U596 ( .A(\knn_comb_/min_val_out[0][14] ), .Z(n610) );
  IV U597 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n608) );
  XOR U598 ( .A(n21), .B(n611), .Z(o[13]) );
  AND U599 ( .A(n30), .B(n612), .Z(n21) );
  XOR U600 ( .A(n22), .B(n611), .Z(n612) );
  XOR U601 ( .A(n613), .B(n614), .Z(n611) );
  AND U602 ( .A(n42), .B(n615), .Z(n614) );
  XOR U603 ( .A(n616), .B(n617), .Z(n22) );
  AND U604 ( .A(n34), .B(n618), .Z(n617) );
  XOR U605 ( .A(p_input[13]), .B(n616), .Z(n618) );
  XNOR U606 ( .A(n619), .B(n620), .Z(n616) );
  AND U607 ( .A(n38), .B(n615), .Z(n620) );
  XNOR U608 ( .A(n619), .B(n613), .Z(n615) );
  XOR U609 ( .A(n621), .B(n622), .Z(n613) );
  AND U610 ( .A(n54), .B(n623), .Z(n622) );
  XNOR U611 ( .A(n624), .B(n625), .Z(n619) );
  AND U612 ( .A(n46), .B(n626), .Z(n625) );
  XOR U613 ( .A(p_input[29]), .B(n624), .Z(n626) );
  XNOR U614 ( .A(n627), .B(n628), .Z(n624) );
  AND U615 ( .A(n50), .B(n623), .Z(n628) );
  XNOR U616 ( .A(n627), .B(n621), .Z(n623) );
  XOR U617 ( .A(n629), .B(n630), .Z(n621) );
  AND U618 ( .A(n65), .B(n631), .Z(n630) );
  XNOR U619 ( .A(n632), .B(n633), .Z(n627) );
  AND U620 ( .A(n57), .B(n634), .Z(n633) );
  XOR U621 ( .A(p_input[45]), .B(n632), .Z(n634) );
  XNOR U622 ( .A(n635), .B(n636), .Z(n632) );
  AND U623 ( .A(n61), .B(n631), .Z(n636) );
  XNOR U624 ( .A(n635), .B(n629), .Z(n631) );
  XOR U625 ( .A(n637), .B(n638), .Z(n629) );
  AND U626 ( .A(n76), .B(n639), .Z(n638) );
  XNOR U627 ( .A(n640), .B(n641), .Z(n635) );
  AND U628 ( .A(n68), .B(n642), .Z(n641) );
  XOR U629 ( .A(p_input[61]), .B(n640), .Z(n642) );
  XNOR U630 ( .A(n643), .B(n644), .Z(n640) );
  AND U631 ( .A(n72), .B(n639), .Z(n644) );
  XNOR U632 ( .A(n643), .B(n637), .Z(n639) );
  XOR U633 ( .A(n645), .B(n646), .Z(n637) );
  AND U634 ( .A(n87), .B(n647), .Z(n646) );
  XNOR U635 ( .A(n648), .B(n649), .Z(n643) );
  AND U636 ( .A(n79), .B(n650), .Z(n649) );
  XOR U637 ( .A(p_input[77]), .B(n648), .Z(n650) );
  XNOR U638 ( .A(n651), .B(n652), .Z(n648) );
  AND U639 ( .A(n83), .B(n647), .Z(n652) );
  XNOR U640 ( .A(n651), .B(n645), .Z(n647) );
  XOR U641 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n653), .Z(n645) );
  AND U642 ( .A(n97), .B(n654), .Z(n653) );
  XNOR U643 ( .A(n655), .B(n656), .Z(n651) );
  AND U644 ( .A(n90), .B(n657), .Z(n656) );
  XOR U645 ( .A(p_input[93]), .B(n655), .Z(n657) );
  XNOR U646 ( .A(n658), .B(n659), .Z(n655) );
  AND U647 ( .A(n94), .B(n654), .Z(n659) );
  XOR U648 ( .A(\knn_comb_/min_val_out[0][13] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n654) );
  XOR U649 ( .A(n23), .B(n660), .Z(o[12]) );
  AND U650 ( .A(n30), .B(n661), .Z(n23) );
  XOR U651 ( .A(n24), .B(n660), .Z(n661) );
  XOR U652 ( .A(n662), .B(n663), .Z(n660) );
  AND U653 ( .A(n42), .B(n664), .Z(n663) );
  XOR U654 ( .A(n665), .B(n666), .Z(n24) );
  AND U655 ( .A(n34), .B(n667), .Z(n666) );
  XOR U656 ( .A(p_input[12]), .B(n665), .Z(n667) );
  XNOR U657 ( .A(n668), .B(n669), .Z(n665) );
  AND U658 ( .A(n38), .B(n664), .Z(n669) );
  XNOR U659 ( .A(n668), .B(n662), .Z(n664) );
  XOR U660 ( .A(n670), .B(n671), .Z(n662) );
  AND U661 ( .A(n54), .B(n672), .Z(n671) );
  XNOR U662 ( .A(n673), .B(n674), .Z(n668) );
  AND U663 ( .A(n46), .B(n675), .Z(n674) );
  XOR U664 ( .A(p_input[28]), .B(n673), .Z(n675) );
  XNOR U665 ( .A(n676), .B(n677), .Z(n673) );
  AND U666 ( .A(n50), .B(n672), .Z(n677) );
  XNOR U667 ( .A(n676), .B(n670), .Z(n672) );
  XOR U668 ( .A(n678), .B(n679), .Z(n670) );
  AND U669 ( .A(n65), .B(n680), .Z(n679) );
  XNOR U670 ( .A(n681), .B(n682), .Z(n676) );
  AND U671 ( .A(n57), .B(n683), .Z(n682) );
  XOR U672 ( .A(p_input[44]), .B(n681), .Z(n683) );
  XNOR U673 ( .A(n684), .B(n685), .Z(n681) );
  AND U674 ( .A(n61), .B(n680), .Z(n685) );
  XNOR U675 ( .A(n684), .B(n678), .Z(n680) );
  XOR U676 ( .A(n686), .B(n687), .Z(n678) );
  AND U677 ( .A(n76), .B(n688), .Z(n687) );
  XNOR U678 ( .A(n689), .B(n690), .Z(n684) );
  AND U679 ( .A(n68), .B(n691), .Z(n690) );
  XOR U680 ( .A(p_input[60]), .B(n689), .Z(n691) );
  XNOR U681 ( .A(n692), .B(n693), .Z(n689) );
  AND U682 ( .A(n72), .B(n688), .Z(n693) );
  XNOR U683 ( .A(n692), .B(n686), .Z(n688) );
  XOR U684 ( .A(n694), .B(n695), .Z(n686) );
  AND U685 ( .A(n87), .B(n696), .Z(n695) );
  XNOR U686 ( .A(n697), .B(n698), .Z(n692) );
  AND U687 ( .A(n79), .B(n699), .Z(n698) );
  XOR U688 ( .A(p_input[76]), .B(n697), .Z(n699) );
  XNOR U689 ( .A(n700), .B(n701), .Z(n697) );
  AND U690 ( .A(n83), .B(n696), .Z(n701) );
  XNOR U691 ( .A(n700), .B(n694), .Z(n696) );
  XOR U692 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n702), .Z(n694) );
  AND U693 ( .A(n97), .B(n703), .Z(n702) );
  XNOR U694 ( .A(n704), .B(n705), .Z(n700) );
  AND U695 ( .A(n90), .B(n706), .Z(n705) );
  XOR U696 ( .A(p_input[92]), .B(n704), .Z(n706) );
  XNOR U697 ( .A(n707), .B(n708), .Z(n704) );
  AND U698 ( .A(n94), .B(n703), .Z(n708) );
  XOR U699 ( .A(\knn_comb_/min_val_out[0][12] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n703) );
  XOR U700 ( .A(n25), .B(n709), .Z(o[11]) );
  AND U701 ( .A(n30), .B(n710), .Z(n25) );
  XOR U702 ( .A(n26), .B(n709), .Z(n710) );
  XOR U703 ( .A(n711), .B(n712), .Z(n709) );
  AND U704 ( .A(n42), .B(n713), .Z(n712) );
  XOR U705 ( .A(n714), .B(n715), .Z(n26) );
  AND U706 ( .A(n34), .B(n716), .Z(n715) );
  XOR U707 ( .A(p_input[11]), .B(n714), .Z(n716) );
  XNOR U708 ( .A(n717), .B(n718), .Z(n714) );
  AND U709 ( .A(n38), .B(n713), .Z(n718) );
  XNOR U710 ( .A(n717), .B(n711), .Z(n713) );
  XOR U711 ( .A(n719), .B(n720), .Z(n711) );
  AND U712 ( .A(n54), .B(n721), .Z(n720) );
  XNOR U713 ( .A(n722), .B(n723), .Z(n717) );
  AND U714 ( .A(n46), .B(n724), .Z(n723) );
  XOR U715 ( .A(p_input[27]), .B(n722), .Z(n724) );
  XNOR U716 ( .A(n725), .B(n726), .Z(n722) );
  AND U717 ( .A(n50), .B(n721), .Z(n726) );
  XNOR U718 ( .A(n725), .B(n719), .Z(n721) );
  XOR U719 ( .A(n727), .B(n728), .Z(n719) );
  AND U720 ( .A(n65), .B(n729), .Z(n728) );
  XNOR U721 ( .A(n730), .B(n731), .Z(n725) );
  AND U722 ( .A(n57), .B(n732), .Z(n731) );
  XOR U723 ( .A(p_input[43]), .B(n730), .Z(n732) );
  XNOR U724 ( .A(n733), .B(n734), .Z(n730) );
  AND U725 ( .A(n61), .B(n729), .Z(n734) );
  XNOR U726 ( .A(n733), .B(n727), .Z(n729) );
  XOR U727 ( .A(n735), .B(n736), .Z(n727) );
  AND U728 ( .A(n76), .B(n737), .Z(n736) );
  XNOR U729 ( .A(n738), .B(n739), .Z(n733) );
  AND U730 ( .A(n68), .B(n740), .Z(n739) );
  XOR U731 ( .A(p_input[59]), .B(n738), .Z(n740) );
  XNOR U732 ( .A(n741), .B(n742), .Z(n738) );
  AND U733 ( .A(n72), .B(n737), .Z(n742) );
  XNOR U734 ( .A(n741), .B(n735), .Z(n737) );
  XOR U735 ( .A(n743), .B(n744), .Z(n735) );
  AND U736 ( .A(n87), .B(n745), .Z(n744) );
  XNOR U737 ( .A(n746), .B(n747), .Z(n741) );
  AND U738 ( .A(n79), .B(n748), .Z(n747) );
  XOR U739 ( .A(p_input[75]), .B(n746), .Z(n748) );
  XNOR U740 ( .A(n749), .B(n750), .Z(n746) );
  AND U741 ( .A(n83), .B(n745), .Z(n750) );
  XNOR U742 ( .A(n749), .B(n743), .Z(n745) );
  XOR U743 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n751), .Z(n743) );
  AND U744 ( .A(n97), .B(n752), .Z(n751) );
  XNOR U745 ( .A(n753), .B(n754), .Z(n749) );
  AND U746 ( .A(n90), .B(n755), .Z(n754) );
  XOR U747 ( .A(p_input[91]), .B(n753), .Z(n755) );
  XNOR U748 ( .A(n756), .B(n757), .Z(n753) );
  AND U749 ( .A(n94), .B(n752), .Z(n757) );
  XOR U750 ( .A(n758), .B(n756), .Z(n752) );
  IV U751 ( .A(\knn_comb_/min_val_out[0][11] ), .Z(n758) );
  IV U752 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n756) );
  XOR U753 ( .A(n27), .B(n759), .Z(o[10]) );
  AND U754 ( .A(n30), .B(n760), .Z(n27) );
  XOR U755 ( .A(n28), .B(n759), .Z(n760) );
  XOR U756 ( .A(n761), .B(n762), .Z(n759) );
  AND U757 ( .A(n42), .B(n763), .Z(n762) );
  XOR U758 ( .A(n764), .B(n765), .Z(n28) );
  AND U759 ( .A(n34), .B(n766), .Z(n765) );
  XOR U760 ( .A(p_input[10]), .B(n764), .Z(n766) );
  XNOR U761 ( .A(n767), .B(n768), .Z(n764) );
  AND U762 ( .A(n38), .B(n763), .Z(n768) );
  XNOR U763 ( .A(n767), .B(n761), .Z(n763) );
  XOR U764 ( .A(n769), .B(n770), .Z(n761) );
  AND U765 ( .A(n54), .B(n771), .Z(n770) );
  XNOR U766 ( .A(n772), .B(n773), .Z(n767) );
  AND U767 ( .A(n46), .B(n774), .Z(n773) );
  XOR U768 ( .A(p_input[26]), .B(n772), .Z(n774) );
  XNOR U769 ( .A(n775), .B(n776), .Z(n772) );
  AND U770 ( .A(n50), .B(n771), .Z(n776) );
  XNOR U771 ( .A(n775), .B(n769), .Z(n771) );
  XOR U772 ( .A(n777), .B(n778), .Z(n769) );
  AND U773 ( .A(n65), .B(n779), .Z(n778) );
  XNOR U774 ( .A(n780), .B(n781), .Z(n775) );
  AND U775 ( .A(n57), .B(n782), .Z(n781) );
  XOR U776 ( .A(p_input[42]), .B(n780), .Z(n782) );
  XNOR U777 ( .A(n783), .B(n784), .Z(n780) );
  AND U778 ( .A(n61), .B(n779), .Z(n784) );
  XNOR U779 ( .A(n783), .B(n777), .Z(n779) );
  XOR U780 ( .A(n785), .B(n786), .Z(n777) );
  AND U781 ( .A(n76), .B(n787), .Z(n786) );
  XNOR U782 ( .A(n788), .B(n789), .Z(n783) );
  AND U783 ( .A(n68), .B(n790), .Z(n789) );
  XOR U784 ( .A(p_input[58]), .B(n788), .Z(n790) );
  XNOR U785 ( .A(n791), .B(n792), .Z(n788) );
  AND U786 ( .A(n72), .B(n787), .Z(n792) );
  XNOR U787 ( .A(n791), .B(n785), .Z(n787) );
  XOR U788 ( .A(n793), .B(n794), .Z(n785) );
  AND U789 ( .A(n87), .B(n795), .Z(n794) );
  XNOR U790 ( .A(n796), .B(n797), .Z(n791) );
  AND U791 ( .A(n79), .B(n798), .Z(n797) );
  XOR U792 ( .A(p_input[74]), .B(n796), .Z(n798) );
  XNOR U793 ( .A(n799), .B(n800), .Z(n796) );
  AND U794 ( .A(n83), .B(n795), .Z(n800) );
  XNOR U795 ( .A(n799), .B(n793), .Z(n795) );
  XOR U796 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n801), .Z(n793) );
  AND U797 ( .A(n97), .B(n802), .Z(n801) );
  XNOR U798 ( .A(n803), .B(n804), .Z(n799) );
  AND U799 ( .A(n90), .B(n805), .Z(n804) );
  XOR U800 ( .A(p_input[90]), .B(n803), .Z(n805) );
  XNOR U801 ( .A(n806), .B(n807), .Z(n803) );
  AND U802 ( .A(n94), .B(n802), .Z(n807) );
  XOR U803 ( .A(\knn_comb_/min_val_out[0][10] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n802) );
  XOR U804 ( .A(n509), .B(n808), .Z(o[0]) );
  AND U805 ( .A(n30), .B(n809), .Z(n509) );
  XOR U806 ( .A(n510), .B(n808), .Z(n809) );
  XOR U807 ( .A(n810), .B(n811), .Z(n808) );
  AND U808 ( .A(n42), .B(n812), .Z(n811) );
  XOR U809 ( .A(n813), .B(n814), .Z(n510) );
  AND U810 ( .A(n34), .B(n815), .Z(n814) );
  XOR U811 ( .A(p_input[0]), .B(n813), .Z(n815) );
  XNOR U812 ( .A(n816), .B(n817), .Z(n813) );
  AND U813 ( .A(n38), .B(n812), .Z(n817) );
  XNOR U814 ( .A(n816), .B(n810), .Z(n812) );
  XOR U815 ( .A(n818), .B(n819), .Z(n810) );
  AND U816 ( .A(n54), .B(n820), .Z(n819) );
  XNOR U817 ( .A(n821), .B(n822), .Z(n816) );
  AND U818 ( .A(n46), .B(n823), .Z(n822) );
  XOR U819 ( .A(p_input[16]), .B(n821), .Z(n823) );
  XNOR U820 ( .A(n824), .B(n825), .Z(n821) );
  AND U821 ( .A(n50), .B(n820), .Z(n825) );
  XNOR U822 ( .A(n824), .B(n818), .Z(n820) );
  XOR U823 ( .A(n826), .B(n827), .Z(n818) );
  AND U824 ( .A(n65), .B(n828), .Z(n827) );
  XNOR U825 ( .A(n829), .B(n830), .Z(n824) );
  AND U826 ( .A(n57), .B(n831), .Z(n830) );
  XOR U827 ( .A(p_input[32]), .B(n829), .Z(n831) );
  XNOR U828 ( .A(n832), .B(n833), .Z(n829) );
  AND U829 ( .A(n61), .B(n828), .Z(n833) );
  XNOR U830 ( .A(n832), .B(n826), .Z(n828) );
  XOR U831 ( .A(n834), .B(n835), .Z(n826) );
  AND U832 ( .A(n76), .B(n836), .Z(n835) );
  XNOR U833 ( .A(n837), .B(n838), .Z(n832) );
  AND U834 ( .A(n68), .B(n839), .Z(n838) );
  XOR U835 ( .A(p_input[48]), .B(n837), .Z(n839) );
  XNOR U836 ( .A(n840), .B(n841), .Z(n837) );
  AND U837 ( .A(n72), .B(n836), .Z(n841) );
  XNOR U838 ( .A(n840), .B(n834), .Z(n836) );
  XOR U839 ( .A(n842), .B(n843), .Z(n834) );
  AND U840 ( .A(n87), .B(n844), .Z(n843) );
  XNOR U841 ( .A(n845), .B(n846), .Z(n840) );
  AND U842 ( .A(n79), .B(n847), .Z(n846) );
  XOR U843 ( .A(p_input[64]), .B(n845), .Z(n847) );
  XNOR U844 ( .A(n848), .B(n849), .Z(n845) );
  AND U845 ( .A(n83), .B(n844), .Z(n849) );
  XNOR U846 ( .A(n848), .B(n842), .Z(n844) );
  XOR U847 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n850), .Z(n842) );
  AND U848 ( .A(n97), .B(n851), .Z(n850) );
  XNOR U849 ( .A(n852), .B(n853), .Z(n848) );
  AND U850 ( .A(n90), .B(n854), .Z(n853) );
  XOR U851 ( .A(p_input[80]), .B(n852), .Z(n854) );
  XNOR U852 ( .A(n855), .B(n856), .Z(n852) );
  AND U853 ( .A(n94), .B(n851), .Z(n856) );
  XOR U854 ( .A(\knn_comb_/min_val_out[0][0] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n851) );
  IV U855 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n855) );
  XNOR U856 ( .A(n857), .B(n858), .Z(n30) );
  AND U857 ( .A(n859), .B(n860), .Z(n858) );
  XNOR U858 ( .A(n857), .B(n861), .Z(n860) );
  XOR U859 ( .A(n862), .B(n863), .Z(n861) );
  AND U860 ( .A(n34), .B(n864), .Z(n863) );
  XNOR U861 ( .A(n862), .B(n865), .Z(n864) );
  XNOR U862 ( .A(n857), .B(n866), .Z(n859) );
  XOR U863 ( .A(n867), .B(n868), .Z(n866) );
  AND U864 ( .A(n42), .B(n869), .Z(n868) );
  XOR U865 ( .A(n870), .B(n871), .Z(n857) );
  AND U866 ( .A(n872), .B(n873), .Z(n871) );
  XOR U867 ( .A(n874), .B(n870), .Z(n873) );
  XOR U868 ( .A(n875), .B(n876), .Z(n874) );
  AND U869 ( .A(n34), .B(n877), .Z(n876) );
  XOR U870 ( .A(n878), .B(n875), .Z(n877) );
  XNOR U871 ( .A(n870), .B(n879), .Z(n872) );
  XOR U872 ( .A(n880), .B(n881), .Z(n879) );
  AND U873 ( .A(n42), .B(n882), .Z(n881) );
  XOR U874 ( .A(n883), .B(n884), .Z(n870) );
  AND U875 ( .A(n885), .B(n886), .Z(n884) );
  XOR U876 ( .A(n887), .B(n883), .Z(n886) );
  XOR U877 ( .A(n888), .B(n889), .Z(n887) );
  AND U878 ( .A(n34), .B(n890), .Z(n889) );
  XNOR U879 ( .A(n891), .B(n888), .Z(n890) );
  XNOR U880 ( .A(n883), .B(n892), .Z(n885) );
  XOR U881 ( .A(n893), .B(n894), .Z(n892) );
  AND U882 ( .A(n42), .B(n895), .Z(n894) );
  XOR U883 ( .A(n896), .B(n897), .Z(n883) );
  AND U884 ( .A(n898), .B(n899), .Z(n897) );
  XOR U885 ( .A(n896), .B(n900), .Z(n899) );
  XOR U886 ( .A(n901), .B(n902), .Z(n900) );
  AND U887 ( .A(n34), .B(n903), .Z(n902) );
  XOR U888 ( .A(n904), .B(n901), .Z(n903) );
  XNOR U889 ( .A(n905), .B(n896), .Z(n898) );
  XNOR U890 ( .A(n906), .B(n907), .Z(n905) );
  AND U891 ( .A(n42), .B(n908), .Z(n907) );
  AND U892 ( .A(n909), .B(n910), .Z(n896) );
  XNOR U893 ( .A(n911), .B(n912), .Z(n910) );
  AND U894 ( .A(n34), .B(n913), .Z(n912) );
  XNOR U895 ( .A(n914), .B(n911), .Z(n913) );
  XNOR U896 ( .A(n915), .B(n916), .Z(n34) );
  AND U897 ( .A(n917), .B(n918), .Z(n916) );
  XOR U898 ( .A(n865), .B(n915), .Z(n918) );
  AND U899 ( .A(n919), .B(n920), .Z(n865) );
  XOR U900 ( .A(n915), .B(n862), .Z(n917) );
  XOR U901 ( .A(n921), .B(n922), .Z(n862) );
  AND U902 ( .A(n38), .B(n869), .Z(n922) );
  XNOR U903 ( .A(n921), .B(n867), .Z(n869) );
  XOR U904 ( .A(n923), .B(n924), .Z(n915) );
  AND U905 ( .A(n925), .B(n926), .Z(n924) );
  XNOR U906 ( .A(n923), .B(n919), .Z(n926) );
  IV U907 ( .A(n878), .Z(n919) );
  XOR U908 ( .A(n927), .B(n928), .Z(n878) );
  XOR U909 ( .A(n929), .B(n920), .Z(n928) );
  AND U910 ( .A(n891), .B(n930), .Z(n920) );
  AND U911 ( .A(n931), .B(n932), .Z(n929) );
  XOR U912 ( .A(n933), .B(n927), .Z(n931) );
  XNOR U913 ( .A(n875), .B(n923), .Z(n925) );
  XNOR U914 ( .A(n934), .B(n935), .Z(n875) );
  AND U915 ( .A(n38), .B(n882), .Z(n935) );
  XOR U916 ( .A(n934), .B(n936), .Z(n882) );
  XOR U917 ( .A(n937), .B(n938), .Z(n923) );
  AND U918 ( .A(n939), .B(n940), .Z(n938) );
  XNOR U919 ( .A(n937), .B(n891), .Z(n940) );
  XOR U920 ( .A(n941), .B(n932), .Z(n891) );
  XNOR U921 ( .A(n942), .B(n927), .Z(n932) );
  XOR U922 ( .A(n943), .B(n944), .Z(n927) );
  AND U923 ( .A(n945), .B(n946), .Z(n944) );
  XOR U924 ( .A(n947), .B(n943), .Z(n945) );
  XNOR U925 ( .A(n948), .B(n949), .Z(n942) );
  AND U926 ( .A(n950), .B(n951), .Z(n949) );
  XOR U927 ( .A(n948), .B(n952), .Z(n950) );
  XNOR U928 ( .A(n933), .B(n930), .Z(n941) );
  AND U929 ( .A(n953), .B(n954), .Z(n930) );
  XOR U930 ( .A(n955), .B(n956), .Z(n933) );
  AND U931 ( .A(n957), .B(n958), .Z(n956) );
  XOR U932 ( .A(n955), .B(n959), .Z(n957) );
  XNOR U933 ( .A(n888), .B(n937), .Z(n939) );
  XNOR U934 ( .A(n960), .B(n961), .Z(n888) );
  AND U935 ( .A(n38), .B(n895), .Z(n961) );
  XOR U936 ( .A(n960), .B(n962), .Z(n895) );
  XOR U937 ( .A(n963), .B(n964), .Z(n937) );
  AND U938 ( .A(n965), .B(n966), .Z(n964) );
  XNOR U939 ( .A(n963), .B(n953), .Z(n966) );
  IV U940 ( .A(n904), .Z(n953) );
  XNOR U941 ( .A(n967), .B(n946), .Z(n904) );
  XNOR U942 ( .A(n968), .B(n952), .Z(n946) );
  XNOR U943 ( .A(n969), .B(n970), .Z(n952) );
  NOR U944 ( .A(n971), .B(n972), .Z(n970) );
  XOR U945 ( .A(n969), .B(n973), .Z(n971) );
  XNOR U946 ( .A(n951), .B(n943), .Z(n968) );
  XOR U947 ( .A(n974), .B(n975), .Z(n943) );
  AND U948 ( .A(n976), .B(n977), .Z(n975) );
  XNOR U949 ( .A(n974), .B(n978), .Z(n976) );
  XNOR U950 ( .A(n979), .B(n948), .Z(n951) );
  XOR U951 ( .A(n980), .B(n981), .Z(n948) );
  AND U952 ( .A(n982), .B(n983), .Z(n981) );
  XOR U953 ( .A(n980), .B(n984), .Z(n982) );
  XNOR U954 ( .A(n985), .B(n986), .Z(n979) );
  NOR U955 ( .A(n987), .B(n988), .Z(n986) );
  XOR U956 ( .A(n985), .B(n989), .Z(n987) );
  XNOR U957 ( .A(n947), .B(n954), .Z(n967) );
  NOR U958 ( .A(n914), .B(n990), .Z(n954) );
  XOR U959 ( .A(n959), .B(n958), .Z(n947) );
  XNOR U960 ( .A(n991), .B(n955), .Z(n958) );
  XOR U961 ( .A(n992), .B(n993), .Z(n955) );
  AND U962 ( .A(n994), .B(n995), .Z(n993) );
  XOR U963 ( .A(n992), .B(n996), .Z(n994) );
  XNOR U964 ( .A(n997), .B(n998), .Z(n991) );
  NOR U965 ( .A(n999), .B(n1000), .Z(n998) );
  XNOR U966 ( .A(n997), .B(n1001), .Z(n999) );
  XOR U967 ( .A(n1002), .B(n1003), .Z(n959) );
  NOR U968 ( .A(n1004), .B(n1005), .Z(n1003) );
  XNOR U969 ( .A(n1002), .B(n1006), .Z(n1004) );
  XNOR U970 ( .A(n901), .B(n963), .Z(n965) );
  XNOR U971 ( .A(n1007), .B(n1008), .Z(n901) );
  AND U972 ( .A(n38), .B(n908), .Z(n1008) );
  XOR U973 ( .A(n1007), .B(n906), .Z(n908) );
  AND U974 ( .A(n911), .B(n914), .Z(n963) );
  XOR U975 ( .A(n1009), .B(n990), .Z(n914) );
  XNOR U976 ( .A(p_input[0]), .B(p_input[128]), .Z(n990) );
  XOR U977 ( .A(n978), .B(n977), .Z(n1009) );
  XNOR U978 ( .A(n1010), .B(n984), .Z(n977) );
  XNOR U979 ( .A(n973), .B(n972), .Z(n984) );
  XOR U980 ( .A(n1011), .B(n1012), .Z(n972) );
  IV U981 ( .A(n969), .Z(n1012) );
  XNOR U982 ( .A(p_input[10]), .B(p_input[138]), .Z(n969) );
  XOR U983 ( .A(p_input[11]), .B(n1013), .Z(n1011) );
  XOR U984 ( .A(p_input[12]), .B(p_input[140]), .Z(n973) );
  XNOR U985 ( .A(n983), .B(n974), .Z(n1010) );
  XOR U986 ( .A(p_input[129]), .B(p_input[1]), .Z(n974) );
  XOR U987 ( .A(n1014), .B(n989), .Z(n983) );
  XNOR U988 ( .A(p_input[143]), .B(p_input[15]), .Z(n989) );
  XOR U989 ( .A(n980), .B(n988), .Z(n1014) );
  XOR U990 ( .A(n1015), .B(n985), .Z(n988) );
  XOR U991 ( .A(p_input[13]), .B(p_input[141]), .Z(n985) );
  XNOR U992 ( .A(p_input[142]), .B(p_input[14]), .Z(n1015) );
  XOR U993 ( .A(p_input[137]), .B(p_input[9]), .Z(n980) );
  XNOR U994 ( .A(n996), .B(n995), .Z(n978) );
  XNOR U995 ( .A(n1016), .B(n1001), .Z(n995) );
  XOR U996 ( .A(p_input[136]), .B(p_input[8]), .Z(n1001) );
  XOR U997 ( .A(n992), .B(n1000), .Z(n1016) );
  XOR U998 ( .A(n1017), .B(n997), .Z(n1000) );
  XOR U999 ( .A(p_input[134]), .B(p_input[6]), .Z(n997) );
  XNOR U1000 ( .A(p_input[135]), .B(p_input[7]), .Z(n1017) );
  XOR U1001 ( .A(p_input[130]), .B(p_input[2]), .Z(n992) );
  XNOR U1002 ( .A(n1006), .B(n1005), .Z(n996) );
  XOR U1003 ( .A(n1018), .B(n1002), .Z(n1005) );
  XOR U1004 ( .A(p_input[131]), .B(p_input[3]), .Z(n1002) );
  XNOR U1005 ( .A(p_input[132]), .B(p_input[4]), .Z(n1018) );
  XOR U1006 ( .A(p_input[133]), .B(p_input[5]), .Z(n1006) );
  XNOR U1007 ( .A(n1019), .B(n1020), .Z(n911) );
  AND U1008 ( .A(n38), .B(n1021), .Z(n1020) );
  XNOR U1009 ( .A(n1022), .B(n1023), .Z(n38) );
  AND U1010 ( .A(n1024), .B(n1025), .Z(n1023) );
  XNOR U1011 ( .A(n1022), .B(n921), .Z(n1025) );
  XNOR U1012 ( .A(n1022), .B(n867), .Z(n1024) );
  XOR U1013 ( .A(n1026), .B(n1027), .Z(n1022) );
  AND U1014 ( .A(n1028), .B(n1029), .Z(n1027) );
  XNOR U1015 ( .A(n934), .B(n1026), .Z(n1029) );
  XOR U1016 ( .A(n1026), .B(n936), .Z(n1028) );
  XOR U1017 ( .A(n1030), .B(n1031), .Z(n1026) );
  AND U1018 ( .A(n1032), .B(n1033), .Z(n1031) );
  XOR U1019 ( .A(n1030), .B(n962), .Z(n1032) );
  IV U1020 ( .A(n893), .Z(n962) );
  XOR U1021 ( .A(n1034), .B(n1035), .Z(n909) );
  AND U1022 ( .A(n42), .B(n1021), .Z(n1035) );
  XNOR U1023 ( .A(n1019), .B(n1034), .Z(n1021) );
  XNOR U1024 ( .A(n1036), .B(n1037), .Z(n42) );
  AND U1025 ( .A(n1038), .B(n1039), .Z(n1037) );
  XNOR U1026 ( .A(n921), .B(n1036), .Z(n1039) );
  XOR U1027 ( .A(n1040), .B(n1041), .Z(n921) );
  AND U1028 ( .A(n1042), .B(n46), .Z(n1041) );
  NOR U1029 ( .A(n1043), .B(n1040), .Z(n1042) );
  XNOR U1030 ( .A(n1036), .B(n867), .Z(n1038) );
  AND U1031 ( .A(n1044), .B(n1045), .Z(n867) );
  XOR U1032 ( .A(n1046), .B(n1047), .Z(n1036) );
  AND U1033 ( .A(n1048), .B(n1049), .Z(n1047) );
  XNOR U1034 ( .A(n1046), .B(n934), .Z(n1049) );
  XNOR U1035 ( .A(n1050), .B(n1051), .Z(n934) );
  AND U1036 ( .A(n46), .B(n1052), .Z(n1051) );
  XOR U1037 ( .A(n1053), .B(n1050), .Z(n1052) );
  XNOR U1038 ( .A(n880), .B(n1046), .Z(n1048) );
  IV U1039 ( .A(n936), .Z(n880) );
  XOR U1040 ( .A(n1054), .B(n1055), .Z(n936) );
  AND U1041 ( .A(n54), .B(n1056), .Z(n1055) );
  XOR U1042 ( .A(n1030), .B(n1057), .Z(n1046) );
  AND U1043 ( .A(n1058), .B(n1033), .Z(n1057) );
  XNOR U1044 ( .A(n960), .B(n1030), .Z(n1033) );
  XNOR U1045 ( .A(n1059), .B(n1060), .Z(n960) );
  AND U1046 ( .A(n46), .B(n1061), .Z(n1060) );
  XNOR U1047 ( .A(n1062), .B(n1059), .Z(n1061) );
  XNOR U1048 ( .A(n893), .B(n1030), .Z(n1058) );
  XNOR U1049 ( .A(n1063), .B(n1064), .Z(n893) );
  AND U1050 ( .A(n54), .B(n1065), .Z(n1064) );
  XOR U1051 ( .A(n1066), .B(n1067), .Z(n1030) );
  AND U1052 ( .A(n1068), .B(n1069), .Z(n1067) );
  XNOR U1053 ( .A(n1066), .B(n1007), .Z(n1069) );
  XNOR U1054 ( .A(n1070), .B(n1071), .Z(n1007) );
  AND U1055 ( .A(n46), .B(n1072), .Z(n1071) );
  XOR U1056 ( .A(n1073), .B(n1070), .Z(n1072) );
  XNOR U1057 ( .A(n1074), .B(n1066), .Z(n1068) );
  IV U1058 ( .A(n906), .Z(n1074) );
  XOR U1059 ( .A(n1075), .B(n1076), .Z(n906) );
  AND U1060 ( .A(n54), .B(n1077), .Z(n1076) );
  AND U1061 ( .A(n1034), .B(n1019), .Z(n1066) );
  XNOR U1062 ( .A(n1078), .B(n1079), .Z(n1019) );
  AND U1063 ( .A(n46), .B(n1080), .Z(n1079) );
  XNOR U1064 ( .A(n1081), .B(n1078), .Z(n1080) );
  XNOR U1065 ( .A(n1082), .B(n1083), .Z(n46) );
  AND U1066 ( .A(n1084), .B(n1085), .Z(n1083) );
  XOR U1067 ( .A(n1043), .B(n1082), .Z(n1085) );
  AND U1068 ( .A(n1086), .B(n1087), .Z(n1043) );
  XOR U1069 ( .A(n1040), .B(n1082), .Z(n1084) );
  NOR U1070 ( .A(n1044), .B(n1045), .Z(n1040) );
  XOR U1071 ( .A(n1088), .B(n1089), .Z(n1082) );
  AND U1072 ( .A(n1090), .B(n1091), .Z(n1089) );
  XNOR U1073 ( .A(n1088), .B(n1086), .Z(n1091) );
  IV U1074 ( .A(n1053), .Z(n1086) );
  XOR U1075 ( .A(n1092), .B(n1093), .Z(n1053) );
  XOR U1076 ( .A(n1094), .B(n1087), .Z(n1093) );
  AND U1077 ( .A(n1062), .B(n1095), .Z(n1087) );
  AND U1078 ( .A(n1096), .B(n1097), .Z(n1094) );
  XOR U1079 ( .A(n1098), .B(n1092), .Z(n1096) );
  XNOR U1080 ( .A(n1050), .B(n1088), .Z(n1090) );
  XNOR U1081 ( .A(n1099), .B(n1100), .Z(n1050) );
  AND U1082 ( .A(n50), .B(n1056), .Z(n1100) );
  XOR U1083 ( .A(n1099), .B(n1054), .Z(n1056) );
  XOR U1084 ( .A(n1101), .B(n1102), .Z(n1088) );
  AND U1085 ( .A(n1103), .B(n1104), .Z(n1102) );
  XNOR U1086 ( .A(n1101), .B(n1062), .Z(n1104) );
  XOR U1087 ( .A(n1105), .B(n1097), .Z(n1062) );
  XNOR U1088 ( .A(n1106), .B(n1092), .Z(n1097) );
  XOR U1089 ( .A(n1107), .B(n1108), .Z(n1092) );
  AND U1090 ( .A(n1109), .B(n1110), .Z(n1108) );
  XOR U1091 ( .A(n1111), .B(n1107), .Z(n1109) );
  XNOR U1092 ( .A(n1112), .B(n1113), .Z(n1106) );
  AND U1093 ( .A(n1114), .B(n1115), .Z(n1113) );
  XOR U1094 ( .A(n1112), .B(n1116), .Z(n1114) );
  XNOR U1095 ( .A(n1098), .B(n1095), .Z(n1105) );
  AND U1096 ( .A(n1117), .B(n1118), .Z(n1095) );
  XOR U1097 ( .A(n1119), .B(n1120), .Z(n1098) );
  AND U1098 ( .A(n1121), .B(n1122), .Z(n1120) );
  XOR U1099 ( .A(n1119), .B(n1123), .Z(n1121) );
  XNOR U1100 ( .A(n1059), .B(n1101), .Z(n1103) );
  XNOR U1101 ( .A(n1124), .B(n1125), .Z(n1059) );
  AND U1102 ( .A(n50), .B(n1065), .Z(n1125) );
  XOR U1103 ( .A(n1124), .B(n1063), .Z(n1065) );
  XOR U1104 ( .A(n1126), .B(n1127), .Z(n1101) );
  AND U1105 ( .A(n1128), .B(n1129), .Z(n1127) );
  XNOR U1106 ( .A(n1126), .B(n1117), .Z(n1129) );
  IV U1107 ( .A(n1073), .Z(n1117) );
  XNOR U1108 ( .A(n1130), .B(n1110), .Z(n1073) );
  XNOR U1109 ( .A(n1131), .B(n1116), .Z(n1110) );
  XOR U1110 ( .A(n1132), .B(n1133), .Z(n1116) );
  NOR U1111 ( .A(n1134), .B(n1135), .Z(n1133) );
  XNOR U1112 ( .A(n1132), .B(n1136), .Z(n1134) );
  XNOR U1113 ( .A(n1115), .B(n1107), .Z(n1131) );
  XOR U1114 ( .A(n1137), .B(n1138), .Z(n1107) );
  AND U1115 ( .A(n1139), .B(n1140), .Z(n1138) );
  XNOR U1116 ( .A(n1137), .B(n1141), .Z(n1139) );
  XNOR U1117 ( .A(n1142), .B(n1112), .Z(n1115) );
  XOR U1118 ( .A(n1143), .B(n1144), .Z(n1112) );
  AND U1119 ( .A(n1145), .B(n1146), .Z(n1144) );
  XOR U1120 ( .A(n1143), .B(n1147), .Z(n1145) );
  XNOR U1121 ( .A(n1148), .B(n1149), .Z(n1142) );
  NOR U1122 ( .A(n1150), .B(n1151), .Z(n1149) );
  XOR U1123 ( .A(n1148), .B(n1152), .Z(n1150) );
  XNOR U1124 ( .A(n1111), .B(n1118), .Z(n1130) );
  NOR U1125 ( .A(n1081), .B(n1153), .Z(n1118) );
  XOR U1126 ( .A(n1123), .B(n1122), .Z(n1111) );
  XNOR U1127 ( .A(n1154), .B(n1119), .Z(n1122) );
  XOR U1128 ( .A(n1155), .B(n1156), .Z(n1119) );
  AND U1129 ( .A(n1157), .B(n1158), .Z(n1156) );
  XOR U1130 ( .A(n1155), .B(n1159), .Z(n1157) );
  XNOR U1131 ( .A(n1160), .B(n1161), .Z(n1154) );
  NOR U1132 ( .A(n1162), .B(n1163), .Z(n1161) );
  XNOR U1133 ( .A(n1160), .B(n1164), .Z(n1162) );
  XOR U1134 ( .A(n1165), .B(n1166), .Z(n1123) );
  NOR U1135 ( .A(n1167), .B(n1168), .Z(n1166) );
  XNOR U1136 ( .A(n1165), .B(n1169), .Z(n1167) );
  XNOR U1137 ( .A(n1070), .B(n1126), .Z(n1128) );
  XNOR U1138 ( .A(n1170), .B(n1171), .Z(n1070) );
  AND U1139 ( .A(n50), .B(n1077), .Z(n1171) );
  XOR U1140 ( .A(n1170), .B(n1075), .Z(n1077) );
  AND U1141 ( .A(n1078), .B(n1081), .Z(n1126) );
  XOR U1142 ( .A(n1172), .B(n1153), .Z(n1081) );
  XNOR U1143 ( .A(p_input[128]), .B(p_input[16]), .Z(n1153) );
  XOR U1144 ( .A(n1141), .B(n1140), .Z(n1172) );
  XNOR U1145 ( .A(n1173), .B(n1147), .Z(n1140) );
  XNOR U1146 ( .A(n1136), .B(n1135), .Z(n1147) );
  XOR U1147 ( .A(n1174), .B(n1132), .Z(n1135) );
  XOR U1148 ( .A(p_input[138]), .B(p_input[26]), .Z(n1132) );
  XNOR U1149 ( .A(p_input[139]), .B(p_input[27]), .Z(n1174) );
  XOR U1150 ( .A(p_input[140]), .B(p_input[28]), .Z(n1136) );
  XNOR U1151 ( .A(n1146), .B(n1137), .Z(n1173) );
  XOR U1152 ( .A(p_input[129]), .B(p_input[17]), .Z(n1137) );
  XOR U1153 ( .A(n1175), .B(n1152), .Z(n1146) );
  XNOR U1154 ( .A(p_input[143]), .B(p_input[31]), .Z(n1152) );
  XOR U1155 ( .A(n1143), .B(n1151), .Z(n1175) );
  XOR U1156 ( .A(n1176), .B(n1148), .Z(n1151) );
  XOR U1157 ( .A(p_input[141]), .B(p_input[29]), .Z(n1148) );
  XNOR U1158 ( .A(p_input[142]), .B(p_input[30]), .Z(n1176) );
  XOR U1159 ( .A(p_input[137]), .B(p_input[25]), .Z(n1143) );
  XNOR U1160 ( .A(n1159), .B(n1158), .Z(n1141) );
  XNOR U1161 ( .A(n1177), .B(n1164), .Z(n1158) );
  XOR U1162 ( .A(p_input[136]), .B(p_input[24]), .Z(n1164) );
  XOR U1163 ( .A(n1155), .B(n1163), .Z(n1177) );
  XOR U1164 ( .A(n1178), .B(n1160), .Z(n1163) );
  XOR U1165 ( .A(p_input[134]), .B(p_input[22]), .Z(n1160) );
  XNOR U1166 ( .A(p_input[135]), .B(p_input[23]), .Z(n1178) );
  XOR U1167 ( .A(p_input[130]), .B(p_input[18]), .Z(n1155) );
  XNOR U1168 ( .A(n1169), .B(n1168), .Z(n1159) );
  XOR U1169 ( .A(n1179), .B(n1165), .Z(n1168) );
  XOR U1170 ( .A(p_input[131]), .B(p_input[19]), .Z(n1165) );
  XNOR U1171 ( .A(p_input[132]), .B(p_input[20]), .Z(n1179) );
  XOR U1172 ( .A(p_input[133]), .B(p_input[21]), .Z(n1169) );
  XNOR U1173 ( .A(n1180), .B(n1181), .Z(n1078) );
  AND U1174 ( .A(n50), .B(n1182), .Z(n1181) );
  XNOR U1175 ( .A(n1183), .B(n1184), .Z(n50) );
  NOR U1176 ( .A(n1185), .B(n1186), .Z(n1184) );
  XOR U1177 ( .A(n1045), .B(n1183), .Z(n1186) );
  NOR U1178 ( .A(n1183), .B(n1044), .Z(n1185) );
  XOR U1179 ( .A(n1187), .B(n1188), .Z(n1183) );
  AND U1180 ( .A(n1189), .B(n1190), .Z(n1188) );
  XOR U1181 ( .A(n1187), .B(n1054), .Z(n1189) );
  XOR U1182 ( .A(n1191), .B(n1192), .Z(n1034) );
  AND U1183 ( .A(n54), .B(n1182), .Z(n1192) );
  XNOR U1184 ( .A(n1180), .B(n1191), .Z(n1182) );
  XNOR U1185 ( .A(n1193), .B(n1194), .Z(n54) );
  NOR U1186 ( .A(n1195), .B(n1196), .Z(n1194) );
  XNOR U1187 ( .A(n1045), .B(n1197), .Z(n1196) );
  IV U1188 ( .A(n1193), .Z(n1197) );
  AND U1189 ( .A(n1198), .B(n1199), .Z(n1045) );
  NOR U1190 ( .A(n1193), .B(n1044), .Z(n1195) );
  AND U1191 ( .A(n1200), .B(n1201), .Z(n1044) );
  IV U1192 ( .A(n1202), .Z(n1200) );
  XOR U1193 ( .A(n1187), .B(n1203), .Z(n1193) );
  AND U1194 ( .A(n1204), .B(n1190), .Z(n1203) );
  XNOR U1195 ( .A(n1099), .B(n1187), .Z(n1190) );
  XNOR U1196 ( .A(n1205), .B(n1206), .Z(n1099) );
  AND U1197 ( .A(n57), .B(n1207), .Z(n1206) );
  XOR U1198 ( .A(n1208), .B(n1205), .Z(n1207) );
  XNOR U1199 ( .A(n1209), .B(n1187), .Z(n1204) );
  IV U1200 ( .A(n1054), .Z(n1209) );
  XOR U1201 ( .A(n1210), .B(n1211), .Z(n1054) );
  AND U1202 ( .A(n65), .B(n1212), .Z(n1211) );
  XOR U1203 ( .A(n1213), .B(n1214), .Z(n1187) );
  AND U1204 ( .A(n1215), .B(n1216), .Z(n1214) );
  XNOR U1205 ( .A(n1124), .B(n1213), .Z(n1216) );
  XNOR U1206 ( .A(n1217), .B(n1218), .Z(n1124) );
  AND U1207 ( .A(n57), .B(n1219), .Z(n1218) );
  XNOR U1208 ( .A(n1220), .B(n1217), .Z(n1219) );
  XOR U1209 ( .A(n1213), .B(n1063), .Z(n1215) );
  XOR U1210 ( .A(n1221), .B(n1222), .Z(n1063) );
  AND U1211 ( .A(n65), .B(n1223), .Z(n1222) );
  XOR U1212 ( .A(n1224), .B(n1225), .Z(n1213) );
  AND U1213 ( .A(n1226), .B(n1227), .Z(n1225) );
  XNOR U1214 ( .A(n1224), .B(n1170), .Z(n1227) );
  XNOR U1215 ( .A(n1228), .B(n1229), .Z(n1170) );
  AND U1216 ( .A(n57), .B(n1230), .Z(n1229) );
  XOR U1217 ( .A(n1231), .B(n1228), .Z(n1230) );
  XNOR U1218 ( .A(n1232), .B(n1224), .Z(n1226) );
  IV U1219 ( .A(n1075), .Z(n1232) );
  XOR U1220 ( .A(n1233), .B(n1234), .Z(n1075) );
  AND U1221 ( .A(n65), .B(n1235), .Z(n1234) );
  AND U1222 ( .A(n1191), .B(n1180), .Z(n1224) );
  XNOR U1223 ( .A(n1236), .B(n1237), .Z(n1180) );
  AND U1224 ( .A(n57), .B(n1238), .Z(n1237) );
  XNOR U1225 ( .A(n1239), .B(n1236), .Z(n1238) );
  XNOR U1226 ( .A(n1240), .B(n1241), .Z(n57) );
  NOR U1227 ( .A(n1242), .B(n1243), .Z(n1241) );
  XNOR U1228 ( .A(n1240), .B(n1202), .Z(n1243) );
  NOR U1229 ( .A(n1198), .B(n1199), .Z(n1202) );
  NOR U1230 ( .A(n1240), .B(n1201), .Z(n1242) );
  AND U1231 ( .A(n1244), .B(n1245), .Z(n1201) );
  XOR U1232 ( .A(n1246), .B(n1247), .Z(n1240) );
  AND U1233 ( .A(n1248), .B(n1249), .Z(n1247) );
  XNOR U1234 ( .A(n1246), .B(n1244), .Z(n1249) );
  IV U1235 ( .A(n1208), .Z(n1244) );
  XOR U1236 ( .A(n1250), .B(n1251), .Z(n1208) );
  XOR U1237 ( .A(n1252), .B(n1245), .Z(n1251) );
  AND U1238 ( .A(n1220), .B(n1253), .Z(n1245) );
  AND U1239 ( .A(n1254), .B(n1255), .Z(n1252) );
  XOR U1240 ( .A(n1256), .B(n1250), .Z(n1254) );
  XNOR U1241 ( .A(n1205), .B(n1246), .Z(n1248) );
  XNOR U1242 ( .A(n1257), .B(n1258), .Z(n1205) );
  AND U1243 ( .A(n61), .B(n1212), .Z(n1258) );
  XOR U1244 ( .A(n1257), .B(n1210), .Z(n1212) );
  XOR U1245 ( .A(n1259), .B(n1260), .Z(n1246) );
  AND U1246 ( .A(n1261), .B(n1262), .Z(n1260) );
  XNOR U1247 ( .A(n1259), .B(n1220), .Z(n1262) );
  XOR U1248 ( .A(n1263), .B(n1255), .Z(n1220) );
  XNOR U1249 ( .A(n1264), .B(n1250), .Z(n1255) );
  XOR U1250 ( .A(n1265), .B(n1266), .Z(n1250) );
  AND U1251 ( .A(n1267), .B(n1268), .Z(n1266) );
  XOR U1252 ( .A(n1269), .B(n1265), .Z(n1267) );
  XNOR U1253 ( .A(n1270), .B(n1271), .Z(n1264) );
  AND U1254 ( .A(n1272), .B(n1273), .Z(n1271) );
  XOR U1255 ( .A(n1270), .B(n1274), .Z(n1272) );
  XNOR U1256 ( .A(n1256), .B(n1253), .Z(n1263) );
  AND U1257 ( .A(n1275), .B(n1276), .Z(n1253) );
  XOR U1258 ( .A(n1277), .B(n1278), .Z(n1256) );
  AND U1259 ( .A(n1279), .B(n1280), .Z(n1278) );
  XOR U1260 ( .A(n1277), .B(n1281), .Z(n1279) );
  XNOR U1261 ( .A(n1217), .B(n1259), .Z(n1261) );
  XNOR U1262 ( .A(n1282), .B(n1283), .Z(n1217) );
  AND U1263 ( .A(n61), .B(n1223), .Z(n1283) );
  XOR U1264 ( .A(n1282), .B(n1221), .Z(n1223) );
  XOR U1265 ( .A(n1284), .B(n1285), .Z(n1259) );
  AND U1266 ( .A(n1286), .B(n1287), .Z(n1285) );
  XNOR U1267 ( .A(n1284), .B(n1275), .Z(n1287) );
  IV U1268 ( .A(n1231), .Z(n1275) );
  XNOR U1269 ( .A(n1288), .B(n1268), .Z(n1231) );
  XNOR U1270 ( .A(n1289), .B(n1274), .Z(n1268) );
  XOR U1271 ( .A(n1290), .B(n1291), .Z(n1274) );
  NOR U1272 ( .A(n1292), .B(n1293), .Z(n1291) );
  XNOR U1273 ( .A(n1290), .B(n1294), .Z(n1292) );
  XNOR U1274 ( .A(n1273), .B(n1265), .Z(n1289) );
  XOR U1275 ( .A(n1295), .B(n1296), .Z(n1265) );
  AND U1276 ( .A(n1297), .B(n1298), .Z(n1296) );
  XNOR U1277 ( .A(n1295), .B(n1299), .Z(n1297) );
  XNOR U1278 ( .A(n1300), .B(n1270), .Z(n1273) );
  XOR U1279 ( .A(n1301), .B(n1302), .Z(n1270) );
  AND U1280 ( .A(n1303), .B(n1304), .Z(n1302) );
  XOR U1281 ( .A(n1301), .B(n1305), .Z(n1303) );
  XNOR U1282 ( .A(n1306), .B(n1307), .Z(n1300) );
  NOR U1283 ( .A(n1308), .B(n1309), .Z(n1307) );
  XOR U1284 ( .A(n1306), .B(n1310), .Z(n1308) );
  XNOR U1285 ( .A(n1269), .B(n1276), .Z(n1288) );
  NOR U1286 ( .A(n1239), .B(n1311), .Z(n1276) );
  XOR U1287 ( .A(n1281), .B(n1280), .Z(n1269) );
  XNOR U1288 ( .A(n1312), .B(n1277), .Z(n1280) );
  XOR U1289 ( .A(n1313), .B(n1314), .Z(n1277) );
  AND U1290 ( .A(n1315), .B(n1316), .Z(n1314) );
  XOR U1291 ( .A(n1313), .B(n1317), .Z(n1315) );
  XNOR U1292 ( .A(n1318), .B(n1319), .Z(n1312) );
  NOR U1293 ( .A(n1320), .B(n1321), .Z(n1319) );
  XNOR U1294 ( .A(n1318), .B(n1322), .Z(n1320) );
  XOR U1295 ( .A(n1323), .B(n1324), .Z(n1281) );
  NOR U1296 ( .A(n1325), .B(n1326), .Z(n1324) );
  XNOR U1297 ( .A(n1323), .B(n1327), .Z(n1325) );
  XNOR U1298 ( .A(n1228), .B(n1284), .Z(n1286) );
  XNOR U1299 ( .A(n1328), .B(n1329), .Z(n1228) );
  AND U1300 ( .A(n61), .B(n1235), .Z(n1329) );
  XOR U1301 ( .A(n1328), .B(n1233), .Z(n1235) );
  AND U1302 ( .A(n1236), .B(n1239), .Z(n1284) );
  XOR U1303 ( .A(n1330), .B(n1311), .Z(n1239) );
  XNOR U1304 ( .A(p_input[128]), .B(p_input[32]), .Z(n1311) );
  XOR U1305 ( .A(n1299), .B(n1298), .Z(n1330) );
  XNOR U1306 ( .A(n1331), .B(n1305), .Z(n1298) );
  XNOR U1307 ( .A(n1294), .B(n1293), .Z(n1305) );
  XOR U1308 ( .A(n1332), .B(n1290), .Z(n1293) );
  XOR U1309 ( .A(p_input[138]), .B(p_input[42]), .Z(n1290) );
  XNOR U1310 ( .A(p_input[139]), .B(p_input[43]), .Z(n1332) );
  XOR U1311 ( .A(p_input[140]), .B(p_input[44]), .Z(n1294) );
  XNOR U1312 ( .A(n1304), .B(n1295), .Z(n1331) );
  XOR U1313 ( .A(p_input[129]), .B(p_input[33]), .Z(n1295) );
  XOR U1314 ( .A(n1333), .B(n1310), .Z(n1304) );
  XNOR U1315 ( .A(p_input[143]), .B(p_input[47]), .Z(n1310) );
  XOR U1316 ( .A(n1301), .B(n1309), .Z(n1333) );
  XOR U1317 ( .A(n1334), .B(n1306), .Z(n1309) );
  XOR U1318 ( .A(p_input[141]), .B(p_input[45]), .Z(n1306) );
  XNOR U1319 ( .A(p_input[142]), .B(p_input[46]), .Z(n1334) );
  XOR U1320 ( .A(p_input[137]), .B(p_input[41]), .Z(n1301) );
  XNOR U1321 ( .A(n1317), .B(n1316), .Z(n1299) );
  XNOR U1322 ( .A(n1335), .B(n1322), .Z(n1316) );
  XOR U1323 ( .A(p_input[136]), .B(p_input[40]), .Z(n1322) );
  XOR U1324 ( .A(n1313), .B(n1321), .Z(n1335) );
  XOR U1325 ( .A(n1336), .B(n1318), .Z(n1321) );
  XOR U1326 ( .A(p_input[134]), .B(p_input[38]), .Z(n1318) );
  XNOR U1327 ( .A(p_input[135]), .B(p_input[39]), .Z(n1336) );
  XOR U1328 ( .A(p_input[130]), .B(p_input[34]), .Z(n1313) );
  XNOR U1329 ( .A(n1327), .B(n1326), .Z(n1317) );
  XOR U1330 ( .A(n1337), .B(n1323), .Z(n1326) );
  XOR U1331 ( .A(p_input[131]), .B(p_input[35]), .Z(n1323) );
  XNOR U1332 ( .A(p_input[132]), .B(p_input[36]), .Z(n1337) );
  XOR U1333 ( .A(p_input[133]), .B(p_input[37]), .Z(n1327) );
  XNOR U1334 ( .A(n1338), .B(n1339), .Z(n1236) );
  AND U1335 ( .A(n61), .B(n1340), .Z(n1339) );
  XNOR U1336 ( .A(n1341), .B(n1342), .Z(n61) );
  NOR U1337 ( .A(n1343), .B(n1344), .Z(n1342) );
  XOR U1338 ( .A(n1199), .B(n1341), .Z(n1344) );
  NOR U1339 ( .A(n1341), .B(n1198), .Z(n1343) );
  XOR U1340 ( .A(n1345), .B(n1346), .Z(n1341) );
  AND U1341 ( .A(n1347), .B(n1348), .Z(n1346) );
  XOR U1342 ( .A(n1345), .B(n1210), .Z(n1347) );
  XOR U1343 ( .A(n1349), .B(n1350), .Z(n1191) );
  AND U1344 ( .A(n65), .B(n1340), .Z(n1350) );
  XNOR U1345 ( .A(n1338), .B(n1349), .Z(n1340) );
  XNOR U1346 ( .A(n1351), .B(n1352), .Z(n65) );
  NOR U1347 ( .A(n1353), .B(n1354), .Z(n1352) );
  XNOR U1348 ( .A(n1199), .B(n1355), .Z(n1354) );
  IV U1349 ( .A(n1351), .Z(n1355) );
  AND U1350 ( .A(n1356), .B(n1357), .Z(n1199) );
  NOR U1351 ( .A(n1351), .B(n1198), .Z(n1353) );
  AND U1352 ( .A(n1358), .B(n1359), .Z(n1198) );
  IV U1353 ( .A(n1360), .Z(n1358) );
  XOR U1354 ( .A(n1345), .B(n1361), .Z(n1351) );
  AND U1355 ( .A(n1362), .B(n1348), .Z(n1361) );
  XNOR U1356 ( .A(n1257), .B(n1345), .Z(n1348) );
  XNOR U1357 ( .A(n1363), .B(n1364), .Z(n1257) );
  AND U1358 ( .A(n68), .B(n1365), .Z(n1364) );
  XOR U1359 ( .A(n1366), .B(n1363), .Z(n1365) );
  XNOR U1360 ( .A(n1367), .B(n1345), .Z(n1362) );
  IV U1361 ( .A(n1210), .Z(n1367) );
  XOR U1362 ( .A(n1368), .B(n1369), .Z(n1210) );
  AND U1363 ( .A(n76), .B(n1370), .Z(n1369) );
  XOR U1364 ( .A(n1371), .B(n1372), .Z(n1345) );
  AND U1365 ( .A(n1373), .B(n1374), .Z(n1372) );
  XNOR U1366 ( .A(n1282), .B(n1371), .Z(n1374) );
  XNOR U1367 ( .A(n1375), .B(n1376), .Z(n1282) );
  AND U1368 ( .A(n68), .B(n1377), .Z(n1376) );
  XNOR U1369 ( .A(n1378), .B(n1375), .Z(n1377) );
  XOR U1370 ( .A(n1371), .B(n1221), .Z(n1373) );
  XOR U1371 ( .A(n1379), .B(n1380), .Z(n1221) );
  AND U1372 ( .A(n76), .B(n1381), .Z(n1380) );
  XOR U1373 ( .A(n1382), .B(n1383), .Z(n1371) );
  AND U1374 ( .A(n1384), .B(n1385), .Z(n1383) );
  XNOR U1375 ( .A(n1382), .B(n1328), .Z(n1385) );
  XNOR U1376 ( .A(n1386), .B(n1387), .Z(n1328) );
  AND U1377 ( .A(n68), .B(n1388), .Z(n1387) );
  XOR U1378 ( .A(n1389), .B(n1386), .Z(n1388) );
  XNOR U1379 ( .A(n1390), .B(n1382), .Z(n1384) );
  IV U1380 ( .A(n1233), .Z(n1390) );
  XOR U1381 ( .A(n1391), .B(n1392), .Z(n1233) );
  AND U1382 ( .A(n76), .B(n1393), .Z(n1392) );
  AND U1383 ( .A(n1349), .B(n1338), .Z(n1382) );
  XNOR U1384 ( .A(n1394), .B(n1395), .Z(n1338) );
  AND U1385 ( .A(n68), .B(n1396), .Z(n1395) );
  XNOR U1386 ( .A(n1397), .B(n1394), .Z(n1396) );
  XNOR U1387 ( .A(n1398), .B(n1399), .Z(n68) );
  NOR U1388 ( .A(n1400), .B(n1401), .Z(n1399) );
  XNOR U1389 ( .A(n1398), .B(n1360), .Z(n1401) );
  NOR U1390 ( .A(n1356), .B(n1357), .Z(n1360) );
  NOR U1391 ( .A(n1398), .B(n1359), .Z(n1400) );
  AND U1392 ( .A(n1402), .B(n1403), .Z(n1359) );
  XOR U1393 ( .A(n1404), .B(n1405), .Z(n1398) );
  AND U1394 ( .A(n1406), .B(n1407), .Z(n1405) );
  XNOR U1395 ( .A(n1404), .B(n1402), .Z(n1407) );
  IV U1396 ( .A(n1366), .Z(n1402) );
  XOR U1397 ( .A(n1408), .B(n1409), .Z(n1366) );
  XOR U1398 ( .A(n1410), .B(n1403), .Z(n1409) );
  AND U1399 ( .A(n1378), .B(n1411), .Z(n1403) );
  AND U1400 ( .A(n1412), .B(n1413), .Z(n1410) );
  XOR U1401 ( .A(n1414), .B(n1408), .Z(n1412) );
  XNOR U1402 ( .A(n1363), .B(n1404), .Z(n1406) );
  XNOR U1403 ( .A(n1415), .B(n1416), .Z(n1363) );
  AND U1404 ( .A(n72), .B(n1370), .Z(n1416) );
  XOR U1405 ( .A(n1415), .B(n1368), .Z(n1370) );
  XOR U1406 ( .A(n1417), .B(n1418), .Z(n1404) );
  AND U1407 ( .A(n1419), .B(n1420), .Z(n1418) );
  XNOR U1408 ( .A(n1417), .B(n1378), .Z(n1420) );
  XOR U1409 ( .A(n1421), .B(n1413), .Z(n1378) );
  XNOR U1410 ( .A(n1422), .B(n1408), .Z(n1413) );
  XOR U1411 ( .A(n1423), .B(n1424), .Z(n1408) );
  AND U1412 ( .A(n1425), .B(n1426), .Z(n1424) );
  XOR U1413 ( .A(n1427), .B(n1423), .Z(n1425) );
  XNOR U1414 ( .A(n1428), .B(n1429), .Z(n1422) );
  AND U1415 ( .A(n1430), .B(n1431), .Z(n1429) );
  XOR U1416 ( .A(n1428), .B(n1432), .Z(n1430) );
  XNOR U1417 ( .A(n1414), .B(n1411), .Z(n1421) );
  AND U1418 ( .A(n1433), .B(n1434), .Z(n1411) );
  XOR U1419 ( .A(n1435), .B(n1436), .Z(n1414) );
  AND U1420 ( .A(n1437), .B(n1438), .Z(n1436) );
  XOR U1421 ( .A(n1435), .B(n1439), .Z(n1437) );
  XNOR U1422 ( .A(n1375), .B(n1417), .Z(n1419) );
  XNOR U1423 ( .A(n1440), .B(n1441), .Z(n1375) );
  AND U1424 ( .A(n72), .B(n1381), .Z(n1441) );
  XOR U1425 ( .A(n1440), .B(n1379), .Z(n1381) );
  XOR U1426 ( .A(n1442), .B(n1443), .Z(n1417) );
  AND U1427 ( .A(n1444), .B(n1445), .Z(n1443) );
  XNOR U1428 ( .A(n1442), .B(n1433), .Z(n1445) );
  IV U1429 ( .A(n1389), .Z(n1433) );
  XNOR U1430 ( .A(n1446), .B(n1426), .Z(n1389) );
  XNOR U1431 ( .A(n1447), .B(n1432), .Z(n1426) );
  XOR U1432 ( .A(n1448), .B(n1449), .Z(n1432) );
  NOR U1433 ( .A(n1450), .B(n1451), .Z(n1449) );
  XNOR U1434 ( .A(n1448), .B(n1452), .Z(n1450) );
  XNOR U1435 ( .A(n1431), .B(n1423), .Z(n1447) );
  XOR U1436 ( .A(n1453), .B(n1454), .Z(n1423) );
  AND U1437 ( .A(n1455), .B(n1456), .Z(n1454) );
  XNOR U1438 ( .A(n1453), .B(n1457), .Z(n1455) );
  XNOR U1439 ( .A(n1458), .B(n1428), .Z(n1431) );
  XOR U1440 ( .A(n1459), .B(n1460), .Z(n1428) );
  AND U1441 ( .A(n1461), .B(n1462), .Z(n1460) );
  XOR U1442 ( .A(n1459), .B(n1463), .Z(n1461) );
  XNOR U1443 ( .A(n1464), .B(n1465), .Z(n1458) );
  NOR U1444 ( .A(n1466), .B(n1467), .Z(n1465) );
  XOR U1445 ( .A(n1464), .B(n1468), .Z(n1466) );
  XNOR U1446 ( .A(n1427), .B(n1434), .Z(n1446) );
  NOR U1447 ( .A(n1397), .B(n1469), .Z(n1434) );
  XOR U1448 ( .A(n1439), .B(n1438), .Z(n1427) );
  XNOR U1449 ( .A(n1470), .B(n1435), .Z(n1438) );
  XOR U1450 ( .A(n1471), .B(n1472), .Z(n1435) );
  AND U1451 ( .A(n1473), .B(n1474), .Z(n1472) );
  XOR U1452 ( .A(n1471), .B(n1475), .Z(n1473) );
  XNOR U1453 ( .A(n1476), .B(n1477), .Z(n1470) );
  NOR U1454 ( .A(n1478), .B(n1479), .Z(n1477) );
  XNOR U1455 ( .A(n1476), .B(n1480), .Z(n1478) );
  XOR U1456 ( .A(n1481), .B(n1482), .Z(n1439) );
  NOR U1457 ( .A(n1483), .B(n1484), .Z(n1482) );
  XNOR U1458 ( .A(n1481), .B(n1485), .Z(n1483) );
  XNOR U1459 ( .A(n1386), .B(n1442), .Z(n1444) );
  XNOR U1460 ( .A(n1486), .B(n1487), .Z(n1386) );
  AND U1461 ( .A(n72), .B(n1393), .Z(n1487) );
  XOR U1462 ( .A(n1486), .B(n1391), .Z(n1393) );
  AND U1463 ( .A(n1394), .B(n1397), .Z(n1442) );
  XOR U1464 ( .A(n1488), .B(n1469), .Z(n1397) );
  XNOR U1465 ( .A(p_input[128]), .B(p_input[48]), .Z(n1469) );
  XOR U1466 ( .A(n1457), .B(n1456), .Z(n1488) );
  XNOR U1467 ( .A(n1489), .B(n1463), .Z(n1456) );
  XNOR U1468 ( .A(n1452), .B(n1451), .Z(n1463) );
  XOR U1469 ( .A(n1490), .B(n1448), .Z(n1451) );
  XOR U1470 ( .A(p_input[138]), .B(p_input[58]), .Z(n1448) );
  XNOR U1471 ( .A(p_input[139]), .B(p_input[59]), .Z(n1490) );
  XOR U1472 ( .A(p_input[140]), .B(p_input[60]), .Z(n1452) );
  XNOR U1473 ( .A(n1462), .B(n1453), .Z(n1489) );
  XOR U1474 ( .A(p_input[129]), .B(p_input[49]), .Z(n1453) );
  XOR U1475 ( .A(n1491), .B(n1468), .Z(n1462) );
  XNOR U1476 ( .A(p_input[143]), .B(p_input[63]), .Z(n1468) );
  XOR U1477 ( .A(n1459), .B(n1467), .Z(n1491) );
  XOR U1478 ( .A(n1492), .B(n1464), .Z(n1467) );
  XOR U1479 ( .A(p_input[141]), .B(p_input[61]), .Z(n1464) );
  XNOR U1480 ( .A(p_input[142]), .B(p_input[62]), .Z(n1492) );
  XOR U1481 ( .A(p_input[137]), .B(p_input[57]), .Z(n1459) );
  XNOR U1482 ( .A(n1475), .B(n1474), .Z(n1457) );
  XNOR U1483 ( .A(n1493), .B(n1480), .Z(n1474) );
  XOR U1484 ( .A(p_input[136]), .B(p_input[56]), .Z(n1480) );
  XOR U1485 ( .A(n1471), .B(n1479), .Z(n1493) );
  XOR U1486 ( .A(n1494), .B(n1476), .Z(n1479) );
  XOR U1487 ( .A(p_input[134]), .B(p_input[54]), .Z(n1476) );
  XNOR U1488 ( .A(p_input[135]), .B(p_input[55]), .Z(n1494) );
  XOR U1489 ( .A(p_input[130]), .B(p_input[50]), .Z(n1471) );
  XNOR U1490 ( .A(n1485), .B(n1484), .Z(n1475) );
  XOR U1491 ( .A(n1495), .B(n1481), .Z(n1484) );
  XOR U1492 ( .A(p_input[131]), .B(p_input[51]), .Z(n1481) );
  XNOR U1493 ( .A(p_input[132]), .B(p_input[52]), .Z(n1495) );
  XOR U1494 ( .A(p_input[133]), .B(p_input[53]), .Z(n1485) );
  XNOR U1495 ( .A(n1496), .B(n1497), .Z(n1394) );
  AND U1496 ( .A(n72), .B(n1498), .Z(n1497) );
  XNOR U1497 ( .A(n1499), .B(n1500), .Z(n72) );
  NOR U1498 ( .A(n1501), .B(n1502), .Z(n1500) );
  XOR U1499 ( .A(n1357), .B(n1499), .Z(n1502) );
  NOR U1500 ( .A(n1499), .B(n1356), .Z(n1501) );
  XOR U1501 ( .A(n1503), .B(n1504), .Z(n1499) );
  AND U1502 ( .A(n1505), .B(n1506), .Z(n1504) );
  XOR U1503 ( .A(n1503), .B(n1368), .Z(n1505) );
  XOR U1504 ( .A(n1507), .B(n1508), .Z(n1349) );
  AND U1505 ( .A(n76), .B(n1498), .Z(n1508) );
  XNOR U1506 ( .A(n1496), .B(n1507), .Z(n1498) );
  XNOR U1507 ( .A(n1509), .B(n1510), .Z(n76) );
  NOR U1508 ( .A(n1511), .B(n1512), .Z(n1510) );
  XNOR U1509 ( .A(n1357), .B(n1513), .Z(n1512) );
  IV U1510 ( .A(n1509), .Z(n1513) );
  AND U1511 ( .A(n1514), .B(n1515), .Z(n1357) );
  NOR U1512 ( .A(n1509), .B(n1356), .Z(n1511) );
  AND U1513 ( .A(n1516), .B(n1517), .Z(n1356) );
  IV U1514 ( .A(n1518), .Z(n1516) );
  XOR U1515 ( .A(n1503), .B(n1519), .Z(n1509) );
  AND U1516 ( .A(n1520), .B(n1506), .Z(n1519) );
  XNOR U1517 ( .A(n1415), .B(n1503), .Z(n1506) );
  XNOR U1518 ( .A(n1521), .B(n1522), .Z(n1415) );
  AND U1519 ( .A(n79), .B(n1523), .Z(n1522) );
  XOR U1520 ( .A(n1524), .B(n1521), .Z(n1523) );
  XNOR U1521 ( .A(n1525), .B(n1503), .Z(n1520) );
  IV U1522 ( .A(n1368), .Z(n1525) );
  XOR U1523 ( .A(n1526), .B(n1527), .Z(n1368) );
  AND U1524 ( .A(n87), .B(n1528), .Z(n1527) );
  XOR U1525 ( .A(n1529), .B(n1530), .Z(n1503) );
  AND U1526 ( .A(n1531), .B(n1532), .Z(n1530) );
  XNOR U1527 ( .A(n1440), .B(n1529), .Z(n1532) );
  XNOR U1528 ( .A(n1533), .B(n1534), .Z(n1440) );
  AND U1529 ( .A(n79), .B(n1535), .Z(n1534) );
  XNOR U1530 ( .A(n1536), .B(n1533), .Z(n1535) );
  XOR U1531 ( .A(n1529), .B(n1379), .Z(n1531) );
  XOR U1532 ( .A(n1537), .B(n1538), .Z(n1379) );
  AND U1533 ( .A(n87), .B(n1539), .Z(n1538) );
  XOR U1534 ( .A(n1540), .B(n1541), .Z(n1529) );
  AND U1535 ( .A(n1542), .B(n1543), .Z(n1541) );
  XNOR U1536 ( .A(n1540), .B(n1486), .Z(n1543) );
  XNOR U1537 ( .A(n1544), .B(n1545), .Z(n1486) );
  AND U1538 ( .A(n79), .B(n1546), .Z(n1545) );
  XOR U1539 ( .A(n1547), .B(n1544), .Z(n1546) );
  XNOR U1540 ( .A(n1548), .B(n1540), .Z(n1542) );
  IV U1541 ( .A(n1391), .Z(n1548) );
  XOR U1542 ( .A(n1549), .B(n1550), .Z(n1391) );
  AND U1543 ( .A(n87), .B(n1551), .Z(n1550) );
  AND U1544 ( .A(n1507), .B(n1496), .Z(n1540) );
  XNOR U1545 ( .A(n1552), .B(n1553), .Z(n1496) );
  AND U1546 ( .A(n79), .B(n1554), .Z(n1553) );
  XNOR U1547 ( .A(n1555), .B(n1552), .Z(n1554) );
  XNOR U1548 ( .A(n1556), .B(n1557), .Z(n79) );
  NOR U1549 ( .A(n1558), .B(n1559), .Z(n1557) );
  XNOR U1550 ( .A(n1556), .B(n1518), .Z(n1559) );
  NOR U1551 ( .A(n1514), .B(n1515), .Z(n1518) );
  NOR U1552 ( .A(n1556), .B(n1517), .Z(n1558) );
  AND U1553 ( .A(n1560), .B(n1561), .Z(n1517) );
  XOR U1554 ( .A(n1562), .B(n1563), .Z(n1556) );
  AND U1555 ( .A(n1564), .B(n1565), .Z(n1563) );
  XNOR U1556 ( .A(n1562), .B(n1560), .Z(n1565) );
  IV U1557 ( .A(n1524), .Z(n1560) );
  XOR U1558 ( .A(n1566), .B(n1567), .Z(n1524) );
  XOR U1559 ( .A(n1568), .B(n1561), .Z(n1567) );
  AND U1560 ( .A(n1536), .B(n1569), .Z(n1561) );
  AND U1561 ( .A(n1570), .B(n1571), .Z(n1568) );
  XOR U1562 ( .A(n1572), .B(n1566), .Z(n1570) );
  XNOR U1563 ( .A(n1521), .B(n1562), .Z(n1564) );
  XNOR U1564 ( .A(n1573), .B(n1574), .Z(n1521) );
  AND U1565 ( .A(n83), .B(n1528), .Z(n1574) );
  XOR U1566 ( .A(n1573), .B(n1526), .Z(n1528) );
  XOR U1567 ( .A(n1575), .B(n1576), .Z(n1562) );
  AND U1568 ( .A(n1577), .B(n1578), .Z(n1576) );
  XNOR U1569 ( .A(n1575), .B(n1536), .Z(n1578) );
  XOR U1570 ( .A(n1579), .B(n1571), .Z(n1536) );
  XNOR U1571 ( .A(n1580), .B(n1566), .Z(n1571) );
  XOR U1572 ( .A(n1581), .B(n1582), .Z(n1566) );
  AND U1573 ( .A(n1583), .B(n1584), .Z(n1582) );
  XOR U1574 ( .A(n1585), .B(n1581), .Z(n1583) );
  XNOR U1575 ( .A(n1586), .B(n1587), .Z(n1580) );
  AND U1576 ( .A(n1588), .B(n1589), .Z(n1587) );
  XOR U1577 ( .A(n1586), .B(n1590), .Z(n1588) );
  XNOR U1578 ( .A(n1572), .B(n1569), .Z(n1579) );
  AND U1579 ( .A(n1591), .B(n1592), .Z(n1569) );
  XOR U1580 ( .A(n1593), .B(n1594), .Z(n1572) );
  AND U1581 ( .A(n1595), .B(n1596), .Z(n1594) );
  XOR U1582 ( .A(n1593), .B(n1597), .Z(n1595) );
  XNOR U1583 ( .A(n1533), .B(n1575), .Z(n1577) );
  XNOR U1584 ( .A(n1598), .B(n1599), .Z(n1533) );
  AND U1585 ( .A(n83), .B(n1539), .Z(n1599) );
  XOR U1586 ( .A(n1598), .B(n1537), .Z(n1539) );
  XOR U1587 ( .A(n1600), .B(n1601), .Z(n1575) );
  AND U1588 ( .A(n1602), .B(n1603), .Z(n1601) );
  XNOR U1589 ( .A(n1600), .B(n1591), .Z(n1603) );
  IV U1590 ( .A(n1547), .Z(n1591) );
  XNOR U1591 ( .A(n1604), .B(n1584), .Z(n1547) );
  XNOR U1592 ( .A(n1605), .B(n1590), .Z(n1584) );
  XOR U1593 ( .A(n1606), .B(n1607), .Z(n1590) );
  NOR U1594 ( .A(n1608), .B(n1609), .Z(n1607) );
  XNOR U1595 ( .A(n1606), .B(n1610), .Z(n1608) );
  XNOR U1596 ( .A(n1589), .B(n1581), .Z(n1605) );
  XOR U1597 ( .A(n1611), .B(n1612), .Z(n1581) );
  AND U1598 ( .A(n1613), .B(n1614), .Z(n1612) );
  XNOR U1599 ( .A(n1611), .B(n1615), .Z(n1613) );
  XNOR U1600 ( .A(n1616), .B(n1586), .Z(n1589) );
  XOR U1601 ( .A(n1617), .B(n1618), .Z(n1586) );
  AND U1602 ( .A(n1619), .B(n1620), .Z(n1618) );
  XOR U1603 ( .A(n1617), .B(n1621), .Z(n1619) );
  XNOR U1604 ( .A(n1622), .B(n1623), .Z(n1616) );
  NOR U1605 ( .A(n1624), .B(n1625), .Z(n1623) );
  XOR U1606 ( .A(n1622), .B(n1626), .Z(n1624) );
  XNOR U1607 ( .A(n1585), .B(n1592), .Z(n1604) );
  NOR U1608 ( .A(n1555), .B(n1627), .Z(n1592) );
  XOR U1609 ( .A(n1597), .B(n1596), .Z(n1585) );
  XNOR U1610 ( .A(n1628), .B(n1593), .Z(n1596) );
  XOR U1611 ( .A(n1629), .B(n1630), .Z(n1593) );
  AND U1612 ( .A(n1631), .B(n1632), .Z(n1630) );
  XOR U1613 ( .A(n1629), .B(n1633), .Z(n1631) );
  XNOR U1614 ( .A(n1634), .B(n1635), .Z(n1628) );
  NOR U1615 ( .A(n1636), .B(n1637), .Z(n1635) );
  XNOR U1616 ( .A(n1634), .B(n1638), .Z(n1636) );
  XOR U1617 ( .A(n1639), .B(n1640), .Z(n1597) );
  NOR U1618 ( .A(n1641), .B(n1642), .Z(n1640) );
  XNOR U1619 ( .A(n1639), .B(n1643), .Z(n1641) );
  XNOR U1620 ( .A(n1544), .B(n1600), .Z(n1602) );
  XNOR U1621 ( .A(n1644), .B(n1645), .Z(n1544) );
  AND U1622 ( .A(n83), .B(n1551), .Z(n1645) );
  XOR U1623 ( .A(n1644), .B(n1549), .Z(n1551) );
  AND U1624 ( .A(n1552), .B(n1555), .Z(n1600) );
  XOR U1625 ( .A(n1646), .B(n1627), .Z(n1555) );
  XNOR U1626 ( .A(p_input[128]), .B(p_input[64]), .Z(n1627) );
  XOR U1627 ( .A(n1615), .B(n1614), .Z(n1646) );
  XNOR U1628 ( .A(n1647), .B(n1621), .Z(n1614) );
  XNOR U1629 ( .A(n1610), .B(n1609), .Z(n1621) );
  XOR U1630 ( .A(n1648), .B(n1606), .Z(n1609) );
  XOR U1631 ( .A(p_input[138]), .B(p_input[74]), .Z(n1606) );
  XNOR U1632 ( .A(p_input[139]), .B(p_input[75]), .Z(n1648) );
  XOR U1633 ( .A(p_input[140]), .B(p_input[76]), .Z(n1610) );
  XNOR U1634 ( .A(n1620), .B(n1611), .Z(n1647) );
  XOR U1635 ( .A(p_input[129]), .B(p_input[65]), .Z(n1611) );
  XOR U1636 ( .A(n1649), .B(n1626), .Z(n1620) );
  XNOR U1637 ( .A(p_input[143]), .B(p_input[79]), .Z(n1626) );
  XOR U1638 ( .A(n1617), .B(n1625), .Z(n1649) );
  XOR U1639 ( .A(n1650), .B(n1622), .Z(n1625) );
  XOR U1640 ( .A(p_input[141]), .B(p_input[77]), .Z(n1622) );
  XNOR U1641 ( .A(p_input[142]), .B(p_input[78]), .Z(n1650) );
  XOR U1642 ( .A(p_input[137]), .B(p_input[73]), .Z(n1617) );
  XNOR U1643 ( .A(n1633), .B(n1632), .Z(n1615) );
  XNOR U1644 ( .A(n1651), .B(n1638), .Z(n1632) );
  XOR U1645 ( .A(p_input[136]), .B(p_input[72]), .Z(n1638) );
  XOR U1646 ( .A(n1629), .B(n1637), .Z(n1651) );
  XOR U1647 ( .A(n1652), .B(n1634), .Z(n1637) );
  XOR U1648 ( .A(p_input[134]), .B(p_input[70]), .Z(n1634) );
  XNOR U1649 ( .A(p_input[135]), .B(p_input[71]), .Z(n1652) );
  XOR U1650 ( .A(p_input[130]), .B(p_input[66]), .Z(n1629) );
  XNOR U1651 ( .A(n1643), .B(n1642), .Z(n1633) );
  XOR U1652 ( .A(n1653), .B(n1639), .Z(n1642) );
  XOR U1653 ( .A(p_input[131]), .B(p_input[67]), .Z(n1639) );
  XNOR U1654 ( .A(p_input[132]), .B(p_input[68]), .Z(n1653) );
  XOR U1655 ( .A(p_input[133]), .B(p_input[69]), .Z(n1643) );
  XNOR U1656 ( .A(n1654), .B(n1655), .Z(n1552) );
  AND U1657 ( .A(n83), .B(n1656), .Z(n1655) );
  XNOR U1658 ( .A(n1657), .B(n1658), .Z(n83) );
  NOR U1659 ( .A(n1659), .B(n1660), .Z(n1658) );
  XOR U1660 ( .A(n1515), .B(n1657), .Z(n1660) );
  NOR U1661 ( .A(n1657), .B(n1514), .Z(n1659) );
  XOR U1662 ( .A(n1661), .B(n1662), .Z(n1657) );
  AND U1663 ( .A(n1663), .B(n1664), .Z(n1662) );
  XOR U1664 ( .A(n1661), .B(n1526), .Z(n1663) );
  XOR U1665 ( .A(n1665), .B(n1666), .Z(n1507) );
  AND U1666 ( .A(n87), .B(n1656), .Z(n1666) );
  XNOR U1667 ( .A(n1654), .B(n1665), .Z(n1656) );
  XNOR U1668 ( .A(n1667), .B(n1668), .Z(n87) );
  NOR U1669 ( .A(n1669), .B(n1670), .Z(n1668) );
  XNOR U1670 ( .A(n1515), .B(n1671), .Z(n1670) );
  IV U1671 ( .A(n1667), .Z(n1671) );
  AND U1672 ( .A(n1672), .B(n1673), .Z(n1515) );
  NOR U1673 ( .A(n1667), .B(n1514), .Z(n1669) );
  AND U1674 ( .A(n1674), .B(n1675), .Z(n1514) );
  IV U1675 ( .A(n1676), .Z(n1674) );
  XOR U1676 ( .A(n1661), .B(n1677), .Z(n1667) );
  AND U1677 ( .A(n1678), .B(n1664), .Z(n1677) );
  XNOR U1678 ( .A(n1573), .B(n1661), .Z(n1664) );
  XNOR U1679 ( .A(n1679), .B(n1680), .Z(n1573) );
  AND U1680 ( .A(n90), .B(n1681), .Z(n1680) );
  XOR U1681 ( .A(n1682), .B(n1679), .Z(n1681) );
  XNOR U1682 ( .A(n1683), .B(n1661), .Z(n1678) );
  IV U1683 ( .A(n1526), .Z(n1683) );
  XOR U1684 ( .A(n1684), .B(n1685), .Z(n1526) );
  AND U1685 ( .A(n97), .B(n1686), .Z(n1685) );
  XOR U1686 ( .A(n1687), .B(n1688), .Z(n1661) );
  AND U1687 ( .A(n1689), .B(n1690), .Z(n1688) );
  XNOR U1688 ( .A(n1598), .B(n1687), .Z(n1690) );
  XNOR U1689 ( .A(n1691), .B(n1692), .Z(n1598) );
  AND U1690 ( .A(n90), .B(n1693), .Z(n1692) );
  XNOR U1691 ( .A(n1694), .B(n1691), .Z(n1693) );
  XOR U1692 ( .A(n1687), .B(n1537), .Z(n1689) );
  XOR U1693 ( .A(n1695), .B(n1696), .Z(n1537) );
  AND U1694 ( .A(n97), .B(n1697), .Z(n1696) );
  XOR U1695 ( .A(n1698), .B(n1699), .Z(n1687) );
  AND U1696 ( .A(n1700), .B(n1701), .Z(n1699) );
  XNOR U1697 ( .A(n1698), .B(n1644), .Z(n1701) );
  XNOR U1698 ( .A(n1702), .B(n1703), .Z(n1644) );
  AND U1699 ( .A(n90), .B(n1704), .Z(n1703) );
  XOR U1700 ( .A(n1705), .B(n1702), .Z(n1704) );
  XNOR U1701 ( .A(n1706), .B(n1698), .Z(n1700) );
  IV U1702 ( .A(n1549), .Z(n1706) );
  XOR U1703 ( .A(n1707), .B(n1708), .Z(n1549) );
  AND U1704 ( .A(n97), .B(n1709), .Z(n1708) );
  AND U1705 ( .A(n1665), .B(n1654), .Z(n1698) );
  XNOR U1706 ( .A(n1710), .B(n1711), .Z(n1654) );
  AND U1707 ( .A(n90), .B(n1712), .Z(n1711) );
  XNOR U1708 ( .A(n1713), .B(n1710), .Z(n1712) );
  XNOR U1709 ( .A(n1714), .B(n1715), .Z(n90) );
  NOR U1710 ( .A(n1716), .B(n1717), .Z(n1715) );
  XNOR U1711 ( .A(n1714), .B(n1676), .Z(n1717) );
  NOR U1712 ( .A(n1672), .B(n1673), .Z(n1676) );
  NOR U1713 ( .A(n1714), .B(n1675), .Z(n1716) );
  AND U1714 ( .A(n1718), .B(n1719), .Z(n1675) );
  XOR U1715 ( .A(n1720), .B(n1721), .Z(n1714) );
  AND U1716 ( .A(n1722), .B(n1723), .Z(n1721) );
  XNOR U1717 ( .A(n1720), .B(n1718), .Z(n1723) );
  IV U1718 ( .A(n1682), .Z(n1718) );
  XOR U1719 ( .A(n1724), .B(n1725), .Z(n1682) );
  XOR U1720 ( .A(n1726), .B(n1719), .Z(n1725) );
  AND U1721 ( .A(n1694), .B(n1727), .Z(n1719) );
  AND U1722 ( .A(n1728), .B(n1729), .Z(n1726) );
  XOR U1723 ( .A(n1730), .B(n1724), .Z(n1728) );
  XNOR U1724 ( .A(n1679), .B(n1720), .Z(n1722) );
  XNOR U1725 ( .A(n1731), .B(n1732), .Z(n1679) );
  AND U1726 ( .A(n94), .B(n1686), .Z(n1732) );
  XOR U1727 ( .A(n1731), .B(n1684), .Z(n1686) );
  XOR U1728 ( .A(n1733), .B(n1734), .Z(n1720) );
  AND U1729 ( .A(n1735), .B(n1736), .Z(n1734) );
  XNOR U1730 ( .A(n1733), .B(n1694), .Z(n1736) );
  XOR U1731 ( .A(n1737), .B(n1729), .Z(n1694) );
  XNOR U1732 ( .A(n1738), .B(n1724), .Z(n1729) );
  XOR U1733 ( .A(n1739), .B(n1740), .Z(n1724) );
  AND U1734 ( .A(n1741), .B(n1742), .Z(n1740) );
  XOR U1735 ( .A(n1743), .B(n1739), .Z(n1741) );
  XNOR U1736 ( .A(n1744), .B(n1745), .Z(n1738) );
  AND U1737 ( .A(n1746), .B(n1747), .Z(n1745) );
  XOR U1738 ( .A(n1744), .B(n1748), .Z(n1746) );
  XNOR U1739 ( .A(n1730), .B(n1727), .Z(n1737) );
  AND U1740 ( .A(n1749), .B(n1750), .Z(n1727) );
  XOR U1741 ( .A(n1751), .B(n1752), .Z(n1730) );
  AND U1742 ( .A(n1753), .B(n1754), .Z(n1752) );
  XOR U1743 ( .A(n1751), .B(n1755), .Z(n1753) );
  XNOR U1744 ( .A(n1691), .B(n1733), .Z(n1735) );
  XNOR U1745 ( .A(n1756), .B(n1757), .Z(n1691) );
  AND U1746 ( .A(n94), .B(n1697), .Z(n1757) );
  XOR U1747 ( .A(n1756), .B(n1695), .Z(n1697) );
  XOR U1748 ( .A(n1758), .B(n1759), .Z(n1733) );
  AND U1749 ( .A(n1760), .B(n1761), .Z(n1759) );
  XNOR U1750 ( .A(n1758), .B(n1749), .Z(n1761) );
  IV U1751 ( .A(n1705), .Z(n1749) );
  XNOR U1752 ( .A(n1762), .B(n1742), .Z(n1705) );
  XNOR U1753 ( .A(n1763), .B(n1748), .Z(n1742) );
  XOR U1754 ( .A(n1764), .B(n1765), .Z(n1748) );
  NOR U1755 ( .A(n1766), .B(n1767), .Z(n1765) );
  XNOR U1756 ( .A(n1764), .B(n1768), .Z(n1766) );
  XNOR U1757 ( .A(n1747), .B(n1739), .Z(n1763) );
  XOR U1758 ( .A(n1769), .B(n1770), .Z(n1739) );
  AND U1759 ( .A(n1771), .B(n1772), .Z(n1770) );
  XNOR U1760 ( .A(n1769), .B(n1773), .Z(n1771) );
  XNOR U1761 ( .A(n1774), .B(n1744), .Z(n1747) );
  XOR U1762 ( .A(n1775), .B(n1776), .Z(n1744) );
  AND U1763 ( .A(n1777), .B(n1778), .Z(n1776) );
  XOR U1764 ( .A(n1775), .B(n1779), .Z(n1777) );
  XNOR U1765 ( .A(n1780), .B(n1781), .Z(n1774) );
  NOR U1766 ( .A(n1782), .B(n1783), .Z(n1781) );
  XOR U1767 ( .A(n1780), .B(n1784), .Z(n1782) );
  XNOR U1768 ( .A(n1743), .B(n1750), .Z(n1762) );
  NOR U1769 ( .A(n1713), .B(n1785), .Z(n1750) );
  XOR U1770 ( .A(n1755), .B(n1754), .Z(n1743) );
  XNOR U1771 ( .A(n1786), .B(n1751), .Z(n1754) );
  XOR U1772 ( .A(n1787), .B(n1788), .Z(n1751) );
  AND U1773 ( .A(n1789), .B(n1790), .Z(n1788) );
  XOR U1774 ( .A(n1787), .B(n1791), .Z(n1789) );
  XNOR U1775 ( .A(n1792), .B(n1793), .Z(n1786) );
  NOR U1776 ( .A(n1794), .B(n1795), .Z(n1793) );
  XNOR U1777 ( .A(n1792), .B(n1796), .Z(n1794) );
  XOR U1778 ( .A(n1797), .B(n1798), .Z(n1755) );
  NOR U1779 ( .A(n1799), .B(n1800), .Z(n1798) );
  XNOR U1780 ( .A(n1797), .B(n1801), .Z(n1799) );
  XNOR U1781 ( .A(n1702), .B(n1758), .Z(n1760) );
  XNOR U1782 ( .A(n1802), .B(n1803), .Z(n1702) );
  AND U1783 ( .A(n94), .B(n1709), .Z(n1803) );
  XOR U1784 ( .A(n1802), .B(n1707), .Z(n1709) );
  AND U1785 ( .A(n1710), .B(n1713), .Z(n1758) );
  XOR U1786 ( .A(n1804), .B(n1785), .Z(n1713) );
  XNOR U1787 ( .A(p_input[128]), .B(p_input[80]), .Z(n1785) );
  XOR U1788 ( .A(n1773), .B(n1772), .Z(n1804) );
  XNOR U1789 ( .A(n1805), .B(n1779), .Z(n1772) );
  XNOR U1790 ( .A(n1768), .B(n1767), .Z(n1779) );
  XOR U1791 ( .A(n1806), .B(n1764), .Z(n1767) );
  XOR U1792 ( .A(p_input[138]), .B(p_input[90]), .Z(n1764) );
  XNOR U1793 ( .A(p_input[139]), .B(p_input[91]), .Z(n1806) );
  XOR U1794 ( .A(p_input[140]), .B(p_input[92]), .Z(n1768) );
  XNOR U1795 ( .A(n1778), .B(n1769), .Z(n1805) );
  XOR U1796 ( .A(p_input[129]), .B(p_input[81]), .Z(n1769) );
  XOR U1797 ( .A(n1807), .B(n1784), .Z(n1778) );
  XNOR U1798 ( .A(p_input[143]), .B(p_input[95]), .Z(n1784) );
  XOR U1799 ( .A(n1775), .B(n1783), .Z(n1807) );
  XOR U1800 ( .A(n1808), .B(n1780), .Z(n1783) );
  XOR U1801 ( .A(p_input[141]), .B(p_input[93]), .Z(n1780) );
  XNOR U1802 ( .A(p_input[142]), .B(p_input[94]), .Z(n1808) );
  XOR U1803 ( .A(p_input[137]), .B(p_input[89]), .Z(n1775) );
  XNOR U1804 ( .A(n1791), .B(n1790), .Z(n1773) );
  XNOR U1805 ( .A(n1809), .B(n1796), .Z(n1790) );
  XOR U1806 ( .A(p_input[136]), .B(p_input[88]), .Z(n1796) );
  XOR U1807 ( .A(n1787), .B(n1795), .Z(n1809) );
  XOR U1808 ( .A(n1810), .B(n1792), .Z(n1795) );
  XOR U1809 ( .A(p_input[134]), .B(p_input[86]), .Z(n1792) );
  XNOR U1810 ( .A(p_input[135]), .B(p_input[87]), .Z(n1810) );
  XOR U1811 ( .A(p_input[130]), .B(p_input[82]), .Z(n1787) );
  XNOR U1812 ( .A(n1801), .B(n1800), .Z(n1791) );
  XOR U1813 ( .A(n1811), .B(n1797), .Z(n1800) );
  XOR U1814 ( .A(p_input[131]), .B(p_input[83]), .Z(n1797) );
  XNOR U1815 ( .A(p_input[132]), .B(p_input[84]), .Z(n1811) );
  XOR U1816 ( .A(p_input[133]), .B(p_input[85]), .Z(n1801) );
  XNOR U1817 ( .A(n1812), .B(n1813), .Z(n1710) );
  AND U1818 ( .A(n94), .B(n1814), .Z(n1813) );
  XNOR U1819 ( .A(n1815), .B(n1816), .Z(n94) );
  NOR U1820 ( .A(n1817), .B(n1818), .Z(n1816) );
  XOR U1821 ( .A(n1673), .B(n1815), .Z(n1818) );
  NOR U1822 ( .A(n1815), .B(n1672), .Z(n1817) );
  XOR U1823 ( .A(n1819), .B(n1820), .Z(n1815) );
  AND U1824 ( .A(n1821), .B(n1822), .Z(n1820) );
  XOR U1825 ( .A(n1819), .B(n1684), .Z(n1821) );
  XOR U1826 ( .A(n1823), .B(n1824), .Z(n1665) );
  AND U1827 ( .A(n97), .B(n1814), .Z(n1824) );
  XOR U1828 ( .A(n1825), .B(n1823), .Z(n1814) );
  XNOR U1829 ( .A(n1826), .B(n1827), .Z(n97) );
  NOR U1830 ( .A(n1828), .B(n1829), .Z(n1827) );
  XNOR U1831 ( .A(n1673), .B(n1830), .Z(n1829) );
  IV U1832 ( .A(n1826), .Z(n1830) );
  AND U1833 ( .A(n1684), .B(n1831), .Z(n1673) );
  NOR U1834 ( .A(n1826), .B(n1672), .Z(n1828) );
  AND U1835 ( .A(n1731), .B(n1832), .Z(n1672) );
  XOR U1836 ( .A(n1819), .B(n1833), .Z(n1826) );
  AND U1837 ( .A(n1834), .B(n1822), .Z(n1833) );
  XNOR U1838 ( .A(n1731), .B(n1819), .Z(n1822) );
  XNOR U1839 ( .A(n1835), .B(n1836), .Z(n1731) );
  XOR U1840 ( .A(n1837), .B(n1832), .Z(n1836) );
  AND U1841 ( .A(n1756), .B(n1838), .Z(n1832) );
  AND U1842 ( .A(n1839), .B(n1840), .Z(n1837) );
  XOR U1843 ( .A(n1841), .B(n1835), .Z(n1839) );
  XNOR U1844 ( .A(n1842), .B(n1819), .Z(n1834) );
  IV U1845 ( .A(n1684), .Z(n1842) );
  XNOR U1846 ( .A(n1843), .B(n1844), .Z(n1684) );
  XOR U1847 ( .A(n1845), .B(n1831), .Z(n1844) );
  AND U1848 ( .A(n1695), .B(n1846), .Z(n1831) );
  AND U1849 ( .A(n1847), .B(n1848), .Z(n1845) );
  XNOR U1850 ( .A(n1843), .B(n1849), .Z(n1847) );
  XOR U1851 ( .A(n1850), .B(n1851), .Z(n1819) );
  AND U1852 ( .A(n1852), .B(n1853), .Z(n1851) );
  XNOR U1853 ( .A(n1756), .B(n1850), .Z(n1853) );
  XOR U1854 ( .A(n1854), .B(n1840), .Z(n1756) );
  XNOR U1855 ( .A(n1855), .B(n1835), .Z(n1840) );
  XOR U1856 ( .A(n1856), .B(n1857), .Z(n1835) );
  AND U1857 ( .A(n1858), .B(n1859), .Z(n1857) );
  XOR U1858 ( .A(n1860), .B(n1856), .Z(n1858) );
  XNOR U1859 ( .A(n1861), .B(n1862), .Z(n1855) );
  AND U1860 ( .A(n1863), .B(n1864), .Z(n1862) );
  XOR U1861 ( .A(n1861), .B(n1865), .Z(n1863) );
  XNOR U1862 ( .A(n1841), .B(n1838), .Z(n1854) );
  AND U1863 ( .A(n1802), .B(n1866), .Z(n1838) );
  XOR U1864 ( .A(n1867), .B(n1868), .Z(n1841) );
  AND U1865 ( .A(n1869), .B(n1870), .Z(n1868) );
  XOR U1866 ( .A(n1867), .B(n1871), .Z(n1869) );
  XOR U1867 ( .A(n1850), .B(n1695), .Z(n1852) );
  XNOR U1868 ( .A(n1872), .B(n1849), .Z(n1695) );
  XNOR U1869 ( .A(n1873), .B(n1874), .Z(n1849) );
  AND U1870 ( .A(n1875), .B(n1876), .Z(n1874) );
  XOR U1871 ( .A(n1873), .B(n1877), .Z(n1875) );
  XNOR U1872 ( .A(n1848), .B(n1846), .Z(n1872) );
  AND U1873 ( .A(n1707), .B(n1878), .Z(n1846) );
  XNOR U1874 ( .A(n1879), .B(n1843), .Z(n1848) );
  XOR U1875 ( .A(n1880), .B(n1881), .Z(n1843) );
  AND U1876 ( .A(n1882), .B(n1883), .Z(n1881) );
  XOR U1877 ( .A(n1880), .B(n1884), .Z(n1882) );
  XNOR U1878 ( .A(n1885), .B(n1886), .Z(n1879) );
  AND U1879 ( .A(n1887), .B(n1888), .Z(n1886) );
  XNOR U1880 ( .A(n1885), .B(n1889), .Z(n1887) );
  XOR U1881 ( .A(n1890), .B(n1891), .Z(n1850) );
  AND U1882 ( .A(n1892), .B(n1893), .Z(n1891) );
  XNOR U1883 ( .A(n1890), .B(n1802), .Z(n1893) );
  XOR U1884 ( .A(n1894), .B(n1859), .Z(n1802) );
  XNOR U1885 ( .A(n1895), .B(n1865), .Z(n1859) );
  XOR U1886 ( .A(n1896), .B(n1897), .Z(n1865) );
  NOR U1887 ( .A(n1898), .B(n1899), .Z(n1897) );
  XNOR U1888 ( .A(n1896), .B(n1900), .Z(n1898) );
  XNOR U1889 ( .A(n1864), .B(n1856), .Z(n1895) );
  XOR U1890 ( .A(n1901), .B(n1902), .Z(n1856) );
  AND U1891 ( .A(n1903), .B(n1904), .Z(n1902) );
  XNOR U1892 ( .A(n1901), .B(n1905), .Z(n1903) );
  XNOR U1893 ( .A(n1906), .B(n1861), .Z(n1864) );
  XOR U1894 ( .A(n1907), .B(n1908), .Z(n1861) );
  AND U1895 ( .A(n1909), .B(n1910), .Z(n1908) );
  XNOR U1896 ( .A(n1911), .B(n1912), .Z(n1909) );
  XNOR U1897 ( .A(n1913), .B(n1914), .Z(n1906) );
  NOR U1898 ( .A(n1915), .B(n1916), .Z(n1914) );
  XOR U1899 ( .A(n1913), .B(n1917), .Z(n1915) );
  XNOR U1900 ( .A(n1860), .B(n1866), .Z(n1894) );
  AND U1901 ( .A(n1825), .B(n1918), .Z(n1866) );
  IV U1902 ( .A(n1812), .Z(n1825) );
  XOR U1903 ( .A(n1871), .B(n1870), .Z(n1860) );
  XNOR U1904 ( .A(n1919), .B(n1867), .Z(n1870) );
  XOR U1905 ( .A(n1920), .B(n1921), .Z(n1867) );
  AND U1906 ( .A(n1922), .B(n1923), .Z(n1921) );
  XNOR U1907 ( .A(n1924), .B(n1925), .Z(n1922) );
  XNOR U1908 ( .A(n1926), .B(n1927), .Z(n1919) );
  AND U1909 ( .A(n1928), .B(n1929), .Z(n1927) );
  XNOR U1910 ( .A(n1926), .B(n1930), .Z(n1928) );
  XOR U1911 ( .A(n1931), .B(n1932), .Z(n1871) );
  AND U1912 ( .A(n1933), .B(n1934), .Z(n1932) );
  XOR U1913 ( .A(n1931), .B(n1935), .Z(n1933) );
  XNOR U1914 ( .A(n1936), .B(n1890), .Z(n1892) );
  IV U1915 ( .A(n1707), .Z(n1936) );
  XOR U1916 ( .A(n1937), .B(n1884), .Z(n1707) );
  XOR U1917 ( .A(n1877), .B(n1876), .Z(n1884) );
  XNOR U1918 ( .A(n1938), .B(n1873), .Z(n1876) );
  XOR U1919 ( .A(n1939), .B(n1940), .Z(n1873) );
  AND U1920 ( .A(n1941), .B(n1942), .Z(n1940) );
  XOR U1921 ( .A(n1939), .B(n1943), .Z(n1941) );
  XNOR U1922 ( .A(n1944), .B(n1945), .Z(n1938) );
  NOR U1923 ( .A(n1946), .B(n1947), .Z(n1945) );
  XNOR U1924 ( .A(n1944), .B(n1948), .Z(n1946) );
  XOR U1925 ( .A(n1949), .B(n1950), .Z(n1877) );
  NOR U1926 ( .A(n1951), .B(n1952), .Z(n1950) );
  XNOR U1927 ( .A(n1949), .B(n1953), .Z(n1951) );
  XNOR U1928 ( .A(n1883), .B(n1878), .Z(n1937) );
  AND U1929 ( .A(n1823), .B(n1954), .Z(n1878) );
  XOR U1930 ( .A(n1955), .B(n1889), .Z(n1883) );
  XNOR U1931 ( .A(n1956), .B(n1957), .Z(n1889) );
  NOR U1932 ( .A(n1958), .B(n1959), .Z(n1957) );
  XNOR U1933 ( .A(n1956), .B(n1960), .Z(n1958) );
  XNOR U1934 ( .A(n1888), .B(n1880), .Z(n1955) );
  XOR U1935 ( .A(n1961), .B(n1962), .Z(n1880) );
  AND U1936 ( .A(n1963), .B(n1964), .Z(n1962) );
  XOR U1937 ( .A(n1961), .B(n1965), .Z(n1963) );
  XNOR U1938 ( .A(n1966), .B(n1885), .Z(n1888) );
  XOR U1939 ( .A(n1967), .B(n1968), .Z(n1885) );
  AND U1940 ( .A(n1969), .B(n1970), .Z(n1968) );
  XOR U1941 ( .A(n1967), .B(n1971), .Z(n1969) );
  XNOR U1942 ( .A(n1972), .B(n1973), .Z(n1966) );
  NOR U1943 ( .A(n1974), .B(n1975), .Z(n1973) );
  XOR U1944 ( .A(n1972), .B(n1976), .Z(n1974) );
  AND U1945 ( .A(n1823), .B(n1812), .Z(n1890) );
  XNOR U1946 ( .A(n1977), .B(n1918), .Z(n1812) );
  XOR U1947 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(
        p_input[128]), .Z(n1918) );
  XOR U1948 ( .A(n1905), .B(n1904), .Z(n1977) );
  XNOR U1949 ( .A(n1978), .B(n1912), .Z(n1904) );
  XNOR U1950 ( .A(n1900), .B(n1899), .Z(n1912) );
  XOR U1951 ( .A(n1979), .B(n1896), .Z(n1899) );
  XNOR U1952 ( .A(n806), .B(p_input[138]), .Z(n1896) );
  IV U1953 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n806) );
  XOR U1954 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n1013), 
        .Z(n1979) );
  XNOR U1955 ( .A(n707), .B(p_input[140]), .Z(n1900) );
  IV U1956 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n707) );
  XNOR U1957 ( .A(n1910), .B(n1901), .Z(n1978) );
  XOR U1958 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(
        p_input[129]), .Z(n1901) );
  XOR U1959 ( .A(n1980), .B(n1917), .Z(n1910) );
  XOR U1960 ( .A(n558), .B(p_input[143]), .Z(n1917) );
  IV U1961 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .Z(n558) );
  XOR U1962 ( .A(n1907), .B(n1916), .Z(n1980) );
  XOR U1963 ( .A(n1981), .B(n1913), .Z(n1916) );
  XNOR U1964 ( .A(n658), .B(p_input[141]), .Z(n1913) );
  IV U1965 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n658) );
  XNOR U1966 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(
        p_input[142]), .Z(n1981) );
  IV U1967 ( .A(n1911), .Z(n1907) );
  XOR U1968 ( .A(n92), .B(p_input[137]), .Z(n1911) );
  IV U1969 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .Z(n92) );
  XNOR U1970 ( .A(n1925), .B(n1923), .Z(n1905) );
  XOR U1971 ( .A(n1982), .B(n1930), .Z(n1923) );
  XOR U1972 ( .A(n145), .B(p_input[136]), .Z(n1930) );
  IV U1973 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .Z(n145) );
  XNOR U1974 ( .A(n1920), .B(n1929), .Z(n1982) );
  XNOR U1975 ( .A(n1983), .B(n1926), .Z(n1929) );
  XOR U1976 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .B(
        p_input[134]), .Z(n1926) );
  XNOR U1977 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(
        p_input[135]), .Z(n1983) );
  IV U1978 ( .A(n1924), .Z(n1920) );
  XOR U1979 ( .A(n453), .B(p_input[130]), .Z(n1924) );
  IV U1980 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n453) );
  XOR U1981 ( .A(n1935), .B(n1934), .Z(n1925) );
  XNOR U1982 ( .A(n1984), .B(n1931), .Z(n1934) );
  XOR U1983 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .B(
        p_input[131]), .Z(n1931) );
  XNOR U1984 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(
        p_input[132]), .Z(n1984) );
  XOR U1985 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(
        p_input[133]), .Z(n1935) );
  XOR U1986 ( .A(n1985), .B(n1965), .Z(n1823) );
  XOR U1987 ( .A(n1943), .B(n1942), .Z(n1965) );
  XNOR U1988 ( .A(n1986), .B(n1948), .Z(n1942) );
  XNOR U1989 ( .A(n149), .B(p_input[136]), .Z(n1948) );
  IV U1990 ( .A(\knn_comb_/min_val_out[0][8] ), .Z(n149) );
  XOR U1991 ( .A(n1939), .B(n1947), .Z(n1986) );
  XOR U1992 ( .A(n1987), .B(n1944), .Z(n1947) );
  XNOR U1993 ( .A(n251), .B(p_input[134]), .Z(n1944) );
  IV U1994 ( .A(\knn_comb_/min_val_out[0][6] ), .Z(n251) );
  XNOR U1995 ( .A(\knn_comb_/min_val_out[0][7] ), .B(p_input[135]), .Z(n1987)
         );
  XNOR U1996 ( .A(n457), .B(p_input[130]), .Z(n1939) );
  IV U1997 ( .A(\knn_comb_/min_val_out[0][2] ), .Z(n457) );
  XNOR U1998 ( .A(n1953), .B(n1952), .Z(n1943) );
  XOR U1999 ( .A(n1988), .B(n1949), .Z(n1952) );
  XNOR U2000 ( .A(n406), .B(p_input[131]), .Z(n1949) );
  IV U2001 ( .A(\knn_comb_/min_val_out[0][3] ), .Z(n406) );
  XNOR U2002 ( .A(\knn_comb_/min_val_out[0][4] ), .B(p_input[132]), .Z(n1988)
         );
  XNOR U2003 ( .A(n302), .B(p_input[133]), .Z(n1953) );
  IV U2004 ( .A(\knn_comb_/min_val_out[0][5] ), .Z(n302) );
  XNOR U2005 ( .A(n1964), .B(n1954), .Z(n1985) );
  XOR U2006 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[128]), .Z(n1954)
         );
  XNOR U2007 ( .A(n1989), .B(n1971), .Z(n1964) );
  XNOR U2008 ( .A(n1960), .B(n1959), .Z(n1971) );
  XOR U2009 ( .A(n1990), .B(n1956), .Z(n1959) );
  XOR U2010 ( .A(\knn_comb_/min_val_out[0][10] ), .B(p_input[138]), .Z(n1956)
         );
  XOR U2011 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n1013), .Z(n1990) );
  IV U2012 ( .A(p_input[139]), .Z(n1013) );
  XOR U2013 ( .A(\knn_comb_/min_val_out[0][12] ), .B(p_input[140]), .Z(n1960)
         );
  XNOR U2014 ( .A(n1970), .B(n1961), .Z(n1989) );
  XNOR U2015 ( .A(n508), .B(p_input[129]), .Z(n1961) );
  IV U2016 ( .A(\knn_comb_/min_val_out[0][1] ), .Z(n508) );
  XOR U2017 ( .A(n1991), .B(n1976), .Z(n1970) );
  XNOR U2018 ( .A(\knn_comb_/min_val_out[0][15] ), .B(p_input[143]), .Z(n1976)
         );
  XOR U2019 ( .A(n1967), .B(n1975), .Z(n1991) );
  XOR U2020 ( .A(n1992), .B(n1972), .Z(n1975) );
  XOR U2021 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[141]), .Z(n1972)
         );
  XNOR U2022 ( .A(\knn_comb_/min_val_out[0][14] ), .B(p_input[142]), .Z(n1992)
         );
  XNOR U2023 ( .A(n98), .B(p_input[137]), .Z(n1967) );
  IV U2024 ( .A(\knn_comb_/min_val_out[0][9] ), .Z(n98) );
endmodule

