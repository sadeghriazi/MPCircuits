
module knn_comb_BMR_W16_K2_N16 ( p_input, o );
  input [271:0] p_input;
  output [31:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][15] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369;
  assign \knn_comb_/min_val_out[0][0]  = p_input[240];
  assign \knn_comb_/min_val_out[0][1]  = p_input[241];
  assign \knn_comb_/min_val_out[0][2]  = p_input[242];
  assign \knn_comb_/min_val_out[0][3]  = p_input[243];
  assign \knn_comb_/min_val_out[0][4]  = p_input[244];
  assign \knn_comb_/min_val_out[0][5]  = p_input[245];
  assign \knn_comb_/min_val_out[0][6]  = p_input[246];
  assign \knn_comb_/min_val_out[0][7]  = p_input[247];
  assign \knn_comb_/min_val_out[0][8]  = p_input[248];
  assign \knn_comb_/min_val_out[0][9]  = p_input[249];
  assign \knn_comb_/min_val_out[0][10]  = p_input[250];
  assign \knn_comb_/min_val_out[0][11]  = p_input[251];
  assign \knn_comb_/min_val_out[0][12]  = p_input[252];
  assign \knn_comb_/min_val_out[0][13]  = p_input[253];
  assign \knn_comb_/min_val_out[0][14]  = p_input[254];
  assign \knn_comb_/min_val_out[0][15]  = p_input[255];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][0]  = p_input[224];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][1]  = p_input[225];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][2]  = p_input[226];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][3]  = p_input[227];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][4]  = p_input[228];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][5]  = p_input[229];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][6]  = p_input[230];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][7]  = p_input[231];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][8]  = p_input[232];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][9]  = p_input[233];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][10]  = p_input[234];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][11]  = p_input[235];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][12]  = p_input[236];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][13]  = p_input[237];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][14]  = p_input[238];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][15]  = p_input[239];

  XOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  XOR U2 ( .A(n3), .B(n4), .Z(o[8]) );
  XOR U3 ( .A(n5), .B(n6), .Z(o[7]) );
  XOR U4 ( .A(n7), .B(n8), .Z(o[6]) );
  XOR U5 ( .A(n9), .B(n10), .Z(o[5]) );
  XOR U6 ( .A(n11), .B(n12), .Z(o[4]) );
  XOR U7 ( .A(n13), .B(n14), .Z(o[3]) );
  XOR U8 ( .A(n15), .B(n16), .Z(o[31]) );
  XOR U9 ( .A(n17), .B(n18), .Z(o[30]) );
  XOR U10 ( .A(n19), .B(n20), .Z(o[2]) );
  XOR U11 ( .A(n21), .B(n22), .Z(o[29]) );
  XOR U12 ( .A(n23), .B(n24), .Z(o[28]) );
  XOR U13 ( .A(n25), .B(n26), .Z(o[27]) );
  XOR U14 ( .A(n27), .B(n28), .Z(o[26]) );
  XOR U15 ( .A(n1), .B(n29), .Z(o[25]) );
  AND U16 ( .A(n30), .B(n31), .Z(n1) );
  XOR U17 ( .A(n2), .B(n29), .Z(n31) );
  XOR U18 ( .A(n32), .B(n33), .Z(n29) );
  AND U19 ( .A(n34), .B(n35), .Z(n33) );
  XOR U20 ( .A(p_input[9]), .B(n32), .Z(n35) );
  XOR U21 ( .A(n36), .B(n37), .Z(n32) );
  AND U22 ( .A(n38), .B(n39), .Z(n37) );
  XOR U23 ( .A(n40), .B(n41), .Z(n2) );
  AND U24 ( .A(n42), .B(n39), .Z(n41) );
  XNOR U25 ( .A(n43), .B(n36), .Z(n39) );
  XOR U26 ( .A(n44), .B(n45), .Z(n36) );
  AND U27 ( .A(n46), .B(n47), .Z(n45) );
  XOR U28 ( .A(p_input[25]), .B(n44), .Z(n47) );
  XOR U29 ( .A(n48), .B(n49), .Z(n44) );
  AND U30 ( .A(n50), .B(n51), .Z(n49) );
  IV U31 ( .A(n40), .Z(n43) );
  XNOR U32 ( .A(n52), .B(n53), .Z(n40) );
  AND U33 ( .A(n54), .B(n51), .Z(n53) );
  XNOR U34 ( .A(n52), .B(n48), .Z(n51) );
  XOR U35 ( .A(n55), .B(n56), .Z(n48) );
  AND U36 ( .A(n57), .B(n58), .Z(n56) );
  XOR U37 ( .A(p_input[41]), .B(n55), .Z(n58) );
  XOR U38 ( .A(n59), .B(n60), .Z(n55) );
  AND U39 ( .A(n61), .B(n62), .Z(n60) );
  XOR U40 ( .A(n63), .B(n64), .Z(n52) );
  AND U41 ( .A(n65), .B(n62), .Z(n64) );
  XNOR U42 ( .A(n63), .B(n59), .Z(n62) );
  XOR U43 ( .A(n66), .B(n67), .Z(n59) );
  AND U44 ( .A(n68), .B(n69), .Z(n67) );
  XOR U45 ( .A(p_input[57]), .B(n66), .Z(n69) );
  XOR U46 ( .A(n70), .B(n71), .Z(n66) );
  AND U47 ( .A(n72), .B(n73), .Z(n71) );
  XOR U48 ( .A(n74), .B(n75), .Z(n63) );
  AND U49 ( .A(n76), .B(n73), .Z(n75) );
  XNOR U50 ( .A(n74), .B(n70), .Z(n73) );
  XOR U51 ( .A(n77), .B(n78), .Z(n70) );
  AND U52 ( .A(n79), .B(n80), .Z(n78) );
  XOR U53 ( .A(p_input[73]), .B(n77), .Z(n80) );
  XOR U54 ( .A(n81), .B(n82), .Z(n77) );
  AND U55 ( .A(n83), .B(n84), .Z(n82) );
  XOR U56 ( .A(n85), .B(n86), .Z(n74) );
  AND U57 ( .A(n87), .B(n84), .Z(n86) );
  XNOR U58 ( .A(n85), .B(n81), .Z(n84) );
  XOR U59 ( .A(n88), .B(n89), .Z(n81) );
  AND U60 ( .A(n90), .B(n91), .Z(n89) );
  XOR U61 ( .A(p_input[89]), .B(n88), .Z(n91) );
  XOR U62 ( .A(n92), .B(n93), .Z(n88) );
  AND U63 ( .A(n94), .B(n95), .Z(n93) );
  XOR U64 ( .A(n96), .B(n97), .Z(n85) );
  AND U65 ( .A(n98), .B(n95), .Z(n97) );
  XNOR U66 ( .A(n96), .B(n92), .Z(n95) );
  XOR U67 ( .A(n99), .B(n100), .Z(n92) );
  AND U68 ( .A(n101), .B(n102), .Z(n100) );
  XOR U69 ( .A(p_input[105]), .B(n99), .Z(n102) );
  XOR U70 ( .A(n103), .B(n104), .Z(n99) );
  AND U71 ( .A(n105), .B(n106), .Z(n104) );
  XOR U72 ( .A(n107), .B(n108), .Z(n96) );
  AND U73 ( .A(n109), .B(n106), .Z(n108) );
  XNOR U74 ( .A(n107), .B(n103), .Z(n106) );
  XOR U75 ( .A(n110), .B(n111), .Z(n103) );
  AND U76 ( .A(n112), .B(n113), .Z(n111) );
  XOR U77 ( .A(p_input[121]), .B(n110), .Z(n113) );
  XOR U78 ( .A(n114), .B(n115), .Z(n110) );
  AND U79 ( .A(n116), .B(n117), .Z(n115) );
  XOR U80 ( .A(n118), .B(n119), .Z(n107) );
  AND U81 ( .A(n120), .B(n117), .Z(n119) );
  XNOR U82 ( .A(n118), .B(n114), .Z(n117) );
  XOR U83 ( .A(n121), .B(n122), .Z(n114) );
  AND U84 ( .A(n123), .B(n124), .Z(n122) );
  XOR U85 ( .A(p_input[137]), .B(n121), .Z(n124) );
  XOR U86 ( .A(n125), .B(n126), .Z(n121) );
  AND U87 ( .A(n127), .B(n128), .Z(n126) );
  XOR U88 ( .A(n129), .B(n130), .Z(n118) );
  AND U89 ( .A(n131), .B(n128), .Z(n130) );
  XNOR U90 ( .A(n129), .B(n125), .Z(n128) );
  XOR U91 ( .A(n132), .B(n133), .Z(n125) );
  AND U92 ( .A(n134), .B(n135), .Z(n133) );
  XOR U93 ( .A(p_input[153]), .B(n132), .Z(n135) );
  XOR U94 ( .A(n136), .B(n137), .Z(n132) );
  AND U95 ( .A(n138), .B(n139), .Z(n137) );
  XOR U96 ( .A(n140), .B(n141), .Z(n129) );
  AND U97 ( .A(n142), .B(n139), .Z(n141) );
  XNOR U98 ( .A(n140), .B(n136), .Z(n139) );
  XOR U99 ( .A(n143), .B(n144), .Z(n136) );
  AND U100 ( .A(n145), .B(n146), .Z(n144) );
  XOR U101 ( .A(p_input[169]), .B(n143), .Z(n146) );
  XOR U102 ( .A(n147), .B(n148), .Z(n143) );
  AND U103 ( .A(n149), .B(n150), .Z(n148) );
  XOR U104 ( .A(n151), .B(n152), .Z(n140) );
  AND U105 ( .A(n153), .B(n150), .Z(n152) );
  XNOR U106 ( .A(n151), .B(n147), .Z(n150) );
  XOR U107 ( .A(n154), .B(n155), .Z(n147) );
  AND U108 ( .A(n156), .B(n157), .Z(n155) );
  XOR U109 ( .A(p_input[185]), .B(n154), .Z(n157) );
  XOR U110 ( .A(n158), .B(n159), .Z(n154) );
  AND U111 ( .A(n160), .B(n161), .Z(n159) );
  XOR U112 ( .A(n162), .B(n163), .Z(n151) );
  AND U113 ( .A(n164), .B(n161), .Z(n163) );
  XNOR U114 ( .A(n162), .B(n158), .Z(n161) );
  XOR U115 ( .A(n165), .B(n166), .Z(n158) );
  AND U116 ( .A(n167), .B(n168), .Z(n166) );
  XOR U117 ( .A(p_input[201]), .B(n165), .Z(n168) );
  XOR U118 ( .A(n169), .B(n170), .Z(n165) );
  AND U119 ( .A(n171), .B(n172), .Z(n170) );
  XOR U120 ( .A(n173), .B(n174), .Z(n162) );
  AND U121 ( .A(n175), .B(n172), .Z(n174) );
  XNOR U122 ( .A(n173), .B(n169), .Z(n172) );
  XOR U123 ( .A(n176), .B(n177), .Z(n169) );
  AND U124 ( .A(n178), .B(n179), .Z(n177) );
  XOR U125 ( .A(p_input[217]), .B(n176), .Z(n179) );
  XNOR U126 ( .A(n180), .B(n181), .Z(n176) );
  AND U127 ( .A(n182), .B(n183), .Z(n181) );
  XNOR U128 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n184), .Z(n173) );
  AND U129 ( .A(n185), .B(n183), .Z(n184) );
  XOR U130 ( .A(n186), .B(n180), .Z(n183) );
  XOR U131 ( .A(n3), .B(n187), .Z(o[24]) );
  AND U132 ( .A(n30), .B(n188), .Z(n3) );
  XOR U133 ( .A(n4), .B(n187), .Z(n188) );
  XOR U134 ( .A(n189), .B(n190), .Z(n187) );
  AND U135 ( .A(n34), .B(n191), .Z(n190) );
  XOR U136 ( .A(p_input[8]), .B(n189), .Z(n191) );
  XOR U137 ( .A(n192), .B(n193), .Z(n189) );
  AND U138 ( .A(n38), .B(n194), .Z(n193) );
  XOR U139 ( .A(n195), .B(n196), .Z(n4) );
  AND U140 ( .A(n42), .B(n194), .Z(n196) );
  XNOR U141 ( .A(n197), .B(n192), .Z(n194) );
  XOR U142 ( .A(n198), .B(n199), .Z(n192) );
  AND U143 ( .A(n46), .B(n200), .Z(n199) );
  XOR U144 ( .A(p_input[24]), .B(n198), .Z(n200) );
  XOR U145 ( .A(n201), .B(n202), .Z(n198) );
  AND U146 ( .A(n50), .B(n203), .Z(n202) );
  IV U147 ( .A(n195), .Z(n197) );
  XNOR U148 ( .A(n204), .B(n205), .Z(n195) );
  AND U149 ( .A(n54), .B(n203), .Z(n205) );
  XNOR U150 ( .A(n204), .B(n201), .Z(n203) );
  XOR U151 ( .A(n206), .B(n207), .Z(n201) );
  AND U152 ( .A(n57), .B(n208), .Z(n207) );
  XOR U153 ( .A(p_input[40]), .B(n206), .Z(n208) );
  XOR U154 ( .A(n209), .B(n210), .Z(n206) );
  AND U155 ( .A(n61), .B(n211), .Z(n210) );
  XOR U156 ( .A(n212), .B(n213), .Z(n204) );
  AND U157 ( .A(n65), .B(n211), .Z(n213) );
  XNOR U158 ( .A(n212), .B(n209), .Z(n211) );
  XOR U159 ( .A(n214), .B(n215), .Z(n209) );
  AND U160 ( .A(n68), .B(n216), .Z(n215) );
  XOR U161 ( .A(p_input[56]), .B(n214), .Z(n216) );
  XOR U162 ( .A(n217), .B(n218), .Z(n214) );
  AND U163 ( .A(n72), .B(n219), .Z(n218) );
  XOR U164 ( .A(n220), .B(n221), .Z(n212) );
  AND U165 ( .A(n76), .B(n219), .Z(n221) );
  XNOR U166 ( .A(n220), .B(n217), .Z(n219) );
  XOR U167 ( .A(n222), .B(n223), .Z(n217) );
  AND U168 ( .A(n79), .B(n224), .Z(n223) );
  XOR U169 ( .A(p_input[72]), .B(n222), .Z(n224) );
  XOR U170 ( .A(n225), .B(n226), .Z(n222) );
  AND U171 ( .A(n83), .B(n227), .Z(n226) );
  XOR U172 ( .A(n228), .B(n229), .Z(n220) );
  AND U173 ( .A(n87), .B(n227), .Z(n229) );
  XNOR U174 ( .A(n228), .B(n225), .Z(n227) );
  XOR U175 ( .A(n230), .B(n231), .Z(n225) );
  AND U176 ( .A(n90), .B(n232), .Z(n231) );
  XOR U177 ( .A(p_input[88]), .B(n230), .Z(n232) );
  XOR U178 ( .A(n233), .B(n234), .Z(n230) );
  AND U179 ( .A(n94), .B(n235), .Z(n234) );
  XOR U180 ( .A(n236), .B(n237), .Z(n228) );
  AND U181 ( .A(n98), .B(n235), .Z(n237) );
  XNOR U182 ( .A(n236), .B(n233), .Z(n235) );
  XOR U183 ( .A(n238), .B(n239), .Z(n233) );
  AND U184 ( .A(n101), .B(n240), .Z(n239) );
  XOR U185 ( .A(p_input[104]), .B(n238), .Z(n240) );
  XOR U186 ( .A(n241), .B(n242), .Z(n238) );
  AND U187 ( .A(n105), .B(n243), .Z(n242) );
  XOR U188 ( .A(n244), .B(n245), .Z(n236) );
  AND U189 ( .A(n109), .B(n243), .Z(n245) );
  XNOR U190 ( .A(n244), .B(n241), .Z(n243) );
  XOR U191 ( .A(n246), .B(n247), .Z(n241) );
  AND U192 ( .A(n112), .B(n248), .Z(n247) );
  XOR U193 ( .A(p_input[120]), .B(n246), .Z(n248) );
  XOR U194 ( .A(n249), .B(n250), .Z(n246) );
  AND U195 ( .A(n116), .B(n251), .Z(n250) );
  XOR U196 ( .A(n252), .B(n253), .Z(n244) );
  AND U197 ( .A(n120), .B(n251), .Z(n253) );
  XNOR U198 ( .A(n252), .B(n249), .Z(n251) );
  XOR U199 ( .A(n254), .B(n255), .Z(n249) );
  AND U200 ( .A(n123), .B(n256), .Z(n255) );
  XOR U201 ( .A(p_input[136]), .B(n254), .Z(n256) );
  XOR U202 ( .A(n257), .B(n258), .Z(n254) );
  AND U203 ( .A(n127), .B(n259), .Z(n258) );
  XOR U204 ( .A(n260), .B(n261), .Z(n252) );
  AND U205 ( .A(n131), .B(n259), .Z(n261) );
  XNOR U206 ( .A(n260), .B(n257), .Z(n259) );
  XOR U207 ( .A(n262), .B(n263), .Z(n257) );
  AND U208 ( .A(n134), .B(n264), .Z(n263) );
  XOR U209 ( .A(p_input[152]), .B(n262), .Z(n264) );
  XOR U210 ( .A(n265), .B(n266), .Z(n262) );
  AND U211 ( .A(n138), .B(n267), .Z(n266) );
  XOR U212 ( .A(n268), .B(n269), .Z(n260) );
  AND U213 ( .A(n142), .B(n267), .Z(n269) );
  XNOR U214 ( .A(n268), .B(n265), .Z(n267) );
  XOR U215 ( .A(n270), .B(n271), .Z(n265) );
  AND U216 ( .A(n145), .B(n272), .Z(n271) );
  XOR U217 ( .A(p_input[168]), .B(n270), .Z(n272) );
  XOR U218 ( .A(n273), .B(n274), .Z(n270) );
  AND U219 ( .A(n149), .B(n275), .Z(n274) );
  XOR U220 ( .A(n276), .B(n277), .Z(n268) );
  AND U221 ( .A(n153), .B(n275), .Z(n277) );
  XNOR U222 ( .A(n276), .B(n273), .Z(n275) );
  XOR U223 ( .A(n278), .B(n279), .Z(n273) );
  AND U224 ( .A(n156), .B(n280), .Z(n279) );
  XOR U225 ( .A(p_input[184]), .B(n278), .Z(n280) );
  XOR U226 ( .A(n281), .B(n282), .Z(n278) );
  AND U227 ( .A(n160), .B(n283), .Z(n282) );
  XOR U228 ( .A(n284), .B(n285), .Z(n276) );
  AND U229 ( .A(n164), .B(n283), .Z(n285) );
  XNOR U230 ( .A(n284), .B(n281), .Z(n283) );
  XOR U231 ( .A(n286), .B(n287), .Z(n281) );
  AND U232 ( .A(n167), .B(n288), .Z(n287) );
  XOR U233 ( .A(p_input[200]), .B(n286), .Z(n288) );
  XOR U234 ( .A(n289), .B(n290), .Z(n286) );
  AND U235 ( .A(n171), .B(n291), .Z(n290) );
  XOR U236 ( .A(n292), .B(n293), .Z(n284) );
  AND U237 ( .A(n175), .B(n291), .Z(n293) );
  XNOR U238 ( .A(n292), .B(n289), .Z(n291) );
  XOR U239 ( .A(n294), .B(n295), .Z(n289) );
  AND U240 ( .A(n178), .B(n296), .Z(n295) );
  XOR U241 ( .A(p_input[216]), .B(n294), .Z(n296) );
  XNOR U242 ( .A(n297), .B(n298), .Z(n294) );
  AND U243 ( .A(n182), .B(n299), .Z(n298) );
  XNOR U244 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n300), .Z(n292) );
  AND U245 ( .A(n185), .B(n299), .Z(n300) );
  XOR U246 ( .A(n301), .B(n297), .Z(n299) );
  XOR U247 ( .A(n5), .B(n302), .Z(o[23]) );
  AND U248 ( .A(n30), .B(n303), .Z(n5) );
  XOR U249 ( .A(n6), .B(n302), .Z(n303) );
  XOR U250 ( .A(n304), .B(n305), .Z(n302) );
  AND U251 ( .A(n34), .B(n306), .Z(n305) );
  XOR U252 ( .A(p_input[7]), .B(n304), .Z(n306) );
  XOR U253 ( .A(n307), .B(n308), .Z(n304) );
  AND U254 ( .A(n38), .B(n309), .Z(n308) );
  XOR U255 ( .A(n310), .B(n311), .Z(n6) );
  AND U256 ( .A(n42), .B(n309), .Z(n311) );
  XNOR U257 ( .A(n312), .B(n307), .Z(n309) );
  XOR U258 ( .A(n313), .B(n314), .Z(n307) );
  AND U259 ( .A(n46), .B(n315), .Z(n314) );
  XOR U260 ( .A(p_input[23]), .B(n313), .Z(n315) );
  XOR U261 ( .A(n316), .B(n317), .Z(n313) );
  AND U262 ( .A(n50), .B(n318), .Z(n317) );
  IV U263 ( .A(n310), .Z(n312) );
  XNOR U264 ( .A(n319), .B(n320), .Z(n310) );
  AND U265 ( .A(n54), .B(n318), .Z(n320) );
  XNOR U266 ( .A(n319), .B(n316), .Z(n318) );
  XOR U267 ( .A(n321), .B(n322), .Z(n316) );
  AND U268 ( .A(n57), .B(n323), .Z(n322) );
  XOR U269 ( .A(p_input[39]), .B(n321), .Z(n323) );
  XOR U270 ( .A(n324), .B(n325), .Z(n321) );
  AND U271 ( .A(n61), .B(n326), .Z(n325) );
  XOR U272 ( .A(n327), .B(n328), .Z(n319) );
  AND U273 ( .A(n65), .B(n326), .Z(n328) );
  XNOR U274 ( .A(n327), .B(n324), .Z(n326) );
  XOR U275 ( .A(n329), .B(n330), .Z(n324) );
  AND U276 ( .A(n68), .B(n331), .Z(n330) );
  XOR U277 ( .A(p_input[55]), .B(n329), .Z(n331) );
  XOR U278 ( .A(n332), .B(n333), .Z(n329) );
  AND U279 ( .A(n72), .B(n334), .Z(n333) );
  XOR U280 ( .A(n335), .B(n336), .Z(n327) );
  AND U281 ( .A(n76), .B(n334), .Z(n336) );
  XNOR U282 ( .A(n335), .B(n332), .Z(n334) );
  XOR U283 ( .A(n337), .B(n338), .Z(n332) );
  AND U284 ( .A(n79), .B(n339), .Z(n338) );
  XOR U285 ( .A(p_input[71]), .B(n337), .Z(n339) );
  XOR U286 ( .A(n340), .B(n341), .Z(n337) );
  AND U287 ( .A(n83), .B(n342), .Z(n341) );
  XOR U288 ( .A(n343), .B(n344), .Z(n335) );
  AND U289 ( .A(n87), .B(n342), .Z(n344) );
  XNOR U290 ( .A(n343), .B(n340), .Z(n342) );
  XOR U291 ( .A(n345), .B(n346), .Z(n340) );
  AND U292 ( .A(n90), .B(n347), .Z(n346) );
  XOR U293 ( .A(p_input[87]), .B(n345), .Z(n347) );
  XOR U294 ( .A(n348), .B(n349), .Z(n345) );
  AND U295 ( .A(n94), .B(n350), .Z(n349) );
  XOR U296 ( .A(n351), .B(n352), .Z(n343) );
  AND U297 ( .A(n98), .B(n350), .Z(n352) );
  XNOR U298 ( .A(n351), .B(n348), .Z(n350) );
  XOR U299 ( .A(n353), .B(n354), .Z(n348) );
  AND U300 ( .A(n101), .B(n355), .Z(n354) );
  XOR U301 ( .A(p_input[103]), .B(n353), .Z(n355) );
  XOR U302 ( .A(n356), .B(n357), .Z(n353) );
  AND U303 ( .A(n105), .B(n358), .Z(n357) );
  XOR U304 ( .A(n359), .B(n360), .Z(n351) );
  AND U305 ( .A(n109), .B(n358), .Z(n360) );
  XNOR U306 ( .A(n359), .B(n356), .Z(n358) );
  XOR U307 ( .A(n361), .B(n362), .Z(n356) );
  AND U308 ( .A(n112), .B(n363), .Z(n362) );
  XOR U309 ( .A(p_input[119]), .B(n361), .Z(n363) );
  XOR U310 ( .A(n364), .B(n365), .Z(n361) );
  AND U311 ( .A(n116), .B(n366), .Z(n365) );
  XOR U312 ( .A(n367), .B(n368), .Z(n359) );
  AND U313 ( .A(n120), .B(n366), .Z(n368) );
  XNOR U314 ( .A(n367), .B(n364), .Z(n366) );
  XOR U315 ( .A(n369), .B(n370), .Z(n364) );
  AND U316 ( .A(n123), .B(n371), .Z(n370) );
  XOR U317 ( .A(p_input[135]), .B(n369), .Z(n371) );
  XOR U318 ( .A(n372), .B(n373), .Z(n369) );
  AND U319 ( .A(n127), .B(n374), .Z(n373) );
  XOR U320 ( .A(n375), .B(n376), .Z(n367) );
  AND U321 ( .A(n131), .B(n374), .Z(n376) );
  XNOR U322 ( .A(n375), .B(n372), .Z(n374) );
  XOR U323 ( .A(n377), .B(n378), .Z(n372) );
  AND U324 ( .A(n134), .B(n379), .Z(n378) );
  XOR U325 ( .A(p_input[151]), .B(n377), .Z(n379) );
  XOR U326 ( .A(n380), .B(n381), .Z(n377) );
  AND U327 ( .A(n138), .B(n382), .Z(n381) );
  XOR U328 ( .A(n383), .B(n384), .Z(n375) );
  AND U329 ( .A(n142), .B(n382), .Z(n384) );
  XNOR U330 ( .A(n383), .B(n380), .Z(n382) );
  XOR U331 ( .A(n385), .B(n386), .Z(n380) );
  AND U332 ( .A(n145), .B(n387), .Z(n386) );
  XOR U333 ( .A(p_input[167]), .B(n385), .Z(n387) );
  XOR U334 ( .A(n388), .B(n389), .Z(n385) );
  AND U335 ( .A(n149), .B(n390), .Z(n389) );
  XOR U336 ( .A(n391), .B(n392), .Z(n383) );
  AND U337 ( .A(n153), .B(n390), .Z(n392) );
  XNOR U338 ( .A(n391), .B(n388), .Z(n390) );
  XOR U339 ( .A(n393), .B(n394), .Z(n388) );
  AND U340 ( .A(n156), .B(n395), .Z(n394) );
  XOR U341 ( .A(p_input[183]), .B(n393), .Z(n395) );
  XOR U342 ( .A(n396), .B(n397), .Z(n393) );
  AND U343 ( .A(n160), .B(n398), .Z(n397) );
  XOR U344 ( .A(n399), .B(n400), .Z(n391) );
  AND U345 ( .A(n164), .B(n398), .Z(n400) );
  XNOR U346 ( .A(n399), .B(n396), .Z(n398) );
  XOR U347 ( .A(n401), .B(n402), .Z(n396) );
  AND U348 ( .A(n167), .B(n403), .Z(n402) );
  XOR U349 ( .A(p_input[199]), .B(n401), .Z(n403) );
  XOR U350 ( .A(n404), .B(n405), .Z(n401) );
  AND U351 ( .A(n171), .B(n406), .Z(n405) );
  XOR U352 ( .A(n407), .B(n408), .Z(n399) );
  AND U353 ( .A(n175), .B(n406), .Z(n408) );
  XNOR U354 ( .A(n407), .B(n404), .Z(n406) );
  XOR U355 ( .A(n409), .B(n410), .Z(n404) );
  AND U356 ( .A(n178), .B(n411), .Z(n410) );
  XOR U357 ( .A(p_input[215]), .B(n409), .Z(n411) );
  XNOR U358 ( .A(n412), .B(n413), .Z(n409) );
  AND U359 ( .A(n182), .B(n414), .Z(n413) );
  XNOR U360 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n415), .Z(n407) );
  AND U361 ( .A(n185), .B(n414), .Z(n415) );
  XOR U362 ( .A(n416), .B(n412), .Z(n414) );
  IV U363 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .Z(n412) );
  IV U364 ( .A(\knn_comb_/min_val_out[0][7] ), .Z(n416) );
  XOR U365 ( .A(n7), .B(n417), .Z(o[22]) );
  AND U366 ( .A(n30), .B(n418), .Z(n7) );
  XOR U367 ( .A(n8), .B(n417), .Z(n418) );
  XOR U368 ( .A(n419), .B(n420), .Z(n417) );
  AND U369 ( .A(n34), .B(n421), .Z(n420) );
  XOR U370 ( .A(p_input[6]), .B(n419), .Z(n421) );
  XOR U371 ( .A(n422), .B(n423), .Z(n419) );
  AND U372 ( .A(n38), .B(n424), .Z(n423) );
  XOR U373 ( .A(n425), .B(n426), .Z(n8) );
  AND U374 ( .A(n42), .B(n424), .Z(n426) );
  XNOR U375 ( .A(n427), .B(n422), .Z(n424) );
  XOR U376 ( .A(n428), .B(n429), .Z(n422) );
  AND U377 ( .A(n46), .B(n430), .Z(n429) );
  XOR U378 ( .A(p_input[22]), .B(n428), .Z(n430) );
  XOR U379 ( .A(n431), .B(n432), .Z(n428) );
  AND U380 ( .A(n50), .B(n433), .Z(n432) );
  IV U381 ( .A(n425), .Z(n427) );
  XNOR U382 ( .A(n434), .B(n435), .Z(n425) );
  AND U383 ( .A(n54), .B(n433), .Z(n435) );
  XNOR U384 ( .A(n434), .B(n431), .Z(n433) );
  XOR U385 ( .A(n436), .B(n437), .Z(n431) );
  AND U386 ( .A(n57), .B(n438), .Z(n437) );
  XOR U387 ( .A(p_input[38]), .B(n436), .Z(n438) );
  XOR U388 ( .A(n439), .B(n440), .Z(n436) );
  AND U389 ( .A(n61), .B(n441), .Z(n440) );
  XOR U390 ( .A(n442), .B(n443), .Z(n434) );
  AND U391 ( .A(n65), .B(n441), .Z(n443) );
  XNOR U392 ( .A(n442), .B(n439), .Z(n441) );
  XOR U393 ( .A(n444), .B(n445), .Z(n439) );
  AND U394 ( .A(n68), .B(n446), .Z(n445) );
  XOR U395 ( .A(p_input[54]), .B(n444), .Z(n446) );
  XOR U396 ( .A(n447), .B(n448), .Z(n444) );
  AND U397 ( .A(n72), .B(n449), .Z(n448) );
  XOR U398 ( .A(n450), .B(n451), .Z(n442) );
  AND U399 ( .A(n76), .B(n449), .Z(n451) );
  XNOR U400 ( .A(n450), .B(n447), .Z(n449) );
  XOR U401 ( .A(n452), .B(n453), .Z(n447) );
  AND U402 ( .A(n79), .B(n454), .Z(n453) );
  XOR U403 ( .A(p_input[70]), .B(n452), .Z(n454) );
  XOR U404 ( .A(n455), .B(n456), .Z(n452) );
  AND U405 ( .A(n83), .B(n457), .Z(n456) );
  XOR U406 ( .A(n458), .B(n459), .Z(n450) );
  AND U407 ( .A(n87), .B(n457), .Z(n459) );
  XNOR U408 ( .A(n458), .B(n455), .Z(n457) );
  XOR U409 ( .A(n460), .B(n461), .Z(n455) );
  AND U410 ( .A(n90), .B(n462), .Z(n461) );
  XOR U411 ( .A(p_input[86]), .B(n460), .Z(n462) );
  XOR U412 ( .A(n463), .B(n464), .Z(n460) );
  AND U413 ( .A(n94), .B(n465), .Z(n464) );
  XOR U414 ( .A(n466), .B(n467), .Z(n458) );
  AND U415 ( .A(n98), .B(n465), .Z(n467) );
  XNOR U416 ( .A(n466), .B(n463), .Z(n465) );
  XOR U417 ( .A(n468), .B(n469), .Z(n463) );
  AND U418 ( .A(n101), .B(n470), .Z(n469) );
  XOR U419 ( .A(p_input[102]), .B(n468), .Z(n470) );
  XOR U420 ( .A(n471), .B(n472), .Z(n468) );
  AND U421 ( .A(n105), .B(n473), .Z(n472) );
  XOR U422 ( .A(n474), .B(n475), .Z(n466) );
  AND U423 ( .A(n109), .B(n473), .Z(n475) );
  XNOR U424 ( .A(n474), .B(n471), .Z(n473) );
  XOR U425 ( .A(n476), .B(n477), .Z(n471) );
  AND U426 ( .A(n112), .B(n478), .Z(n477) );
  XOR U427 ( .A(p_input[118]), .B(n476), .Z(n478) );
  XOR U428 ( .A(n479), .B(n480), .Z(n476) );
  AND U429 ( .A(n116), .B(n481), .Z(n480) );
  XOR U430 ( .A(n482), .B(n483), .Z(n474) );
  AND U431 ( .A(n120), .B(n481), .Z(n483) );
  XNOR U432 ( .A(n482), .B(n479), .Z(n481) );
  XOR U433 ( .A(n484), .B(n485), .Z(n479) );
  AND U434 ( .A(n123), .B(n486), .Z(n485) );
  XOR U435 ( .A(p_input[134]), .B(n484), .Z(n486) );
  XOR U436 ( .A(n487), .B(n488), .Z(n484) );
  AND U437 ( .A(n127), .B(n489), .Z(n488) );
  XOR U438 ( .A(n490), .B(n491), .Z(n482) );
  AND U439 ( .A(n131), .B(n489), .Z(n491) );
  XNOR U440 ( .A(n490), .B(n487), .Z(n489) );
  XOR U441 ( .A(n492), .B(n493), .Z(n487) );
  AND U442 ( .A(n134), .B(n494), .Z(n493) );
  XOR U443 ( .A(p_input[150]), .B(n492), .Z(n494) );
  XOR U444 ( .A(n495), .B(n496), .Z(n492) );
  AND U445 ( .A(n138), .B(n497), .Z(n496) );
  XOR U446 ( .A(n498), .B(n499), .Z(n490) );
  AND U447 ( .A(n142), .B(n497), .Z(n499) );
  XNOR U448 ( .A(n498), .B(n495), .Z(n497) );
  XOR U449 ( .A(n500), .B(n501), .Z(n495) );
  AND U450 ( .A(n145), .B(n502), .Z(n501) );
  XOR U451 ( .A(p_input[166]), .B(n500), .Z(n502) );
  XOR U452 ( .A(n503), .B(n504), .Z(n500) );
  AND U453 ( .A(n149), .B(n505), .Z(n504) );
  XOR U454 ( .A(n506), .B(n507), .Z(n498) );
  AND U455 ( .A(n153), .B(n505), .Z(n507) );
  XNOR U456 ( .A(n506), .B(n503), .Z(n505) );
  XOR U457 ( .A(n508), .B(n509), .Z(n503) );
  AND U458 ( .A(n156), .B(n510), .Z(n509) );
  XOR U459 ( .A(p_input[182]), .B(n508), .Z(n510) );
  XOR U460 ( .A(n511), .B(n512), .Z(n508) );
  AND U461 ( .A(n160), .B(n513), .Z(n512) );
  XOR U462 ( .A(n514), .B(n515), .Z(n506) );
  AND U463 ( .A(n164), .B(n513), .Z(n515) );
  XNOR U464 ( .A(n514), .B(n511), .Z(n513) );
  XOR U465 ( .A(n516), .B(n517), .Z(n511) );
  AND U466 ( .A(n167), .B(n518), .Z(n517) );
  XOR U467 ( .A(p_input[198]), .B(n516), .Z(n518) );
  XOR U468 ( .A(n519), .B(n520), .Z(n516) );
  AND U469 ( .A(n171), .B(n521), .Z(n520) );
  XOR U470 ( .A(n522), .B(n523), .Z(n514) );
  AND U471 ( .A(n175), .B(n521), .Z(n523) );
  XNOR U472 ( .A(n522), .B(n519), .Z(n521) );
  XOR U473 ( .A(n524), .B(n525), .Z(n519) );
  AND U474 ( .A(n178), .B(n526), .Z(n525) );
  XOR U475 ( .A(p_input[214]), .B(n524), .Z(n526) );
  XNOR U476 ( .A(n527), .B(n528), .Z(n524) );
  AND U477 ( .A(n182), .B(n529), .Z(n528) );
  XNOR U478 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n530), .Z(n522) );
  AND U479 ( .A(n185), .B(n529), .Z(n530) );
  XOR U480 ( .A(n531), .B(n527), .Z(n529) );
  XOR U481 ( .A(n9), .B(n532), .Z(o[21]) );
  AND U482 ( .A(n30), .B(n533), .Z(n9) );
  XOR U483 ( .A(n10), .B(n532), .Z(n533) );
  XOR U484 ( .A(n534), .B(n535), .Z(n532) );
  AND U485 ( .A(n34), .B(n536), .Z(n535) );
  XOR U486 ( .A(p_input[5]), .B(n534), .Z(n536) );
  XOR U487 ( .A(n537), .B(n538), .Z(n534) );
  AND U488 ( .A(n38), .B(n539), .Z(n538) );
  XOR U489 ( .A(n540), .B(n541), .Z(n10) );
  AND U490 ( .A(n42), .B(n539), .Z(n541) );
  XNOR U491 ( .A(n542), .B(n537), .Z(n539) );
  XOR U492 ( .A(n543), .B(n544), .Z(n537) );
  AND U493 ( .A(n46), .B(n545), .Z(n544) );
  XOR U494 ( .A(p_input[21]), .B(n543), .Z(n545) );
  XOR U495 ( .A(n546), .B(n547), .Z(n543) );
  AND U496 ( .A(n50), .B(n548), .Z(n547) );
  IV U497 ( .A(n540), .Z(n542) );
  XNOR U498 ( .A(n549), .B(n550), .Z(n540) );
  AND U499 ( .A(n54), .B(n548), .Z(n550) );
  XNOR U500 ( .A(n549), .B(n546), .Z(n548) );
  XOR U501 ( .A(n551), .B(n552), .Z(n546) );
  AND U502 ( .A(n57), .B(n553), .Z(n552) );
  XOR U503 ( .A(p_input[37]), .B(n551), .Z(n553) );
  XOR U504 ( .A(n554), .B(n555), .Z(n551) );
  AND U505 ( .A(n61), .B(n556), .Z(n555) );
  XOR U506 ( .A(n557), .B(n558), .Z(n549) );
  AND U507 ( .A(n65), .B(n556), .Z(n558) );
  XNOR U508 ( .A(n557), .B(n554), .Z(n556) );
  XOR U509 ( .A(n559), .B(n560), .Z(n554) );
  AND U510 ( .A(n68), .B(n561), .Z(n560) );
  XOR U511 ( .A(p_input[53]), .B(n559), .Z(n561) );
  XOR U512 ( .A(n562), .B(n563), .Z(n559) );
  AND U513 ( .A(n72), .B(n564), .Z(n563) );
  XOR U514 ( .A(n565), .B(n566), .Z(n557) );
  AND U515 ( .A(n76), .B(n564), .Z(n566) );
  XNOR U516 ( .A(n565), .B(n562), .Z(n564) );
  XOR U517 ( .A(n567), .B(n568), .Z(n562) );
  AND U518 ( .A(n79), .B(n569), .Z(n568) );
  XOR U519 ( .A(p_input[69]), .B(n567), .Z(n569) );
  XOR U520 ( .A(n570), .B(n571), .Z(n567) );
  AND U521 ( .A(n83), .B(n572), .Z(n571) );
  XOR U522 ( .A(n573), .B(n574), .Z(n565) );
  AND U523 ( .A(n87), .B(n572), .Z(n574) );
  XNOR U524 ( .A(n573), .B(n570), .Z(n572) );
  XOR U525 ( .A(n575), .B(n576), .Z(n570) );
  AND U526 ( .A(n90), .B(n577), .Z(n576) );
  XOR U527 ( .A(p_input[85]), .B(n575), .Z(n577) );
  XOR U528 ( .A(n578), .B(n579), .Z(n575) );
  AND U529 ( .A(n94), .B(n580), .Z(n579) );
  XOR U530 ( .A(n581), .B(n582), .Z(n573) );
  AND U531 ( .A(n98), .B(n580), .Z(n582) );
  XNOR U532 ( .A(n581), .B(n578), .Z(n580) );
  XOR U533 ( .A(n583), .B(n584), .Z(n578) );
  AND U534 ( .A(n101), .B(n585), .Z(n584) );
  XOR U535 ( .A(p_input[101]), .B(n583), .Z(n585) );
  XOR U536 ( .A(n586), .B(n587), .Z(n583) );
  AND U537 ( .A(n105), .B(n588), .Z(n587) );
  XOR U538 ( .A(n589), .B(n590), .Z(n581) );
  AND U539 ( .A(n109), .B(n588), .Z(n590) );
  XNOR U540 ( .A(n589), .B(n586), .Z(n588) );
  XOR U541 ( .A(n591), .B(n592), .Z(n586) );
  AND U542 ( .A(n112), .B(n593), .Z(n592) );
  XOR U543 ( .A(p_input[117]), .B(n591), .Z(n593) );
  XOR U544 ( .A(n594), .B(n595), .Z(n591) );
  AND U545 ( .A(n116), .B(n596), .Z(n595) );
  XOR U546 ( .A(n597), .B(n598), .Z(n589) );
  AND U547 ( .A(n120), .B(n596), .Z(n598) );
  XNOR U548 ( .A(n597), .B(n594), .Z(n596) );
  XOR U549 ( .A(n599), .B(n600), .Z(n594) );
  AND U550 ( .A(n123), .B(n601), .Z(n600) );
  XOR U551 ( .A(p_input[133]), .B(n599), .Z(n601) );
  XOR U552 ( .A(n602), .B(n603), .Z(n599) );
  AND U553 ( .A(n127), .B(n604), .Z(n603) );
  XOR U554 ( .A(n605), .B(n606), .Z(n597) );
  AND U555 ( .A(n131), .B(n604), .Z(n606) );
  XNOR U556 ( .A(n605), .B(n602), .Z(n604) );
  XOR U557 ( .A(n607), .B(n608), .Z(n602) );
  AND U558 ( .A(n134), .B(n609), .Z(n608) );
  XOR U559 ( .A(p_input[149]), .B(n607), .Z(n609) );
  XOR U560 ( .A(n610), .B(n611), .Z(n607) );
  AND U561 ( .A(n138), .B(n612), .Z(n611) );
  XOR U562 ( .A(n613), .B(n614), .Z(n605) );
  AND U563 ( .A(n142), .B(n612), .Z(n614) );
  XNOR U564 ( .A(n613), .B(n610), .Z(n612) );
  XOR U565 ( .A(n615), .B(n616), .Z(n610) );
  AND U566 ( .A(n145), .B(n617), .Z(n616) );
  XOR U567 ( .A(p_input[165]), .B(n615), .Z(n617) );
  XOR U568 ( .A(n618), .B(n619), .Z(n615) );
  AND U569 ( .A(n149), .B(n620), .Z(n619) );
  XOR U570 ( .A(n621), .B(n622), .Z(n613) );
  AND U571 ( .A(n153), .B(n620), .Z(n622) );
  XNOR U572 ( .A(n621), .B(n618), .Z(n620) );
  XOR U573 ( .A(n623), .B(n624), .Z(n618) );
  AND U574 ( .A(n156), .B(n625), .Z(n624) );
  XOR U575 ( .A(p_input[181]), .B(n623), .Z(n625) );
  XOR U576 ( .A(n626), .B(n627), .Z(n623) );
  AND U577 ( .A(n160), .B(n628), .Z(n627) );
  XOR U578 ( .A(n629), .B(n630), .Z(n621) );
  AND U579 ( .A(n164), .B(n628), .Z(n630) );
  XNOR U580 ( .A(n629), .B(n626), .Z(n628) );
  XOR U581 ( .A(n631), .B(n632), .Z(n626) );
  AND U582 ( .A(n167), .B(n633), .Z(n632) );
  XOR U583 ( .A(p_input[197]), .B(n631), .Z(n633) );
  XOR U584 ( .A(n634), .B(n635), .Z(n631) );
  AND U585 ( .A(n171), .B(n636), .Z(n635) );
  XOR U586 ( .A(n637), .B(n638), .Z(n629) );
  AND U587 ( .A(n175), .B(n636), .Z(n638) );
  XNOR U588 ( .A(n637), .B(n634), .Z(n636) );
  XOR U589 ( .A(n639), .B(n640), .Z(n634) );
  AND U590 ( .A(n178), .B(n641), .Z(n640) );
  XOR U591 ( .A(p_input[213]), .B(n639), .Z(n641) );
  XNOR U592 ( .A(n642), .B(n643), .Z(n639) );
  AND U593 ( .A(n182), .B(n644), .Z(n643) );
  XNOR U594 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n645), .Z(n637) );
  AND U595 ( .A(n185), .B(n644), .Z(n645) );
  XOR U596 ( .A(n646), .B(n642), .Z(n644) );
  XOR U597 ( .A(n11), .B(n647), .Z(o[20]) );
  AND U598 ( .A(n30), .B(n648), .Z(n11) );
  XOR U599 ( .A(n12), .B(n647), .Z(n648) );
  XOR U600 ( .A(n649), .B(n650), .Z(n647) );
  AND U601 ( .A(n34), .B(n651), .Z(n650) );
  XOR U602 ( .A(p_input[4]), .B(n649), .Z(n651) );
  XOR U603 ( .A(n652), .B(n653), .Z(n649) );
  AND U604 ( .A(n38), .B(n654), .Z(n653) );
  XOR U605 ( .A(n655), .B(n656), .Z(n12) );
  AND U606 ( .A(n42), .B(n654), .Z(n656) );
  XNOR U607 ( .A(n657), .B(n652), .Z(n654) );
  XOR U608 ( .A(n658), .B(n659), .Z(n652) );
  AND U609 ( .A(n46), .B(n660), .Z(n659) );
  XOR U610 ( .A(p_input[20]), .B(n658), .Z(n660) );
  XOR U611 ( .A(n661), .B(n662), .Z(n658) );
  AND U612 ( .A(n50), .B(n663), .Z(n662) );
  IV U613 ( .A(n655), .Z(n657) );
  XNOR U614 ( .A(n664), .B(n665), .Z(n655) );
  AND U615 ( .A(n54), .B(n663), .Z(n665) );
  XNOR U616 ( .A(n664), .B(n661), .Z(n663) );
  XOR U617 ( .A(n666), .B(n667), .Z(n661) );
  AND U618 ( .A(n57), .B(n668), .Z(n667) );
  XOR U619 ( .A(p_input[36]), .B(n666), .Z(n668) );
  XOR U620 ( .A(n669), .B(n670), .Z(n666) );
  AND U621 ( .A(n61), .B(n671), .Z(n670) );
  XOR U622 ( .A(n672), .B(n673), .Z(n664) );
  AND U623 ( .A(n65), .B(n671), .Z(n673) );
  XNOR U624 ( .A(n672), .B(n669), .Z(n671) );
  XOR U625 ( .A(n674), .B(n675), .Z(n669) );
  AND U626 ( .A(n68), .B(n676), .Z(n675) );
  XOR U627 ( .A(p_input[52]), .B(n674), .Z(n676) );
  XOR U628 ( .A(n677), .B(n678), .Z(n674) );
  AND U629 ( .A(n72), .B(n679), .Z(n678) );
  XOR U630 ( .A(n680), .B(n681), .Z(n672) );
  AND U631 ( .A(n76), .B(n679), .Z(n681) );
  XNOR U632 ( .A(n680), .B(n677), .Z(n679) );
  XOR U633 ( .A(n682), .B(n683), .Z(n677) );
  AND U634 ( .A(n79), .B(n684), .Z(n683) );
  XOR U635 ( .A(p_input[68]), .B(n682), .Z(n684) );
  XOR U636 ( .A(n685), .B(n686), .Z(n682) );
  AND U637 ( .A(n83), .B(n687), .Z(n686) );
  XOR U638 ( .A(n688), .B(n689), .Z(n680) );
  AND U639 ( .A(n87), .B(n687), .Z(n689) );
  XNOR U640 ( .A(n688), .B(n685), .Z(n687) );
  XOR U641 ( .A(n690), .B(n691), .Z(n685) );
  AND U642 ( .A(n90), .B(n692), .Z(n691) );
  XOR U643 ( .A(p_input[84]), .B(n690), .Z(n692) );
  XOR U644 ( .A(n693), .B(n694), .Z(n690) );
  AND U645 ( .A(n94), .B(n695), .Z(n694) );
  XOR U646 ( .A(n696), .B(n697), .Z(n688) );
  AND U647 ( .A(n98), .B(n695), .Z(n697) );
  XNOR U648 ( .A(n696), .B(n693), .Z(n695) );
  XOR U649 ( .A(n698), .B(n699), .Z(n693) );
  AND U650 ( .A(n101), .B(n700), .Z(n699) );
  XOR U651 ( .A(p_input[100]), .B(n698), .Z(n700) );
  XOR U652 ( .A(n701), .B(n702), .Z(n698) );
  AND U653 ( .A(n105), .B(n703), .Z(n702) );
  XOR U654 ( .A(n704), .B(n705), .Z(n696) );
  AND U655 ( .A(n109), .B(n703), .Z(n705) );
  XNOR U656 ( .A(n704), .B(n701), .Z(n703) );
  XOR U657 ( .A(n706), .B(n707), .Z(n701) );
  AND U658 ( .A(n112), .B(n708), .Z(n707) );
  XOR U659 ( .A(p_input[116]), .B(n706), .Z(n708) );
  XOR U660 ( .A(n709), .B(n710), .Z(n706) );
  AND U661 ( .A(n116), .B(n711), .Z(n710) );
  XOR U662 ( .A(n712), .B(n713), .Z(n704) );
  AND U663 ( .A(n120), .B(n711), .Z(n713) );
  XNOR U664 ( .A(n712), .B(n709), .Z(n711) );
  XOR U665 ( .A(n714), .B(n715), .Z(n709) );
  AND U666 ( .A(n123), .B(n716), .Z(n715) );
  XOR U667 ( .A(p_input[132]), .B(n714), .Z(n716) );
  XOR U668 ( .A(n717), .B(n718), .Z(n714) );
  AND U669 ( .A(n127), .B(n719), .Z(n718) );
  XOR U670 ( .A(n720), .B(n721), .Z(n712) );
  AND U671 ( .A(n131), .B(n719), .Z(n721) );
  XNOR U672 ( .A(n720), .B(n717), .Z(n719) );
  XOR U673 ( .A(n722), .B(n723), .Z(n717) );
  AND U674 ( .A(n134), .B(n724), .Z(n723) );
  XOR U675 ( .A(p_input[148]), .B(n722), .Z(n724) );
  XOR U676 ( .A(n725), .B(n726), .Z(n722) );
  AND U677 ( .A(n138), .B(n727), .Z(n726) );
  XOR U678 ( .A(n728), .B(n729), .Z(n720) );
  AND U679 ( .A(n142), .B(n727), .Z(n729) );
  XNOR U680 ( .A(n728), .B(n725), .Z(n727) );
  XOR U681 ( .A(n730), .B(n731), .Z(n725) );
  AND U682 ( .A(n145), .B(n732), .Z(n731) );
  XOR U683 ( .A(p_input[164]), .B(n730), .Z(n732) );
  XOR U684 ( .A(n733), .B(n734), .Z(n730) );
  AND U685 ( .A(n149), .B(n735), .Z(n734) );
  XOR U686 ( .A(n736), .B(n737), .Z(n728) );
  AND U687 ( .A(n153), .B(n735), .Z(n737) );
  XNOR U688 ( .A(n736), .B(n733), .Z(n735) );
  XOR U689 ( .A(n738), .B(n739), .Z(n733) );
  AND U690 ( .A(n156), .B(n740), .Z(n739) );
  XOR U691 ( .A(p_input[180]), .B(n738), .Z(n740) );
  XOR U692 ( .A(n741), .B(n742), .Z(n738) );
  AND U693 ( .A(n160), .B(n743), .Z(n742) );
  XOR U694 ( .A(n744), .B(n745), .Z(n736) );
  AND U695 ( .A(n164), .B(n743), .Z(n745) );
  XNOR U696 ( .A(n744), .B(n741), .Z(n743) );
  XOR U697 ( .A(n746), .B(n747), .Z(n741) );
  AND U698 ( .A(n167), .B(n748), .Z(n747) );
  XOR U699 ( .A(p_input[196]), .B(n746), .Z(n748) );
  XOR U700 ( .A(n749), .B(n750), .Z(n746) );
  AND U701 ( .A(n171), .B(n751), .Z(n750) );
  XOR U702 ( .A(n752), .B(n753), .Z(n744) );
  AND U703 ( .A(n175), .B(n751), .Z(n753) );
  XNOR U704 ( .A(n752), .B(n749), .Z(n751) );
  XOR U705 ( .A(n754), .B(n755), .Z(n749) );
  AND U706 ( .A(n178), .B(n756), .Z(n755) );
  XOR U707 ( .A(p_input[212]), .B(n754), .Z(n756) );
  XNOR U708 ( .A(n757), .B(n758), .Z(n754) );
  AND U709 ( .A(n182), .B(n759), .Z(n758) );
  XNOR U710 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n760), .Z(n752) );
  AND U711 ( .A(n185), .B(n759), .Z(n760) );
  XOR U712 ( .A(n761), .B(n757), .Z(n759) );
  IV U713 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .Z(n757) );
  IV U714 ( .A(\knn_comb_/min_val_out[0][4] ), .Z(n761) );
  XOR U715 ( .A(n762), .B(n763), .Z(o[1]) );
  XOR U716 ( .A(n13), .B(n764), .Z(o[19]) );
  AND U717 ( .A(n30), .B(n765), .Z(n13) );
  XOR U718 ( .A(n14), .B(n764), .Z(n765) );
  XOR U719 ( .A(n766), .B(n767), .Z(n764) );
  AND U720 ( .A(n34), .B(n768), .Z(n767) );
  XOR U721 ( .A(p_input[3]), .B(n766), .Z(n768) );
  XOR U722 ( .A(n769), .B(n770), .Z(n766) );
  AND U723 ( .A(n38), .B(n771), .Z(n770) );
  XOR U724 ( .A(n772), .B(n773), .Z(n14) );
  AND U725 ( .A(n42), .B(n771), .Z(n773) );
  XNOR U726 ( .A(n774), .B(n769), .Z(n771) );
  XOR U727 ( .A(n775), .B(n776), .Z(n769) );
  AND U728 ( .A(n46), .B(n777), .Z(n776) );
  XOR U729 ( .A(p_input[19]), .B(n775), .Z(n777) );
  XOR U730 ( .A(n778), .B(n779), .Z(n775) );
  AND U731 ( .A(n50), .B(n780), .Z(n779) );
  IV U732 ( .A(n772), .Z(n774) );
  XNOR U733 ( .A(n781), .B(n782), .Z(n772) );
  AND U734 ( .A(n54), .B(n780), .Z(n782) );
  XNOR U735 ( .A(n781), .B(n778), .Z(n780) );
  XOR U736 ( .A(n783), .B(n784), .Z(n778) );
  AND U737 ( .A(n57), .B(n785), .Z(n784) );
  XOR U738 ( .A(p_input[35]), .B(n783), .Z(n785) );
  XOR U739 ( .A(n786), .B(n787), .Z(n783) );
  AND U740 ( .A(n61), .B(n788), .Z(n787) );
  XOR U741 ( .A(n789), .B(n790), .Z(n781) );
  AND U742 ( .A(n65), .B(n788), .Z(n790) );
  XNOR U743 ( .A(n789), .B(n786), .Z(n788) );
  XOR U744 ( .A(n791), .B(n792), .Z(n786) );
  AND U745 ( .A(n68), .B(n793), .Z(n792) );
  XOR U746 ( .A(p_input[51]), .B(n791), .Z(n793) );
  XOR U747 ( .A(n794), .B(n795), .Z(n791) );
  AND U748 ( .A(n72), .B(n796), .Z(n795) );
  XOR U749 ( .A(n797), .B(n798), .Z(n789) );
  AND U750 ( .A(n76), .B(n796), .Z(n798) );
  XNOR U751 ( .A(n797), .B(n794), .Z(n796) );
  XOR U752 ( .A(n799), .B(n800), .Z(n794) );
  AND U753 ( .A(n79), .B(n801), .Z(n800) );
  XOR U754 ( .A(p_input[67]), .B(n799), .Z(n801) );
  XOR U755 ( .A(n802), .B(n803), .Z(n799) );
  AND U756 ( .A(n83), .B(n804), .Z(n803) );
  XOR U757 ( .A(n805), .B(n806), .Z(n797) );
  AND U758 ( .A(n87), .B(n804), .Z(n806) );
  XNOR U759 ( .A(n805), .B(n802), .Z(n804) );
  XOR U760 ( .A(n807), .B(n808), .Z(n802) );
  AND U761 ( .A(n90), .B(n809), .Z(n808) );
  XOR U762 ( .A(p_input[83]), .B(n807), .Z(n809) );
  XOR U763 ( .A(n810), .B(n811), .Z(n807) );
  AND U764 ( .A(n94), .B(n812), .Z(n811) );
  XOR U765 ( .A(n813), .B(n814), .Z(n805) );
  AND U766 ( .A(n98), .B(n812), .Z(n814) );
  XNOR U767 ( .A(n813), .B(n810), .Z(n812) );
  XOR U768 ( .A(n815), .B(n816), .Z(n810) );
  AND U769 ( .A(n101), .B(n817), .Z(n816) );
  XOR U770 ( .A(p_input[99]), .B(n815), .Z(n817) );
  XOR U771 ( .A(n818), .B(n819), .Z(n815) );
  AND U772 ( .A(n105), .B(n820), .Z(n819) );
  XOR U773 ( .A(n821), .B(n822), .Z(n813) );
  AND U774 ( .A(n109), .B(n820), .Z(n822) );
  XNOR U775 ( .A(n821), .B(n818), .Z(n820) );
  XOR U776 ( .A(n823), .B(n824), .Z(n818) );
  AND U777 ( .A(n112), .B(n825), .Z(n824) );
  XOR U778 ( .A(p_input[115]), .B(n823), .Z(n825) );
  XOR U779 ( .A(n826), .B(n827), .Z(n823) );
  AND U780 ( .A(n116), .B(n828), .Z(n827) );
  XOR U781 ( .A(n829), .B(n830), .Z(n821) );
  AND U782 ( .A(n120), .B(n828), .Z(n830) );
  XNOR U783 ( .A(n829), .B(n826), .Z(n828) );
  XOR U784 ( .A(n831), .B(n832), .Z(n826) );
  AND U785 ( .A(n123), .B(n833), .Z(n832) );
  XOR U786 ( .A(p_input[131]), .B(n831), .Z(n833) );
  XOR U787 ( .A(n834), .B(n835), .Z(n831) );
  AND U788 ( .A(n127), .B(n836), .Z(n835) );
  XOR U789 ( .A(n837), .B(n838), .Z(n829) );
  AND U790 ( .A(n131), .B(n836), .Z(n838) );
  XNOR U791 ( .A(n837), .B(n834), .Z(n836) );
  XOR U792 ( .A(n839), .B(n840), .Z(n834) );
  AND U793 ( .A(n134), .B(n841), .Z(n840) );
  XOR U794 ( .A(p_input[147]), .B(n839), .Z(n841) );
  XOR U795 ( .A(n842), .B(n843), .Z(n839) );
  AND U796 ( .A(n138), .B(n844), .Z(n843) );
  XOR U797 ( .A(n845), .B(n846), .Z(n837) );
  AND U798 ( .A(n142), .B(n844), .Z(n846) );
  XNOR U799 ( .A(n845), .B(n842), .Z(n844) );
  XOR U800 ( .A(n847), .B(n848), .Z(n842) );
  AND U801 ( .A(n145), .B(n849), .Z(n848) );
  XOR U802 ( .A(p_input[163]), .B(n847), .Z(n849) );
  XOR U803 ( .A(n850), .B(n851), .Z(n847) );
  AND U804 ( .A(n149), .B(n852), .Z(n851) );
  XOR U805 ( .A(n853), .B(n854), .Z(n845) );
  AND U806 ( .A(n153), .B(n852), .Z(n854) );
  XNOR U807 ( .A(n853), .B(n850), .Z(n852) );
  XOR U808 ( .A(n855), .B(n856), .Z(n850) );
  AND U809 ( .A(n156), .B(n857), .Z(n856) );
  XOR U810 ( .A(p_input[179]), .B(n855), .Z(n857) );
  XOR U811 ( .A(n858), .B(n859), .Z(n855) );
  AND U812 ( .A(n160), .B(n860), .Z(n859) );
  XOR U813 ( .A(n861), .B(n862), .Z(n853) );
  AND U814 ( .A(n164), .B(n860), .Z(n862) );
  XNOR U815 ( .A(n861), .B(n858), .Z(n860) );
  XOR U816 ( .A(n863), .B(n864), .Z(n858) );
  AND U817 ( .A(n167), .B(n865), .Z(n864) );
  XOR U818 ( .A(p_input[195]), .B(n863), .Z(n865) );
  XOR U819 ( .A(n866), .B(n867), .Z(n863) );
  AND U820 ( .A(n171), .B(n868), .Z(n867) );
  XOR U821 ( .A(n869), .B(n870), .Z(n861) );
  AND U822 ( .A(n175), .B(n868), .Z(n870) );
  XNOR U823 ( .A(n869), .B(n866), .Z(n868) );
  XOR U824 ( .A(n871), .B(n872), .Z(n866) );
  AND U825 ( .A(n178), .B(n873), .Z(n872) );
  XOR U826 ( .A(p_input[211]), .B(n871), .Z(n873) );
  XNOR U827 ( .A(n874), .B(n875), .Z(n871) );
  AND U828 ( .A(n182), .B(n876), .Z(n875) );
  XNOR U829 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n877), .Z(n869) );
  AND U830 ( .A(n185), .B(n876), .Z(n877) );
  XOR U831 ( .A(n878), .B(n874), .Z(n876) );
  XOR U832 ( .A(n19), .B(n879), .Z(o[18]) );
  AND U833 ( .A(n30), .B(n880), .Z(n19) );
  XOR U834 ( .A(n20), .B(n879), .Z(n880) );
  XOR U835 ( .A(n881), .B(n882), .Z(n879) );
  AND U836 ( .A(n34), .B(n883), .Z(n882) );
  XOR U837 ( .A(p_input[2]), .B(n881), .Z(n883) );
  XOR U838 ( .A(n884), .B(n885), .Z(n881) );
  AND U839 ( .A(n38), .B(n886), .Z(n885) );
  XOR U840 ( .A(n887), .B(n888), .Z(n20) );
  AND U841 ( .A(n42), .B(n886), .Z(n888) );
  XNOR U842 ( .A(n889), .B(n884), .Z(n886) );
  XOR U843 ( .A(n890), .B(n891), .Z(n884) );
  AND U844 ( .A(n46), .B(n892), .Z(n891) );
  XOR U845 ( .A(p_input[18]), .B(n890), .Z(n892) );
  XOR U846 ( .A(n893), .B(n894), .Z(n890) );
  AND U847 ( .A(n50), .B(n895), .Z(n894) );
  IV U848 ( .A(n887), .Z(n889) );
  XNOR U849 ( .A(n896), .B(n897), .Z(n887) );
  AND U850 ( .A(n54), .B(n895), .Z(n897) );
  XNOR U851 ( .A(n896), .B(n893), .Z(n895) );
  XOR U852 ( .A(n898), .B(n899), .Z(n893) );
  AND U853 ( .A(n57), .B(n900), .Z(n899) );
  XOR U854 ( .A(p_input[34]), .B(n898), .Z(n900) );
  XOR U855 ( .A(n901), .B(n902), .Z(n898) );
  AND U856 ( .A(n61), .B(n903), .Z(n902) );
  XOR U857 ( .A(n904), .B(n905), .Z(n896) );
  AND U858 ( .A(n65), .B(n903), .Z(n905) );
  XNOR U859 ( .A(n904), .B(n901), .Z(n903) );
  XOR U860 ( .A(n906), .B(n907), .Z(n901) );
  AND U861 ( .A(n68), .B(n908), .Z(n907) );
  XOR U862 ( .A(p_input[50]), .B(n906), .Z(n908) );
  XOR U863 ( .A(n909), .B(n910), .Z(n906) );
  AND U864 ( .A(n72), .B(n911), .Z(n910) );
  XOR U865 ( .A(n912), .B(n913), .Z(n904) );
  AND U866 ( .A(n76), .B(n911), .Z(n913) );
  XNOR U867 ( .A(n912), .B(n909), .Z(n911) );
  XOR U868 ( .A(n914), .B(n915), .Z(n909) );
  AND U869 ( .A(n79), .B(n916), .Z(n915) );
  XOR U870 ( .A(p_input[66]), .B(n914), .Z(n916) );
  XOR U871 ( .A(n917), .B(n918), .Z(n914) );
  AND U872 ( .A(n83), .B(n919), .Z(n918) );
  XOR U873 ( .A(n920), .B(n921), .Z(n912) );
  AND U874 ( .A(n87), .B(n919), .Z(n921) );
  XNOR U875 ( .A(n920), .B(n917), .Z(n919) );
  XOR U876 ( .A(n922), .B(n923), .Z(n917) );
  AND U877 ( .A(n90), .B(n924), .Z(n923) );
  XOR U878 ( .A(p_input[82]), .B(n922), .Z(n924) );
  XOR U879 ( .A(n925), .B(n926), .Z(n922) );
  AND U880 ( .A(n94), .B(n927), .Z(n926) );
  XOR U881 ( .A(n928), .B(n929), .Z(n920) );
  AND U882 ( .A(n98), .B(n927), .Z(n929) );
  XNOR U883 ( .A(n928), .B(n925), .Z(n927) );
  XOR U884 ( .A(n930), .B(n931), .Z(n925) );
  AND U885 ( .A(n101), .B(n932), .Z(n931) );
  XOR U886 ( .A(p_input[98]), .B(n930), .Z(n932) );
  XOR U887 ( .A(n933), .B(n934), .Z(n930) );
  AND U888 ( .A(n105), .B(n935), .Z(n934) );
  XOR U889 ( .A(n936), .B(n937), .Z(n928) );
  AND U890 ( .A(n109), .B(n935), .Z(n937) );
  XNOR U891 ( .A(n936), .B(n933), .Z(n935) );
  XOR U892 ( .A(n938), .B(n939), .Z(n933) );
  AND U893 ( .A(n112), .B(n940), .Z(n939) );
  XOR U894 ( .A(p_input[114]), .B(n938), .Z(n940) );
  XOR U895 ( .A(n941), .B(n942), .Z(n938) );
  AND U896 ( .A(n116), .B(n943), .Z(n942) );
  XOR U897 ( .A(n944), .B(n945), .Z(n936) );
  AND U898 ( .A(n120), .B(n943), .Z(n945) );
  XNOR U899 ( .A(n944), .B(n941), .Z(n943) );
  XOR U900 ( .A(n946), .B(n947), .Z(n941) );
  AND U901 ( .A(n123), .B(n948), .Z(n947) );
  XOR U902 ( .A(p_input[130]), .B(n946), .Z(n948) );
  XOR U903 ( .A(n949), .B(n950), .Z(n946) );
  AND U904 ( .A(n127), .B(n951), .Z(n950) );
  XOR U905 ( .A(n952), .B(n953), .Z(n944) );
  AND U906 ( .A(n131), .B(n951), .Z(n953) );
  XNOR U907 ( .A(n952), .B(n949), .Z(n951) );
  XOR U908 ( .A(n954), .B(n955), .Z(n949) );
  AND U909 ( .A(n134), .B(n956), .Z(n955) );
  XOR U910 ( .A(p_input[146]), .B(n954), .Z(n956) );
  XOR U911 ( .A(n957), .B(n958), .Z(n954) );
  AND U912 ( .A(n138), .B(n959), .Z(n958) );
  XOR U913 ( .A(n960), .B(n961), .Z(n952) );
  AND U914 ( .A(n142), .B(n959), .Z(n961) );
  XNOR U915 ( .A(n960), .B(n957), .Z(n959) );
  XOR U916 ( .A(n962), .B(n963), .Z(n957) );
  AND U917 ( .A(n145), .B(n964), .Z(n963) );
  XOR U918 ( .A(p_input[162]), .B(n962), .Z(n964) );
  XOR U919 ( .A(n965), .B(n966), .Z(n962) );
  AND U920 ( .A(n149), .B(n967), .Z(n966) );
  XOR U921 ( .A(n968), .B(n969), .Z(n960) );
  AND U922 ( .A(n153), .B(n967), .Z(n969) );
  XNOR U923 ( .A(n968), .B(n965), .Z(n967) );
  XOR U924 ( .A(n970), .B(n971), .Z(n965) );
  AND U925 ( .A(n156), .B(n972), .Z(n971) );
  XOR U926 ( .A(p_input[178]), .B(n970), .Z(n972) );
  XOR U927 ( .A(n973), .B(n974), .Z(n970) );
  AND U928 ( .A(n160), .B(n975), .Z(n974) );
  XOR U929 ( .A(n976), .B(n977), .Z(n968) );
  AND U930 ( .A(n164), .B(n975), .Z(n977) );
  XNOR U931 ( .A(n976), .B(n973), .Z(n975) );
  XOR U932 ( .A(n978), .B(n979), .Z(n973) );
  AND U933 ( .A(n167), .B(n980), .Z(n979) );
  XOR U934 ( .A(p_input[194]), .B(n978), .Z(n980) );
  XOR U935 ( .A(n981), .B(n982), .Z(n978) );
  AND U936 ( .A(n171), .B(n983), .Z(n982) );
  XOR U937 ( .A(n984), .B(n985), .Z(n976) );
  AND U938 ( .A(n175), .B(n983), .Z(n985) );
  XNOR U939 ( .A(n984), .B(n981), .Z(n983) );
  XOR U940 ( .A(n986), .B(n987), .Z(n981) );
  AND U941 ( .A(n178), .B(n988), .Z(n987) );
  XOR U942 ( .A(p_input[210]), .B(n986), .Z(n988) );
  XNOR U943 ( .A(n989), .B(n990), .Z(n986) );
  AND U944 ( .A(n182), .B(n991), .Z(n990) );
  XNOR U945 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n992), .Z(n984) );
  AND U946 ( .A(n185), .B(n991), .Z(n992) );
  XOR U947 ( .A(n993), .B(n989), .Z(n991) );
  XOR U948 ( .A(n762), .B(n994), .Z(o[17]) );
  AND U949 ( .A(n30), .B(n995), .Z(n762) );
  XOR U950 ( .A(n763), .B(n994), .Z(n995) );
  XOR U951 ( .A(n996), .B(n997), .Z(n994) );
  AND U952 ( .A(n34), .B(n998), .Z(n997) );
  XOR U953 ( .A(p_input[1]), .B(n996), .Z(n998) );
  XOR U954 ( .A(n999), .B(n1000), .Z(n996) );
  AND U955 ( .A(n38), .B(n1001), .Z(n1000) );
  XOR U956 ( .A(n1002), .B(n1003), .Z(n763) );
  AND U957 ( .A(n42), .B(n1001), .Z(n1003) );
  XNOR U958 ( .A(n1004), .B(n999), .Z(n1001) );
  XOR U959 ( .A(n1005), .B(n1006), .Z(n999) );
  AND U960 ( .A(n46), .B(n1007), .Z(n1006) );
  XOR U961 ( .A(p_input[17]), .B(n1005), .Z(n1007) );
  XOR U962 ( .A(n1008), .B(n1009), .Z(n1005) );
  AND U963 ( .A(n50), .B(n1010), .Z(n1009) );
  IV U964 ( .A(n1002), .Z(n1004) );
  XNOR U965 ( .A(n1011), .B(n1012), .Z(n1002) );
  AND U966 ( .A(n54), .B(n1010), .Z(n1012) );
  XNOR U967 ( .A(n1011), .B(n1008), .Z(n1010) );
  XOR U968 ( .A(n1013), .B(n1014), .Z(n1008) );
  AND U969 ( .A(n57), .B(n1015), .Z(n1014) );
  XOR U970 ( .A(p_input[33]), .B(n1013), .Z(n1015) );
  XOR U971 ( .A(n1016), .B(n1017), .Z(n1013) );
  AND U972 ( .A(n61), .B(n1018), .Z(n1017) );
  XOR U973 ( .A(n1019), .B(n1020), .Z(n1011) );
  AND U974 ( .A(n65), .B(n1018), .Z(n1020) );
  XNOR U975 ( .A(n1019), .B(n1016), .Z(n1018) );
  XOR U976 ( .A(n1021), .B(n1022), .Z(n1016) );
  AND U977 ( .A(n68), .B(n1023), .Z(n1022) );
  XOR U978 ( .A(p_input[49]), .B(n1021), .Z(n1023) );
  XOR U979 ( .A(n1024), .B(n1025), .Z(n1021) );
  AND U980 ( .A(n72), .B(n1026), .Z(n1025) );
  XOR U981 ( .A(n1027), .B(n1028), .Z(n1019) );
  AND U982 ( .A(n76), .B(n1026), .Z(n1028) );
  XNOR U983 ( .A(n1027), .B(n1024), .Z(n1026) );
  XOR U984 ( .A(n1029), .B(n1030), .Z(n1024) );
  AND U985 ( .A(n79), .B(n1031), .Z(n1030) );
  XOR U986 ( .A(p_input[65]), .B(n1029), .Z(n1031) );
  XOR U987 ( .A(n1032), .B(n1033), .Z(n1029) );
  AND U988 ( .A(n83), .B(n1034), .Z(n1033) );
  XOR U989 ( .A(n1035), .B(n1036), .Z(n1027) );
  AND U990 ( .A(n87), .B(n1034), .Z(n1036) );
  XNOR U991 ( .A(n1035), .B(n1032), .Z(n1034) );
  XOR U992 ( .A(n1037), .B(n1038), .Z(n1032) );
  AND U993 ( .A(n90), .B(n1039), .Z(n1038) );
  XOR U994 ( .A(p_input[81]), .B(n1037), .Z(n1039) );
  XOR U995 ( .A(n1040), .B(n1041), .Z(n1037) );
  AND U996 ( .A(n94), .B(n1042), .Z(n1041) );
  XOR U997 ( .A(n1043), .B(n1044), .Z(n1035) );
  AND U998 ( .A(n98), .B(n1042), .Z(n1044) );
  XNOR U999 ( .A(n1043), .B(n1040), .Z(n1042) );
  XOR U1000 ( .A(n1045), .B(n1046), .Z(n1040) );
  AND U1001 ( .A(n101), .B(n1047), .Z(n1046) );
  XOR U1002 ( .A(p_input[97]), .B(n1045), .Z(n1047) );
  XOR U1003 ( .A(n1048), .B(n1049), .Z(n1045) );
  AND U1004 ( .A(n105), .B(n1050), .Z(n1049) );
  XOR U1005 ( .A(n1051), .B(n1052), .Z(n1043) );
  AND U1006 ( .A(n109), .B(n1050), .Z(n1052) );
  XNOR U1007 ( .A(n1051), .B(n1048), .Z(n1050) );
  XOR U1008 ( .A(n1053), .B(n1054), .Z(n1048) );
  AND U1009 ( .A(n112), .B(n1055), .Z(n1054) );
  XOR U1010 ( .A(p_input[113]), .B(n1053), .Z(n1055) );
  XOR U1011 ( .A(n1056), .B(n1057), .Z(n1053) );
  AND U1012 ( .A(n116), .B(n1058), .Z(n1057) );
  XOR U1013 ( .A(n1059), .B(n1060), .Z(n1051) );
  AND U1014 ( .A(n120), .B(n1058), .Z(n1060) );
  XNOR U1015 ( .A(n1059), .B(n1056), .Z(n1058) );
  XOR U1016 ( .A(n1061), .B(n1062), .Z(n1056) );
  AND U1017 ( .A(n123), .B(n1063), .Z(n1062) );
  XOR U1018 ( .A(p_input[129]), .B(n1061), .Z(n1063) );
  XOR U1019 ( .A(n1064), .B(n1065), .Z(n1061) );
  AND U1020 ( .A(n127), .B(n1066), .Z(n1065) );
  XOR U1021 ( .A(n1067), .B(n1068), .Z(n1059) );
  AND U1022 ( .A(n131), .B(n1066), .Z(n1068) );
  XNOR U1023 ( .A(n1067), .B(n1064), .Z(n1066) );
  XOR U1024 ( .A(n1069), .B(n1070), .Z(n1064) );
  AND U1025 ( .A(n134), .B(n1071), .Z(n1070) );
  XOR U1026 ( .A(p_input[145]), .B(n1069), .Z(n1071) );
  XOR U1027 ( .A(n1072), .B(n1073), .Z(n1069) );
  AND U1028 ( .A(n138), .B(n1074), .Z(n1073) );
  XOR U1029 ( .A(n1075), .B(n1076), .Z(n1067) );
  AND U1030 ( .A(n142), .B(n1074), .Z(n1076) );
  XNOR U1031 ( .A(n1075), .B(n1072), .Z(n1074) );
  XOR U1032 ( .A(n1077), .B(n1078), .Z(n1072) );
  AND U1033 ( .A(n145), .B(n1079), .Z(n1078) );
  XOR U1034 ( .A(p_input[161]), .B(n1077), .Z(n1079) );
  XOR U1035 ( .A(n1080), .B(n1081), .Z(n1077) );
  AND U1036 ( .A(n149), .B(n1082), .Z(n1081) );
  XOR U1037 ( .A(n1083), .B(n1084), .Z(n1075) );
  AND U1038 ( .A(n153), .B(n1082), .Z(n1084) );
  XNOR U1039 ( .A(n1083), .B(n1080), .Z(n1082) );
  XOR U1040 ( .A(n1085), .B(n1086), .Z(n1080) );
  AND U1041 ( .A(n156), .B(n1087), .Z(n1086) );
  XOR U1042 ( .A(p_input[177]), .B(n1085), .Z(n1087) );
  XOR U1043 ( .A(n1088), .B(n1089), .Z(n1085) );
  AND U1044 ( .A(n160), .B(n1090), .Z(n1089) );
  XOR U1045 ( .A(n1091), .B(n1092), .Z(n1083) );
  AND U1046 ( .A(n164), .B(n1090), .Z(n1092) );
  XNOR U1047 ( .A(n1091), .B(n1088), .Z(n1090) );
  XOR U1048 ( .A(n1093), .B(n1094), .Z(n1088) );
  AND U1049 ( .A(n167), .B(n1095), .Z(n1094) );
  XOR U1050 ( .A(p_input[193]), .B(n1093), .Z(n1095) );
  XOR U1051 ( .A(n1096), .B(n1097), .Z(n1093) );
  AND U1052 ( .A(n171), .B(n1098), .Z(n1097) );
  XOR U1053 ( .A(n1099), .B(n1100), .Z(n1091) );
  AND U1054 ( .A(n175), .B(n1098), .Z(n1100) );
  XNOR U1055 ( .A(n1099), .B(n1096), .Z(n1098) );
  XOR U1056 ( .A(n1101), .B(n1102), .Z(n1096) );
  AND U1057 ( .A(n178), .B(n1103), .Z(n1102) );
  XOR U1058 ( .A(p_input[209]), .B(n1101), .Z(n1103) );
  XNOR U1059 ( .A(n1104), .B(n1105), .Z(n1101) );
  AND U1060 ( .A(n182), .B(n1106), .Z(n1105) );
  XNOR U1061 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n1107), .Z(n1099) );
  AND U1062 ( .A(n185), .B(n1106), .Z(n1107) );
  XOR U1063 ( .A(n1108), .B(n1104), .Z(n1106) );
  XOR U1064 ( .A(n1109), .B(n1110), .Z(o[16]) );
  XOR U1065 ( .A(n15), .B(n1111), .Z(o[15]) );
  AND U1066 ( .A(n30), .B(n1112), .Z(n15) );
  XOR U1067 ( .A(n16), .B(n1111), .Z(n1112) );
  XOR U1068 ( .A(n1113), .B(n1114), .Z(n1111) );
  AND U1069 ( .A(n42), .B(n1115), .Z(n1114) );
  XOR U1070 ( .A(n1116), .B(n1117), .Z(n16) );
  AND U1071 ( .A(n34), .B(n1118), .Z(n1117) );
  XOR U1072 ( .A(p_input[15]), .B(n1116), .Z(n1118) );
  XNOR U1073 ( .A(n1119), .B(n1120), .Z(n1116) );
  AND U1074 ( .A(n38), .B(n1115), .Z(n1120) );
  XNOR U1075 ( .A(n1119), .B(n1113), .Z(n1115) );
  XOR U1076 ( .A(n1121), .B(n1122), .Z(n1113) );
  AND U1077 ( .A(n54), .B(n1123), .Z(n1122) );
  XNOR U1078 ( .A(n1124), .B(n1125), .Z(n1119) );
  AND U1079 ( .A(n46), .B(n1126), .Z(n1125) );
  XOR U1080 ( .A(p_input[31]), .B(n1124), .Z(n1126) );
  XNOR U1081 ( .A(n1127), .B(n1128), .Z(n1124) );
  AND U1082 ( .A(n50), .B(n1123), .Z(n1128) );
  XNOR U1083 ( .A(n1127), .B(n1121), .Z(n1123) );
  XOR U1084 ( .A(n1129), .B(n1130), .Z(n1121) );
  AND U1085 ( .A(n65), .B(n1131), .Z(n1130) );
  XNOR U1086 ( .A(n1132), .B(n1133), .Z(n1127) );
  AND U1087 ( .A(n57), .B(n1134), .Z(n1133) );
  XOR U1088 ( .A(p_input[47]), .B(n1132), .Z(n1134) );
  XNOR U1089 ( .A(n1135), .B(n1136), .Z(n1132) );
  AND U1090 ( .A(n61), .B(n1131), .Z(n1136) );
  XNOR U1091 ( .A(n1135), .B(n1129), .Z(n1131) );
  XOR U1092 ( .A(n1137), .B(n1138), .Z(n1129) );
  AND U1093 ( .A(n76), .B(n1139), .Z(n1138) );
  XNOR U1094 ( .A(n1140), .B(n1141), .Z(n1135) );
  AND U1095 ( .A(n68), .B(n1142), .Z(n1141) );
  XOR U1096 ( .A(p_input[63]), .B(n1140), .Z(n1142) );
  XNOR U1097 ( .A(n1143), .B(n1144), .Z(n1140) );
  AND U1098 ( .A(n72), .B(n1139), .Z(n1144) );
  XNOR U1099 ( .A(n1143), .B(n1137), .Z(n1139) );
  XOR U1100 ( .A(n1145), .B(n1146), .Z(n1137) );
  AND U1101 ( .A(n87), .B(n1147), .Z(n1146) );
  XNOR U1102 ( .A(n1148), .B(n1149), .Z(n1143) );
  AND U1103 ( .A(n79), .B(n1150), .Z(n1149) );
  XOR U1104 ( .A(p_input[79]), .B(n1148), .Z(n1150) );
  XNOR U1105 ( .A(n1151), .B(n1152), .Z(n1148) );
  AND U1106 ( .A(n83), .B(n1147), .Z(n1152) );
  XNOR U1107 ( .A(n1151), .B(n1145), .Z(n1147) );
  XOR U1108 ( .A(n1153), .B(n1154), .Z(n1145) );
  AND U1109 ( .A(n98), .B(n1155), .Z(n1154) );
  XNOR U1110 ( .A(n1156), .B(n1157), .Z(n1151) );
  AND U1111 ( .A(n90), .B(n1158), .Z(n1157) );
  XOR U1112 ( .A(p_input[95]), .B(n1156), .Z(n1158) );
  XNOR U1113 ( .A(n1159), .B(n1160), .Z(n1156) );
  AND U1114 ( .A(n94), .B(n1155), .Z(n1160) );
  XNOR U1115 ( .A(n1159), .B(n1153), .Z(n1155) );
  XOR U1116 ( .A(n1161), .B(n1162), .Z(n1153) );
  AND U1117 ( .A(n109), .B(n1163), .Z(n1162) );
  XNOR U1118 ( .A(n1164), .B(n1165), .Z(n1159) );
  AND U1119 ( .A(n101), .B(n1166), .Z(n1165) );
  XOR U1120 ( .A(p_input[111]), .B(n1164), .Z(n1166) );
  XNOR U1121 ( .A(n1167), .B(n1168), .Z(n1164) );
  AND U1122 ( .A(n105), .B(n1163), .Z(n1168) );
  XNOR U1123 ( .A(n1167), .B(n1161), .Z(n1163) );
  XOR U1124 ( .A(n1169), .B(n1170), .Z(n1161) );
  AND U1125 ( .A(n120), .B(n1171), .Z(n1170) );
  XNOR U1126 ( .A(n1172), .B(n1173), .Z(n1167) );
  AND U1127 ( .A(n112), .B(n1174), .Z(n1173) );
  XOR U1128 ( .A(p_input[127]), .B(n1172), .Z(n1174) );
  XNOR U1129 ( .A(n1175), .B(n1176), .Z(n1172) );
  AND U1130 ( .A(n116), .B(n1171), .Z(n1176) );
  XNOR U1131 ( .A(n1175), .B(n1169), .Z(n1171) );
  XOR U1132 ( .A(n1177), .B(n1178), .Z(n1169) );
  AND U1133 ( .A(n131), .B(n1179), .Z(n1178) );
  XNOR U1134 ( .A(n1180), .B(n1181), .Z(n1175) );
  AND U1135 ( .A(n123), .B(n1182), .Z(n1181) );
  XOR U1136 ( .A(p_input[143]), .B(n1180), .Z(n1182) );
  XNOR U1137 ( .A(n1183), .B(n1184), .Z(n1180) );
  AND U1138 ( .A(n127), .B(n1179), .Z(n1184) );
  XNOR U1139 ( .A(n1183), .B(n1177), .Z(n1179) );
  XOR U1140 ( .A(n1185), .B(n1186), .Z(n1177) );
  AND U1141 ( .A(n142), .B(n1187), .Z(n1186) );
  XNOR U1142 ( .A(n1188), .B(n1189), .Z(n1183) );
  AND U1143 ( .A(n134), .B(n1190), .Z(n1189) );
  XOR U1144 ( .A(p_input[159]), .B(n1188), .Z(n1190) );
  XNOR U1145 ( .A(n1191), .B(n1192), .Z(n1188) );
  AND U1146 ( .A(n138), .B(n1187), .Z(n1192) );
  XNOR U1147 ( .A(n1191), .B(n1185), .Z(n1187) );
  XOR U1148 ( .A(n1193), .B(n1194), .Z(n1185) );
  AND U1149 ( .A(n153), .B(n1195), .Z(n1194) );
  XNOR U1150 ( .A(n1196), .B(n1197), .Z(n1191) );
  AND U1151 ( .A(n145), .B(n1198), .Z(n1197) );
  XOR U1152 ( .A(p_input[175]), .B(n1196), .Z(n1198) );
  XNOR U1153 ( .A(n1199), .B(n1200), .Z(n1196) );
  AND U1154 ( .A(n149), .B(n1195), .Z(n1200) );
  XNOR U1155 ( .A(n1199), .B(n1193), .Z(n1195) );
  XOR U1156 ( .A(n1201), .B(n1202), .Z(n1193) );
  AND U1157 ( .A(n164), .B(n1203), .Z(n1202) );
  XNOR U1158 ( .A(n1204), .B(n1205), .Z(n1199) );
  AND U1159 ( .A(n156), .B(n1206), .Z(n1205) );
  XOR U1160 ( .A(p_input[191]), .B(n1204), .Z(n1206) );
  XNOR U1161 ( .A(n1207), .B(n1208), .Z(n1204) );
  AND U1162 ( .A(n160), .B(n1203), .Z(n1208) );
  XNOR U1163 ( .A(n1207), .B(n1201), .Z(n1203) );
  XOR U1164 ( .A(n1209), .B(n1210), .Z(n1201) );
  AND U1165 ( .A(n175), .B(n1211), .Z(n1210) );
  XNOR U1166 ( .A(n1212), .B(n1213), .Z(n1207) );
  AND U1167 ( .A(n167), .B(n1214), .Z(n1213) );
  XOR U1168 ( .A(p_input[207]), .B(n1212), .Z(n1214) );
  XNOR U1169 ( .A(n1215), .B(n1216), .Z(n1212) );
  AND U1170 ( .A(n171), .B(n1211), .Z(n1216) );
  XNOR U1171 ( .A(n1215), .B(n1209), .Z(n1211) );
  XOR U1172 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n1217), .Z(n1209) );
  AND U1173 ( .A(n185), .B(n1218), .Z(n1217) );
  XNOR U1174 ( .A(n1219), .B(n1220), .Z(n1215) );
  AND U1175 ( .A(n178), .B(n1221), .Z(n1220) );
  XOR U1176 ( .A(p_input[223]), .B(n1219), .Z(n1221) );
  XNOR U1177 ( .A(n1222), .B(n1223), .Z(n1219) );
  AND U1178 ( .A(n182), .B(n1218), .Z(n1223) );
  XOR U1179 ( .A(n1224), .B(n1222), .Z(n1218) );
  IV U1180 ( .A(\knn_comb_/min_val_out[0][15] ), .Z(n1224) );
  IV U1181 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .Z(n1222) );
  XOR U1182 ( .A(n17), .B(n1225), .Z(o[14]) );
  AND U1183 ( .A(n30), .B(n1226), .Z(n17) );
  XOR U1184 ( .A(n18), .B(n1225), .Z(n1226) );
  XOR U1185 ( .A(n1227), .B(n1228), .Z(n1225) );
  AND U1186 ( .A(n42), .B(n1229), .Z(n1228) );
  XOR U1187 ( .A(n1230), .B(n1231), .Z(n18) );
  AND U1188 ( .A(n34), .B(n1232), .Z(n1231) );
  XOR U1189 ( .A(p_input[14]), .B(n1230), .Z(n1232) );
  XNOR U1190 ( .A(n1233), .B(n1234), .Z(n1230) );
  AND U1191 ( .A(n38), .B(n1229), .Z(n1234) );
  XNOR U1192 ( .A(n1233), .B(n1227), .Z(n1229) );
  XOR U1193 ( .A(n1235), .B(n1236), .Z(n1227) );
  AND U1194 ( .A(n54), .B(n1237), .Z(n1236) );
  XNOR U1195 ( .A(n1238), .B(n1239), .Z(n1233) );
  AND U1196 ( .A(n46), .B(n1240), .Z(n1239) );
  XOR U1197 ( .A(p_input[30]), .B(n1238), .Z(n1240) );
  XNOR U1198 ( .A(n1241), .B(n1242), .Z(n1238) );
  AND U1199 ( .A(n50), .B(n1237), .Z(n1242) );
  XNOR U1200 ( .A(n1241), .B(n1235), .Z(n1237) );
  XOR U1201 ( .A(n1243), .B(n1244), .Z(n1235) );
  AND U1202 ( .A(n65), .B(n1245), .Z(n1244) );
  XNOR U1203 ( .A(n1246), .B(n1247), .Z(n1241) );
  AND U1204 ( .A(n57), .B(n1248), .Z(n1247) );
  XOR U1205 ( .A(p_input[46]), .B(n1246), .Z(n1248) );
  XNOR U1206 ( .A(n1249), .B(n1250), .Z(n1246) );
  AND U1207 ( .A(n61), .B(n1245), .Z(n1250) );
  XNOR U1208 ( .A(n1249), .B(n1243), .Z(n1245) );
  XOR U1209 ( .A(n1251), .B(n1252), .Z(n1243) );
  AND U1210 ( .A(n76), .B(n1253), .Z(n1252) );
  XNOR U1211 ( .A(n1254), .B(n1255), .Z(n1249) );
  AND U1212 ( .A(n68), .B(n1256), .Z(n1255) );
  XOR U1213 ( .A(p_input[62]), .B(n1254), .Z(n1256) );
  XNOR U1214 ( .A(n1257), .B(n1258), .Z(n1254) );
  AND U1215 ( .A(n72), .B(n1253), .Z(n1258) );
  XNOR U1216 ( .A(n1257), .B(n1251), .Z(n1253) );
  XOR U1217 ( .A(n1259), .B(n1260), .Z(n1251) );
  AND U1218 ( .A(n87), .B(n1261), .Z(n1260) );
  XNOR U1219 ( .A(n1262), .B(n1263), .Z(n1257) );
  AND U1220 ( .A(n79), .B(n1264), .Z(n1263) );
  XOR U1221 ( .A(p_input[78]), .B(n1262), .Z(n1264) );
  XNOR U1222 ( .A(n1265), .B(n1266), .Z(n1262) );
  AND U1223 ( .A(n83), .B(n1261), .Z(n1266) );
  XNOR U1224 ( .A(n1265), .B(n1259), .Z(n1261) );
  XOR U1225 ( .A(n1267), .B(n1268), .Z(n1259) );
  AND U1226 ( .A(n98), .B(n1269), .Z(n1268) );
  XNOR U1227 ( .A(n1270), .B(n1271), .Z(n1265) );
  AND U1228 ( .A(n90), .B(n1272), .Z(n1271) );
  XOR U1229 ( .A(p_input[94]), .B(n1270), .Z(n1272) );
  XNOR U1230 ( .A(n1273), .B(n1274), .Z(n1270) );
  AND U1231 ( .A(n94), .B(n1269), .Z(n1274) );
  XNOR U1232 ( .A(n1273), .B(n1267), .Z(n1269) );
  XOR U1233 ( .A(n1275), .B(n1276), .Z(n1267) );
  AND U1234 ( .A(n109), .B(n1277), .Z(n1276) );
  XNOR U1235 ( .A(n1278), .B(n1279), .Z(n1273) );
  AND U1236 ( .A(n101), .B(n1280), .Z(n1279) );
  XOR U1237 ( .A(p_input[110]), .B(n1278), .Z(n1280) );
  XNOR U1238 ( .A(n1281), .B(n1282), .Z(n1278) );
  AND U1239 ( .A(n105), .B(n1277), .Z(n1282) );
  XNOR U1240 ( .A(n1281), .B(n1275), .Z(n1277) );
  XOR U1241 ( .A(n1283), .B(n1284), .Z(n1275) );
  AND U1242 ( .A(n120), .B(n1285), .Z(n1284) );
  XNOR U1243 ( .A(n1286), .B(n1287), .Z(n1281) );
  AND U1244 ( .A(n112), .B(n1288), .Z(n1287) );
  XOR U1245 ( .A(p_input[126]), .B(n1286), .Z(n1288) );
  XNOR U1246 ( .A(n1289), .B(n1290), .Z(n1286) );
  AND U1247 ( .A(n116), .B(n1285), .Z(n1290) );
  XNOR U1248 ( .A(n1289), .B(n1283), .Z(n1285) );
  XOR U1249 ( .A(n1291), .B(n1292), .Z(n1283) );
  AND U1250 ( .A(n131), .B(n1293), .Z(n1292) );
  XNOR U1251 ( .A(n1294), .B(n1295), .Z(n1289) );
  AND U1252 ( .A(n123), .B(n1296), .Z(n1295) );
  XOR U1253 ( .A(p_input[142]), .B(n1294), .Z(n1296) );
  XNOR U1254 ( .A(n1297), .B(n1298), .Z(n1294) );
  AND U1255 ( .A(n127), .B(n1293), .Z(n1298) );
  XNOR U1256 ( .A(n1297), .B(n1291), .Z(n1293) );
  XOR U1257 ( .A(n1299), .B(n1300), .Z(n1291) );
  AND U1258 ( .A(n142), .B(n1301), .Z(n1300) );
  XNOR U1259 ( .A(n1302), .B(n1303), .Z(n1297) );
  AND U1260 ( .A(n134), .B(n1304), .Z(n1303) );
  XOR U1261 ( .A(p_input[158]), .B(n1302), .Z(n1304) );
  XNOR U1262 ( .A(n1305), .B(n1306), .Z(n1302) );
  AND U1263 ( .A(n138), .B(n1301), .Z(n1306) );
  XNOR U1264 ( .A(n1305), .B(n1299), .Z(n1301) );
  XOR U1265 ( .A(n1307), .B(n1308), .Z(n1299) );
  AND U1266 ( .A(n153), .B(n1309), .Z(n1308) );
  XNOR U1267 ( .A(n1310), .B(n1311), .Z(n1305) );
  AND U1268 ( .A(n145), .B(n1312), .Z(n1311) );
  XOR U1269 ( .A(p_input[174]), .B(n1310), .Z(n1312) );
  XNOR U1270 ( .A(n1313), .B(n1314), .Z(n1310) );
  AND U1271 ( .A(n149), .B(n1309), .Z(n1314) );
  XNOR U1272 ( .A(n1313), .B(n1307), .Z(n1309) );
  XOR U1273 ( .A(n1315), .B(n1316), .Z(n1307) );
  AND U1274 ( .A(n164), .B(n1317), .Z(n1316) );
  XNOR U1275 ( .A(n1318), .B(n1319), .Z(n1313) );
  AND U1276 ( .A(n156), .B(n1320), .Z(n1319) );
  XOR U1277 ( .A(p_input[190]), .B(n1318), .Z(n1320) );
  XNOR U1278 ( .A(n1321), .B(n1322), .Z(n1318) );
  AND U1279 ( .A(n160), .B(n1317), .Z(n1322) );
  XNOR U1280 ( .A(n1321), .B(n1315), .Z(n1317) );
  XOR U1281 ( .A(n1323), .B(n1324), .Z(n1315) );
  AND U1282 ( .A(n175), .B(n1325), .Z(n1324) );
  XNOR U1283 ( .A(n1326), .B(n1327), .Z(n1321) );
  AND U1284 ( .A(n167), .B(n1328), .Z(n1327) );
  XOR U1285 ( .A(p_input[206]), .B(n1326), .Z(n1328) );
  XNOR U1286 ( .A(n1329), .B(n1330), .Z(n1326) );
  AND U1287 ( .A(n171), .B(n1325), .Z(n1330) );
  XNOR U1288 ( .A(n1329), .B(n1323), .Z(n1325) );
  XOR U1289 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n1331), .Z(n1323) );
  AND U1290 ( .A(n185), .B(n1332), .Z(n1331) );
  XNOR U1291 ( .A(n1333), .B(n1334), .Z(n1329) );
  AND U1292 ( .A(n178), .B(n1335), .Z(n1334) );
  XOR U1293 ( .A(p_input[222]), .B(n1333), .Z(n1335) );
  XNOR U1294 ( .A(n1336), .B(n1337), .Z(n1333) );
  AND U1295 ( .A(n182), .B(n1332), .Z(n1337) );
  XOR U1296 ( .A(n1338), .B(n1336), .Z(n1332) );
  IV U1297 ( .A(\knn_comb_/min_val_out[0][14] ), .Z(n1338) );
  IV U1298 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n1336) );
  XOR U1299 ( .A(n21), .B(n1339), .Z(o[13]) );
  AND U1300 ( .A(n30), .B(n1340), .Z(n21) );
  XOR U1301 ( .A(n22), .B(n1339), .Z(n1340) );
  XOR U1302 ( .A(n1341), .B(n1342), .Z(n1339) );
  AND U1303 ( .A(n42), .B(n1343), .Z(n1342) );
  XOR U1304 ( .A(n1344), .B(n1345), .Z(n22) );
  AND U1305 ( .A(n34), .B(n1346), .Z(n1345) );
  XOR U1306 ( .A(p_input[13]), .B(n1344), .Z(n1346) );
  XNOR U1307 ( .A(n1347), .B(n1348), .Z(n1344) );
  AND U1308 ( .A(n38), .B(n1343), .Z(n1348) );
  XNOR U1309 ( .A(n1347), .B(n1341), .Z(n1343) );
  XOR U1310 ( .A(n1349), .B(n1350), .Z(n1341) );
  AND U1311 ( .A(n54), .B(n1351), .Z(n1350) );
  XNOR U1312 ( .A(n1352), .B(n1353), .Z(n1347) );
  AND U1313 ( .A(n46), .B(n1354), .Z(n1353) );
  XOR U1314 ( .A(p_input[29]), .B(n1352), .Z(n1354) );
  XNOR U1315 ( .A(n1355), .B(n1356), .Z(n1352) );
  AND U1316 ( .A(n50), .B(n1351), .Z(n1356) );
  XNOR U1317 ( .A(n1355), .B(n1349), .Z(n1351) );
  XOR U1318 ( .A(n1357), .B(n1358), .Z(n1349) );
  AND U1319 ( .A(n65), .B(n1359), .Z(n1358) );
  XNOR U1320 ( .A(n1360), .B(n1361), .Z(n1355) );
  AND U1321 ( .A(n57), .B(n1362), .Z(n1361) );
  XOR U1322 ( .A(p_input[45]), .B(n1360), .Z(n1362) );
  XNOR U1323 ( .A(n1363), .B(n1364), .Z(n1360) );
  AND U1324 ( .A(n61), .B(n1359), .Z(n1364) );
  XNOR U1325 ( .A(n1363), .B(n1357), .Z(n1359) );
  XOR U1326 ( .A(n1365), .B(n1366), .Z(n1357) );
  AND U1327 ( .A(n76), .B(n1367), .Z(n1366) );
  XNOR U1328 ( .A(n1368), .B(n1369), .Z(n1363) );
  AND U1329 ( .A(n68), .B(n1370), .Z(n1369) );
  XOR U1330 ( .A(p_input[61]), .B(n1368), .Z(n1370) );
  XNOR U1331 ( .A(n1371), .B(n1372), .Z(n1368) );
  AND U1332 ( .A(n72), .B(n1367), .Z(n1372) );
  XNOR U1333 ( .A(n1371), .B(n1365), .Z(n1367) );
  XOR U1334 ( .A(n1373), .B(n1374), .Z(n1365) );
  AND U1335 ( .A(n87), .B(n1375), .Z(n1374) );
  XNOR U1336 ( .A(n1376), .B(n1377), .Z(n1371) );
  AND U1337 ( .A(n79), .B(n1378), .Z(n1377) );
  XOR U1338 ( .A(p_input[77]), .B(n1376), .Z(n1378) );
  XNOR U1339 ( .A(n1379), .B(n1380), .Z(n1376) );
  AND U1340 ( .A(n83), .B(n1375), .Z(n1380) );
  XNOR U1341 ( .A(n1379), .B(n1373), .Z(n1375) );
  XOR U1342 ( .A(n1381), .B(n1382), .Z(n1373) );
  AND U1343 ( .A(n98), .B(n1383), .Z(n1382) );
  XNOR U1344 ( .A(n1384), .B(n1385), .Z(n1379) );
  AND U1345 ( .A(n90), .B(n1386), .Z(n1385) );
  XOR U1346 ( .A(p_input[93]), .B(n1384), .Z(n1386) );
  XNOR U1347 ( .A(n1387), .B(n1388), .Z(n1384) );
  AND U1348 ( .A(n94), .B(n1383), .Z(n1388) );
  XNOR U1349 ( .A(n1387), .B(n1381), .Z(n1383) );
  XOR U1350 ( .A(n1389), .B(n1390), .Z(n1381) );
  AND U1351 ( .A(n109), .B(n1391), .Z(n1390) );
  XNOR U1352 ( .A(n1392), .B(n1393), .Z(n1387) );
  AND U1353 ( .A(n101), .B(n1394), .Z(n1393) );
  XOR U1354 ( .A(p_input[109]), .B(n1392), .Z(n1394) );
  XNOR U1355 ( .A(n1395), .B(n1396), .Z(n1392) );
  AND U1356 ( .A(n105), .B(n1391), .Z(n1396) );
  XNOR U1357 ( .A(n1395), .B(n1389), .Z(n1391) );
  XOR U1358 ( .A(n1397), .B(n1398), .Z(n1389) );
  AND U1359 ( .A(n120), .B(n1399), .Z(n1398) );
  XNOR U1360 ( .A(n1400), .B(n1401), .Z(n1395) );
  AND U1361 ( .A(n112), .B(n1402), .Z(n1401) );
  XOR U1362 ( .A(p_input[125]), .B(n1400), .Z(n1402) );
  XNOR U1363 ( .A(n1403), .B(n1404), .Z(n1400) );
  AND U1364 ( .A(n116), .B(n1399), .Z(n1404) );
  XNOR U1365 ( .A(n1403), .B(n1397), .Z(n1399) );
  XOR U1366 ( .A(n1405), .B(n1406), .Z(n1397) );
  AND U1367 ( .A(n131), .B(n1407), .Z(n1406) );
  XNOR U1368 ( .A(n1408), .B(n1409), .Z(n1403) );
  AND U1369 ( .A(n123), .B(n1410), .Z(n1409) );
  XOR U1370 ( .A(p_input[141]), .B(n1408), .Z(n1410) );
  XNOR U1371 ( .A(n1411), .B(n1412), .Z(n1408) );
  AND U1372 ( .A(n127), .B(n1407), .Z(n1412) );
  XNOR U1373 ( .A(n1411), .B(n1405), .Z(n1407) );
  XOR U1374 ( .A(n1413), .B(n1414), .Z(n1405) );
  AND U1375 ( .A(n142), .B(n1415), .Z(n1414) );
  XNOR U1376 ( .A(n1416), .B(n1417), .Z(n1411) );
  AND U1377 ( .A(n134), .B(n1418), .Z(n1417) );
  XOR U1378 ( .A(p_input[157]), .B(n1416), .Z(n1418) );
  XNOR U1379 ( .A(n1419), .B(n1420), .Z(n1416) );
  AND U1380 ( .A(n138), .B(n1415), .Z(n1420) );
  XNOR U1381 ( .A(n1419), .B(n1413), .Z(n1415) );
  XOR U1382 ( .A(n1421), .B(n1422), .Z(n1413) );
  AND U1383 ( .A(n153), .B(n1423), .Z(n1422) );
  XNOR U1384 ( .A(n1424), .B(n1425), .Z(n1419) );
  AND U1385 ( .A(n145), .B(n1426), .Z(n1425) );
  XOR U1386 ( .A(p_input[173]), .B(n1424), .Z(n1426) );
  XNOR U1387 ( .A(n1427), .B(n1428), .Z(n1424) );
  AND U1388 ( .A(n149), .B(n1423), .Z(n1428) );
  XNOR U1389 ( .A(n1427), .B(n1421), .Z(n1423) );
  XOR U1390 ( .A(n1429), .B(n1430), .Z(n1421) );
  AND U1391 ( .A(n164), .B(n1431), .Z(n1430) );
  XNOR U1392 ( .A(n1432), .B(n1433), .Z(n1427) );
  AND U1393 ( .A(n156), .B(n1434), .Z(n1433) );
  XOR U1394 ( .A(p_input[189]), .B(n1432), .Z(n1434) );
  XNOR U1395 ( .A(n1435), .B(n1436), .Z(n1432) );
  AND U1396 ( .A(n160), .B(n1431), .Z(n1436) );
  XNOR U1397 ( .A(n1435), .B(n1429), .Z(n1431) );
  XOR U1398 ( .A(n1437), .B(n1438), .Z(n1429) );
  AND U1399 ( .A(n175), .B(n1439), .Z(n1438) );
  XNOR U1400 ( .A(n1440), .B(n1441), .Z(n1435) );
  AND U1401 ( .A(n167), .B(n1442), .Z(n1441) );
  XOR U1402 ( .A(p_input[205]), .B(n1440), .Z(n1442) );
  XNOR U1403 ( .A(n1443), .B(n1444), .Z(n1440) );
  AND U1404 ( .A(n171), .B(n1439), .Z(n1444) );
  XNOR U1405 ( .A(n1443), .B(n1437), .Z(n1439) );
  XOR U1406 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n1445), .Z(n1437) );
  AND U1407 ( .A(n185), .B(n1446), .Z(n1445) );
  XNOR U1408 ( .A(n1447), .B(n1448), .Z(n1443) );
  AND U1409 ( .A(n178), .B(n1449), .Z(n1448) );
  XOR U1410 ( .A(p_input[221]), .B(n1447), .Z(n1449) );
  XNOR U1411 ( .A(n1450), .B(n1451), .Z(n1447) );
  AND U1412 ( .A(n182), .B(n1446), .Z(n1451) );
  XOR U1413 ( .A(\knn_comb_/min_val_out[0][13] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n1446) );
  XOR U1414 ( .A(n23), .B(n1452), .Z(o[12]) );
  AND U1415 ( .A(n30), .B(n1453), .Z(n23) );
  XOR U1416 ( .A(n24), .B(n1452), .Z(n1453) );
  XOR U1417 ( .A(n1454), .B(n1455), .Z(n1452) );
  AND U1418 ( .A(n42), .B(n1456), .Z(n1455) );
  XOR U1419 ( .A(n1457), .B(n1458), .Z(n24) );
  AND U1420 ( .A(n34), .B(n1459), .Z(n1458) );
  XOR U1421 ( .A(p_input[12]), .B(n1457), .Z(n1459) );
  XNOR U1422 ( .A(n1460), .B(n1461), .Z(n1457) );
  AND U1423 ( .A(n38), .B(n1456), .Z(n1461) );
  XNOR U1424 ( .A(n1460), .B(n1454), .Z(n1456) );
  XOR U1425 ( .A(n1462), .B(n1463), .Z(n1454) );
  AND U1426 ( .A(n54), .B(n1464), .Z(n1463) );
  XNOR U1427 ( .A(n1465), .B(n1466), .Z(n1460) );
  AND U1428 ( .A(n46), .B(n1467), .Z(n1466) );
  XOR U1429 ( .A(p_input[28]), .B(n1465), .Z(n1467) );
  XNOR U1430 ( .A(n1468), .B(n1469), .Z(n1465) );
  AND U1431 ( .A(n50), .B(n1464), .Z(n1469) );
  XNOR U1432 ( .A(n1468), .B(n1462), .Z(n1464) );
  XOR U1433 ( .A(n1470), .B(n1471), .Z(n1462) );
  AND U1434 ( .A(n65), .B(n1472), .Z(n1471) );
  XNOR U1435 ( .A(n1473), .B(n1474), .Z(n1468) );
  AND U1436 ( .A(n57), .B(n1475), .Z(n1474) );
  XOR U1437 ( .A(p_input[44]), .B(n1473), .Z(n1475) );
  XNOR U1438 ( .A(n1476), .B(n1477), .Z(n1473) );
  AND U1439 ( .A(n61), .B(n1472), .Z(n1477) );
  XNOR U1440 ( .A(n1476), .B(n1470), .Z(n1472) );
  XOR U1441 ( .A(n1478), .B(n1479), .Z(n1470) );
  AND U1442 ( .A(n76), .B(n1480), .Z(n1479) );
  XNOR U1443 ( .A(n1481), .B(n1482), .Z(n1476) );
  AND U1444 ( .A(n68), .B(n1483), .Z(n1482) );
  XOR U1445 ( .A(p_input[60]), .B(n1481), .Z(n1483) );
  XNOR U1446 ( .A(n1484), .B(n1485), .Z(n1481) );
  AND U1447 ( .A(n72), .B(n1480), .Z(n1485) );
  XNOR U1448 ( .A(n1484), .B(n1478), .Z(n1480) );
  XOR U1449 ( .A(n1486), .B(n1487), .Z(n1478) );
  AND U1450 ( .A(n87), .B(n1488), .Z(n1487) );
  XNOR U1451 ( .A(n1489), .B(n1490), .Z(n1484) );
  AND U1452 ( .A(n79), .B(n1491), .Z(n1490) );
  XOR U1453 ( .A(p_input[76]), .B(n1489), .Z(n1491) );
  XNOR U1454 ( .A(n1492), .B(n1493), .Z(n1489) );
  AND U1455 ( .A(n83), .B(n1488), .Z(n1493) );
  XNOR U1456 ( .A(n1492), .B(n1486), .Z(n1488) );
  XOR U1457 ( .A(n1494), .B(n1495), .Z(n1486) );
  AND U1458 ( .A(n98), .B(n1496), .Z(n1495) );
  XNOR U1459 ( .A(n1497), .B(n1498), .Z(n1492) );
  AND U1460 ( .A(n90), .B(n1499), .Z(n1498) );
  XOR U1461 ( .A(p_input[92]), .B(n1497), .Z(n1499) );
  XNOR U1462 ( .A(n1500), .B(n1501), .Z(n1497) );
  AND U1463 ( .A(n94), .B(n1496), .Z(n1501) );
  XNOR U1464 ( .A(n1500), .B(n1494), .Z(n1496) );
  XOR U1465 ( .A(n1502), .B(n1503), .Z(n1494) );
  AND U1466 ( .A(n109), .B(n1504), .Z(n1503) );
  XNOR U1467 ( .A(n1505), .B(n1506), .Z(n1500) );
  AND U1468 ( .A(n101), .B(n1507), .Z(n1506) );
  XOR U1469 ( .A(p_input[108]), .B(n1505), .Z(n1507) );
  XNOR U1470 ( .A(n1508), .B(n1509), .Z(n1505) );
  AND U1471 ( .A(n105), .B(n1504), .Z(n1509) );
  XNOR U1472 ( .A(n1508), .B(n1502), .Z(n1504) );
  XOR U1473 ( .A(n1510), .B(n1511), .Z(n1502) );
  AND U1474 ( .A(n120), .B(n1512), .Z(n1511) );
  XNOR U1475 ( .A(n1513), .B(n1514), .Z(n1508) );
  AND U1476 ( .A(n112), .B(n1515), .Z(n1514) );
  XOR U1477 ( .A(p_input[124]), .B(n1513), .Z(n1515) );
  XNOR U1478 ( .A(n1516), .B(n1517), .Z(n1513) );
  AND U1479 ( .A(n116), .B(n1512), .Z(n1517) );
  XNOR U1480 ( .A(n1516), .B(n1510), .Z(n1512) );
  XOR U1481 ( .A(n1518), .B(n1519), .Z(n1510) );
  AND U1482 ( .A(n131), .B(n1520), .Z(n1519) );
  XNOR U1483 ( .A(n1521), .B(n1522), .Z(n1516) );
  AND U1484 ( .A(n123), .B(n1523), .Z(n1522) );
  XOR U1485 ( .A(p_input[140]), .B(n1521), .Z(n1523) );
  XNOR U1486 ( .A(n1524), .B(n1525), .Z(n1521) );
  AND U1487 ( .A(n127), .B(n1520), .Z(n1525) );
  XNOR U1488 ( .A(n1524), .B(n1518), .Z(n1520) );
  XOR U1489 ( .A(n1526), .B(n1527), .Z(n1518) );
  AND U1490 ( .A(n142), .B(n1528), .Z(n1527) );
  XNOR U1491 ( .A(n1529), .B(n1530), .Z(n1524) );
  AND U1492 ( .A(n134), .B(n1531), .Z(n1530) );
  XOR U1493 ( .A(p_input[156]), .B(n1529), .Z(n1531) );
  XNOR U1494 ( .A(n1532), .B(n1533), .Z(n1529) );
  AND U1495 ( .A(n138), .B(n1528), .Z(n1533) );
  XNOR U1496 ( .A(n1532), .B(n1526), .Z(n1528) );
  XOR U1497 ( .A(n1534), .B(n1535), .Z(n1526) );
  AND U1498 ( .A(n153), .B(n1536), .Z(n1535) );
  XNOR U1499 ( .A(n1537), .B(n1538), .Z(n1532) );
  AND U1500 ( .A(n145), .B(n1539), .Z(n1538) );
  XOR U1501 ( .A(p_input[172]), .B(n1537), .Z(n1539) );
  XNOR U1502 ( .A(n1540), .B(n1541), .Z(n1537) );
  AND U1503 ( .A(n149), .B(n1536), .Z(n1541) );
  XNOR U1504 ( .A(n1540), .B(n1534), .Z(n1536) );
  XOR U1505 ( .A(n1542), .B(n1543), .Z(n1534) );
  AND U1506 ( .A(n164), .B(n1544), .Z(n1543) );
  XNOR U1507 ( .A(n1545), .B(n1546), .Z(n1540) );
  AND U1508 ( .A(n156), .B(n1547), .Z(n1546) );
  XOR U1509 ( .A(p_input[188]), .B(n1545), .Z(n1547) );
  XNOR U1510 ( .A(n1548), .B(n1549), .Z(n1545) );
  AND U1511 ( .A(n160), .B(n1544), .Z(n1549) );
  XNOR U1512 ( .A(n1548), .B(n1542), .Z(n1544) );
  XOR U1513 ( .A(n1550), .B(n1551), .Z(n1542) );
  AND U1514 ( .A(n175), .B(n1552), .Z(n1551) );
  XNOR U1515 ( .A(n1553), .B(n1554), .Z(n1548) );
  AND U1516 ( .A(n167), .B(n1555), .Z(n1554) );
  XOR U1517 ( .A(p_input[204]), .B(n1553), .Z(n1555) );
  XNOR U1518 ( .A(n1556), .B(n1557), .Z(n1553) );
  AND U1519 ( .A(n171), .B(n1552), .Z(n1557) );
  XNOR U1520 ( .A(n1556), .B(n1550), .Z(n1552) );
  XOR U1521 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n1558), .Z(n1550) );
  AND U1522 ( .A(n185), .B(n1559), .Z(n1558) );
  XNOR U1523 ( .A(n1560), .B(n1561), .Z(n1556) );
  AND U1524 ( .A(n178), .B(n1562), .Z(n1561) );
  XOR U1525 ( .A(p_input[220]), .B(n1560), .Z(n1562) );
  XNOR U1526 ( .A(n1563), .B(n1564), .Z(n1560) );
  AND U1527 ( .A(n182), .B(n1559), .Z(n1564) );
  XOR U1528 ( .A(\knn_comb_/min_val_out[0][12] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n1559) );
  XOR U1529 ( .A(n25), .B(n1565), .Z(o[11]) );
  AND U1530 ( .A(n30), .B(n1566), .Z(n25) );
  XOR U1531 ( .A(n26), .B(n1565), .Z(n1566) );
  XOR U1532 ( .A(n1567), .B(n1568), .Z(n1565) );
  AND U1533 ( .A(n42), .B(n1569), .Z(n1568) );
  XOR U1534 ( .A(n1570), .B(n1571), .Z(n26) );
  AND U1535 ( .A(n34), .B(n1572), .Z(n1571) );
  XOR U1536 ( .A(p_input[11]), .B(n1570), .Z(n1572) );
  XNOR U1537 ( .A(n1573), .B(n1574), .Z(n1570) );
  AND U1538 ( .A(n38), .B(n1569), .Z(n1574) );
  XNOR U1539 ( .A(n1573), .B(n1567), .Z(n1569) );
  XOR U1540 ( .A(n1575), .B(n1576), .Z(n1567) );
  AND U1541 ( .A(n54), .B(n1577), .Z(n1576) );
  XNOR U1542 ( .A(n1578), .B(n1579), .Z(n1573) );
  AND U1543 ( .A(n46), .B(n1580), .Z(n1579) );
  XOR U1544 ( .A(p_input[27]), .B(n1578), .Z(n1580) );
  XNOR U1545 ( .A(n1581), .B(n1582), .Z(n1578) );
  AND U1546 ( .A(n50), .B(n1577), .Z(n1582) );
  XNOR U1547 ( .A(n1581), .B(n1575), .Z(n1577) );
  XOR U1548 ( .A(n1583), .B(n1584), .Z(n1575) );
  AND U1549 ( .A(n65), .B(n1585), .Z(n1584) );
  XNOR U1550 ( .A(n1586), .B(n1587), .Z(n1581) );
  AND U1551 ( .A(n57), .B(n1588), .Z(n1587) );
  XOR U1552 ( .A(p_input[43]), .B(n1586), .Z(n1588) );
  XNOR U1553 ( .A(n1589), .B(n1590), .Z(n1586) );
  AND U1554 ( .A(n61), .B(n1585), .Z(n1590) );
  XNOR U1555 ( .A(n1589), .B(n1583), .Z(n1585) );
  XOR U1556 ( .A(n1591), .B(n1592), .Z(n1583) );
  AND U1557 ( .A(n76), .B(n1593), .Z(n1592) );
  XNOR U1558 ( .A(n1594), .B(n1595), .Z(n1589) );
  AND U1559 ( .A(n68), .B(n1596), .Z(n1595) );
  XOR U1560 ( .A(p_input[59]), .B(n1594), .Z(n1596) );
  XNOR U1561 ( .A(n1597), .B(n1598), .Z(n1594) );
  AND U1562 ( .A(n72), .B(n1593), .Z(n1598) );
  XNOR U1563 ( .A(n1597), .B(n1591), .Z(n1593) );
  XOR U1564 ( .A(n1599), .B(n1600), .Z(n1591) );
  AND U1565 ( .A(n87), .B(n1601), .Z(n1600) );
  XNOR U1566 ( .A(n1602), .B(n1603), .Z(n1597) );
  AND U1567 ( .A(n79), .B(n1604), .Z(n1603) );
  XOR U1568 ( .A(p_input[75]), .B(n1602), .Z(n1604) );
  XNOR U1569 ( .A(n1605), .B(n1606), .Z(n1602) );
  AND U1570 ( .A(n83), .B(n1601), .Z(n1606) );
  XNOR U1571 ( .A(n1605), .B(n1599), .Z(n1601) );
  XOR U1572 ( .A(n1607), .B(n1608), .Z(n1599) );
  AND U1573 ( .A(n98), .B(n1609), .Z(n1608) );
  XNOR U1574 ( .A(n1610), .B(n1611), .Z(n1605) );
  AND U1575 ( .A(n90), .B(n1612), .Z(n1611) );
  XOR U1576 ( .A(p_input[91]), .B(n1610), .Z(n1612) );
  XNOR U1577 ( .A(n1613), .B(n1614), .Z(n1610) );
  AND U1578 ( .A(n94), .B(n1609), .Z(n1614) );
  XNOR U1579 ( .A(n1613), .B(n1607), .Z(n1609) );
  XOR U1580 ( .A(n1615), .B(n1616), .Z(n1607) );
  AND U1581 ( .A(n109), .B(n1617), .Z(n1616) );
  XNOR U1582 ( .A(n1618), .B(n1619), .Z(n1613) );
  AND U1583 ( .A(n101), .B(n1620), .Z(n1619) );
  XOR U1584 ( .A(p_input[107]), .B(n1618), .Z(n1620) );
  XNOR U1585 ( .A(n1621), .B(n1622), .Z(n1618) );
  AND U1586 ( .A(n105), .B(n1617), .Z(n1622) );
  XNOR U1587 ( .A(n1621), .B(n1615), .Z(n1617) );
  XOR U1588 ( .A(n1623), .B(n1624), .Z(n1615) );
  AND U1589 ( .A(n120), .B(n1625), .Z(n1624) );
  XNOR U1590 ( .A(n1626), .B(n1627), .Z(n1621) );
  AND U1591 ( .A(n112), .B(n1628), .Z(n1627) );
  XOR U1592 ( .A(p_input[123]), .B(n1626), .Z(n1628) );
  XNOR U1593 ( .A(n1629), .B(n1630), .Z(n1626) );
  AND U1594 ( .A(n116), .B(n1625), .Z(n1630) );
  XNOR U1595 ( .A(n1629), .B(n1623), .Z(n1625) );
  XOR U1596 ( .A(n1631), .B(n1632), .Z(n1623) );
  AND U1597 ( .A(n131), .B(n1633), .Z(n1632) );
  XNOR U1598 ( .A(n1634), .B(n1635), .Z(n1629) );
  AND U1599 ( .A(n123), .B(n1636), .Z(n1635) );
  XOR U1600 ( .A(p_input[139]), .B(n1634), .Z(n1636) );
  XNOR U1601 ( .A(n1637), .B(n1638), .Z(n1634) );
  AND U1602 ( .A(n127), .B(n1633), .Z(n1638) );
  XNOR U1603 ( .A(n1637), .B(n1631), .Z(n1633) );
  XOR U1604 ( .A(n1639), .B(n1640), .Z(n1631) );
  AND U1605 ( .A(n142), .B(n1641), .Z(n1640) );
  XNOR U1606 ( .A(n1642), .B(n1643), .Z(n1637) );
  AND U1607 ( .A(n134), .B(n1644), .Z(n1643) );
  XOR U1608 ( .A(p_input[155]), .B(n1642), .Z(n1644) );
  XNOR U1609 ( .A(n1645), .B(n1646), .Z(n1642) );
  AND U1610 ( .A(n138), .B(n1641), .Z(n1646) );
  XNOR U1611 ( .A(n1645), .B(n1639), .Z(n1641) );
  XOR U1612 ( .A(n1647), .B(n1648), .Z(n1639) );
  AND U1613 ( .A(n153), .B(n1649), .Z(n1648) );
  XNOR U1614 ( .A(n1650), .B(n1651), .Z(n1645) );
  AND U1615 ( .A(n145), .B(n1652), .Z(n1651) );
  XOR U1616 ( .A(p_input[171]), .B(n1650), .Z(n1652) );
  XNOR U1617 ( .A(n1653), .B(n1654), .Z(n1650) );
  AND U1618 ( .A(n149), .B(n1649), .Z(n1654) );
  XNOR U1619 ( .A(n1653), .B(n1647), .Z(n1649) );
  XOR U1620 ( .A(n1655), .B(n1656), .Z(n1647) );
  AND U1621 ( .A(n164), .B(n1657), .Z(n1656) );
  XNOR U1622 ( .A(n1658), .B(n1659), .Z(n1653) );
  AND U1623 ( .A(n156), .B(n1660), .Z(n1659) );
  XOR U1624 ( .A(p_input[187]), .B(n1658), .Z(n1660) );
  XNOR U1625 ( .A(n1661), .B(n1662), .Z(n1658) );
  AND U1626 ( .A(n160), .B(n1657), .Z(n1662) );
  XNOR U1627 ( .A(n1661), .B(n1655), .Z(n1657) );
  XOR U1628 ( .A(n1663), .B(n1664), .Z(n1655) );
  AND U1629 ( .A(n175), .B(n1665), .Z(n1664) );
  XNOR U1630 ( .A(n1666), .B(n1667), .Z(n1661) );
  AND U1631 ( .A(n167), .B(n1668), .Z(n1667) );
  XOR U1632 ( .A(p_input[203]), .B(n1666), .Z(n1668) );
  XNOR U1633 ( .A(n1669), .B(n1670), .Z(n1666) );
  AND U1634 ( .A(n171), .B(n1665), .Z(n1670) );
  XNOR U1635 ( .A(n1669), .B(n1663), .Z(n1665) );
  XOR U1636 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n1671), .Z(n1663) );
  AND U1637 ( .A(n185), .B(n1672), .Z(n1671) );
  XNOR U1638 ( .A(n1673), .B(n1674), .Z(n1669) );
  AND U1639 ( .A(n178), .B(n1675), .Z(n1674) );
  XOR U1640 ( .A(p_input[219]), .B(n1673), .Z(n1675) );
  XNOR U1641 ( .A(n1676), .B(n1677), .Z(n1673) );
  AND U1642 ( .A(n182), .B(n1672), .Z(n1677) );
  XOR U1643 ( .A(n1678), .B(n1676), .Z(n1672) );
  IV U1644 ( .A(\knn_comb_/min_val_out[0][11] ), .Z(n1678) );
  IV U1645 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n1676) );
  XOR U1646 ( .A(n27), .B(n1679), .Z(o[10]) );
  AND U1647 ( .A(n30), .B(n1680), .Z(n27) );
  XOR U1648 ( .A(n28), .B(n1679), .Z(n1680) );
  XOR U1649 ( .A(n1681), .B(n1682), .Z(n1679) );
  AND U1650 ( .A(n42), .B(n1683), .Z(n1682) );
  XOR U1651 ( .A(n1684), .B(n1685), .Z(n28) );
  AND U1652 ( .A(n34), .B(n1686), .Z(n1685) );
  XOR U1653 ( .A(p_input[10]), .B(n1684), .Z(n1686) );
  XNOR U1654 ( .A(n1687), .B(n1688), .Z(n1684) );
  AND U1655 ( .A(n38), .B(n1683), .Z(n1688) );
  XNOR U1656 ( .A(n1687), .B(n1681), .Z(n1683) );
  XOR U1657 ( .A(n1689), .B(n1690), .Z(n1681) );
  AND U1658 ( .A(n54), .B(n1691), .Z(n1690) );
  XNOR U1659 ( .A(n1692), .B(n1693), .Z(n1687) );
  AND U1660 ( .A(n46), .B(n1694), .Z(n1693) );
  XOR U1661 ( .A(p_input[26]), .B(n1692), .Z(n1694) );
  XNOR U1662 ( .A(n1695), .B(n1696), .Z(n1692) );
  AND U1663 ( .A(n50), .B(n1691), .Z(n1696) );
  XNOR U1664 ( .A(n1695), .B(n1689), .Z(n1691) );
  XOR U1665 ( .A(n1697), .B(n1698), .Z(n1689) );
  AND U1666 ( .A(n65), .B(n1699), .Z(n1698) );
  XNOR U1667 ( .A(n1700), .B(n1701), .Z(n1695) );
  AND U1668 ( .A(n57), .B(n1702), .Z(n1701) );
  XOR U1669 ( .A(p_input[42]), .B(n1700), .Z(n1702) );
  XNOR U1670 ( .A(n1703), .B(n1704), .Z(n1700) );
  AND U1671 ( .A(n61), .B(n1699), .Z(n1704) );
  XNOR U1672 ( .A(n1703), .B(n1697), .Z(n1699) );
  XOR U1673 ( .A(n1705), .B(n1706), .Z(n1697) );
  AND U1674 ( .A(n76), .B(n1707), .Z(n1706) );
  XNOR U1675 ( .A(n1708), .B(n1709), .Z(n1703) );
  AND U1676 ( .A(n68), .B(n1710), .Z(n1709) );
  XOR U1677 ( .A(p_input[58]), .B(n1708), .Z(n1710) );
  XNOR U1678 ( .A(n1711), .B(n1712), .Z(n1708) );
  AND U1679 ( .A(n72), .B(n1707), .Z(n1712) );
  XNOR U1680 ( .A(n1711), .B(n1705), .Z(n1707) );
  XOR U1681 ( .A(n1713), .B(n1714), .Z(n1705) );
  AND U1682 ( .A(n87), .B(n1715), .Z(n1714) );
  XNOR U1683 ( .A(n1716), .B(n1717), .Z(n1711) );
  AND U1684 ( .A(n79), .B(n1718), .Z(n1717) );
  XOR U1685 ( .A(p_input[74]), .B(n1716), .Z(n1718) );
  XNOR U1686 ( .A(n1719), .B(n1720), .Z(n1716) );
  AND U1687 ( .A(n83), .B(n1715), .Z(n1720) );
  XNOR U1688 ( .A(n1719), .B(n1713), .Z(n1715) );
  XOR U1689 ( .A(n1721), .B(n1722), .Z(n1713) );
  AND U1690 ( .A(n98), .B(n1723), .Z(n1722) );
  XNOR U1691 ( .A(n1724), .B(n1725), .Z(n1719) );
  AND U1692 ( .A(n90), .B(n1726), .Z(n1725) );
  XOR U1693 ( .A(p_input[90]), .B(n1724), .Z(n1726) );
  XNOR U1694 ( .A(n1727), .B(n1728), .Z(n1724) );
  AND U1695 ( .A(n94), .B(n1723), .Z(n1728) );
  XNOR U1696 ( .A(n1727), .B(n1721), .Z(n1723) );
  XOR U1697 ( .A(n1729), .B(n1730), .Z(n1721) );
  AND U1698 ( .A(n109), .B(n1731), .Z(n1730) );
  XNOR U1699 ( .A(n1732), .B(n1733), .Z(n1727) );
  AND U1700 ( .A(n101), .B(n1734), .Z(n1733) );
  XOR U1701 ( .A(p_input[106]), .B(n1732), .Z(n1734) );
  XNOR U1702 ( .A(n1735), .B(n1736), .Z(n1732) );
  AND U1703 ( .A(n105), .B(n1731), .Z(n1736) );
  XNOR U1704 ( .A(n1735), .B(n1729), .Z(n1731) );
  XOR U1705 ( .A(n1737), .B(n1738), .Z(n1729) );
  AND U1706 ( .A(n120), .B(n1739), .Z(n1738) );
  XNOR U1707 ( .A(n1740), .B(n1741), .Z(n1735) );
  AND U1708 ( .A(n112), .B(n1742), .Z(n1741) );
  XOR U1709 ( .A(p_input[122]), .B(n1740), .Z(n1742) );
  XNOR U1710 ( .A(n1743), .B(n1744), .Z(n1740) );
  AND U1711 ( .A(n116), .B(n1739), .Z(n1744) );
  XNOR U1712 ( .A(n1743), .B(n1737), .Z(n1739) );
  XOR U1713 ( .A(n1745), .B(n1746), .Z(n1737) );
  AND U1714 ( .A(n131), .B(n1747), .Z(n1746) );
  XNOR U1715 ( .A(n1748), .B(n1749), .Z(n1743) );
  AND U1716 ( .A(n123), .B(n1750), .Z(n1749) );
  XOR U1717 ( .A(p_input[138]), .B(n1748), .Z(n1750) );
  XNOR U1718 ( .A(n1751), .B(n1752), .Z(n1748) );
  AND U1719 ( .A(n127), .B(n1747), .Z(n1752) );
  XNOR U1720 ( .A(n1751), .B(n1745), .Z(n1747) );
  XOR U1721 ( .A(n1753), .B(n1754), .Z(n1745) );
  AND U1722 ( .A(n142), .B(n1755), .Z(n1754) );
  XNOR U1723 ( .A(n1756), .B(n1757), .Z(n1751) );
  AND U1724 ( .A(n134), .B(n1758), .Z(n1757) );
  XOR U1725 ( .A(p_input[154]), .B(n1756), .Z(n1758) );
  XNOR U1726 ( .A(n1759), .B(n1760), .Z(n1756) );
  AND U1727 ( .A(n138), .B(n1755), .Z(n1760) );
  XNOR U1728 ( .A(n1759), .B(n1753), .Z(n1755) );
  XOR U1729 ( .A(n1761), .B(n1762), .Z(n1753) );
  AND U1730 ( .A(n153), .B(n1763), .Z(n1762) );
  XNOR U1731 ( .A(n1764), .B(n1765), .Z(n1759) );
  AND U1732 ( .A(n145), .B(n1766), .Z(n1765) );
  XOR U1733 ( .A(p_input[170]), .B(n1764), .Z(n1766) );
  XNOR U1734 ( .A(n1767), .B(n1768), .Z(n1764) );
  AND U1735 ( .A(n149), .B(n1763), .Z(n1768) );
  XNOR U1736 ( .A(n1767), .B(n1761), .Z(n1763) );
  XOR U1737 ( .A(n1769), .B(n1770), .Z(n1761) );
  AND U1738 ( .A(n164), .B(n1771), .Z(n1770) );
  XNOR U1739 ( .A(n1772), .B(n1773), .Z(n1767) );
  AND U1740 ( .A(n156), .B(n1774), .Z(n1773) );
  XOR U1741 ( .A(p_input[186]), .B(n1772), .Z(n1774) );
  XNOR U1742 ( .A(n1775), .B(n1776), .Z(n1772) );
  AND U1743 ( .A(n160), .B(n1771), .Z(n1776) );
  XNOR U1744 ( .A(n1775), .B(n1769), .Z(n1771) );
  XOR U1745 ( .A(n1777), .B(n1778), .Z(n1769) );
  AND U1746 ( .A(n175), .B(n1779), .Z(n1778) );
  XNOR U1747 ( .A(n1780), .B(n1781), .Z(n1775) );
  AND U1748 ( .A(n167), .B(n1782), .Z(n1781) );
  XOR U1749 ( .A(p_input[202]), .B(n1780), .Z(n1782) );
  XNOR U1750 ( .A(n1783), .B(n1784), .Z(n1780) );
  AND U1751 ( .A(n171), .B(n1779), .Z(n1784) );
  XNOR U1752 ( .A(n1783), .B(n1777), .Z(n1779) );
  XOR U1753 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n1785), .Z(n1777) );
  AND U1754 ( .A(n185), .B(n1786), .Z(n1785) );
  XNOR U1755 ( .A(n1787), .B(n1788), .Z(n1783) );
  AND U1756 ( .A(n178), .B(n1789), .Z(n1788) );
  XOR U1757 ( .A(p_input[218]), .B(n1787), .Z(n1789) );
  XNOR U1758 ( .A(n1790), .B(n1791), .Z(n1787) );
  AND U1759 ( .A(n182), .B(n1786), .Z(n1791) );
  XOR U1760 ( .A(\knn_comb_/min_val_out[0][10] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n1786) );
  XOR U1761 ( .A(n1109), .B(n1792), .Z(o[0]) );
  AND U1762 ( .A(n30), .B(n1793), .Z(n1109) );
  XOR U1763 ( .A(n1110), .B(n1792), .Z(n1793) );
  XOR U1764 ( .A(n1794), .B(n1795), .Z(n1792) );
  AND U1765 ( .A(n42), .B(n1796), .Z(n1795) );
  XOR U1766 ( .A(n1797), .B(n1798), .Z(n1110) );
  AND U1767 ( .A(n34), .B(n1799), .Z(n1798) );
  XOR U1768 ( .A(p_input[0]), .B(n1797), .Z(n1799) );
  XNOR U1769 ( .A(n1800), .B(n1801), .Z(n1797) );
  AND U1770 ( .A(n38), .B(n1796), .Z(n1801) );
  XNOR U1771 ( .A(n1800), .B(n1794), .Z(n1796) );
  XOR U1772 ( .A(n1802), .B(n1803), .Z(n1794) );
  AND U1773 ( .A(n54), .B(n1804), .Z(n1803) );
  XNOR U1774 ( .A(n1805), .B(n1806), .Z(n1800) );
  AND U1775 ( .A(n46), .B(n1807), .Z(n1806) );
  XOR U1776 ( .A(p_input[16]), .B(n1805), .Z(n1807) );
  XNOR U1777 ( .A(n1808), .B(n1809), .Z(n1805) );
  AND U1778 ( .A(n50), .B(n1804), .Z(n1809) );
  XNOR U1779 ( .A(n1808), .B(n1802), .Z(n1804) );
  XOR U1780 ( .A(n1810), .B(n1811), .Z(n1802) );
  AND U1781 ( .A(n65), .B(n1812), .Z(n1811) );
  XNOR U1782 ( .A(n1813), .B(n1814), .Z(n1808) );
  AND U1783 ( .A(n57), .B(n1815), .Z(n1814) );
  XOR U1784 ( .A(p_input[32]), .B(n1813), .Z(n1815) );
  XNOR U1785 ( .A(n1816), .B(n1817), .Z(n1813) );
  AND U1786 ( .A(n61), .B(n1812), .Z(n1817) );
  XNOR U1787 ( .A(n1816), .B(n1810), .Z(n1812) );
  XOR U1788 ( .A(n1818), .B(n1819), .Z(n1810) );
  AND U1789 ( .A(n76), .B(n1820), .Z(n1819) );
  XNOR U1790 ( .A(n1821), .B(n1822), .Z(n1816) );
  AND U1791 ( .A(n68), .B(n1823), .Z(n1822) );
  XOR U1792 ( .A(p_input[48]), .B(n1821), .Z(n1823) );
  XNOR U1793 ( .A(n1824), .B(n1825), .Z(n1821) );
  AND U1794 ( .A(n72), .B(n1820), .Z(n1825) );
  XNOR U1795 ( .A(n1824), .B(n1818), .Z(n1820) );
  XOR U1796 ( .A(n1826), .B(n1827), .Z(n1818) );
  AND U1797 ( .A(n87), .B(n1828), .Z(n1827) );
  XNOR U1798 ( .A(n1829), .B(n1830), .Z(n1824) );
  AND U1799 ( .A(n79), .B(n1831), .Z(n1830) );
  XOR U1800 ( .A(p_input[64]), .B(n1829), .Z(n1831) );
  XNOR U1801 ( .A(n1832), .B(n1833), .Z(n1829) );
  AND U1802 ( .A(n83), .B(n1828), .Z(n1833) );
  XNOR U1803 ( .A(n1832), .B(n1826), .Z(n1828) );
  XOR U1804 ( .A(n1834), .B(n1835), .Z(n1826) );
  AND U1805 ( .A(n98), .B(n1836), .Z(n1835) );
  XNOR U1806 ( .A(n1837), .B(n1838), .Z(n1832) );
  AND U1807 ( .A(n90), .B(n1839), .Z(n1838) );
  XOR U1808 ( .A(p_input[80]), .B(n1837), .Z(n1839) );
  XNOR U1809 ( .A(n1840), .B(n1841), .Z(n1837) );
  AND U1810 ( .A(n94), .B(n1836), .Z(n1841) );
  XNOR U1811 ( .A(n1840), .B(n1834), .Z(n1836) );
  XOR U1812 ( .A(n1842), .B(n1843), .Z(n1834) );
  AND U1813 ( .A(n109), .B(n1844), .Z(n1843) );
  XNOR U1814 ( .A(n1845), .B(n1846), .Z(n1840) );
  AND U1815 ( .A(n101), .B(n1847), .Z(n1846) );
  XOR U1816 ( .A(p_input[96]), .B(n1845), .Z(n1847) );
  XNOR U1817 ( .A(n1848), .B(n1849), .Z(n1845) );
  AND U1818 ( .A(n105), .B(n1844), .Z(n1849) );
  XNOR U1819 ( .A(n1848), .B(n1842), .Z(n1844) );
  XOR U1820 ( .A(n1850), .B(n1851), .Z(n1842) );
  AND U1821 ( .A(n120), .B(n1852), .Z(n1851) );
  XNOR U1822 ( .A(n1853), .B(n1854), .Z(n1848) );
  AND U1823 ( .A(n112), .B(n1855), .Z(n1854) );
  XOR U1824 ( .A(p_input[112]), .B(n1853), .Z(n1855) );
  XNOR U1825 ( .A(n1856), .B(n1857), .Z(n1853) );
  AND U1826 ( .A(n116), .B(n1852), .Z(n1857) );
  XNOR U1827 ( .A(n1856), .B(n1850), .Z(n1852) );
  XOR U1828 ( .A(n1858), .B(n1859), .Z(n1850) );
  AND U1829 ( .A(n131), .B(n1860), .Z(n1859) );
  XNOR U1830 ( .A(n1861), .B(n1862), .Z(n1856) );
  AND U1831 ( .A(n123), .B(n1863), .Z(n1862) );
  XOR U1832 ( .A(p_input[128]), .B(n1861), .Z(n1863) );
  XNOR U1833 ( .A(n1864), .B(n1865), .Z(n1861) );
  AND U1834 ( .A(n127), .B(n1860), .Z(n1865) );
  XNOR U1835 ( .A(n1864), .B(n1858), .Z(n1860) );
  XOR U1836 ( .A(n1866), .B(n1867), .Z(n1858) );
  AND U1837 ( .A(n142), .B(n1868), .Z(n1867) );
  XNOR U1838 ( .A(n1869), .B(n1870), .Z(n1864) );
  AND U1839 ( .A(n134), .B(n1871), .Z(n1870) );
  XOR U1840 ( .A(p_input[144]), .B(n1869), .Z(n1871) );
  XNOR U1841 ( .A(n1872), .B(n1873), .Z(n1869) );
  AND U1842 ( .A(n138), .B(n1868), .Z(n1873) );
  XNOR U1843 ( .A(n1872), .B(n1866), .Z(n1868) );
  XOR U1844 ( .A(n1874), .B(n1875), .Z(n1866) );
  AND U1845 ( .A(n153), .B(n1876), .Z(n1875) );
  XNOR U1846 ( .A(n1877), .B(n1878), .Z(n1872) );
  AND U1847 ( .A(n145), .B(n1879), .Z(n1878) );
  XOR U1848 ( .A(p_input[160]), .B(n1877), .Z(n1879) );
  XNOR U1849 ( .A(n1880), .B(n1881), .Z(n1877) );
  AND U1850 ( .A(n149), .B(n1876), .Z(n1881) );
  XNOR U1851 ( .A(n1880), .B(n1874), .Z(n1876) );
  XOR U1852 ( .A(n1882), .B(n1883), .Z(n1874) );
  AND U1853 ( .A(n164), .B(n1884), .Z(n1883) );
  XNOR U1854 ( .A(n1885), .B(n1886), .Z(n1880) );
  AND U1855 ( .A(n156), .B(n1887), .Z(n1886) );
  XOR U1856 ( .A(p_input[176]), .B(n1885), .Z(n1887) );
  XNOR U1857 ( .A(n1888), .B(n1889), .Z(n1885) );
  AND U1858 ( .A(n160), .B(n1884), .Z(n1889) );
  XNOR U1859 ( .A(n1888), .B(n1882), .Z(n1884) );
  XOR U1860 ( .A(n1890), .B(n1891), .Z(n1882) );
  AND U1861 ( .A(n175), .B(n1892), .Z(n1891) );
  XNOR U1862 ( .A(n1893), .B(n1894), .Z(n1888) );
  AND U1863 ( .A(n167), .B(n1895), .Z(n1894) );
  XOR U1864 ( .A(p_input[192]), .B(n1893), .Z(n1895) );
  XNOR U1865 ( .A(n1896), .B(n1897), .Z(n1893) );
  AND U1866 ( .A(n171), .B(n1892), .Z(n1897) );
  XNOR U1867 ( .A(n1896), .B(n1890), .Z(n1892) );
  XOR U1868 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n1898), .Z(n1890) );
  AND U1869 ( .A(n185), .B(n1899), .Z(n1898) );
  XNOR U1870 ( .A(n1900), .B(n1901), .Z(n1896) );
  AND U1871 ( .A(n178), .B(n1902), .Z(n1901) );
  XOR U1872 ( .A(p_input[208]), .B(n1900), .Z(n1902) );
  XNOR U1873 ( .A(n1903), .B(n1904), .Z(n1900) );
  AND U1874 ( .A(n182), .B(n1899), .Z(n1904) );
  XOR U1875 ( .A(\knn_comb_/min_val_out[0][0] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n1899) );
  IV U1876 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n1903) );
  XNOR U1877 ( .A(n1905), .B(n1906), .Z(n30) );
  AND U1878 ( .A(n1907), .B(n1908), .Z(n1906) );
  XNOR U1879 ( .A(n1905), .B(n1909), .Z(n1908) );
  XOR U1880 ( .A(n1910), .B(n1911), .Z(n1909) );
  AND U1881 ( .A(n34), .B(n1912), .Z(n1911) );
  XNOR U1882 ( .A(n1910), .B(n1913), .Z(n1912) );
  XNOR U1883 ( .A(n1905), .B(n1914), .Z(n1907) );
  XOR U1884 ( .A(n1915), .B(n1916), .Z(n1914) );
  AND U1885 ( .A(n42), .B(n1917), .Z(n1916) );
  XOR U1886 ( .A(n1918), .B(n1919), .Z(n1905) );
  AND U1887 ( .A(n1920), .B(n1921), .Z(n1919) );
  XOR U1888 ( .A(n1922), .B(n1918), .Z(n1921) );
  XOR U1889 ( .A(n1923), .B(n1924), .Z(n1922) );
  AND U1890 ( .A(n34), .B(n1925), .Z(n1924) );
  XOR U1891 ( .A(n1926), .B(n1923), .Z(n1925) );
  XNOR U1892 ( .A(n1918), .B(n1927), .Z(n1920) );
  XOR U1893 ( .A(n1928), .B(n1929), .Z(n1927) );
  AND U1894 ( .A(n42), .B(n1930), .Z(n1929) );
  XOR U1895 ( .A(n1931), .B(n1932), .Z(n1918) );
  AND U1896 ( .A(n1933), .B(n1934), .Z(n1932) );
  XOR U1897 ( .A(n1935), .B(n1931), .Z(n1934) );
  XOR U1898 ( .A(n1936), .B(n1937), .Z(n1935) );
  AND U1899 ( .A(n34), .B(n1938), .Z(n1937) );
  XNOR U1900 ( .A(n1939), .B(n1936), .Z(n1938) );
  XNOR U1901 ( .A(n1931), .B(n1940), .Z(n1933) );
  XOR U1902 ( .A(n1941), .B(n1942), .Z(n1940) );
  AND U1903 ( .A(n42), .B(n1943), .Z(n1942) );
  XOR U1904 ( .A(n1944), .B(n1945), .Z(n1931) );
  AND U1905 ( .A(n1946), .B(n1947), .Z(n1945) );
  XOR U1906 ( .A(n1944), .B(n1948), .Z(n1947) );
  XOR U1907 ( .A(n1949), .B(n1950), .Z(n1948) );
  AND U1908 ( .A(n34), .B(n1951), .Z(n1950) );
  XOR U1909 ( .A(n1952), .B(n1949), .Z(n1951) );
  XNOR U1910 ( .A(n1953), .B(n1944), .Z(n1946) );
  XNOR U1911 ( .A(n1954), .B(n1955), .Z(n1953) );
  AND U1912 ( .A(n42), .B(n1956), .Z(n1955) );
  AND U1913 ( .A(n1957), .B(n1958), .Z(n1944) );
  XNOR U1914 ( .A(n1959), .B(n1960), .Z(n1958) );
  AND U1915 ( .A(n34), .B(n1961), .Z(n1960) );
  XNOR U1916 ( .A(n1962), .B(n1959), .Z(n1961) );
  XNOR U1917 ( .A(n1963), .B(n1964), .Z(n34) );
  AND U1918 ( .A(n1965), .B(n1966), .Z(n1964) );
  XOR U1919 ( .A(n1913), .B(n1963), .Z(n1966) );
  AND U1920 ( .A(n1967), .B(n1968), .Z(n1913) );
  XOR U1921 ( .A(n1963), .B(n1910), .Z(n1965) );
  XNOR U1922 ( .A(n1969), .B(n1970), .Z(n1910) );
  AND U1923 ( .A(n38), .B(n1917), .Z(n1970) );
  XOR U1924 ( .A(n1915), .B(n1969), .Z(n1917) );
  XOR U1925 ( .A(n1971), .B(n1972), .Z(n1963) );
  AND U1926 ( .A(n1973), .B(n1974), .Z(n1972) );
  XNOR U1927 ( .A(n1971), .B(n1967), .Z(n1974) );
  IV U1928 ( .A(n1926), .Z(n1967) );
  XOR U1929 ( .A(n1975), .B(n1976), .Z(n1926) );
  XOR U1930 ( .A(n1977), .B(n1968), .Z(n1976) );
  AND U1931 ( .A(n1939), .B(n1978), .Z(n1968) );
  AND U1932 ( .A(n1979), .B(n1980), .Z(n1977) );
  XOR U1933 ( .A(n1981), .B(n1975), .Z(n1979) );
  XNOR U1934 ( .A(n1923), .B(n1971), .Z(n1973) );
  XNOR U1935 ( .A(n1982), .B(n1983), .Z(n1923) );
  AND U1936 ( .A(n38), .B(n1930), .Z(n1983) );
  XOR U1937 ( .A(n1982), .B(n1984), .Z(n1930) );
  XOR U1938 ( .A(n1985), .B(n1986), .Z(n1971) );
  AND U1939 ( .A(n1987), .B(n1988), .Z(n1986) );
  XNOR U1940 ( .A(n1985), .B(n1939), .Z(n1988) );
  XOR U1941 ( .A(n1989), .B(n1980), .Z(n1939) );
  XNOR U1942 ( .A(n1990), .B(n1975), .Z(n1980) );
  XOR U1943 ( .A(n1991), .B(n1992), .Z(n1975) );
  AND U1944 ( .A(n1993), .B(n1994), .Z(n1992) );
  XOR U1945 ( .A(n1995), .B(n1991), .Z(n1993) );
  XNOR U1946 ( .A(n1996), .B(n1997), .Z(n1990) );
  AND U1947 ( .A(n1998), .B(n1999), .Z(n1997) );
  XOR U1948 ( .A(n1996), .B(n2000), .Z(n1998) );
  XNOR U1949 ( .A(n1981), .B(n1978), .Z(n1989) );
  AND U1950 ( .A(n2001), .B(n2002), .Z(n1978) );
  XOR U1951 ( .A(n2003), .B(n2004), .Z(n1981) );
  AND U1952 ( .A(n2005), .B(n2006), .Z(n2004) );
  XOR U1953 ( .A(n2003), .B(n2007), .Z(n2005) );
  XNOR U1954 ( .A(n1936), .B(n1985), .Z(n1987) );
  XNOR U1955 ( .A(n2008), .B(n2009), .Z(n1936) );
  AND U1956 ( .A(n38), .B(n1943), .Z(n2009) );
  XOR U1957 ( .A(n2008), .B(n2010), .Z(n1943) );
  XOR U1958 ( .A(n2011), .B(n2012), .Z(n1985) );
  AND U1959 ( .A(n2013), .B(n2014), .Z(n2012) );
  XNOR U1960 ( .A(n2011), .B(n2001), .Z(n2014) );
  IV U1961 ( .A(n1952), .Z(n2001) );
  XNOR U1962 ( .A(n2015), .B(n1994), .Z(n1952) );
  XNOR U1963 ( .A(n2016), .B(n2000), .Z(n1994) );
  XNOR U1964 ( .A(n2017), .B(n2018), .Z(n2000) );
  NOR U1965 ( .A(n2019), .B(n2020), .Z(n2018) );
  XOR U1966 ( .A(n2017), .B(n2021), .Z(n2019) );
  XNOR U1967 ( .A(n1999), .B(n1991), .Z(n2016) );
  XOR U1968 ( .A(n2022), .B(n2023), .Z(n1991) );
  AND U1969 ( .A(n2024), .B(n2025), .Z(n2023) );
  XNOR U1970 ( .A(n2022), .B(n2026), .Z(n2024) );
  XNOR U1971 ( .A(n2027), .B(n1996), .Z(n1999) );
  XOR U1972 ( .A(n2028), .B(n2029), .Z(n1996) );
  AND U1973 ( .A(n2030), .B(n2031), .Z(n2029) );
  XOR U1974 ( .A(n2028), .B(n2032), .Z(n2030) );
  XNOR U1975 ( .A(n2033), .B(n2034), .Z(n2027) );
  NOR U1976 ( .A(n2035), .B(n2036), .Z(n2034) );
  XNOR U1977 ( .A(n2033), .B(n2037), .Z(n2035) );
  XNOR U1978 ( .A(n1995), .B(n2002), .Z(n2015) );
  NOR U1979 ( .A(n1962), .B(n2038), .Z(n2002) );
  XOR U1980 ( .A(n2007), .B(n2006), .Z(n1995) );
  XNOR U1981 ( .A(n2039), .B(n2003), .Z(n2006) );
  XOR U1982 ( .A(n2040), .B(n2041), .Z(n2003) );
  AND U1983 ( .A(n2042), .B(n2043), .Z(n2041) );
  XOR U1984 ( .A(n2040), .B(n2044), .Z(n2042) );
  XNOR U1985 ( .A(n2045), .B(n2046), .Z(n2039) );
  NOR U1986 ( .A(n2047), .B(n2048), .Z(n2046) );
  XNOR U1987 ( .A(n2045), .B(n2049), .Z(n2047) );
  XOR U1988 ( .A(n2050), .B(n2051), .Z(n2007) );
  NOR U1989 ( .A(n2052), .B(n2053), .Z(n2051) );
  XNOR U1990 ( .A(n2050), .B(n2054), .Z(n2052) );
  XNOR U1991 ( .A(n1949), .B(n2011), .Z(n2013) );
  XNOR U1992 ( .A(n2055), .B(n2056), .Z(n1949) );
  AND U1993 ( .A(n38), .B(n1956), .Z(n2056) );
  XOR U1994 ( .A(n2055), .B(n1954), .Z(n1956) );
  AND U1995 ( .A(n1959), .B(n1962), .Z(n2011) );
  XOR U1996 ( .A(n2057), .B(n2038), .Z(n1962) );
  XNOR U1997 ( .A(p_input[0]), .B(p_input[256]), .Z(n2038) );
  XOR U1998 ( .A(n2026), .B(n2025), .Z(n2057) );
  XNOR U1999 ( .A(n2058), .B(n2032), .Z(n2025) );
  XNOR U2000 ( .A(n2021), .B(n2020), .Z(n2032) );
  XNOR U2001 ( .A(n2059), .B(n2017), .Z(n2020) );
  XNOR U2002 ( .A(p_input[10]), .B(p_input[266]), .Z(n2017) );
  XOR U2003 ( .A(p_input[11]), .B(n2060), .Z(n2059) );
  XOR U2004 ( .A(p_input[12]), .B(p_input[268]), .Z(n2021) );
  XOR U2005 ( .A(n2031), .B(n2061), .Z(n2058) );
  IV U2006 ( .A(n2022), .Z(n2061) );
  XOR U2007 ( .A(p_input[1]), .B(p_input[257]), .Z(n2022) );
  XNOR U2008 ( .A(n2062), .B(n2037), .Z(n2031) );
  XNOR U2009 ( .A(p_input[15]), .B(n2063), .Z(n2037) );
  XOR U2010 ( .A(n2028), .B(n2036), .Z(n2062) );
  XOR U2011 ( .A(n2064), .B(n2033), .Z(n2036) );
  XOR U2012 ( .A(p_input[13]), .B(p_input[269]), .Z(n2033) );
  XOR U2013 ( .A(p_input[14]), .B(n2065), .Z(n2064) );
  XNOR U2014 ( .A(n2066), .B(p_input[9]), .Z(n2028) );
  XNOR U2015 ( .A(n2044), .B(n2043), .Z(n2026) );
  XNOR U2016 ( .A(n2067), .B(n2049), .Z(n2043) );
  XOR U2017 ( .A(p_input[264]), .B(p_input[8]), .Z(n2049) );
  XOR U2018 ( .A(n2040), .B(n2048), .Z(n2067) );
  XOR U2019 ( .A(n2068), .B(n2045), .Z(n2048) );
  XOR U2020 ( .A(p_input[262]), .B(p_input[6]), .Z(n2045) );
  XNOR U2021 ( .A(p_input[263]), .B(p_input[7]), .Z(n2068) );
  XNOR U2022 ( .A(n2069), .B(p_input[2]), .Z(n2040) );
  XNOR U2023 ( .A(n2054), .B(n2053), .Z(n2044) );
  XOR U2024 ( .A(n2070), .B(n2050), .Z(n2053) );
  XOR U2025 ( .A(p_input[259]), .B(p_input[3]), .Z(n2050) );
  XNOR U2026 ( .A(p_input[260]), .B(p_input[4]), .Z(n2070) );
  XOR U2027 ( .A(p_input[261]), .B(p_input[5]), .Z(n2054) );
  XNOR U2028 ( .A(n2071), .B(n2072), .Z(n1959) );
  AND U2029 ( .A(n38), .B(n2073), .Z(n2072) );
  XNOR U2030 ( .A(n2074), .B(n2075), .Z(n38) );
  AND U2031 ( .A(n2076), .B(n2077), .Z(n2075) );
  XOR U2032 ( .A(n2074), .B(n1969), .Z(n2077) );
  XNOR U2033 ( .A(n2074), .B(n1915), .Z(n2076) );
  XOR U2034 ( .A(n2078), .B(n2079), .Z(n2074) );
  AND U2035 ( .A(n2080), .B(n2081), .Z(n2079) );
  XNOR U2036 ( .A(n1982), .B(n2078), .Z(n2081) );
  XOR U2037 ( .A(n2078), .B(n1984), .Z(n2080) );
  XOR U2038 ( .A(n2082), .B(n2083), .Z(n2078) );
  AND U2039 ( .A(n2084), .B(n2085), .Z(n2083) );
  XOR U2040 ( .A(n2082), .B(n2010), .Z(n2084) );
  IV U2041 ( .A(n1941), .Z(n2010) );
  XOR U2042 ( .A(n2086), .B(n2087), .Z(n1957) );
  AND U2043 ( .A(n42), .B(n2073), .Z(n2087) );
  XNOR U2044 ( .A(n2071), .B(n2086), .Z(n2073) );
  XNOR U2045 ( .A(n2088), .B(n2089), .Z(n42) );
  AND U2046 ( .A(n2090), .B(n2091), .Z(n2089) );
  XNOR U2047 ( .A(n2092), .B(n2088), .Z(n2091) );
  IV U2048 ( .A(n1969), .Z(n2092) );
  XNOR U2049 ( .A(n2093), .B(n2094), .Z(n1969) );
  AND U2050 ( .A(n46), .B(n2095), .Z(n2094) );
  XNOR U2051 ( .A(n2093), .B(n2096), .Z(n2095) );
  XNOR U2052 ( .A(n1915), .B(n2088), .Z(n2090) );
  XOR U2053 ( .A(n2097), .B(n2098), .Z(n1915) );
  AND U2054 ( .A(n54), .B(n2099), .Z(n2098) );
  XOR U2055 ( .A(n2100), .B(n2101), .Z(n2088) );
  AND U2056 ( .A(n2102), .B(n2103), .Z(n2101) );
  XNOR U2057 ( .A(n2100), .B(n1982), .Z(n2103) );
  XNOR U2058 ( .A(n2104), .B(n2105), .Z(n1982) );
  AND U2059 ( .A(n46), .B(n2106), .Z(n2105) );
  XOR U2060 ( .A(n2107), .B(n2104), .Z(n2106) );
  XNOR U2061 ( .A(n1928), .B(n2100), .Z(n2102) );
  IV U2062 ( .A(n1984), .Z(n1928) );
  XOR U2063 ( .A(n2108), .B(n2109), .Z(n1984) );
  AND U2064 ( .A(n54), .B(n2110), .Z(n2109) );
  XOR U2065 ( .A(n2082), .B(n2111), .Z(n2100) );
  AND U2066 ( .A(n2112), .B(n2085), .Z(n2111) );
  XNOR U2067 ( .A(n2008), .B(n2082), .Z(n2085) );
  XNOR U2068 ( .A(n2113), .B(n2114), .Z(n2008) );
  AND U2069 ( .A(n46), .B(n2115), .Z(n2114) );
  XNOR U2070 ( .A(n2116), .B(n2113), .Z(n2115) );
  XNOR U2071 ( .A(n1941), .B(n2082), .Z(n2112) );
  XNOR U2072 ( .A(n2117), .B(n2118), .Z(n1941) );
  AND U2073 ( .A(n54), .B(n2119), .Z(n2118) );
  XOR U2074 ( .A(n2120), .B(n2121), .Z(n2082) );
  AND U2075 ( .A(n2122), .B(n2123), .Z(n2121) );
  XNOR U2076 ( .A(n2120), .B(n2055), .Z(n2123) );
  XNOR U2077 ( .A(n2124), .B(n2125), .Z(n2055) );
  AND U2078 ( .A(n46), .B(n2126), .Z(n2125) );
  XOR U2079 ( .A(n2127), .B(n2124), .Z(n2126) );
  XNOR U2080 ( .A(n2128), .B(n2120), .Z(n2122) );
  IV U2081 ( .A(n1954), .Z(n2128) );
  XOR U2082 ( .A(n2129), .B(n2130), .Z(n1954) );
  AND U2083 ( .A(n54), .B(n2131), .Z(n2130) );
  AND U2084 ( .A(n2086), .B(n2071), .Z(n2120) );
  XNOR U2085 ( .A(n2132), .B(n2133), .Z(n2071) );
  AND U2086 ( .A(n46), .B(n2134), .Z(n2133) );
  XNOR U2087 ( .A(n2135), .B(n2132), .Z(n2134) );
  XNOR U2088 ( .A(n2136), .B(n2137), .Z(n46) );
  AND U2089 ( .A(n2138), .B(n2139), .Z(n2137) );
  XOR U2090 ( .A(n2096), .B(n2136), .Z(n2139) );
  AND U2091 ( .A(n2140), .B(n2141), .Z(n2096) );
  XOR U2092 ( .A(n2136), .B(n2093), .Z(n2138) );
  XNOR U2093 ( .A(n2142), .B(n2143), .Z(n2093) );
  AND U2094 ( .A(n50), .B(n2099), .Z(n2143) );
  XOR U2095 ( .A(n2097), .B(n2142), .Z(n2099) );
  XOR U2096 ( .A(n2144), .B(n2145), .Z(n2136) );
  AND U2097 ( .A(n2146), .B(n2147), .Z(n2145) );
  XNOR U2098 ( .A(n2144), .B(n2140), .Z(n2147) );
  IV U2099 ( .A(n2107), .Z(n2140) );
  XOR U2100 ( .A(n2148), .B(n2149), .Z(n2107) );
  XOR U2101 ( .A(n2150), .B(n2141), .Z(n2149) );
  AND U2102 ( .A(n2116), .B(n2151), .Z(n2141) );
  AND U2103 ( .A(n2152), .B(n2153), .Z(n2150) );
  XOR U2104 ( .A(n2154), .B(n2148), .Z(n2152) );
  XNOR U2105 ( .A(n2104), .B(n2144), .Z(n2146) );
  XNOR U2106 ( .A(n2155), .B(n2156), .Z(n2104) );
  AND U2107 ( .A(n50), .B(n2110), .Z(n2156) );
  XOR U2108 ( .A(n2155), .B(n2108), .Z(n2110) );
  XOR U2109 ( .A(n2157), .B(n2158), .Z(n2144) );
  AND U2110 ( .A(n2159), .B(n2160), .Z(n2158) );
  XNOR U2111 ( .A(n2157), .B(n2116), .Z(n2160) );
  XOR U2112 ( .A(n2161), .B(n2153), .Z(n2116) );
  XNOR U2113 ( .A(n2162), .B(n2148), .Z(n2153) );
  XOR U2114 ( .A(n2163), .B(n2164), .Z(n2148) );
  AND U2115 ( .A(n2165), .B(n2166), .Z(n2164) );
  XOR U2116 ( .A(n2167), .B(n2163), .Z(n2165) );
  XNOR U2117 ( .A(n2168), .B(n2169), .Z(n2162) );
  AND U2118 ( .A(n2170), .B(n2171), .Z(n2169) );
  XOR U2119 ( .A(n2168), .B(n2172), .Z(n2170) );
  XNOR U2120 ( .A(n2154), .B(n2151), .Z(n2161) );
  AND U2121 ( .A(n2173), .B(n2174), .Z(n2151) );
  XOR U2122 ( .A(n2175), .B(n2176), .Z(n2154) );
  AND U2123 ( .A(n2177), .B(n2178), .Z(n2176) );
  XOR U2124 ( .A(n2175), .B(n2179), .Z(n2177) );
  XNOR U2125 ( .A(n2113), .B(n2157), .Z(n2159) );
  XNOR U2126 ( .A(n2180), .B(n2181), .Z(n2113) );
  AND U2127 ( .A(n50), .B(n2119), .Z(n2181) );
  XOR U2128 ( .A(n2180), .B(n2117), .Z(n2119) );
  XOR U2129 ( .A(n2182), .B(n2183), .Z(n2157) );
  AND U2130 ( .A(n2184), .B(n2185), .Z(n2183) );
  XNOR U2131 ( .A(n2182), .B(n2173), .Z(n2185) );
  IV U2132 ( .A(n2127), .Z(n2173) );
  XNOR U2133 ( .A(n2186), .B(n2166), .Z(n2127) );
  XNOR U2134 ( .A(n2187), .B(n2172), .Z(n2166) );
  XOR U2135 ( .A(n2188), .B(n2189), .Z(n2172) );
  NOR U2136 ( .A(n2190), .B(n2191), .Z(n2189) );
  XNOR U2137 ( .A(n2188), .B(n2192), .Z(n2190) );
  XNOR U2138 ( .A(n2171), .B(n2163), .Z(n2187) );
  XOR U2139 ( .A(n2193), .B(n2194), .Z(n2163) );
  AND U2140 ( .A(n2195), .B(n2196), .Z(n2194) );
  XOR U2141 ( .A(n2193), .B(n2197), .Z(n2195) );
  XNOR U2142 ( .A(n2198), .B(n2168), .Z(n2171) );
  XOR U2143 ( .A(n2199), .B(n2200), .Z(n2168) );
  AND U2144 ( .A(n2201), .B(n2202), .Z(n2200) );
  XNOR U2145 ( .A(n2203), .B(n2204), .Z(n2201) );
  IV U2146 ( .A(n2199), .Z(n2203) );
  XNOR U2147 ( .A(n2205), .B(n2206), .Z(n2198) );
  NOR U2148 ( .A(n2207), .B(n2208), .Z(n2206) );
  XOR U2149 ( .A(n2205), .B(n2209), .Z(n2207) );
  XNOR U2150 ( .A(n2167), .B(n2174), .Z(n2186) );
  NOR U2151 ( .A(n2135), .B(n2210), .Z(n2174) );
  XOR U2152 ( .A(n2179), .B(n2178), .Z(n2167) );
  XNOR U2153 ( .A(n2211), .B(n2175), .Z(n2178) );
  XOR U2154 ( .A(n2212), .B(n2213), .Z(n2175) );
  AND U2155 ( .A(n2214), .B(n2215), .Z(n2213) );
  XNOR U2156 ( .A(n2216), .B(n2217), .Z(n2214) );
  IV U2157 ( .A(n2212), .Z(n2216) );
  XNOR U2158 ( .A(n2218), .B(n2219), .Z(n2211) );
  NOR U2159 ( .A(n2220), .B(n2221), .Z(n2219) );
  XNOR U2160 ( .A(n2218), .B(n2222), .Z(n2220) );
  XOR U2161 ( .A(n2223), .B(n2224), .Z(n2179) );
  NOR U2162 ( .A(n2225), .B(n2226), .Z(n2224) );
  XNOR U2163 ( .A(n2223), .B(n2227), .Z(n2225) );
  XNOR U2164 ( .A(n2124), .B(n2182), .Z(n2184) );
  XNOR U2165 ( .A(n2228), .B(n2229), .Z(n2124) );
  AND U2166 ( .A(n50), .B(n2131), .Z(n2229) );
  XOR U2167 ( .A(n2228), .B(n2129), .Z(n2131) );
  AND U2168 ( .A(n2132), .B(n2135), .Z(n2182) );
  XOR U2169 ( .A(n2230), .B(n2210), .Z(n2135) );
  XNOR U2170 ( .A(p_input[16]), .B(p_input[256]), .Z(n2210) );
  XNOR U2171 ( .A(n2197), .B(n2196), .Z(n2230) );
  XNOR U2172 ( .A(n2231), .B(n2204), .Z(n2196) );
  XNOR U2173 ( .A(n2192), .B(n2191), .Z(n2204) );
  XOR U2174 ( .A(n2232), .B(n2188), .Z(n2191) );
  XNOR U2175 ( .A(n2233), .B(p_input[26]), .Z(n2188) );
  XNOR U2176 ( .A(p_input[267]), .B(p_input[27]), .Z(n2232) );
  XOR U2177 ( .A(p_input[268]), .B(p_input[28]), .Z(n2192) );
  XOR U2178 ( .A(n2202), .B(n2234), .Z(n2231) );
  IV U2179 ( .A(n2193), .Z(n2234) );
  XOR U2180 ( .A(p_input[17]), .B(p_input[257]), .Z(n2193) );
  XOR U2181 ( .A(n2235), .B(n2209), .Z(n2202) );
  XNOR U2182 ( .A(p_input[271]), .B(p_input[31]), .Z(n2209) );
  XOR U2183 ( .A(n2199), .B(n2208), .Z(n2235) );
  XOR U2184 ( .A(n2236), .B(n2205), .Z(n2208) );
  XOR U2185 ( .A(p_input[269]), .B(p_input[29]), .Z(n2205) );
  XNOR U2186 ( .A(p_input[270]), .B(p_input[30]), .Z(n2236) );
  XOR U2187 ( .A(p_input[25]), .B(p_input[265]), .Z(n2199) );
  XOR U2188 ( .A(n2217), .B(n2215), .Z(n2197) );
  XNOR U2189 ( .A(n2237), .B(n2222), .Z(n2215) );
  XOR U2190 ( .A(p_input[24]), .B(p_input[264]), .Z(n2222) );
  XOR U2191 ( .A(n2212), .B(n2221), .Z(n2237) );
  XOR U2192 ( .A(n2238), .B(n2218), .Z(n2221) );
  XOR U2193 ( .A(p_input[22]), .B(p_input[262]), .Z(n2218) );
  XOR U2194 ( .A(p_input[23]), .B(n2239), .Z(n2238) );
  XOR U2195 ( .A(p_input[18]), .B(p_input[258]), .Z(n2212) );
  XNOR U2196 ( .A(n2227), .B(n2226), .Z(n2217) );
  XOR U2197 ( .A(n2240), .B(n2223), .Z(n2226) );
  XOR U2198 ( .A(p_input[19]), .B(p_input[259]), .Z(n2223) );
  XOR U2199 ( .A(p_input[20]), .B(n2241), .Z(n2240) );
  XOR U2200 ( .A(p_input[21]), .B(p_input[261]), .Z(n2227) );
  XNOR U2201 ( .A(n2242), .B(n2243), .Z(n2132) );
  AND U2202 ( .A(n50), .B(n2244), .Z(n2243) );
  XNOR U2203 ( .A(n2245), .B(n2246), .Z(n50) );
  AND U2204 ( .A(n2247), .B(n2248), .Z(n2246) );
  XOR U2205 ( .A(n2245), .B(n2142), .Z(n2248) );
  XNOR U2206 ( .A(n2245), .B(n2097), .Z(n2247) );
  XOR U2207 ( .A(n2249), .B(n2250), .Z(n2245) );
  AND U2208 ( .A(n2251), .B(n2252), .Z(n2250) );
  XOR U2209 ( .A(n2249), .B(n2108), .Z(n2251) );
  XOR U2210 ( .A(n2253), .B(n2254), .Z(n2086) );
  AND U2211 ( .A(n54), .B(n2244), .Z(n2254) );
  XNOR U2212 ( .A(n2242), .B(n2253), .Z(n2244) );
  XNOR U2213 ( .A(n2255), .B(n2256), .Z(n54) );
  AND U2214 ( .A(n2257), .B(n2258), .Z(n2256) );
  XNOR U2215 ( .A(n2259), .B(n2255), .Z(n2258) );
  IV U2216 ( .A(n2142), .Z(n2259) );
  XNOR U2217 ( .A(n2260), .B(n2261), .Z(n2142) );
  AND U2218 ( .A(n57), .B(n2262), .Z(n2261) );
  XNOR U2219 ( .A(n2260), .B(n2263), .Z(n2262) );
  XNOR U2220 ( .A(n2097), .B(n2255), .Z(n2257) );
  XOR U2221 ( .A(n2264), .B(n2265), .Z(n2097) );
  AND U2222 ( .A(n65), .B(n2266), .Z(n2265) );
  XOR U2223 ( .A(n2249), .B(n2267), .Z(n2255) );
  AND U2224 ( .A(n2268), .B(n2252), .Z(n2267) );
  XNOR U2225 ( .A(n2155), .B(n2249), .Z(n2252) );
  XNOR U2226 ( .A(n2269), .B(n2270), .Z(n2155) );
  AND U2227 ( .A(n57), .B(n2271), .Z(n2270) );
  XOR U2228 ( .A(n2272), .B(n2269), .Z(n2271) );
  XNOR U2229 ( .A(n2273), .B(n2249), .Z(n2268) );
  IV U2230 ( .A(n2108), .Z(n2273) );
  XOR U2231 ( .A(n2274), .B(n2275), .Z(n2108) );
  AND U2232 ( .A(n65), .B(n2276), .Z(n2275) );
  XOR U2233 ( .A(n2277), .B(n2278), .Z(n2249) );
  AND U2234 ( .A(n2279), .B(n2280), .Z(n2278) );
  XNOR U2235 ( .A(n2180), .B(n2277), .Z(n2280) );
  XNOR U2236 ( .A(n2281), .B(n2282), .Z(n2180) );
  AND U2237 ( .A(n57), .B(n2283), .Z(n2282) );
  XNOR U2238 ( .A(n2284), .B(n2281), .Z(n2283) );
  XOR U2239 ( .A(n2277), .B(n2117), .Z(n2279) );
  XOR U2240 ( .A(n2285), .B(n2286), .Z(n2117) );
  AND U2241 ( .A(n65), .B(n2287), .Z(n2286) );
  XOR U2242 ( .A(n2288), .B(n2289), .Z(n2277) );
  AND U2243 ( .A(n2290), .B(n2291), .Z(n2289) );
  XNOR U2244 ( .A(n2288), .B(n2228), .Z(n2291) );
  XNOR U2245 ( .A(n2292), .B(n2293), .Z(n2228) );
  AND U2246 ( .A(n57), .B(n2294), .Z(n2293) );
  XOR U2247 ( .A(n2295), .B(n2292), .Z(n2294) );
  XNOR U2248 ( .A(n2296), .B(n2288), .Z(n2290) );
  IV U2249 ( .A(n2129), .Z(n2296) );
  XOR U2250 ( .A(n2297), .B(n2298), .Z(n2129) );
  AND U2251 ( .A(n65), .B(n2299), .Z(n2298) );
  AND U2252 ( .A(n2253), .B(n2242), .Z(n2288) );
  XNOR U2253 ( .A(n2300), .B(n2301), .Z(n2242) );
  AND U2254 ( .A(n57), .B(n2302), .Z(n2301) );
  XNOR U2255 ( .A(n2303), .B(n2300), .Z(n2302) );
  XNOR U2256 ( .A(n2304), .B(n2305), .Z(n57) );
  AND U2257 ( .A(n2306), .B(n2307), .Z(n2305) );
  XOR U2258 ( .A(n2263), .B(n2304), .Z(n2307) );
  AND U2259 ( .A(n2308), .B(n2309), .Z(n2263) );
  XOR U2260 ( .A(n2304), .B(n2260), .Z(n2306) );
  XNOR U2261 ( .A(n2310), .B(n2311), .Z(n2260) );
  AND U2262 ( .A(n61), .B(n2266), .Z(n2311) );
  XOR U2263 ( .A(n2264), .B(n2310), .Z(n2266) );
  XOR U2264 ( .A(n2312), .B(n2313), .Z(n2304) );
  AND U2265 ( .A(n2314), .B(n2315), .Z(n2313) );
  XNOR U2266 ( .A(n2312), .B(n2308), .Z(n2315) );
  IV U2267 ( .A(n2272), .Z(n2308) );
  XOR U2268 ( .A(n2316), .B(n2317), .Z(n2272) );
  XOR U2269 ( .A(n2318), .B(n2309), .Z(n2317) );
  AND U2270 ( .A(n2284), .B(n2319), .Z(n2309) );
  AND U2271 ( .A(n2320), .B(n2321), .Z(n2318) );
  XOR U2272 ( .A(n2322), .B(n2316), .Z(n2320) );
  XNOR U2273 ( .A(n2269), .B(n2312), .Z(n2314) );
  XNOR U2274 ( .A(n2323), .B(n2324), .Z(n2269) );
  AND U2275 ( .A(n61), .B(n2276), .Z(n2324) );
  XOR U2276 ( .A(n2323), .B(n2274), .Z(n2276) );
  XOR U2277 ( .A(n2325), .B(n2326), .Z(n2312) );
  AND U2278 ( .A(n2327), .B(n2328), .Z(n2326) );
  XNOR U2279 ( .A(n2325), .B(n2284), .Z(n2328) );
  XOR U2280 ( .A(n2329), .B(n2321), .Z(n2284) );
  XNOR U2281 ( .A(n2330), .B(n2316), .Z(n2321) );
  XOR U2282 ( .A(n2331), .B(n2332), .Z(n2316) );
  AND U2283 ( .A(n2333), .B(n2334), .Z(n2332) );
  XOR U2284 ( .A(n2335), .B(n2331), .Z(n2333) );
  XNOR U2285 ( .A(n2336), .B(n2337), .Z(n2330) );
  AND U2286 ( .A(n2338), .B(n2339), .Z(n2337) );
  XOR U2287 ( .A(n2336), .B(n2340), .Z(n2338) );
  XNOR U2288 ( .A(n2322), .B(n2319), .Z(n2329) );
  AND U2289 ( .A(n2341), .B(n2342), .Z(n2319) );
  XOR U2290 ( .A(n2343), .B(n2344), .Z(n2322) );
  AND U2291 ( .A(n2345), .B(n2346), .Z(n2344) );
  XOR U2292 ( .A(n2343), .B(n2347), .Z(n2345) );
  XNOR U2293 ( .A(n2281), .B(n2325), .Z(n2327) );
  XNOR U2294 ( .A(n2348), .B(n2349), .Z(n2281) );
  AND U2295 ( .A(n61), .B(n2287), .Z(n2349) );
  XOR U2296 ( .A(n2348), .B(n2285), .Z(n2287) );
  XOR U2297 ( .A(n2350), .B(n2351), .Z(n2325) );
  AND U2298 ( .A(n2352), .B(n2353), .Z(n2351) );
  XNOR U2299 ( .A(n2350), .B(n2341), .Z(n2353) );
  IV U2300 ( .A(n2295), .Z(n2341) );
  XNOR U2301 ( .A(n2354), .B(n2334), .Z(n2295) );
  XNOR U2302 ( .A(n2355), .B(n2340), .Z(n2334) );
  XOR U2303 ( .A(n2356), .B(n2357), .Z(n2340) );
  NOR U2304 ( .A(n2358), .B(n2359), .Z(n2357) );
  XNOR U2305 ( .A(n2356), .B(n2360), .Z(n2358) );
  XNOR U2306 ( .A(n2339), .B(n2331), .Z(n2355) );
  XOR U2307 ( .A(n2361), .B(n2362), .Z(n2331) );
  AND U2308 ( .A(n2363), .B(n2364), .Z(n2362) );
  XNOR U2309 ( .A(n2361), .B(n2365), .Z(n2363) );
  XNOR U2310 ( .A(n2366), .B(n2336), .Z(n2339) );
  XOR U2311 ( .A(n2367), .B(n2368), .Z(n2336) );
  AND U2312 ( .A(n2369), .B(n2370), .Z(n2368) );
  XOR U2313 ( .A(n2367), .B(n2371), .Z(n2369) );
  XNOR U2314 ( .A(n2372), .B(n2373), .Z(n2366) );
  NOR U2315 ( .A(n2374), .B(n2375), .Z(n2373) );
  XOR U2316 ( .A(n2372), .B(n2376), .Z(n2374) );
  XNOR U2317 ( .A(n2335), .B(n2342), .Z(n2354) );
  NOR U2318 ( .A(n2303), .B(n2377), .Z(n2342) );
  XOR U2319 ( .A(n2347), .B(n2346), .Z(n2335) );
  XNOR U2320 ( .A(n2378), .B(n2343), .Z(n2346) );
  XOR U2321 ( .A(n2379), .B(n2380), .Z(n2343) );
  AND U2322 ( .A(n2381), .B(n2382), .Z(n2380) );
  XOR U2323 ( .A(n2379), .B(n2383), .Z(n2381) );
  XNOR U2324 ( .A(n2384), .B(n2385), .Z(n2378) );
  NOR U2325 ( .A(n2386), .B(n2387), .Z(n2385) );
  XNOR U2326 ( .A(n2384), .B(n2388), .Z(n2386) );
  XOR U2327 ( .A(n2389), .B(n2390), .Z(n2347) );
  NOR U2328 ( .A(n2391), .B(n2392), .Z(n2390) );
  XNOR U2329 ( .A(n2389), .B(n2393), .Z(n2391) );
  XNOR U2330 ( .A(n2292), .B(n2350), .Z(n2352) );
  XNOR U2331 ( .A(n2394), .B(n2395), .Z(n2292) );
  AND U2332 ( .A(n61), .B(n2299), .Z(n2395) );
  XOR U2333 ( .A(n2394), .B(n2297), .Z(n2299) );
  AND U2334 ( .A(n2300), .B(n2303), .Z(n2350) );
  XOR U2335 ( .A(n2396), .B(n2377), .Z(n2303) );
  XNOR U2336 ( .A(p_input[256]), .B(p_input[32]), .Z(n2377) );
  XOR U2337 ( .A(n2365), .B(n2364), .Z(n2396) );
  XNOR U2338 ( .A(n2397), .B(n2371), .Z(n2364) );
  XNOR U2339 ( .A(n2360), .B(n2359), .Z(n2371) );
  XOR U2340 ( .A(n2398), .B(n2356), .Z(n2359) );
  XNOR U2341 ( .A(n2233), .B(p_input[42]), .Z(n2356) );
  XNOR U2342 ( .A(p_input[267]), .B(p_input[43]), .Z(n2398) );
  XOR U2343 ( .A(p_input[268]), .B(p_input[44]), .Z(n2360) );
  XNOR U2344 ( .A(n2370), .B(n2361), .Z(n2397) );
  XNOR U2345 ( .A(n2399), .B(p_input[33]), .Z(n2361) );
  XOR U2346 ( .A(n2400), .B(n2376), .Z(n2370) );
  XNOR U2347 ( .A(p_input[271]), .B(p_input[47]), .Z(n2376) );
  XOR U2348 ( .A(n2367), .B(n2375), .Z(n2400) );
  XOR U2349 ( .A(n2401), .B(n2372), .Z(n2375) );
  XOR U2350 ( .A(p_input[269]), .B(p_input[45]), .Z(n2372) );
  XNOR U2351 ( .A(p_input[270]), .B(p_input[46]), .Z(n2401) );
  XNOR U2352 ( .A(n2066), .B(p_input[41]), .Z(n2367) );
  XNOR U2353 ( .A(n2383), .B(n2382), .Z(n2365) );
  XNOR U2354 ( .A(n2402), .B(n2388), .Z(n2382) );
  XOR U2355 ( .A(p_input[264]), .B(p_input[40]), .Z(n2388) );
  XOR U2356 ( .A(n2379), .B(n2387), .Z(n2402) );
  XOR U2357 ( .A(n2403), .B(n2384), .Z(n2387) );
  XOR U2358 ( .A(p_input[262]), .B(p_input[38]), .Z(n2384) );
  XNOR U2359 ( .A(p_input[263]), .B(p_input[39]), .Z(n2403) );
  XNOR U2360 ( .A(n2069), .B(p_input[34]), .Z(n2379) );
  XNOR U2361 ( .A(n2393), .B(n2392), .Z(n2383) );
  XOR U2362 ( .A(n2404), .B(n2389), .Z(n2392) );
  XOR U2363 ( .A(p_input[259]), .B(p_input[35]), .Z(n2389) );
  XNOR U2364 ( .A(p_input[260]), .B(p_input[36]), .Z(n2404) );
  XOR U2365 ( .A(p_input[261]), .B(p_input[37]), .Z(n2393) );
  XNOR U2366 ( .A(n2405), .B(n2406), .Z(n2300) );
  AND U2367 ( .A(n61), .B(n2407), .Z(n2406) );
  XNOR U2368 ( .A(n2408), .B(n2409), .Z(n61) );
  AND U2369 ( .A(n2410), .B(n2411), .Z(n2409) );
  XOR U2370 ( .A(n2408), .B(n2310), .Z(n2411) );
  XNOR U2371 ( .A(n2408), .B(n2264), .Z(n2410) );
  XOR U2372 ( .A(n2412), .B(n2413), .Z(n2408) );
  AND U2373 ( .A(n2414), .B(n2415), .Z(n2413) );
  XOR U2374 ( .A(n2412), .B(n2274), .Z(n2414) );
  XOR U2375 ( .A(n2416), .B(n2417), .Z(n2253) );
  AND U2376 ( .A(n65), .B(n2407), .Z(n2417) );
  XNOR U2377 ( .A(n2405), .B(n2416), .Z(n2407) );
  XNOR U2378 ( .A(n2418), .B(n2419), .Z(n65) );
  AND U2379 ( .A(n2420), .B(n2421), .Z(n2419) );
  XNOR U2380 ( .A(n2422), .B(n2418), .Z(n2421) );
  IV U2381 ( .A(n2310), .Z(n2422) );
  XNOR U2382 ( .A(n2423), .B(n2424), .Z(n2310) );
  AND U2383 ( .A(n68), .B(n2425), .Z(n2424) );
  XNOR U2384 ( .A(n2423), .B(n2426), .Z(n2425) );
  XNOR U2385 ( .A(n2264), .B(n2418), .Z(n2420) );
  XOR U2386 ( .A(n2427), .B(n2428), .Z(n2264) );
  AND U2387 ( .A(n76), .B(n2429), .Z(n2428) );
  XOR U2388 ( .A(n2412), .B(n2430), .Z(n2418) );
  AND U2389 ( .A(n2431), .B(n2415), .Z(n2430) );
  XNOR U2390 ( .A(n2323), .B(n2412), .Z(n2415) );
  XNOR U2391 ( .A(n2432), .B(n2433), .Z(n2323) );
  AND U2392 ( .A(n68), .B(n2434), .Z(n2433) );
  XOR U2393 ( .A(n2435), .B(n2432), .Z(n2434) );
  XNOR U2394 ( .A(n2436), .B(n2412), .Z(n2431) );
  IV U2395 ( .A(n2274), .Z(n2436) );
  XOR U2396 ( .A(n2437), .B(n2438), .Z(n2274) );
  AND U2397 ( .A(n76), .B(n2439), .Z(n2438) );
  XOR U2398 ( .A(n2440), .B(n2441), .Z(n2412) );
  AND U2399 ( .A(n2442), .B(n2443), .Z(n2441) );
  XNOR U2400 ( .A(n2348), .B(n2440), .Z(n2443) );
  XNOR U2401 ( .A(n2444), .B(n2445), .Z(n2348) );
  AND U2402 ( .A(n68), .B(n2446), .Z(n2445) );
  XNOR U2403 ( .A(n2447), .B(n2444), .Z(n2446) );
  XOR U2404 ( .A(n2440), .B(n2285), .Z(n2442) );
  XOR U2405 ( .A(n2448), .B(n2449), .Z(n2285) );
  AND U2406 ( .A(n76), .B(n2450), .Z(n2449) );
  XOR U2407 ( .A(n2451), .B(n2452), .Z(n2440) );
  AND U2408 ( .A(n2453), .B(n2454), .Z(n2452) );
  XNOR U2409 ( .A(n2451), .B(n2394), .Z(n2454) );
  XNOR U2410 ( .A(n2455), .B(n2456), .Z(n2394) );
  AND U2411 ( .A(n68), .B(n2457), .Z(n2456) );
  XOR U2412 ( .A(n2458), .B(n2455), .Z(n2457) );
  XNOR U2413 ( .A(n2459), .B(n2451), .Z(n2453) );
  IV U2414 ( .A(n2297), .Z(n2459) );
  XOR U2415 ( .A(n2460), .B(n2461), .Z(n2297) );
  AND U2416 ( .A(n76), .B(n2462), .Z(n2461) );
  AND U2417 ( .A(n2416), .B(n2405), .Z(n2451) );
  XNOR U2418 ( .A(n2463), .B(n2464), .Z(n2405) );
  AND U2419 ( .A(n68), .B(n2465), .Z(n2464) );
  XNOR U2420 ( .A(n2466), .B(n2463), .Z(n2465) );
  XNOR U2421 ( .A(n2467), .B(n2468), .Z(n68) );
  AND U2422 ( .A(n2469), .B(n2470), .Z(n2468) );
  XOR U2423 ( .A(n2426), .B(n2467), .Z(n2470) );
  AND U2424 ( .A(n2471), .B(n2472), .Z(n2426) );
  XOR U2425 ( .A(n2467), .B(n2423), .Z(n2469) );
  XNOR U2426 ( .A(n2473), .B(n2474), .Z(n2423) );
  AND U2427 ( .A(n72), .B(n2429), .Z(n2474) );
  XOR U2428 ( .A(n2427), .B(n2473), .Z(n2429) );
  XOR U2429 ( .A(n2475), .B(n2476), .Z(n2467) );
  AND U2430 ( .A(n2477), .B(n2478), .Z(n2476) );
  XNOR U2431 ( .A(n2475), .B(n2471), .Z(n2478) );
  IV U2432 ( .A(n2435), .Z(n2471) );
  XOR U2433 ( .A(n2479), .B(n2480), .Z(n2435) );
  XOR U2434 ( .A(n2481), .B(n2472), .Z(n2480) );
  AND U2435 ( .A(n2447), .B(n2482), .Z(n2472) );
  AND U2436 ( .A(n2483), .B(n2484), .Z(n2481) );
  XOR U2437 ( .A(n2485), .B(n2479), .Z(n2483) );
  XNOR U2438 ( .A(n2432), .B(n2475), .Z(n2477) );
  XNOR U2439 ( .A(n2486), .B(n2487), .Z(n2432) );
  AND U2440 ( .A(n72), .B(n2439), .Z(n2487) );
  XOR U2441 ( .A(n2486), .B(n2437), .Z(n2439) );
  XOR U2442 ( .A(n2488), .B(n2489), .Z(n2475) );
  AND U2443 ( .A(n2490), .B(n2491), .Z(n2489) );
  XNOR U2444 ( .A(n2488), .B(n2447), .Z(n2491) );
  XOR U2445 ( .A(n2492), .B(n2484), .Z(n2447) );
  XNOR U2446 ( .A(n2493), .B(n2479), .Z(n2484) );
  XOR U2447 ( .A(n2494), .B(n2495), .Z(n2479) );
  AND U2448 ( .A(n2496), .B(n2497), .Z(n2495) );
  XOR U2449 ( .A(n2498), .B(n2494), .Z(n2496) );
  XNOR U2450 ( .A(n2499), .B(n2500), .Z(n2493) );
  AND U2451 ( .A(n2501), .B(n2502), .Z(n2500) );
  XOR U2452 ( .A(n2499), .B(n2503), .Z(n2501) );
  XNOR U2453 ( .A(n2485), .B(n2482), .Z(n2492) );
  AND U2454 ( .A(n2504), .B(n2505), .Z(n2482) );
  XOR U2455 ( .A(n2506), .B(n2507), .Z(n2485) );
  AND U2456 ( .A(n2508), .B(n2509), .Z(n2507) );
  XOR U2457 ( .A(n2506), .B(n2510), .Z(n2508) );
  XNOR U2458 ( .A(n2444), .B(n2488), .Z(n2490) );
  XNOR U2459 ( .A(n2511), .B(n2512), .Z(n2444) );
  AND U2460 ( .A(n72), .B(n2450), .Z(n2512) );
  XOR U2461 ( .A(n2511), .B(n2448), .Z(n2450) );
  XOR U2462 ( .A(n2513), .B(n2514), .Z(n2488) );
  AND U2463 ( .A(n2515), .B(n2516), .Z(n2514) );
  XNOR U2464 ( .A(n2513), .B(n2504), .Z(n2516) );
  IV U2465 ( .A(n2458), .Z(n2504) );
  XNOR U2466 ( .A(n2517), .B(n2497), .Z(n2458) );
  XNOR U2467 ( .A(n2518), .B(n2503), .Z(n2497) );
  XOR U2468 ( .A(n2519), .B(n2520), .Z(n2503) );
  NOR U2469 ( .A(n2521), .B(n2522), .Z(n2520) );
  XNOR U2470 ( .A(n2519), .B(n2523), .Z(n2521) );
  XNOR U2471 ( .A(n2502), .B(n2494), .Z(n2518) );
  XOR U2472 ( .A(n2524), .B(n2525), .Z(n2494) );
  AND U2473 ( .A(n2526), .B(n2527), .Z(n2525) );
  XNOR U2474 ( .A(n2524), .B(n2528), .Z(n2526) );
  XNOR U2475 ( .A(n2529), .B(n2499), .Z(n2502) );
  XOR U2476 ( .A(n2530), .B(n2531), .Z(n2499) );
  AND U2477 ( .A(n2532), .B(n2533), .Z(n2531) );
  XOR U2478 ( .A(n2530), .B(n2534), .Z(n2532) );
  XNOR U2479 ( .A(n2535), .B(n2536), .Z(n2529) );
  NOR U2480 ( .A(n2537), .B(n2538), .Z(n2536) );
  XOR U2481 ( .A(n2535), .B(n2539), .Z(n2537) );
  XNOR U2482 ( .A(n2498), .B(n2505), .Z(n2517) );
  NOR U2483 ( .A(n2466), .B(n2540), .Z(n2505) );
  XOR U2484 ( .A(n2510), .B(n2509), .Z(n2498) );
  XNOR U2485 ( .A(n2541), .B(n2506), .Z(n2509) );
  XOR U2486 ( .A(n2542), .B(n2543), .Z(n2506) );
  AND U2487 ( .A(n2544), .B(n2545), .Z(n2543) );
  XOR U2488 ( .A(n2542), .B(n2546), .Z(n2544) );
  XNOR U2489 ( .A(n2547), .B(n2548), .Z(n2541) );
  NOR U2490 ( .A(n2549), .B(n2550), .Z(n2548) );
  XNOR U2491 ( .A(n2547), .B(n2551), .Z(n2549) );
  XOR U2492 ( .A(n2552), .B(n2553), .Z(n2510) );
  NOR U2493 ( .A(n2554), .B(n2555), .Z(n2553) );
  XNOR U2494 ( .A(n2552), .B(n2556), .Z(n2554) );
  XNOR U2495 ( .A(n2455), .B(n2513), .Z(n2515) );
  XNOR U2496 ( .A(n2557), .B(n2558), .Z(n2455) );
  AND U2497 ( .A(n72), .B(n2462), .Z(n2558) );
  XOR U2498 ( .A(n2557), .B(n2460), .Z(n2462) );
  AND U2499 ( .A(n2463), .B(n2466), .Z(n2513) );
  XOR U2500 ( .A(n2559), .B(n2540), .Z(n2466) );
  XNOR U2501 ( .A(p_input[256]), .B(p_input[48]), .Z(n2540) );
  XOR U2502 ( .A(n2528), .B(n2527), .Z(n2559) );
  XNOR U2503 ( .A(n2560), .B(n2534), .Z(n2527) );
  XNOR U2504 ( .A(n2523), .B(n2522), .Z(n2534) );
  XOR U2505 ( .A(n2561), .B(n2519), .Z(n2522) );
  XNOR U2506 ( .A(n2233), .B(p_input[58]), .Z(n2519) );
  XNOR U2507 ( .A(p_input[267]), .B(p_input[59]), .Z(n2561) );
  XOR U2508 ( .A(p_input[268]), .B(p_input[60]), .Z(n2523) );
  XNOR U2509 ( .A(n2533), .B(n2524), .Z(n2560) );
  XNOR U2510 ( .A(n2399), .B(p_input[49]), .Z(n2524) );
  XOR U2511 ( .A(n2562), .B(n2539), .Z(n2533) );
  XNOR U2512 ( .A(p_input[271]), .B(p_input[63]), .Z(n2539) );
  XOR U2513 ( .A(n2530), .B(n2538), .Z(n2562) );
  XOR U2514 ( .A(n2563), .B(n2535), .Z(n2538) );
  XOR U2515 ( .A(p_input[269]), .B(p_input[61]), .Z(n2535) );
  XNOR U2516 ( .A(p_input[270]), .B(p_input[62]), .Z(n2563) );
  XNOR U2517 ( .A(n2066), .B(p_input[57]), .Z(n2530) );
  XNOR U2518 ( .A(n2546), .B(n2545), .Z(n2528) );
  XNOR U2519 ( .A(n2564), .B(n2551), .Z(n2545) );
  XOR U2520 ( .A(p_input[264]), .B(p_input[56]), .Z(n2551) );
  XOR U2521 ( .A(n2542), .B(n2550), .Z(n2564) );
  XOR U2522 ( .A(n2565), .B(n2547), .Z(n2550) );
  XOR U2523 ( .A(p_input[262]), .B(p_input[54]), .Z(n2547) );
  XNOR U2524 ( .A(p_input[263]), .B(p_input[55]), .Z(n2565) );
  XNOR U2525 ( .A(n2069), .B(p_input[50]), .Z(n2542) );
  XNOR U2526 ( .A(n2556), .B(n2555), .Z(n2546) );
  XOR U2527 ( .A(n2566), .B(n2552), .Z(n2555) );
  XOR U2528 ( .A(p_input[259]), .B(p_input[51]), .Z(n2552) );
  XNOR U2529 ( .A(p_input[260]), .B(p_input[52]), .Z(n2566) );
  XOR U2530 ( .A(p_input[261]), .B(p_input[53]), .Z(n2556) );
  XNOR U2531 ( .A(n2567), .B(n2568), .Z(n2463) );
  AND U2532 ( .A(n72), .B(n2569), .Z(n2568) );
  XNOR U2533 ( .A(n2570), .B(n2571), .Z(n72) );
  AND U2534 ( .A(n2572), .B(n2573), .Z(n2571) );
  XOR U2535 ( .A(n2570), .B(n2473), .Z(n2573) );
  XNOR U2536 ( .A(n2570), .B(n2427), .Z(n2572) );
  XOR U2537 ( .A(n2574), .B(n2575), .Z(n2570) );
  AND U2538 ( .A(n2576), .B(n2577), .Z(n2575) );
  XOR U2539 ( .A(n2574), .B(n2437), .Z(n2576) );
  XOR U2540 ( .A(n2578), .B(n2579), .Z(n2416) );
  AND U2541 ( .A(n76), .B(n2569), .Z(n2579) );
  XNOR U2542 ( .A(n2567), .B(n2578), .Z(n2569) );
  XNOR U2543 ( .A(n2580), .B(n2581), .Z(n76) );
  AND U2544 ( .A(n2582), .B(n2583), .Z(n2581) );
  XNOR U2545 ( .A(n2584), .B(n2580), .Z(n2583) );
  IV U2546 ( .A(n2473), .Z(n2584) );
  XNOR U2547 ( .A(n2585), .B(n2586), .Z(n2473) );
  AND U2548 ( .A(n79), .B(n2587), .Z(n2586) );
  XNOR U2549 ( .A(n2585), .B(n2588), .Z(n2587) );
  XNOR U2550 ( .A(n2427), .B(n2580), .Z(n2582) );
  XOR U2551 ( .A(n2589), .B(n2590), .Z(n2427) );
  AND U2552 ( .A(n87), .B(n2591), .Z(n2590) );
  XOR U2553 ( .A(n2574), .B(n2592), .Z(n2580) );
  AND U2554 ( .A(n2593), .B(n2577), .Z(n2592) );
  XNOR U2555 ( .A(n2486), .B(n2574), .Z(n2577) );
  XNOR U2556 ( .A(n2594), .B(n2595), .Z(n2486) );
  AND U2557 ( .A(n79), .B(n2596), .Z(n2595) );
  XOR U2558 ( .A(n2597), .B(n2594), .Z(n2596) );
  XNOR U2559 ( .A(n2598), .B(n2574), .Z(n2593) );
  IV U2560 ( .A(n2437), .Z(n2598) );
  XOR U2561 ( .A(n2599), .B(n2600), .Z(n2437) );
  AND U2562 ( .A(n87), .B(n2601), .Z(n2600) );
  XOR U2563 ( .A(n2602), .B(n2603), .Z(n2574) );
  AND U2564 ( .A(n2604), .B(n2605), .Z(n2603) );
  XNOR U2565 ( .A(n2511), .B(n2602), .Z(n2605) );
  XNOR U2566 ( .A(n2606), .B(n2607), .Z(n2511) );
  AND U2567 ( .A(n79), .B(n2608), .Z(n2607) );
  XNOR U2568 ( .A(n2609), .B(n2606), .Z(n2608) );
  XOR U2569 ( .A(n2602), .B(n2448), .Z(n2604) );
  XOR U2570 ( .A(n2610), .B(n2611), .Z(n2448) );
  AND U2571 ( .A(n87), .B(n2612), .Z(n2611) );
  XOR U2572 ( .A(n2613), .B(n2614), .Z(n2602) );
  AND U2573 ( .A(n2615), .B(n2616), .Z(n2614) );
  XNOR U2574 ( .A(n2613), .B(n2557), .Z(n2616) );
  XNOR U2575 ( .A(n2617), .B(n2618), .Z(n2557) );
  AND U2576 ( .A(n79), .B(n2619), .Z(n2618) );
  XOR U2577 ( .A(n2620), .B(n2617), .Z(n2619) );
  XNOR U2578 ( .A(n2621), .B(n2613), .Z(n2615) );
  IV U2579 ( .A(n2460), .Z(n2621) );
  XOR U2580 ( .A(n2622), .B(n2623), .Z(n2460) );
  AND U2581 ( .A(n87), .B(n2624), .Z(n2623) );
  AND U2582 ( .A(n2578), .B(n2567), .Z(n2613) );
  XNOR U2583 ( .A(n2625), .B(n2626), .Z(n2567) );
  AND U2584 ( .A(n79), .B(n2627), .Z(n2626) );
  XNOR U2585 ( .A(n2628), .B(n2625), .Z(n2627) );
  XNOR U2586 ( .A(n2629), .B(n2630), .Z(n79) );
  AND U2587 ( .A(n2631), .B(n2632), .Z(n2630) );
  XOR U2588 ( .A(n2588), .B(n2629), .Z(n2632) );
  AND U2589 ( .A(n2633), .B(n2634), .Z(n2588) );
  XOR U2590 ( .A(n2629), .B(n2585), .Z(n2631) );
  XNOR U2591 ( .A(n2635), .B(n2636), .Z(n2585) );
  AND U2592 ( .A(n83), .B(n2591), .Z(n2636) );
  XOR U2593 ( .A(n2589), .B(n2635), .Z(n2591) );
  XOR U2594 ( .A(n2637), .B(n2638), .Z(n2629) );
  AND U2595 ( .A(n2639), .B(n2640), .Z(n2638) );
  XNOR U2596 ( .A(n2637), .B(n2633), .Z(n2640) );
  IV U2597 ( .A(n2597), .Z(n2633) );
  XOR U2598 ( .A(n2641), .B(n2642), .Z(n2597) );
  XOR U2599 ( .A(n2643), .B(n2634), .Z(n2642) );
  AND U2600 ( .A(n2609), .B(n2644), .Z(n2634) );
  AND U2601 ( .A(n2645), .B(n2646), .Z(n2643) );
  XOR U2602 ( .A(n2647), .B(n2641), .Z(n2645) );
  XNOR U2603 ( .A(n2594), .B(n2637), .Z(n2639) );
  XNOR U2604 ( .A(n2648), .B(n2649), .Z(n2594) );
  AND U2605 ( .A(n83), .B(n2601), .Z(n2649) );
  XOR U2606 ( .A(n2648), .B(n2599), .Z(n2601) );
  XOR U2607 ( .A(n2650), .B(n2651), .Z(n2637) );
  AND U2608 ( .A(n2652), .B(n2653), .Z(n2651) );
  XNOR U2609 ( .A(n2650), .B(n2609), .Z(n2653) );
  XOR U2610 ( .A(n2654), .B(n2646), .Z(n2609) );
  XNOR U2611 ( .A(n2655), .B(n2641), .Z(n2646) );
  XOR U2612 ( .A(n2656), .B(n2657), .Z(n2641) );
  AND U2613 ( .A(n2658), .B(n2659), .Z(n2657) );
  XOR U2614 ( .A(n2660), .B(n2656), .Z(n2658) );
  XNOR U2615 ( .A(n2661), .B(n2662), .Z(n2655) );
  AND U2616 ( .A(n2663), .B(n2664), .Z(n2662) );
  XOR U2617 ( .A(n2661), .B(n2665), .Z(n2663) );
  XNOR U2618 ( .A(n2647), .B(n2644), .Z(n2654) );
  AND U2619 ( .A(n2666), .B(n2667), .Z(n2644) );
  XOR U2620 ( .A(n2668), .B(n2669), .Z(n2647) );
  AND U2621 ( .A(n2670), .B(n2671), .Z(n2669) );
  XOR U2622 ( .A(n2668), .B(n2672), .Z(n2670) );
  XNOR U2623 ( .A(n2606), .B(n2650), .Z(n2652) );
  XNOR U2624 ( .A(n2673), .B(n2674), .Z(n2606) );
  AND U2625 ( .A(n83), .B(n2612), .Z(n2674) );
  XOR U2626 ( .A(n2673), .B(n2610), .Z(n2612) );
  XOR U2627 ( .A(n2675), .B(n2676), .Z(n2650) );
  AND U2628 ( .A(n2677), .B(n2678), .Z(n2676) );
  XNOR U2629 ( .A(n2675), .B(n2666), .Z(n2678) );
  IV U2630 ( .A(n2620), .Z(n2666) );
  XNOR U2631 ( .A(n2679), .B(n2659), .Z(n2620) );
  XNOR U2632 ( .A(n2680), .B(n2665), .Z(n2659) );
  XOR U2633 ( .A(n2681), .B(n2682), .Z(n2665) );
  NOR U2634 ( .A(n2683), .B(n2684), .Z(n2682) );
  XNOR U2635 ( .A(n2681), .B(n2685), .Z(n2683) );
  XNOR U2636 ( .A(n2664), .B(n2656), .Z(n2680) );
  XOR U2637 ( .A(n2686), .B(n2687), .Z(n2656) );
  AND U2638 ( .A(n2688), .B(n2689), .Z(n2687) );
  XNOR U2639 ( .A(n2686), .B(n2690), .Z(n2688) );
  XNOR U2640 ( .A(n2691), .B(n2661), .Z(n2664) );
  XOR U2641 ( .A(n2692), .B(n2693), .Z(n2661) );
  AND U2642 ( .A(n2694), .B(n2695), .Z(n2693) );
  XOR U2643 ( .A(n2692), .B(n2696), .Z(n2694) );
  XNOR U2644 ( .A(n2697), .B(n2698), .Z(n2691) );
  NOR U2645 ( .A(n2699), .B(n2700), .Z(n2698) );
  XOR U2646 ( .A(n2697), .B(n2701), .Z(n2699) );
  XNOR U2647 ( .A(n2660), .B(n2667), .Z(n2679) );
  NOR U2648 ( .A(n2628), .B(n2702), .Z(n2667) );
  XOR U2649 ( .A(n2672), .B(n2671), .Z(n2660) );
  XNOR U2650 ( .A(n2703), .B(n2668), .Z(n2671) );
  XOR U2651 ( .A(n2704), .B(n2705), .Z(n2668) );
  AND U2652 ( .A(n2706), .B(n2707), .Z(n2705) );
  XOR U2653 ( .A(n2704), .B(n2708), .Z(n2706) );
  XNOR U2654 ( .A(n2709), .B(n2710), .Z(n2703) );
  NOR U2655 ( .A(n2711), .B(n2712), .Z(n2710) );
  XNOR U2656 ( .A(n2709), .B(n2713), .Z(n2711) );
  XOR U2657 ( .A(n2714), .B(n2715), .Z(n2672) );
  NOR U2658 ( .A(n2716), .B(n2717), .Z(n2715) );
  XNOR U2659 ( .A(n2714), .B(n2718), .Z(n2716) );
  XNOR U2660 ( .A(n2617), .B(n2675), .Z(n2677) );
  XNOR U2661 ( .A(n2719), .B(n2720), .Z(n2617) );
  AND U2662 ( .A(n83), .B(n2624), .Z(n2720) );
  XOR U2663 ( .A(n2719), .B(n2622), .Z(n2624) );
  AND U2664 ( .A(n2625), .B(n2628), .Z(n2675) );
  XOR U2665 ( .A(n2721), .B(n2702), .Z(n2628) );
  XNOR U2666 ( .A(p_input[256]), .B(p_input[64]), .Z(n2702) );
  XOR U2667 ( .A(n2690), .B(n2689), .Z(n2721) );
  XNOR U2668 ( .A(n2722), .B(n2696), .Z(n2689) );
  XNOR U2669 ( .A(n2685), .B(n2684), .Z(n2696) );
  XOR U2670 ( .A(n2723), .B(n2681), .Z(n2684) );
  XNOR U2671 ( .A(n2233), .B(p_input[74]), .Z(n2681) );
  XNOR U2672 ( .A(p_input[267]), .B(p_input[75]), .Z(n2723) );
  XOR U2673 ( .A(p_input[268]), .B(p_input[76]), .Z(n2685) );
  XNOR U2674 ( .A(n2695), .B(n2686), .Z(n2722) );
  XNOR U2675 ( .A(n2399), .B(p_input[65]), .Z(n2686) );
  XOR U2676 ( .A(n2724), .B(n2701), .Z(n2695) );
  XNOR U2677 ( .A(p_input[271]), .B(p_input[79]), .Z(n2701) );
  XOR U2678 ( .A(n2692), .B(n2700), .Z(n2724) );
  XOR U2679 ( .A(n2725), .B(n2697), .Z(n2700) );
  XOR U2680 ( .A(p_input[269]), .B(p_input[77]), .Z(n2697) );
  XNOR U2681 ( .A(p_input[270]), .B(p_input[78]), .Z(n2725) );
  XNOR U2682 ( .A(n2066), .B(p_input[73]), .Z(n2692) );
  XNOR U2683 ( .A(n2708), .B(n2707), .Z(n2690) );
  XNOR U2684 ( .A(n2726), .B(n2713), .Z(n2707) );
  XOR U2685 ( .A(p_input[264]), .B(p_input[72]), .Z(n2713) );
  XOR U2686 ( .A(n2704), .B(n2712), .Z(n2726) );
  XOR U2687 ( .A(n2727), .B(n2709), .Z(n2712) );
  XOR U2688 ( .A(p_input[262]), .B(p_input[70]), .Z(n2709) );
  XNOR U2689 ( .A(p_input[263]), .B(p_input[71]), .Z(n2727) );
  XNOR U2690 ( .A(n2069), .B(p_input[66]), .Z(n2704) );
  XNOR U2691 ( .A(n2718), .B(n2717), .Z(n2708) );
  XOR U2692 ( .A(n2728), .B(n2714), .Z(n2717) );
  XOR U2693 ( .A(p_input[259]), .B(p_input[67]), .Z(n2714) );
  XNOR U2694 ( .A(p_input[260]), .B(p_input[68]), .Z(n2728) );
  XOR U2695 ( .A(p_input[261]), .B(p_input[69]), .Z(n2718) );
  XNOR U2696 ( .A(n2729), .B(n2730), .Z(n2625) );
  AND U2697 ( .A(n83), .B(n2731), .Z(n2730) );
  XNOR U2698 ( .A(n2732), .B(n2733), .Z(n83) );
  AND U2699 ( .A(n2734), .B(n2735), .Z(n2733) );
  XOR U2700 ( .A(n2732), .B(n2635), .Z(n2735) );
  XNOR U2701 ( .A(n2732), .B(n2589), .Z(n2734) );
  XOR U2702 ( .A(n2736), .B(n2737), .Z(n2732) );
  AND U2703 ( .A(n2738), .B(n2739), .Z(n2737) );
  XOR U2704 ( .A(n2736), .B(n2599), .Z(n2738) );
  XOR U2705 ( .A(n2740), .B(n2741), .Z(n2578) );
  AND U2706 ( .A(n87), .B(n2731), .Z(n2741) );
  XNOR U2707 ( .A(n2729), .B(n2740), .Z(n2731) );
  XNOR U2708 ( .A(n2742), .B(n2743), .Z(n87) );
  AND U2709 ( .A(n2744), .B(n2745), .Z(n2743) );
  XNOR U2710 ( .A(n2746), .B(n2742), .Z(n2745) );
  IV U2711 ( .A(n2635), .Z(n2746) );
  XNOR U2712 ( .A(n2747), .B(n2748), .Z(n2635) );
  AND U2713 ( .A(n90), .B(n2749), .Z(n2748) );
  XNOR U2714 ( .A(n2747), .B(n2750), .Z(n2749) );
  XNOR U2715 ( .A(n2589), .B(n2742), .Z(n2744) );
  XOR U2716 ( .A(n2751), .B(n2752), .Z(n2589) );
  AND U2717 ( .A(n98), .B(n2753), .Z(n2752) );
  XOR U2718 ( .A(n2736), .B(n2754), .Z(n2742) );
  AND U2719 ( .A(n2755), .B(n2739), .Z(n2754) );
  XNOR U2720 ( .A(n2648), .B(n2736), .Z(n2739) );
  XNOR U2721 ( .A(n2756), .B(n2757), .Z(n2648) );
  AND U2722 ( .A(n90), .B(n2758), .Z(n2757) );
  XOR U2723 ( .A(n2759), .B(n2756), .Z(n2758) );
  XNOR U2724 ( .A(n2760), .B(n2736), .Z(n2755) );
  IV U2725 ( .A(n2599), .Z(n2760) );
  XOR U2726 ( .A(n2761), .B(n2762), .Z(n2599) );
  AND U2727 ( .A(n98), .B(n2763), .Z(n2762) );
  XOR U2728 ( .A(n2764), .B(n2765), .Z(n2736) );
  AND U2729 ( .A(n2766), .B(n2767), .Z(n2765) );
  XNOR U2730 ( .A(n2673), .B(n2764), .Z(n2767) );
  XNOR U2731 ( .A(n2768), .B(n2769), .Z(n2673) );
  AND U2732 ( .A(n90), .B(n2770), .Z(n2769) );
  XNOR U2733 ( .A(n2771), .B(n2768), .Z(n2770) );
  XOR U2734 ( .A(n2764), .B(n2610), .Z(n2766) );
  XOR U2735 ( .A(n2772), .B(n2773), .Z(n2610) );
  AND U2736 ( .A(n98), .B(n2774), .Z(n2773) );
  XOR U2737 ( .A(n2775), .B(n2776), .Z(n2764) );
  AND U2738 ( .A(n2777), .B(n2778), .Z(n2776) );
  XNOR U2739 ( .A(n2775), .B(n2719), .Z(n2778) );
  XNOR U2740 ( .A(n2779), .B(n2780), .Z(n2719) );
  AND U2741 ( .A(n90), .B(n2781), .Z(n2780) );
  XOR U2742 ( .A(n2782), .B(n2779), .Z(n2781) );
  XNOR U2743 ( .A(n2783), .B(n2775), .Z(n2777) );
  IV U2744 ( .A(n2622), .Z(n2783) );
  XOR U2745 ( .A(n2784), .B(n2785), .Z(n2622) );
  AND U2746 ( .A(n98), .B(n2786), .Z(n2785) );
  AND U2747 ( .A(n2740), .B(n2729), .Z(n2775) );
  XNOR U2748 ( .A(n2787), .B(n2788), .Z(n2729) );
  AND U2749 ( .A(n90), .B(n2789), .Z(n2788) );
  XNOR U2750 ( .A(n2790), .B(n2787), .Z(n2789) );
  XNOR U2751 ( .A(n2791), .B(n2792), .Z(n90) );
  AND U2752 ( .A(n2793), .B(n2794), .Z(n2792) );
  XOR U2753 ( .A(n2750), .B(n2791), .Z(n2794) );
  AND U2754 ( .A(n2795), .B(n2796), .Z(n2750) );
  XOR U2755 ( .A(n2791), .B(n2747), .Z(n2793) );
  XNOR U2756 ( .A(n2797), .B(n2798), .Z(n2747) );
  AND U2757 ( .A(n94), .B(n2753), .Z(n2798) );
  XOR U2758 ( .A(n2751), .B(n2797), .Z(n2753) );
  XOR U2759 ( .A(n2799), .B(n2800), .Z(n2791) );
  AND U2760 ( .A(n2801), .B(n2802), .Z(n2800) );
  XNOR U2761 ( .A(n2799), .B(n2795), .Z(n2802) );
  IV U2762 ( .A(n2759), .Z(n2795) );
  XOR U2763 ( .A(n2803), .B(n2804), .Z(n2759) );
  XOR U2764 ( .A(n2805), .B(n2796), .Z(n2804) );
  AND U2765 ( .A(n2771), .B(n2806), .Z(n2796) );
  AND U2766 ( .A(n2807), .B(n2808), .Z(n2805) );
  XOR U2767 ( .A(n2809), .B(n2803), .Z(n2807) );
  XNOR U2768 ( .A(n2756), .B(n2799), .Z(n2801) );
  XNOR U2769 ( .A(n2810), .B(n2811), .Z(n2756) );
  AND U2770 ( .A(n94), .B(n2763), .Z(n2811) );
  XOR U2771 ( .A(n2810), .B(n2761), .Z(n2763) );
  XOR U2772 ( .A(n2812), .B(n2813), .Z(n2799) );
  AND U2773 ( .A(n2814), .B(n2815), .Z(n2813) );
  XNOR U2774 ( .A(n2812), .B(n2771), .Z(n2815) );
  XOR U2775 ( .A(n2816), .B(n2808), .Z(n2771) );
  XNOR U2776 ( .A(n2817), .B(n2803), .Z(n2808) );
  XOR U2777 ( .A(n2818), .B(n2819), .Z(n2803) );
  AND U2778 ( .A(n2820), .B(n2821), .Z(n2819) );
  XOR U2779 ( .A(n2822), .B(n2818), .Z(n2820) );
  XNOR U2780 ( .A(n2823), .B(n2824), .Z(n2817) );
  AND U2781 ( .A(n2825), .B(n2826), .Z(n2824) );
  XOR U2782 ( .A(n2823), .B(n2827), .Z(n2825) );
  XNOR U2783 ( .A(n2809), .B(n2806), .Z(n2816) );
  AND U2784 ( .A(n2828), .B(n2829), .Z(n2806) );
  XOR U2785 ( .A(n2830), .B(n2831), .Z(n2809) );
  AND U2786 ( .A(n2832), .B(n2833), .Z(n2831) );
  XOR U2787 ( .A(n2830), .B(n2834), .Z(n2832) );
  XNOR U2788 ( .A(n2768), .B(n2812), .Z(n2814) );
  XNOR U2789 ( .A(n2835), .B(n2836), .Z(n2768) );
  AND U2790 ( .A(n94), .B(n2774), .Z(n2836) );
  XOR U2791 ( .A(n2835), .B(n2772), .Z(n2774) );
  XOR U2792 ( .A(n2837), .B(n2838), .Z(n2812) );
  AND U2793 ( .A(n2839), .B(n2840), .Z(n2838) );
  XNOR U2794 ( .A(n2837), .B(n2828), .Z(n2840) );
  IV U2795 ( .A(n2782), .Z(n2828) );
  XNOR U2796 ( .A(n2841), .B(n2821), .Z(n2782) );
  XNOR U2797 ( .A(n2842), .B(n2827), .Z(n2821) );
  XOR U2798 ( .A(n2843), .B(n2844), .Z(n2827) );
  NOR U2799 ( .A(n2845), .B(n2846), .Z(n2844) );
  XNOR U2800 ( .A(n2843), .B(n2847), .Z(n2845) );
  XNOR U2801 ( .A(n2826), .B(n2818), .Z(n2842) );
  XOR U2802 ( .A(n2848), .B(n2849), .Z(n2818) );
  AND U2803 ( .A(n2850), .B(n2851), .Z(n2849) );
  XNOR U2804 ( .A(n2848), .B(n2852), .Z(n2850) );
  XNOR U2805 ( .A(n2853), .B(n2823), .Z(n2826) );
  XOR U2806 ( .A(n2854), .B(n2855), .Z(n2823) );
  AND U2807 ( .A(n2856), .B(n2857), .Z(n2855) );
  XOR U2808 ( .A(n2854), .B(n2858), .Z(n2856) );
  XNOR U2809 ( .A(n2859), .B(n2860), .Z(n2853) );
  NOR U2810 ( .A(n2861), .B(n2862), .Z(n2860) );
  XOR U2811 ( .A(n2859), .B(n2863), .Z(n2861) );
  XNOR U2812 ( .A(n2822), .B(n2829), .Z(n2841) );
  NOR U2813 ( .A(n2790), .B(n2864), .Z(n2829) );
  XOR U2814 ( .A(n2834), .B(n2833), .Z(n2822) );
  XNOR U2815 ( .A(n2865), .B(n2830), .Z(n2833) );
  XOR U2816 ( .A(n2866), .B(n2867), .Z(n2830) );
  AND U2817 ( .A(n2868), .B(n2869), .Z(n2867) );
  XOR U2818 ( .A(n2866), .B(n2870), .Z(n2868) );
  XNOR U2819 ( .A(n2871), .B(n2872), .Z(n2865) );
  NOR U2820 ( .A(n2873), .B(n2874), .Z(n2872) );
  XNOR U2821 ( .A(n2871), .B(n2875), .Z(n2873) );
  XOR U2822 ( .A(n2876), .B(n2877), .Z(n2834) );
  NOR U2823 ( .A(n2878), .B(n2879), .Z(n2877) );
  XNOR U2824 ( .A(n2876), .B(n2880), .Z(n2878) );
  XNOR U2825 ( .A(n2779), .B(n2837), .Z(n2839) );
  XNOR U2826 ( .A(n2881), .B(n2882), .Z(n2779) );
  AND U2827 ( .A(n94), .B(n2786), .Z(n2882) );
  XOR U2828 ( .A(n2881), .B(n2784), .Z(n2786) );
  AND U2829 ( .A(n2787), .B(n2790), .Z(n2837) );
  XOR U2830 ( .A(n2883), .B(n2864), .Z(n2790) );
  XNOR U2831 ( .A(p_input[256]), .B(p_input[80]), .Z(n2864) );
  XOR U2832 ( .A(n2852), .B(n2851), .Z(n2883) );
  XNOR U2833 ( .A(n2884), .B(n2858), .Z(n2851) );
  XNOR U2834 ( .A(n2847), .B(n2846), .Z(n2858) );
  XOR U2835 ( .A(n2885), .B(n2843), .Z(n2846) );
  XNOR U2836 ( .A(n2233), .B(p_input[90]), .Z(n2843) );
  XNOR U2837 ( .A(p_input[267]), .B(p_input[91]), .Z(n2885) );
  XOR U2838 ( .A(p_input[268]), .B(p_input[92]), .Z(n2847) );
  XNOR U2839 ( .A(n2857), .B(n2848), .Z(n2884) );
  XNOR U2840 ( .A(n2399), .B(p_input[81]), .Z(n2848) );
  XOR U2841 ( .A(n2886), .B(n2863), .Z(n2857) );
  XNOR U2842 ( .A(p_input[271]), .B(p_input[95]), .Z(n2863) );
  XOR U2843 ( .A(n2854), .B(n2862), .Z(n2886) );
  XOR U2844 ( .A(n2887), .B(n2859), .Z(n2862) );
  XOR U2845 ( .A(p_input[269]), .B(p_input[93]), .Z(n2859) );
  XNOR U2846 ( .A(p_input[270]), .B(p_input[94]), .Z(n2887) );
  XNOR U2847 ( .A(n2066), .B(p_input[89]), .Z(n2854) );
  IV U2848 ( .A(p_input[265]), .Z(n2066) );
  XNOR U2849 ( .A(n2870), .B(n2869), .Z(n2852) );
  XNOR U2850 ( .A(n2888), .B(n2875), .Z(n2869) );
  XOR U2851 ( .A(p_input[264]), .B(p_input[88]), .Z(n2875) );
  XOR U2852 ( .A(n2866), .B(n2874), .Z(n2888) );
  XOR U2853 ( .A(n2889), .B(n2871), .Z(n2874) );
  XOR U2854 ( .A(p_input[262]), .B(p_input[86]), .Z(n2871) );
  XNOR U2855 ( .A(p_input[263]), .B(p_input[87]), .Z(n2889) );
  XNOR U2856 ( .A(n2069), .B(p_input[82]), .Z(n2866) );
  XNOR U2857 ( .A(n2880), .B(n2879), .Z(n2870) );
  XOR U2858 ( .A(n2890), .B(n2876), .Z(n2879) );
  XOR U2859 ( .A(p_input[259]), .B(p_input[83]), .Z(n2876) );
  XNOR U2860 ( .A(p_input[260]), .B(p_input[84]), .Z(n2890) );
  XOR U2861 ( .A(p_input[261]), .B(p_input[85]), .Z(n2880) );
  XNOR U2862 ( .A(n2891), .B(n2892), .Z(n2787) );
  AND U2863 ( .A(n94), .B(n2893), .Z(n2892) );
  XNOR U2864 ( .A(n2894), .B(n2895), .Z(n94) );
  AND U2865 ( .A(n2896), .B(n2897), .Z(n2895) );
  XOR U2866 ( .A(n2894), .B(n2797), .Z(n2897) );
  XNOR U2867 ( .A(n2894), .B(n2751), .Z(n2896) );
  XOR U2868 ( .A(n2898), .B(n2899), .Z(n2894) );
  AND U2869 ( .A(n2900), .B(n2901), .Z(n2899) );
  XOR U2870 ( .A(n2898), .B(n2761), .Z(n2900) );
  XOR U2871 ( .A(n2902), .B(n2903), .Z(n2740) );
  AND U2872 ( .A(n98), .B(n2893), .Z(n2903) );
  XNOR U2873 ( .A(n2891), .B(n2902), .Z(n2893) );
  XNOR U2874 ( .A(n2904), .B(n2905), .Z(n98) );
  AND U2875 ( .A(n2906), .B(n2907), .Z(n2905) );
  XNOR U2876 ( .A(n2908), .B(n2904), .Z(n2907) );
  IV U2877 ( .A(n2797), .Z(n2908) );
  XNOR U2878 ( .A(n2909), .B(n2910), .Z(n2797) );
  AND U2879 ( .A(n101), .B(n2911), .Z(n2910) );
  XNOR U2880 ( .A(n2909), .B(n2912), .Z(n2911) );
  XNOR U2881 ( .A(n2751), .B(n2904), .Z(n2906) );
  XOR U2882 ( .A(n2913), .B(n2914), .Z(n2751) );
  AND U2883 ( .A(n109), .B(n2915), .Z(n2914) );
  XOR U2884 ( .A(n2898), .B(n2916), .Z(n2904) );
  AND U2885 ( .A(n2917), .B(n2901), .Z(n2916) );
  XNOR U2886 ( .A(n2810), .B(n2898), .Z(n2901) );
  XNOR U2887 ( .A(n2918), .B(n2919), .Z(n2810) );
  AND U2888 ( .A(n101), .B(n2920), .Z(n2919) );
  XOR U2889 ( .A(n2921), .B(n2918), .Z(n2920) );
  XNOR U2890 ( .A(n2922), .B(n2898), .Z(n2917) );
  IV U2891 ( .A(n2761), .Z(n2922) );
  XOR U2892 ( .A(n2923), .B(n2924), .Z(n2761) );
  AND U2893 ( .A(n109), .B(n2925), .Z(n2924) );
  XOR U2894 ( .A(n2926), .B(n2927), .Z(n2898) );
  AND U2895 ( .A(n2928), .B(n2929), .Z(n2927) );
  XNOR U2896 ( .A(n2835), .B(n2926), .Z(n2929) );
  XNOR U2897 ( .A(n2930), .B(n2931), .Z(n2835) );
  AND U2898 ( .A(n101), .B(n2932), .Z(n2931) );
  XNOR U2899 ( .A(n2933), .B(n2930), .Z(n2932) );
  XOR U2900 ( .A(n2926), .B(n2772), .Z(n2928) );
  XOR U2901 ( .A(n2934), .B(n2935), .Z(n2772) );
  AND U2902 ( .A(n109), .B(n2936), .Z(n2935) );
  XOR U2903 ( .A(n2937), .B(n2938), .Z(n2926) );
  AND U2904 ( .A(n2939), .B(n2940), .Z(n2938) );
  XNOR U2905 ( .A(n2937), .B(n2881), .Z(n2940) );
  XNOR U2906 ( .A(n2941), .B(n2942), .Z(n2881) );
  AND U2907 ( .A(n101), .B(n2943), .Z(n2942) );
  XOR U2908 ( .A(n2944), .B(n2941), .Z(n2943) );
  XNOR U2909 ( .A(n2945), .B(n2937), .Z(n2939) );
  IV U2910 ( .A(n2784), .Z(n2945) );
  XOR U2911 ( .A(n2946), .B(n2947), .Z(n2784) );
  AND U2912 ( .A(n109), .B(n2948), .Z(n2947) );
  AND U2913 ( .A(n2902), .B(n2891), .Z(n2937) );
  XNOR U2914 ( .A(n2949), .B(n2950), .Z(n2891) );
  AND U2915 ( .A(n101), .B(n2951), .Z(n2950) );
  XNOR U2916 ( .A(n2952), .B(n2949), .Z(n2951) );
  XNOR U2917 ( .A(n2953), .B(n2954), .Z(n101) );
  AND U2918 ( .A(n2955), .B(n2956), .Z(n2954) );
  XOR U2919 ( .A(n2912), .B(n2953), .Z(n2956) );
  AND U2920 ( .A(n2957), .B(n2958), .Z(n2912) );
  XOR U2921 ( .A(n2953), .B(n2909), .Z(n2955) );
  XNOR U2922 ( .A(n2959), .B(n2960), .Z(n2909) );
  AND U2923 ( .A(n105), .B(n2915), .Z(n2960) );
  XOR U2924 ( .A(n2913), .B(n2959), .Z(n2915) );
  XOR U2925 ( .A(n2961), .B(n2962), .Z(n2953) );
  AND U2926 ( .A(n2963), .B(n2964), .Z(n2962) );
  XNOR U2927 ( .A(n2961), .B(n2957), .Z(n2964) );
  IV U2928 ( .A(n2921), .Z(n2957) );
  XOR U2929 ( .A(n2965), .B(n2966), .Z(n2921) );
  XOR U2930 ( .A(n2967), .B(n2958), .Z(n2966) );
  AND U2931 ( .A(n2933), .B(n2968), .Z(n2958) );
  AND U2932 ( .A(n2969), .B(n2970), .Z(n2967) );
  XOR U2933 ( .A(n2971), .B(n2965), .Z(n2969) );
  XNOR U2934 ( .A(n2918), .B(n2961), .Z(n2963) );
  XNOR U2935 ( .A(n2972), .B(n2973), .Z(n2918) );
  AND U2936 ( .A(n105), .B(n2925), .Z(n2973) );
  XOR U2937 ( .A(n2972), .B(n2923), .Z(n2925) );
  XOR U2938 ( .A(n2974), .B(n2975), .Z(n2961) );
  AND U2939 ( .A(n2976), .B(n2977), .Z(n2975) );
  XNOR U2940 ( .A(n2974), .B(n2933), .Z(n2977) );
  XOR U2941 ( .A(n2978), .B(n2970), .Z(n2933) );
  XNOR U2942 ( .A(n2979), .B(n2965), .Z(n2970) );
  XOR U2943 ( .A(n2980), .B(n2981), .Z(n2965) );
  AND U2944 ( .A(n2982), .B(n2983), .Z(n2981) );
  XOR U2945 ( .A(n2984), .B(n2980), .Z(n2982) );
  XNOR U2946 ( .A(n2985), .B(n2986), .Z(n2979) );
  AND U2947 ( .A(n2987), .B(n2988), .Z(n2986) );
  XOR U2948 ( .A(n2985), .B(n2989), .Z(n2987) );
  XNOR U2949 ( .A(n2971), .B(n2968), .Z(n2978) );
  AND U2950 ( .A(n2990), .B(n2991), .Z(n2968) );
  XOR U2951 ( .A(n2992), .B(n2993), .Z(n2971) );
  AND U2952 ( .A(n2994), .B(n2995), .Z(n2993) );
  XOR U2953 ( .A(n2992), .B(n2996), .Z(n2994) );
  XNOR U2954 ( .A(n2930), .B(n2974), .Z(n2976) );
  XNOR U2955 ( .A(n2997), .B(n2998), .Z(n2930) );
  AND U2956 ( .A(n105), .B(n2936), .Z(n2998) );
  XOR U2957 ( .A(n2997), .B(n2934), .Z(n2936) );
  XOR U2958 ( .A(n2999), .B(n3000), .Z(n2974) );
  AND U2959 ( .A(n3001), .B(n3002), .Z(n3000) );
  XNOR U2960 ( .A(n2999), .B(n2990), .Z(n3002) );
  IV U2961 ( .A(n2944), .Z(n2990) );
  XNOR U2962 ( .A(n3003), .B(n2983), .Z(n2944) );
  XNOR U2963 ( .A(n3004), .B(n2989), .Z(n2983) );
  XNOR U2964 ( .A(n3005), .B(n3006), .Z(n2989) );
  NOR U2965 ( .A(n3007), .B(n3008), .Z(n3006) );
  XOR U2966 ( .A(n3005), .B(n3009), .Z(n3007) );
  XNOR U2967 ( .A(n2988), .B(n2980), .Z(n3004) );
  XOR U2968 ( .A(n3010), .B(n3011), .Z(n2980) );
  AND U2969 ( .A(n3012), .B(n3013), .Z(n3011) );
  XOR U2970 ( .A(n3010), .B(n3014), .Z(n3012) );
  XNOR U2971 ( .A(n3015), .B(n2985), .Z(n2988) );
  XOR U2972 ( .A(n3016), .B(n3017), .Z(n2985) );
  AND U2973 ( .A(n3018), .B(n3019), .Z(n3017) );
  XNOR U2974 ( .A(n3020), .B(n3021), .Z(n3018) );
  IV U2975 ( .A(n3016), .Z(n3020) );
  XNOR U2976 ( .A(n3022), .B(n3023), .Z(n3015) );
  NOR U2977 ( .A(n3024), .B(n3025), .Z(n3023) );
  XNOR U2978 ( .A(n3022), .B(n3026), .Z(n3024) );
  XNOR U2979 ( .A(n2984), .B(n2991), .Z(n3003) );
  NOR U2980 ( .A(n2952), .B(n3027), .Z(n2991) );
  XOR U2981 ( .A(n2996), .B(n2995), .Z(n2984) );
  XNOR U2982 ( .A(n3028), .B(n2992), .Z(n2995) );
  XOR U2983 ( .A(n3029), .B(n3030), .Z(n2992) );
  AND U2984 ( .A(n3031), .B(n3032), .Z(n3030) );
  XOR U2985 ( .A(n3029), .B(n3033), .Z(n3031) );
  XNOR U2986 ( .A(n3034), .B(n3035), .Z(n3028) );
  NOR U2987 ( .A(n3036), .B(n3037), .Z(n3035) );
  XNOR U2988 ( .A(n3034), .B(n3038), .Z(n3036) );
  XOR U2989 ( .A(n3039), .B(n3040), .Z(n2996) );
  NOR U2990 ( .A(n3041), .B(n3042), .Z(n3040) );
  XNOR U2991 ( .A(n3039), .B(n3043), .Z(n3041) );
  XNOR U2992 ( .A(n2941), .B(n2999), .Z(n3001) );
  XNOR U2993 ( .A(n3044), .B(n3045), .Z(n2941) );
  AND U2994 ( .A(n105), .B(n2948), .Z(n3045) );
  XOR U2995 ( .A(n3044), .B(n2946), .Z(n2948) );
  AND U2996 ( .A(n2949), .B(n2952), .Z(n2999) );
  XOR U2997 ( .A(n3046), .B(n3027), .Z(n2952) );
  XNOR U2998 ( .A(p_input[256]), .B(p_input[96]), .Z(n3027) );
  XNOR U2999 ( .A(n3014), .B(n3013), .Z(n3046) );
  XNOR U3000 ( .A(n3047), .B(n3021), .Z(n3013) );
  XNOR U3001 ( .A(n3009), .B(n3008), .Z(n3021) );
  XNOR U3002 ( .A(n3048), .B(n3005), .Z(n3008) );
  XNOR U3003 ( .A(p_input[106]), .B(p_input[266]), .Z(n3005) );
  XOR U3004 ( .A(p_input[107]), .B(n2060), .Z(n3048) );
  XOR U3005 ( .A(p_input[108]), .B(p_input[268]), .Z(n3009) );
  XNOR U3006 ( .A(n3019), .B(n3010), .Z(n3047) );
  XNOR U3007 ( .A(n2399), .B(p_input[97]), .Z(n3010) );
  IV U3008 ( .A(p_input[257]), .Z(n2399) );
  XNOR U3009 ( .A(n3049), .B(n3026), .Z(n3019) );
  XNOR U3010 ( .A(p_input[111]), .B(n2063), .Z(n3026) );
  XOR U3011 ( .A(n3016), .B(n3025), .Z(n3049) );
  XOR U3012 ( .A(n3050), .B(n3022), .Z(n3025) );
  XOR U3013 ( .A(p_input[109]), .B(p_input[269]), .Z(n3022) );
  XOR U3014 ( .A(p_input[110]), .B(n2065), .Z(n3050) );
  XOR U3015 ( .A(p_input[105]), .B(p_input[265]), .Z(n3016) );
  XOR U3016 ( .A(n3033), .B(n3032), .Z(n3014) );
  XNOR U3017 ( .A(n3051), .B(n3038), .Z(n3032) );
  XOR U3018 ( .A(p_input[104]), .B(p_input[264]), .Z(n3038) );
  XOR U3019 ( .A(n3029), .B(n3037), .Z(n3051) );
  XOR U3020 ( .A(n3052), .B(n3034), .Z(n3037) );
  XOR U3021 ( .A(p_input[102]), .B(p_input[262]), .Z(n3034) );
  XOR U3022 ( .A(p_input[103]), .B(n2239), .Z(n3052) );
  XNOR U3023 ( .A(n2069), .B(p_input[98]), .Z(n3029) );
  IV U3024 ( .A(p_input[258]), .Z(n2069) );
  XNOR U3025 ( .A(n3043), .B(n3042), .Z(n3033) );
  XOR U3026 ( .A(n3053), .B(n3039), .Z(n3042) );
  XOR U3027 ( .A(p_input[259]), .B(p_input[99]), .Z(n3039) );
  XOR U3028 ( .A(p_input[100]), .B(n2241), .Z(n3053) );
  XOR U3029 ( .A(p_input[101]), .B(p_input[261]), .Z(n3043) );
  XNOR U3030 ( .A(n3054), .B(n3055), .Z(n2949) );
  AND U3031 ( .A(n105), .B(n3056), .Z(n3055) );
  XNOR U3032 ( .A(n3057), .B(n3058), .Z(n105) );
  AND U3033 ( .A(n3059), .B(n3060), .Z(n3058) );
  XOR U3034 ( .A(n3057), .B(n2959), .Z(n3060) );
  XNOR U3035 ( .A(n3057), .B(n2913), .Z(n3059) );
  XOR U3036 ( .A(n3061), .B(n3062), .Z(n3057) );
  AND U3037 ( .A(n3063), .B(n3064), .Z(n3062) );
  XOR U3038 ( .A(n3061), .B(n2923), .Z(n3063) );
  XOR U3039 ( .A(n3065), .B(n3066), .Z(n2902) );
  AND U3040 ( .A(n109), .B(n3056), .Z(n3066) );
  XNOR U3041 ( .A(n3054), .B(n3065), .Z(n3056) );
  XNOR U3042 ( .A(n3067), .B(n3068), .Z(n109) );
  AND U3043 ( .A(n3069), .B(n3070), .Z(n3068) );
  XNOR U3044 ( .A(n3071), .B(n3067), .Z(n3070) );
  IV U3045 ( .A(n2959), .Z(n3071) );
  XNOR U3046 ( .A(n3072), .B(n3073), .Z(n2959) );
  AND U3047 ( .A(n112), .B(n3074), .Z(n3073) );
  XNOR U3048 ( .A(n3072), .B(n3075), .Z(n3074) );
  XNOR U3049 ( .A(n2913), .B(n3067), .Z(n3069) );
  XOR U3050 ( .A(n3076), .B(n3077), .Z(n2913) );
  AND U3051 ( .A(n120), .B(n3078), .Z(n3077) );
  XOR U3052 ( .A(n3061), .B(n3079), .Z(n3067) );
  AND U3053 ( .A(n3080), .B(n3064), .Z(n3079) );
  XNOR U3054 ( .A(n2972), .B(n3061), .Z(n3064) );
  XNOR U3055 ( .A(n3081), .B(n3082), .Z(n2972) );
  AND U3056 ( .A(n112), .B(n3083), .Z(n3082) );
  XOR U3057 ( .A(n3084), .B(n3081), .Z(n3083) );
  XNOR U3058 ( .A(n3085), .B(n3061), .Z(n3080) );
  IV U3059 ( .A(n2923), .Z(n3085) );
  XOR U3060 ( .A(n3086), .B(n3087), .Z(n2923) );
  AND U3061 ( .A(n120), .B(n3088), .Z(n3087) );
  XOR U3062 ( .A(n3089), .B(n3090), .Z(n3061) );
  AND U3063 ( .A(n3091), .B(n3092), .Z(n3090) );
  XNOR U3064 ( .A(n2997), .B(n3089), .Z(n3092) );
  XNOR U3065 ( .A(n3093), .B(n3094), .Z(n2997) );
  AND U3066 ( .A(n112), .B(n3095), .Z(n3094) );
  XNOR U3067 ( .A(n3096), .B(n3093), .Z(n3095) );
  XOR U3068 ( .A(n3089), .B(n2934), .Z(n3091) );
  XOR U3069 ( .A(n3097), .B(n3098), .Z(n2934) );
  AND U3070 ( .A(n120), .B(n3099), .Z(n3098) );
  XOR U3071 ( .A(n3100), .B(n3101), .Z(n3089) );
  AND U3072 ( .A(n3102), .B(n3103), .Z(n3101) );
  XNOR U3073 ( .A(n3100), .B(n3044), .Z(n3103) );
  XNOR U3074 ( .A(n3104), .B(n3105), .Z(n3044) );
  AND U3075 ( .A(n112), .B(n3106), .Z(n3105) );
  XOR U3076 ( .A(n3107), .B(n3104), .Z(n3106) );
  XNOR U3077 ( .A(n3108), .B(n3100), .Z(n3102) );
  IV U3078 ( .A(n2946), .Z(n3108) );
  XOR U3079 ( .A(n3109), .B(n3110), .Z(n2946) );
  AND U3080 ( .A(n120), .B(n3111), .Z(n3110) );
  AND U3081 ( .A(n3065), .B(n3054), .Z(n3100) );
  XNOR U3082 ( .A(n3112), .B(n3113), .Z(n3054) );
  AND U3083 ( .A(n112), .B(n3114), .Z(n3113) );
  XNOR U3084 ( .A(n3115), .B(n3112), .Z(n3114) );
  XNOR U3085 ( .A(n3116), .B(n3117), .Z(n112) );
  AND U3086 ( .A(n3118), .B(n3119), .Z(n3117) );
  XOR U3087 ( .A(n3075), .B(n3116), .Z(n3119) );
  AND U3088 ( .A(n3120), .B(n3121), .Z(n3075) );
  XOR U3089 ( .A(n3116), .B(n3072), .Z(n3118) );
  XNOR U3090 ( .A(n3122), .B(n3123), .Z(n3072) );
  AND U3091 ( .A(n116), .B(n3078), .Z(n3123) );
  XOR U3092 ( .A(n3076), .B(n3122), .Z(n3078) );
  XOR U3093 ( .A(n3124), .B(n3125), .Z(n3116) );
  AND U3094 ( .A(n3126), .B(n3127), .Z(n3125) );
  XNOR U3095 ( .A(n3124), .B(n3120), .Z(n3127) );
  IV U3096 ( .A(n3084), .Z(n3120) );
  XOR U3097 ( .A(n3128), .B(n3129), .Z(n3084) );
  XOR U3098 ( .A(n3130), .B(n3121), .Z(n3129) );
  AND U3099 ( .A(n3096), .B(n3131), .Z(n3121) );
  AND U3100 ( .A(n3132), .B(n3133), .Z(n3130) );
  XOR U3101 ( .A(n3134), .B(n3128), .Z(n3132) );
  XNOR U3102 ( .A(n3081), .B(n3124), .Z(n3126) );
  XNOR U3103 ( .A(n3135), .B(n3136), .Z(n3081) );
  AND U3104 ( .A(n116), .B(n3088), .Z(n3136) );
  XOR U3105 ( .A(n3135), .B(n3086), .Z(n3088) );
  XOR U3106 ( .A(n3137), .B(n3138), .Z(n3124) );
  AND U3107 ( .A(n3139), .B(n3140), .Z(n3138) );
  XNOR U3108 ( .A(n3137), .B(n3096), .Z(n3140) );
  XOR U3109 ( .A(n3141), .B(n3133), .Z(n3096) );
  XNOR U3110 ( .A(n3142), .B(n3128), .Z(n3133) );
  XOR U3111 ( .A(n3143), .B(n3144), .Z(n3128) );
  AND U3112 ( .A(n3145), .B(n3146), .Z(n3144) );
  XOR U3113 ( .A(n3147), .B(n3143), .Z(n3145) );
  XNOR U3114 ( .A(n3148), .B(n3149), .Z(n3142) );
  AND U3115 ( .A(n3150), .B(n3151), .Z(n3149) );
  XOR U3116 ( .A(n3148), .B(n3152), .Z(n3150) );
  XNOR U3117 ( .A(n3134), .B(n3131), .Z(n3141) );
  AND U3118 ( .A(n3153), .B(n3154), .Z(n3131) );
  XOR U3119 ( .A(n3155), .B(n3156), .Z(n3134) );
  AND U3120 ( .A(n3157), .B(n3158), .Z(n3156) );
  XOR U3121 ( .A(n3155), .B(n3159), .Z(n3157) );
  XNOR U3122 ( .A(n3093), .B(n3137), .Z(n3139) );
  XNOR U3123 ( .A(n3160), .B(n3161), .Z(n3093) );
  AND U3124 ( .A(n116), .B(n3099), .Z(n3161) );
  XOR U3125 ( .A(n3160), .B(n3097), .Z(n3099) );
  XOR U3126 ( .A(n3162), .B(n3163), .Z(n3137) );
  AND U3127 ( .A(n3164), .B(n3165), .Z(n3163) );
  XNOR U3128 ( .A(n3162), .B(n3153), .Z(n3165) );
  IV U3129 ( .A(n3107), .Z(n3153) );
  XNOR U3130 ( .A(n3166), .B(n3146), .Z(n3107) );
  XNOR U3131 ( .A(n3167), .B(n3152), .Z(n3146) );
  XNOR U3132 ( .A(n3168), .B(n3169), .Z(n3152) );
  NOR U3133 ( .A(n3170), .B(n3171), .Z(n3169) );
  XOR U3134 ( .A(n3168), .B(n3172), .Z(n3170) );
  XNOR U3135 ( .A(n3151), .B(n3143), .Z(n3167) );
  XOR U3136 ( .A(n3173), .B(n3174), .Z(n3143) );
  AND U3137 ( .A(n3175), .B(n3176), .Z(n3174) );
  XOR U3138 ( .A(n3173), .B(n3177), .Z(n3175) );
  XNOR U3139 ( .A(n3178), .B(n3148), .Z(n3151) );
  XOR U3140 ( .A(n3179), .B(n3180), .Z(n3148) );
  AND U3141 ( .A(n3181), .B(n3182), .Z(n3180) );
  XNOR U3142 ( .A(n3183), .B(n3184), .Z(n3181) );
  IV U3143 ( .A(n3179), .Z(n3183) );
  XNOR U3144 ( .A(n3185), .B(n3186), .Z(n3178) );
  NOR U3145 ( .A(n3187), .B(n3188), .Z(n3186) );
  XNOR U3146 ( .A(n3185), .B(n3189), .Z(n3187) );
  XNOR U3147 ( .A(n3147), .B(n3154), .Z(n3166) );
  NOR U3148 ( .A(n3115), .B(n3190), .Z(n3154) );
  XOR U3149 ( .A(n3159), .B(n3158), .Z(n3147) );
  XNOR U3150 ( .A(n3191), .B(n3155), .Z(n3158) );
  XOR U3151 ( .A(n3192), .B(n3193), .Z(n3155) );
  AND U3152 ( .A(n3194), .B(n3195), .Z(n3193) );
  XNOR U3153 ( .A(n3196), .B(n3197), .Z(n3194) );
  IV U3154 ( .A(n3192), .Z(n3196) );
  XNOR U3155 ( .A(n3198), .B(n3199), .Z(n3191) );
  NOR U3156 ( .A(n3200), .B(n3201), .Z(n3199) );
  XNOR U3157 ( .A(n3198), .B(n3202), .Z(n3200) );
  XOR U3158 ( .A(n3203), .B(n3204), .Z(n3159) );
  NOR U3159 ( .A(n3205), .B(n3206), .Z(n3204) );
  XNOR U3160 ( .A(n3203), .B(n3207), .Z(n3205) );
  XNOR U3161 ( .A(n3104), .B(n3162), .Z(n3164) );
  XNOR U3162 ( .A(n3208), .B(n3209), .Z(n3104) );
  AND U3163 ( .A(n116), .B(n3111), .Z(n3209) );
  XOR U3164 ( .A(n3208), .B(n3109), .Z(n3111) );
  AND U3165 ( .A(n3112), .B(n3115), .Z(n3162) );
  XOR U3166 ( .A(n3210), .B(n3190), .Z(n3115) );
  XNOR U3167 ( .A(p_input[112]), .B(p_input[256]), .Z(n3190) );
  XNOR U3168 ( .A(n3177), .B(n3176), .Z(n3210) );
  XNOR U3169 ( .A(n3211), .B(n3184), .Z(n3176) );
  XNOR U3170 ( .A(n3172), .B(n3171), .Z(n3184) );
  XNOR U3171 ( .A(n3212), .B(n3168), .Z(n3171) );
  XNOR U3172 ( .A(p_input[122]), .B(p_input[266]), .Z(n3168) );
  XOR U3173 ( .A(p_input[123]), .B(n2060), .Z(n3212) );
  XOR U3174 ( .A(p_input[124]), .B(p_input[268]), .Z(n3172) );
  XOR U3175 ( .A(n3182), .B(n3213), .Z(n3211) );
  IV U3176 ( .A(n3173), .Z(n3213) );
  XOR U3177 ( .A(p_input[113]), .B(p_input[257]), .Z(n3173) );
  XNOR U3178 ( .A(n3214), .B(n3189), .Z(n3182) );
  XNOR U3179 ( .A(p_input[127]), .B(n2063), .Z(n3189) );
  XOR U3180 ( .A(n3179), .B(n3188), .Z(n3214) );
  XOR U3181 ( .A(n3215), .B(n3185), .Z(n3188) );
  XOR U3182 ( .A(p_input[125]), .B(p_input[269]), .Z(n3185) );
  XOR U3183 ( .A(p_input[126]), .B(n2065), .Z(n3215) );
  XOR U3184 ( .A(p_input[121]), .B(p_input[265]), .Z(n3179) );
  XOR U3185 ( .A(n3197), .B(n3195), .Z(n3177) );
  XNOR U3186 ( .A(n3216), .B(n3202), .Z(n3195) );
  XOR U3187 ( .A(p_input[120]), .B(p_input[264]), .Z(n3202) );
  XOR U3188 ( .A(n3192), .B(n3201), .Z(n3216) );
  XOR U3189 ( .A(n3217), .B(n3198), .Z(n3201) );
  XOR U3190 ( .A(p_input[118]), .B(p_input[262]), .Z(n3198) );
  XOR U3191 ( .A(p_input[119]), .B(n2239), .Z(n3217) );
  XOR U3192 ( .A(p_input[114]), .B(p_input[258]), .Z(n3192) );
  XNOR U3193 ( .A(n3207), .B(n3206), .Z(n3197) );
  XOR U3194 ( .A(n3218), .B(n3203), .Z(n3206) );
  XOR U3195 ( .A(p_input[115]), .B(p_input[259]), .Z(n3203) );
  XOR U3196 ( .A(p_input[116]), .B(n2241), .Z(n3218) );
  XOR U3197 ( .A(p_input[117]), .B(p_input[261]), .Z(n3207) );
  XNOR U3198 ( .A(n3219), .B(n3220), .Z(n3112) );
  AND U3199 ( .A(n116), .B(n3221), .Z(n3220) );
  XNOR U3200 ( .A(n3222), .B(n3223), .Z(n116) );
  AND U3201 ( .A(n3224), .B(n3225), .Z(n3223) );
  XOR U3202 ( .A(n3222), .B(n3122), .Z(n3225) );
  XNOR U3203 ( .A(n3222), .B(n3076), .Z(n3224) );
  XOR U3204 ( .A(n3226), .B(n3227), .Z(n3222) );
  AND U3205 ( .A(n3228), .B(n3229), .Z(n3227) );
  XOR U3206 ( .A(n3226), .B(n3086), .Z(n3228) );
  XOR U3207 ( .A(n3230), .B(n3231), .Z(n3065) );
  AND U3208 ( .A(n120), .B(n3221), .Z(n3231) );
  XNOR U3209 ( .A(n3219), .B(n3230), .Z(n3221) );
  XNOR U3210 ( .A(n3232), .B(n3233), .Z(n120) );
  AND U3211 ( .A(n3234), .B(n3235), .Z(n3233) );
  XNOR U3212 ( .A(n3236), .B(n3232), .Z(n3235) );
  IV U3213 ( .A(n3122), .Z(n3236) );
  XNOR U3214 ( .A(n3237), .B(n3238), .Z(n3122) );
  AND U3215 ( .A(n123), .B(n3239), .Z(n3238) );
  XNOR U3216 ( .A(n3237), .B(n3240), .Z(n3239) );
  XNOR U3217 ( .A(n3076), .B(n3232), .Z(n3234) );
  XNOR U3218 ( .A(n3241), .B(n3242), .Z(n3076) );
  AND U3219 ( .A(n131), .B(n3243), .Z(n3242) );
  XNOR U3220 ( .A(n3244), .B(n3245), .Z(n3243) );
  XOR U3221 ( .A(n3226), .B(n3246), .Z(n3232) );
  AND U3222 ( .A(n3247), .B(n3229), .Z(n3246) );
  XNOR U3223 ( .A(n3135), .B(n3226), .Z(n3229) );
  XNOR U3224 ( .A(n3248), .B(n3249), .Z(n3135) );
  AND U3225 ( .A(n123), .B(n3250), .Z(n3249) );
  XOR U3226 ( .A(n3251), .B(n3248), .Z(n3250) );
  XNOR U3227 ( .A(n3252), .B(n3226), .Z(n3247) );
  IV U3228 ( .A(n3086), .Z(n3252) );
  XOR U3229 ( .A(n3253), .B(n3254), .Z(n3086) );
  AND U3230 ( .A(n131), .B(n3255), .Z(n3254) );
  XOR U3231 ( .A(n3256), .B(n3257), .Z(n3226) );
  AND U3232 ( .A(n3258), .B(n3259), .Z(n3257) );
  XNOR U3233 ( .A(n3160), .B(n3256), .Z(n3259) );
  XNOR U3234 ( .A(n3260), .B(n3261), .Z(n3160) );
  AND U3235 ( .A(n123), .B(n3262), .Z(n3261) );
  XNOR U3236 ( .A(n3263), .B(n3260), .Z(n3262) );
  XOR U3237 ( .A(n3256), .B(n3097), .Z(n3258) );
  XOR U3238 ( .A(n3264), .B(n3265), .Z(n3097) );
  AND U3239 ( .A(n131), .B(n3266), .Z(n3265) );
  XOR U3240 ( .A(n3267), .B(n3268), .Z(n3256) );
  AND U3241 ( .A(n3269), .B(n3270), .Z(n3268) );
  XNOR U3242 ( .A(n3267), .B(n3208), .Z(n3270) );
  XNOR U3243 ( .A(n3271), .B(n3272), .Z(n3208) );
  AND U3244 ( .A(n123), .B(n3273), .Z(n3272) );
  XOR U3245 ( .A(n3274), .B(n3271), .Z(n3273) );
  XNOR U3246 ( .A(n3275), .B(n3267), .Z(n3269) );
  IV U3247 ( .A(n3109), .Z(n3275) );
  XOR U3248 ( .A(n3276), .B(n3277), .Z(n3109) );
  AND U3249 ( .A(n131), .B(n3278), .Z(n3277) );
  AND U3250 ( .A(n3230), .B(n3219), .Z(n3267) );
  XNOR U3251 ( .A(n3279), .B(n3280), .Z(n3219) );
  AND U3252 ( .A(n123), .B(n3281), .Z(n3280) );
  XNOR U3253 ( .A(n3282), .B(n3279), .Z(n3281) );
  XNOR U3254 ( .A(n3283), .B(n3284), .Z(n123) );
  AND U3255 ( .A(n3285), .B(n3286), .Z(n3284) );
  XOR U3256 ( .A(n3240), .B(n3283), .Z(n3286) );
  AND U3257 ( .A(n3287), .B(n3288), .Z(n3240) );
  XOR U3258 ( .A(n3283), .B(n3237), .Z(n3285) );
  XOR U3259 ( .A(n3244), .B(n3289), .Z(n3237) );
  AND U3260 ( .A(n127), .B(n3290), .Z(n3289) );
  XOR U3261 ( .A(n3244), .B(n3241), .Z(n3290) );
  XOR U3262 ( .A(n3291), .B(n3292), .Z(n3283) );
  AND U3263 ( .A(n3293), .B(n3294), .Z(n3292) );
  XNOR U3264 ( .A(n3291), .B(n3287), .Z(n3294) );
  IV U3265 ( .A(n3251), .Z(n3287) );
  XOR U3266 ( .A(n3295), .B(n3296), .Z(n3251) );
  XOR U3267 ( .A(n3297), .B(n3288), .Z(n3296) );
  AND U3268 ( .A(n3263), .B(n3298), .Z(n3288) );
  AND U3269 ( .A(n3299), .B(n3300), .Z(n3297) );
  XOR U3270 ( .A(n3301), .B(n3295), .Z(n3299) );
  XNOR U3271 ( .A(n3248), .B(n3291), .Z(n3293) );
  XNOR U3272 ( .A(n3302), .B(n3303), .Z(n3248) );
  AND U3273 ( .A(n127), .B(n3255), .Z(n3303) );
  XOR U3274 ( .A(n3302), .B(n3253), .Z(n3255) );
  XOR U3275 ( .A(n3304), .B(n3305), .Z(n3291) );
  AND U3276 ( .A(n3306), .B(n3307), .Z(n3305) );
  XNOR U3277 ( .A(n3304), .B(n3263), .Z(n3307) );
  XOR U3278 ( .A(n3308), .B(n3300), .Z(n3263) );
  XNOR U3279 ( .A(n3309), .B(n3295), .Z(n3300) );
  XOR U3280 ( .A(n3310), .B(n3311), .Z(n3295) );
  AND U3281 ( .A(n3312), .B(n3313), .Z(n3311) );
  XOR U3282 ( .A(n3314), .B(n3310), .Z(n3312) );
  XNOR U3283 ( .A(n3315), .B(n3316), .Z(n3309) );
  AND U3284 ( .A(n3317), .B(n3318), .Z(n3316) );
  XOR U3285 ( .A(n3315), .B(n3319), .Z(n3317) );
  XNOR U3286 ( .A(n3301), .B(n3298), .Z(n3308) );
  AND U3287 ( .A(n3320), .B(n3321), .Z(n3298) );
  XOR U3288 ( .A(n3322), .B(n3323), .Z(n3301) );
  AND U3289 ( .A(n3324), .B(n3325), .Z(n3323) );
  XOR U3290 ( .A(n3322), .B(n3326), .Z(n3324) );
  XNOR U3291 ( .A(n3260), .B(n3304), .Z(n3306) );
  XNOR U3292 ( .A(n3327), .B(n3328), .Z(n3260) );
  AND U3293 ( .A(n127), .B(n3266), .Z(n3328) );
  XOR U3294 ( .A(n3327), .B(n3264), .Z(n3266) );
  XOR U3295 ( .A(n3329), .B(n3330), .Z(n3304) );
  AND U3296 ( .A(n3331), .B(n3332), .Z(n3330) );
  XNOR U3297 ( .A(n3329), .B(n3320), .Z(n3332) );
  IV U3298 ( .A(n3274), .Z(n3320) );
  XNOR U3299 ( .A(n3333), .B(n3313), .Z(n3274) );
  XNOR U3300 ( .A(n3334), .B(n3319), .Z(n3313) );
  XNOR U3301 ( .A(n3335), .B(n3336), .Z(n3319) );
  NOR U3302 ( .A(n3337), .B(n3338), .Z(n3336) );
  XOR U3303 ( .A(n3335), .B(n3339), .Z(n3337) );
  XNOR U3304 ( .A(n3318), .B(n3310), .Z(n3334) );
  XOR U3305 ( .A(n3340), .B(n3341), .Z(n3310) );
  AND U3306 ( .A(n3342), .B(n3343), .Z(n3341) );
  XOR U3307 ( .A(n3340), .B(n3344), .Z(n3342) );
  XNOR U3308 ( .A(n3345), .B(n3315), .Z(n3318) );
  XOR U3309 ( .A(n3346), .B(n3347), .Z(n3315) );
  AND U3310 ( .A(n3348), .B(n3349), .Z(n3347) );
  XNOR U3311 ( .A(n3350), .B(n3351), .Z(n3348) );
  IV U3312 ( .A(n3346), .Z(n3350) );
  XNOR U3313 ( .A(n3352), .B(n3353), .Z(n3345) );
  NOR U3314 ( .A(n3354), .B(n3355), .Z(n3353) );
  XNOR U3315 ( .A(n3352), .B(n3356), .Z(n3354) );
  XNOR U3316 ( .A(n3314), .B(n3321), .Z(n3333) );
  NOR U3317 ( .A(n3282), .B(n3357), .Z(n3321) );
  XOR U3318 ( .A(n3326), .B(n3325), .Z(n3314) );
  XNOR U3319 ( .A(n3358), .B(n3322), .Z(n3325) );
  XOR U3320 ( .A(n3359), .B(n3360), .Z(n3322) );
  AND U3321 ( .A(n3361), .B(n3362), .Z(n3360) );
  XNOR U3322 ( .A(n3363), .B(n3364), .Z(n3361) );
  IV U3323 ( .A(n3359), .Z(n3363) );
  XNOR U3324 ( .A(n3365), .B(n3366), .Z(n3358) );
  NOR U3325 ( .A(n3367), .B(n3368), .Z(n3366) );
  XNOR U3326 ( .A(n3365), .B(n3369), .Z(n3367) );
  XOR U3327 ( .A(n3370), .B(n3371), .Z(n3326) );
  NOR U3328 ( .A(n3372), .B(n3373), .Z(n3371) );
  XNOR U3329 ( .A(n3370), .B(n3374), .Z(n3372) );
  XNOR U3330 ( .A(n3271), .B(n3329), .Z(n3331) );
  XNOR U3331 ( .A(n3375), .B(n3376), .Z(n3271) );
  AND U3332 ( .A(n127), .B(n3278), .Z(n3376) );
  XOR U3333 ( .A(n3375), .B(n3276), .Z(n3278) );
  AND U3334 ( .A(n3279), .B(n3282), .Z(n3329) );
  XOR U3335 ( .A(n3377), .B(n3357), .Z(n3282) );
  XNOR U3336 ( .A(p_input[128]), .B(p_input[256]), .Z(n3357) );
  XNOR U3337 ( .A(n3344), .B(n3343), .Z(n3377) );
  XNOR U3338 ( .A(n3378), .B(n3351), .Z(n3343) );
  XNOR U3339 ( .A(n3339), .B(n3338), .Z(n3351) );
  XNOR U3340 ( .A(n3379), .B(n3335), .Z(n3338) );
  XNOR U3341 ( .A(p_input[138]), .B(p_input[266]), .Z(n3335) );
  XOR U3342 ( .A(p_input[139]), .B(n2060), .Z(n3379) );
  XOR U3343 ( .A(p_input[140]), .B(p_input[268]), .Z(n3339) );
  XOR U3344 ( .A(n3349), .B(n3380), .Z(n3378) );
  IV U3345 ( .A(n3340), .Z(n3380) );
  XOR U3346 ( .A(p_input[129]), .B(p_input[257]), .Z(n3340) );
  XNOR U3347 ( .A(n3381), .B(n3356), .Z(n3349) );
  XNOR U3348 ( .A(p_input[143]), .B(n2063), .Z(n3356) );
  XOR U3349 ( .A(n3346), .B(n3355), .Z(n3381) );
  XOR U3350 ( .A(n3382), .B(n3352), .Z(n3355) );
  XOR U3351 ( .A(p_input[141]), .B(p_input[269]), .Z(n3352) );
  XOR U3352 ( .A(p_input[142]), .B(n2065), .Z(n3382) );
  XOR U3353 ( .A(p_input[137]), .B(p_input[265]), .Z(n3346) );
  XOR U3354 ( .A(n3364), .B(n3362), .Z(n3344) );
  XNOR U3355 ( .A(n3383), .B(n3369), .Z(n3362) );
  XOR U3356 ( .A(p_input[136]), .B(p_input[264]), .Z(n3369) );
  XOR U3357 ( .A(n3359), .B(n3368), .Z(n3383) );
  XOR U3358 ( .A(n3384), .B(n3365), .Z(n3368) );
  XOR U3359 ( .A(p_input[134]), .B(p_input[262]), .Z(n3365) );
  XOR U3360 ( .A(p_input[135]), .B(n2239), .Z(n3384) );
  XOR U3361 ( .A(p_input[130]), .B(p_input[258]), .Z(n3359) );
  XNOR U3362 ( .A(n3374), .B(n3373), .Z(n3364) );
  XOR U3363 ( .A(n3385), .B(n3370), .Z(n3373) );
  XOR U3364 ( .A(p_input[131]), .B(p_input[259]), .Z(n3370) );
  XOR U3365 ( .A(p_input[132]), .B(n2241), .Z(n3385) );
  XOR U3366 ( .A(p_input[133]), .B(p_input[261]), .Z(n3374) );
  XNOR U3367 ( .A(n3386), .B(n3387), .Z(n3279) );
  AND U3368 ( .A(n127), .B(n3388), .Z(n3387) );
  XNOR U3369 ( .A(n3389), .B(n3390), .Z(n127) );
  AND U3370 ( .A(n3391), .B(n3392), .Z(n3390) );
  XNOR U3371 ( .A(n3389), .B(n3244), .Z(n3392) );
  XOR U3372 ( .A(n3389), .B(n3241), .Z(n3391) );
  XOR U3373 ( .A(n3393), .B(n3394), .Z(n3389) );
  AND U3374 ( .A(n3395), .B(n3396), .Z(n3394) );
  XOR U3375 ( .A(n3393), .B(n3253), .Z(n3395) );
  XOR U3376 ( .A(n3397), .B(n3398), .Z(n3230) );
  AND U3377 ( .A(n131), .B(n3388), .Z(n3398) );
  XNOR U3378 ( .A(n3386), .B(n3397), .Z(n3388) );
  XNOR U3379 ( .A(n3399), .B(n3400), .Z(n131) );
  AND U3380 ( .A(n3401), .B(n3402), .Z(n3400) );
  XNOR U3381 ( .A(n3244), .B(n3399), .Z(n3402) );
  XOR U3382 ( .A(n3403), .B(n3404), .Z(n3244) );
  AND U3383 ( .A(n3405), .B(n134), .Z(n3404) );
  NOR U3384 ( .A(n3406), .B(n3403), .Z(n3405) );
  XOR U3385 ( .A(n3399), .B(n3241), .Z(n3401) );
  IV U3386 ( .A(n3245), .Z(n3241) );
  AND U3387 ( .A(n3407), .B(n3408), .Z(n3245) );
  XOR U3388 ( .A(n3393), .B(n3409), .Z(n3399) );
  AND U3389 ( .A(n3410), .B(n3396), .Z(n3409) );
  XNOR U3390 ( .A(n3302), .B(n3393), .Z(n3396) );
  XNOR U3391 ( .A(n3411), .B(n3412), .Z(n3302) );
  AND U3392 ( .A(n134), .B(n3413), .Z(n3412) );
  XOR U3393 ( .A(n3414), .B(n3411), .Z(n3413) );
  XNOR U3394 ( .A(n3415), .B(n3393), .Z(n3410) );
  IV U3395 ( .A(n3253), .Z(n3415) );
  XOR U3396 ( .A(n3416), .B(n3417), .Z(n3253) );
  AND U3397 ( .A(n142), .B(n3418), .Z(n3417) );
  XOR U3398 ( .A(n3419), .B(n3420), .Z(n3393) );
  AND U3399 ( .A(n3421), .B(n3422), .Z(n3420) );
  XNOR U3400 ( .A(n3327), .B(n3419), .Z(n3422) );
  XNOR U3401 ( .A(n3423), .B(n3424), .Z(n3327) );
  AND U3402 ( .A(n134), .B(n3425), .Z(n3424) );
  XNOR U3403 ( .A(n3426), .B(n3423), .Z(n3425) );
  XOR U3404 ( .A(n3419), .B(n3264), .Z(n3421) );
  XOR U3405 ( .A(n3427), .B(n3428), .Z(n3264) );
  AND U3406 ( .A(n142), .B(n3429), .Z(n3428) );
  XOR U3407 ( .A(n3430), .B(n3431), .Z(n3419) );
  AND U3408 ( .A(n3432), .B(n3433), .Z(n3431) );
  XNOR U3409 ( .A(n3430), .B(n3375), .Z(n3433) );
  XNOR U3410 ( .A(n3434), .B(n3435), .Z(n3375) );
  AND U3411 ( .A(n134), .B(n3436), .Z(n3435) );
  XOR U3412 ( .A(n3437), .B(n3434), .Z(n3436) );
  XNOR U3413 ( .A(n3438), .B(n3430), .Z(n3432) );
  IV U3414 ( .A(n3276), .Z(n3438) );
  XOR U3415 ( .A(n3439), .B(n3440), .Z(n3276) );
  AND U3416 ( .A(n142), .B(n3441), .Z(n3440) );
  AND U3417 ( .A(n3397), .B(n3386), .Z(n3430) );
  XNOR U3418 ( .A(n3442), .B(n3443), .Z(n3386) );
  AND U3419 ( .A(n134), .B(n3444), .Z(n3443) );
  XNOR U3420 ( .A(n3445), .B(n3442), .Z(n3444) );
  XNOR U3421 ( .A(n3446), .B(n3447), .Z(n134) );
  AND U3422 ( .A(n3448), .B(n3449), .Z(n3447) );
  XOR U3423 ( .A(n3406), .B(n3446), .Z(n3449) );
  AND U3424 ( .A(n3450), .B(n3451), .Z(n3406) );
  XOR U3425 ( .A(n3403), .B(n3446), .Z(n3448) );
  NOR U3426 ( .A(n3407), .B(n3408), .Z(n3403) );
  XOR U3427 ( .A(n3452), .B(n3453), .Z(n3446) );
  AND U3428 ( .A(n3454), .B(n3455), .Z(n3453) );
  XNOR U3429 ( .A(n3452), .B(n3450), .Z(n3455) );
  IV U3430 ( .A(n3414), .Z(n3450) );
  XOR U3431 ( .A(n3456), .B(n3457), .Z(n3414) );
  XOR U3432 ( .A(n3458), .B(n3451), .Z(n3457) );
  AND U3433 ( .A(n3426), .B(n3459), .Z(n3451) );
  AND U3434 ( .A(n3460), .B(n3461), .Z(n3458) );
  XOR U3435 ( .A(n3462), .B(n3456), .Z(n3460) );
  XNOR U3436 ( .A(n3411), .B(n3452), .Z(n3454) );
  XNOR U3437 ( .A(n3463), .B(n3464), .Z(n3411) );
  AND U3438 ( .A(n138), .B(n3418), .Z(n3464) );
  XOR U3439 ( .A(n3463), .B(n3416), .Z(n3418) );
  XOR U3440 ( .A(n3465), .B(n3466), .Z(n3452) );
  AND U3441 ( .A(n3467), .B(n3468), .Z(n3466) );
  XNOR U3442 ( .A(n3465), .B(n3426), .Z(n3468) );
  XOR U3443 ( .A(n3469), .B(n3461), .Z(n3426) );
  XNOR U3444 ( .A(n3470), .B(n3456), .Z(n3461) );
  XOR U3445 ( .A(n3471), .B(n3472), .Z(n3456) );
  AND U3446 ( .A(n3473), .B(n3474), .Z(n3472) );
  XOR U3447 ( .A(n3475), .B(n3471), .Z(n3473) );
  XNOR U3448 ( .A(n3476), .B(n3477), .Z(n3470) );
  AND U3449 ( .A(n3478), .B(n3479), .Z(n3477) );
  XOR U3450 ( .A(n3476), .B(n3480), .Z(n3478) );
  XNOR U3451 ( .A(n3462), .B(n3459), .Z(n3469) );
  AND U3452 ( .A(n3481), .B(n3482), .Z(n3459) );
  XOR U3453 ( .A(n3483), .B(n3484), .Z(n3462) );
  AND U3454 ( .A(n3485), .B(n3486), .Z(n3484) );
  XOR U3455 ( .A(n3483), .B(n3487), .Z(n3485) );
  XNOR U3456 ( .A(n3423), .B(n3465), .Z(n3467) );
  XNOR U3457 ( .A(n3488), .B(n3489), .Z(n3423) );
  AND U3458 ( .A(n138), .B(n3429), .Z(n3489) );
  XOR U3459 ( .A(n3488), .B(n3427), .Z(n3429) );
  XOR U3460 ( .A(n3490), .B(n3491), .Z(n3465) );
  AND U3461 ( .A(n3492), .B(n3493), .Z(n3491) );
  XNOR U3462 ( .A(n3490), .B(n3481), .Z(n3493) );
  IV U3463 ( .A(n3437), .Z(n3481) );
  XNOR U3464 ( .A(n3494), .B(n3474), .Z(n3437) );
  XNOR U3465 ( .A(n3495), .B(n3480), .Z(n3474) );
  XNOR U3466 ( .A(n3496), .B(n3497), .Z(n3480) );
  NOR U3467 ( .A(n3498), .B(n3499), .Z(n3497) );
  XOR U3468 ( .A(n3496), .B(n3500), .Z(n3498) );
  XNOR U3469 ( .A(n3479), .B(n3471), .Z(n3495) );
  XOR U3470 ( .A(n3501), .B(n3502), .Z(n3471) );
  AND U3471 ( .A(n3503), .B(n3504), .Z(n3502) );
  XOR U3472 ( .A(n3501), .B(n3505), .Z(n3503) );
  XNOR U3473 ( .A(n3506), .B(n3476), .Z(n3479) );
  XOR U3474 ( .A(n3507), .B(n3508), .Z(n3476) );
  AND U3475 ( .A(n3509), .B(n3510), .Z(n3508) );
  XNOR U3476 ( .A(n3511), .B(n3512), .Z(n3509) );
  IV U3477 ( .A(n3507), .Z(n3511) );
  XNOR U3478 ( .A(n3513), .B(n3514), .Z(n3506) );
  NOR U3479 ( .A(n3515), .B(n3516), .Z(n3514) );
  XNOR U3480 ( .A(n3513), .B(n3517), .Z(n3515) );
  XNOR U3481 ( .A(n3475), .B(n3482), .Z(n3494) );
  NOR U3482 ( .A(n3445), .B(n3518), .Z(n3482) );
  XOR U3483 ( .A(n3487), .B(n3486), .Z(n3475) );
  XNOR U3484 ( .A(n3519), .B(n3483), .Z(n3486) );
  XOR U3485 ( .A(n3520), .B(n3521), .Z(n3483) );
  AND U3486 ( .A(n3522), .B(n3523), .Z(n3521) );
  XNOR U3487 ( .A(n3524), .B(n3525), .Z(n3522) );
  IV U3488 ( .A(n3520), .Z(n3524) );
  XNOR U3489 ( .A(n3526), .B(n3527), .Z(n3519) );
  NOR U3490 ( .A(n3528), .B(n3529), .Z(n3527) );
  XNOR U3491 ( .A(n3526), .B(n3530), .Z(n3528) );
  XOR U3492 ( .A(n3531), .B(n3532), .Z(n3487) );
  NOR U3493 ( .A(n3533), .B(n3534), .Z(n3532) );
  XNOR U3494 ( .A(n3531), .B(n3535), .Z(n3533) );
  XNOR U3495 ( .A(n3434), .B(n3490), .Z(n3492) );
  XNOR U3496 ( .A(n3536), .B(n3537), .Z(n3434) );
  AND U3497 ( .A(n138), .B(n3441), .Z(n3537) );
  XOR U3498 ( .A(n3536), .B(n3439), .Z(n3441) );
  AND U3499 ( .A(n3442), .B(n3445), .Z(n3490) );
  XOR U3500 ( .A(n3538), .B(n3518), .Z(n3445) );
  XNOR U3501 ( .A(p_input[144]), .B(p_input[256]), .Z(n3518) );
  XNOR U3502 ( .A(n3505), .B(n3504), .Z(n3538) );
  XNOR U3503 ( .A(n3539), .B(n3512), .Z(n3504) );
  XNOR U3504 ( .A(n3500), .B(n3499), .Z(n3512) );
  XNOR U3505 ( .A(n3540), .B(n3496), .Z(n3499) );
  XNOR U3506 ( .A(p_input[154]), .B(p_input[266]), .Z(n3496) );
  XOR U3507 ( .A(p_input[155]), .B(n2060), .Z(n3540) );
  XOR U3508 ( .A(p_input[156]), .B(p_input[268]), .Z(n3500) );
  XOR U3509 ( .A(n3510), .B(n3541), .Z(n3539) );
  IV U3510 ( .A(n3501), .Z(n3541) );
  XOR U3511 ( .A(p_input[145]), .B(p_input[257]), .Z(n3501) );
  XNOR U3512 ( .A(n3542), .B(n3517), .Z(n3510) );
  XNOR U3513 ( .A(p_input[159]), .B(n2063), .Z(n3517) );
  XOR U3514 ( .A(n3507), .B(n3516), .Z(n3542) );
  XOR U3515 ( .A(n3543), .B(n3513), .Z(n3516) );
  XOR U3516 ( .A(p_input[157]), .B(p_input[269]), .Z(n3513) );
  XOR U3517 ( .A(p_input[158]), .B(n2065), .Z(n3543) );
  XOR U3518 ( .A(p_input[153]), .B(p_input[265]), .Z(n3507) );
  XOR U3519 ( .A(n3525), .B(n3523), .Z(n3505) );
  XNOR U3520 ( .A(n3544), .B(n3530), .Z(n3523) );
  XOR U3521 ( .A(p_input[152]), .B(p_input[264]), .Z(n3530) );
  XOR U3522 ( .A(n3520), .B(n3529), .Z(n3544) );
  XOR U3523 ( .A(n3545), .B(n3526), .Z(n3529) );
  XOR U3524 ( .A(p_input[150]), .B(p_input[262]), .Z(n3526) );
  XOR U3525 ( .A(p_input[151]), .B(n2239), .Z(n3545) );
  XOR U3526 ( .A(p_input[146]), .B(p_input[258]), .Z(n3520) );
  XNOR U3527 ( .A(n3535), .B(n3534), .Z(n3525) );
  XOR U3528 ( .A(n3546), .B(n3531), .Z(n3534) );
  XOR U3529 ( .A(p_input[147]), .B(p_input[259]), .Z(n3531) );
  XOR U3530 ( .A(p_input[148]), .B(n2241), .Z(n3546) );
  XOR U3531 ( .A(p_input[149]), .B(p_input[261]), .Z(n3535) );
  XNOR U3532 ( .A(n3547), .B(n3548), .Z(n3442) );
  AND U3533 ( .A(n138), .B(n3549), .Z(n3548) );
  XNOR U3534 ( .A(n3550), .B(n3551), .Z(n138) );
  NOR U3535 ( .A(n3552), .B(n3553), .Z(n3551) );
  XOR U3536 ( .A(n3408), .B(n3550), .Z(n3553) );
  NOR U3537 ( .A(n3550), .B(n3407), .Z(n3552) );
  XOR U3538 ( .A(n3554), .B(n3555), .Z(n3550) );
  AND U3539 ( .A(n3556), .B(n3557), .Z(n3555) );
  XOR U3540 ( .A(n3554), .B(n3416), .Z(n3556) );
  XOR U3541 ( .A(n3558), .B(n3559), .Z(n3397) );
  AND U3542 ( .A(n142), .B(n3549), .Z(n3559) );
  XNOR U3543 ( .A(n3547), .B(n3558), .Z(n3549) );
  XNOR U3544 ( .A(n3560), .B(n3561), .Z(n142) );
  NOR U3545 ( .A(n3562), .B(n3563), .Z(n3561) );
  XNOR U3546 ( .A(n3408), .B(n3564), .Z(n3563) );
  IV U3547 ( .A(n3560), .Z(n3564) );
  AND U3548 ( .A(n3565), .B(n3566), .Z(n3408) );
  NOR U3549 ( .A(n3560), .B(n3407), .Z(n3562) );
  AND U3550 ( .A(n3567), .B(n3568), .Z(n3407) );
  IV U3551 ( .A(n3569), .Z(n3567) );
  XOR U3552 ( .A(n3554), .B(n3570), .Z(n3560) );
  AND U3553 ( .A(n3571), .B(n3557), .Z(n3570) );
  XNOR U3554 ( .A(n3463), .B(n3554), .Z(n3557) );
  XNOR U3555 ( .A(n3572), .B(n3573), .Z(n3463) );
  AND U3556 ( .A(n145), .B(n3574), .Z(n3573) );
  XOR U3557 ( .A(n3575), .B(n3572), .Z(n3574) );
  XNOR U3558 ( .A(n3576), .B(n3554), .Z(n3571) );
  IV U3559 ( .A(n3416), .Z(n3576) );
  XOR U3560 ( .A(n3577), .B(n3578), .Z(n3416) );
  AND U3561 ( .A(n153), .B(n3579), .Z(n3578) );
  XOR U3562 ( .A(n3580), .B(n3581), .Z(n3554) );
  AND U3563 ( .A(n3582), .B(n3583), .Z(n3581) );
  XNOR U3564 ( .A(n3488), .B(n3580), .Z(n3583) );
  XNOR U3565 ( .A(n3584), .B(n3585), .Z(n3488) );
  AND U3566 ( .A(n145), .B(n3586), .Z(n3585) );
  XNOR U3567 ( .A(n3587), .B(n3584), .Z(n3586) );
  XOR U3568 ( .A(n3580), .B(n3427), .Z(n3582) );
  XOR U3569 ( .A(n3588), .B(n3589), .Z(n3427) );
  AND U3570 ( .A(n153), .B(n3590), .Z(n3589) );
  XOR U3571 ( .A(n3591), .B(n3592), .Z(n3580) );
  AND U3572 ( .A(n3593), .B(n3594), .Z(n3592) );
  XNOR U3573 ( .A(n3591), .B(n3536), .Z(n3594) );
  XNOR U3574 ( .A(n3595), .B(n3596), .Z(n3536) );
  AND U3575 ( .A(n145), .B(n3597), .Z(n3596) );
  XOR U3576 ( .A(n3598), .B(n3595), .Z(n3597) );
  XNOR U3577 ( .A(n3599), .B(n3591), .Z(n3593) );
  IV U3578 ( .A(n3439), .Z(n3599) );
  XOR U3579 ( .A(n3600), .B(n3601), .Z(n3439) );
  AND U3580 ( .A(n153), .B(n3602), .Z(n3601) );
  AND U3581 ( .A(n3558), .B(n3547), .Z(n3591) );
  XNOR U3582 ( .A(n3603), .B(n3604), .Z(n3547) );
  AND U3583 ( .A(n145), .B(n3605), .Z(n3604) );
  XNOR U3584 ( .A(n3606), .B(n3603), .Z(n3605) );
  XNOR U3585 ( .A(n3607), .B(n3608), .Z(n145) );
  NOR U3586 ( .A(n3609), .B(n3610), .Z(n3608) );
  XNOR U3587 ( .A(n3607), .B(n3569), .Z(n3610) );
  NOR U3588 ( .A(n3565), .B(n3566), .Z(n3569) );
  NOR U3589 ( .A(n3607), .B(n3568), .Z(n3609) );
  AND U3590 ( .A(n3611), .B(n3612), .Z(n3568) );
  XOR U3591 ( .A(n3613), .B(n3614), .Z(n3607) );
  AND U3592 ( .A(n3615), .B(n3616), .Z(n3614) );
  XNOR U3593 ( .A(n3613), .B(n3611), .Z(n3616) );
  IV U3594 ( .A(n3575), .Z(n3611) );
  XOR U3595 ( .A(n3617), .B(n3618), .Z(n3575) );
  XOR U3596 ( .A(n3619), .B(n3612), .Z(n3618) );
  AND U3597 ( .A(n3587), .B(n3620), .Z(n3612) );
  AND U3598 ( .A(n3621), .B(n3622), .Z(n3619) );
  XOR U3599 ( .A(n3623), .B(n3617), .Z(n3621) );
  XNOR U3600 ( .A(n3572), .B(n3613), .Z(n3615) );
  XNOR U3601 ( .A(n3624), .B(n3625), .Z(n3572) );
  AND U3602 ( .A(n149), .B(n3579), .Z(n3625) );
  XOR U3603 ( .A(n3624), .B(n3577), .Z(n3579) );
  XOR U3604 ( .A(n3626), .B(n3627), .Z(n3613) );
  AND U3605 ( .A(n3628), .B(n3629), .Z(n3627) );
  XNOR U3606 ( .A(n3626), .B(n3587), .Z(n3629) );
  XOR U3607 ( .A(n3630), .B(n3622), .Z(n3587) );
  XNOR U3608 ( .A(n3631), .B(n3617), .Z(n3622) );
  XOR U3609 ( .A(n3632), .B(n3633), .Z(n3617) );
  AND U3610 ( .A(n3634), .B(n3635), .Z(n3633) );
  XOR U3611 ( .A(n3636), .B(n3632), .Z(n3634) );
  XNOR U3612 ( .A(n3637), .B(n3638), .Z(n3631) );
  AND U3613 ( .A(n3639), .B(n3640), .Z(n3638) );
  XOR U3614 ( .A(n3637), .B(n3641), .Z(n3639) );
  XNOR U3615 ( .A(n3623), .B(n3620), .Z(n3630) );
  AND U3616 ( .A(n3642), .B(n3643), .Z(n3620) );
  XOR U3617 ( .A(n3644), .B(n3645), .Z(n3623) );
  AND U3618 ( .A(n3646), .B(n3647), .Z(n3645) );
  XOR U3619 ( .A(n3644), .B(n3648), .Z(n3646) );
  XNOR U3620 ( .A(n3584), .B(n3626), .Z(n3628) );
  XNOR U3621 ( .A(n3649), .B(n3650), .Z(n3584) );
  AND U3622 ( .A(n149), .B(n3590), .Z(n3650) );
  XOR U3623 ( .A(n3649), .B(n3588), .Z(n3590) );
  XOR U3624 ( .A(n3651), .B(n3652), .Z(n3626) );
  AND U3625 ( .A(n3653), .B(n3654), .Z(n3652) );
  XNOR U3626 ( .A(n3651), .B(n3642), .Z(n3654) );
  IV U3627 ( .A(n3598), .Z(n3642) );
  XNOR U3628 ( .A(n3655), .B(n3635), .Z(n3598) );
  XNOR U3629 ( .A(n3656), .B(n3641), .Z(n3635) );
  XNOR U3630 ( .A(n3657), .B(n3658), .Z(n3641) );
  NOR U3631 ( .A(n3659), .B(n3660), .Z(n3658) );
  XOR U3632 ( .A(n3657), .B(n3661), .Z(n3659) );
  XNOR U3633 ( .A(n3640), .B(n3632), .Z(n3656) );
  XOR U3634 ( .A(n3662), .B(n3663), .Z(n3632) );
  AND U3635 ( .A(n3664), .B(n3665), .Z(n3663) );
  XOR U3636 ( .A(n3662), .B(n3666), .Z(n3664) );
  XNOR U3637 ( .A(n3667), .B(n3637), .Z(n3640) );
  XOR U3638 ( .A(n3668), .B(n3669), .Z(n3637) );
  AND U3639 ( .A(n3670), .B(n3671), .Z(n3669) );
  XNOR U3640 ( .A(n3672), .B(n3673), .Z(n3670) );
  IV U3641 ( .A(n3668), .Z(n3672) );
  XNOR U3642 ( .A(n3674), .B(n3675), .Z(n3667) );
  NOR U3643 ( .A(n3676), .B(n3677), .Z(n3675) );
  XNOR U3644 ( .A(n3674), .B(n3678), .Z(n3676) );
  XNOR U3645 ( .A(n3636), .B(n3643), .Z(n3655) );
  NOR U3646 ( .A(n3606), .B(n3679), .Z(n3643) );
  XOR U3647 ( .A(n3648), .B(n3647), .Z(n3636) );
  XNOR U3648 ( .A(n3680), .B(n3644), .Z(n3647) );
  XOR U3649 ( .A(n3681), .B(n3682), .Z(n3644) );
  AND U3650 ( .A(n3683), .B(n3684), .Z(n3682) );
  XNOR U3651 ( .A(n3685), .B(n3686), .Z(n3683) );
  IV U3652 ( .A(n3681), .Z(n3685) );
  XNOR U3653 ( .A(n3687), .B(n3688), .Z(n3680) );
  NOR U3654 ( .A(n3689), .B(n3690), .Z(n3688) );
  XNOR U3655 ( .A(n3687), .B(n3691), .Z(n3689) );
  XOR U3656 ( .A(n3692), .B(n3693), .Z(n3648) );
  NOR U3657 ( .A(n3694), .B(n3695), .Z(n3693) );
  XNOR U3658 ( .A(n3692), .B(n3696), .Z(n3694) );
  XNOR U3659 ( .A(n3595), .B(n3651), .Z(n3653) );
  XNOR U3660 ( .A(n3697), .B(n3698), .Z(n3595) );
  AND U3661 ( .A(n149), .B(n3602), .Z(n3698) );
  XOR U3662 ( .A(n3697), .B(n3600), .Z(n3602) );
  AND U3663 ( .A(n3603), .B(n3606), .Z(n3651) );
  XOR U3664 ( .A(n3699), .B(n3679), .Z(n3606) );
  XNOR U3665 ( .A(p_input[160]), .B(p_input[256]), .Z(n3679) );
  XNOR U3666 ( .A(n3666), .B(n3665), .Z(n3699) );
  XNOR U3667 ( .A(n3700), .B(n3673), .Z(n3665) );
  XNOR U3668 ( .A(n3661), .B(n3660), .Z(n3673) );
  XNOR U3669 ( .A(n3701), .B(n3657), .Z(n3660) );
  XNOR U3670 ( .A(p_input[170]), .B(p_input[266]), .Z(n3657) );
  XOR U3671 ( .A(p_input[171]), .B(n2060), .Z(n3701) );
  XOR U3672 ( .A(p_input[172]), .B(p_input[268]), .Z(n3661) );
  XOR U3673 ( .A(n3671), .B(n3702), .Z(n3700) );
  IV U3674 ( .A(n3662), .Z(n3702) );
  XOR U3675 ( .A(p_input[161]), .B(p_input[257]), .Z(n3662) );
  XNOR U3676 ( .A(n3703), .B(n3678), .Z(n3671) );
  XNOR U3677 ( .A(p_input[175]), .B(n2063), .Z(n3678) );
  XOR U3678 ( .A(n3668), .B(n3677), .Z(n3703) );
  XOR U3679 ( .A(n3704), .B(n3674), .Z(n3677) );
  XOR U3680 ( .A(p_input[173]), .B(p_input[269]), .Z(n3674) );
  XOR U3681 ( .A(p_input[174]), .B(n2065), .Z(n3704) );
  XOR U3682 ( .A(p_input[169]), .B(p_input[265]), .Z(n3668) );
  XOR U3683 ( .A(n3686), .B(n3684), .Z(n3666) );
  XNOR U3684 ( .A(n3705), .B(n3691), .Z(n3684) );
  XOR U3685 ( .A(p_input[168]), .B(p_input[264]), .Z(n3691) );
  XOR U3686 ( .A(n3681), .B(n3690), .Z(n3705) );
  XOR U3687 ( .A(n3706), .B(n3687), .Z(n3690) );
  XOR U3688 ( .A(p_input[166]), .B(p_input[262]), .Z(n3687) );
  XOR U3689 ( .A(p_input[167]), .B(n2239), .Z(n3706) );
  XOR U3690 ( .A(p_input[162]), .B(p_input[258]), .Z(n3681) );
  XNOR U3691 ( .A(n3696), .B(n3695), .Z(n3686) );
  XOR U3692 ( .A(n3707), .B(n3692), .Z(n3695) );
  XOR U3693 ( .A(p_input[163]), .B(p_input[259]), .Z(n3692) );
  XOR U3694 ( .A(p_input[164]), .B(n2241), .Z(n3707) );
  XOR U3695 ( .A(p_input[165]), .B(p_input[261]), .Z(n3696) );
  XNOR U3696 ( .A(n3708), .B(n3709), .Z(n3603) );
  AND U3697 ( .A(n149), .B(n3710), .Z(n3709) );
  XNOR U3698 ( .A(n3711), .B(n3712), .Z(n149) );
  NOR U3699 ( .A(n3713), .B(n3714), .Z(n3712) );
  XOR U3700 ( .A(n3566), .B(n3711), .Z(n3714) );
  NOR U3701 ( .A(n3711), .B(n3565), .Z(n3713) );
  XOR U3702 ( .A(n3715), .B(n3716), .Z(n3711) );
  AND U3703 ( .A(n3717), .B(n3718), .Z(n3716) );
  XOR U3704 ( .A(n3715), .B(n3577), .Z(n3717) );
  XOR U3705 ( .A(n3719), .B(n3720), .Z(n3558) );
  AND U3706 ( .A(n153), .B(n3710), .Z(n3720) );
  XNOR U3707 ( .A(n3708), .B(n3719), .Z(n3710) );
  XNOR U3708 ( .A(n3721), .B(n3722), .Z(n153) );
  NOR U3709 ( .A(n3723), .B(n3724), .Z(n3722) );
  XNOR U3710 ( .A(n3566), .B(n3725), .Z(n3724) );
  IV U3711 ( .A(n3721), .Z(n3725) );
  AND U3712 ( .A(n3726), .B(n3727), .Z(n3566) );
  NOR U3713 ( .A(n3721), .B(n3565), .Z(n3723) );
  AND U3714 ( .A(n3728), .B(n3729), .Z(n3565) );
  IV U3715 ( .A(n3730), .Z(n3728) );
  XOR U3716 ( .A(n3715), .B(n3731), .Z(n3721) );
  AND U3717 ( .A(n3732), .B(n3718), .Z(n3731) );
  XNOR U3718 ( .A(n3624), .B(n3715), .Z(n3718) );
  XNOR U3719 ( .A(n3733), .B(n3734), .Z(n3624) );
  AND U3720 ( .A(n156), .B(n3735), .Z(n3734) );
  XOR U3721 ( .A(n3736), .B(n3733), .Z(n3735) );
  XNOR U3722 ( .A(n3737), .B(n3715), .Z(n3732) );
  IV U3723 ( .A(n3577), .Z(n3737) );
  XOR U3724 ( .A(n3738), .B(n3739), .Z(n3577) );
  AND U3725 ( .A(n164), .B(n3740), .Z(n3739) );
  XOR U3726 ( .A(n3741), .B(n3742), .Z(n3715) );
  AND U3727 ( .A(n3743), .B(n3744), .Z(n3742) );
  XNOR U3728 ( .A(n3649), .B(n3741), .Z(n3744) );
  XNOR U3729 ( .A(n3745), .B(n3746), .Z(n3649) );
  AND U3730 ( .A(n156), .B(n3747), .Z(n3746) );
  XNOR U3731 ( .A(n3748), .B(n3745), .Z(n3747) );
  XOR U3732 ( .A(n3741), .B(n3588), .Z(n3743) );
  XOR U3733 ( .A(n3749), .B(n3750), .Z(n3588) );
  AND U3734 ( .A(n164), .B(n3751), .Z(n3750) );
  XOR U3735 ( .A(n3752), .B(n3753), .Z(n3741) );
  AND U3736 ( .A(n3754), .B(n3755), .Z(n3753) );
  XNOR U3737 ( .A(n3752), .B(n3697), .Z(n3755) );
  XNOR U3738 ( .A(n3756), .B(n3757), .Z(n3697) );
  AND U3739 ( .A(n156), .B(n3758), .Z(n3757) );
  XOR U3740 ( .A(n3759), .B(n3756), .Z(n3758) );
  XNOR U3741 ( .A(n3760), .B(n3752), .Z(n3754) );
  IV U3742 ( .A(n3600), .Z(n3760) );
  XOR U3743 ( .A(n3761), .B(n3762), .Z(n3600) );
  AND U3744 ( .A(n164), .B(n3763), .Z(n3762) );
  AND U3745 ( .A(n3719), .B(n3708), .Z(n3752) );
  XNOR U3746 ( .A(n3764), .B(n3765), .Z(n3708) );
  AND U3747 ( .A(n156), .B(n3766), .Z(n3765) );
  XNOR U3748 ( .A(n3767), .B(n3764), .Z(n3766) );
  XNOR U3749 ( .A(n3768), .B(n3769), .Z(n156) );
  NOR U3750 ( .A(n3770), .B(n3771), .Z(n3769) );
  XNOR U3751 ( .A(n3768), .B(n3730), .Z(n3771) );
  NOR U3752 ( .A(n3726), .B(n3727), .Z(n3730) );
  NOR U3753 ( .A(n3768), .B(n3729), .Z(n3770) );
  AND U3754 ( .A(n3772), .B(n3773), .Z(n3729) );
  XOR U3755 ( .A(n3774), .B(n3775), .Z(n3768) );
  AND U3756 ( .A(n3776), .B(n3777), .Z(n3775) );
  XNOR U3757 ( .A(n3774), .B(n3772), .Z(n3777) );
  IV U3758 ( .A(n3736), .Z(n3772) );
  XOR U3759 ( .A(n3778), .B(n3779), .Z(n3736) );
  XOR U3760 ( .A(n3780), .B(n3773), .Z(n3779) );
  AND U3761 ( .A(n3748), .B(n3781), .Z(n3773) );
  AND U3762 ( .A(n3782), .B(n3783), .Z(n3780) );
  XOR U3763 ( .A(n3784), .B(n3778), .Z(n3782) );
  XNOR U3764 ( .A(n3733), .B(n3774), .Z(n3776) );
  XNOR U3765 ( .A(n3785), .B(n3786), .Z(n3733) );
  AND U3766 ( .A(n160), .B(n3740), .Z(n3786) );
  XOR U3767 ( .A(n3785), .B(n3738), .Z(n3740) );
  XOR U3768 ( .A(n3787), .B(n3788), .Z(n3774) );
  AND U3769 ( .A(n3789), .B(n3790), .Z(n3788) );
  XNOR U3770 ( .A(n3787), .B(n3748), .Z(n3790) );
  XOR U3771 ( .A(n3791), .B(n3783), .Z(n3748) );
  XNOR U3772 ( .A(n3792), .B(n3778), .Z(n3783) );
  XOR U3773 ( .A(n3793), .B(n3794), .Z(n3778) );
  AND U3774 ( .A(n3795), .B(n3796), .Z(n3794) );
  XOR U3775 ( .A(n3797), .B(n3793), .Z(n3795) );
  XNOR U3776 ( .A(n3798), .B(n3799), .Z(n3792) );
  AND U3777 ( .A(n3800), .B(n3801), .Z(n3799) );
  XOR U3778 ( .A(n3798), .B(n3802), .Z(n3800) );
  XNOR U3779 ( .A(n3784), .B(n3781), .Z(n3791) );
  AND U3780 ( .A(n3803), .B(n3804), .Z(n3781) );
  XOR U3781 ( .A(n3805), .B(n3806), .Z(n3784) );
  AND U3782 ( .A(n3807), .B(n3808), .Z(n3806) );
  XOR U3783 ( .A(n3805), .B(n3809), .Z(n3807) );
  XNOR U3784 ( .A(n3745), .B(n3787), .Z(n3789) );
  XNOR U3785 ( .A(n3810), .B(n3811), .Z(n3745) );
  AND U3786 ( .A(n160), .B(n3751), .Z(n3811) );
  XOR U3787 ( .A(n3810), .B(n3749), .Z(n3751) );
  XOR U3788 ( .A(n3812), .B(n3813), .Z(n3787) );
  AND U3789 ( .A(n3814), .B(n3815), .Z(n3813) );
  XNOR U3790 ( .A(n3812), .B(n3803), .Z(n3815) );
  IV U3791 ( .A(n3759), .Z(n3803) );
  XNOR U3792 ( .A(n3816), .B(n3796), .Z(n3759) );
  XNOR U3793 ( .A(n3817), .B(n3802), .Z(n3796) );
  XNOR U3794 ( .A(n3818), .B(n3819), .Z(n3802) );
  NOR U3795 ( .A(n3820), .B(n3821), .Z(n3819) );
  XOR U3796 ( .A(n3818), .B(n3822), .Z(n3820) );
  XNOR U3797 ( .A(n3801), .B(n3793), .Z(n3817) );
  XOR U3798 ( .A(n3823), .B(n3824), .Z(n3793) );
  AND U3799 ( .A(n3825), .B(n3826), .Z(n3824) );
  XOR U3800 ( .A(n3823), .B(n3827), .Z(n3825) );
  XNOR U3801 ( .A(n3828), .B(n3798), .Z(n3801) );
  XOR U3802 ( .A(n3829), .B(n3830), .Z(n3798) );
  AND U3803 ( .A(n3831), .B(n3832), .Z(n3830) );
  XNOR U3804 ( .A(n3833), .B(n3834), .Z(n3831) );
  IV U3805 ( .A(n3829), .Z(n3833) );
  XNOR U3806 ( .A(n3835), .B(n3836), .Z(n3828) );
  NOR U3807 ( .A(n3837), .B(n3838), .Z(n3836) );
  XNOR U3808 ( .A(n3835), .B(n3839), .Z(n3837) );
  XNOR U3809 ( .A(n3797), .B(n3804), .Z(n3816) );
  NOR U3810 ( .A(n3767), .B(n3840), .Z(n3804) );
  XOR U3811 ( .A(n3809), .B(n3808), .Z(n3797) );
  XNOR U3812 ( .A(n3841), .B(n3805), .Z(n3808) );
  XOR U3813 ( .A(n3842), .B(n3843), .Z(n3805) );
  AND U3814 ( .A(n3844), .B(n3845), .Z(n3843) );
  XNOR U3815 ( .A(n3846), .B(n3847), .Z(n3844) );
  IV U3816 ( .A(n3842), .Z(n3846) );
  XNOR U3817 ( .A(n3848), .B(n3849), .Z(n3841) );
  NOR U3818 ( .A(n3850), .B(n3851), .Z(n3849) );
  XNOR U3819 ( .A(n3848), .B(n3852), .Z(n3850) );
  XOR U3820 ( .A(n3853), .B(n3854), .Z(n3809) );
  NOR U3821 ( .A(n3855), .B(n3856), .Z(n3854) );
  XNOR U3822 ( .A(n3853), .B(n3857), .Z(n3855) );
  XNOR U3823 ( .A(n3756), .B(n3812), .Z(n3814) );
  XNOR U3824 ( .A(n3858), .B(n3859), .Z(n3756) );
  AND U3825 ( .A(n160), .B(n3763), .Z(n3859) );
  XOR U3826 ( .A(n3858), .B(n3761), .Z(n3763) );
  AND U3827 ( .A(n3764), .B(n3767), .Z(n3812) );
  XOR U3828 ( .A(n3860), .B(n3840), .Z(n3767) );
  XNOR U3829 ( .A(p_input[176]), .B(p_input[256]), .Z(n3840) );
  XNOR U3830 ( .A(n3827), .B(n3826), .Z(n3860) );
  XNOR U3831 ( .A(n3861), .B(n3834), .Z(n3826) );
  XNOR U3832 ( .A(n3822), .B(n3821), .Z(n3834) );
  XNOR U3833 ( .A(n3862), .B(n3818), .Z(n3821) );
  XNOR U3834 ( .A(p_input[186]), .B(p_input[266]), .Z(n3818) );
  XOR U3835 ( .A(p_input[187]), .B(n2060), .Z(n3862) );
  XOR U3836 ( .A(p_input[188]), .B(p_input[268]), .Z(n3822) );
  XOR U3837 ( .A(n3832), .B(n3863), .Z(n3861) );
  IV U3838 ( .A(n3823), .Z(n3863) );
  XOR U3839 ( .A(p_input[177]), .B(p_input[257]), .Z(n3823) );
  XNOR U3840 ( .A(n3864), .B(n3839), .Z(n3832) );
  XNOR U3841 ( .A(p_input[191]), .B(n2063), .Z(n3839) );
  XOR U3842 ( .A(n3829), .B(n3838), .Z(n3864) );
  XOR U3843 ( .A(n3865), .B(n3835), .Z(n3838) );
  XOR U3844 ( .A(p_input[189]), .B(p_input[269]), .Z(n3835) );
  XOR U3845 ( .A(p_input[190]), .B(n2065), .Z(n3865) );
  XOR U3846 ( .A(p_input[185]), .B(p_input[265]), .Z(n3829) );
  XOR U3847 ( .A(n3847), .B(n3845), .Z(n3827) );
  XNOR U3848 ( .A(n3866), .B(n3852), .Z(n3845) );
  XOR U3849 ( .A(p_input[184]), .B(p_input[264]), .Z(n3852) );
  XOR U3850 ( .A(n3842), .B(n3851), .Z(n3866) );
  XOR U3851 ( .A(n3867), .B(n3848), .Z(n3851) );
  XOR U3852 ( .A(p_input[182]), .B(p_input[262]), .Z(n3848) );
  XOR U3853 ( .A(p_input[183]), .B(n2239), .Z(n3867) );
  XOR U3854 ( .A(p_input[178]), .B(p_input[258]), .Z(n3842) );
  XNOR U3855 ( .A(n3857), .B(n3856), .Z(n3847) );
  XOR U3856 ( .A(n3868), .B(n3853), .Z(n3856) );
  XOR U3857 ( .A(p_input[179]), .B(p_input[259]), .Z(n3853) );
  XOR U3858 ( .A(p_input[180]), .B(n2241), .Z(n3868) );
  XOR U3859 ( .A(p_input[181]), .B(p_input[261]), .Z(n3857) );
  XNOR U3860 ( .A(n3869), .B(n3870), .Z(n3764) );
  AND U3861 ( .A(n160), .B(n3871), .Z(n3870) );
  XNOR U3862 ( .A(n3872), .B(n3873), .Z(n160) );
  NOR U3863 ( .A(n3874), .B(n3875), .Z(n3873) );
  XOR U3864 ( .A(n3727), .B(n3872), .Z(n3875) );
  NOR U3865 ( .A(n3872), .B(n3726), .Z(n3874) );
  XOR U3866 ( .A(n3876), .B(n3877), .Z(n3872) );
  AND U3867 ( .A(n3878), .B(n3879), .Z(n3877) );
  XOR U3868 ( .A(n3876), .B(n3738), .Z(n3878) );
  XOR U3869 ( .A(n3880), .B(n3881), .Z(n3719) );
  AND U3870 ( .A(n164), .B(n3871), .Z(n3881) );
  XNOR U3871 ( .A(n3869), .B(n3880), .Z(n3871) );
  XNOR U3872 ( .A(n3882), .B(n3883), .Z(n164) );
  NOR U3873 ( .A(n3884), .B(n3885), .Z(n3883) );
  XNOR U3874 ( .A(n3727), .B(n3886), .Z(n3885) );
  IV U3875 ( .A(n3882), .Z(n3886) );
  AND U3876 ( .A(n3887), .B(n3888), .Z(n3727) );
  NOR U3877 ( .A(n3882), .B(n3726), .Z(n3884) );
  AND U3878 ( .A(n3889), .B(n3890), .Z(n3726) );
  IV U3879 ( .A(n3891), .Z(n3889) );
  XOR U3880 ( .A(n3876), .B(n3892), .Z(n3882) );
  AND U3881 ( .A(n3893), .B(n3879), .Z(n3892) );
  XNOR U3882 ( .A(n3785), .B(n3876), .Z(n3879) );
  XNOR U3883 ( .A(n3894), .B(n3895), .Z(n3785) );
  AND U3884 ( .A(n167), .B(n3896), .Z(n3895) );
  XOR U3885 ( .A(n3897), .B(n3894), .Z(n3896) );
  XNOR U3886 ( .A(n3898), .B(n3876), .Z(n3893) );
  IV U3887 ( .A(n3738), .Z(n3898) );
  XOR U3888 ( .A(n3899), .B(n3900), .Z(n3738) );
  AND U3889 ( .A(n175), .B(n3901), .Z(n3900) );
  XOR U3890 ( .A(n3902), .B(n3903), .Z(n3876) );
  AND U3891 ( .A(n3904), .B(n3905), .Z(n3903) );
  XNOR U3892 ( .A(n3810), .B(n3902), .Z(n3905) );
  XNOR U3893 ( .A(n3906), .B(n3907), .Z(n3810) );
  AND U3894 ( .A(n167), .B(n3908), .Z(n3907) );
  XNOR U3895 ( .A(n3909), .B(n3906), .Z(n3908) );
  XOR U3896 ( .A(n3902), .B(n3749), .Z(n3904) );
  XOR U3897 ( .A(n3910), .B(n3911), .Z(n3749) );
  AND U3898 ( .A(n175), .B(n3912), .Z(n3911) );
  XOR U3899 ( .A(n3913), .B(n3914), .Z(n3902) );
  AND U3900 ( .A(n3915), .B(n3916), .Z(n3914) );
  XNOR U3901 ( .A(n3913), .B(n3858), .Z(n3916) );
  XNOR U3902 ( .A(n3917), .B(n3918), .Z(n3858) );
  AND U3903 ( .A(n167), .B(n3919), .Z(n3918) );
  XOR U3904 ( .A(n3920), .B(n3917), .Z(n3919) );
  XNOR U3905 ( .A(n3921), .B(n3913), .Z(n3915) );
  IV U3906 ( .A(n3761), .Z(n3921) );
  XOR U3907 ( .A(n3922), .B(n3923), .Z(n3761) );
  AND U3908 ( .A(n175), .B(n3924), .Z(n3923) );
  AND U3909 ( .A(n3880), .B(n3869), .Z(n3913) );
  XNOR U3910 ( .A(n3925), .B(n3926), .Z(n3869) );
  AND U3911 ( .A(n167), .B(n3927), .Z(n3926) );
  XNOR U3912 ( .A(n3928), .B(n3925), .Z(n3927) );
  XNOR U3913 ( .A(n3929), .B(n3930), .Z(n167) );
  NOR U3914 ( .A(n3931), .B(n3932), .Z(n3930) );
  XNOR U3915 ( .A(n3929), .B(n3891), .Z(n3932) );
  NOR U3916 ( .A(n3887), .B(n3888), .Z(n3891) );
  NOR U3917 ( .A(n3929), .B(n3890), .Z(n3931) );
  AND U3918 ( .A(n3933), .B(n3934), .Z(n3890) );
  XOR U3919 ( .A(n3935), .B(n3936), .Z(n3929) );
  AND U3920 ( .A(n3937), .B(n3938), .Z(n3936) );
  XNOR U3921 ( .A(n3935), .B(n3933), .Z(n3938) );
  IV U3922 ( .A(n3897), .Z(n3933) );
  XOR U3923 ( .A(n3939), .B(n3940), .Z(n3897) );
  XOR U3924 ( .A(n3941), .B(n3934), .Z(n3940) );
  AND U3925 ( .A(n3909), .B(n3942), .Z(n3934) );
  AND U3926 ( .A(n3943), .B(n3944), .Z(n3941) );
  XOR U3927 ( .A(n3945), .B(n3939), .Z(n3943) );
  XNOR U3928 ( .A(n3894), .B(n3935), .Z(n3937) );
  XNOR U3929 ( .A(n3946), .B(n3947), .Z(n3894) );
  AND U3930 ( .A(n171), .B(n3901), .Z(n3947) );
  XOR U3931 ( .A(n3946), .B(n3899), .Z(n3901) );
  XOR U3932 ( .A(n3948), .B(n3949), .Z(n3935) );
  AND U3933 ( .A(n3950), .B(n3951), .Z(n3949) );
  XNOR U3934 ( .A(n3948), .B(n3909), .Z(n3951) );
  XOR U3935 ( .A(n3952), .B(n3944), .Z(n3909) );
  XNOR U3936 ( .A(n3953), .B(n3939), .Z(n3944) );
  XOR U3937 ( .A(n3954), .B(n3955), .Z(n3939) );
  AND U3938 ( .A(n3956), .B(n3957), .Z(n3955) );
  XOR U3939 ( .A(n3958), .B(n3954), .Z(n3956) );
  XNOR U3940 ( .A(n3959), .B(n3960), .Z(n3953) );
  AND U3941 ( .A(n3961), .B(n3962), .Z(n3960) );
  XOR U3942 ( .A(n3959), .B(n3963), .Z(n3961) );
  XNOR U3943 ( .A(n3945), .B(n3942), .Z(n3952) );
  AND U3944 ( .A(n3964), .B(n3965), .Z(n3942) );
  XOR U3945 ( .A(n3966), .B(n3967), .Z(n3945) );
  AND U3946 ( .A(n3968), .B(n3969), .Z(n3967) );
  XOR U3947 ( .A(n3966), .B(n3970), .Z(n3968) );
  XNOR U3948 ( .A(n3906), .B(n3948), .Z(n3950) );
  XNOR U3949 ( .A(n3971), .B(n3972), .Z(n3906) );
  AND U3950 ( .A(n171), .B(n3912), .Z(n3972) );
  XOR U3951 ( .A(n3971), .B(n3910), .Z(n3912) );
  XOR U3952 ( .A(n3973), .B(n3974), .Z(n3948) );
  AND U3953 ( .A(n3975), .B(n3976), .Z(n3974) );
  XNOR U3954 ( .A(n3973), .B(n3964), .Z(n3976) );
  IV U3955 ( .A(n3920), .Z(n3964) );
  XNOR U3956 ( .A(n3977), .B(n3957), .Z(n3920) );
  XNOR U3957 ( .A(n3978), .B(n3963), .Z(n3957) );
  XNOR U3958 ( .A(n3979), .B(n3980), .Z(n3963) );
  NOR U3959 ( .A(n3981), .B(n3982), .Z(n3980) );
  XOR U3960 ( .A(n3979), .B(n3983), .Z(n3981) );
  XNOR U3961 ( .A(n3962), .B(n3954), .Z(n3978) );
  XOR U3962 ( .A(n3984), .B(n3985), .Z(n3954) );
  AND U3963 ( .A(n3986), .B(n3987), .Z(n3985) );
  XOR U3964 ( .A(n3984), .B(n3988), .Z(n3986) );
  XNOR U3965 ( .A(n3989), .B(n3959), .Z(n3962) );
  XOR U3966 ( .A(n3990), .B(n3991), .Z(n3959) );
  AND U3967 ( .A(n3992), .B(n3993), .Z(n3991) );
  XNOR U3968 ( .A(n3994), .B(n3995), .Z(n3992) );
  IV U3969 ( .A(n3990), .Z(n3994) );
  XNOR U3970 ( .A(n3996), .B(n3997), .Z(n3989) );
  NOR U3971 ( .A(n3998), .B(n3999), .Z(n3997) );
  XNOR U3972 ( .A(n3996), .B(n4000), .Z(n3998) );
  XNOR U3973 ( .A(n3958), .B(n3965), .Z(n3977) );
  NOR U3974 ( .A(n3928), .B(n4001), .Z(n3965) );
  XOR U3975 ( .A(n3970), .B(n3969), .Z(n3958) );
  XNOR U3976 ( .A(n4002), .B(n3966), .Z(n3969) );
  XOR U3977 ( .A(n4003), .B(n4004), .Z(n3966) );
  AND U3978 ( .A(n4005), .B(n4006), .Z(n4004) );
  XNOR U3979 ( .A(n4007), .B(n4008), .Z(n4005) );
  IV U3980 ( .A(n4003), .Z(n4007) );
  XNOR U3981 ( .A(n4009), .B(n4010), .Z(n4002) );
  NOR U3982 ( .A(n4011), .B(n4012), .Z(n4010) );
  XNOR U3983 ( .A(n4009), .B(n4013), .Z(n4011) );
  XOR U3984 ( .A(n4014), .B(n4015), .Z(n3970) );
  NOR U3985 ( .A(n4016), .B(n4017), .Z(n4015) );
  XNOR U3986 ( .A(n4014), .B(n4018), .Z(n4016) );
  XNOR U3987 ( .A(n3917), .B(n3973), .Z(n3975) );
  XNOR U3988 ( .A(n4019), .B(n4020), .Z(n3917) );
  AND U3989 ( .A(n171), .B(n3924), .Z(n4020) );
  XOR U3990 ( .A(n4019), .B(n3922), .Z(n3924) );
  AND U3991 ( .A(n3925), .B(n3928), .Z(n3973) );
  XOR U3992 ( .A(n4021), .B(n4001), .Z(n3928) );
  XNOR U3993 ( .A(p_input[192]), .B(p_input[256]), .Z(n4001) );
  XNOR U3994 ( .A(n3988), .B(n3987), .Z(n4021) );
  XNOR U3995 ( .A(n4022), .B(n3995), .Z(n3987) );
  XNOR U3996 ( .A(n3983), .B(n3982), .Z(n3995) );
  XNOR U3997 ( .A(n4023), .B(n3979), .Z(n3982) );
  XNOR U3998 ( .A(p_input[202]), .B(p_input[266]), .Z(n3979) );
  XOR U3999 ( .A(p_input[203]), .B(n2060), .Z(n4023) );
  XOR U4000 ( .A(p_input[204]), .B(p_input[268]), .Z(n3983) );
  XOR U4001 ( .A(n3993), .B(n4024), .Z(n4022) );
  IV U4002 ( .A(n3984), .Z(n4024) );
  XOR U4003 ( .A(p_input[193]), .B(p_input[257]), .Z(n3984) );
  XNOR U4004 ( .A(n4025), .B(n4000), .Z(n3993) );
  XNOR U4005 ( .A(p_input[207]), .B(n2063), .Z(n4000) );
  XOR U4006 ( .A(n3990), .B(n3999), .Z(n4025) );
  XOR U4007 ( .A(n4026), .B(n3996), .Z(n3999) );
  XOR U4008 ( .A(p_input[205]), .B(p_input[269]), .Z(n3996) );
  XOR U4009 ( .A(p_input[206]), .B(n2065), .Z(n4026) );
  XOR U4010 ( .A(p_input[201]), .B(p_input[265]), .Z(n3990) );
  XOR U4011 ( .A(n4008), .B(n4006), .Z(n3988) );
  XNOR U4012 ( .A(n4027), .B(n4013), .Z(n4006) );
  XOR U4013 ( .A(p_input[200]), .B(p_input[264]), .Z(n4013) );
  XOR U4014 ( .A(n4003), .B(n4012), .Z(n4027) );
  XOR U4015 ( .A(n4028), .B(n4009), .Z(n4012) );
  XOR U4016 ( .A(p_input[198]), .B(p_input[262]), .Z(n4009) );
  XOR U4017 ( .A(p_input[199]), .B(n2239), .Z(n4028) );
  XOR U4018 ( .A(p_input[194]), .B(p_input[258]), .Z(n4003) );
  XNOR U4019 ( .A(n4018), .B(n4017), .Z(n4008) );
  XOR U4020 ( .A(n4029), .B(n4014), .Z(n4017) );
  XOR U4021 ( .A(p_input[195]), .B(p_input[259]), .Z(n4014) );
  XOR U4022 ( .A(p_input[196]), .B(n2241), .Z(n4029) );
  XOR U4023 ( .A(p_input[197]), .B(p_input[261]), .Z(n4018) );
  XNOR U4024 ( .A(n4030), .B(n4031), .Z(n3925) );
  AND U4025 ( .A(n171), .B(n4032), .Z(n4031) );
  XNOR U4026 ( .A(n4033), .B(n4034), .Z(n171) );
  NOR U4027 ( .A(n4035), .B(n4036), .Z(n4034) );
  XOR U4028 ( .A(n3888), .B(n4033), .Z(n4036) );
  NOR U4029 ( .A(n4033), .B(n3887), .Z(n4035) );
  XOR U4030 ( .A(n4037), .B(n4038), .Z(n4033) );
  AND U4031 ( .A(n4039), .B(n4040), .Z(n4038) );
  XOR U4032 ( .A(n4037), .B(n3899), .Z(n4039) );
  XOR U4033 ( .A(n4041), .B(n4042), .Z(n3880) );
  AND U4034 ( .A(n175), .B(n4032), .Z(n4042) );
  XNOR U4035 ( .A(n4030), .B(n4041), .Z(n4032) );
  XNOR U4036 ( .A(n4043), .B(n4044), .Z(n175) );
  NOR U4037 ( .A(n4045), .B(n4046), .Z(n4044) );
  XNOR U4038 ( .A(n3888), .B(n4047), .Z(n4046) );
  IV U4039 ( .A(n4043), .Z(n4047) );
  AND U4040 ( .A(n4048), .B(n4049), .Z(n3888) );
  NOR U4041 ( .A(n4043), .B(n3887), .Z(n4045) );
  AND U4042 ( .A(n4050), .B(n4051), .Z(n3887) );
  IV U4043 ( .A(n4052), .Z(n4050) );
  XOR U4044 ( .A(n4037), .B(n4053), .Z(n4043) );
  AND U4045 ( .A(n4054), .B(n4040), .Z(n4053) );
  XNOR U4046 ( .A(n3946), .B(n4037), .Z(n4040) );
  XNOR U4047 ( .A(n4055), .B(n4056), .Z(n3946) );
  AND U4048 ( .A(n178), .B(n4057), .Z(n4056) );
  XOR U4049 ( .A(n4058), .B(n4055), .Z(n4057) );
  XNOR U4050 ( .A(n4059), .B(n4037), .Z(n4054) );
  IV U4051 ( .A(n3899), .Z(n4059) );
  XOR U4052 ( .A(n4060), .B(n4061), .Z(n3899) );
  AND U4053 ( .A(n185), .B(n4062), .Z(n4061) );
  XOR U4054 ( .A(n4063), .B(n4064), .Z(n4037) );
  AND U4055 ( .A(n4065), .B(n4066), .Z(n4064) );
  XNOR U4056 ( .A(n3971), .B(n4063), .Z(n4066) );
  XNOR U4057 ( .A(n4067), .B(n4068), .Z(n3971) );
  AND U4058 ( .A(n178), .B(n4069), .Z(n4068) );
  XNOR U4059 ( .A(n4070), .B(n4067), .Z(n4069) );
  XOR U4060 ( .A(n4063), .B(n3910), .Z(n4065) );
  XOR U4061 ( .A(n4071), .B(n4072), .Z(n3910) );
  AND U4062 ( .A(n185), .B(n4073), .Z(n4072) );
  XOR U4063 ( .A(n4074), .B(n4075), .Z(n4063) );
  AND U4064 ( .A(n4076), .B(n4077), .Z(n4075) );
  XNOR U4065 ( .A(n4074), .B(n4019), .Z(n4077) );
  XNOR U4066 ( .A(n4078), .B(n4079), .Z(n4019) );
  AND U4067 ( .A(n178), .B(n4080), .Z(n4079) );
  XOR U4068 ( .A(n4081), .B(n4078), .Z(n4080) );
  XNOR U4069 ( .A(n4082), .B(n4074), .Z(n4076) );
  IV U4070 ( .A(n3922), .Z(n4082) );
  XOR U4071 ( .A(n4083), .B(n4084), .Z(n3922) );
  AND U4072 ( .A(n185), .B(n4085), .Z(n4084) );
  AND U4073 ( .A(n4041), .B(n4030), .Z(n4074) );
  XNOR U4074 ( .A(n4086), .B(n4087), .Z(n4030) );
  AND U4075 ( .A(n178), .B(n4088), .Z(n4087) );
  XNOR U4076 ( .A(n4089), .B(n4086), .Z(n4088) );
  XNOR U4077 ( .A(n4090), .B(n4091), .Z(n178) );
  NOR U4078 ( .A(n4092), .B(n4093), .Z(n4091) );
  XNOR U4079 ( .A(n4090), .B(n4052), .Z(n4093) );
  NOR U4080 ( .A(n4048), .B(n4049), .Z(n4052) );
  NOR U4081 ( .A(n4090), .B(n4051), .Z(n4092) );
  AND U4082 ( .A(n4094), .B(n4095), .Z(n4051) );
  XOR U4083 ( .A(n4096), .B(n4097), .Z(n4090) );
  AND U4084 ( .A(n4098), .B(n4099), .Z(n4097) );
  XNOR U4085 ( .A(n4096), .B(n4094), .Z(n4099) );
  IV U4086 ( .A(n4058), .Z(n4094) );
  XOR U4087 ( .A(n4100), .B(n4101), .Z(n4058) );
  XOR U4088 ( .A(n4102), .B(n4095), .Z(n4101) );
  AND U4089 ( .A(n4070), .B(n4103), .Z(n4095) );
  AND U4090 ( .A(n4104), .B(n4105), .Z(n4102) );
  XOR U4091 ( .A(n4106), .B(n4100), .Z(n4104) );
  XNOR U4092 ( .A(n4055), .B(n4096), .Z(n4098) );
  XNOR U4093 ( .A(n4107), .B(n4108), .Z(n4055) );
  AND U4094 ( .A(n182), .B(n4062), .Z(n4108) );
  XOR U4095 ( .A(n4107), .B(n4060), .Z(n4062) );
  XOR U4096 ( .A(n4109), .B(n4110), .Z(n4096) );
  AND U4097 ( .A(n4111), .B(n4112), .Z(n4110) );
  XNOR U4098 ( .A(n4109), .B(n4070), .Z(n4112) );
  XOR U4099 ( .A(n4113), .B(n4105), .Z(n4070) );
  XNOR U4100 ( .A(n4114), .B(n4100), .Z(n4105) );
  XOR U4101 ( .A(n4115), .B(n4116), .Z(n4100) );
  AND U4102 ( .A(n4117), .B(n4118), .Z(n4116) );
  XOR U4103 ( .A(n4119), .B(n4115), .Z(n4117) );
  XNOR U4104 ( .A(n4120), .B(n4121), .Z(n4114) );
  AND U4105 ( .A(n4122), .B(n4123), .Z(n4121) );
  XOR U4106 ( .A(n4120), .B(n4124), .Z(n4122) );
  XNOR U4107 ( .A(n4106), .B(n4103), .Z(n4113) );
  AND U4108 ( .A(n4125), .B(n4126), .Z(n4103) );
  XOR U4109 ( .A(n4127), .B(n4128), .Z(n4106) );
  AND U4110 ( .A(n4129), .B(n4130), .Z(n4128) );
  XOR U4111 ( .A(n4127), .B(n4131), .Z(n4129) );
  XNOR U4112 ( .A(n4067), .B(n4109), .Z(n4111) );
  XNOR U4113 ( .A(n4132), .B(n4133), .Z(n4067) );
  AND U4114 ( .A(n182), .B(n4073), .Z(n4133) );
  XOR U4115 ( .A(n4132), .B(n4071), .Z(n4073) );
  XOR U4116 ( .A(n4134), .B(n4135), .Z(n4109) );
  AND U4117 ( .A(n4136), .B(n4137), .Z(n4135) );
  XNOR U4118 ( .A(n4134), .B(n4125), .Z(n4137) );
  IV U4119 ( .A(n4081), .Z(n4125) );
  XNOR U4120 ( .A(n4138), .B(n4118), .Z(n4081) );
  XNOR U4121 ( .A(n4139), .B(n4124), .Z(n4118) );
  XNOR U4122 ( .A(n4140), .B(n4141), .Z(n4124) );
  NOR U4123 ( .A(n4142), .B(n4143), .Z(n4141) );
  XOR U4124 ( .A(n4140), .B(n4144), .Z(n4142) );
  XNOR U4125 ( .A(n4123), .B(n4115), .Z(n4139) );
  XOR U4126 ( .A(n4145), .B(n4146), .Z(n4115) );
  AND U4127 ( .A(n4147), .B(n4148), .Z(n4146) );
  XOR U4128 ( .A(n4145), .B(n4149), .Z(n4147) );
  XNOR U4129 ( .A(n4150), .B(n4120), .Z(n4123) );
  XOR U4130 ( .A(n4151), .B(n4152), .Z(n4120) );
  AND U4131 ( .A(n4153), .B(n4154), .Z(n4152) );
  XNOR U4132 ( .A(n4155), .B(n4156), .Z(n4153) );
  IV U4133 ( .A(n4151), .Z(n4155) );
  XNOR U4134 ( .A(n4157), .B(n4158), .Z(n4150) );
  NOR U4135 ( .A(n4159), .B(n4160), .Z(n4158) );
  XNOR U4136 ( .A(n4157), .B(n4161), .Z(n4159) );
  XNOR U4137 ( .A(n4119), .B(n4126), .Z(n4138) );
  NOR U4138 ( .A(n4089), .B(n4162), .Z(n4126) );
  XOR U4139 ( .A(n4131), .B(n4130), .Z(n4119) );
  XNOR U4140 ( .A(n4163), .B(n4127), .Z(n4130) );
  XOR U4141 ( .A(n4164), .B(n4165), .Z(n4127) );
  AND U4142 ( .A(n4166), .B(n4167), .Z(n4165) );
  XNOR U4143 ( .A(n4168), .B(n4169), .Z(n4166) );
  IV U4144 ( .A(n4164), .Z(n4168) );
  XNOR U4145 ( .A(n4170), .B(n4171), .Z(n4163) );
  NOR U4146 ( .A(n4172), .B(n4173), .Z(n4171) );
  XNOR U4147 ( .A(n4170), .B(n4174), .Z(n4172) );
  XOR U4148 ( .A(n4175), .B(n4176), .Z(n4131) );
  NOR U4149 ( .A(n4177), .B(n4178), .Z(n4176) );
  XNOR U4150 ( .A(n4175), .B(n4179), .Z(n4177) );
  XNOR U4151 ( .A(n4078), .B(n4134), .Z(n4136) );
  XNOR U4152 ( .A(n4180), .B(n4181), .Z(n4078) );
  AND U4153 ( .A(n182), .B(n4085), .Z(n4181) );
  XOR U4154 ( .A(n4180), .B(n4083), .Z(n4085) );
  AND U4155 ( .A(n4086), .B(n4089), .Z(n4134) );
  XOR U4156 ( .A(n4182), .B(n4162), .Z(n4089) );
  XNOR U4157 ( .A(p_input[208]), .B(p_input[256]), .Z(n4162) );
  XNOR U4158 ( .A(n4149), .B(n4148), .Z(n4182) );
  XNOR U4159 ( .A(n4183), .B(n4156), .Z(n4148) );
  XNOR U4160 ( .A(n4144), .B(n4143), .Z(n4156) );
  XNOR U4161 ( .A(n4184), .B(n4140), .Z(n4143) );
  XNOR U4162 ( .A(p_input[218]), .B(p_input[266]), .Z(n4140) );
  XOR U4163 ( .A(p_input[219]), .B(n2060), .Z(n4184) );
  XOR U4164 ( .A(p_input[220]), .B(p_input[268]), .Z(n4144) );
  XOR U4165 ( .A(n4154), .B(n4185), .Z(n4183) );
  IV U4166 ( .A(n4145), .Z(n4185) );
  XOR U4167 ( .A(p_input[209]), .B(p_input[257]), .Z(n4145) );
  XNOR U4168 ( .A(n4186), .B(n4161), .Z(n4154) );
  XNOR U4169 ( .A(p_input[223]), .B(n2063), .Z(n4161) );
  IV U4170 ( .A(p_input[271]), .Z(n2063) );
  XOR U4171 ( .A(n4151), .B(n4160), .Z(n4186) );
  XOR U4172 ( .A(n4187), .B(n4157), .Z(n4160) );
  XOR U4173 ( .A(p_input[221]), .B(p_input[269]), .Z(n4157) );
  XOR U4174 ( .A(p_input[222]), .B(n2065), .Z(n4187) );
  XOR U4175 ( .A(p_input[217]), .B(p_input[265]), .Z(n4151) );
  XOR U4176 ( .A(n4169), .B(n4167), .Z(n4149) );
  XNOR U4177 ( .A(n4188), .B(n4174), .Z(n4167) );
  XOR U4178 ( .A(p_input[216]), .B(p_input[264]), .Z(n4174) );
  XOR U4179 ( .A(n4164), .B(n4173), .Z(n4188) );
  XOR U4180 ( .A(n4189), .B(n4170), .Z(n4173) );
  XOR U4181 ( .A(p_input[214]), .B(p_input[262]), .Z(n4170) );
  XOR U4182 ( .A(p_input[215]), .B(n2239), .Z(n4189) );
  XOR U4183 ( .A(p_input[210]), .B(p_input[258]), .Z(n4164) );
  XNOR U4184 ( .A(n4179), .B(n4178), .Z(n4169) );
  XOR U4185 ( .A(n4190), .B(n4175), .Z(n4178) );
  XOR U4186 ( .A(p_input[211]), .B(p_input[259]), .Z(n4175) );
  XOR U4187 ( .A(p_input[212]), .B(n2241), .Z(n4190) );
  XOR U4188 ( .A(p_input[213]), .B(p_input[261]), .Z(n4179) );
  XNOR U4189 ( .A(n4191), .B(n4192), .Z(n4086) );
  AND U4190 ( .A(n182), .B(n4193), .Z(n4192) );
  XNOR U4191 ( .A(n4194), .B(n4195), .Z(n182) );
  NOR U4192 ( .A(n4196), .B(n4197), .Z(n4195) );
  XOR U4193 ( .A(n4049), .B(n4194), .Z(n4197) );
  NOR U4194 ( .A(n4194), .B(n4048), .Z(n4196) );
  XOR U4195 ( .A(n4198), .B(n4199), .Z(n4194) );
  AND U4196 ( .A(n4200), .B(n4201), .Z(n4199) );
  XOR U4197 ( .A(n4198), .B(n4060), .Z(n4200) );
  XOR U4198 ( .A(n4202), .B(n4203), .Z(n4041) );
  AND U4199 ( .A(n185), .B(n4193), .Z(n4203) );
  XOR U4200 ( .A(n4204), .B(n4202), .Z(n4193) );
  XNOR U4201 ( .A(n4205), .B(n4206), .Z(n185) );
  NOR U4202 ( .A(n4207), .B(n4208), .Z(n4206) );
  XNOR U4203 ( .A(n4049), .B(n4209), .Z(n4208) );
  IV U4204 ( .A(n4205), .Z(n4209) );
  AND U4205 ( .A(n4060), .B(n4210), .Z(n4049) );
  NOR U4206 ( .A(n4205), .B(n4048), .Z(n4207) );
  AND U4207 ( .A(n4107), .B(n4211), .Z(n4048) );
  XOR U4208 ( .A(n4198), .B(n4212), .Z(n4205) );
  AND U4209 ( .A(n4213), .B(n4201), .Z(n4212) );
  XNOR U4210 ( .A(n4107), .B(n4198), .Z(n4201) );
  XNOR U4211 ( .A(n4214), .B(n4215), .Z(n4107) );
  XOR U4212 ( .A(n4216), .B(n4211), .Z(n4215) );
  AND U4213 ( .A(n4132), .B(n4217), .Z(n4211) );
  AND U4214 ( .A(n4218), .B(n4219), .Z(n4216) );
  XOR U4215 ( .A(n4220), .B(n4214), .Z(n4218) );
  XNOR U4216 ( .A(n4221), .B(n4198), .Z(n4213) );
  IV U4217 ( .A(n4060), .Z(n4221) );
  XNOR U4218 ( .A(n4222), .B(n4223), .Z(n4060) );
  XOR U4219 ( .A(n4224), .B(n4210), .Z(n4223) );
  AND U4220 ( .A(n4071), .B(n4225), .Z(n4210) );
  AND U4221 ( .A(n4226), .B(n4227), .Z(n4224) );
  XNOR U4222 ( .A(n4222), .B(n4228), .Z(n4226) );
  XOR U4223 ( .A(n4229), .B(n4230), .Z(n4198) );
  AND U4224 ( .A(n4231), .B(n4232), .Z(n4230) );
  XNOR U4225 ( .A(n4132), .B(n4229), .Z(n4232) );
  XOR U4226 ( .A(n4233), .B(n4219), .Z(n4132) );
  XNOR U4227 ( .A(n4234), .B(n4214), .Z(n4219) );
  XOR U4228 ( .A(n4235), .B(n4236), .Z(n4214) );
  AND U4229 ( .A(n4237), .B(n4238), .Z(n4236) );
  XOR U4230 ( .A(n4239), .B(n4235), .Z(n4237) );
  XNOR U4231 ( .A(n4240), .B(n4241), .Z(n4234) );
  AND U4232 ( .A(n4242), .B(n4243), .Z(n4241) );
  XOR U4233 ( .A(n4240), .B(n4244), .Z(n4242) );
  XNOR U4234 ( .A(n4220), .B(n4217), .Z(n4233) );
  AND U4235 ( .A(n4180), .B(n4245), .Z(n4217) );
  XOR U4236 ( .A(n4246), .B(n4247), .Z(n4220) );
  AND U4237 ( .A(n4248), .B(n4249), .Z(n4247) );
  XOR U4238 ( .A(n4246), .B(n4250), .Z(n4248) );
  XOR U4239 ( .A(n4229), .B(n4071), .Z(n4231) );
  XNOR U4240 ( .A(n4251), .B(n4228), .Z(n4071) );
  XNOR U4241 ( .A(n4252), .B(n4253), .Z(n4228) );
  AND U4242 ( .A(n4254), .B(n4255), .Z(n4253) );
  XOR U4243 ( .A(n4252), .B(n4256), .Z(n4254) );
  XNOR U4244 ( .A(n4227), .B(n4225), .Z(n4251) );
  AND U4245 ( .A(n4083), .B(n4257), .Z(n4225) );
  XNOR U4246 ( .A(n4258), .B(n4222), .Z(n4227) );
  XOR U4247 ( .A(n4259), .B(n4260), .Z(n4222) );
  AND U4248 ( .A(n4261), .B(n4262), .Z(n4260) );
  XOR U4249 ( .A(n4259), .B(n4263), .Z(n4261) );
  XNOR U4250 ( .A(n4264), .B(n4265), .Z(n4258) );
  AND U4251 ( .A(n4266), .B(n4267), .Z(n4265) );
  XNOR U4252 ( .A(n4264), .B(n4268), .Z(n4266) );
  XOR U4253 ( .A(n4269), .B(n4270), .Z(n4229) );
  AND U4254 ( .A(n4271), .B(n4272), .Z(n4270) );
  XNOR U4255 ( .A(n4269), .B(n4180), .Z(n4272) );
  XOR U4256 ( .A(n4273), .B(n4238), .Z(n4180) );
  XNOR U4257 ( .A(n4274), .B(n4244), .Z(n4238) );
  XOR U4258 ( .A(n4275), .B(n4276), .Z(n4244) );
  NOR U4259 ( .A(n4277), .B(n4278), .Z(n4276) );
  XNOR U4260 ( .A(n4275), .B(n4279), .Z(n4277) );
  XNOR U4261 ( .A(n4243), .B(n4235), .Z(n4274) );
  XOR U4262 ( .A(n4280), .B(n4281), .Z(n4235) );
  AND U4263 ( .A(n4282), .B(n4283), .Z(n4281) );
  XNOR U4264 ( .A(n4280), .B(n4284), .Z(n4282) );
  XNOR U4265 ( .A(n4285), .B(n4240), .Z(n4243) );
  XOR U4266 ( .A(n4286), .B(n4287), .Z(n4240) );
  AND U4267 ( .A(n4288), .B(n4289), .Z(n4287) );
  XOR U4268 ( .A(n4286), .B(n4290), .Z(n4288) );
  XNOR U4269 ( .A(n4291), .B(n4292), .Z(n4285) );
  NOR U4270 ( .A(n4293), .B(n4294), .Z(n4292) );
  XOR U4271 ( .A(n4291), .B(n4295), .Z(n4293) );
  XNOR U4272 ( .A(n4239), .B(n4245), .Z(n4273) );
  AND U4273 ( .A(n4204), .B(n4296), .Z(n4245) );
  IV U4274 ( .A(n4191), .Z(n4204) );
  XOR U4275 ( .A(n4250), .B(n4249), .Z(n4239) );
  XNOR U4276 ( .A(n4297), .B(n4246), .Z(n4249) );
  XOR U4277 ( .A(n4298), .B(n4299), .Z(n4246) );
  AND U4278 ( .A(n4300), .B(n4301), .Z(n4299) );
  XOR U4279 ( .A(n4298), .B(n4302), .Z(n4300) );
  XNOR U4280 ( .A(n4303), .B(n4304), .Z(n4297) );
  NOR U4281 ( .A(n4305), .B(n4306), .Z(n4304) );
  XNOR U4282 ( .A(n4303), .B(n4307), .Z(n4305) );
  XOR U4283 ( .A(n4308), .B(n4309), .Z(n4250) );
  NOR U4284 ( .A(n4310), .B(n4311), .Z(n4309) );
  XNOR U4285 ( .A(n4308), .B(n4312), .Z(n4310) );
  XNOR U4286 ( .A(n4313), .B(n4269), .Z(n4271) );
  IV U4287 ( .A(n4083), .Z(n4313) );
  XOR U4288 ( .A(n4314), .B(n4263), .Z(n4083) );
  XOR U4289 ( .A(n4256), .B(n4255), .Z(n4263) );
  XNOR U4290 ( .A(n4315), .B(n4252), .Z(n4255) );
  XOR U4291 ( .A(n4316), .B(n4317), .Z(n4252) );
  AND U4292 ( .A(n4318), .B(n4319), .Z(n4317) );
  XOR U4293 ( .A(n4316), .B(n4320), .Z(n4318) );
  XNOR U4294 ( .A(n4321), .B(n4322), .Z(n4315) );
  NOR U4295 ( .A(n4323), .B(n4324), .Z(n4322) );
  XNOR U4296 ( .A(n4321), .B(n4325), .Z(n4323) );
  XOR U4297 ( .A(n4326), .B(n4327), .Z(n4256) );
  NOR U4298 ( .A(n4328), .B(n4329), .Z(n4327) );
  XNOR U4299 ( .A(n4326), .B(n4330), .Z(n4328) );
  XNOR U4300 ( .A(n4262), .B(n4257), .Z(n4314) );
  AND U4301 ( .A(n4202), .B(n4331), .Z(n4257) );
  XOR U4302 ( .A(n4332), .B(n4268), .Z(n4262) );
  XNOR U4303 ( .A(n4333), .B(n4334), .Z(n4268) );
  NOR U4304 ( .A(n4335), .B(n4336), .Z(n4334) );
  XNOR U4305 ( .A(n4333), .B(n4337), .Z(n4335) );
  XNOR U4306 ( .A(n4267), .B(n4259), .Z(n4332) );
  XOR U4307 ( .A(n4338), .B(n4339), .Z(n4259) );
  AND U4308 ( .A(n4340), .B(n4341), .Z(n4339) );
  XOR U4309 ( .A(n4338), .B(n4342), .Z(n4340) );
  XNOR U4310 ( .A(n4343), .B(n4264), .Z(n4267) );
  XOR U4311 ( .A(n4344), .B(n4345), .Z(n4264) );
  AND U4312 ( .A(n4346), .B(n4347), .Z(n4345) );
  XOR U4313 ( .A(n4344), .B(n4348), .Z(n4346) );
  XNOR U4314 ( .A(n4349), .B(n4350), .Z(n4343) );
  NOR U4315 ( .A(n4351), .B(n4352), .Z(n4350) );
  XOR U4316 ( .A(n4349), .B(n4353), .Z(n4351) );
  AND U4317 ( .A(n4202), .B(n4191), .Z(n4269) );
  XNOR U4318 ( .A(n4354), .B(n4296), .Z(n4191) );
  XOR U4319 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(
        p_input[256]), .Z(n4296) );
  XOR U4320 ( .A(n4284), .B(n4283), .Z(n4354) );
  XNOR U4321 ( .A(n4355), .B(n4290), .Z(n4283) );
  XNOR U4322 ( .A(n4279), .B(n4278), .Z(n4290) );
  XOR U4323 ( .A(n4356), .B(n4275), .Z(n4278) );
  XNOR U4324 ( .A(n1790), .B(p_input[266]), .Z(n4275) );
  IV U4325 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n1790) );
  XOR U4326 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n2060), 
        .Z(n4356) );
  XNOR U4327 ( .A(n1563), .B(p_input[268]), .Z(n4279) );
  IV U4328 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n1563) );
  XNOR U4329 ( .A(n4289), .B(n4280), .Z(n4355) );
  XNOR U4330 ( .A(n1104), .B(p_input[257]), .Z(n4280) );
  IV U4331 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n1104) );
  XOR U4332 ( .A(n4357), .B(n4295), .Z(n4289) );
  XNOR U4333 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(
        p_input[271]), .Z(n4295) );
  XOR U4334 ( .A(n4286), .B(n4294), .Z(n4357) );
  XOR U4335 ( .A(n4358), .B(n4291), .Z(n4294) );
  XNOR U4336 ( .A(n1450), .B(p_input[269]), .Z(n4291) );
  IV U4337 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n1450) );
  XOR U4338 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(n2065), 
        .Z(n4358) );
  XNOR U4339 ( .A(n180), .B(p_input[265]), .Z(n4286) );
  IV U4340 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .Z(n180) );
  XNOR U4341 ( .A(n4302), .B(n4301), .Z(n4284) );
  XNOR U4342 ( .A(n4359), .B(n4307), .Z(n4301) );
  XNOR U4343 ( .A(n297), .B(p_input[264]), .Z(n4307) );
  IV U4344 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .Z(n297) );
  XOR U4345 ( .A(n4298), .B(n4306), .Z(n4359) );
  XOR U4346 ( .A(n4360), .B(n4303), .Z(n4306) );
  XNOR U4347 ( .A(n527), .B(p_input[262]), .Z(n4303) );
  IV U4348 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .Z(n527) );
  XOR U4349 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(n2239), 
        .Z(n4360) );
  XNOR U4350 ( .A(n989), .B(p_input[258]), .Z(n4298) );
  IV U4351 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n989) );
  XNOR U4352 ( .A(n4312), .B(n4311), .Z(n4302) );
  XOR U4353 ( .A(n4361), .B(n4308), .Z(n4311) );
  XNOR U4354 ( .A(n874), .B(p_input[259]), .Z(n4308) );
  IV U4355 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .Z(n874) );
  XOR U4356 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(n2241), 
        .Z(n4361) );
  XNOR U4357 ( .A(n642), .B(p_input[261]), .Z(n4312) );
  IV U4358 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .Z(n642) );
  XOR U4359 ( .A(n4362), .B(n4342), .Z(n4202) );
  XOR U4360 ( .A(n4320), .B(n4319), .Z(n4342) );
  XNOR U4361 ( .A(n4363), .B(n4325), .Z(n4319) );
  XNOR U4362 ( .A(n301), .B(p_input[264]), .Z(n4325) );
  IV U4363 ( .A(\knn_comb_/min_val_out[0][8] ), .Z(n301) );
  XOR U4364 ( .A(n4316), .B(n4324), .Z(n4363) );
  XOR U4365 ( .A(n4364), .B(n4321), .Z(n4324) );
  XNOR U4366 ( .A(n531), .B(p_input[262]), .Z(n4321) );
  IV U4367 ( .A(\knn_comb_/min_val_out[0][6] ), .Z(n531) );
  XOR U4368 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n2239), .Z(n4364) );
  IV U4369 ( .A(p_input[263]), .Z(n2239) );
  XNOR U4370 ( .A(n993), .B(p_input[258]), .Z(n4316) );
  IV U4371 ( .A(\knn_comb_/min_val_out[0][2] ), .Z(n993) );
  XNOR U4372 ( .A(n4330), .B(n4329), .Z(n4320) );
  XOR U4373 ( .A(n4365), .B(n4326), .Z(n4329) );
  XNOR U4374 ( .A(n878), .B(p_input[259]), .Z(n4326) );
  IV U4375 ( .A(\knn_comb_/min_val_out[0][3] ), .Z(n878) );
  XOR U4376 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n2241), .Z(n4365) );
  IV U4377 ( .A(p_input[260]), .Z(n2241) );
  XNOR U4378 ( .A(n646), .B(p_input[261]), .Z(n4330) );
  IV U4379 ( .A(\knn_comb_/min_val_out[0][5] ), .Z(n646) );
  XNOR U4380 ( .A(n4341), .B(n4331), .Z(n4362) );
  XOR U4381 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[256]), .Z(n4331)
         );
  XNOR U4382 ( .A(n4366), .B(n4348), .Z(n4341) );
  XNOR U4383 ( .A(n4337), .B(n4336), .Z(n4348) );
  XOR U4384 ( .A(n4367), .B(n4333), .Z(n4336) );
  XNOR U4385 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n2233), .Z(n4333) );
  IV U4386 ( .A(p_input[266]), .Z(n2233) );
  XOR U4387 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n2060), .Z(n4367) );
  IV U4388 ( .A(p_input[267]), .Z(n2060) );
  XOR U4389 ( .A(\knn_comb_/min_val_out[0][12] ), .B(p_input[268]), .Z(n4337)
         );
  XNOR U4390 ( .A(n4347), .B(n4338), .Z(n4366) );
  XNOR U4391 ( .A(n1108), .B(p_input[257]), .Z(n4338) );
  IV U4392 ( .A(\knn_comb_/min_val_out[0][1] ), .Z(n1108) );
  XOR U4393 ( .A(n4368), .B(n4353), .Z(n4347) );
  XNOR U4394 ( .A(\knn_comb_/min_val_out[0][15] ), .B(p_input[271]), .Z(n4353)
         );
  XOR U4395 ( .A(n4344), .B(n4352), .Z(n4368) );
  XOR U4396 ( .A(n4369), .B(n4349), .Z(n4352) );
  XOR U4397 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[269]), .Z(n4349)
         );
  XOR U4398 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n2065), .Z(n4369) );
  IV U4399 ( .A(p_input[270]), .Z(n2065) );
  XNOR U4400 ( .A(n186), .B(p_input[265]), .Z(n4344) );
  IV U4401 ( .A(\knn_comb_/min_val_out[0][9] ), .Z(n186) );
endmodule

