
module knn_comb_BMR_W32_K3_N16 ( p_input, o );
  input [543:0] p_input;
  output [95:0] o;
  wire   \knn_comb_/min_val_out[0][0] , \knn_comb_/min_val_out[0][1] ,
         \knn_comb_/min_val_out[0][2] , \knn_comb_/min_val_out[0][3] ,
         \knn_comb_/min_val_out[0][4] , \knn_comb_/min_val_out[0][5] ,
         \knn_comb_/min_val_out[0][6] , \knn_comb_/min_val_out[0][7] ,
         \knn_comb_/min_val_out[0][8] , \knn_comb_/min_val_out[0][9] ,
         \knn_comb_/min_val_out[0][10] , \knn_comb_/min_val_out[0][11] ,
         \knn_comb_/min_val_out[0][12] , \knn_comb_/min_val_out[0][13] ,
         \knn_comb_/min_val_out[0][14] , \knn_comb_/min_val_out[0][15] ,
         \knn_comb_/min_val_out[0][16] , \knn_comb_/min_val_out[0][17] ,
         \knn_comb_/min_val_out[0][18] , \knn_comb_/min_val_out[0][19] ,
         \knn_comb_/min_val_out[0][20] , \knn_comb_/min_val_out[0][21] ,
         \knn_comb_/min_val_out[0][22] , \knn_comb_/min_val_out[0][23] ,
         \knn_comb_/min_val_out[0][24] , \knn_comb_/min_val_out[0][25] ,
         \knn_comb_/min_val_out[0][26] , \knn_comb_/min_val_out[0][27] ,
         \knn_comb_/min_val_out[0][28] , \knn_comb_/min_val_out[0][29] ,
         \knn_comb_/min_val_out[0][30] , \knn_comb_/min_val_out[0][31] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][16] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][17] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][18] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][19] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][20] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][21] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][22] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][23] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][24] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][25] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][26] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][27] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][28] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][29] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][30] ,
         \knn_comb_/ASN_1[2].knn_/local_min_val[2][31] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ,
         \knn_comb_/ASN_1[1].knn_/local_min_val[1][31] , n1, n2, n3, n4, n5,
         n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444,
         n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454,
         n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464,
         n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474,
         n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483, n2484,
         n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494,
         n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503, n2504,
         n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513, n2514,
         n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523, n2524,
         n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574,
         n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583, n2584,
         n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593, n2594,
         n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603, n2604,
         n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613, n2614,
         n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623, n2624,
         n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634,
         n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644,
         n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654,
         n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674,
         n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684,
         n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694,
         n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704,
         n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714,
         n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724,
         n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734,
         n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744,
         n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754,
         n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764,
         n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774,
         n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784,
         n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814,
         n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824,
         n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834,
         n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844,
         n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854,
         n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864,
         n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874,
         n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884,
         n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894,
         n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904,
         n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914,
         n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944,
         n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954,
         n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964,
         n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974,
         n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984,
         n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994,
         n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064,
         n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074,
         n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084,
         n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094,
         n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104,
         n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114,
         n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124,
         n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134,
         n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144,
         n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154,
         n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164,
         n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174,
         n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184,
         n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194,
         n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204,
         n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214,
         n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224,
         n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234,
         n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244,
         n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254,
         n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264,
         n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274,
         n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284,
         n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294,
         n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304,
         n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314,
         n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324,
         n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334,
         n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344,
         n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354,
         n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364,
         n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374,
         n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384,
         n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394,
         n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404,
         n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414,
         n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424,
         n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434,
         n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444,
         n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454,
         n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464,
         n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474,
         n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484,
         n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494,
         n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504,
         n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514,
         n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764,
         n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774,
         n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784,
         n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794,
         n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804,
         n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814,
         n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824,
         n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834,
         n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844,
         n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854,
         n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864,
         n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874,
         n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884,
         n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894,
         n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903, n3904,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943, n3944,
         n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954,
         n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963, n3964,
         n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973, n3974,
         n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984,
         n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994,
         n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004,
         n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014,
         n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024,
         n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034,
         n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044,
         n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054,
         n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064,
         n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074,
         n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084,
         n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094,
         n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104,
         n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114,
         n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124,
         n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134,
         n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144,
         n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154,
         n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164,
         n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174,
         n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184,
         n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194,
         n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204,
         n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684,
         n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10891,
         n10892, n10893, n10894, n10895, n10896, n10897, n10898, n10899,
         n10900, n10901, n10902, n10903, n10904, n10905, n10906, n10907,
         n10908, n10909, n10910, n10911, n10912, n10913, n10914, n10915,
         n10916, n10917, n10918, n10919, n10920, n10921, n10922, n10923,
         n10924, n10925, n10926, n10927, n10928, n10929, n10930, n10931,
         n10932, n10933, n10934, n10935, n10936, n10937, n10938, n10939,
         n10940, n10941, n10942, n10943, n10944, n10945, n10946, n10947,
         n10948, n10949, n10950, n10951, n10952, n10953, n10954, n10955,
         n10956, n10957, n10958, n10959, n10960, n10961, n10962, n10963,
         n10964, n10965, n10966, n10967, n10968, n10969, n10970, n10971,
         n10972, n10973, n10974, n10975, n10976, n10977, n10978, n10979,
         n10980, n10981, n10982, n10983, n10984, n10985, n10986, n10987,
         n10988, n10989, n10990, n10991, n10992, n10993, n10994, n10995,
         n10996, n10997, n10998, n10999, n11000, n11001, n11002, n11003,
         n11004, n11005, n11006, n11007, n11008, n11009, n11010, n11011,
         n11012, n11013, n11014, n11015, n11016, n11017, n11018, n11019,
         n11020, n11021, n11022, n11023, n11024, n11025, n11026, n11027,
         n11028, n11029, n11030, n11031, n11032, n11033, n11034, n11035,
         n11036, n11037, n11038, n11039, n11040, n11041, n11042, n11043,
         n11044, n11045, n11046, n11047, n11048, n11049, n11050, n11051,
         n11052, n11053, n11054, n11055, n11056, n11057, n11058, n11059,
         n11060, n11061, n11062, n11063, n11064, n11065, n11066, n11067,
         n11068, n11069, n11070, n11071, n11072, n11073, n11074, n11075,
         n11076, n11077, n11078, n11079, n11080, n11081, n11082, n11083,
         n11084, n11085, n11086, n11087, n11088, n11089, n11090, n11091,
         n11092, n11093, n11094, n11095, n11096, n11097, n11098, n11099,
         n11100, n11101, n11102, n11103, n11104, n11105, n11106, n11107,
         n11108, n11109, n11110, n11111, n11112, n11113, n11114, n11115,
         n11116, n11117, n11118, n11119, n11120, n11121, n11122, n11123,
         n11124, n11125, n11126, n11127, n11128, n11129, n11130, n11131,
         n11132, n11133, n11134, n11135, n11136, n11137, n11138, n11139,
         n11140, n11141, n11142, n11143, n11144, n11145, n11146, n11147,
         n11148, n11149, n11150, n11151, n11152, n11153, n11154, n11155,
         n11156, n11157, n11158, n11159, n11160, n11161, n11162, n11163,
         n11164, n11165, n11166, n11167, n11168, n11169, n11170, n11171,
         n11172, n11173, n11174, n11175, n11176, n11177, n11178, n11179,
         n11180, n11181, n11182, n11183, n11184, n11185, n11186, n11187,
         n11188, n11189, n11190, n11191, n11192, n11193, n11194, n11195,
         n11196, n11197, n11198, n11199, n11200, n11201, n11202, n11203,
         n11204, n11205, n11206, n11207, n11208, n11209, n11210, n11211,
         n11212, n11213, n11214, n11215, n11216, n11217, n11218, n11219,
         n11220, n11221, n11222, n11223, n11224, n11225, n11226, n11227,
         n11228, n11229, n11230, n11231, n11232, n11233, n11234, n11235,
         n11236, n11237, n11238, n11239, n11240, n11241, n11242, n11243,
         n11244, n11245, n11246, n11247, n11248, n11249, n11250, n11251,
         n11252, n11253, n11254, n11255, n11256, n11257, n11258, n11259,
         n11260, n11261, n11262, n11263, n11264, n11265, n11266, n11267,
         n11268, n11269, n11270, n11271, n11272, n11273, n11274, n11275,
         n11276, n11277, n11278, n11279, n11280, n11281, n11282, n11283,
         n11284, n11285, n11286, n11287, n11288, n11289, n11290, n11291,
         n11292, n11293, n11294, n11295, n11296, n11297, n11298, n11299,
         n11300, n11301, n11302, n11303, n11304, n11305, n11306, n11307,
         n11308, n11309, n11310, n11311, n11312, n11313, n11314, n11315,
         n11316, n11317, n11318, n11319, n11320, n11321, n11322, n11323,
         n11324, n11325, n11326, n11327, n11328, n11329, n11330, n11331,
         n11332, n11333, n11334, n11335, n11336, n11337, n11338, n11339,
         n11340, n11341, n11342, n11343, n11344, n11345, n11346, n11347,
         n11348, n11349, n11350, n11351, n11352, n11353, n11354, n11355,
         n11356, n11357, n11358, n11359, n11360, n11361, n11362, n11363,
         n11364, n11365, n11366, n11367, n11368, n11369, n11370, n11371,
         n11372, n11373, n11374, n11375, n11376, n11377, n11378, n11379,
         n11380, n11381, n11382, n11383, n11384, n11385, n11386, n11387,
         n11388, n11389, n11390, n11391, n11392, n11393, n11394, n11395,
         n11396, n11397, n11398, n11399, n11400, n11401, n11402, n11403,
         n11404, n11405, n11406, n11407, n11408, n11409, n11410, n11411,
         n11412, n11413, n11414, n11415, n11416, n11417, n11418, n11419,
         n11420, n11421, n11422, n11423, n11424, n11425, n11426, n11427,
         n11428, n11429, n11430, n11431, n11432, n11433, n11434, n11435,
         n11436, n11437, n11438, n11439, n11440, n11441, n11442, n11443,
         n11444, n11445, n11446, n11447, n11448, n11449, n11450, n11451,
         n11452, n11453, n11454, n11455, n11456, n11457, n11458, n11459,
         n11460, n11461, n11462, n11463, n11464, n11465, n11466, n11467,
         n11468, n11469, n11470, n11471, n11472, n11473, n11474, n11475,
         n11476, n11477, n11478, n11479, n11480, n11481, n11482, n11483,
         n11484, n11485, n11486, n11487, n11488, n11489, n11490, n11491,
         n11492, n11493, n11494, n11495, n11496, n11497, n11498, n11499,
         n11500, n11501, n11502, n11503, n11504, n11505, n11506, n11507,
         n11508, n11509, n11510, n11511, n11512, n11513, n11514, n11515,
         n11516, n11517, n11518, n11519, n11520, n11521, n11522, n11523,
         n11524, n11525, n11526, n11527, n11528, n11529, n11530, n11531,
         n11532, n11533, n11534, n11535, n11536, n11537, n11538, n11539,
         n11540, n11541, n11542, n11543, n11544, n11545, n11546, n11547,
         n11548, n11549, n11550, n11551, n11552, n11553, n11554, n11555,
         n11556, n11557, n11558, n11559, n11560, n11561, n11562, n11563,
         n11564, n11565, n11566, n11567, n11568, n11569, n11570, n11571,
         n11572, n11573, n11574, n11575, n11576, n11577, n11578, n11579,
         n11580, n11581, n11582, n11583, n11584, n11585, n11586, n11587,
         n11588, n11589, n11590, n11591, n11592, n11593, n11594, n11595,
         n11596, n11597, n11598, n11599, n11600, n11601, n11602, n11603,
         n11604;
  assign \knn_comb_/min_val_out[0][0]  = p_input[480];
  assign \knn_comb_/min_val_out[0][1]  = p_input[481];
  assign \knn_comb_/min_val_out[0][2]  = p_input[482];
  assign \knn_comb_/min_val_out[0][3]  = p_input[483];
  assign \knn_comb_/min_val_out[0][4]  = p_input[484];
  assign \knn_comb_/min_val_out[0][5]  = p_input[485];
  assign \knn_comb_/min_val_out[0][6]  = p_input[486];
  assign \knn_comb_/min_val_out[0][7]  = p_input[487];
  assign \knn_comb_/min_val_out[0][8]  = p_input[488];
  assign \knn_comb_/min_val_out[0][9]  = p_input[489];
  assign \knn_comb_/min_val_out[0][10]  = p_input[490];
  assign \knn_comb_/min_val_out[0][11]  = p_input[491];
  assign \knn_comb_/min_val_out[0][12]  = p_input[492];
  assign \knn_comb_/min_val_out[0][13]  = p_input[493];
  assign \knn_comb_/min_val_out[0][14]  = p_input[494];
  assign \knn_comb_/min_val_out[0][15]  = p_input[495];
  assign \knn_comb_/min_val_out[0][16]  = p_input[496];
  assign \knn_comb_/min_val_out[0][17]  = p_input[497];
  assign \knn_comb_/min_val_out[0][18]  = p_input[498];
  assign \knn_comb_/min_val_out[0][19]  = p_input[499];
  assign \knn_comb_/min_val_out[0][20]  = p_input[500];
  assign \knn_comb_/min_val_out[0][21]  = p_input[501];
  assign \knn_comb_/min_val_out[0][22]  = p_input[502];
  assign \knn_comb_/min_val_out[0][23]  = p_input[503];
  assign \knn_comb_/min_val_out[0][24]  = p_input[504];
  assign \knn_comb_/min_val_out[0][25]  = p_input[505];
  assign \knn_comb_/min_val_out[0][26]  = p_input[506];
  assign \knn_comb_/min_val_out[0][27]  = p_input[507];
  assign \knn_comb_/min_val_out[0][28]  = p_input[508];
  assign \knn_comb_/min_val_out[0][29]  = p_input[509];
  assign \knn_comb_/min_val_out[0][30]  = p_input[510];
  assign \knn_comb_/min_val_out[0][31]  = p_input[511];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][0]  = p_input[416];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][1]  = p_input[417];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][2]  = p_input[418];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][3]  = p_input[419];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][4]  = p_input[420];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][5]  = p_input[421];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][6]  = p_input[422];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][7]  = p_input[423];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][8]  = p_input[424];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][9]  = p_input[425];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][10]  = p_input[426];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][11]  = p_input[427];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][12]  = p_input[428];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][13]  = p_input[429];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][14]  = p_input[430];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][15]  = p_input[431];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][16]  = p_input[432];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][17]  = p_input[433];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][18]  = p_input[434];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][19]  = p_input[435];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][20]  = p_input[436];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][21]  = p_input[437];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][22]  = p_input[438];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][23]  = p_input[439];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][24]  = p_input[440];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][25]  = p_input[441];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][26]  = p_input[442];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][27]  = p_input[443];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][28]  = p_input[444];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][29]  = p_input[445];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][30]  = p_input[446];
  assign \knn_comb_/ASN_1[2].knn_/local_min_val[2][31]  = p_input[447];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][0]  = p_input[448];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][1]  = p_input[449];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][2]  = p_input[450];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][3]  = p_input[451];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][4]  = p_input[452];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][5]  = p_input[453];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][6]  = p_input[454];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][7]  = p_input[455];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][8]  = p_input[456];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][9]  = p_input[457];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][10]  = p_input[458];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][11]  = p_input[459];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][12]  = p_input[460];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][13]  = p_input[461];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][14]  = p_input[462];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][15]  = p_input[463];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][16]  = p_input[464];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][17]  = p_input[465];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][18]  = p_input[466];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][19]  = p_input[467];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][20]  = p_input[468];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][21]  = p_input[469];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][22]  = p_input[470];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][23]  = p_input[471];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][24]  = p_input[472];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][25]  = p_input[473];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][26]  = p_input[474];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][27]  = p_input[475];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][28]  = p_input[476];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][29]  = p_input[477];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][30]  = p_input[478];
  assign \knn_comb_/ASN_1[1].knn_/local_min_val[1][31]  = p_input[479];

  XOR U1 ( .A(n1), .B(n2), .Z(o[9]) );
  XOR U2 ( .A(n3), .B(n4), .Z(o[95]) );
  XOR U3 ( .A(n5), .B(n6), .Z(o[94]) );
  XOR U4 ( .A(n7), .B(n8), .Z(o[93]) );
  XOR U5 ( .A(n9), .B(n10), .Z(o[92]) );
  XOR U6 ( .A(n11), .B(n12), .Z(o[91]) );
  XOR U7 ( .A(n13), .B(n14), .Z(o[90]) );
  XOR U8 ( .A(n15), .B(n16), .Z(o[8]) );
  XOR U9 ( .A(n17), .B(n18), .Z(o[89]) );
  XOR U10 ( .A(n19), .B(n20), .Z(o[88]) );
  XOR U11 ( .A(n21), .B(n22), .Z(o[87]) );
  XOR U12 ( .A(n23), .B(n24), .Z(o[86]) );
  XOR U13 ( .A(n25), .B(n26), .Z(o[85]) );
  XOR U14 ( .A(n27), .B(n28), .Z(o[84]) );
  XOR U15 ( .A(n29), .B(n30), .Z(o[83]) );
  XOR U16 ( .A(n31), .B(n32), .Z(o[82]) );
  XOR U17 ( .A(n33), .B(n34), .Z(o[81]) );
  XOR U18 ( .A(n35), .B(n36), .Z(o[80]) );
  XOR U19 ( .A(n37), .B(n38), .Z(o[7]) );
  XOR U20 ( .A(n39), .B(n40), .Z(o[79]) );
  XOR U21 ( .A(n41), .B(n42), .Z(o[78]) );
  XOR U22 ( .A(n43), .B(n44), .Z(o[77]) );
  XOR U23 ( .A(n45), .B(n46), .Z(o[76]) );
  XOR U24 ( .A(n47), .B(n48), .Z(o[75]) );
  XOR U25 ( .A(n49), .B(n50), .Z(o[74]) );
  XOR U26 ( .A(n51), .B(n52), .Z(o[73]) );
  XOR U27 ( .A(n53), .B(n54), .Z(o[72]) );
  XOR U28 ( .A(n55), .B(n56), .Z(o[71]) );
  XOR U29 ( .A(n57), .B(n58), .Z(o[70]) );
  XOR U30 ( .A(n59), .B(n60), .Z(o[6]) );
  XOR U31 ( .A(n61), .B(n62), .Z(o[69]) );
  XOR U32 ( .A(n63), .B(n64), .Z(o[68]) );
  XOR U33 ( .A(n65), .B(n66), .Z(o[67]) );
  XOR U34 ( .A(n67), .B(n68), .Z(o[66]) );
  XOR U35 ( .A(n69), .B(n70), .Z(o[65]) );
  XOR U36 ( .A(n71), .B(n72), .Z(o[64]) );
  XOR U37 ( .A(n73), .B(n74), .Z(o[63]) );
  XOR U38 ( .A(n75), .B(n76), .Z(o[62]) );
  XOR U39 ( .A(n77), .B(n78), .Z(o[61]) );
  XOR U40 ( .A(n79), .B(n80), .Z(o[60]) );
  XOR U41 ( .A(n81), .B(n82), .Z(o[5]) );
  XOR U42 ( .A(n83), .B(n84), .Z(o[59]) );
  XOR U43 ( .A(n85), .B(n86), .Z(o[58]) );
  XOR U44 ( .A(n87), .B(n88), .Z(o[57]) );
  XOR U45 ( .A(n89), .B(n90), .Z(o[56]) );
  XOR U46 ( .A(n91), .B(n92), .Z(o[55]) );
  XOR U47 ( .A(n93), .B(n94), .Z(o[54]) );
  XOR U48 ( .A(n95), .B(n96), .Z(o[53]) );
  XOR U49 ( .A(n97), .B(n98), .Z(o[52]) );
  XOR U50 ( .A(n99), .B(n100), .Z(o[51]) );
  XOR U51 ( .A(n101), .B(n102), .Z(o[50]) );
  XOR U52 ( .A(n103), .B(n104), .Z(o[4]) );
  XOR U53 ( .A(n105), .B(n106), .Z(o[49]) );
  XOR U54 ( .A(n107), .B(n108), .Z(o[48]) );
  XOR U55 ( .A(n109), .B(n110), .Z(o[47]) );
  XOR U56 ( .A(n111), .B(n112), .Z(o[46]) );
  XOR U57 ( .A(n113), .B(n114), .Z(o[45]) );
  XOR U58 ( .A(n115), .B(n116), .Z(o[44]) );
  XOR U59 ( .A(n117), .B(n118), .Z(o[43]) );
  XOR U60 ( .A(n119), .B(n120), .Z(o[42]) );
  XOR U61 ( .A(n1), .B(n121), .Z(o[41]) );
  AND U62 ( .A(n122), .B(n123), .Z(n1) );
  XOR U63 ( .A(n2), .B(n121), .Z(n123) );
  XOR U64 ( .A(n124), .B(n51), .Z(n121) );
  AND U65 ( .A(n125), .B(n126), .Z(n51) );
  XNOR U66 ( .A(n127), .B(n52), .Z(n126) );
  XOR U67 ( .A(n128), .B(n129), .Z(n52) );
  AND U68 ( .A(n130), .B(n131), .Z(n129) );
  XOR U69 ( .A(p_input[9]), .B(n128), .Z(n131) );
  XOR U70 ( .A(n132), .B(n133), .Z(n128) );
  AND U71 ( .A(n134), .B(n135), .Z(n133) );
  IV U72 ( .A(n124), .Z(n127) );
  XOR U73 ( .A(n136), .B(n137), .Z(n124) );
  AND U74 ( .A(n138), .B(n139), .Z(n137) );
  XOR U75 ( .A(n140), .B(n141), .Z(n2) );
  AND U76 ( .A(n142), .B(n139), .Z(n141) );
  XNOR U77 ( .A(n143), .B(n136), .Z(n139) );
  XOR U78 ( .A(n144), .B(n145), .Z(n136) );
  AND U79 ( .A(n146), .B(n135), .Z(n145) );
  XNOR U80 ( .A(n147), .B(n132), .Z(n135) );
  XOR U81 ( .A(n148), .B(n149), .Z(n132) );
  AND U82 ( .A(n150), .B(n151), .Z(n149) );
  XOR U83 ( .A(p_input[41]), .B(n148), .Z(n151) );
  XOR U84 ( .A(n152), .B(n153), .Z(n148) );
  AND U85 ( .A(n154), .B(n155), .Z(n153) );
  IV U86 ( .A(n144), .Z(n147) );
  XOR U87 ( .A(n156), .B(n157), .Z(n144) );
  AND U88 ( .A(n158), .B(n159), .Z(n157) );
  IV U89 ( .A(n140), .Z(n143) );
  XNOR U90 ( .A(n160), .B(n161), .Z(n140) );
  AND U91 ( .A(n162), .B(n159), .Z(n161) );
  XNOR U92 ( .A(n160), .B(n156), .Z(n159) );
  XOR U93 ( .A(n163), .B(n164), .Z(n156) );
  AND U94 ( .A(n165), .B(n155), .Z(n164) );
  XNOR U95 ( .A(n166), .B(n152), .Z(n155) );
  XOR U96 ( .A(n167), .B(n168), .Z(n152) );
  AND U97 ( .A(n169), .B(n170), .Z(n168) );
  XOR U98 ( .A(p_input[73]), .B(n167), .Z(n170) );
  XOR U99 ( .A(n171), .B(n172), .Z(n167) );
  AND U100 ( .A(n173), .B(n174), .Z(n172) );
  IV U101 ( .A(n163), .Z(n166) );
  XOR U102 ( .A(n175), .B(n176), .Z(n163) );
  AND U103 ( .A(n177), .B(n178), .Z(n176) );
  XOR U104 ( .A(n179), .B(n180), .Z(n160) );
  AND U105 ( .A(n181), .B(n178), .Z(n180) );
  XNOR U106 ( .A(n179), .B(n175), .Z(n178) );
  XOR U107 ( .A(n182), .B(n183), .Z(n175) );
  AND U108 ( .A(n184), .B(n174), .Z(n183) );
  XNOR U109 ( .A(n185), .B(n171), .Z(n174) );
  XOR U110 ( .A(n186), .B(n187), .Z(n171) );
  AND U111 ( .A(n188), .B(n189), .Z(n187) );
  XOR U112 ( .A(p_input[105]), .B(n186), .Z(n189) );
  XOR U113 ( .A(n190), .B(n191), .Z(n186) );
  AND U114 ( .A(n192), .B(n193), .Z(n191) );
  IV U115 ( .A(n182), .Z(n185) );
  XOR U116 ( .A(n194), .B(n195), .Z(n182) );
  AND U117 ( .A(n196), .B(n197), .Z(n195) );
  XOR U118 ( .A(n198), .B(n199), .Z(n179) );
  AND U119 ( .A(n200), .B(n197), .Z(n199) );
  XNOR U120 ( .A(n198), .B(n194), .Z(n197) );
  XOR U121 ( .A(n201), .B(n202), .Z(n194) );
  AND U122 ( .A(n203), .B(n193), .Z(n202) );
  XNOR U123 ( .A(n204), .B(n190), .Z(n193) );
  XOR U124 ( .A(n205), .B(n206), .Z(n190) );
  AND U125 ( .A(n207), .B(n208), .Z(n206) );
  XOR U126 ( .A(p_input[137]), .B(n205), .Z(n208) );
  XOR U127 ( .A(n209), .B(n210), .Z(n205) );
  AND U128 ( .A(n211), .B(n212), .Z(n210) );
  IV U129 ( .A(n201), .Z(n204) );
  XOR U130 ( .A(n213), .B(n214), .Z(n201) );
  AND U131 ( .A(n215), .B(n216), .Z(n214) );
  XOR U132 ( .A(n217), .B(n218), .Z(n198) );
  AND U133 ( .A(n219), .B(n216), .Z(n218) );
  XNOR U134 ( .A(n217), .B(n213), .Z(n216) );
  XOR U135 ( .A(n220), .B(n221), .Z(n213) );
  AND U136 ( .A(n222), .B(n212), .Z(n221) );
  XNOR U137 ( .A(n223), .B(n209), .Z(n212) );
  XOR U138 ( .A(n224), .B(n225), .Z(n209) );
  AND U139 ( .A(n226), .B(n227), .Z(n225) );
  XOR U140 ( .A(p_input[169]), .B(n224), .Z(n227) );
  XOR U141 ( .A(n228), .B(n229), .Z(n224) );
  AND U142 ( .A(n230), .B(n231), .Z(n229) );
  IV U143 ( .A(n220), .Z(n223) );
  XOR U144 ( .A(n232), .B(n233), .Z(n220) );
  AND U145 ( .A(n234), .B(n235), .Z(n233) );
  XOR U146 ( .A(n236), .B(n237), .Z(n217) );
  AND U147 ( .A(n238), .B(n235), .Z(n237) );
  XNOR U148 ( .A(n236), .B(n232), .Z(n235) );
  XOR U149 ( .A(n239), .B(n240), .Z(n232) );
  AND U150 ( .A(n241), .B(n231), .Z(n240) );
  XNOR U151 ( .A(n242), .B(n228), .Z(n231) );
  XOR U152 ( .A(n243), .B(n244), .Z(n228) );
  AND U153 ( .A(n245), .B(n246), .Z(n244) );
  XOR U154 ( .A(p_input[201]), .B(n243), .Z(n246) );
  XOR U155 ( .A(n247), .B(n248), .Z(n243) );
  AND U156 ( .A(n249), .B(n250), .Z(n248) );
  IV U157 ( .A(n239), .Z(n242) );
  XOR U158 ( .A(n251), .B(n252), .Z(n239) );
  AND U159 ( .A(n253), .B(n254), .Z(n252) );
  XOR U160 ( .A(n255), .B(n256), .Z(n236) );
  AND U161 ( .A(n257), .B(n254), .Z(n256) );
  XNOR U162 ( .A(n255), .B(n251), .Z(n254) );
  XOR U163 ( .A(n258), .B(n259), .Z(n251) );
  AND U164 ( .A(n260), .B(n250), .Z(n259) );
  XNOR U165 ( .A(n261), .B(n247), .Z(n250) );
  XOR U166 ( .A(n262), .B(n263), .Z(n247) );
  AND U167 ( .A(n264), .B(n265), .Z(n263) );
  XOR U168 ( .A(p_input[233]), .B(n262), .Z(n265) );
  XOR U169 ( .A(n266), .B(n267), .Z(n262) );
  AND U170 ( .A(n268), .B(n269), .Z(n267) );
  IV U171 ( .A(n258), .Z(n261) );
  XOR U172 ( .A(n270), .B(n271), .Z(n258) );
  AND U173 ( .A(n272), .B(n273), .Z(n271) );
  XOR U174 ( .A(n274), .B(n275), .Z(n255) );
  AND U175 ( .A(n276), .B(n273), .Z(n275) );
  XNOR U176 ( .A(n274), .B(n270), .Z(n273) );
  XOR U177 ( .A(n277), .B(n278), .Z(n270) );
  AND U178 ( .A(n279), .B(n269), .Z(n278) );
  XNOR U179 ( .A(n280), .B(n266), .Z(n269) );
  XOR U180 ( .A(n281), .B(n282), .Z(n266) );
  AND U181 ( .A(n283), .B(n284), .Z(n282) );
  XOR U182 ( .A(p_input[265]), .B(n281), .Z(n284) );
  XOR U183 ( .A(n285), .B(n286), .Z(n281) );
  AND U184 ( .A(n287), .B(n288), .Z(n286) );
  IV U185 ( .A(n277), .Z(n280) );
  XOR U186 ( .A(n289), .B(n290), .Z(n277) );
  AND U187 ( .A(n291), .B(n292), .Z(n290) );
  XOR U188 ( .A(n293), .B(n294), .Z(n274) );
  AND U189 ( .A(n295), .B(n292), .Z(n294) );
  XNOR U190 ( .A(n293), .B(n289), .Z(n292) );
  XOR U191 ( .A(n296), .B(n297), .Z(n289) );
  AND U192 ( .A(n298), .B(n288), .Z(n297) );
  XNOR U193 ( .A(n299), .B(n285), .Z(n288) );
  XOR U194 ( .A(n300), .B(n301), .Z(n285) );
  AND U195 ( .A(n302), .B(n303), .Z(n301) );
  XOR U196 ( .A(p_input[297]), .B(n300), .Z(n303) );
  XOR U197 ( .A(n304), .B(n305), .Z(n300) );
  AND U198 ( .A(n306), .B(n307), .Z(n305) );
  IV U199 ( .A(n296), .Z(n299) );
  XOR U200 ( .A(n308), .B(n309), .Z(n296) );
  AND U201 ( .A(n310), .B(n311), .Z(n309) );
  XOR U202 ( .A(n312), .B(n313), .Z(n293) );
  AND U203 ( .A(n314), .B(n311), .Z(n313) );
  XNOR U204 ( .A(n312), .B(n308), .Z(n311) );
  XOR U205 ( .A(n315), .B(n316), .Z(n308) );
  AND U206 ( .A(n317), .B(n307), .Z(n316) );
  XNOR U207 ( .A(n318), .B(n304), .Z(n307) );
  XOR U208 ( .A(n319), .B(n320), .Z(n304) );
  AND U209 ( .A(n321), .B(n322), .Z(n320) );
  XOR U210 ( .A(p_input[329]), .B(n319), .Z(n322) );
  XOR U211 ( .A(n323), .B(n324), .Z(n319) );
  AND U212 ( .A(n325), .B(n326), .Z(n324) );
  IV U213 ( .A(n315), .Z(n318) );
  XOR U214 ( .A(n327), .B(n328), .Z(n315) );
  AND U215 ( .A(n329), .B(n330), .Z(n328) );
  XOR U216 ( .A(n331), .B(n332), .Z(n312) );
  AND U217 ( .A(n333), .B(n330), .Z(n332) );
  XNOR U218 ( .A(n331), .B(n327), .Z(n330) );
  XOR U219 ( .A(n334), .B(n335), .Z(n327) );
  AND U220 ( .A(n336), .B(n326), .Z(n335) );
  XNOR U221 ( .A(n337), .B(n323), .Z(n326) );
  XOR U222 ( .A(n338), .B(n339), .Z(n323) );
  AND U223 ( .A(n340), .B(n341), .Z(n339) );
  XOR U224 ( .A(p_input[361]), .B(n338), .Z(n341) );
  XOR U225 ( .A(n342), .B(n343), .Z(n338) );
  AND U226 ( .A(n344), .B(n345), .Z(n343) );
  IV U227 ( .A(n334), .Z(n337) );
  XOR U228 ( .A(n346), .B(n347), .Z(n334) );
  AND U229 ( .A(n348), .B(n349), .Z(n347) );
  XOR U230 ( .A(n350), .B(n351), .Z(n331) );
  AND U231 ( .A(n352), .B(n349), .Z(n351) );
  XNOR U232 ( .A(n350), .B(n346), .Z(n349) );
  XOR U233 ( .A(n353), .B(n354), .Z(n346) );
  AND U234 ( .A(n355), .B(n345), .Z(n354) );
  XNOR U235 ( .A(n356), .B(n342), .Z(n345) );
  XOR U236 ( .A(n357), .B(n358), .Z(n342) );
  AND U237 ( .A(n359), .B(n360), .Z(n358) );
  XOR U238 ( .A(p_input[393]), .B(n357), .Z(n360) );
  XOR U239 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(n361), .Z(
        n357) );
  AND U240 ( .A(n362), .B(n363), .Z(n361) );
  IV U241 ( .A(n353), .Z(n356) );
  XOR U242 ( .A(n364), .B(n365), .Z(n353) );
  AND U243 ( .A(n366), .B(n367), .Z(n365) );
  XOR U244 ( .A(n368), .B(n369), .Z(n350) );
  AND U245 ( .A(n370), .B(n367), .Z(n369) );
  XNOR U246 ( .A(n368), .B(n364), .Z(n367) );
  XNOR U247 ( .A(n371), .B(n372), .Z(n364) );
  AND U248 ( .A(n373), .B(n363), .Z(n372) );
  XNOR U249 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(n371), .Z(
        n363) );
  XNOR U250 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .B(n374), .Z(
        n371) );
  AND U251 ( .A(n375), .B(n376), .Z(n374) );
  XNOR U252 ( .A(\knn_comb_/min_val_out[0][9] ), .B(n377), .Z(n368) );
  AND U253 ( .A(n378), .B(n376), .Z(n377) );
  XOR U254 ( .A(n379), .B(n380), .Z(n376) );
  XOR U255 ( .A(n15), .B(n381), .Z(o[40]) );
  AND U256 ( .A(n122), .B(n382), .Z(n15) );
  XOR U257 ( .A(n16), .B(n381), .Z(n382) );
  XOR U258 ( .A(n383), .B(n53), .Z(n381) );
  AND U259 ( .A(n125), .B(n384), .Z(n53) );
  XNOR U260 ( .A(n385), .B(n54), .Z(n384) );
  XOR U261 ( .A(n386), .B(n387), .Z(n54) );
  AND U262 ( .A(n130), .B(n388), .Z(n387) );
  XOR U263 ( .A(p_input[8]), .B(n386), .Z(n388) );
  XOR U264 ( .A(n389), .B(n390), .Z(n386) );
  AND U265 ( .A(n134), .B(n391), .Z(n390) );
  IV U266 ( .A(n383), .Z(n385) );
  XOR U267 ( .A(n392), .B(n393), .Z(n383) );
  AND U268 ( .A(n138), .B(n394), .Z(n393) );
  XOR U269 ( .A(n395), .B(n396), .Z(n16) );
  AND U270 ( .A(n142), .B(n394), .Z(n396) );
  XNOR U271 ( .A(n397), .B(n392), .Z(n394) );
  XOR U272 ( .A(n398), .B(n399), .Z(n392) );
  AND U273 ( .A(n146), .B(n391), .Z(n399) );
  XNOR U274 ( .A(n400), .B(n389), .Z(n391) );
  XOR U275 ( .A(n401), .B(n402), .Z(n389) );
  AND U276 ( .A(n150), .B(n403), .Z(n402) );
  XOR U277 ( .A(p_input[40]), .B(n401), .Z(n403) );
  XOR U278 ( .A(n404), .B(n405), .Z(n401) );
  AND U279 ( .A(n154), .B(n406), .Z(n405) );
  IV U280 ( .A(n398), .Z(n400) );
  XOR U281 ( .A(n407), .B(n408), .Z(n398) );
  AND U282 ( .A(n158), .B(n409), .Z(n408) );
  IV U283 ( .A(n395), .Z(n397) );
  XNOR U284 ( .A(n410), .B(n411), .Z(n395) );
  AND U285 ( .A(n162), .B(n409), .Z(n411) );
  XNOR U286 ( .A(n410), .B(n407), .Z(n409) );
  XOR U287 ( .A(n412), .B(n413), .Z(n407) );
  AND U288 ( .A(n165), .B(n406), .Z(n413) );
  XNOR U289 ( .A(n414), .B(n404), .Z(n406) );
  XOR U290 ( .A(n415), .B(n416), .Z(n404) );
  AND U291 ( .A(n169), .B(n417), .Z(n416) );
  XOR U292 ( .A(p_input[72]), .B(n415), .Z(n417) );
  XOR U293 ( .A(n418), .B(n419), .Z(n415) );
  AND U294 ( .A(n173), .B(n420), .Z(n419) );
  IV U295 ( .A(n412), .Z(n414) );
  XOR U296 ( .A(n421), .B(n422), .Z(n412) );
  AND U297 ( .A(n177), .B(n423), .Z(n422) );
  XOR U298 ( .A(n424), .B(n425), .Z(n410) );
  AND U299 ( .A(n181), .B(n423), .Z(n425) );
  XNOR U300 ( .A(n424), .B(n421), .Z(n423) );
  XOR U301 ( .A(n426), .B(n427), .Z(n421) );
  AND U302 ( .A(n184), .B(n420), .Z(n427) );
  XNOR U303 ( .A(n428), .B(n418), .Z(n420) );
  XOR U304 ( .A(n429), .B(n430), .Z(n418) );
  AND U305 ( .A(n188), .B(n431), .Z(n430) );
  XOR U306 ( .A(p_input[104]), .B(n429), .Z(n431) );
  XOR U307 ( .A(n432), .B(n433), .Z(n429) );
  AND U308 ( .A(n192), .B(n434), .Z(n433) );
  IV U309 ( .A(n426), .Z(n428) );
  XOR U310 ( .A(n435), .B(n436), .Z(n426) );
  AND U311 ( .A(n196), .B(n437), .Z(n436) );
  XOR U312 ( .A(n438), .B(n439), .Z(n424) );
  AND U313 ( .A(n200), .B(n437), .Z(n439) );
  XNOR U314 ( .A(n438), .B(n435), .Z(n437) );
  XOR U315 ( .A(n440), .B(n441), .Z(n435) );
  AND U316 ( .A(n203), .B(n434), .Z(n441) );
  XNOR U317 ( .A(n442), .B(n432), .Z(n434) );
  XOR U318 ( .A(n443), .B(n444), .Z(n432) );
  AND U319 ( .A(n207), .B(n445), .Z(n444) );
  XOR U320 ( .A(p_input[136]), .B(n443), .Z(n445) );
  XOR U321 ( .A(n446), .B(n447), .Z(n443) );
  AND U322 ( .A(n211), .B(n448), .Z(n447) );
  IV U323 ( .A(n440), .Z(n442) );
  XOR U324 ( .A(n449), .B(n450), .Z(n440) );
  AND U325 ( .A(n215), .B(n451), .Z(n450) );
  XOR U326 ( .A(n452), .B(n453), .Z(n438) );
  AND U327 ( .A(n219), .B(n451), .Z(n453) );
  XNOR U328 ( .A(n452), .B(n449), .Z(n451) );
  XOR U329 ( .A(n454), .B(n455), .Z(n449) );
  AND U330 ( .A(n222), .B(n448), .Z(n455) );
  XNOR U331 ( .A(n456), .B(n446), .Z(n448) );
  XOR U332 ( .A(n457), .B(n458), .Z(n446) );
  AND U333 ( .A(n226), .B(n459), .Z(n458) );
  XOR U334 ( .A(p_input[168]), .B(n457), .Z(n459) );
  XOR U335 ( .A(n460), .B(n461), .Z(n457) );
  AND U336 ( .A(n230), .B(n462), .Z(n461) );
  IV U337 ( .A(n454), .Z(n456) );
  XOR U338 ( .A(n463), .B(n464), .Z(n454) );
  AND U339 ( .A(n234), .B(n465), .Z(n464) );
  XOR U340 ( .A(n466), .B(n467), .Z(n452) );
  AND U341 ( .A(n238), .B(n465), .Z(n467) );
  XNOR U342 ( .A(n466), .B(n463), .Z(n465) );
  XOR U343 ( .A(n468), .B(n469), .Z(n463) );
  AND U344 ( .A(n241), .B(n462), .Z(n469) );
  XNOR U345 ( .A(n470), .B(n460), .Z(n462) );
  XOR U346 ( .A(n471), .B(n472), .Z(n460) );
  AND U347 ( .A(n245), .B(n473), .Z(n472) );
  XOR U348 ( .A(p_input[200]), .B(n471), .Z(n473) );
  XOR U349 ( .A(n474), .B(n475), .Z(n471) );
  AND U350 ( .A(n249), .B(n476), .Z(n475) );
  IV U351 ( .A(n468), .Z(n470) );
  XOR U352 ( .A(n477), .B(n478), .Z(n468) );
  AND U353 ( .A(n253), .B(n479), .Z(n478) );
  XOR U354 ( .A(n480), .B(n481), .Z(n466) );
  AND U355 ( .A(n257), .B(n479), .Z(n481) );
  XNOR U356 ( .A(n480), .B(n477), .Z(n479) );
  XOR U357 ( .A(n482), .B(n483), .Z(n477) );
  AND U358 ( .A(n260), .B(n476), .Z(n483) );
  XNOR U359 ( .A(n484), .B(n474), .Z(n476) );
  XOR U360 ( .A(n485), .B(n486), .Z(n474) );
  AND U361 ( .A(n264), .B(n487), .Z(n486) );
  XOR U362 ( .A(p_input[232]), .B(n485), .Z(n487) );
  XOR U363 ( .A(n488), .B(n489), .Z(n485) );
  AND U364 ( .A(n268), .B(n490), .Z(n489) );
  IV U365 ( .A(n482), .Z(n484) );
  XOR U366 ( .A(n491), .B(n492), .Z(n482) );
  AND U367 ( .A(n272), .B(n493), .Z(n492) );
  XOR U368 ( .A(n494), .B(n495), .Z(n480) );
  AND U369 ( .A(n276), .B(n493), .Z(n495) );
  XNOR U370 ( .A(n494), .B(n491), .Z(n493) );
  XOR U371 ( .A(n496), .B(n497), .Z(n491) );
  AND U372 ( .A(n279), .B(n490), .Z(n497) );
  XNOR U373 ( .A(n498), .B(n488), .Z(n490) );
  XOR U374 ( .A(n499), .B(n500), .Z(n488) );
  AND U375 ( .A(n283), .B(n501), .Z(n500) );
  XOR U376 ( .A(p_input[264]), .B(n499), .Z(n501) );
  XOR U377 ( .A(n502), .B(n503), .Z(n499) );
  AND U378 ( .A(n287), .B(n504), .Z(n503) );
  IV U379 ( .A(n496), .Z(n498) );
  XOR U380 ( .A(n505), .B(n506), .Z(n496) );
  AND U381 ( .A(n291), .B(n507), .Z(n506) );
  XOR U382 ( .A(n508), .B(n509), .Z(n494) );
  AND U383 ( .A(n295), .B(n507), .Z(n509) );
  XNOR U384 ( .A(n508), .B(n505), .Z(n507) );
  XOR U385 ( .A(n510), .B(n511), .Z(n505) );
  AND U386 ( .A(n298), .B(n504), .Z(n511) );
  XNOR U387 ( .A(n512), .B(n502), .Z(n504) );
  XOR U388 ( .A(n513), .B(n514), .Z(n502) );
  AND U389 ( .A(n302), .B(n515), .Z(n514) );
  XOR U390 ( .A(p_input[296]), .B(n513), .Z(n515) );
  XOR U391 ( .A(n516), .B(n517), .Z(n513) );
  AND U392 ( .A(n306), .B(n518), .Z(n517) );
  IV U393 ( .A(n510), .Z(n512) );
  XOR U394 ( .A(n519), .B(n520), .Z(n510) );
  AND U395 ( .A(n310), .B(n521), .Z(n520) );
  XOR U396 ( .A(n522), .B(n523), .Z(n508) );
  AND U397 ( .A(n314), .B(n521), .Z(n523) );
  XNOR U398 ( .A(n522), .B(n519), .Z(n521) );
  XOR U399 ( .A(n524), .B(n525), .Z(n519) );
  AND U400 ( .A(n317), .B(n518), .Z(n525) );
  XNOR U401 ( .A(n526), .B(n516), .Z(n518) );
  XOR U402 ( .A(n527), .B(n528), .Z(n516) );
  AND U403 ( .A(n321), .B(n529), .Z(n528) );
  XOR U404 ( .A(p_input[328]), .B(n527), .Z(n529) );
  XOR U405 ( .A(n530), .B(n531), .Z(n527) );
  AND U406 ( .A(n325), .B(n532), .Z(n531) );
  IV U407 ( .A(n524), .Z(n526) );
  XOR U408 ( .A(n533), .B(n534), .Z(n524) );
  AND U409 ( .A(n329), .B(n535), .Z(n534) );
  XOR U410 ( .A(n536), .B(n537), .Z(n522) );
  AND U411 ( .A(n333), .B(n535), .Z(n537) );
  XNOR U412 ( .A(n536), .B(n533), .Z(n535) );
  XOR U413 ( .A(n538), .B(n539), .Z(n533) );
  AND U414 ( .A(n336), .B(n532), .Z(n539) );
  XNOR U415 ( .A(n540), .B(n530), .Z(n532) );
  XOR U416 ( .A(n541), .B(n542), .Z(n530) );
  AND U417 ( .A(n340), .B(n543), .Z(n542) );
  XOR U418 ( .A(p_input[360]), .B(n541), .Z(n543) );
  XOR U419 ( .A(n544), .B(n545), .Z(n541) );
  AND U420 ( .A(n344), .B(n546), .Z(n545) );
  IV U421 ( .A(n538), .Z(n540) );
  XOR U422 ( .A(n547), .B(n548), .Z(n538) );
  AND U423 ( .A(n348), .B(n549), .Z(n548) );
  XOR U424 ( .A(n550), .B(n551), .Z(n536) );
  AND U425 ( .A(n352), .B(n549), .Z(n551) );
  XNOR U426 ( .A(n550), .B(n547), .Z(n549) );
  XOR U427 ( .A(n552), .B(n553), .Z(n547) );
  AND U428 ( .A(n355), .B(n546), .Z(n553) );
  XNOR U429 ( .A(n554), .B(n544), .Z(n546) );
  XOR U430 ( .A(n555), .B(n556), .Z(n544) );
  AND U431 ( .A(n359), .B(n557), .Z(n556) );
  XOR U432 ( .A(p_input[392]), .B(n555), .Z(n557) );
  XOR U433 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n558), .Z(
        n555) );
  AND U434 ( .A(n362), .B(n559), .Z(n558) );
  IV U435 ( .A(n552), .Z(n554) );
  XOR U436 ( .A(n560), .B(n561), .Z(n552) );
  AND U437 ( .A(n366), .B(n562), .Z(n561) );
  XOR U438 ( .A(n563), .B(n564), .Z(n550) );
  AND U439 ( .A(n370), .B(n562), .Z(n564) );
  XNOR U440 ( .A(n563), .B(n560), .Z(n562) );
  XNOR U441 ( .A(n565), .B(n566), .Z(n560) );
  AND U442 ( .A(n373), .B(n559), .Z(n566) );
  XNOR U443 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n565), .Z(
        n559) );
  XNOR U444 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .B(n567), .Z(
        n565) );
  AND U445 ( .A(n375), .B(n568), .Z(n567) );
  XNOR U446 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n569), .Z(n563) );
  AND U447 ( .A(n378), .B(n568), .Z(n569) );
  XOR U448 ( .A(n570), .B(n571), .Z(n568) );
  IV U449 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .Z(n571) );
  IV U450 ( .A(\knn_comb_/min_val_out[0][8] ), .Z(n570) );
  XOR U451 ( .A(n572), .B(n573), .Z(o[3]) );
  XOR U452 ( .A(n37), .B(n574), .Z(o[39]) );
  AND U453 ( .A(n122), .B(n575), .Z(n37) );
  XOR U454 ( .A(n38), .B(n574), .Z(n575) );
  XOR U455 ( .A(n576), .B(n55), .Z(n574) );
  AND U456 ( .A(n125), .B(n577), .Z(n55) );
  XNOR U457 ( .A(n578), .B(n56), .Z(n577) );
  XOR U458 ( .A(n579), .B(n580), .Z(n56) );
  AND U459 ( .A(n130), .B(n581), .Z(n580) );
  XOR U460 ( .A(p_input[7]), .B(n579), .Z(n581) );
  XOR U461 ( .A(n582), .B(n583), .Z(n579) );
  AND U462 ( .A(n134), .B(n584), .Z(n583) );
  IV U463 ( .A(n576), .Z(n578) );
  XOR U464 ( .A(n585), .B(n586), .Z(n576) );
  AND U465 ( .A(n138), .B(n587), .Z(n586) );
  XOR U466 ( .A(n588), .B(n589), .Z(n38) );
  AND U467 ( .A(n142), .B(n587), .Z(n589) );
  XNOR U468 ( .A(n590), .B(n585), .Z(n587) );
  XOR U469 ( .A(n591), .B(n592), .Z(n585) );
  AND U470 ( .A(n146), .B(n584), .Z(n592) );
  XNOR U471 ( .A(n593), .B(n582), .Z(n584) );
  XOR U472 ( .A(n594), .B(n595), .Z(n582) );
  AND U473 ( .A(n150), .B(n596), .Z(n595) );
  XOR U474 ( .A(p_input[39]), .B(n594), .Z(n596) );
  XOR U475 ( .A(n597), .B(n598), .Z(n594) );
  AND U476 ( .A(n154), .B(n599), .Z(n598) );
  IV U477 ( .A(n591), .Z(n593) );
  XOR U478 ( .A(n600), .B(n601), .Z(n591) );
  AND U479 ( .A(n158), .B(n602), .Z(n601) );
  IV U480 ( .A(n588), .Z(n590) );
  XNOR U481 ( .A(n603), .B(n604), .Z(n588) );
  AND U482 ( .A(n162), .B(n602), .Z(n604) );
  XNOR U483 ( .A(n603), .B(n600), .Z(n602) );
  XOR U484 ( .A(n605), .B(n606), .Z(n600) );
  AND U485 ( .A(n165), .B(n599), .Z(n606) );
  XNOR U486 ( .A(n607), .B(n597), .Z(n599) );
  XOR U487 ( .A(n608), .B(n609), .Z(n597) );
  AND U488 ( .A(n169), .B(n610), .Z(n609) );
  XOR U489 ( .A(p_input[71]), .B(n608), .Z(n610) );
  XOR U490 ( .A(n611), .B(n612), .Z(n608) );
  AND U491 ( .A(n173), .B(n613), .Z(n612) );
  IV U492 ( .A(n605), .Z(n607) );
  XOR U493 ( .A(n614), .B(n615), .Z(n605) );
  AND U494 ( .A(n177), .B(n616), .Z(n615) );
  XOR U495 ( .A(n617), .B(n618), .Z(n603) );
  AND U496 ( .A(n181), .B(n616), .Z(n618) );
  XNOR U497 ( .A(n617), .B(n614), .Z(n616) );
  XOR U498 ( .A(n619), .B(n620), .Z(n614) );
  AND U499 ( .A(n184), .B(n613), .Z(n620) );
  XNOR U500 ( .A(n621), .B(n611), .Z(n613) );
  XOR U501 ( .A(n622), .B(n623), .Z(n611) );
  AND U502 ( .A(n188), .B(n624), .Z(n623) );
  XOR U503 ( .A(p_input[103]), .B(n622), .Z(n624) );
  XOR U504 ( .A(n625), .B(n626), .Z(n622) );
  AND U505 ( .A(n192), .B(n627), .Z(n626) );
  IV U506 ( .A(n619), .Z(n621) );
  XOR U507 ( .A(n628), .B(n629), .Z(n619) );
  AND U508 ( .A(n196), .B(n630), .Z(n629) );
  XOR U509 ( .A(n631), .B(n632), .Z(n617) );
  AND U510 ( .A(n200), .B(n630), .Z(n632) );
  XNOR U511 ( .A(n631), .B(n628), .Z(n630) );
  XOR U512 ( .A(n633), .B(n634), .Z(n628) );
  AND U513 ( .A(n203), .B(n627), .Z(n634) );
  XNOR U514 ( .A(n635), .B(n625), .Z(n627) );
  XOR U515 ( .A(n636), .B(n637), .Z(n625) );
  AND U516 ( .A(n207), .B(n638), .Z(n637) );
  XOR U517 ( .A(p_input[135]), .B(n636), .Z(n638) );
  XOR U518 ( .A(n639), .B(n640), .Z(n636) );
  AND U519 ( .A(n211), .B(n641), .Z(n640) );
  IV U520 ( .A(n633), .Z(n635) );
  XOR U521 ( .A(n642), .B(n643), .Z(n633) );
  AND U522 ( .A(n215), .B(n644), .Z(n643) );
  XOR U523 ( .A(n645), .B(n646), .Z(n631) );
  AND U524 ( .A(n219), .B(n644), .Z(n646) );
  XNOR U525 ( .A(n645), .B(n642), .Z(n644) );
  XOR U526 ( .A(n647), .B(n648), .Z(n642) );
  AND U527 ( .A(n222), .B(n641), .Z(n648) );
  XNOR U528 ( .A(n649), .B(n639), .Z(n641) );
  XOR U529 ( .A(n650), .B(n651), .Z(n639) );
  AND U530 ( .A(n226), .B(n652), .Z(n651) );
  XOR U531 ( .A(p_input[167]), .B(n650), .Z(n652) );
  XOR U532 ( .A(n653), .B(n654), .Z(n650) );
  AND U533 ( .A(n230), .B(n655), .Z(n654) );
  IV U534 ( .A(n647), .Z(n649) );
  XOR U535 ( .A(n656), .B(n657), .Z(n647) );
  AND U536 ( .A(n234), .B(n658), .Z(n657) );
  XOR U537 ( .A(n659), .B(n660), .Z(n645) );
  AND U538 ( .A(n238), .B(n658), .Z(n660) );
  XNOR U539 ( .A(n659), .B(n656), .Z(n658) );
  XOR U540 ( .A(n661), .B(n662), .Z(n656) );
  AND U541 ( .A(n241), .B(n655), .Z(n662) );
  XNOR U542 ( .A(n663), .B(n653), .Z(n655) );
  XOR U543 ( .A(n664), .B(n665), .Z(n653) );
  AND U544 ( .A(n245), .B(n666), .Z(n665) );
  XOR U545 ( .A(p_input[199]), .B(n664), .Z(n666) );
  XOR U546 ( .A(n667), .B(n668), .Z(n664) );
  AND U547 ( .A(n249), .B(n669), .Z(n668) );
  IV U548 ( .A(n661), .Z(n663) );
  XOR U549 ( .A(n670), .B(n671), .Z(n661) );
  AND U550 ( .A(n253), .B(n672), .Z(n671) );
  XOR U551 ( .A(n673), .B(n674), .Z(n659) );
  AND U552 ( .A(n257), .B(n672), .Z(n674) );
  XNOR U553 ( .A(n673), .B(n670), .Z(n672) );
  XOR U554 ( .A(n675), .B(n676), .Z(n670) );
  AND U555 ( .A(n260), .B(n669), .Z(n676) );
  XNOR U556 ( .A(n677), .B(n667), .Z(n669) );
  XOR U557 ( .A(n678), .B(n679), .Z(n667) );
  AND U558 ( .A(n264), .B(n680), .Z(n679) );
  XOR U559 ( .A(p_input[231]), .B(n678), .Z(n680) );
  XOR U560 ( .A(n681), .B(n682), .Z(n678) );
  AND U561 ( .A(n268), .B(n683), .Z(n682) );
  IV U562 ( .A(n675), .Z(n677) );
  XOR U563 ( .A(n684), .B(n685), .Z(n675) );
  AND U564 ( .A(n272), .B(n686), .Z(n685) );
  XOR U565 ( .A(n687), .B(n688), .Z(n673) );
  AND U566 ( .A(n276), .B(n686), .Z(n688) );
  XNOR U567 ( .A(n687), .B(n684), .Z(n686) );
  XOR U568 ( .A(n689), .B(n690), .Z(n684) );
  AND U569 ( .A(n279), .B(n683), .Z(n690) );
  XNOR U570 ( .A(n691), .B(n681), .Z(n683) );
  XOR U571 ( .A(n692), .B(n693), .Z(n681) );
  AND U572 ( .A(n283), .B(n694), .Z(n693) );
  XOR U573 ( .A(p_input[263]), .B(n692), .Z(n694) );
  XOR U574 ( .A(n695), .B(n696), .Z(n692) );
  AND U575 ( .A(n287), .B(n697), .Z(n696) );
  IV U576 ( .A(n689), .Z(n691) );
  XOR U577 ( .A(n698), .B(n699), .Z(n689) );
  AND U578 ( .A(n291), .B(n700), .Z(n699) );
  XOR U579 ( .A(n701), .B(n702), .Z(n687) );
  AND U580 ( .A(n295), .B(n700), .Z(n702) );
  XNOR U581 ( .A(n701), .B(n698), .Z(n700) );
  XOR U582 ( .A(n703), .B(n704), .Z(n698) );
  AND U583 ( .A(n298), .B(n697), .Z(n704) );
  XNOR U584 ( .A(n705), .B(n695), .Z(n697) );
  XOR U585 ( .A(n706), .B(n707), .Z(n695) );
  AND U586 ( .A(n302), .B(n708), .Z(n707) );
  XOR U587 ( .A(p_input[295]), .B(n706), .Z(n708) );
  XOR U588 ( .A(n709), .B(n710), .Z(n706) );
  AND U589 ( .A(n306), .B(n711), .Z(n710) );
  IV U590 ( .A(n703), .Z(n705) );
  XOR U591 ( .A(n712), .B(n713), .Z(n703) );
  AND U592 ( .A(n310), .B(n714), .Z(n713) );
  XOR U593 ( .A(n715), .B(n716), .Z(n701) );
  AND U594 ( .A(n314), .B(n714), .Z(n716) );
  XNOR U595 ( .A(n715), .B(n712), .Z(n714) );
  XOR U596 ( .A(n717), .B(n718), .Z(n712) );
  AND U597 ( .A(n317), .B(n711), .Z(n718) );
  XNOR U598 ( .A(n719), .B(n709), .Z(n711) );
  XOR U599 ( .A(n720), .B(n721), .Z(n709) );
  AND U600 ( .A(n321), .B(n722), .Z(n721) );
  XOR U601 ( .A(p_input[327]), .B(n720), .Z(n722) );
  XOR U602 ( .A(n723), .B(n724), .Z(n720) );
  AND U603 ( .A(n325), .B(n725), .Z(n724) );
  IV U604 ( .A(n717), .Z(n719) );
  XOR U605 ( .A(n726), .B(n727), .Z(n717) );
  AND U606 ( .A(n329), .B(n728), .Z(n727) );
  XOR U607 ( .A(n729), .B(n730), .Z(n715) );
  AND U608 ( .A(n333), .B(n728), .Z(n730) );
  XNOR U609 ( .A(n729), .B(n726), .Z(n728) );
  XOR U610 ( .A(n731), .B(n732), .Z(n726) );
  AND U611 ( .A(n336), .B(n725), .Z(n732) );
  XNOR U612 ( .A(n733), .B(n723), .Z(n725) );
  XOR U613 ( .A(n734), .B(n735), .Z(n723) );
  AND U614 ( .A(n340), .B(n736), .Z(n735) );
  XOR U615 ( .A(p_input[359]), .B(n734), .Z(n736) );
  XOR U616 ( .A(n737), .B(n738), .Z(n734) );
  AND U617 ( .A(n344), .B(n739), .Z(n738) );
  IV U618 ( .A(n731), .Z(n733) );
  XOR U619 ( .A(n740), .B(n741), .Z(n731) );
  AND U620 ( .A(n348), .B(n742), .Z(n741) );
  XOR U621 ( .A(n743), .B(n744), .Z(n729) );
  AND U622 ( .A(n352), .B(n742), .Z(n744) );
  XNOR U623 ( .A(n743), .B(n740), .Z(n742) );
  XOR U624 ( .A(n745), .B(n746), .Z(n740) );
  AND U625 ( .A(n355), .B(n739), .Z(n746) );
  XNOR U626 ( .A(n747), .B(n737), .Z(n739) );
  XOR U627 ( .A(n748), .B(n749), .Z(n737) );
  AND U628 ( .A(n359), .B(n750), .Z(n749) );
  XOR U629 ( .A(p_input[391]), .B(n748), .Z(n750) );
  XOR U630 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(n751), .Z(
        n748) );
  AND U631 ( .A(n362), .B(n752), .Z(n751) );
  IV U632 ( .A(n745), .Z(n747) );
  XOR U633 ( .A(n753), .B(n754), .Z(n745) );
  AND U634 ( .A(n366), .B(n755), .Z(n754) );
  XOR U635 ( .A(n756), .B(n757), .Z(n743) );
  AND U636 ( .A(n370), .B(n755), .Z(n757) );
  XNOR U637 ( .A(n756), .B(n753), .Z(n755) );
  XNOR U638 ( .A(n758), .B(n759), .Z(n753) );
  AND U639 ( .A(n373), .B(n752), .Z(n759) );
  XNOR U640 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(n758), .Z(
        n752) );
  XNOR U641 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .B(n760), .Z(
        n758) );
  AND U642 ( .A(n375), .B(n761), .Z(n760) );
  XNOR U643 ( .A(\knn_comb_/min_val_out[0][7] ), .B(n762), .Z(n756) );
  AND U644 ( .A(n378), .B(n761), .Z(n762) );
  XOR U645 ( .A(n763), .B(n764), .Z(n761) );
  XOR U646 ( .A(n59), .B(n765), .Z(o[38]) );
  AND U647 ( .A(n122), .B(n766), .Z(n59) );
  XOR U648 ( .A(n60), .B(n765), .Z(n766) );
  XOR U649 ( .A(n767), .B(n57), .Z(n765) );
  AND U650 ( .A(n125), .B(n768), .Z(n57) );
  XOR U651 ( .A(n58), .B(n767), .Z(n768) );
  XOR U652 ( .A(n769), .B(n770), .Z(n58) );
  AND U653 ( .A(n130), .B(n771), .Z(n770) );
  XOR U654 ( .A(p_input[6]), .B(n769), .Z(n771) );
  XNOR U655 ( .A(n772), .B(n773), .Z(n769) );
  AND U656 ( .A(n134), .B(n774), .Z(n773) );
  XOR U657 ( .A(n775), .B(n776), .Z(n767) );
  AND U658 ( .A(n138), .B(n777), .Z(n776) );
  XOR U659 ( .A(n778), .B(n779), .Z(n60) );
  AND U660 ( .A(n142), .B(n777), .Z(n779) );
  XNOR U661 ( .A(n780), .B(n778), .Z(n777) );
  IV U662 ( .A(n775), .Z(n780) );
  XOR U663 ( .A(n781), .B(n782), .Z(n775) );
  AND U664 ( .A(n146), .B(n774), .Z(n782) );
  XNOR U665 ( .A(n772), .B(n781), .Z(n774) );
  XNOR U666 ( .A(n783), .B(n784), .Z(n772) );
  AND U667 ( .A(n150), .B(n785), .Z(n784) );
  XOR U668 ( .A(p_input[38]), .B(n783), .Z(n785) );
  XNOR U669 ( .A(n786), .B(n787), .Z(n783) );
  AND U670 ( .A(n154), .B(n788), .Z(n787) );
  XOR U671 ( .A(n789), .B(n790), .Z(n781) );
  AND U672 ( .A(n158), .B(n791), .Z(n790) );
  XOR U673 ( .A(n792), .B(n793), .Z(n778) );
  AND U674 ( .A(n162), .B(n791), .Z(n793) );
  XNOR U675 ( .A(n794), .B(n792), .Z(n791) );
  IV U676 ( .A(n789), .Z(n794) );
  XOR U677 ( .A(n795), .B(n796), .Z(n789) );
  AND U678 ( .A(n165), .B(n788), .Z(n796) );
  XNOR U679 ( .A(n786), .B(n795), .Z(n788) );
  XNOR U680 ( .A(n797), .B(n798), .Z(n786) );
  AND U681 ( .A(n169), .B(n799), .Z(n798) );
  XOR U682 ( .A(p_input[70]), .B(n797), .Z(n799) );
  XNOR U683 ( .A(n800), .B(n801), .Z(n797) );
  AND U684 ( .A(n173), .B(n802), .Z(n801) );
  XOR U685 ( .A(n803), .B(n804), .Z(n795) );
  AND U686 ( .A(n177), .B(n805), .Z(n804) );
  XOR U687 ( .A(n806), .B(n807), .Z(n792) );
  AND U688 ( .A(n181), .B(n805), .Z(n807) );
  XNOR U689 ( .A(n808), .B(n806), .Z(n805) );
  IV U690 ( .A(n803), .Z(n808) );
  XOR U691 ( .A(n809), .B(n810), .Z(n803) );
  AND U692 ( .A(n184), .B(n802), .Z(n810) );
  XNOR U693 ( .A(n800), .B(n809), .Z(n802) );
  XNOR U694 ( .A(n811), .B(n812), .Z(n800) );
  AND U695 ( .A(n188), .B(n813), .Z(n812) );
  XOR U696 ( .A(p_input[102]), .B(n811), .Z(n813) );
  XNOR U697 ( .A(n814), .B(n815), .Z(n811) );
  AND U698 ( .A(n192), .B(n816), .Z(n815) );
  XOR U699 ( .A(n817), .B(n818), .Z(n809) );
  AND U700 ( .A(n196), .B(n819), .Z(n818) );
  XOR U701 ( .A(n820), .B(n821), .Z(n806) );
  AND U702 ( .A(n200), .B(n819), .Z(n821) );
  XNOR U703 ( .A(n822), .B(n820), .Z(n819) );
  IV U704 ( .A(n817), .Z(n822) );
  XOR U705 ( .A(n823), .B(n824), .Z(n817) );
  AND U706 ( .A(n203), .B(n816), .Z(n824) );
  XNOR U707 ( .A(n814), .B(n823), .Z(n816) );
  XNOR U708 ( .A(n825), .B(n826), .Z(n814) );
  AND U709 ( .A(n207), .B(n827), .Z(n826) );
  XOR U710 ( .A(p_input[134]), .B(n825), .Z(n827) );
  XNOR U711 ( .A(n828), .B(n829), .Z(n825) );
  AND U712 ( .A(n211), .B(n830), .Z(n829) );
  XOR U713 ( .A(n831), .B(n832), .Z(n823) );
  AND U714 ( .A(n215), .B(n833), .Z(n832) );
  XOR U715 ( .A(n834), .B(n835), .Z(n820) );
  AND U716 ( .A(n219), .B(n833), .Z(n835) );
  XNOR U717 ( .A(n836), .B(n834), .Z(n833) );
  IV U718 ( .A(n831), .Z(n836) );
  XOR U719 ( .A(n837), .B(n838), .Z(n831) );
  AND U720 ( .A(n222), .B(n830), .Z(n838) );
  XNOR U721 ( .A(n828), .B(n837), .Z(n830) );
  XNOR U722 ( .A(n839), .B(n840), .Z(n828) );
  AND U723 ( .A(n226), .B(n841), .Z(n840) );
  XOR U724 ( .A(p_input[166]), .B(n839), .Z(n841) );
  XNOR U725 ( .A(n842), .B(n843), .Z(n839) );
  AND U726 ( .A(n230), .B(n844), .Z(n843) );
  XOR U727 ( .A(n845), .B(n846), .Z(n837) );
  AND U728 ( .A(n234), .B(n847), .Z(n846) );
  XOR U729 ( .A(n848), .B(n849), .Z(n834) );
  AND U730 ( .A(n238), .B(n847), .Z(n849) );
  XNOR U731 ( .A(n850), .B(n848), .Z(n847) );
  IV U732 ( .A(n845), .Z(n850) );
  XOR U733 ( .A(n851), .B(n852), .Z(n845) );
  AND U734 ( .A(n241), .B(n844), .Z(n852) );
  XNOR U735 ( .A(n842), .B(n851), .Z(n844) );
  XNOR U736 ( .A(n853), .B(n854), .Z(n842) );
  AND U737 ( .A(n245), .B(n855), .Z(n854) );
  XOR U738 ( .A(p_input[198]), .B(n853), .Z(n855) );
  XNOR U739 ( .A(n856), .B(n857), .Z(n853) );
  AND U740 ( .A(n249), .B(n858), .Z(n857) );
  XOR U741 ( .A(n859), .B(n860), .Z(n851) );
  AND U742 ( .A(n253), .B(n861), .Z(n860) );
  XOR U743 ( .A(n862), .B(n863), .Z(n848) );
  AND U744 ( .A(n257), .B(n861), .Z(n863) );
  XNOR U745 ( .A(n864), .B(n862), .Z(n861) );
  IV U746 ( .A(n859), .Z(n864) );
  XOR U747 ( .A(n865), .B(n866), .Z(n859) );
  AND U748 ( .A(n260), .B(n858), .Z(n866) );
  XNOR U749 ( .A(n856), .B(n865), .Z(n858) );
  XNOR U750 ( .A(n867), .B(n868), .Z(n856) );
  AND U751 ( .A(n264), .B(n869), .Z(n868) );
  XOR U752 ( .A(p_input[230]), .B(n867), .Z(n869) );
  XNOR U753 ( .A(n870), .B(n871), .Z(n867) );
  AND U754 ( .A(n268), .B(n872), .Z(n871) );
  XOR U755 ( .A(n873), .B(n874), .Z(n865) );
  AND U756 ( .A(n272), .B(n875), .Z(n874) );
  XOR U757 ( .A(n876), .B(n877), .Z(n862) );
  AND U758 ( .A(n276), .B(n875), .Z(n877) );
  XNOR U759 ( .A(n878), .B(n876), .Z(n875) );
  IV U760 ( .A(n873), .Z(n878) );
  XOR U761 ( .A(n879), .B(n880), .Z(n873) );
  AND U762 ( .A(n279), .B(n872), .Z(n880) );
  XNOR U763 ( .A(n870), .B(n879), .Z(n872) );
  XNOR U764 ( .A(n881), .B(n882), .Z(n870) );
  AND U765 ( .A(n283), .B(n883), .Z(n882) );
  XOR U766 ( .A(p_input[262]), .B(n881), .Z(n883) );
  XNOR U767 ( .A(n884), .B(n885), .Z(n881) );
  AND U768 ( .A(n287), .B(n886), .Z(n885) );
  XOR U769 ( .A(n887), .B(n888), .Z(n879) );
  AND U770 ( .A(n291), .B(n889), .Z(n888) );
  XOR U771 ( .A(n890), .B(n891), .Z(n876) );
  AND U772 ( .A(n295), .B(n889), .Z(n891) );
  XNOR U773 ( .A(n892), .B(n890), .Z(n889) );
  IV U774 ( .A(n887), .Z(n892) );
  XOR U775 ( .A(n893), .B(n894), .Z(n887) );
  AND U776 ( .A(n298), .B(n886), .Z(n894) );
  XNOR U777 ( .A(n884), .B(n893), .Z(n886) );
  XNOR U778 ( .A(n895), .B(n896), .Z(n884) );
  AND U779 ( .A(n302), .B(n897), .Z(n896) );
  XOR U780 ( .A(p_input[294]), .B(n895), .Z(n897) );
  XNOR U781 ( .A(n898), .B(n899), .Z(n895) );
  AND U782 ( .A(n306), .B(n900), .Z(n899) );
  XOR U783 ( .A(n901), .B(n902), .Z(n893) );
  AND U784 ( .A(n310), .B(n903), .Z(n902) );
  XOR U785 ( .A(n904), .B(n905), .Z(n890) );
  AND U786 ( .A(n314), .B(n903), .Z(n905) );
  XNOR U787 ( .A(n906), .B(n904), .Z(n903) );
  IV U788 ( .A(n901), .Z(n906) );
  XOR U789 ( .A(n907), .B(n908), .Z(n901) );
  AND U790 ( .A(n317), .B(n900), .Z(n908) );
  XNOR U791 ( .A(n898), .B(n907), .Z(n900) );
  XNOR U792 ( .A(n909), .B(n910), .Z(n898) );
  AND U793 ( .A(n321), .B(n911), .Z(n910) );
  XOR U794 ( .A(p_input[326]), .B(n909), .Z(n911) );
  XNOR U795 ( .A(n912), .B(n913), .Z(n909) );
  AND U796 ( .A(n325), .B(n914), .Z(n913) );
  XOR U797 ( .A(n915), .B(n916), .Z(n907) );
  AND U798 ( .A(n329), .B(n917), .Z(n916) );
  XOR U799 ( .A(n918), .B(n919), .Z(n904) );
  AND U800 ( .A(n333), .B(n917), .Z(n919) );
  XNOR U801 ( .A(n920), .B(n918), .Z(n917) );
  IV U802 ( .A(n915), .Z(n920) );
  XOR U803 ( .A(n921), .B(n922), .Z(n915) );
  AND U804 ( .A(n336), .B(n914), .Z(n922) );
  XNOR U805 ( .A(n912), .B(n921), .Z(n914) );
  XNOR U806 ( .A(n923), .B(n924), .Z(n912) );
  AND U807 ( .A(n340), .B(n925), .Z(n924) );
  XOR U808 ( .A(p_input[358]), .B(n923), .Z(n925) );
  XNOR U809 ( .A(n926), .B(n927), .Z(n923) );
  AND U810 ( .A(n344), .B(n928), .Z(n927) );
  XOR U811 ( .A(n929), .B(n930), .Z(n921) );
  AND U812 ( .A(n348), .B(n931), .Z(n930) );
  XOR U813 ( .A(n932), .B(n933), .Z(n918) );
  AND U814 ( .A(n352), .B(n931), .Z(n933) );
  XNOR U815 ( .A(n934), .B(n932), .Z(n931) );
  IV U816 ( .A(n929), .Z(n934) );
  XOR U817 ( .A(n935), .B(n936), .Z(n929) );
  AND U818 ( .A(n355), .B(n928), .Z(n936) );
  XNOR U819 ( .A(n926), .B(n935), .Z(n928) );
  XNOR U820 ( .A(n937), .B(n938), .Z(n926) );
  AND U821 ( .A(n359), .B(n939), .Z(n938) );
  XOR U822 ( .A(p_input[390]), .B(n937), .Z(n939) );
  XOR U823 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(n940), .Z(
        n937) );
  AND U824 ( .A(n362), .B(n941), .Z(n940) );
  XOR U825 ( .A(n942), .B(n943), .Z(n935) );
  AND U826 ( .A(n366), .B(n944), .Z(n943) );
  XOR U827 ( .A(n945), .B(n946), .Z(n932) );
  AND U828 ( .A(n370), .B(n944), .Z(n946) );
  XNOR U829 ( .A(n947), .B(n945), .Z(n944) );
  IV U830 ( .A(n942), .Z(n947) );
  XOR U831 ( .A(n948), .B(n949), .Z(n942) );
  AND U832 ( .A(n373), .B(n941), .Z(n949) );
  XOR U833 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(n948), .Z(
        n941) );
  XOR U834 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .B(n950), .Z(
        n948) );
  AND U835 ( .A(n375), .B(n951), .Z(n950) );
  XOR U836 ( .A(\knn_comb_/min_val_out[0][6] ), .B(n952), .Z(n945) );
  AND U837 ( .A(n378), .B(n951), .Z(n952) );
  XOR U838 ( .A(\knn_comb_/min_val_out[0][6] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .Z(n951) );
  XOR U839 ( .A(n81), .B(n953), .Z(o[37]) );
  AND U840 ( .A(n122), .B(n954), .Z(n81) );
  XOR U841 ( .A(n82), .B(n953), .Z(n954) );
  XOR U842 ( .A(n955), .B(n61), .Z(n953) );
  AND U843 ( .A(n125), .B(n956), .Z(n61) );
  XOR U844 ( .A(n62), .B(n955), .Z(n956) );
  XOR U845 ( .A(n957), .B(n958), .Z(n62) );
  AND U846 ( .A(n130), .B(n959), .Z(n958) );
  XOR U847 ( .A(p_input[5]), .B(n957), .Z(n959) );
  XNOR U848 ( .A(n960), .B(n961), .Z(n957) );
  AND U849 ( .A(n134), .B(n962), .Z(n961) );
  XOR U850 ( .A(n963), .B(n964), .Z(n955) );
  AND U851 ( .A(n138), .B(n965), .Z(n964) );
  XOR U852 ( .A(n966), .B(n967), .Z(n82) );
  AND U853 ( .A(n142), .B(n965), .Z(n967) );
  XNOR U854 ( .A(n968), .B(n966), .Z(n965) );
  IV U855 ( .A(n963), .Z(n968) );
  XOR U856 ( .A(n969), .B(n970), .Z(n963) );
  AND U857 ( .A(n146), .B(n962), .Z(n970) );
  XNOR U858 ( .A(n960), .B(n969), .Z(n962) );
  XNOR U859 ( .A(n971), .B(n972), .Z(n960) );
  AND U860 ( .A(n150), .B(n973), .Z(n972) );
  XOR U861 ( .A(p_input[37]), .B(n971), .Z(n973) );
  XNOR U862 ( .A(n974), .B(n975), .Z(n971) );
  AND U863 ( .A(n154), .B(n976), .Z(n975) );
  XOR U864 ( .A(n977), .B(n978), .Z(n969) );
  AND U865 ( .A(n158), .B(n979), .Z(n978) );
  XOR U866 ( .A(n980), .B(n981), .Z(n966) );
  AND U867 ( .A(n162), .B(n979), .Z(n981) );
  XNOR U868 ( .A(n982), .B(n980), .Z(n979) );
  IV U869 ( .A(n977), .Z(n982) );
  XOR U870 ( .A(n983), .B(n984), .Z(n977) );
  AND U871 ( .A(n165), .B(n976), .Z(n984) );
  XNOR U872 ( .A(n974), .B(n983), .Z(n976) );
  XNOR U873 ( .A(n985), .B(n986), .Z(n974) );
  AND U874 ( .A(n169), .B(n987), .Z(n986) );
  XOR U875 ( .A(p_input[69]), .B(n985), .Z(n987) );
  XNOR U876 ( .A(n988), .B(n989), .Z(n985) );
  AND U877 ( .A(n173), .B(n990), .Z(n989) );
  XOR U878 ( .A(n991), .B(n992), .Z(n983) );
  AND U879 ( .A(n177), .B(n993), .Z(n992) );
  XOR U880 ( .A(n994), .B(n995), .Z(n980) );
  AND U881 ( .A(n181), .B(n993), .Z(n995) );
  XNOR U882 ( .A(n996), .B(n994), .Z(n993) );
  IV U883 ( .A(n991), .Z(n996) );
  XOR U884 ( .A(n997), .B(n998), .Z(n991) );
  AND U885 ( .A(n184), .B(n990), .Z(n998) );
  XNOR U886 ( .A(n988), .B(n997), .Z(n990) );
  XNOR U887 ( .A(n999), .B(n1000), .Z(n988) );
  AND U888 ( .A(n188), .B(n1001), .Z(n1000) );
  XOR U889 ( .A(p_input[101]), .B(n999), .Z(n1001) );
  XNOR U890 ( .A(n1002), .B(n1003), .Z(n999) );
  AND U891 ( .A(n192), .B(n1004), .Z(n1003) );
  XOR U892 ( .A(n1005), .B(n1006), .Z(n997) );
  AND U893 ( .A(n196), .B(n1007), .Z(n1006) );
  XOR U894 ( .A(n1008), .B(n1009), .Z(n994) );
  AND U895 ( .A(n200), .B(n1007), .Z(n1009) );
  XNOR U896 ( .A(n1010), .B(n1008), .Z(n1007) );
  IV U897 ( .A(n1005), .Z(n1010) );
  XOR U898 ( .A(n1011), .B(n1012), .Z(n1005) );
  AND U899 ( .A(n203), .B(n1004), .Z(n1012) );
  XNOR U900 ( .A(n1002), .B(n1011), .Z(n1004) );
  XNOR U901 ( .A(n1013), .B(n1014), .Z(n1002) );
  AND U902 ( .A(n207), .B(n1015), .Z(n1014) );
  XOR U903 ( .A(p_input[133]), .B(n1013), .Z(n1015) );
  XNOR U904 ( .A(n1016), .B(n1017), .Z(n1013) );
  AND U905 ( .A(n211), .B(n1018), .Z(n1017) );
  XOR U906 ( .A(n1019), .B(n1020), .Z(n1011) );
  AND U907 ( .A(n215), .B(n1021), .Z(n1020) );
  XOR U908 ( .A(n1022), .B(n1023), .Z(n1008) );
  AND U909 ( .A(n219), .B(n1021), .Z(n1023) );
  XNOR U910 ( .A(n1024), .B(n1022), .Z(n1021) );
  IV U911 ( .A(n1019), .Z(n1024) );
  XOR U912 ( .A(n1025), .B(n1026), .Z(n1019) );
  AND U913 ( .A(n222), .B(n1018), .Z(n1026) );
  XNOR U914 ( .A(n1016), .B(n1025), .Z(n1018) );
  XNOR U915 ( .A(n1027), .B(n1028), .Z(n1016) );
  AND U916 ( .A(n226), .B(n1029), .Z(n1028) );
  XOR U917 ( .A(p_input[165]), .B(n1027), .Z(n1029) );
  XNOR U918 ( .A(n1030), .B(n1031), .Z(n1027) );
  AND U919 ( .A(n230), .B(n1032), .Z(n1031) );
  XOR U920 ( .A(n1033), .B(n1034), .Z(n1025) );
  AND U921 ( .A(n234), .B(n1035), .Z(n1034) );
  XOR U922 ( .A(n1036), .B(n1037), .Z(n1022) );
  AND U923 ( .A(n238), .B(n1035), .Z(n1037) );
  XNOR U924 ( .A(n1038), .B(n1036), .Z(n1035) );
  IV U925 ( .A(n1033), .Z(n1038) );
  XOR U926 ( .A(n1039), .B(n1040), .Z(n1033) );
  AND U927 ( .A(n241), .B(n1032), .Z(n1040) );
  XNOR U928 ( .A(n1030), .B(n1039), .Z(n1032) );
  XNOR U929 ( .A(n1041), .B(n1042), .Z(n1030) );
  AND U930 ( .A(n245), .B(n1043), .Z(n1042) );
  XOR U931 ( .A(p_input[197]), .B(n1041), .Z(n1043) );
  XNOR U932 ( .A(n1044), .B(n1045), .Z(n1041) );
  AND U933 ( .A(n249), .B(n1046), .Z(n1045) );
  XOR U934 ( .A(n1047), .B(n1048), .Z(n1039) );
  AND U935 ( .A(n253), .B(n1049), .Z(n1048) );
  XOR U936 ( .A(n1050), .B(n1051), .Z(n1036) );
  AND U937 ( .A(n257), .B(n1049), .Z(n1051) );
  XNOR U938 ( .A(n1052), .B(n1050), .Z(n1049) );
  IV U939 ( .A(n1047), .Z(n1052) );
  XOR U940 ( .A(n1053), .B(n1054), .Z(n1047) );
  AND U941 ( .A(n260), .B(n1046), .Z(n1054) );
  XNOR U942 ( .A(n1044), .B(n1053), .Z(n1046) );
  XNOR U943 ( .A(n1055), .B(n1056), .Z(n1044) );
  AND U944 ( .A(n264), .B(n1057), .Z(n1056) );
  XOR U945 ( .A(p_input[229]), .B(n1055), .Z(n1057) );
  XNOR U946 ( .A(n1058), .B(n1059), .Z(n1055) );
  AND U947 ( .A(n268), .B(n1060), .Z(n1059) );
  XOR U948 ( .A(n1061), .B(n1062), .Z(n1053) );
  AND U949 ( .A(n272), .B(n1063), .Z(n1062) );
  XOR U950 ( .A(n1064), .B(n1065), .Z(n1050) );
  AND U951 ( .A(n276), .B(n1063), .Z(n1065) );
  XNOR U952 ( .A(n1066), .B(n1064), .Z(n1063) );
  IV U953 ( .A(n1061), .Z(n1066) );
  XOR U954 ( .A(n1067), .B(n1068), .Z(n1061) );
  AND U955 ( .A(n279), .B(n1060), .Z(n1068) );
  XNOR U956 ( .A(n1058), .B(n1067), .Z(n1060) );
  XNOR U957 ( .A(n1069), .B(n1070), .Z(n1058) );
  AND U958 ( .A(n283), .B(n1071), .Z(n1070) );
  XOR U959 ( .A(p_input[261]), .B(n1069), .Z(n1071) );
  XNOR U960 ( .A(n1072), .B(n1073), .Z(n1069) );
  AND U961 ( .A(n287), .B(n1074), .Z(n1073) );
  XOR U962 ( .A(n1075), .B(n1076), .Z(n1067) );
  AND U963 ( .A(n291), .B(n1077), .Z(n1076) );
  XOR U964 ( .A(n1078), .B(n1079), .Z(n1064) );
  AND U965 ( .A(n295), .B(n1077), .Z(n1079) );
  XNOR U966 ( .A(n1080), .B(n1078), .Z(n1077) );
  IV U967 ( .A(n1075), .Z(n1080) );
  XOR U968 ( .A(n1081), .B(n1082), .Z(n1075) );
  AND U969 ( .A(n298), .B(n1074), .Z(n1082) );
  XNOR U970 ( .A(n1072), .B(n1081), .Z(n1074) );
  XNOR U971 ( .A(n1083), .B(n1084), .Z(n1072) );
  AND U972 ( .A(n302), .B(n1085), .Z(n1084) );
  XOR U973 ( .A(p_input[293]), .B(n1083), .Z(n1085) );
  XNOR U974 ( .A(n1086), .B(n1087), .Z(n1083) );
  AND U975 ( .A(n306), .B(n1088), .Z(n1087) );
  XOR U976 ( .A(n1089), .B(n1090), .Z(n1081) );
  AND U977 ( .A(n310), .B(n1091), .Z(n1090) );
  XOR U978 ( .A(n1092), .B(n1093), .Z(n1078) );
  AND U979 ( .A(n314), .B(n1091), .Z(n1093) );
  XNOR U980 ( .A(n1094), .B(n1092), .Z(n1091) );
  IV U981 ( .A(n1089), .Z(n1094) );
  XOR U982 ( .A(n1095), .B(n1096), .Z(n1089) );
  AND U983 ( .A(n317), .B(n1088), .Z(n1096) );
  XNOR U984 ( .A(n1086), .B(n1095), .Z(n1088) );
  XNOR U985 ( .A(n1097), .B(n1098), .Z(n1086) );
  AND U986 ( .A(n321), .B(n1099), .Z(n1098) );
  XOR U987 ( .A(p_input[325]), .B(n1097), .Z(n1099) );
  XNOR U988 ( .A(n1100), .B(n1101), .Z(n1097) );
  AND U989 ( .A(n325), .B(n1102), .Z(n1101) );
  XOR U990 ( .A(n1103), .B(n1104), .Z(n1095) );
  AND U991 ( .A(n329), .B(n1105), .Z(n1104) );
  XOR U992 ( .A(n1106), .B(n1107), .Z(n1092) );
  AND U993 ( .A(n333), .B(n1105), .Z(n1107) );
  XNOR U994 ( .A(n1108), .B(n1106), .Z(n1105) );
  IV U995 ( .A(n1103), .Z(n1108) );
  XOR U996 ( .A(n1109), .B(n1110), .Z(n1103) );
  AND U997 ( .A(n336), .B(n1102), .Z(n1110) );
  XNOR U998 ( .A(n1100), .B(n1109), .Z(n1102) );
  XNOR U999 ( .A(n1111), .B(n1112), .Z(n1100) );
  AND U1000 ( .A(n340), .B(n1113), .Z(n1112) );
  XOR U1001 ( .A(p_input[357]), .B(n1111), .Z(n1113) );
  XNOR U1002 ( .A(n1114), .B(n1115), .Z(n1111) );
  AND U1003 ( .A(n344), .B(n1116), .Z(n1115) );
  XOR U1004 ( .A(n1117), .B(n1118), .Z(n1109) );
  AND U1005 ( .A(n348), .B(n1119), .Z(n1118) );
  XOR U1006 ( .A(n1120), .B(n1121), .Z(n1106) );
  AND U1007 ( .A(n352), .B(n1119), .Z(n1121) );
  XNOR U1008 ( .A(n1122), .B(n1120), .Z(n1119) );
  IV U1009 ( .A(n1117), .Z(n1122) );
  XOR U1010 ( .A(n1123), .B(n1124), .Z(n1117) );
  AND U1011 ( .A(n355), .B(n1116), .Z(n1124) );
  XNOR U1012 ( .A(n1114), .B(n1123), .Z(n1116) );
  XNOR U1013 ( .A(n1125), .B(n1126), .Z(n1114) );
  AND U1014 ( .A(n359), .B(n1127), .Z(n1126) );
  XOR U1015 ( .A(p_input[389]), .B(n1125), .Z(n1127) );
  XOR U1016 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n1128), 
        .Z(n1125) );
  AND U1017 ( .A(n362), .B(n1129), .Z(n1128) );
  XOR U1018 ( .A(n1130), .B(n1131), .Z(n1123) );
  AND U1019 ( .A(n366), .B(n1132), .Z(n1131) );
  XOR U1020 ( .A(n1133), .B(n1134), .Z(n1120) );
  AND U1021 ( .A(n370), .B(n1132), .Z(n1134) );
  XNOR U1022 ( .A(n1135), .B(n1133), .Z(n1132) );
  IV U1023 ( .A(n1130), .Z(n1135) );
  XOR U1024 ( .A(n1136), .B(n1137), .Z(n1130) );
  AND U1025 ( .A(n373), .B(n1129), .Z(n1137) );
  XOR U1026 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n1136), 
        .Z(n1129) );
  XOR U1027 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(n1138), 
        .Z(n1136) );
  AND U1028 ( .A(n375), .B(n1139), .Z(n1138) );
  XOR U1029 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n1140), .Z(n1133) );
  AND U1030 ( .A(n378), .B(n1139), .Z(n1140) );
  XOR U1031 ( .A(n1141), .B(n1142), .Z(n1139) );
  IV U1032 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .Z(n1142) );
  IV U1033 ( .A(\knn_comb_/min_val_out[0][5] ), .Z(n1141) );
  XOR U1034 ( .A(n103), .B(n1143), .Z(o[36]) );
  AND U1035 ( .A(n122), .B(n1144), .Z(n103) );
  XOR U1036 ( .A(n104), .B(n1143), .Z(n1144) );
  XOR U1037 ( .A(n1145), .B(n63), .Z(n1143) );
  AND U1038 ( .A(n125), .B(n1146), .Z(n63) );
  XOR U1039 ( .A(n64), .B(n1145), .Z(n1146) );
  XOR U1040 ( .A(n1147), .B(n1148), .Z(n64) );
  AND U1041 ( .A(n130), .B(n1149), .Z(n1148) );
  XOR U1042 ( .A(p_input[4]), .B(n1147), .Z(n1149) );
  XNOR U1043 ( .A(n1150), .B(n1151), .Z(n1147) );
  AND U1044 ( .A(n134), .B(n1152), .Z(n1151) );
  XOR U1045 ( .A(n1153), .B(n1154), .Z(n1145) );
  AND U1046 ( .A(n138), .B(n1155), .Z(n1154) );
  XOR U1047 ( .A(n1156), .B(n1157), .Z(n104) );
  AND U1048 ( .A(n142), .B(n1155), .Z(n1157) );
  XNOR U1049 ( .A(n1158), .B(n1156), .Z(n1155) );
  IV U1050 ( .A(n1153), .Z(n1158) );
  XOR U1051 ( .A(n1159), .B(n1160), .Z(n1153) );
  AND U1052 ( .A(n146), .B(n1152), .Z(n1160) );
  XNOR U1053 ( .A(n1150), .B(n1159), .Z(n1152) );
  XNOR U1054 ( .A(n1161), .B(n1162), .Z(n1150) );
  AND U1055 ( .A(n150), .B(n1163), .Z(n1162) );
  XOR U1056 ( .A(p_input[36]), .B(n1161), .Z(n1163) );
  XNOR U1057 ( .A(n1164), .B(n1165), .Z(n1161) );
  AND U1058 ( .A(n154), .B(n1166), .Z(n1165) );
  XOR U1059 ( .A(n1167), .B(n1168), .Z(n1159) );
  AND U1060 ( .A(n158), .B(n1169), .Z(n1168) );
  XOR U1061 ( .A(n1170), .B(n1171), .Z(n1156) );
  AND U1062 ( .A(n162), .B(n1169), .Z(n1171) );
  XNOR U1063 ( .A(n1172), .B(n1170), .Z(n1169) );
  IV U1064 ( .A(n1167), .Z(n1172) );
  XOR U1065 ( .A(n1173), .B(n1174), .Z(n1167) );
  AND U1066 ( .A(n165), .B(n1166), .Z(n1174) );
  XNOR U1067 ( .A(n1164), .B(n1173), .Z(n1166) );
  XNOR U1068 ( .A(n1175), .B(n1176), .Z(n1164) );
  AND U1069 ( .A(n169), .B(n1177), .Z(n1176) );
  XOR U1070 ( .A(p_input[68]), .B(n1175), .Z(n1177) );
  XNOR U1071 ( .A(n1178), .B(n1179), .Z(n1175) );
  AND U1072 ( .A(n173), .B(n1180), .Z(n1179) );
  XOR U1073 ( .A(n1181), .B(n1182), .Z(n1173) );
  AND U1074 ( .A(n177), .B(n1183), .Z(n1182) );
  XOR U1075 ( .A(n1184), .B(n1185), .Z(n1170) );
  AND U1076 ( .A(n181), .B(n1183), .Z(n1185) );
  XNOR U1077 ( .A(n1186), .B(n1184), .Z(n1183) );
  IV U1078 ( .A(n1181), .Z(n1186) );
  XOR U1079 ( .A(n1187), .B(n1188), .Z(n1181) );
  AND U1080 ( .A(n184), .B(n1180), .Z(n1188) );
  XNOR U1081 ( .A(n1178), .B(n1187), .Z(n1180) );
  XNOR U1082 ( .A(n1189), .B(n1190), .Z(n1178) );
  AND U1083 ( .A(n188), .B(n1191), .Z(n1190) );
  XOR U1084 ( .A(p_input[100]), .B(n1189), .Z(n1191) );
  XNOR U1085 ( .A(n1192), .B(n1193), .Z(n1189) );
  AND U1086 ( .A(n192), .B(n1194), .Z(n1193) );
  XOR U1087 ( .A(n1195), .B(n1196), .Z(n1187) );
  AND U1088 ( .A(n196), .B(n1197), .Z(n1196) );
  XOR U1089 ( .A(n1198), .B(n1199), .Z(n1184) );
  AND U1090 ( .A(n200), .B(n1197), .Z(n1199) );
  XNOR U1091 ( .A(n1200), .B(n1198), .Z(n1197) );
  IV U1092 ( .A(n1195), .Z(n1200) );
  XOR U1093 ( .A(n1201), .B(n1202), .Z(n1195) );
  AND U1094 ( .A(n203), .B(n1194), .Z(n1202) );
  XNOR U1095 ( .A(n1192), .B(n1201), .Z(n1194) );
  XNOR U1096 ( .A(n1203), .B(n1204), .Z(n1192) );
  AND U1097 ( .A(n207), .B(n1205), .Z(n1204) );
  XOR U1098 ( .A(p_input[132]), .B(n1203), .Z(n1205) );
  XNOR U1099 ( .A(n1206), .B(n1207), .Z(n1203) );
  AND U1100 ( .A(n211), .B(n1208), .Z(n1207) );
  XOR U1101 ( .A(n1209), .B(n1210), .Z(n1201) );
  AND U1102 ( .A(n215), .B(n1211), .Z(n1210) );
  XOR U1103 ( .A(n1212), .B(n1213), .Z(n1198) );
  AND U1104 ( .A(n219), .B(n1211), .Z(n1213) );
  XNOR U1105 ( .A(n1214), .B(n1212), .Z(n1211) );
  IV U1106 ( .A(n1209), .Z(n1214) );
  XOR U1107 ( .A(n1215), .B(n1216), .Z(n1209) );
  AND U1108 ( .A(n222), .B(n1208), .Z(n1216) );
  XNOR U1109 ( .A(n1206), .B(n1215), .Z(n1208) );
  XNOR U1110 ( .A(n1217), .B(n1218), .Z(n1206) );
  AND U1111 ( .A(n226), .B(n1219), .Z(n1218) );
  XOR U1112 ( .A(p_input[164]), .B(n1217), .Z(n1219) );
  XNOR U1113 ( .A(n1220), .B(n1221), .Z(n1217) );
  AND U1114 ( .A(n230), .B(n1222), .Z(n1221) );
  XOR U1115 ( .A(n1223), .B(n1224), .Z(n1215) );
  AND U1116 ( .A(n234), .B(n1225), .Z(n1224) );
  XOR U1117 ( .A(n1226), .B(n1227), .Z(n1212) );
  AND U1118 ( .A(n238), .B(n1225), .Z(n1227) );
  XNOR U1119 ( .A(n1228), .B(n1226), .Z(n1225) );
  IV U1120 ( .A(n1223), .Z(n1228) );
  XOR U1121 ( .A(n1229), .B(n1230), .Z(n1223) );
  AND U1122 ( .A(n241), .B(n1222), .Z(n1230) );
  XNOR U1123 ( .A(n1220), .B(n1229), .Z(n1222) );
  XNOR U1124 ( .A(n1231), .B(n1232), .Z(n1220) );
  AND U1125 ( .A(n245), .B(n1233), .Z(n1232) );
  XOR U1126 ( .A(p_input[196]), .B(n1231), .Z(n1233) );
  XNOR U1127 ( .A(n1234), .B(n1235), .Z(n1231) );
  AND U1128 ( .A(n249), .B(n1236), .Z(n1235) );
  XOR U1129 ( .A(n1237), .B(n1238), .Z(n1229) );
  AND U1130 ( .A(n253), .B(n1239), .Z(n1238) );
  XOR U1131 ( .A(n1240), .B(n1241), .Z(n1226) );
  AND U1132 ( .A(n257), .B(n1239), .Z(n1241) );
  XNOR U1133 ( .A(n1242), .B(n1240), .Z(n1239) );
  IV U1134 ( .A(n1237), .Z(n1242) );
  XOR U1135 ( .A(n1243), .B(n1244), .Z(n1237) );
  AND U1136 ( .A(n260), .B(n1236), .Z(n1244) );
  XNOR U1137 ( .A(n1234), .B(n1243), .Z(n1236) );
  XNOR U1138 ( .A(n1245), .B(n1246), .Z(n1234) );
  AND U1139 ( .A(n264), .B(n1247), .Z(n1246) );
  XOR U1140 ( .A(p_input[228]), .B(n1245), .Z(n1247) );
  XNOR U1141 ( .A(n1248), .B(n1249), .Z(n1245) );
  AND U1142 ( .A(n268), .B(n1250), .Z(n1249) );
  XOR U1143 ( .A(n1251), .B(n1252), .Z(n1243) );
  AND U1144 ( .A(n272), .B(n1253), .Z(n1252) );
  XOR U1145 ( .A(n1254), .B(n1255), .Z(n1240) );
  AND U1146 ( .A(n276), .B(n1253), .Z(n1255) );
  XNOR U1147 ( .A(n1256), .B(n1254), .Z(n1253) );
  IV U1148 ( .A(n1251), .Z(n1256) );
  XOR U1149 ( .A(n1257), .B(n1258), .Z(n1251) );
  AND U1150 ( .A(n279), .B(n1250), .Z(n1258) );
  XNOR U1151 ( .A(n1248), .B(n1257), .Z(n1250) );
  XNOR U1152 ( .A(n1259), .B(n1260), .Z(n1248) );
  AND U1153 ( .A(n283), .B(n1261), .Z(n1260) );
  XOR U1154 ( .A(p_input[260]), .B(n1259), .Z(n1261) );
  XNOR U1155 ( .A(n1262), .B(n1263), .Z(n1259) );
  AND U1156 ( .A(n287), .B(n1264), .Z(n1263) );
  XOR U1157 ( .A(n1265), .B(n1266), .Z(n1257) );
  AND U1158 ( .A(n291), .B(n1267), .Z(n1266) );
  XOR U1159 ( .A(n1268), .B(n1269), .Z(n1254) );
  AND U1160 ( .A(n295), .B(n1267), .Z(n1269) );
  XNOR U1161 ( .A(n1270), .B(n1268), .Z(n1267) );
  IV U1162 ( .A(n1265), .Z(n1270) );
  XOR U1163 ( .A(n1271), .B(n1272), .Z(n1265) );
  AND U1164 ( .A(n298), .B(n1264), .Z(n1272) );
  XNOR U1165 ( .A(n1262), .B(n1271), .Z(n1264) );
  XNOR U1166 ( .A(n1273), .B(n1274), .Z(n1262) );
  AND U1167 ( .A(n302), .B(n1275), .Z(n1274) );
  XOR U1168 ( .A(p_input[292]), .B(n1273), .Z(n1275) );
  XNOR U1169 ( .A(n1276), .B(n1277), .Z(n1273) );
  AND U1170 ( .A(n306), .B(n1278), .Z(n1277) );
  XOR U1171 ( .A(n1279), .B(n1280), .Z(n1271) );
  AND U1172 ( .A(n310), .B(n1281), .Z(n1280) );
  XOR U1173 ( .A(n1282), .B(n1283), .Z(n1268) );
  AND U1174 ( .A(n314), .B(n1281), .Z(n1283) );
  XNOR U1175 ( .A(n1284), .B(n1282), .Z(n1281) );
  IV U1176 ( .A(n1279), .Z(n1284) );
  XOR U1177 ( .A(n1285), .B(n1286), .Z(n1279) );
  AND U1178 ( .A(n317), .B(n1278), .Z(n1286) );
  XNOR U1179 ( .A(n1276), .B(n1285), .Z(n1278) );
  XNOR U1180 ( .A(n1287), .B(n1288), .Z(n1276) );
  AND U1181 ( .A(n321), .B(n1289), .Z(n1288) );
  XOR U1182 ( .A(p_input[324]), .B(n1287), .Z(n1289) );
  XNOR U1183 ( .A(n1290), .B(n1291), .Z(n1287) );
  AND U1184 ( .A(n325), .B(n1292), .Z(n1291) );
  XOR U1185 ( .A(n1293), .B(n1294), .Z(n1285) );
  AND U1186 ( .A(n329), .B(n1295), .Z(n1294) );
  XOR U1187 ( .A(n1296), .B(n1297), .Z(n1282) );
  AND U1188 ( .A(n333), .B(n1295), .Z(n1297) );
  XNOR U1189 ( .A(n1298), .B(n1296), .Z(n1295) );
  IV U1190 ( .A(n1293), .Z(n1298) );
  XOR U1191 ( .A(n1299), .B(n1300), .Z(n1293) );
  AND U1192 ( .A(n336), .B(n1292), .Z(n1300) );
  XNOR U1193 ( .A(n1290), .B(n1299), .Z(n1292) );
  XNOR U1194 ( .A(n1301), .B(n1302), .Z(n1290) );
  AND U1195 ( .A(n340), .B(n1303), .Z(n1302) );
  XOR U1196 ( .A(p_input[356]), .B(n1301), .Z(n1303) );
  XNOR U1197 ( .A(n1304), .B(n1305), .Z(n1301) );
  AND U1198 ( .A(n344), .B(n1306), .Z(n1305) );
  XOR U1199 ( .A(n1307), .B(n1308), .Z(n1299) );
  AND U1200 ( .A(n348), .B(n1309), .Z(n1308) );
  XOR U1201 ( .A(n1310), .B(n1311), .Z(n1296) );
  AND U1202 ( .A(n352), .B(n1309), .Z(n1311) );
  XNOR U1203 ( .A(n1312), .B(n1310), .Z(n1309) );
  IV U1204 ( .A(n1307), .Z(n1312) );
  XOR U1205 ( .A(n1313), .B(n1314), .Z(n1307) );
  AND U1206 ( .A(n355), .B(n1306), .Z(n1314) );
  XNOR U1207 ( .A(n1304), .B(n1313), .Z(n1306) );
  XNOR U1208 ( .A(n1315), .B(n1316), .Z(n1304) );
  AND U1209 ( .A(n359), .B(n1317), .Z(n1316) );
  XOR U1210 ( .A(p_input[388]), .B(n1315), .Z(n1317) );
  XOR U1211 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(n1318), 
        .Z(n1315) );
  AND U1212 ( .A(n362), .B(n1319), .Z(n1318) );
  XOR U1213 ( .A(n1320), .B(n1321), .Z(n1313) );
  AND U1214 ( .A(n366), .B(n1322), .Z(n1321) );
  XOR U1215 ( .A(n1323), .B(n1324), .Z(n1310) );
  AND U1216 ( .A(n370), .B(n1322), .Z(n1324) );
  XNOR U1217 ( .A(n1325), .B(n1323), .Z(n1322) );
  IV U1218 ( .A(n1320), .Z(n1325) );
  XOR U1219 ( .A(n1326), .B(n1327), .Z(n1320) );
  AND U1220 ( .A(n373), .B(n1319), .Z(n1327) );
  XOR U1221 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(n1326), 
        .Z(n1319) );
  XOR U1222 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(n1328), 
        .Z(n1326) );
  AND U1223 ( .A(n375), .B(n1329), .Z(n1328) );
  XOR U1224 ( .A(\knn_comb_/min_val_out[0][4] ), .B(n1330), .Z(n1323) );
  AND U1225 ( .A(n378), .B(n1329), .Z(n1330) );
  XOR U1226 ( .A(\knn_comb_/min_val_out[0][4] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .Z(n1329) );
  XOR U1227 ( .A(n572), .B(n1331), .Z(o[35]) );
  AND U1228 ( .A(n122), .B(n1332), .Z(n572) );
  XOR U1229 ( .A(n573), .B(n1331), .Z(n1332) );
  XOR U1230 ( .A(n1333), .B(n65), .Z(n1331) );
  AND U1231 ( .A(n125), .B(n1334), .Z(n65) );
  XOR U1232 ( .A(n66), .B(n1333), .Z(n1334) );
  XOR U1233 ( .A(n1335), .B(n1336), .Z(n66) );
  AND U1234 ( .A(n130), .B(n1337), .Z(n1336) );
  XOR U1235 ( .A(p_input[3]), .B(n1335), .Z(n1337) );
  XNOR U1236 ( .A(n1338), .B(n1339), .Z(n1335) );
  AND U1237 ( .A(n134), .B(n1340), .Z(n1339) );
  XOR U1238 ( .A(n1341), .B(n1342), .Z(n1333) );
  AND U1239 ( .A(n138), .B(n1343), .Z(n1342) );
  XOR U1240 ( .A(n1344), .B(n1345), .Z(n573) );
  AND U1241 ( .A(n142), .B(n1343), .Z(n1345) );
  XNOR U1242 ( .A(n1346), .B(n1344), .Z(n1343) );
  IV U1243 ( .A(n1341), .Z(n1346) );
  XOR U1244 ( .A(n1347), .B(n1348), .Z(n1341) );
  AND U1245 ( .A(n146), .B(n1340), .Z(n1348) );
  XNOR U1246 ( .A(n1338), .B(n1347), .Z(n1340) );
  XNOR U1247 ( .A(n1349), .B(n1350), .Z(n1338) );
  AND U1248 ( .A(n150), .B(n1351), .Z(n1350) );
  XOR U1249 ( .A(p_input[35]), .B(n1349), .Z(n1351) );
  XNOR U1250 ( .A(n1352), .B(n1353), .Z(n1349) );
  AND U1251 ( .A(n154), .B(n1354), .Z(n1353) );
  XOR U1252 ( .A(n1355), .B(n1356), .Z(n1347) );
  AND U1253 ( .A(n158), .B(n1357), .Z(n1356) );
  XOR U1254 ( .A(n1358), .B(n1359), .Z(n1344) );
  AND U1255 ( .A(n162), .B(n1357), .Z(n1359) );
  XNOR U1256 ( .A(n1360), .B(n1358), .Z(n1357) );
  IV U1257 ( .A(n1355), .Z(n1360) );
  XOR U1258 ( .A(n1361), .B(n1362), .Z(n1355) );
  AND U1259 ( .A(n165), .B(n1354), .Z(n1362) );
  XNOR U1260 ( .A(n1352), .B(n1361), .Z(n1354) );
  XNOR U1261 ( .A(n1363), .B(n1364), .Z(n1352) );
  AND U1262 ( .A(n169), .B(n1365), .Z(n1364) );
  XOR U1263 ( .A(p_input[67]), .B(n1363), .Z(n1365) );
  XNOR U1264 ( .A(n1366), .B(n1367), .Z(n1363) );
  AND U1265 ( .A(n173), .B(n1368), .Z(n1367) );
  XOR U1266 ( .A(n1369), .B(n1370), .Z(n1361) );
  AND U1267 ( .A(n177), .B(n1371), .Z(n1370) );
  XOR U1268 ( .A(n1372), .B(n1373), .Z(n1358) );
  AND U1269 ( .A(n181), .B(n1371), .Z(n1373) );
  XNOR U1270 ( .A(n1374), .B(n1372), .Z(n1371) );
  IV U1271 ( .A(n1369), .Z(n1374) );
  XOR U1272 ( .A(n1375), .B(n1376), .Z(n1369) );
  AND U1273 ( .A(n184), .B(n1368), .Z(n1376) );
  XNOR U1274 ( .A(n1366), .B(n1375), .Z(n1368) );
  XNOR U1275 ( .A(n1377), .B(n1378), .Z(n1366) );
  AND U1276 ( .A(n188), .B(n1379), .Z(n1378) );
  XOR U1277 ( .A(p_input[99]), .B(n1377), .Z(n1379) );
  XNOR U1278 ( .A(n1380), .B(n1381), .Z(n1377) );
  AND U1279 ( .A(n192), .B(n1382), .Z(n1381) );
  XOR U1280 ( .A(n1383), .B(n1384), .Z(n1375) );
  AND U1281 ( .A(n196), .B(n1385), .Z(n1384) );
  XOR U1282 ( .A(n1386), .B(n1387), .Z(n1372) );
  AND U1283 ( .A(n200), .B(n1385), .Z(n1387) );
  XNOR U1284 ( .A(n1388), .B(n1386), .Z(n1385) );
  IV U1285 ( .A(n1383), .Z(n1388) );
  XOR U1286 ( .A(n1389), .B(n1390), .Z(n1383) );
  AND U1287 ( .A(n203), .B(n1382), .Z(n1390) );
  XNOR U1288 ( .A(n1380), .B(n1389), .Z(n1382) );
  XNOR U1289 ( .A(n1391), .B(n1392), .Z(n1380) );
  AND U1290 ( .A(n207), .B(n1393), .Z(n1392) );
  XOR U1291 ( .A(p_input[131]), .B(n1391), .Z(n1393) );
  XNOR U1292 ( .A(n1394), .B(n1395), .Z(n1391) );
  AND U1293 ( .A(n211), .B(n1396), .Z(n1395) );
  XOR U1294 ( .A(n1397), .B(n1398), .Z(n1389) );
  AND U1295 ( .A(n215), .B(n1399), .Z(n1398) );
  XOR U1296 ( .A(n1400), .B(n1401), .Z(n1386) );
  AND U1297 ( .A(n219), .B(n1399), .Z(n1401) );
  XNOR U1298 ( .A(n1402), .B(n1400), .Z(n1399) );
  IV U1299 ( .A(n1397), .Z(n1402) );
  XOR U1300 ( .A(n1403), .B(n1404), .Z(n1397) );
  AND U1301 ( .A(n222), .B(n1396), .Z(n1404) );
  XNOR U1302 ( .A(n1394), .B(n1403), .Z(n1396) );
  XNOR U1303 ( .A(n1405), .B(n1406), .Z(n1394) );
  AND U1304 ( .A(n226), .B(n1407), .Z(n1406) );
  XOR U1305 ( .A(p_input[163]), .B(n1405), .Z(n1407) );
  XNOR U1306 ( .A(n1408), .B(n1409), .Z(n1405) );
  AND U1307 ( .A(n230), .B(n1410), .Z(n1409) );
  XOR U1308 ( .A(n1411), .B(n1412), .Z(n1403) );
  AND U1309 ( .A(n234), .B(n1413), .Z(n1412) );
  XOR U1310 ( .A(n1414), .B(n1415), .Z(n1400) );
  AND U1311 ( .A(n238), .B(n1413), .Z(n1415) );
  XNOR U1312 ( .A(n1416), .B(n1414), .Z(n1413) );
  IV U1313 ( .A(n1411), .Z(n1416) );
  XOR U1314 ( .A(n1417), .B(n1418), .Z(n1411) );
  AND U1315 ( .A(n241), .B(n1410), .Z(n1418) );
  XNOR U1316 ( .A(n1408), .B(n1417), .Z(n1410) );
  XNOR U1317 ( .A(n1419), .B(n1420), .Z(n1408) );
  AND U1318 ( .A(n245), .B(n1421), .Z(n1420) );
  XOR U1319 ( .A(p_input[195]), .B(n1419), .Z(n1421) );
  XNOR U1320 ( .A(n1422), .B(n1423), .Z(n1419) );
  AND U1321 ( .A(n249), .B(n1424), .Z(n1423) );
  XOR U1322 ( .A(n1425), .B(n1426), .Z(n1417) );
  AND U1323 ( .A(n253), .B(n1427), .Z(n1426) );
  XOR U1324 ( .A(n1428), .B(n1429), .Z(n1414) );
  AND U1325 ( .A(n257), .B(n1427), .Z(n1429) );
  XNOR U1326 ( .A(n1430), .B(n1428), .Z(n1427) );
  IV U1327 ( .A(n1425), .Z(n1430) );
  XOR U1328 ( .A(n1431), .B(n1432), .Z(n1425) );
  AND U1329 ( .A(n260), .B(n1424), .Z(n1432) );
  XNOR U1330 ( .A(n1422), .B(n1431), .Z(n1424) );
  XNOR U1331 ( .A(n1433), .B(n1434), .Z(n1422) );
  AND U1332 ( .A(n264), .B(n1435), .Z(n1434) );
  XOR U1333 ( .A(p_input[227]), .B(n1433), .Z(n1435) );
  XNOR U1334 ( .A(n1436), .B(n1437), .Z(n1433) );
  AND U1335 ( .A(n268), .B(n1438), .Z(n1437) );
  XOR U1336 ( .A(n1439), .B(n1440), .Z(n1431) );
  AND U1337 ( .A(n272), .B(n1441), .Z(n1440) );
  XOR U1338 ( .A(n1442), .B(n1443), .Z(n1428) );
  AND U1339 ( .A(n276), .B(n1441), .Z(n1443) );
  XNOR U1340 ( .A(n1444), .B(n1442), .Z(n1441) );
  IV U1341 ( .A(n1439), .Z(n1444) );
  XOR U1342 ( .A(n1445), .B(n1446), .Z(n1439) );
  AND U1343 ( .A(n279), .B(n1438), .Z(n1446) );
  XNOR U1344 ( .A(n1436), .B(n1445), .Z(n1438) );
  XNOR U1345 ( .A(n1447), .B(n1448), .Z(n1436) );
  AND U1346 ( .A(n283), .B(n1449), .Z(n1448) );
  XOR U1347 ( .A(p_input[259]), .B(n1447), .Z(n1449) );
  XNOR U1348 ( .A(n1450), .B(n1451), .Z(n1447) );
  AND U1349 ( .A(n287), .B(n1452), .Z(n1451) );
  XOR U1350 ( .A(n1453), .B(n1454), .Z(n1445) );
  AND U1351 ( .A(n291), .B(n1455), .Z(n1454) );
  XOR U1352 ( .A(n1456), .B(n1457), .Z(n1442) );
  AND U1353 ( .A(n295), .B(n1455), .Z(n1457) );
  XNOR U1354 ( .A(n1458), .B(n1456), .Z(n1455) );
  IV U1355 ( .A(n1453), .Z(n1458) );
  XOR U1356 ( .A(n1459), .B(n1460), .Z(n1453) );
  AND U1357 ( .A(n298), .B(n1452), .Z(n1460) );
  XNOR U1358 ( .A(n1450), .B(n1459), .Z(n1452) );
  XNOR U1359 ( .A(n1461), .B(n1462), .Z(n1450) );
  AND U1360 ( .A(n302), .B(n1463), .Z(n1462) );
  XOR U1361 ( .A(p_input[291]), .B(n1461), .Z(n1463) );
  XNOR U1362 ( .A(n1464), .B(n1465), .Z(n1461) );
  AND U1363 ( .A(n306), .B(n1466), .Z(n1465) );
  XOR U1364 ( .A(n1467), .B(n1468), .Z(n1459) );
  AND U1365 ( .A(n310), .B(n1469), .Z(n1468) );
  XOR U1366 ( .A(n1470), .B(n1471), .Z(n1456) );
  AND U1367 ( .A(n314), .B(n1469), .Z(n1471) );
  XNOR U1368 ( .A(n1472), .B(n1470), .Z(n1469) );
  IV U1369 ( .A(n1467), .Z(n1472) );
  XOR U1370 ( .A(n1473), .B(n1474), .Z(n1467) );
  AND U1371 ( .A(n317), .B(n1466), .Z(n1474) );
  XNOR U1372 ( .A(n1464), .B(n1473), .Z(n1466) );
  XNOR U1373 ( .A(n1475), .B(n1476), .Z(n1464) );
  AND U1374 ( .A(n321), .B(n1477), .Z(n1476) );
  XOR U1375 ( .A(p_input[323]), .B(n1475), .Z(n1477) );
  XNOR U1376 ( .A(n1478), .B(n1479), .Z(n1475) );
  AND U1377 ( .A(n325), .B(n1480), .Z(n1479) );
  XOR U1378 ( .A(n1481), .B(n1482), .Z(n1473) );
  AND U1379 ( .A(n329), .B(n1483), .Z(n1482) );
  XOR U1380 ( .A(n1484), .B(n1485), .Z(n1470) );
  AND U1381 ( .A(n333), .B(n1483), .Z(n1485) );
  XNOR U1382 ( .A(n1486), .B(n1484), .Z(n1483) );
  IV U1383 ( .A(n1481), .Z(n1486) );
  XOR U1384 ( .A(n1487), .B(n1488), .Z(n1481) );
  AND U1385 ( .A(n336), .B(n1480), .Z(n1488) );
  XNOR U1386 ( .A(n1478), .B(n1487), .Z(n1480) );
  XNOR U1387 ( .A(n1489), .B(n1490), .Z(n1478) );
  AND U1388 ( .A(n340), .B(n1491), .Z(n1490) );
  XOR U1389 ( .A(p_input[355]), .B(n1489), .Z(n1491) );
  XNOR U1390 ( .A(n1492), .B(n1493), .Z(n1489) );
  AND U1391 ( .A(n344), .B(n1494), .Z(n1493) );
  XOR U1392 ( .A(n1495), .B(n1496), .Z(n1487) );
  AND U1393 ( .A(n348), .B(n1497), .Z(n1496) );
  XOR U1394 ( .A(n1498), .B(n1499), .Z(n1484) );
  AND U1395 ( .A(n352), .B(n1497), .Z(n1499) );
  XNOR U1396 ( .A(n1500), .B(n1498), .Z(n1497) );
  IV U1397 ( .A(n1495), .Z(n1500) );
  XOR U1398 ( .A(n1501), .B(n1502), .Z(n1495) );
  AND U1399 ( .A(n355), .B(n1494), .Z(n1502) );
  XNOR U1400 ( .A(n1492), .B(n1501), .Z(n1494) );
  XNOR U1401 ( .A(n1503), .B(n1504), .Z(n1492) );
  AND U1402 ( .A(n359), .B(n1505), .Z(n1504) );
  XOR U1403 ( .A(p_input[387]), .B(n1503), .Z(n1505) );
  XOR U1404 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(n1506), 
        .Z(n1503) );
  AND U1405 ( .A(n362), .B(n1507), .Z(n1506) );
  XOR U1406 ( .A(n1508), .B(n1509), .Z(n1501) );
  AND U1407 ( .A(n366), .B(n1510), .Z(n1509) );
  XOR U1408 ( .A(n1511), .B(n1512), .Z(n1498) );
  AND U1409 ( .A(n370), .B(n1510), .Z(n1512) );
  XNOR U1410 ( .A(n1513), .B(n1511), .Z(n1510) );
  IV U1411 ( .A(n1508), .Z(n1513) );
  XOR U1412 ( .A(n1514), .B(n1515), .Z(n1508) );
  AND U1413 ( .A(n373), .B(n1507), .Z(n1515) );
  XOR U1414 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(n1514), 
        .Z(n1507) );
  XOR U1415 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .B(n1516), 
        .Z(n1514) );
  AND U1416 ( .A(n375), .B(n1517), .Z(n1516) );
  XOR U1417 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n1518), .Z(n1511) );
  AND U1418 ( .A(n378), .B(n1517), .Z(n1518) );
  XOR U1419 ( .A(\knn_comb_/min_val_out[0][3] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .Z(n1517) );
  XOR U1420 ( .A(n1519), .B(n1520), .Z(o[34]) );
  XOR U1421 ( .A(n1521), .B(n1522), .Z(o[33]) );
  XOR U1422 ( .A(n1523), .B(n1524), .Z(o[32]) );
  XOR U1423 ( .A(n73), .B(n1525), .Z(o[31]) );
  AND U1424 ( .A(n122), .B(n1526), .Z(n73) );
  XOR U1425 ( .A(n74), .B(n1525), .Z(n1526) );
  XOR U1426 ( .A(n1527), .B(n1528), .Z(n1525) );
  AND U1427 ( .A(n142), .B(n1529), .Z(n1528) );
  XOR U1428 ( .A(n1530), .B(n3), .Z(n74) );
  AND U1429 ( .A(n125), .B(n1531), .Z(n3) );
  XOR U1430 ( .A(n4), .B(n1530), .Z(n1531) );
  XOR U1431 ( .A(n1532), .B(n1533), .Z(n4) );
  AND U1432 ( .A(n130), .B(n1534), .Z(n1533) );
  XOR U1433 ( .A(p_input[31]), .B(n1532), .Z(n1534) );
  XNOR U1434 ( .A(n1535), .B(n1536), .Z(n1532) );
  AND U1435 ( .A(n134), .B(n1537), .Z(n1536) );
  XOR U1436 ( .A(n1538), .B(n1539), .Z(n1530) );
  AND U1437 ( .A(n138), .B(n1529), .Z(n1539) );
  XNOR U1438 ( .A(n1540), .B(n1527), .Z(n1529) );
  XOR U1439 ( .A(n1541), .B(n1542), .Z(n1527) );
  AND U1440 ( .A(n162), .B(n1543), .Z(n1542) );
  IV U1441 ( .A(n1538), .Z(n1540) );
  XOR U1442 ( .A(n1544), .B(n1545), .Z(n1538) );
  AND U1443 ( .A(n146), .B(n1537), .Z(n1545) );
  XNOR U1444 ( .A(n1535), .B(n1544), .Z(n1537) );
  XNOR U1445 ( .A(n1546), .B(n1547), .Z(n1535) );
  AND U1446 ( .A(n150), .B(n1548), .Z(n1547) );
  XOR U1447 ( .A(p_input[63]), .B(n1546), .Z(n1548) );
  XNOR U1448 ( .A(n1549), .B(n1550), .Z(n1546) );
  AND U1449 ( .A(n154), .B(n1551), .Z(n1550) );
  XOR U1450 ( .A(n1552), .B(n1553), .Z(n1544) );
  AND U1451 ( .A(n158), .B(n1543), .Z(n1553) );
  XNOR U1452 ( .A(n1554), .B(n1541), .Z(n1543) );
  XOR U1453 ( .A(n1555), .B(n1556), .Z(n1541) );
  AND U1454 ( .A(n181), .B(n1557), .Z(n1556) );
  IV U1455 ( .A(n1552), .Z(n1554) );
  XOR U1456 ( .A(n1558), .B(n1559), .Z(n1552) );
  AND U1457 ( .A(n165), .B(n1551), .Z(n1559) );
  XNOR U1458 ( .A(n1549), .B(n1558), .Z(n1551) );
  XNOR U1459 ( .A(n1560), .B(n1561), .Z(n1549) );
  AND U1460 ( .A(n169), .B(n1562), .Z(n1561) );
  XOR U1461 ( .A(p_input[95]), .B(n1560), .Z(n1562) );
  XNOR U1462 ( .A(n1563), .B(n1564), .Z(n1560) );
  AND U1463 ( .A(n173), .B(n1565), .Z(n1564) );
  XOR U1464 ( .A(n1566), .B(n1567), .Z(n1558) );
  AND U1465 ( .A(n177), .B(n1557), .Z(n1567) );
  XNOR U1466 ( .A(n1568), .B(n1555), .Z(n1557) );
  XOR U1467 ( .A(n1569), .B(n1570), .Z(n1555) );
  AND U1468 ( .A(n200), .B(n1571), .Z(n1570) );
  IV U1469 ( .A(n1566), .Z(n1568) );
  XOR U1470 ( .A(n1572), .B(n1573), .Z(n1566) );
  AND U1471 ( .A(n184), .B(n1565), .Z(n1573) );
  XNOR U1472 ( .A(n1563), .B(n1572), .Z(n1565) );
  XNOR U1473 ( .A(n1574), .B(n1575), .Z(n1563) );
  AND U1474 ( .A(n188), .B(n1576), .Z(n1575) );
  XOR U1475 ( .A(p_input[127]), .B(n1574), .Z(n1576) );
  XNOR U1476 ( .A(n1577), .B(n1578), .Z(n1574) );
  AND U1477 ( .A(n192), .B(n1579), .Z(n1578) );
  XOR U1478 ( .A(n1580), .B(n1581), .Z(n1572) );
  AND U1479 ( .A(n196), .B(n1571), .Z(n1581) );
  XNOR U1480 ( .A(n1582), .B(n1569), .Z(n1571) );
  XOR U1481 ( .A(n1583), .B(n1584), .Z(n1569) );
  AND U1482 ( .A(n219), .B(n1585), .Z(n1584) );
  IV U1483 ( .A(n1580), .Z(n1582) );
  XOR U1484 ( .A(n1586), .B(n1587), .Z(n1580) );
  AND U1485 ( .A(n203), .B(n1579), .Z(n1587) );
  XNOR U1486 ( .A(n1577), .B(n1586), .Z(n1579) );
  XNOR U1487 ( .A(n1588), .B(n1589), .Z(n1577) );
  AND U1488 ( .A(n207), .B(n1590), .Z(n1589) );
  XOR U1489 ( .A(p_input[159]), .B(n1588), .Z(n1590) );
  XNOR U1490 ( .A(n1591), .B(n1592), .Z(n1588) );
  AND U1491 ( .A(n211), .B(n1593), .Z(n1592) );
  XOR U1492 ( .A(n1594), .B(n1595), .Z(n1586) );
  AND U1493 ( .A(n215), .B(n1585), .Z(n1595) );
  XNOR U1494 ( .A(n1596), .B(n1583), .Z(n1585) );
  XOR U1495 ( .A(n1597), .B(n1598), .Z(n1583) );
  AND U1496 ( .A(n238), .B(n1599), .Z(n1598) );
  IV U1497 ( .A(n1594), .Z(n1596) );
  XOR U1498 ( .A(n1600), .B(n1601), .Z(n1594) );
  AND U1499 ( .A(n222), .B(n1593), .Z(n1601) );
  XNOR U1500 ( .A(n1591), .B(n1600), .Z(n1593) );
  XNOR U1501 ( .A(n1602), .B(n1603), .Z(n1591) );
  AND U1502 ( .A(n226), .B(n1604), .Z(n1603) );
  XOR U1503 ( .A(p_input[191]), .B(n1602), .Z(n1604) );
  XNOR U1504 ( .A(n1605), .B(n1606), .Z(n1602) );
  AND U1505 ( .A(n230), .B(n1607), .Z(n1606) );
  XOR U1506 ( .A(n1608), .B(n1609), .Z(n1600) );
  AND U1507 ( .A(n234), .B(n1599), .Z(n1609) );
  XNOR U1508 ( .A(n1610), .B(n1597), .Z(n1599) );
  XOR U1509 ( .A(n1611), .B(n1612), .Z(n1597) );
  AND U1510 ( .A(n257), .B(n1613), .Z(n1612) );
  IV U1511 ( .A(n1608), .Z(n1610) );
  XOR U1512 ( .A(n1614), .B(n1615), .Z(n1608) );
  AND U1513 ( .A(n241), .B(n1607), .Z(n1615) );
  XNOR U1514 ( .A(n1605), .B(n1614), .Z(n1607) );
  XNOR U1515 ( .A(n1616), .B(n1617), .Z(n1605) );
  AND U1516 ( .A(n245), .B(n1618), .Z(n1617) );
  XOR U1517 ( .A(p_input[223]), .B(n1616), .Z(n1618) );
  XNOR U1518 ( .A(n1619), .B(n1620), .Z(n1616) );
  AND U1519 ( .A(n249), .B(n1621), .Z(n1620) );
  XOR U1520 ( .A(n1622), .B(n1623), .Z(n1614) );
  AND U1521 ( .A(n253), .B(n1613), .Z(n1623) );
  XNOR U1522 ( .A(n1624), .B(n1611), .Z(n1613) );
  XOR U1523 ( .A(n1625), .B(n1626), .Z(n1611) );
  AND U1524 ( .A(n276), .B(n1627), .Z(n1626) );
  IV U1525 ( .A(n1622), .Z(n1624) );
  XOR U1526 ( .A(n1628), .B(n1629), .Z(n1622) );
  AND U1527 ( .A(n260), .B(n1621), .Z(n1629) );
  XNOR U1528 ( .A(n1619), .B(n1628), .Z(n1621) );
  XNOR U1529 ( .A(n1630), .B(n1631), .Z(n1619) );
  AND U1530 ( .A(n264), .B(n1632), .Z(n1631) );
  XOR U1531 ( .A(p_input[255]), .B(n1630), .Z(n1632) );
  XNOR U1532 ( .A(n1633), .B(n1634), .Z(n1630) );
  AND U1533 ( .A(n268), .B(n1635), .Z(n1634) );
  XOR U1534 ( .A(n1636), .B(n1637), .Z(n1628) );
  AND U1535 ( .A(n272), .B(n1627), .Z(n1637) );
  XNOR U1536 ( .A(n1638), .B(n1625), .Z(n1627) );
  XOR U1537 ( .A(n1639), .B(n1640), .Z(n1625) );
  AND U1538 ( .A(n295), .B(n1641), .Z(n1640) );
  IV U1539 ( .A(n1636), .Z(n1638) );
  XOR U1540 ( .A(n1642), .B(n1643), .Z(n1636) );
  AND U1541 ( .A(n279), .B(n1635), .Z(n1643) );
  XNOR U1542 ( .A(n1633), .B(n1642), .Z(n1635) );
  XNOR U1543 ( .A(n1644), .B(n1645), .Z(n1633) );
  AND U1544 ( .A(n283), .B(n1646), .Z(n1645) );
  XOR U1545 ( .A(p_input[287]), .B(n1644), .Z(n1646) );
  XNOR U1546 ( .A(n1647), .B(n1648), .Z(n1644) );
  AND U1547 ( .A(n287), .B(n1649), .Z(n1648) );
  XOR U1548 ( .A(n1650), .B(n1651), .Z(n1642) );
  AND U1549 ( .A(n291), .B(n1641), .Z(n1651) );
  XNOR U1550 ( .A(n1652), .B(n1639), .Z(n1641) );
  XOR U1551 ( .A(n1653), .B(n1654), .Z(n1639) );
  AND U1552 ( .A(n314), .B(n1655), .Z(n1654) );
  IV U1553 ( .A(n1650), .Z(n1652) );
  XOR U1554 ( .A(n1656), .B(n1657), .Z(n1650) );
  AND U1555 ( .A(n298), .B(n1649), .Z(n1657) );
  XNOR U1556 ( .A(n1647), .B(n1656), .Z(n1649) );
  XNOR U1557 ( .A(n1658), .B(n1659), .Z(n1647) );
  AND U1558 ( .A(n302), .B(n1660), .Z(n1659) );
  XOR U1559 ( .A(p_input[319]), .B(n1658), .Z(n1660) );
  XNOR U1560 ( .A(n1661), .B(n1662), .Z(n1658) );
  AND U1561 ( .A(n306), .B(n1663), .Z(n1662) );
  XOR U1562 ( .A(n1664), .B(n1665), .Z(n1656) );
  AND U1563 ( .A(n310), .B(n1655), .Z(n1665) );
  XNOR U1564 ( .A(n1666), .B(n1653), .Z(n1655) );
  XOR U1565 ( .A(n1667), .B(n1668), .Z(n1653) );
  AND U1566 ( .A(n333), .B(n1669), .Z(n1668) );
  IV U1567 ( .A(n1664), .Z(n1666) );
  XOR U1568 ( .A(n1670), .B(n1671), .Z(n1664) );
  AND U1569 ( .A(n317), .B(n1663), .Z(n1671) );
  XNOR U1570 ( .A(n1661), .B(n1670), .Z(n1663) );
  XNOR U1571 ( .A(n1672), .B(n1673), .Z(n1661) );
  AND U1572 ( .A(n321), .B(n1674), .Z(n1673) );
  XOR U1573 ( .A(p_input[351]), .B(n1672), .Z(n1674) );
  XNOR U1574 ( .A(n1675), .B(n1676), .Z(n1672) );
  AND U1575 ( .A(n325), .B(n1677), .Z(n1676) );
  XOR U1576 ( .A(n1678), .B(n1679), .Z(n1670) );
  AND U1577 ( .A(n329), .B(n1669), .Z(n1679) );
  XNOR U1578 ( .A(n1680), .B(n1667), .Z(n1669) );
  XOR U1579 ( .A(n1681), .B(n1682), .Z(n1667) );
  AND U1580 ( .A(n352), .B(n1683), .Z(n1682) );
  IV U1581 ( .A(n1678), .Z(n1680) );
  XOR U1582 ( .A(n1684), .B(n1685), .Z(n1678) );
  AND U1583 ( .A(n336), .B(n1677), .Z(n1685) );
  XNOR U1584 ( .A(n1675), .B(n1684), .Z(n1677) );
  XNOR U1585 ( .A(n1686), .B(n1687), .Z(n1675) );
  AND U1586 ( .A(n340), .B(n1688), .Z(n1687) );
  XOR U1587 ( .A(p_input[383]), .B(n1686), .Z(n1688) );
  XNOR U1588 ( .A(n1689), .B(n1690), .Z(n1686) );
  AND U1589 ( .A(n344), .B(n1691), .Z(n1690) );
  XOR U1590 ( .A(n1692), .B(n1693), .Z(n1684) );
  AND U1591 ( .A(n348), .B(n1683), .Z(n1693) );
  XNOR U1592 ( .A(n1694), .B(n1681), .Z(n1683) );
  XOR U1593 ( .A(n1695), .B(n1696), .Z(n1681) );
  AND U1594 ( .A(n370), .B(n1697), .Z(n1696) );
  IV U1595 ( .A(n1692), .Z(n1694) );
  XOR U1596 ( .A(n1698), .B(n1699), .Z(n1692) );
  AND U1597 ( .A(n355), .B(n1691), .Z(n1699) );
  XNOR U1598 ( .A(n1689), .B(n1698), .Z(n1691) );
  XNOR U1599 ( .A(n1700), .B(n1701), .Z(n1689) );
  AND U1600 ( .A(n359), .B(n1702), .Z(n1701) );
  XOR U1601 ( .A(p_input[415]), .B(n1700), .Z(n1702) );
  XOR U1602 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][31] ), .B(n1703), 
        .Z(n1700) );
  AND U1603 ( .A(n362), .B(n1704), .Z(n1703) );
  XOR U1604 ( .A(n1705), .B(n1706), .Z(n1698) );
  AND U1605 ( .A(n366), .B(n1697), .Z(n1706) );
  XNOR U1606 ( .A(n1707), .B(n1695), .Z(n1697) );
  XOR U1607 ( .A(\knn_comb_/min_val_out[0][31] ), .B(n1708), .Z(n1695) );
  AND U1608 ( .A(n378), .B(n1709), .Z(n1708) );
  IV U1609 ( .A(n1705), .Z(n1707) );
  XOR U1610 ( .A(n1710), .B(n1711), .Z(n1705) );
  AND U1611 ( .A(n373), .B(n1704), .Z(n1711) );
  XOR U1612 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][31] ), .B(n1710), 
        .Z(n1704) );
  XOR U1613 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .B(n1712), 
        .Z(n1710) );
  AND U1614 ( .A(n375), .B(n1709), .Z(n1712) );
  XOR U1615 ( .A(n1713), .B(n1714), .Z(n1709) );
  IV U1616 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .Z(n1714) );
  IV U1617 ( .A(\knn_comb_/min_val_out[0][31] ), .Z(n1713) );
  XOR U1618 ( .A(n75), .B(n1715), .Z(o[30]) );
  AND U1619 ( .A(n122), .B(n1716), .Z(n75) );
  XOR U1620 ( .A(n76), .B(n1715), .Z(n1716) );
  XOR U1621 ( .A(n1717), .B(n1718), .Z(n1715) );
  AND U1622 ( .A(n142), .B(n1719), .Z(n1718) );
  XOR U1623 ( .A(n1720), .B(n5), .Z(n76) );
  AND U1624 ( .A(n125), .B(n1721), .Z(n5) );
  XOR U1625 ( .A(n6), .B(n1720), .Z(n1721) );
  XOR U1626 ( .A(n1722), .B(n1723), .Z(n6) );
  AND U1627 ( .A(n130), .B(n1724), .Z(n1723) );
  XOR U1628 ( .A(p_input[30]), .B(n1722), .Z(n1724) );
  XNOR U1629 ( .A(n1725), .B(n1726), .Z(n1722) );
  AND U1630 ( .A(n134), .B(n1727), .Z(n1726) );
  XOR U1631 ( .A(n1728), .B(n1729), .Z(n1720) );
  AND U1632 ( .A(n138), .B(n1719), .Z(n1729) );
  XNOR U1633 ( .A(n1730), .B(n1717), .Z(n1719) );
  XOR U1634 ( .A(n1731), .B(n1732), .Z(n1717) );
  AND U1635 ( .A(n162), .B(n1733), .Z(n1732) );
  IV U1636 ( .A(n1728), .Z(n1730) );
  XOR U1637 ( .A(n1734), .B(n1735), .Z(n1728) );
  AND U1638 ( .A(n146), .B(n1727), .Z(n1735) );
  XNOR U1639 ( .A(n1725), .B(n1734), .Z(n1727) );
  XNOR U1640 ( .A(n1736), .B(n1737), .Z(n1725) );
  AND U1641 ( .A(n150), .B(n1738), .Z(n1737) );
  XOR U1642 ( .A(p_input[62]), .B(n1736), .Z(n1738) );
  XNOR U1643 ( .A(n1739), .B(n1740), .Z(n1736) );
  AND U1644 ( .A(n154), .B(n1741), .Z(n1740) );
  XOR U1645 ( .A(n1742), .B(n1743), .Z(n1734) );
  AND U1646 ( .A(n158), .B(n1733), .Z(n1743) );
  XNOR U1647 ( .A(n1744), .B(n1731), .Z(n1733) );
  XOR U1648 ( .A(n1745), .B(n1746), .Z(n1731) );
  AND U1649 ( .A(n181), .B(n1747), .Z(n1746) );
  IV U1650 ( .A(n1742), .Z(n1744) );
  XOR U1651 ( .A(n1748), .B(n1749), .Z(n1742) );
  AND U1652 ( .A(n165), .B(n1741), .Z(n1749) );
  XNOR U1653 ( .A(n1739), .B(n1748), .Z(n1741) );
  XNOR U1654 ( .A(n1750), .B(n1751), .Z(n1739) );
  AND U1655 ( .A(n169), .B(n1752), .Z(n1751) );
  XOR U1656 ( .A(p_input[94]), .B(n1750), .Z(n1752) );
  XNOR U1657 ( .A(n1753), .B(n1754), .Z(n1750) );
  AND U1658 ( .A(n173), .B(n1755), .Z(n1754) );
  XOR U1659 ( .A(n1756), .B(n1757), .Z(n1748) );
  AND U1660 ( .A(n177), .B(n1747), .Z(n1757) );
  XNOR U1661 ( .A(n1758), .B(n1745), .Z(n1747) );
  XOR U1662 ( .A(n1759), .B(n1760), .Z(n1745) );
  AND U1663 ( .A(n200), .B(n1761), .Z(n1760) );
  IV U1664 ( .A(n1756), .Z(n1758) );
  XOR U1665 ( .A(n1762), .B(n1763), .Z(n1756) );
  AND U1666 ( .A(n184), .B(n1755), .Z(n1763) );
  XNOR U1667 ( .A(n1753), .B(n1762), .Z(n1755) );
  XNOR U1668 ( .A(n1764), .B(n1765), .Z(n1753) );
  AND U1669 ( .A(n188), .B(n1766), .Z(n1765) );
  XOR U1670 ( .A(p_input[126]), .B(n1764), .Z(n1766) );
  XNOR U1671 ( .A(n1767), .B(n1768), .Z(n1764) );
  AND U1672 ( .A(n192), .B(n1769), .Z(n1768) );
  XOR U1673 ( .A(n1770), .B(n1771), .Z(n1762) );
  AND U1674 ( .A(n196), .B(n1761), .Z(n1771) );
  XNOR U1675 ( .A(n1772), .B(n1759), .Z(n1761) );
  XOR U1676 ( .A(n1773), .B(n1774), .Z(n1759) );
  AND U1677 ( .A(n219), .B(n1775), .Z(n1774) );
  IV U1678 ( .A(n1770), .Z(n1772) );
  XOR U1679 ( .A(n1776), .B(n1777), .Z(n1770) );
  AND U1680 ( .A(n203), .B(n1769), .Z(n1777) );
  XNOR U1681 ( .A(n1767), .B(n1776), .Z(n1769) );
  XNOR U1682 ( .A(n1778), .B(n1779), .Z(n1767) );
  AND U1683 ( .A(n207), .B(n1780), .Z(n1779) );
  XOR U1684 ( .A(p_input[158]), .B(n1778), .Z(n1780) );
  XNOR U1685 ( .A(n1781), .B(n1782), .Z(n1778) );
  AND U1686 ( .A(n211), .B(n1783), .Z(n1782) );
  XOR U1687 ( .A(n1784), .B(n1785), .Z(n1776) );
  AND U1688 ( .A(n215), .B(n1775), .Z(n1785) );
  XNOR U1689 ( .A(n1786), .B(n1773), .Z(n1775) );
  XOR U1690 ( .A(n1787), .B(n1788), .Z(n1773) );
  AND U1691 ( .A(n238), .B(n1789), .Z(n1788) );
  IV U1692 ( .A(n1784), .Z(n1786) );
  XOR U1693 ( .A(n1790), .B(n1791), .Z(n1784) );
  AND U1694 ( .A(n222), .B(n1783), .Z(n1791) );
  XNOR U1695 ( .A(n1781), .B(n1790), .Z(n1783) );
  XNOR U1696 ( .A(n1792), .B(n1793), .Z(n1781) );
  AND U1697 ( .A(n226), .B(n1794), .Z(n1793) );
  XOR U1698 ( .A(p_input[190]), .B(n1792), .Z(n1794) );
  XNOR U1699 ( .A(n1795), .B(n1796), .Z(n1792) );
  AND U1700 ( .A(n230), .B(n1797), .Z(n1796) );
  XOR U1701 ( .A(n1798), .B(n1799), .Z(n1790) );
  AND U1702 ( .A(n234), .B(n1789), .Z(n1799) );
  XNOR U1703 ( .A(n1800), .B(n1787), .Z(n1789) );
  XOR U1704 ( .A(n1801), .B(n1802), .Z(n1787) );
  AND U1705 ( .A(n257), .B(n1803), .Z(n1802) );
  IV U1706 ( .A(n1798), .Z(n1800) );
  XOR U1707 ( .A(n1804), .B(n1805), .Z(n1798) );
  AND U1708 ( .A(n241), .B(n1797), .Z(n1805) );
  XNOR U1709 ( .A(n1795), .B(n1804), .Z(n1797) );
  XNOR U1710 ( .A(n1806), .B(n1807), .Z(n1795) );
  AND U1711 ( .A(n245), .B(n1808), .Z(n1807) );
  XOR U1712 ( .A(p_input[222]), .B(n1806), .Z(n1808) );
  XNOR U1713 ( .A(n1809), .B(n1810), .Z(n1806) );
  AND U1714 ( .A(n249), .B(n1811), .Z(n1810) );
  XOR U1715 ( .A(n1812), .B(n1813), .Z(n1804) );
  AND U1716 ( .A(n253), .B(n1803), .Z(n1813) );
  XNOR U1717 ( .A(n1814), .B(n1801), .Z(n1803) );
  XOR U1718 ( .A(n1815), .B(n1816), .Z(n1801) );
  AND U1719 ( .A(n276), .B(n1817), .Z(n1816) );
  IV U1720 ( .A(n1812), .Z(n1814) );
  XOR U1721 ( .A(n1818), .B(n1819), .Z(n1812) );
  AND U1722 ( .A(n260), .B(n1811), .Z(n1819) );
  XNOR U1723 ( .A(n1809), .B(n1818), .Z(n1811) );
  XNOR U1724 ( .A(n1820), .B(n1821), .Z(n1809) );
  AND U1725 ( .A(n264), .B(n1822), .Z(n1821) );
  XOR U1726 ( .A(p_input[254]), .B(n1820), .Z(n1822) );
  XNOR U1727 ( .A(n1823), .B(n1824), .Z(n1820) );
  AND U1728 ( .A(n268), .B(n1825), .Z(n1824) );
  XOR U1729 ( .A(n1826), .B(n1827), .Z(n1818) );
  AND U1730 ( .A(n272), .B(n1817), .Z(n1827) );
  XNOR U1731 ( .A(n1828), .B(n1815), .Z(n1817) );
  XOR U1732 ( .A(n1829), .B(n1830), .Z(n1815) );
  AND U1733 ( .A(n295), .B(n1831), .Z(n1830) );
  IV U1734 ( .A(n1826), .Z(n1828) );
  XOR U1735 ( .A(n1832), .B(n1833), .Z(n1826) );
  AND U1736 ( .A(n279), .B(n1825), .Z(n1833) );
  XNOR U1737 ( .A(n1823), .B(n1832), .Z(n1825) );
  XNOR U1738 ( .A(n1834), .B(n1835), .Z(n1823) );
  AND U1739 ( .A(n283), .B(n1836), .Z(n1835) );
  XOR U1740 ( .A(p_input[286]), .B(n1834), .Z(n1836) );
  XNOR U1741 ( .A(n1837), .B(n1838), .Z(n1834) );
  AND U1742 ( .A(n287), .B(n1839), .Z(n1838) );
  XOR U1743 ( .A(n1840), .B(n1841), .Z(n1832) );
  AND U1744 ( .A(n291), .B(n1831), .Z(n1841) );
  XNOR U1745 ( .A(n1842), .B(n1829), .Z(n1831) );
  XOR U1746 ( .A(n1843), .B(n1844), .Z(n1829) );
  AND U1747 ( .A(n314), .B(n1845), .Z(n1844) );
  IV U1748 ( .A(n1840), .Z(n1842) );
  XOR U1749 ( .A(n1846), .B(n1847), .Z(n1840) );
  AND U1750 ( .A(n298), .B(n1839), .Z(n1847) );
  XNOR U1751 ( .A(n1837), .B(n1846), .Z(n1839) );
  XNOR U1752 ( .A(n1848), .B(n1849), .Z(n1837) );
  AND U1753 ( .A(n302), .B(n1850), .Z(n1849) );
  XOR U1754 ( .A(p_input[318]), .B(n1848), .Z(n1850) );
  XNOR U1755 ( .A(n1851), .B(n1852), .Z(n1848) );
  AND U1756 ( .A(n306), .B(n1853), .Z(n1852) );
  XOR U1757 ( .A(n1854), .B(n1855), .Z(n1846) );
  AND U1758 ( .A(n310), .B(n1845), .Z(n1855) );
  XNOR U1759 ( .A(n1856), .B(n1843), .Z(n1845) );
  XOR U1760 ( .A(n1857), .B(n1858), .Z(n1843) );
  AND U1761 ( .A(n333), .B(n1859), .Z(n1858) );
  IV U1762 ( .A(n1854), .Z(n1856) );
  XOR U1763 ( .A(n1860), .B(n1861), .Z(n1854) );
  AND U1764 ( .A(n317), .B(n1853), .Z(n1861) );
  XNOR U1765 ( .A(n1851), .B(n1860), .Z(n1853) );
  XNOR U1766 ( .A(n1862), .B(n1863), .Z(n1851) );
  AND U1767 ( .A(n321), .B(n1864), .Z(n1863) );
  XOR U1768 ( .A(p_input[350]), .B(n1862), .Z(n1864) );
  XNOR U1769 ( .A(n1865), .B(n1866), .Z(n1862) );
  AND U1770 ( .A(n325), .B(n1867), .Z(n1866) );
  XOR U1771 ( .A(n1868), .B(n1869), .Z(n1860) );
  AND U1772 ( .A(n329), .B(n1859), .Z(n1869) );
  XNOR U1773 ( .A(n1870), .B(n1857), .Z(n1859) );
  XOR U1774 ( .A(n1871), .B(n1872), .Z(n1857) );
  AND U1775 ( .A(n352), .B(n1873), .Z(n1872) );
  IV U1776 ( .A(n1868), .Z(n1870) );
  XOR U1777 ( .A(n1874), .B(n1875), .Z(n1868) );
  AND U1778 ( .A(n336), .B(n1867), .Z(n1875) );
  XNOR U1779 ( .A(n1865), .B(n1874), .Z(n1867) );
  XNOR U1780 ( .A(n1876), .B(n1877), .Z(n1865) );
  AND U1781 ( .A(n340), .B(n1878), .Z(n1877) );
  XOR U1782 ( .A(p_input[382]), .B(n1876), .Z(n1878) );
  XNOR U1783 ( .A(n1879), .B(n1880), .Z(n1876) );
  AND U1784 ( .A(n344), .B(n1881), .Z(n1880) );
  XOR U1785 ( .A(n1882), .B(n1883), .Z(n1874) );
  AND U1786 ( .A(n348), .B(n1873), .Z(n1883) );
  XNOR U1787 ( .A(n1884), .B(n1871), .Z(n1873) );
  XOR U1788 ( .A(n1885), .B(n1886), .Z(n1871) );
  AND U1789 ( .A(n370), .B(n1887), .Z(n1886) );
  IV U1790 ( .A(n1882), .Z(n1884) );
  XOR U1791 ( .A(n1888), .B(n1889), .Z(n1882) );
  AND U1792 ( .A(n355), .B(n1881), .Z(n1889) );
  XNOR U1793 ( .A(n1879), .B(n1888), .Z(n1881) );
  XNOR U1794 ( .A(n1890), .B(n1891), .Z(n1879) );
  AND U1795 ( .A(n359), .B(n1892), .Z(n1891) );
  XOR U1796 ( .A(p_input[414]), .B(n1890), .Z(n1892) );
  XOR U1797 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][30] ), .B(n1893), 
        .Z(n1890) );
  AND U1798 ( .A(n362), .B(n1894), .Z(n1893) );
  XOR U1799 ( .A(n1895), .B(n1896), .Z(n1888) );
  AND U1800 ( .A(n366), .B(n1887), .Z(n1896) );
  XNOR U1801 ( .A(n1897), .B(n1885), .Z(n1887) );
  XOR U1802 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n1898), .Z(n1885) );
  AND U1803 ( .A(n378), .B(n1899), .Z(n1898) );
  IV U1804 ( .A(n1895), .Z(n1897) );
  XOR U1805 ( .A(n1900), .B(n1901), .Z(n1895) );
  AND U1806 ( .A(n373), .B(n1894), .Z(n1901) );
  XOR U1807 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][30] ), .B(n1900), 
        .Z(n1894) );
  XOR U1808 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .B(n1902), 
        .Z(n1900) );
  AND U1809 ( .A(n375), .B(n1899), .Z(n1902) );
  XOR U1810 ( .A(n1903), .B(n1904), .Z(n1899) );
  IV U1811 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .Z(n1904) );
  IV U1812 ( .A(\knn_comb_/min_val_out[0][30] ), .Z(n1903) );
  XOR U1813 ( .A(n1519), .B(n1905), .Z(o[2]) );
  AND U1814 ( .A(n122), .B(n1906), .Z(n1519) );
  XOR U1815 ( .A(n1520), .B(n1905), .Z(n1906) );
  XOR U1816 ( .A(n1907), .B(n1908), .Z(n1905) );
  AND U1817 ( .A(n142), .B(n1909), .Z(n1908) );
  XOR U1818 ( .A(n1910), .B(n67), .Z(n1520) );
  AND U1819 ( .A(n125), .B(n1911), .Z(n67) );
  XOR U1820 ( .A(n68), .B(n1910), .Z(n1911) );
  XOR U1821 ( .A(n1912), .B(n1913), .Z(n68) );
  AND U1822 ( .A(n130), .B(n1914), .Z(n1913) );
  XOR U1823 ( .A(p_input[2]), .B(n1912), .Z(n1914) );
  XNOR U1824 ( .A(n1915), .B(n1916), .Z(n1912) );
  AND U1825 ( .A(n134), .B(n1917), .Z(n1916) );
  XOR U1826 ( .A(n1918), .B(n1919), .Z(n1910) );
  AND U1827 ( .A(n138), .B(n1909), .Z(n1919) );
  XNOR U1828 ( .A(n1920), .B(n1907), .Z(n1909) );
  XOR U1829 ( .A(n1921), .B(n1922), .Z(n1907) );
  AND U1830 ( .A(n162), .B(n1923), .Z(n1922) );
  IV U1831 ( .A(n1918), .Z(n1920) );
  XOR U1832 ( .A(n1924), .B(n1925), .Z(n1918) );
  AND U1833 ( .A(n146), .B(n1917), .Z(n1925) );
  XNOR U1834 ( .A(n1915), .B(n1924), .Z(n1917) );
  XNOR U1835 ( .A(n1926), .B(n1927), .Z(n1915) );
  AND U1836 ( .A(n150), .B(n1928), .Z(n1927) );
  XOR U1837 ( .A(p_input[34]), .B(n1926), .Z(n1928) );
  XNOR U1838 ( .A(n1929), .B(n1930), .Z(n1926) );
  AND U1839 ( .A(n154), .B(n1931), .Z(n1930) );
  XOR U1840 ( .A(n1932), .B(n1933), .Z(n1924) );
  AND U1841 ( .A(n158), .B(n1923), .Z(n1933) );
  XNOR U1842 ( .A(n1934), .B(n1921), .Z(n1923) );
  XOR U1843 ( .A(n1935), .B(n1936), .Z(n1921) );
  AND U1844 ( .A(n181), .B(n1937), .Z(n1936) );
  IV U1845 ( .A(n1932), .Z(n1934) );
  XOR U1846 ( .A(n1938), .B(n1939), .Z(n1932) );
  AND U1847 ( .A(n165), .B(n1931), .Z(n1939) );
  XNOR U1848 ( .A(n1929), .B(n1938), .Z(n1931) );
  XNOR U1849 ( .A(n1940), .B(n1941), .Z(n1929) );
  AND U1850 ( .A(n169), .B(n1942), .Z(n1941) );
  XOR U1851 ( .A(p_input[66]), .B(n1940), .Z(n1942) );
  XNOR U1852 ( .A(n1943), .B(n1944), .Z(n1940) );
  AND U1853 ( .A(n173), .B(n1945), .Z(n1944) );
  XOR U1854 ( .A(n1946), .B(n1947), .Z(n1938) );
  AND U1855 ( .A(n177), .B(n1937), .Z(n1947) );
  XNOR U1856 ( .A(n1948), .B(n1935), .Z(n1937) );
  XOR U1857 ( .A(n1949), .B(n1950), .Z(n1935) );
  AND U1858 ( .A(n200), .B(n1951), .Z(n1950) );
  IV U1859 ( .A(n1946), .Z(n1948) );
  XOR U1860 ( .A(n1952), .B(n1953), .Z(n1946) );
  AND U1861 ( .A(n184), .B(n1945), .Z(n1953) );
  XNOR U1862 ( .A(n1943), .B(n1952), .Z(n1945) );
  XNOR U1863 ( .A(n1954), .B(n1955), .Z(n1943) );
  AND U1864 ( .A(n188), .B(n1956), .Z(n1955) );
  XOR U1865 ( .A(p_input[98]), .B(n1954), .Z(n1956) );
  XNOR U1866 ( .A(n1957), .B(n1958), .Z(n1954) );
  AND U1867 ( .A(n192), .B(n1959), .Z(n1958) );
  XOR U1868 ( .A(n1960), .B(n1961), .Z(n1952) );
  AND U1869 ( .A(n196), .B(n1951), .Z(n1961) );
  XNOR U1870 ( .A(n1962), .B(n1949), .Z(n1951) );
  XOR U1871 ( .A(n1963), .B(n1964), .Z(n1949) );
  AND U1872 ( .A(n219), .B(n1965), .Z(n1964) );
  IV U1873 ( .A(n1960), .Z(n1962) );
  XOR U1874 ( .A(n1966), .B(n1967), .Z(n1960) );
  AND U1875 ( .A(n203), .B(n1959), .Z(n1967) );
  XNOR U1876 ( .A(n1957), .B(n1966), .Z(n1959) );
  XNOR U1877 ( .A(n1968), .B(n1969), .Z(n1957) );
  AND U1878 ( .A(n207), .B(n1970), .Z(n1969) );
  XOR U1879 ( .A(p_input[130]), .B(n1968), .Z(n1970) );
  XNOR U1880 ( .A(n1971), .B(n1972), .Z(n1968) );
  AND U1881 ( .A(n211), .B(n1973), .Z(n1972) );
  XOR U1882 ( .A(n1974), .B(n1975), .Z(n1966) );
  AND U1883 ( .A(n215), .B(n1965), .Z(n1975) );
  XNOR U1884 ( .A(n1976), .B(n1963), .Z(n1965) );
  XOR U1885 ( .A(n1977), .B(n1978), .Z(n1963) );
  AND U1886 ( .A(n238), .B(n1979), .Z(n1978) );
  IV U1887 ( .A(n1974), .Z(n1976) );
  XOR U1888 ( .A(n1980), .B(n1981), .Z(n1974) );
  AND U1889 ( .A(n222), .B(n1973), .Z(n1981) );
  XNOR U1890 ( .A(n1971), .B(n1980), .Z(n1973) );
  XNOR U1891 ( .A(n1982), .B(n1983), .Z(n1971) );
  AND U1892 ( .A(n226), .B(n1984), .Z(n1983) );
  XOR U1893 ( .A(p_input[162]), .B(n1982), .Z(n1984) );
  XNOR U1894 ( .A(n1985), .B(n1986), .Z(n1982) );
  AND U1895 ( .A(n230), .B(n1987), .Z(n1986) );
  XOR U1896 ( .A(n1988), .B(n1989), .Z(n1980) );
  AND U1897 ( .A(n234), .B(n1979), .Z(n1989) );
  XNOR U1898 ( .A(n1990), .B(n1977), .Z(n1979) );
  XOR U1899 ( .A(n1991), .B(n1992), .Z(n1977) );
  AND U1900 ( .A(n257), .B(n1993), .Z(n1992) );
  IV U1901 ( .A(n1988), .Z(n1990) );
  XOR U1902 ( .A(n1994), .B(n1995), .Z(n1988) );
  AND U1903 ( .A(n241), .B(n1987), .Z(n1995) );
  XNOR U1904 ( .A(n1985), .B(n1994), .Z(n1987) );
  XNOR U1905 ( .A(n1996), .B(n1997), .Z(n1985) );
  AND U1906 ( .A(n245), .B(n1998), .Z(n1997) );
  XOR U1907 ( .A(p_input[194]), .B(n1996), .Z(n1998) );
  XNOR U1908 ( .A(n1999), .B(n2000), .Z(n1996) );
  AND U1909 ( .A(n249), .B(n2001), .Z(n2000) );
  XOR U1910 ( .A(n2002), .B(n2003), .Z(n1994) );
  AND U1911 ( .A(n253), .B(n1993), .Z(n2003) );
  XNOR U1912 ( .A(n2004), .B(n1991), .Z(n1993) );
  XOR U1913 ( .A(n2005), .B(n2006), .Z(n1991) );
  AND U1914 ( .A(n276), .B(n2007), .Z(n2006) );
  IV U1915 ( .A(n2002), .Z(n2004) );
  XOR U1916 ( .A(n2008), .B(n2009), .Z(n2002) );
  AND U1917 ( .A(n260), .B(n2001), .Z(n2009) );
  XNOR U1918 ( .A(n1999), .B(n2008), .Z(n2001) );
  XNOR U1919 ( .A(n2010), .B(n2011), .Z(n1999) );
  AND U1920 ( .A(n264), .B(n2012), .Z(n2011) );
  XOR U1921 ( .A(p_input[226]), .B(n2010), .Z(n2012) );
  XNOR U1922 ( .A(n2013), .B(n2014), .Z(n2010) );
  AND U1923 ( .A(n268), .B(n2015), .Z(n2014) );
  XOR U1924 ( .A(n2016), .B(n2017), .Z(n2008) );
  AND U1925 ( .A(n272), .B(n2007), .Z(n2017) );
  XNOR U1926 ( .A(n2018), .B(n2005), .Z(n2007) );
  XOR U1927 ( .A(n2019), .B(n2020), .Z(n2005) );
  AND U1928 ( .A(n295), .B(n2021), .Z(n2020) );
  IV U1929 ( .A(n2016), .Z(n2018) );
  XOR U1930 ( .A(n2022), .B(n2023), .Z(n2016) );
  AND U1931 ( .A(n279), .B(n2015), .Z(n2023) );
  XNOR U1932 ( .A(n2013), .B(n2022), .Z(n2015) );
  XNOR U1933 ( .A(n2024), .B(n2025), .Z(n2013) );
  AND U1934 ( .A(n283), .B(n2026), .Z(n2025) );
  XOR U1935 ( .A(p_input[258]), .B(n2024), .Z(n2026) );
  XNOR U1936 ( .A(n2027), .B(n2028), .Z(n2024) );
  AND U1937 ( .A(n287), .B(n2029), .Z(n2028) );
  XOR U1938 ( .A(n2030), .B(n2031), .Z(n2022) );
  AND U1939 ( .A(n291), .B(n2021), .Z(n2031) );
  XNOR U1940 ( .A(n2032), .B(n2019), .Z(n2021) );
  XOR U1941 ( .A(n2033), .B(n2034), .Z(n2019) );
  AND U1942 ( .A(n314), .B(n2035), .Z(n2034) );
  IV U1943 ( .A(n2030), .Z(n2032) );
  XOR U1944 ( .A(n2036), .B(n2037), .Z(n2030) );
  AND U1945 ( .A(n298), .B(n2029), .Z(n2037) );
  XNOR U1946 ( .A(n2027), .B(n2036), .Z(n2029) );
  XNOR U1947 ( .A(n2038), .B(n2039), .Z(n2027) );
  AND U1948 ( .A(n302), .B(n2040), .Z(n2039) );
  XOR U1949 ( .A(p_input[290]), .B(n2038), .Z(n2040) );
  XNOR U1950 ( .A(n2041), .B(n2042), .Z(n2038) );
  AND U1951 ( .A(n306), .B(n2043), .Z(n2042) );
  XOR U1952 ( .A(n2044), .B(n2045), .Z(n2036) );
  AND U1953 ( .A(n310), .B(n2035), .Z(n2045) );
  XNOR U1954 ( .A(n2046), .B(n2033), .Z(n2035) );
  XOR U1955 ( .A(n2047), .B(n2048), .Z(n2033) );
  AND U1956 ( .A(n333), .B(n2049), .Z(n2048) );
  IV U1957 ( .A(n2044), .Z(n2046) );
  XOR U1958 ( .A(n2050), .B(n2051), .Z(n2044) );
  AND U1959 ( .A(n317), .B(n2043), .Z(n2051) );
  XNOR U1960 ( .A(n2041), .B(n2050), .Z(n2043) );
  XNOR U1961 ( .A(n2052), .B(n2053), .Z(n2041) );
  AND U1962 ( .A(n321), .B(n2054), .Z(n2053) );
  XOR U1963 ( .A(p_input[322]), .B(n2052), .Z(n2054) );
  XNOR U1964 ( .A(n2055), .B(n2056), .Z(n2052) );
  AND U1965 ( .A(n325), .B(n2057), .Z(n2056) );
  XOR U1966 ( .A(n2058), .B(n2059), .Z(n2050) );
  AND U1967 ( .A(n329), .B(n2049), .Z(n2059) );
  XNOR U1968 ( .A(n2060), .B(n2047), .Z(n2049) );
  XOR U1969 ( .A(n2061), .B(n2062), .Z(n2047) );
  AND U1970 ( .A(n352), .B(n2063), .Z(n2062) );
  IV U1971 ( .A(n2058), .Z(n2060) );
  XOR U1972 ( .A(n2064), .B(n2065), .Z(n2058) );
  AND U1973 ( .A(n336), .B(n2057), .Z(n2065) );
  XNOR U1974 ( .A(n2055), .B(n2064), .Z(n2057) );
  XNOR U1975 ( .A(n2066), .B(n2067), .Z(n2055) );
  AND U1976 ( .A(n340), .B(n2068), .Z(n2067) );
  XOR U1977 ( .A(p_input[354]), .B(n2066), .Z(n2068) );
  XNOR U1978 ( .A(n2069), .B(n2070), .Z(n2066) );
  AND U1979 ( .A(n344), .B(n2071), .Z(n2070) );
  XOR U1980 ( .A(n2072), .B(n2073), .Z(n2064) );
  AND U1981 ( .A(n348), .B(n2063), .Z(n2073) );
  XNOR U1982 ( .A(n2074), .B(n2061), .Z(n2063) );
  XOR U1983 ( .A(n2075), .B(n2076), .Z(n2061) );
  AND U1984 ( .A(n370), .B(n2077), .Z(n2076) );
  IV U1985 ( .A(n2072), .Z(n2074) );
  XOR U1986 ( .A(n2078), .B(n2079), .Z(n2072) );
  AND U1987 ( .A(n355), .B(n2071), .Z(n2079) );
  XNOR U1988 ( .A(n2069), .B(n2078), .Z(n2071) );
  XNOR U1989 ( .A(n2080), .B(n2081), .Z(n2069) );
  AND U1990 ( .A(n359), .B(n2082), .Z(n2081) );
  XOR U1991 ( .A(p_input[386]), .B(n2080), .Z(n2082) );
  XOR U1992 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n2083), 
        .Z(n2080) );
  AND U1993 ( .A(n362), .B(n2084), .Z(n2083) );
  XOR U1994 ( .A(n2085), .B(n2086), .Z(n2078) );
  AND U1995 ( .A(n366), .B(n2077), .Z(n2086) );
  XNOR U1996 ( .A(n2087), .B(n2075), .Z(n2077) );
  XOR U1997 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n2088), .Z(n2075) );
  AND U1998 ( .A(n378), .B(n2089), .Z(n2088) );
  IV U1999 ( .A(n2085), .Z(n2087) );
  XOR U2000 ( .A(n2090), .B(n2091), .Z(n2085) );
  AND U2001 ( .A(n373), .B(n2084), .Z(n2091) );
  XOR U2002 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n2090), 
        .Z(n2084) );
  XOR U2003 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .B(n2092), 
        .Z(n2090) );
  AND U2004 ( .A(n375), .B(n2089), .Z(n2092) );
  XOR U2005 ( .A(\knn_comb_/min_val_out[0][2] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .Z(n2089) );
  XOR U2006 ( .A(n77), .B(n2093), .Z(o[29]) );
  AND U2007 ( .A(n122), .B(n2094), .Z(n77) );
  XOR U2008 ( .A(n78), .B(n2093), .Z(n2094) );
  XOR U2009 ( .A(n2095), .B(n2096), .Z(n2093) );
  AND U2010 ( .A(n142), .B(n2097), .Z(n2096) );
  XOR U2011 ( .A(n2098), .B(n7), .Z(n78) );
  AND U2012 ( .A(n125), .B(n2099), .Z(n7) );
  XOR U2013 ( .A(n8), .B(n2098), .Z(n2099) );
  XOR U2014 ( .A(n2100), .B(n2101), .Z(n8) );
  AND U2015 ( .A(n130), .B(n2102), .Z(n2101) );
  XOR U2016 ( .A(p_input[29]), .B(n2100), .Z(n2102) );
  XNOR U2017 ( .A(n2103), .B(n2104), .Z(n2100) );
  AND U2018 ( .A(n134), .B(n2105), .Z(n2104) );
  XOR U2019 ( .A(n2106), .B(n2107), .Z(n2098) );
  AND U2020 ( .A(n138), .B(n2097), .Z(n2107) );
  XNOR U2021 ( .A(n2108), .B(n2095), .Z(n2097) );
  XOR U2022 ( .A(n2109), .B(n2110), .Z(n2095) );
  AND U2023 ( .A(n162), .B(n2111), .Z(n2110) );
  IV U2024 ( .A(n2106), .Z(n2108) );
  XOR U2025 ( .A(n2112), .B(n2113), .Z(n2106) );
  AND U2026 ( .A(n146), .B(n2105), .Z(n2113) );
  XNOR U2027 ( .A(n2103), .B(n2112), .Z(n2105) );
  XNOR U2028 ( .A(n2114), .B(n2115), .Z(n2103) );
  AND U2029 ( .A(n150), .B(n2116), .Z(n2115) );
  XOR U2030 ( .A(p_input[61]), .B(n2114), .Z(n2116) );
  XNOR U2031 ( .A(n2117), .B(n2118), .Z(n2114) );
  AND U2032 ( .A(n154), .B(n2119), .Z(n2118) );
  XOR U2033 ( .A(n2120), .B(n2121), .Z(n2112) );
  AND U2034 ( .A(n158), .B(n2111), .Z(n2121) );
  XNOR U2035 ( .A(n2122), .B(n2109), .Z(n2111) );
  XOR U2036 ( .A(n2123), .B(n2124), .Z(n2109) );
  AND U2037 ( .A(n181), .B(n2125), .Z(n2124) );
  IV U2038 ( .A(n2120), .Z(n2122) );
  XOR U2039 ( .A(n2126), .B(n2127), .Z(n2120) );
  AND U2040 ( .A(n165), .B(n2119), .Z(n2127) );
  XNOR U2041 ( .A(n2117), .B(n2126), .Z(n2119) );
  XNOR U2042 ( .A(n2128), .B(n2129), .Z(n2117) );
  AND U2043 ( .A(n169), .B(n2130), .Z(n2129) );
  XOR U2044 ( .A(p_input[93]), .B(n2128), .Z(n2130) );
  XNOR U2045 ( .A(n2131), .B(n2132), .Z(n2128) );
  AND U2046 ( .A(n173), .B(n2133), .Z(n2132) );
  XOR U2047 ( .A(n2134), .B(n2135), .Z(n2126) );
  AND U2048 ( .A(n177), .B(n2125), .Z(n2135) );
  XNOR U2049 ( .A(n2136), .B(n2123), .Z(n2125) );
  XOR U2050 ( .A(n2137), .B(n2138), .Z(n2123) );
  AND U2051 ( .A(n200), .B(n2139), .Z(n2138) );
  IV U2052 ( .A(n2134), .Z(n2136) );
  XOR U2053 ( .A(n2140), .B(n2141), .Z(n2134) );
  AND U2054 ( .A(n184), .B(n2133), .Z(n2141) );
  XNOR U2055 ( .A(n2131), .B(n2140), .Z(n2133) );
  XNOR U2056 ( .A(n2142), .B(n2143), .Z(n2131) );
  AND U2057 ( .A(n188), .B(n2144), .Z(n2143) );
  XOR U2058 ( .A(p_input[125]), .B(n2142), .Z(n2144) );
  XNOR U2059 ( .A(n2145), .B(n2146), .Z(n2142) );
  AND U2060 ( .A(n192), .B(n2147), .Z(n2146) );
  XOR U2061 ( .A(n2148), .B(n2149), .Z(n2140) );
  AND U2062 ( .A(n196), .B(n2139), .Z(n2149) );
  XNOR U2063 ( .A(n2150), .B(n2137), .Z(n2139) );
  XOR U2064 ( .A(n2151), .B(n2152), .Z(n2137) );
  AND U2065 ( .A(n219), .B(n2153), .Z(n2152) );
  IV U2066 ( .A(n2148), .Z(n2150) );
  XOR U2067 ( .A(n2154), .B(n2155), .Z(n2148) );
  AND U2068 ( .A(n203), .B(n2147), .Z(n2155) );
  XNOR U2069 ( .A(n2145), .B(n2154), .Z(n2147) );
  XNOR U2070 ( .A(n2156), .B(n2157), .Z(n2145) );
  AND U2071 ( .A(n207), .B(n2158), .Z(n2157) );
  XOR U2072 ( .A(p_input[157]), .B(n2156), .Z(n2158) );
  XNOR U2073 ( .A(n2159), .B(n2160), .Z(n2156) );
  AND U2074 ( .A(n211), .B(n2161), .Z(n2160) );
  XOR U2075 ( .A(n2162), .B(n2163), .Z(n2154) );
  AND U2076 ( .A(n215), .B(n2153), .Z(n2163) );
  XNOR U2077 ( .A(n2164), .B(n2151), .Z(n2153) );
  XOR U2078 ( .A(n2165), .B(n2166), .Z(n2151) );
  AND U2079 ( .A(n238), .B(n2167), .Z(n2166) );
  IV U2080 ( .A(n2162), .Z(n2164) );
  XOR U2081 ( .A(n2168), .B(n2169), .Z(n2162) );
  AND U2082 ( .A(n222), .B(n2161), .Z(n2169) );
  XNOR U2083 ( .A(n2159), .B(n2168), .Z(n2161) );
  XNOR U2084 ( .A(n2170), .B(n2171), .Z(n2159) );
  AND U2085 ( .A(n226), .B(n2172), .Z(n2171) );
  XOR U2086 ( .A(p_input[189]), .B(n2170), .Z(n2172) );
  XNOR U2087 ( .A(n2173), .B(n2174), .Z(n2170) );
  AND U2088 ( .A(n230), .B(n2175), .Z(n2174) );
  XOR U2089 ( .A(n2176), .B(n2177), .Z(n2168) );
  AND U2090 ( .A(n234), .B(n2167), .Z(n2177) );
  XNOR U2091 ( .A(n2178), .B(n2165), .Z(n2167) );
  XOR U2092 ( .A(n2179), .B(n2180), .Z(n2165) );
  AND U2093 ( .A(n257), .B(n2181), .Z(n2180) );
  IV U2094 ( .A(n2176), .Z(n2178) );
  XOR U2095 ( .A(n2182), .B(n2183), .Z(n2176) );
  AND U2096 ( .A(n241), .B(n2175), .Z(n2183) );
  XNOR U2097 ( .A(n2173), .B(n2182), .Z(n2175) );
  XNOR U2098 ( .A(n2184), .B(n2185), .Z(n2173) );
  AND U2099 ( .A(n245), .B(n2186), .Z(n2185) );
  XOR U2100 ( .A(p_input[221]), .B(n2184), .Z(n2186) );
  XNOR U2101 ( .A(n2187), .B(n2188), .Z(n2184) );
  AND U2102 ( .A(n249), .B(n2189), .Z(n2188) );
  XOR U2103 ( .A(n2190), .B(n2191), .Z(n2182) );
  AND U2104 ( .A(n253), .B(n2181), .Z(n2191) );
  XNOR U2105 ( .A(n2192), .B(n2179), .Z(n2181) );
  XOR U2106 ( .A(n2193), .B(n2194), .Z(n2179) );
  AND U2107 ( .A(n276), .B(n2195), .Z(n2194) );
  IV U2108 ( .A(n2190), .Z(n2192) );
  XOR U2109 ( .A(n2196), .B(n2197), .Z(n2190) );
  AND U2110 ( .A(n260), .B(n2189), .Z(n2197) );
  XNOR U2111 ( .A(n2187), .B(n2196), .Z(n2189) );
  XNOR U2112 ( .A(n2198), .B(n2199), .Z(n2187) );
  AND U2113 ( .A(n264), .B(n2200), .Z(n2199) );
  XOR U2114 ( .A(p_input[253]), .B(n2198), .Z(n2200) );
  XNOR U2115 ( .A(n2201), .B(n2202), .Z(n2198) );
  AND U2116 ( .A(n268), .B(n2203), .Z(n2202) );
  XOR U2117 ( .A(n2204), .B(n2205), .Z(n2196) );
  AND U2118 ( .A(n272), .B(n2195), .Z(n2205) );
  XNOR U2119 ( .A(n2206), .B(n2193), .Z(n2195) );
  XOR U2120 ( .A(n2207), .B(n2208), .Z(n2193) );
  AND U2121 ( .A(n295), .B(n2209), .Z(n2208) );
  IV U2122 ( .A(n2204), .Z(n2206) );
  XOR U2123 ( .A(n2210), .B(n2211), .Z(n2204) );
  AND U2124 ( .A(n279), .B(n2203), .Z(n2211) );
  XNOR U2125 ( .A(n2201), .B(n2210), .Z(n2203) );
  XNOR U2126 ( .A(n2212), .B(n2213), .Z(n2201) );
  AND U2127 ( .A(n283), .B(n2214), .Z(n2213) );
  XOR U2128 ( .A(p_input[285]), .B(n2212), .Z(n2214) );
  XNOR U2129 ( .A(n2215), .B(n2216), .Z(n2212) );
  AND U2130 ( .A(n287), .B(n2217), .Z(n2216) );
  XOR U2131 ( .A(n2218), .B(n2219), .Z(n2210) );
  AND U2132 ( .A(n291), .B(n2209), .Z(n2219) );
  XNOR U2133 ( .A(n2220), .B(n2207), .Z(n2209) );
  XOR U2134 ( .A(n2221), .B(n2222), .Z(n2207) );
  AND U2135 ( .A(n314), .B(n2223), .Z(n2222) );
  IV U2136 ( .A(n2218), .Z(n2220) );
  XOR U2137 ( .A(n2224), .B(n2225), .Z(n2218) );
  AND U2138 ( .A(n298), .B(n2217), .Z(n2225) );
  XNOR U2139 ( .A(n2215), .B(n2224), .Z(n2217) );
  XNOR U2140 ( .A(n2226), .B(n2227), .Z(n2215) );
  AND U2141 ( .A(n302), .B(n2228), .Z(n2227) );
  XOR U2142 ( .A(p_input[317]), .B(n2226), .Z(n2228) );
  XNOR U2143 ( .A(n2229), .B(n2230), .Z(n2226) );
  AND U2144 ( .A(n306), .B(n2231), .Z(n2230) );
  XOR U2145 ( .A(n2232), .B(n2233), .Z(n2224) );
  AND U2146 ( .A(n310), .B(n2223), .Z(n2233) );
  XNOR U2147 ( .A(n2234), .B(n2221), .Z(n2223) );
  XOR U2148 ( .A(n2235), .B(n2236), .Z(n2221) );
  AND U2149 ( .A(n333), .B(n2237), .Z(n2236) );
  IV U2150 ( .A(n2232), .Z(n2234) );
  XOR U2151 ( .A(n2238), .B(n2239), .Z(n2232) );
  AND U2152 ( .A(n317), .B(n2231), .Z(n2239) );
  XNOR U2153 ( .A(n2229), .B(n2238), .Z(n2231) );
  XNOR U2154 ( .A(n2240), .B(n2241), .Z(n2229) );
  AND U2155 ( .A(n321), .B(n2242), .Z(n2241) );
  XOR U2156 ( .A(p_input[349]), .B(n2240), .Z(n2242) );
  XNOR U2157 ( .A(n2243), .B(n2244), .Z(n2240) );
  AND U2158 ( .A(n325), .B(n2245), .Z(n2244) );
  XOR U2159 ( .A(n2246), .B(n2247), .Z(n2238) );
  AND U2160 ( .A(n329), .B(n2237), .Z(n2247) );
  XNOR U2161 ( .A(n2248), .B(n2235), .Z(n2237) );
  XOR U2162 ( .A(n2249), .B(n2250), .Z(n2235) );
  AND U2163 ( .A(n352), .B(n2251), .Z(n2250) );
  IV U2164 ( .A(n2246), .Z(n2248) );
  XOR U2165 ( .A(n2252), .B(n2253), .Z(n2246) );
  AND U2166 ( .A(n336), .B(n2245), .Z(n2253) );
  XNOR U2167 ( .A(n2243), .B(n2252), .Z(n2245) );
  XNOR U2168 ( .A(n2254), .B(n2255), .Z(n2243) );
  AND U2169 ( .A(n340), .B(n2256), .Z(n2255) );
  XOR U2170 ( .A(p_input[381]), .B(n2254), .Z(n2256) );
  XNOR U2171 ( .A(n2257), .B(n2258), .Z(n2254) );
  AND U2172 ( .A(n344), .B(n2259), .Z(n2258) );
  XOR U2173 ( .A(n2260), .B(n2261), .Z(n2252) );
  AND U2174 ( .A(n348), .B(n2251), .Z(n2261) );
  XNOR U2175 ( .A(n2262), .B(n2249), .Z(n2251) );
  XOR U2176 ( .A(n2263), .B(n2264), .Z(n2249) );
  AND U2177 ( .A(n370), .B(n2265), .Z(n2264) );
  IV U2178 ( .A(n2260), .Z(n2262) );
  XOR U2179 ( .A(n2266), .B(n2267), .Z(n2260) );
  AND U2180 ( .A(n355), .B(n2259), .Z(n2267) );
  XNOR U2181 ( .A(n2257), .B(n2266), .Z(n2259) );
  XNOR U2182 ( .A(n2268), .B(n2269), .Z(n2257) );
  AND U2183 ( .A(n359), .B(n2270), .Z(n2269) );
  XOR U2184 ( .A(p_input[413]), .B(n2268), .Z(n2270) );
  XOR U2185 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][29] ), .B(n2271), 
        .Z(n2268) );
  AND U2186 ( .A(n362), .B(n2272), .Z(n2271) );
  XOR U2187 ( .A(n2273), .B(n2274), .Z(n2266) );
  AND U2188 ( .A(n366), .B(n2265), .Z(n2274) );
  XNOR U2189 ( .A(n2275), .B(n2263), .Z(n2265) );
  XOR U2190 ( .A(\knn_comb_/min_val_out[0][29] ), .B(n2276), .Z(n2263) );
  AND U2191 ( .A(n378), .B(n2277), .Z(n2276) );
  IV U2192 ( .A(n2273), .Z(n2275) );
  XOR U2193 ( .A(n2278), .B(n2279), .Z(n2273) );
  AND U2194 ( .A(n373), .B(n2272), .Z(n2279) );
  XOR U2195 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][29] ), .B(n2278), 
        .Z(n2272) );
  XOR U2196 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .B(n2280), 
        .Z(n2278) );
  AND U2197 ( .A(n375), .B(n2277), .Z(n2280) );
  XOR U2198 ( .A(\knn_comb_/min_val_out[0][29] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .Z(n2277) );
  XOR U2199 ( .A(n79), .B(n2281), .Z(o[28]) );
  AND U2200 ( .A(n122), .B(n2282), .Z(n79) );
  XOR U2201 ( .A(n80), .B(n2281), .Z(n2282) );
  XOR U2202 ( .A(n2283), .B(n2284), .Z(n2281) );
  AND U2203 ( .A(n142), .B(n2285), .Z(n2284) );
  XOR U2204 ( .A(n2286), .B(n9), .Z(n80) );
  AND U2205 ( .A(n125), .B(n2287), .Z(n9) );
  XOR U2206 ( .A(n10), .B(n2286), .Z(n2287) );
  XOR U2207 ( .A(n2288), .B(n2289), .Z(n10) );
  AND U2208 ( .A(n130), .B(n2290), .Z(n2289) );
  XOR U2209 ( .A(p_input[28]), .B(n2288), .Z(n2290) );
  XNOR U2210 ( .A(n2291), .B(n2292), .Z(n2288) );
  AND U2211 ( .A(n134), .B(n2293), .Z(n2292) );
  XOR U2212 ( .A(n2294), .B(n2295), .Z(n2286) );
  AND U2213 ( .A(n138), .B(n2285), .Z(n2295) );
  XNOR U2214 ( .A(n2296), .B(n2283), .Z(n2285) );
  XOR U2215 ( .A(n2297), .B(n2298), .Z(n2283) );
  AND U2216 ( .A(n162), .B(n2299), .Z(n2298) );
  IV U2217 ( .A(n2294), .Z(n2296) );
  XOR U2218 ( .A(n2300), .B(n2301), .Z(n2294) );
  AND U2219 ( .A(n146), .B(n2293), .Z(n2301) );
  XNOR U2220 ( .A(n2291), .B(n2300), .Z(n2293) );
  XNOR U2221 ( .A(n2302), .B(n2303), .Z(n2291) );
  AND U2222 ( .A(n150), .B(n2304), .Z(n2303) );
  XOR U2223 ( .A(p_input[60]), .B(n2302), .Z(n2304) );
  XNOR U2224 ( .A(n2305), .B(n2306), .Z(n2302) );
  AND U2225 ( .A(n154), .B(n2307), .Z(n2306) );
  XOR U2226 ( .A(n2308), .B(n2309), .Z(n2300) );
  AND U2227 ( .A(n158), .B(n2299), .Z(n2309) );
  XNOR U2228 ( .A(n2310), .B(n2297), .Z(n2299) );
  XOR U2229 ( .A(n2311), .B(n2312), .Z(n2297) );
  AND U2230 ( .A(n181), .B(n2313), .Z(n2312) );
  IV U2231 ( .A(n2308), .Z(n2310) );
  XOR U2232 ( .A(n2314), .B(n2315), .Z(n2308) );
  AND U2233 ( .A(n165), .B(n2307), .Z(n2315) );
  XNOR U2234 ( .A(n2305), .B(n2314), .Z(n2307) );
  XNOR U2235 ( .A(n2316), .B(n2317), .Z(n2305) );
  AND U2236 ( .A(n169), .B(n2318), .Z(n2317) );
  XOR U2237 ( .A(p_input[92]), .B(n2316), .Z(n2318) );
  XNOR U2238 ( .A(n2319), .B(n2320), .Z(n2316) );
  AND U2239 ( .A(n173), .B(n2321), .Z(n2320) );
  XOR U2240 ( .A(n2322), .B(n2323), .Z(n2314) );
  AND U2241 ( .A(n177), .B(n2313), .Z(n2323) );
  XNOR U2242 ( .A(n2324), .B(n2311), .Z(n2313) );
  XOR U2243 ( .A(n2325), .B(n2326), .Z(n2311) );
  AND U2244 ( .A(n200), .B(n2327), .Z(n2326) );
  IV U2245 ( .A(n2322), .Z(n2324) );
  XOR U2246 ( .A(n2328), .B(n2329), .Z(n2322) );
  AND U2247 ( .A(n184), .B(n2321), .Z(n2329) );
  XNOR U2248 ( .A(n2319), .B(n2328), .Z(n2321) );
  XNOR U2249 ( .A(n2330), .B(n2331), .Z(n2319) );
  AND U2250 ( .A(n188), .B(n2332), .Z(n2331) );
  XOR U2251 ( .A(p_input[124]), .B(n2330), .Z(n2332) );
  XNOR U2252 ( .A(n2333), .B(n2334), .Z(n2330) );
  AND U2253 ( .A(n192), .B(n2335), .Z(n2334) );
  XOR U2254 ( .A(n2336), .B(n2337), .Z(n2328) );
  AND U2255 ( .A(n196), .B(n2327), .Z(n2337) );
  XNOR U2256 ( .A(n2338), .B(n2325), .Z(n2327) );
  XOR U2257 ( .A(n2339), .B(n2340), .Z(n2325) );
  AND U2258 ( .A(n219), .B(n2341), .Z(n2340) );
  IV U2259 ( .A(n2336), .Z(n2338) );
  XOR U2260 ( .A(n2342), .B(n2343), .Z(n2336) );
  AND U2261 ( .A(n203), .B(n2335), .Z(n2343) );
  XNOR U2262 ( .A(n2333), .B(n2342), .Z(n2335) );
  XNOR U2263 ( .A(n2344), .B(n2345), .Z(n2333) );
  AND U2264 ( .A(n207), .B(n2346), .Z(n2345) );
  XOR U2265 ( .A(p_input[156]), .B(n2344), .Z(n2346) );
  XNOR U2266 ( .A(n2347), .B(n2348), .Z(n2344) );
  AND U2267 ( .A(n211), .B(n2349), .Z(n2348) );
  XOR U2268 ( .A(n2350), .B(n2351), .Z(n2342) );
  AND U2269 ( .A(n215), .B(n2341), .Z(n2351) );
  XNOR U2270 ( .A(n2352), .B(n2339), .Z(n2341) );
  XOR U2271 ( .A(n2353), .B(n2354), .Z(n2339) );
  AND U2272 ( .A(n238), .B(n2355), .Z(n2354) );
  IV U2273 ( .A(n2350), .Z(n2352) );
  XOR U2274 ( .A(n2356), .B(n2357), .Z(n2350) );
  AND U2275 ( .A(n222), .B(n2349), .Z(n2357) );
  XNOR U2276 ( .A(n2347), .B(n2356), .Z(n2349) );
  XNOR U2277 ( .A(n2358), .B(n2359), .Z(n2347) );
  AND U2278 ( .A(n226), .B(n2360), .Z(n2359) );
  XOR U2279 ( .A(p_input[188]), .B(n2358), .Z(n2360) );
  XNOR U2280 ( .A(n2361), .B(n2362), .Z(n2358) );
  AND U2281 ( .A(n230), .B(n2363), .Z(n2362) );
  XOR U2282 ( .A(n2364), .B(n2365), .Z(n2356) );
  AND U2283 ( .A(n234), .B(n2355), .Z(n2365) );
  XNOR U2284 ( .A(n2366), .B(n2353), .Z(n2355) );
  XOR U2285 ( .A(n2367), .B(n2368), .Z(n2353) );
  AND U2286 ( .A(n257), .B(n2369), .Z(n2368) );
  IV U2287 ( .A(n2364), .Z(n2366) );
  XOR U2288 ( .A(n2370), .B(n2371), .Z(n2364) );
  AND U2289 ( .A(n241), .B(n2363), .Z(n2371) );
  XNOR U2290 ( .A(n2361), .B(n2370), .Z(n2363) );
  XNOR U2291 ( .A(n2372), .B(n2373), .Z(n2361) );
  AND U2292 ( .A(n245), .B(n2374), .Z(n2373) );
  XOR U2293 ( .A(p_input[220]), .B(n2372), .Z(n2374) );
  XNOR U2294 ( .A(n2375), .B(n2376), .Z(n2372) );
  AND U2295 ( .A(n249), .B(n2377), .Z(n2376) );
  XOR U2296 ( .A(n2378), .B(n2379), .Z(n2370) );
  AND U2297 ( .A(n253), .B(n2369), .Z(n2379) );
  XNOR U2298 ( .A(n2380), .B(n2367), .Z(n2369) );
  XOR U2299 ( .A(n2381), .B(n2382), .Z(n2367) );
  AND U2300 ( .A(n276), .B(n2383), .Z(n2382) );
  IV U2301 ( .A(n2378), .Z(n2380) );
  XOR U2302 ( .A(n2384), .B(n2385), .Z(n2378) );
  AND U2303 ( .A(n260), .B(n2377), .Z(n2385) );
  XNOR U2304 ( .A(n2375), .B(n2384), .Z(n2377) );
  XNOR U2305 ( .A(n2386), .B(n2387), .Z(n2375) );
  AND U2306 ( .A(n264), .B(n2388), .Z(n2387) );
  XOR U2307 ( .A(p_input[252]), .B(n2386), .Z(n2388) );
  XNOR U2308 ( .A(n2389), .B(n2390), .Z(n2386) );
  AND U2309 ( .A(n268), .B(n2391), .Z(n2390) );
  XOR U2310 ( .A(n2392), .B(n2393), .Z(n2384) );
  AND U2311 ( .A(n272), .B(n2383), .Z(n2393) );
  XNOR U2312 ( .A(n2394), .B(n2381), .Z(n2383) );
  XOR U2313 ( .A(n2395), .B(n2396), .Z(n2381) );
  AND U2314 ( .A(n295), .B(n2397), .Z(n2396) );
  IV U2315 ( .A(n2392), .Z(n2394) );
  XOR U2316 ( .A(n2398), .B(n2399), .Z(n2392) );
  AND U2317 ( .A(n279), .B(n2391), .Z(n2399) );
  XNOR U2318 ( .A(n2389), .B(n2398), .Z(n2391) );
  XNOR U2319 ( .A(n2400), .B(n2401), .Z(n2389) );
  AND U2320 ( .A(n283), .B(n2402), .Z(n2401) );
  XOR U2321 ( .A(p_input[284]), .B(n2400), .Z(n2402) );
  XNOR U2322 ( .A(n2403), .B(n2404), .Z(n2400) );
  AND U2323 ( .A(n287), .B(n2405), .Z(n2404) );
  XOR U2324 ( .A(n2406), .B(n2407), .Z(n2398) );
  AND U2325 ( .A(n291), .B(n2397), .Z(n2407) );
  XNOR U2326 ( .A(n2408), .B(n2395), .Z(n2397) );
  XOR U2327 ( .A(n2409), .B(n2410), .Z(n2395) );
  AND U2328 ( .A(n314), .B(n2411), .Z(n2410) );
  IV U2329 ( .A(n2406), .Z(n2408) );
  XOR U2330 ( .A(n2412), .B(n2413), .Z(n2406) );
  AND U2331 ( .A(n298), .B(n2405), .Z(n2413) );
  XNOR U2332 ( .A(n2403), .B(n2412), .Z(n2405) );
  XNOR U2333 ( .A(n2414), .B(n2415), .Z(n2403) );
  AND U2334 ( .A(n302), .B(n2416), .Z(n2415) );
  XOR U2335 ( .A(p_input[316]), .B(n2414), .Z(n2416) );
  XNOR U2336 ( .A(n2417), .B(n2418), .Z(n2414) );
  AND U2337 ( .A(n306), .B(n2419), .Z(n2418) );
  XOR U2338 ( .A(n2420), .B(n2421), .Z(n2412) );
  AND U2339 ( .A(n310), .B(n2411), .Z(n2421) );
  XNOR U2340 ( .A(n2422), .B(n2409), .Z(n2411) );
  XOR U2341 ( .A(n2423), .B(n2424), .Z(n2409) );
  AND U2342 ( .A(n333), .B(n2425), .Z(n2424) );
  IV U2343 ( .A(n2420), .Z(n2422) );
  XOR U2344 ( .A(n2426), .B(n2427), .Z(n2420) );
  AND U2345 ( .A(n317), .B(n2419), .Z(n2427) );
  XNOR U2346 ( .A(n2417), .B(n2426), .Z(n2419) );
  XNOR U2347 ( .A(n2428), .B(n2429), .Z(n2417) );
  AND U2348 ( .A(n321), .B(n2430), .Z(n2429) );
  XOR U2349 ( .A(p_input[348]), .B(n2428), .Z(n2430) );
  XNOR U2350 ( .A(n2431), .B(n2432), .Z(n2428) );
  AND U2351 ( .A(n325), .B(n2433), .Z(n2432) );
  XOR U2352 ( .A(n2434), .B(n2435), .Z(n2426) );
  AND U2353 ( .A(n329), .B(n2425), .Z(n2435) );
  XNOR U2354 ( .A(n2436), .B(n2423), .Z(n2425) );
  XOR U2355 ( .A(n2437), .B(n2438), .Z(n2423) );
  AND U2356 ( .A(n352), .B(n2439), .Z(n2438) );
  IV U2357 ( .A(n2434), .Z(n2436) );
  XOR U2358 ( .A(n2440), .B(n2441), .Z(n2434) );
  AND U2359 ( .A(n336), .B(n2433), .Z(n2441) );
  XNOR U2360 ( .A(n2431), .B(n2440), .Z(n2433) );
  XNOR U2361 ( .A(n2442), .B(n2443), .Z(n2431) );
  AND U2362 ( .A(n340), .B(n2444), .Z(n2443) );
  XOR U2363 ( .A(p_input[380]), .B(n2442), .Z(n2444) );
  XNOR U2364 ( .A(n2445), .B(n2446), .Z(n2442) );
  AND U2365 ( .A(n344), .B(n2447), .Z(n2446) );
  XOR U2366 ( .A(n2448), .B(n2449), .Z(n2440) );
  AND U2367 ( .A(n348), .B(n2439), .Z(n2449) );
  XNOR U2368 ( .A(n2450), .B(n2437), .Z(n2439) );
  XOR U2369 ( .A(n2451), .B(n2452), .Z(n2437) );
  AND U2370 ( .A(n370), .B(n2453), .Z(n2452) );
  IV U2371 ( .A(n2448), .Z(n2450) );
  XOR U2372 ( .A(n2454), .B(n2455), .Z(n2448) );
  AND U2373 ( .A(n355), .B(n2447), .Z(n2455) );
  XNOR U2374 ( .A(n2445), .B(n2454), .Z(n2447) );
  XNOR U2375 ( .A(n2456), .B(n2457), .Z(n2445) );
  AND U2376 ( .A(n359), .B(n2458), .Z(n2457) );
  XOR U2377 ( .A(p_input[412]), .B(n2456), .Z(n2458) );
  XOR U2378 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][28] ), .B(n2459), 
        .Z(n2456) );
  AND U2379 ( .A(n362), .B(n2460), .Z(n2459) );
  XOR U2380 ( .A(n2461), .B(n2462), .Z(n2454) );
  AND U2381 ( .A(n366), .B(n2453), .Z(n2462) );
  XNOR U2382 ( .A(n2463), .B(n2451), .Z(n2453) );
  XOR U2383 ( .A(\knn_comb_/min_val_out[0][28] ), .B(n2464), .Z(n2451) );
  AND U2384 ( .A(n378), .B(n2465), .Z(n2464) );
  IV U2385 ( .A(n2461), .Z(n2463) );
  XOR U2386 ( .A(n2466), .B(n2467), .Z(n2461) );
  AND U2387 ( .A(n373), .B(n2460), .Z(n2467) );
  XOR U2388 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][28] ), .B(n2466), 
        .Z(n2460) );
  XOR U2389 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .B(n2468), 
        .Z(n2466) );
  AND U2390 ( .A(n375), .B(n2465), .Z(n2468) );
  XOR U2391 ( .A(\knn_comb_/min_val_out[0][28] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .Z(n2465) );
  XOR U2392 ( .A(n83), .B(n2469), .Z(o[27]) );
  AND U2393 ( .A(n122), .B(n2470), .Z(n83) );
  XOR U2394 ( .A(n84), .B(n2469), .Z(n2470) );
  XOR U2395 ( .A(n2471), .B(n2472), .Z(n2469) );
  AND U2396 ( .A(n142), .B(n2473), .Z(n2472) );
  XOR U2397 ( .A(n2474), .B(n11), .Z(n84) );
  AND U2398 ( .A(n125), .B(n2475), .Z(n11) );
  XOR U2399 ( .A(n12), .B(n2474), .Z(n2475) );
  XOR U2400 ( .A(n2476), .B(n2477), .Z(n12) );
  AND U2401 ( .A(n130), .B(n2478), .Z(n2477) );
  XOR U2402 ( .A(p_input[27]), .B(n2476), .Z(n2478) );
  XNOR U2403 ( .A(n2479), .B(n2480), .Z(n2476) );
  AND U2404 ( .A(n134), .B(n2481), .Z(n2480) );
  XOR U2405 ( .A(n2482), .B(n2483), .Z(n2474) );
  AND U2406 ( .A(n138), .B(n2473), .Z(n2483) );
  XNOR U2407 ( .A(n2484), .B(n2471), .Z(n2473) );
  XOR U2408 ( .A(n2485), .B(n2486), .Z(n2471) );
  AND U2409 ( .A(n162), .B(n2487), .Z(n2486) );
  IV U2410 ( .A(n2482), .Z(n2484) );
  XOR U2411 ( .A(n2488), .B(n2489), .Z(n2482) );
  AND U2412 ( .A(n146), .B(n2481), .Z(n2489) );
  XNOR U2413 ( .A(n2479), .B(n2488), .Z(n2481) );
  XNOR U2414 ( .A(n2490), .B(n2491), .Z(n2479) );
  AND U2415 ( .A(n150), .B(n2492), .Z(n2491) );
  XOR U2416 ( .A(p_input[59]), .B(n2490), .Z(n2492) );
  XNOR U2417 ( .A(n2493), .B(n2494), .Z(n2490) );
  AND U2418 ( .A(n154), .B(n2495), .Z(n2494) );
  XOR U2419 ( .A(n2496), .B(n2497), .Z(n2488) );
  AND U2420 ( .A(n158), .B(n2487), .Z(n2497) );
  XNOR U2421 ( .A(n2498), .B(n2485), .Z(n2487) );
  XOR U2422 ( .A(n2499), .B(n2500), .Z(n2485) );
  AND U2423 ( .A(n181), .B(n2501), .Z(n2500) );
  IV U2424 ( .A(n2496), .Z(n2498) );
  XOR U2425 ( .A(n2502), .B(n2503), .Z(n2496) );
  AND U2426 ( .A(n165), .B(n2495), .Z(n2503) );
  XNOR U2427 ( .A(n2493), .B(n2502), .Z(n2495) );
  XNOR U2428 ( .A(n2504), .B(n2505), .Z(n2493) );
  AND U2429 ( .A(n169), .B(n2506), .Z(n2505) );
  XOR U2430 ( .A(p_input[91]), .B(n2504), .Z(n2506) );
  XNOR U2431 ( .A(n2507), .B(n2508), .Z(n2504) );
  AND U2432 ( .A(n173), .B(n2509), .Z(n2508) );
  XOR U2433 ( .A(n2510), .B(n2511), .Z(n2502) );
  AND U2434 ( .A(n177), .B(n2501), .Z(n2511) );
  XNOR U2435 ( .A(n2512), .B(n2499), .Z(n2501) );
  XOR U2436 ( .A(n2513), .B(n2514), .Z(n2499) );
  AND U2437 ( .A(n200), .B(n2515), .Z(n2514) );
  IV U2438 ( .A(n2510), .Z(n2512) );
  XOR U2439 ( .A(n2516), .B(n2517), .Z(n2510) );
  AND U2440 ( .A(n184), .B(n2509), .Z(n2517) );
  XNOR U2441 ( .A(n2507), .B(n2516), .Z(n2509) );
  XNOR U2442 ( .A(n2518), .B(n2519), .Z(n2507) );
  AND U2443 ( .A(n188), .B(n2520), .Z(n2519) );
  XOR U2444 ( .A(p_input[123]), .B(n2518), .Z(n2520) );
  XNOR U2445 ( .A(n2521), .B(n2522), .Z(n2518) );
  AND U2446 ( .A(n192), .B(n2523), .Z(n2522) );
  XOR U2447 ( .A(n2524), .B(n2525), .Z(n2516) );
  AND U2448 ( .A(n196), .B(n2515), .Z(n2525) );
  XNOR U2449 ( .A(n2526), .B(n2513), .Z(n2515) );
  XOR U2450 ( .A(n2527), .B(n2528), .Z(n2513) );
  AND U2451 ( .A(n219), .B(n2529), .Z(n2528) );
  IV U2452 ( .A(n2524), .Z(n2526) );
  XOR U2453 ( .A(n2530), .B(n2531), .Z(n2524) );
  AND U2454 ( .A(n203), .B(n2523), .Z(n2531) );
  XNOR U2455 ( .A(n2521), .B(n2530), .Z(n2523) );
  XNOR U2456 ( .A(n2532), .B(n2533), .Z(n2521) );
  AND U2457 ( .A(n207), .B(n2534), .Z(n2533) );
  XOR U2458 ( .A(p_input[155]), .B(n2532), .Z(n2534) );
  XNOR U2459 ( .A(n2535), .B(n2536), .Z(n2532) );
  AND U2460 ( .A(n211), .B(n2537), .Z(n2536) );
  XOR U2461 ( .A(n2538), .B(n2539), .Z(n2530) );
  AND U2462 ( .A(n215), .B(n2529), .Z(n2539) );
  XNOR U2463 ( .A(n2540), .B(n2527), .Z(n2529) );
  XOR U2464 ( .A(n2541), .B(n2542), .Z(n2527) );
  AND U2465 ( .A(n238), .B(n2543), .Z(n2542) );
  IV U2466 ( .A(n2538), .Z(n2540) );
  XOR U2467 ( .A(n2544), .B(n2545), .Z(n2538) );
  AND U2468 ( .A(n222), .B(n2537), .Z(n2545) );
  XNOR U2469 ( .A(n2535), .B(n2544), .Z(n2537) );
  XNOR U2470 ( .A(n2546), .B(n2547), .Z(n2535) );
  AND U2471 ( .A(n226), .B(n2548), .Z(n2547) );
  XOR U2472 ( .A(p_input[187]), .B(n2546), .Z(n2548) );
  XNOR U2473 ( .A(n2549), .B(n2550), .Z(n2546) );
  AND U2474 ( .A(n230), .B(n2551), .Z(n2550) );
  XOR U2475 ( .A(n2552), .B(n2553), .Z(n2544) );
  AND U2476 ( .A(n234), .B(n2543), .Z(n2553) );
  XNOR U2477 ( .A(n2554), .B(n2541), .Z(n2543) );
  XOR U2478 ( .A(n2555), .B(n2556), .Z(n2541) );
  AND U2479 ( .A(n257), .B(n2557), .Z(n2556) );
  IV U2480 ( .A(n2552), .Z(n2554) );
  XOR U2481 ( .A(n2558), .B(n2559), .Z(n2552) );
  AND U2482 ( .A(n241), .B(n2551), .Z(n2559) );
  XNOR U2483 ( .A(n2549), .B(n2558), .Z(n2551) );
  XNOR U2484 ( .A(n2560), .B(n2561), .Z(n2549) );
  AND U2485 ( .A(n245), .B(n2562), .Z(n2561) );
  XOR U2486 ( .A(p_input[219]), .B(n2560), .Z(n2562) );
  XNOR U2487 ( .A(n2563), .B(n2564), .Z(n2560) );
  AND U2488 ( .A(n249), .B(n2565), .Z(n2564) );
  XOR U2489 ( .A(n2566), .B(n2567), .Z(n2558) );
  AND U2490 ( .A(n253), .B(n2557), .Z(n2567) );
  XNOR U2491 ( .A(n2568), .B(n2555), .Z(n2557) );
  XOR U2492 ( .A(n2569), .B(n2570), .Z(n2555) );
  AND U2493 ( .A(n276), .B(n2571), .Z(n2570) );
  IV U2494 ( .A(n2566), .Z(n2568) );
  XOR U2495 ( .A(n2572), .B(n2573), .Z(n2566) );
  AND U2496 ( .A(n260), .B(n2565), .Z(n2573) );
  XNOR U2497 ( .A(n2563), .B(n2572), .Z(n2565) );
  XNOR U2498 ( .A(n2574), .B(n2575), .Z(n2563) );
  AND U2499 ( .A(n264), .B(n2576), .Z(n2575) );
  XOR U2500 ( .A(p_input[251]), .B(n2574), .Z(n2576) );
  XNOR U2501 ( .A(n2577), .B(n2578), .Z(n2574) );
  AND U2502 ( .A(n268), .B(n2579), .Z(n2578) );
  XOR U2503 ( .A(n2580), .B(n2581), .Z(n2572) );
  AND U2504 ( .A(n272), .B(n2571), .Z(n2581) );
  XNOR U2505 ( .A(n2582), .B(n2569), .Z(n2571) );
  XOR U2506 ( .A(n2583), .B(n2584), .Z(n2569) );
  AND U2507 ( .A(n295), .B(n2585), .Z(n2584) );
  IV U2508 ( .A(n2580), .Z(n2582) );
  XOR U2509 ( .A(n2586), .B(n2587), .Z(n2580) );
  AND U2510 ( .A(n279), .B(n2579), .Z(n2587) );
  XNOR U2511 ( .A(n2577), .B(n2586), .Z(n2579) );
  XNOR U2512 ( .A(n2588), .B(n2589), .Z(n2577) );
  AND U2513 ( .A(n283), .B(n2590), .Z(n2589) );
  XOR U2514 ( .A(p_input[283]), .B(n2588), .Z(n2590) );
  XNOR U2515 ( .A(n2591), .B(n2592), .Z(n2588) );
  AND U2516 ( .A(n287), .B(n2593), .Z(n2592) );
  XOR U2517 ( .A(n2594), .B(n2595), .Z(n2586) );
  AND U2518 ( .A(n291), .B(n2585), .Z(n2595) );
  XNOR U2519 ( .A(n2596), .B(n2583), .Z(n2585) );
  XOR U2520 ( .A(n2597), .B(n2598), .Z(n2583) );
  AND U2521 ( .A(n314), .B(n2599), .Z(n2598) );
  IV U2522 ( .A(n2594), .Z(n2596) );
  XOR U2523 ( .A(n2600), .B(n2601), .Z(n2594) );
  AND U2524 ( .A(n298), .B(n2593), .Z(n2601) );
  XNOR U2525 ( .A(n2591), .B(n2600), .Z(n2593) );
  XNOR U2526 ( .A(n2602), .B(n2603), .Z(n2591) );
  AND U2527 ( .A(n302), .B(n2604), .Z(n2603) );
  XOR U2528 ( .A(p_input[315]), .B(n2602), .Z(n2604) );
  XNOR U2529 ( .A(n2605), .B(n2606), .Z(n2602) );
  AND U2530 ( .A(n306), .B(n2607), .Z(n2606) );
  XOR U2531 ( .A(n2608), .B(n2609), .Z(n2600) );
  AND U2532 ( .A(n310), .B(n2599), .Z(n2609) );
  XNOR U2533 ( .A(n2610), .B(n2597), .Z(n2599) );
  XOR U2534 ( .A(n2611), .B(n2612), .Z(n2597) );
  AND U2535 ( .A(n333), .B(n2613), .Z(n2612) );
  IV U2536 ( .A(n2608), .Z(n2610) );
  XOR U2537 ( .A(n2614), .B(n2615), .Z(n2608) );
  AND U2538 ( .A(n317), .B(n2607), .Z(n2615) );
  XNOR U2539 ( .A(n2605), .B(n2614), .Z(n2607) );
  XNOR U2540 ( .A(n2616), .B(n2617), .Z(n2605) );
  AND U2541 ( .A(n321), .B(n2618), .Z(n2617) );
  XOR U2542 ( .A(p_input[347]), .B(n2616), .Z(n2618) );
  XNOR U2543 ( .A(n2619), .B(n2620), .Z(n2616) );
  AND U2544 ( .A(n325), .B(n2621), .Z(n2620) );
  XOR U2545 ( .A(n2622), .B(n2623), .Z(n2614) );
  AND U2546 ( .A(n329), .B(n2613), .Z(n2623) );
  XNOR U2547 ( .A(n2624), .B(n2611), .Z(n2613) );
  XOR U2548 ( .A(n2625), .B(n2626), .Z(n2611) );
  AND U2549 ( .A(n352), .B(n2627), .Z(n2626) );
  IV U2550 ( .A(n2622), .Z(n2624) );
  XOR U2551 ( .A(n2628), .B(n2629), .Z(n2622) );
  AND U2552 ( .A(n336), .B(n2621), .Z(n2629) );
  XNOR U2553 ( .A(n2619), .B(n2628), .Z(n2621) );
  XNOR U2554 ( .A(n2630), .B(n2631), .Z(n2619) );
  AND U2555 ( .A(n340), .B(n2632), .Z(n2631) );
  XOR U2556 ( .A(p_input[379]), .B(n2630), .Z(n2632) );
  XNOR U2557 ( .A(n2633), .B(n2634), .Z(n2630) );
  AND U2558 ( .A(n344), .B(n2635), .Z(n2634) );
  XOR U2559 ( .A(n2636), .B(n2637), .Z(n2628) );
  AND U2560 ( .A(n348), .B(n2627), .Z(n2637) );
  XNOR U2561 ( .A(n2638), .B(n2625), .Z(n2627) );
  XOR U2562 ( .A(n2639), .B(n2640), .Z(n2625) );
  AND U2563 ( .A(n370), .B(n2641), .Z(n2640) );
  IV U2564 ( .A(n2636), .Z(n2638) );
  XOR U2565 ( .A(n2642), .B(n2643), .Z(n2636) );
  AND U2566 ( .A(n355), .B(n2635), .Z(n2643) );
  XNOR U2567 ( .A(n2633), .B(n2642), .Z(n2635) );
  XNOR U2568 ( .A(n2644), .B(n2645), .Z(n2633) );
  AND U2569 ( .A(n359), .B(n2646), .Z(n2645) );
  XOR U2570 ( .A(p_input[411]), .B(n2644), .Z(n2646) );
  XOR U2571 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][27] ), .B(n2647), 
        .Z(n2644) );
  AND U2572 ( .A(n362), .B(n2648), .Z(n2647) );
  XOR U2573 ( .A(n2649), .B(n2650), .Z(n2642) );
  AND U2574 ( .A(n366), .B(n2641), .Z(n2650) );
  XNOR U2575 ( .A(n2651), .B(n2639), .Z(n2641) );
  XOR U2576 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n2652), .Z(n2639) );
  AND U2577 ( .A(n378), .B(n2653), .Z(n2652) );
  IV U2578 ( .A(n2649), .Z(n2651) );
  XOR U2579 ( .A(n2654), .B(n2655), .Z(n2649) );
  AND U2580 ( .A(n373), .B(n2648), .Z(n2655) );
  XOR U2581 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][27] ), .B(n2654), 
        .Z(n2648) );
  XOR U2582 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .B(n2656), 
        .Z(n2654) );
  AND U2583 ( .A(n375), .B(n2653), .Z(n2656) );
  XOR U2584 ( .A(n2657), .B(n2658), .Z(n2653) );
  IV U2585 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .Z(n2658) );
  IV U2586 ( .A(\knn_comb_/min_val_out[0][27] ), .Z(n2657) );
  XOR U2587 ( .A(n85), .B(n2659), .Z(o[26]) );
  AND U2588 ( .A(n122), .B(n2660), .Z(n85) );
  XOR U2589 ( .A(n86), .B(n2659), .Z(n2660) );
  XOR U2590 ( .A(n2661), .B(n2662), .Z(n2659) );
  AND U2591 ( .A(n142), .B(n2663), .Z(n2662) );
  XOR U2592 ( .A(n2664), .B(n13), .Z(n86) );
  AND U2593 ( .A(n125), .B(n2665), .Z(n13) );
  XOR U2594 ( .A(n14), .B(n2664), .Z(n2665) );
  XOR U2595 ( .A(n2666), .B(n2667), .Z(n14) );
  AND U2596 ( .A(n130), .B(n2668), .Z(n2667) );
  XOR U2597 ( .A(p_input[26]), .B(n2666), .Z(n2668) );
  XNOR U2598 ( .A(n2669), .B(n2670), .Z(n2666) );
  AND U2599 ( .A(n134), .B(n2671), .Z(n2670) );
  XOR U2600 ( .A(n2672), .B(n2673), .Z(n2664) );
  AND U2601 ( .A(n138), .B(n2663), .Z(n2673) );
  XNOR U2602 ( .A(n2674), .B(n2661), .Z(n2663) );
  XOR U2603 ( .A(n2675), .B(n2676), .Z(n2661) );
  AND U2604 ( .A(n162), .B(n2677), .Z(n2676) );
  IV U2605 ( .A(n2672), .Z(n2674) );
  XOR U2606 ( .A(n2678), .B(n2679), .Z(n2672) );
  AND U2607 ( .A(n146), .B(n2671), .Z(n2679) );
  XNOR U2608 ( .A(n2669), .B(n2678), .Z(n2671) );
  XNOR U2609 ( .A(n2680), .B(n2681), .Z(n2669) );
  AND U2610 ( .A(n150), .B(n2682), .Z(n2681) );
  XOR U2611 ( .A(p_input[58]), .B(n2680), .Z(n2682) );
  XNOR U2612 ( .A(n2683), .B(n2684), .Z(n2680) );
  AND U2613 ( .A(n154), .B(n2685), .Z(n2684) );
  XOR U2614 ( .A(n2686), .B(n2687), .Z(n2678) );
  AND U2615 ( .A(n158), .B(n2677), .Z(n2687) );
  XNOR U2616 ( .A(n2688), .B(n2675), .Z(n2677) );
  XOR U2617 ( .A(n2689), .B(n2690), .Z(n2675) );
  AND U2618 ( .A(n181), .B(n2691), .Z(n2690) );
  IV U2619 ( .A(n2686), .Z(n2688) );
  XOR U2620 ( .A(n2692), .B(n2693), .Z(n2686) );
  AND U2621 ( .A(n165), .B(n2685), .Z(n2693) );
  XNOR U2622 ( .A(n2683), .B(n2692), .Z(n2685) );
  XNOR U2623 ( .A(n2694), .B(n2695), .Z(n2683) );
  AND U2624 ( .A(n169), .B(n2696), .Z(n2695) );
  XOR U2625 ( .A(p_input[90]), .B(n2694), .Z(n2696) );
  XNOR U2626 ( .A(n2697), .B(n2698), .Z(n2694) );
  AND U2627 ( .A(n173), .B(n2699), .Z(n2698) );
  XOR U2628 ( .A(n2700), .B(n2701), .Z(n2692) );
  AND U2629 ( .A(n177), .B(n2691), .Z(n2701) );
  XNOR U2630 ( .A(n2702), .B(n2689), .Z(n2691) );
  XOR U2631 ( .A(n2703), .B(n2704), .Z(n2689) );
  AND U2632 ( .A(n200), .B(n2705), .Z(n2704) );
  IV U2633 ( .A(n2700), .Z(n2702) );
  XOR U2634 ( .A(n2706), .B(n2707), .Z(n2700) );
  AND U2635 ( .A(n184), .B(n2699), .Z(n2707) );
  XNOR U2636 ( .A(n2697), .B(n2706), .Z(n2699) );
  XNOR U2637 ( .A(n2708), .B(n2709), .Z(n2697) );
  AND U2638 ( .A(n188), .B(n2710), .Z(n2709) );
  XOR U2639 ( .A(p_input[122]), .B(n2708), .Z(n2710) );
  XNOR U2640 ( .A(n2711), .B(n2712), .Z(n2708) );
  AND U2641 ( .A(n192), .B(n2713), .Z(n2712) );
  XOR U2642 ( .A(n2714), .B(n2715), .Z(n2706) );
  AND U2643 ( .A(n196), .B(n2705), .Z(n2715) );
  XNOR U2644 ( .A(n2716), .B(n2703), .Z(n2705) );
  XOR U2645 ( .A(n2717), .B(n2718), .Z(n2703) );
  AND U2646 ( .A(n219), .B(n2719), .Z(n2718) );
  IV U2647 ( .A(n2714), .Z(n2716) );
  XOR U2648 ( .A(n2720), .B(n2721), .Z(n2714) );
  AND U2649 ( .A(n203), .B(n2713), .Z(n2721) );
  XNOR U2650 ( .A(n2711), .B(n2720), .Z(n2713) );
  XNOR U2651 ( .A(n2722), .B(n2723), .Z(n2711) );
  AND U2652 ( .A(n207), .B(n2724), .Z(n2723) );
  XOR U2653 ( .A(p_input[154]), .B(n2722), .Z(n2724) );
  XNOR U2654 ( .A(n2725), .B(n2726), .Z(n2722) );
  AND U2655 ( .A(n211), .B(n2727), .Z(n2726) );
  XOR U2656 ( .A(n2728), .B(n2729), .Z(n2720) );
  AND U2657 ( .A(n215), .B(n2719), .Z(n2729) );
  XNOR U2658 ( .A(n2730), .B(n2717), .Z(n2719) );
  XOR U2659 ( .A(n2731), .B(n2732), .Z(n2717) );
  AND U2660 ( .A(n238), .B(n2733), .Z(n2732) );
  IV U2661 ( .A(n2728), .Z(n2730) );
  XOR U2662 ( .A(n2734), .B(n2735), .Z(n2728) );
  AND U2663 ( .A(n222), .B(n2727), .Z(n2735) );
  XNOR U2664 ( .A(n2725), .B(n2734), .Z(n2727) );
  XNOR U2665 ( .A(n2736), .B(n2737), .Z(n2725) );
  AND U2666 ( .A(n226), .B(n2738), .Z(n2737) );
  XOR U2667 ( .A(p_input[186]), .B(n2736), .Z(n2738) );
  XNOR U2668 ( .A(n2739), .B(n2740), .Z(n2736) );
  AND U2669 ( .A(n230), .B(n2741), .Z(n2740) );
  XOR U2670 ( .A(n2742), .B(n2743), .Z(n2734) );
  AND U2671 ( .A(n234), .B(n2733), .Z(n2743) );
  XNOR U2672 ( .A(n2744), .B(n2731), .Z(n2733) );
  XOR U2673 ( .A(n2745), .B(n2746), .Z(n2731) );
  AND U2674 ( .A(n257), .B(n2747), .Z(n2746) );
  IV U2675 ( .A(n2742), .Z(n2744) );
  XOR U2676 ( .A(n2748), .B(n2749), .Z(n2742) );
  AND U2677 ( .A(n241), .B(n2741), .Z(n2749) );
  XNOR U2678 ( .A(n2739), .B(n2748), .Z(n2741) );
  XNOR U2679 ( .A(n2750), .B(n2751), .Z(n2739) );
  AND U2680 ( .A(n245), .B(n2752), .Z(n2751) );
  XOR U2681 ( .A(p_input[218]), .B(n2750), .Z(n2752) );
  XNOR U2682 ( .A(n2753), .B(n2754), .Z(n2750) );
  AND U2683 ( .A(n249), .B(n2755), .Z(n2754) );
  XOR U2684 ( .A(n2756), .B(n2757), .Z(n2748) );
  AND U2685 ( .A(n253), .B(n2747), .Z(n2757) );
  XNOR U2686 ( .A(n2758), .B(n2745), .Z(n2747) );
  XOR U2687 ( .A(n2759), .B(n2760), .Z(n2745) );
  AND U2688 ( .A(n276), .B(n2761), .Z(n2760) );
  IV U2689 ( .A(n2756), .Z(n2758) );
  XOR U2690 ( .A(n2762), .B(n2763), .Z(n2756) );
  AND U2691 ( .A(n260), .B(n2755), .Z(n2763) );
  XNOR U2692 ( .A(n2753), .B(n2762), .Z(n2755) );
  XNOR U2693 ( .A(n2764), .B(n2765), .Z(n2753) );
  AND U2694 ( .A(n264), .B(n2766), .Z(n2765) );
  XOR U2695 ( .A(p_input[250]), .B(n2764), .Z(n2766) );
  XNOR U2696 ( .A(n2767), .B(n2768), .Z(n2764) );
  AND U2697 ( .A(n268), .B(n2769), .Z(n2768) );
  XOR U2698 ( .A(n2770), .B(n2771), .Z(n2762) );
  AND U2699 ( .A(n272), .B(n2761), .Z(n2771) );
  XNOR U2700 ( .A(n2772), .B(n2759), .Z(n2761) );
  XOR U2701 ( .A(n2773), .B(n2774), .Z(n2759) );
  AND U2702 ( .A(n295), .B(n2775), .Z(n2774) );
  IV U2703 ( .A(n2770), .Z(n2772) );
  XOR U2704 ( .A(n2776), .B(n2777), .Z(n2770) );
  AND U2705 ( .A(n279), .B(n2769), .Z(n2777) );
  XNOR U2706 ( .A(n2767), .B(n2776), .Z(n2769) );
  XNOR U2707 ( .A(n2778), .B(n2779), .Z(n2767) );
  AND U2708 ( .A(n283), .B(n2780), .Z(n2779) );
  XOR U2709 ( .A(p_input[282]), .B(n2778), .Z(n2780) );
  XNOR U2710 ( .A(n2781), .B(n2782), .Z(n2778) );
  AND U2711 ( .A(n287), .B(n2783), .Z(n2782) );
  XOR U2712 ( .A(n2784), .B(n2785), .Z(n2776) );
  AND U2713 ( .A(n291), .B(n2775), .Z(n2785) );
  XNOR U2714 ( .A(n2786), .B(n2773), .Z(n2775) );
  XOR U2715 ( .A(n2787), .B(n2788), .Z(n2773) );
  AND U2716 ( .A(n314), .B(n2789), .Z(n2788) );
  IV U2717 ( .A(n2784), .Z(n2786) );
  XOR U2718 ( .A(n2790), .B(n2791), .Z(n2784) );
  AND U2719 ( .A(n298), .B(n2783), .Z(n2791) );
  XNOR U2720 ( .A(n2781), .B(n2790), .Z(n2783) );
  XNOR U2721 ( .A(n2792), .B(n2793), .Z(n2781) );
  AND U2722 ( .A(n302), .B(n2794), .Z(n2793) );
  XOR U2723 ( .A(p_input[314]), .B(n2792), .Z(n2794) );
  XNOR U2724 ( .A(n2795), .B(n2796), .Z(n2792) );
  AND U2725 ( .A(n306), .B(n2797), .Z(n2796) );
  XOR U2726 ( .A(n2798), .B(n2799), .Z(n2790) );
  AND U2727 ( .A(n310), .B(n2789), .Z(n2799) );
  XNOR U2728 ( .A(n2800), .B(n2787), .Z(n2789) );
  XOR U2729 ( .A(n2801), .B(n2802), .Z(n2787) );
  AND U2730 ( .A(n333), .B(n2803), .Z(n2802) );
  IV U2731 ( .A(n2798), .Z(n2800) );
  XOR U2732 ( .A(n2804), .B(n2805), .Z(n2798) );
  AND U2733 ( .A(n317), .B(n2797), .Z(n2805) );
  XNOR U2734 ( .A(n2795), .B(n2804), .Z(n2797) );
  XNOR U2735 ( .A(n2806), .B(n2807), .Z(n2795) );
  AND U2736 ( .A(n321), .B(n2808), .Z(n2807) );
  XOR U2737 ( .A(p_input[346]), .B(n2806), .Z(n2808) );
  XNOR U2738 ( .A(n2809), .B(n2810), .Z(n2806) );
  AND U2739 ( .A(n325), .B(n2811), .Z(n2810) );
  XOR U2740 ( .A(n2812), .B(n2813), .Z(n2804) );
  AND U2741 ( .A(n329), .B(n2803), .Z(n2813) );
  XNOR U2742 ( .A(n2814), .B(n2801), .Z(n2803) );
  XOR U2743 ( .A(n2815), .B(n2816), .Z(n2801) );
  AND U2744 ( .A(n352), .B(n2817), .Z(n2816) );
  IV U2745 ( .A(n2812), .Z(n2814) );
  XOR U2746 ( .A(n2818), .B(n2819), .Z(n2812) );
  AND U2747 ( .A(n336), .B(n2811), .Z(n2819) );
  XNOR U2748 ( .A(n2809), .B(n2818), .Z(n2811) );
  XNOR U2749 ( .A(n2820), .B(n2821), .Z(n2809) );
  AND U2750 ( .A(n340), .B(n2822), .Z(n2821) );
  XOR U2751 ( .A(p_input[378]), .B(n2820), .Z(n2822) );
  XNOR U2752 ( .A(n2823), .B(n2824), .Z(n2820) );
  AND U2753 ( .A(n344), .B(n2825), .Z(n2824) );
  XOR U2754 ( .A(n2826), .B(n2827), .Z(n2818) );
  AND U2755 ( .A(n348), .B(n2817), .Z(n2827) );
  XNOR U2756 ( .A(n2828), .B(n2815), .Z(n2817) );
  XOR U2757 ( .A(n2829), .B(n2830), .Z(n2815) );
  AND U2758 ( .A(n370), .B(n2831), .Z(n2830) );
  IV U2759 ( .A(n2826), .Z(n2828) );
  XOR U2760 ( .A(n2832), .B(n2833), .Z(n2826) );
  AND U2761 ( .A(n355), .B(n2825), .Z(n2833) );
  XNOR U2762 ( .A(n2823), .B(n2832), .Z(n2825) );
  XNOR U2763 ( .A(n2834), .B(n2835), .Z(n2823) );
  AND U2764 ( .A(n359), .B(n2836), .Z(n2835) );
  XOR U2765 ( .A(p_input[410]), .B(n2834), .Z(n2836) );
  XOR U2766 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][26] ), .B(n2837), 
        .Z(n2834) );
  AND U2767 ( .A(n362), .B(n2838), .Z(n2837) );
  XOR U2768 ( .A(n2839), .B(n2840), .Z(n2832) );
  AND U2769 ( .A(n366), .B(n2831), .Z(n2840) );
  XNOR U2770 ( .A(n2841), .B(n2829), .Z(n2831) );
  XOR U2771 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n2842), .Z(n2829) );
  AND U2772 ( .A(n378), .B(n2843), .Z(n2842) );
  IV U2773 ( .A(n2839), .Z(n2841) );
  XOR U2774 ( .A(n2844), .B(n2845), .Z(n2839) );
  AND U2775 ( .A(n373), .B(n2838), .Z(n2845) );
  XOR U2776 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][26] ), .B(n2844), 
        .Z(n2838) );
  XOR U2777 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .B(n2846), 
        .Z(n2844) );
  AND U2778 ( .A(n375), .B(n2843), .Z(n2846) );
  XOR U2779 ( .A(\knn_comb_/min_val_out[0][26] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .Z(n2843) );
  XOR U2780 ( .A(n87), .B(n2847), .Z(o[25]) );
  AND U2781 ( .A(n122), .B(n2848), .Z(n87) );
  XOR U2782 ( .A(n88), .B(n2847), .Z(n2848) );
  XOR U2783 ( .A(n2849), .B(n2850), .Z(n2847) );
  AND U2784 ( .A(n142), .B(n2851), .Z(n2850) );
  XOR U2785 ( .A(n2852), .B(n17), .Z(n88) );
  AND U2786 ( .A(n125), .B(n2853), .Z(n17) );
  XOR U2787 ( .A(n18), .B(n2852), .Z(n2853) );
  XOR U2788 ( .A(n2854), .B(n2855), .Z(n18) );
  AND U2789 ( .A(n130), .B(n2856), .Z(n2855) );
  XOR U2790 ( .A(p_input[25]), .B(n2854), .Z(n2856) );
  XNOR U2791 ( .A(n2857), .B(n2858), .Z(n2854) );
  AND U2792 ( .A(n134), .B(n2859), .Z(n2858) );
  XOR U2793 ( .A(n2860), .B(n2861), .Z(n2852) );
  AND U2794 ( .A(n138), .B(n2851), .Z(n2861) );
  XNOR U2795 ( .A(n2862), .B(n2849), .Z(n2851) );
  XOR U2796 ( .A(n2863), .B(n2864), .Z(n2849) );
  AND U2797 ( .A(n162), .B(n2865), .Z(n2864) );
  IV U2798 ( .A(n2860), .Z(n2862) );
  XOR U2799 ( .A(n2866), .B(n2867), .Z(n2860) );
  AND U2800 ( .A(n146), .B(n2859), .Z(n2867) );
  XNOR U2801 ( .A(n2857), .B(n2866), .Z(n2859) );
  XNOR U2802 ( .A(n2868), .B(n2869), .Z(n2857) );
  AND U2803 ( .A(n150), .B(n2870), .Z(n2869) );
  XOR U2804 ( .A(p_input[57]), .B(n2868), .Z(n2870) );
  XNOR U2805 ( .A(n2871), .B(n2872), .Z(n2868) );
  AND U2806 ( .A(n154), .B(n2873), .Z(n2872) );
  XOR U2807 ( .A(n2874), .B(n2875), .Z(n2866) );
  AND U2808 ( .A(n158), .B(n2865), .Z(n2875) );
  XNOR U2809 ( .A(n2876), .B(n2863), .Z(n2865) );
  XOR U2810 ( .A(n2877), .B(n2878), .Z(n2863) );
  AND U2811 ( .A(n181), .B(n2879), .Z(n2878) );
  IV U2812 ( .A(n2874), .Z(n2876) );
  XOR U2813 ( .A(n2880), .B(n2881), .Z(n2874) );
  AND U2814 ( .A(n165), .B(n2873), .Z(n2881) );
  XNOR U2815 ( .A(n2871), .B(n2880), .Z(n2873) );
  XNOR U2816 ( .A(n2882), .B(n2883), .Z(n2871) );
  AND U2817 ( .A(n169), .B(n2884), .Z(n2883) );
  XOR U2818 ( .A(p_input[89]), .B(n2882), .Z(n2884) );
  XNOR U2819 ( .A(n2885), .B(n2886), .Z(n2882) );
  AND U2820 ( .A(n173), .B(n2887), .Z(n2886) );
  XOR U2821 ( .A(n2888), .B(n2889), .Z(n2880) );
  AND U2822 ( .A(n177), .B(n2879), .Z(n2889) );
  XNOR U2823 ( .A(n2890), .B(n2877), .Z(n2879) );
  XOR U2824 ( .A(n2891), .B(n2892), .Z(n2877) );
  AND U2825 ( .A(n200), .B(n2893), .Z(n2892) );
  IV U2826 ( .A(n2888), .Z(n2890) );
  XOR U2827 ( .A(n2894), .B(n2895), .Z(n2888) );
  AND U2828 ( .A(n184), .B(n2887), .Z(n2895) );
  XNOR U2829 ( .A(n2885), .B(n2894), .Z(n2887) );
  XNOR U2830 ( .A(n2896), .B(n2897), .Z(n2885) );
  AND U2831 ( .A(n188), .B(n2898), .Z(n2897) );
  XOR U2832 ( .A(p_input[121]), .B(n2896), .Z(n2898) );
  XNOR U2833 ( .A(n2899), .B(n2900), .Z(n2896) );
  AND U2834 ( .A(n192), .B(n2901), .Z(n2900) );
  XOR U2835 ( .A(n2902), .B(n2903), .Z(n2894) );
  AND U2836 ( .A(n196), .B(n2893), .Z(n2903) );
  XNOR U2837 ( .A(n2904), .B(n2891), .Z(n2893) );
  XOR U2838 ( .A(n2905), .B(n2906), .Z(n2891) );
  AND U2839 ( .A(n219), .B(n2907), .Z(n2906) );
  IV U2840 ( .A(n2902), .Z(n2904) );
  XOR U2841 ( .A(n2908), .B(n2909), .Z(n2902) );
  AND U2842 ( .A(n203), .B(n2901), .Z(n2909) );
  XNOR U2843 ( .A(n2899), .B(n2908), .Z(n2901) );
  XNOR U2844 ( .A(n2910), .B(n2911), .Z(n2899) );
  AND U2845 ( .A(n207), .B(n2912), .Z(n2911) );
  XOR U2846 ( .A(p_input[153]), .B(n2910), .Z(n2912) );
  XNOR U2847 ( .A(n2913), .B(n2914), .Z(n2910) );
  AND U2848 ( .A(n211), .B(n2915), .Z(n2914) );
  XOR U2849 ( .A(n2916), .B(n2917), .Z(n2908) );
  AND U2850 ( .A(n215), .B(n2907), .Z(n2917) );
  XNOR U2851 ( .A(n2918), .B(n2905), .Z(n2907) );
  XOR U2852 ( .A(n2919), .B(n2920), .Z(n2905) );
  AND U2853 ( .A(n238), .B(n2921), .Z(n2920) );
  IV U2854 ( .A(n2916), .Z(n2918) );
  XOR U2855 ( .A(n2922), .B(n2923), .Z(n2916) );
  AND U2856 ( .A(n222), .B(n2915), .Z(n2923) );
  XNOR U2857 ( .A(n2913), .B(n2922), .Z(n2915) );
  XNOR U2858 ( .A(n2924), .B(n2925), .Z(n2913) );
  AND U2859 ( .A(n226), .B(n2926), .Z(n2925) );
  XOR U2860 ( .A(p_input[185]), .B(n2924), .Z(n2926) );
  XNOR U2861 ( .A(n2927), .B(n2928), .Z(n2924) );
  AND U2862 ( .A(n230), .B(n2929), .Z(n2928) );
  XOR U2863 ( .A(n2930), .B(n2931), .Z(n2922) );
  AND U2864 ( .A(n234), .B(n2921), .Z(n2931) );
  XNOR U2865 ( .A(n2932), .B(n2919), .Z(n2921) );
  XOR U2866 ( .A(n2933), .B(n2934), .Z(n2919) );
  AND U2867 ( .A(n257), .B(n2935), .Z(n2934) );
  IV U2868 ( .A(n2930), .Z(n2932) );
  XOR U2869 ( .A(n2936), .B(n2937), .Z(n2930) );
  AND U2870 ( .A(n241), .B(n2929), .Z(n2937) );
  XNOR U2871 ( .A(n2927), .B(n2936), .Z(n2929) );
  XNOR U2872 ( .A(n2938), .B(n2939), .Z(n2927) );
  AND U2873 ( .A(n245), .B(n2940), .Z(n2939) );
  XOR U2874 ( .A(p_input[217]), .B(n2938), .Z(n2940) );
  XNOR U2875 ( .A(n2941), .B(n2942), .Z(n2938) );
  AND U2876 ( .A(n249), .B(n2943), .Z(n2942) );
  XOR U2877 ( .A(n2944), .B(n2945), .Z(n2936) );
  AND U2878 ( .A(n253), .B(n2935), .Z(n2945) );
  XNOR U2879 ( .A(n2946), .B(n2933), .Z(n2935) );
  XOR U2880 ( .A(n2947), .B(n2948), .Z(n2933) );
  AND U2881 ( .A(n276), .B(n2949), .Z(n2948) );
  IV U2882 ( .A(n2944), .Z(n2946) );
  XOR U2883 ( .A(n2950), .B(n2951), .Z(n2944) );
  AND U2884 ( .A(n260), .B(n2943), .Z(n2951) );
  XNOR U2885 ( .A(n2941), .B(n2950), .Z(n2943) );
  XNOR U2886 ( .A(n2952), .B(n2953), .Z(n2941) );
  AND U2887 ( .A(n264), .B(n2954), .Z(n2953) );
  XOR U2888 ( .A(p_input[249]), .B(n2952), .Z(n2954) );
  XNOR U2889 ( .A(n2955), .B(n2956), .Z(n2952) );
  AND U2890 ( .A(n268), .B(n2957), .Z(n2956) );
  XOR U2891 ( .A(n2958), .B(n2959), .Z(n2950) );
  AND U2892 ( .A(n272), .B(n2949), .Z(n2959) );
  XNOR U2893 ( .A(n2960), .B(n2947), .Z(n2949) );
  XOR U2894 ( .A(n2961), .B(n2962), .Z(n2947) );
  AND U2895 ( .A(n295), .B(n2963), .Z(n2962) );
  IV U2896 ( .A(n2958), .Z(n2960) );
  XOR U2897 ( .A(n2964), .B(n2965), .Z(n2958) );
  AND U2898 ( .A(n279), .B(n2957), .Z(n2965) );
  XNOR U2899 ( .A(n2955), .B(n2964), .Z(n2957) );
  XNOR U2900 ( .A(n2966), .B(n2967), .Z(n2955) );
  AND U2901 ( .A(n283), .B(n2968), .Z(n2967) );
  XOR U2902 ( .A(p_input[281]), .B(n2966), .Z(n2968) );
  XNOR U2903 ( .A(n2969), .B(n2970), .Z(n2966) );
  AND U2904 ( .A(n287), .B(n2971), .Z(n2970) );
  XOR U2905 ( .A(n2972), .B(n2973), .Z(n2964) );
  AND U2906 ( .A(n291), .B(n2963), .Z(n2973) );
  XNOR U2907 ( .A(n2974), .B(n2961), .Z(n2963) );
  XOR U2908 ( .A(n2975), .B(n2976), .Z(n2961) );
  AND U2909 ( .A(n314), .B(n2977), .Z(n2976) );
  IV U2910 ( .A(n2972), .Z(n2974) );
  XOR U2911 ( .A(n2978), .B(n2979), .Z(n2972) );
  AND U2912 ( .A(n298), .B(n2971), .Z(n2979) );
  XNOR U2913 ( .A(n2969), .B(n2978), .Z(n2971) );
  XNOR U2914 ( .A(n2980), .B(n2981), .Z(n2969) );
  AND U2915 ( .A(n302), .B(n2982), .Z(n2981) );
  XOR U2916 ( .A(p_input[313]), .B(n2980), .Z(n2982) );
  XNOR U2917 ( .A(n2983), .B(n2984), .Z(n2980) );
  AND U2918 ( .A(n306), .B(n2985), .Z(n2984) );
  XOR U2919 ( .A(n2986), .B(n2987), .Z(n2978) );
  AND U2920 ( .A(n310), .B(n2977), .Z(n2987) );
  XNOR U2921 ( .A(n2988), .B(n2975), .Z(n2977) );
  XOR U2922 ( .A(n2989), .B(n2990), .Z(n2975) );
  AND U2923 ( .A(n333), .B(n2991), .Z(n2990) );
  IV U2924 ( .A(n2986), .Z(n2988) );
  XOR U2925 ( .A(n2992), .B(n2993), .Z(n2986) );
  AND U2926 ( .A(n317), .B(n2985), .Z(n2993) );
  XNOR U2927 ( .A(n2983), .B(n2992), .Z(n2985) );
  XNOR U2928 ( .A(n2994), .B(n2995), .Z(n2983) );
  AND U2929 ( .A(n321), .B(n2996), .Z(n2995) );
  XOR U2930 ( .A(p_input[345]), .B(n2994), .Z(n2996) );
  XNOR U2931 ( .A(n2997), .B(n2998), .Z(n2994) );
  AND U2932 ( .A(n325), .B(n2999), .Z(n2998) );
  XOR U2933 ( .A(n3000), .B(n3001), .Z(n2992) );
  AND U2934 ( .A(n329), .B(n2991), .Z(n3001) );
  XNOR U2935 ( .A(n3002), .B(n2989), .Z(n2991) );
  XOR U2936 ( .A(n3003), .B(n3004), .Z(n2989) );
  AND U2937 ( .A(n352), .B(n3005), .Z(n3004) );
  IV U2938 ( .A(n3000), .Z(n3002) );
  XOR U2939 ( .A(n3006), .B(n3007), .Z(n3000) );
  AND U2940 ( .A(n336), .B(n2999), .Z(n3007) );
  XNOR U2941 ( .A(n2997), .B(n3006), .Z(n2999) );
  XNOR U2942 ( .A(n3008), .B(n3009), .Z(n2997) );
  AND U2943 ( .A(n340), .B(n3010), .Z(n3009) );
  XOR U2944 ( .A(p_input[377]), .B(n3008), .Z(n3010) );
  XNOR U2945 ( .A(n3011), .B(n3012), .Z(n3008) );
  AND U2946 ( .A(n344), .B(n3013), .Z(n3012) );
  XOR U2947 ( .A(n3014), .B(n3015), .Z(n3006) );
  AND U2948 ( .A(n348), .B(n3005), .Z(n3015) );
  XNOR U2949 ( .A(n3016), .B(n3003), .Z(n3005) );
  XOR U2950 ( .A(n3017), .B(n3018), .Z(n3003) );
  AND U2951 ( .A(n370), .B(n3019), .Z(n3018) );
  IV U2952 ( .A(n3014), .Z(n3016) );
  XOR U2953 ( .A(n3020), .B(n3021), .Z(n3014) );
  AND U2954 ( .A(n355), .B(n3013), .Z(n3021) );
  XNOR U2955 ( .A(n3011), .B(n3020), .Z(n3013) );
  XNOR U2956 ( .A(n3022), .B(n3023), .Z(n3011) );
  AND U2957 ( .A(n359), .B(n3024), .Z(n3023) );
  XOR U2958 ( .A(p_input[409]), .B(n3022), .Z(n3024) );
  XOR U2959 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][25] ), .B(n3025), 
        .Z(n3022) );
  AND U2960 ( .A(n362), .B(n3026), .Z(n3025) );
  XOR U2961 ( .A(n3027), .B(n3028), .Z(n3020) );
  AND U2962 ( .A(n366), .B(n3019), .Z(n3028) );
  XNOR U2963 ( .A(n3029), .B(n3017), .Z(n3019) );
  XOR U2964 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n3030), .Z(n3017) );
  AND U2965 ( .A(n378), .B(n3031), .Z(n3030) );
  IV U2966 ( .A(n3027), .Z(n3029) );
  XOR U2967 ( .A(n3032), .B(n3033), .Z(n3027) );
  AND U2968 ( .A(n373), .B(n3026), .Z(n3033) );
  XOR U2969 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][25] ), .B(n3032), 
        .Z(n3026) );
  XOR U2970 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .B(n3034), 
        .Z(n3032) );
  AND U2971 ( .A(n375), .B(n3031), .Z(n3034) );
  XOR U2972 ( .A(\knn_comb_/min_val_out[0][25] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .Z(n3031) );
  XOR U2973 ( .A(n89), .B(n3035), .Z(o[24]) );
  AND U2974 ( .A(n122), .B(n3036), .Z(n89) );
  XOR U2975 ( .A(n90), .B(n3035), .Z(n3036) );
  XOR U2976 ( .A(n3037), .B(n3038), .Z(n3035) );
  AND U2977 ( .A(n142), .B(n3039), .Z(n3038) );
  XOR U2978 ( .A(n3040), .B(n19), .Z(n90) );
  AND U2979 ( .A(n125), .B(n3041), .Z(n19) );
  XOR U2980 ( .A(n20), .B(n3040), .Z(n3041) );
  XOR U2981 ( .A(n3042), .B(n3043), .Z(n20) );
  AND U2982 ( .A(n130), .B(n3044), .Z(n3043) );
  XOR U2983 ( .A(p_input[24]), .B(n3042), .Z(n3044) );
  XNOR U2984 ( .A(n3045), .B(n3046), .Z(n3042) );
  AND U2985 ( .A(n134), .B(n3047), .Z(n3046) );
  XOR U2986 ( .A(n3048), .B(n3049), .Z(n3040) );
  AND U2987 ( .A(n138), .B(n3039), .Z(n3049) );
  XNOR U2988 ( .A(n3050), .B(n3037), .Z(n3039) );
  XOR U2989 ( .A(n3051), .B(n3052), .Z(n3037) );
  AND U2990 ( .A(n162), .B(n3053), .Z(n3052) );
  IV U2991 ( .A(n3048), .Z(n3050) );
  XOR U2992 ( .A(n3054), .B(n3055), .Z(n3048) );
  AND U2993 ( .A(n146), .B(n3047), .Z(n3055) );
  XNOR U2994 ( .A(n3045), .B(n3054), .Z(n3047) );
  XNOR U2995 ( .A(n3056), .B(n3057), .Z(n3045) );
  AND U2996 ( .A(n150), .B(n3058), .Z(n3057) );
  XOR U2997 ( .A(p_input[56]), .B(n3056), .Z(n3058) );
  XNOR U2998 ( .A(n3059), .B(n3060), .Z(n3056) );
  AND U2999 ( .A(n154), .B(n3061), .Z(n3060) );
  XOR U3000 ( .A(n3062), .B(n3063), .Z(n3054) );
  AND U3001 ( .A(n158), .B(n3053), .Z(n3063) );
  XNOR U3002 ( .A(n3064), .B(n3051), .Z(n3053) );
  XOR U3003 ( .A(n3065), .B(n3066), .Z(n3051) );
  AND U3004 ( .A(n181), .B(n3067), .Z(n3066) );
  IV U3005 ( .A(n3062), .Z(n3064) );
  XOR U3006 ( .A(n3068), .B(n3069), .Z(n3062) );
  AND U3007 ( .A(n165), .B(n3061), .Z(n3069) );
  XNOR U3008 ( .A(n3059), .B(n3068), .Z(n3061) );
  XNOR U3009 ( .A(n3070), .B(n3071), .Z(n3059) );
  AND U3010 ( .A(n169), .B(n3072), .Z(n3071) );
  XOR U3011 ( .A(p_input[88]), .B(n3070), .Z(n3072) );
  XNOR U3012 ( .A(n3073), .B(n3074), .Z(n3070) );
  AND U3013 ( .A(n173), .B(n3075), .Z(n3074) );
  XOR U3014 ( .A(n3076), .B(n3077), .Z(n3068) );
  AND U3015 ( .A(n177), .B(n3067), .Z(n3077) );
  XNOR U3016 ( .A(n3078), .B(n3065), .Z(n3067) );
  XOR U3017 ( .A(n3079), .B(n3080), .Z(n3065) );
  AND U3018 ( .A(n200), .B(n3081), .Z(n3080) );
  IV U3019 ( .A(n3076), .Z(n3078) );
  XOR U3020 ( .A(n3082), .B(n3083), .Z(n3076) );
  AND U3021 ( .A(n184), .B(n3075), .Z(n3083) );
  XNOR U3022 ( .A(n3073), .B(n3082), .Z(n3075) );
  XNOR U3023 ( .A(n3084), .B(n3085), .Z(n3073) );
  AND U3024 ( .A(n188), .B(n3086), .Z(n3085) );
  XOR U3025 ( .A(p_input[120]), .B(n3084), .Z(n3086) );
  XNOR U3026 ( .A(n3087), .B(n3088), .Z(n3084) );
  AND U3027 ( .A(n192), .B(n3089), .Z(n3088) );
  XOR U3028 ( .A(n3090), .B(n3091), .Z(n3082) );
  AND U3029 ( .A(n196), .B(n3081), .Z(n3091) );
  XNOR U3030 ( .A(n3092), .B(n3079), .Z(n3081) );
  XOR U3031 ( .A(n3093), .B(n3094), .Z(n3079) );
  AND U3032 ( .A(n219), .B(n3095), .Z(n3094) );
  IV U3033 ( .A(n3090), .Z(n3092) );
  XOR U3034 ( .A(n3096), .B(n3097), .Z(n3090) );
  AND U3035 ( .A(n203), .B(n3089), .Z(n3097) );
  XNOR U3036 ( .A(n3087), .B(n3096), .Z(n3089) );
  XNOR U3037 ( .A(n3098), .B(n3099), .Z(n3087) );
  AND U3038 ( .A(n207), .B(n3100), .Z(n3099) );
  XOR U3039 ( .A(p_input[152]), .B(n3098), .Z(n3100) );
  XNOR U3040 ( .A(n3101), .B(n3102), .Z(n3098) );
  AND U3041 ( .A(n211), .B(n3103), .Z(n3102) );
  XOR U3042 ( .A(n3104), .B(n3105), .Z(n3096) );
  AND U3043 ( .A(n215), .B(n3095), .Z(n3105) );
  XNOR U3044 ( .A(n3106), .B(n3093), .Z(n3095) );
  XOR U3045 ( .A(n3107), .B(n3108), .Z(n3093) );
  AND U3046 ( .A(n238), .B(n3109), .Z(n3108) );
  IV U3047 ( .A(n3104), .Z(n3106) );
  XOR U3048 ( .A(n3110), .B(n3111), .Z(n3104) );
  AND U3049 ( .A(n222), .B(n3103), .Z(n3111) );
  XNOR U3050 ( .A(n3101), .B(n3110), .Z(n3103) );
  XNOR U3051 ( .A(n3112), .B(n3113), .Z(n3101) );
  AND U3052 ( .A(n226), .B(n3114), .Z(n3113) );
  XOR U3053 ( .A(p_input[184]), .B(n3112), .Z(n3114) );
  XNOR U3054 ( .A(n3115), .B(n3116), .Z(n3112) );
  AND U3055 ( .A(n230), .B(n3117), .Z(n3116) );
  XOR U3056 ( .A(n3118), .B(n3119), .Z(n3110) );
  AND U3057 ( .A(n234), .B(n3109), .Z(n3119) );
  XNOR U3058 ( .A(n3120), .B(n3107), .Z(n3109) );
  XOR U3059 ( .A(n3121), .B(n3122), .Z(n3107) );
  AND U3060 ( .A(n257), .B(n3123), .Z(n3122) );
  IV U3061 ( .A(n3118), .Z(n3120) );
  XOR U3062 ( .A(n3124), .B(n3125), .Z(n3118) );
  AND U3063 ( .A(n241), .B(n3117), .Z(n3125) );
  XNOR U3064 ( .A(n3115), .B(n3124), .Z(n3117) );
  XNOR U3065 ( .A(n3126), .B(n3127), .Z(n3115) );
  AND U3066 ( .A(n245), .B(n3128), .Z(n3127) );
  XOR U3067 ( .A(p_input[216]), .B(n3126), .Z(n3128) );
  XNOR U3068 ( .A(n3129), .B(n3130), .Z(n3126) );
  AND U3069 ( .A(n249), .B(n3131), .Z(n3130) );
  XOR U3070 ( .A(n3132), .B(n3133), .Z(n3124) );
  AND U3071 ( .A(n253), .B(n3123), .Z(n3133) );
  XNOR U3072 ( .A(n3134), .B(n3121), .Z(n3123) );
  XOR U3073 ( .A(n3135), .B(n3136), .Z(n3121) );
  AND U3074 ( .A(n276), .B(n3137), .Z(n3136) );
  IV U3075 ( .A(n3132), .Z(n3134) );
  XOR U3076 ( .A(n3138), .B(n3139), .Z(n3132) );
  AND U3077 ( .A(n260), .B(n3131), .Z(n3139) );
  XNOR U3078 ( .A(n3129), .B(n3138), .Z(n3131) );
  XNOR U3079 ( .A(n3140), .B(n3141), .Z(n3129) );
  AND U3080 ( .A(n264), .B(n3142), .Z(n3141) );
  XOR U3081 ( .A(p_input[248]), .B(n3140), .Z(n3142) );
  XNOR U3082 ( .A(n3143), .B(n3144), .Z(n3140) );
  AND U3083 ( .A(n268), .B(n3145), .Z(n3144) );
  XOR U3084 ( .A(n3146), .B(n3147), .Z(n3138) );
  AND U3085 ( .A(n272), .B(n3137), .Z(n3147) );
  XNOR U3086 ( .A(n3148), .B(n3135), .Z(n3137) );
  XOR U3087 ( .A(n3149), .B(n3150), .Z(n3135) );
  AND U3088 ( .A(n295), .B(n3151), .Z(n3150) );
  IV U3089 ( .A(n3146), .Z(n3148) );
  XOR U3090 ( .A(n3152), .B(n3153), .Z(n3146) );
  AND U3091 ( .A(n279), .B(n3145), .Z(n3153) );
  XNOR U3092 ( .A(n3143), .B(n3152), .Z(n3145) );
  XNOR U3093 ( .A(n3154), .B(n3155), .Z(n3143) );
  AND U3094 ( .A(n283), .B(n3156), .Z(n3155) );
  XOR U3095 ( .A(p_input[280]), .B(n3154), .Z(n3156) );
  XNOR U3096 ( .A(n3157), .B(n3158), .Z(n3154) );
  AND U3097 ( .A(n287), .B(n3159), .Z(n3158) );
  XOR U3098 ( .A(n3160), .B(n3161), .Z(n3152) );
  AND U3099 ( .A(n291), .B(n3151), .Z(n3161) );
  XNOR U3100 ( .A(n3162), .B(n3149), .Z(n3151) );
  XOR U3101 ( .A(n3163), .B(n3164), .Z(n3149) );
  AND U3102 ( .A(n314), .B(n3165), .Z(n3164) );
  IV U3103 ( .A(n3160), .Z(n3162) );
  XOR U3104 ( .A(n3166), .B(n3167), .Z(n3160) );
  AND U3105 ( .A(n298), .B(n3159), .Z(n3167) );
  XNOR U3106 ( .A(n3157), .B(n3166), .Z(n3159) );
  XNOR U3107 ( .A(n3168), .B(n3169), .Z(n3157) );
  AND U3108 ( .A(n302), .B(n3170), .Z(n3169) );
  XOR U3109 ( .A(p_input[312]), .B(n3168), .Z(n3170) );
  XNOR U3110 ( .A(n3171), .B(n3172), .Z(n3168) );
  AND U3111 ( .A(n306), .B(n3173), .Z(n3172) );
  XOR U3112 ( .A(n3174), .B(n3175), .Z(n3166) );
  AND U3113 ( .A(n310), .B(n3165), .Z(n3175) );
  XNOR U3114 ( .A(n3176), .B(n3163), .Z(n3165) );
  XOR U3115 ( .A(n3177), .B(n3178), .Z(n3163) );
  AND U3116 ( .A(n333), .B(n3179), .Z(n3178) );
  IV U3117 ( .A(n3174), .Z(n3176) );
  XOR U3118 ( .A(n3180), .B(n3181), .Z(n3174) );
  AND U3119 ( .A(n317), .B(n3173), .Z(n3181) );
  XNOR U3120 ( .A(n3171), .B(n3180), .Z(n3173) );
  XNOR U3121 ( .A(n3182), .B(n3183), .Z(n3171) );
  AND U3122 ( .A(n321), .B(n3184), .Z(n3183) );
  XOR U3123 ( .A(p_input[344]), .B(n3182), .Z(n3184) );
  XNOR U3124 ( .A(n3185), .B(n3186), .Z(n3182) );
  AND U3125 ( .A(n325), .B(n3187), .Z(n3186) );
  XOR U3126 ( .A(n3188), .B(n3189), .Z(n3180) );
  AND U3127 ( .A(n329), .B(n3179), .Z(n3189) );
  XNOR U3128 ( .A(n3190), .B(n3177), .Z(n3179) );
  XOR U3129 ( .A(n3191), .B(n3192), .Z(n3177) );
  AND U3130 ( .A(n352), .B(n3193), .Z(n3192) );
  IV U3131 ( .A(n3188), .Z(n3190) );
  XOR U3132 ( .A(n3194), .B(n3195), .Z(n3188) );
  AND U3133 ( .A(n336), .B(n3187), .Z(n3195) );
  XNOR U3134 ( .A(n3185), .B(n3194), .Z(n3187) );
  XNOR U3135 ( .A(n3196), .B(n3197), .Z(n3185) );
  AND U3136 ( .A(n340), .B(n3198), .Z(n3197) );
  XOR U3137 ( .A(p_input[376]), .B(n3196), .Z(n3198) );
  XNOR U3138 ( .A(n3199), .B(n3200), .Z(n3196) );
  AND U3139 ( .A(n344), .B(n3201), .Z(n3200) );
  XOR U3140 ( .A(n3202), .B(n3203), .Z(n3194) );
  AND U3141 ( .A(n348), .B(n3193), .Z(n3203) );
  XNOR U3142 ( .A(n3204), .B(n3191), .Z(n3193) );
  XOR U3143 ( .A(n3205), .B(n3206), .Z(n3191) );
  AND U3144 ( .A(n370), .B(n3207), .Z(n3206) );
  IV U3145 ( .A(n3202), .Z(n3204) );
  XOR U3146 ( .A(n3208), .B(n3209), .Z(n3202) );
  AND U3147 ( .A(n355), .B(n3201), .Z(n3209) );
  XNOR U3148 ( .A(n3199), .B(n3208), .Z(n3201) );
  XNOR U3149 ( .A(n3210), .B(n3211), .Z(n3199) );
  AND U3150 ( .A(n359), .B(n3212), .Z(n3211) );
  XOR U3151 ( .A(p_input[408]), .B(n3210), .Z(n3212) );
  XOR U3152 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][24] ), .B(n3213), 
        .Z(n3210) );
  AND U3153 ( .A(n362), .B(n3214), .Z(n3213) );
  XOR U3154 ( .A(n3215), .B(n3216), .Z(n3208) );
  AND U3155 ( .A(n366), .B(n3207), .Z(n3216) );
  XNOR U3156 ( .A(n3217), .B(n3205), .Z(n3207) );
  XOR U3157 ( .A(\knn_comb_/min_val_out[0][24] ), .B(n3218), .Z(n3205) );
  AND U3158 ( .A(n378), .B(n3219), .Z(n3218) );
  IV U3159 ( .A(n3215), .Z(n3217) );
  XOR U3160 ( .A(n3220), .B(n3221), .Z(n3215) );
  AND U3161 ( .A(n373), .B(n3214), .Z(n3221) );
  XOR U3162 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][24] ), .B(n3220), 
        .Z(n3214) );
  XOR U3163 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .B(n3222), 
        .Z(n3220) );
  AND U3164 ( .A(n375), .B(n3219), .Z(n3222) );
  XOR U3165 ( .A(\knn_comb_/min_val_out[0][24] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .Z(n3219) );
  XOR U3166 ( .A(n91), .B(n3223), .Z(o[23]) );
  AND U3167 ( .A(n122), .B(n3224), .Z(n91) );
  XOR U3168 ( .A(n92), .B(n3223), .Z(n3224) );
  XOR U3169 ( .A(n3225), .B(n3226), .Z(n3223) );
  AND U3170 ( .A(n142), .B(n3227), .Z(n3226) );
  XOR U3171 ( .A(n3228), .B(n21), .Z(n92) );
  AND U3172 ( .A(n125), .B(n3229), .Z(n21) );
  XOR U3173 ( .A(n22), .B(n3228), .Z(n3229) );
  XOR U3174 ( .A(n3230), .B(n3231), .Z(n22) );
  AND U3175 ( .A(n130), .B(n3232), .Z(n3231) );
  XOR U3176 ( .A(p_input[23]), .B(n3230), .Z(n3232) );
  XNOR U3177 ( .A(n3233), .B(n3234), .Z(n3230) );
  AND U3178 ( .A(n134), .B(n3235), .Z(n3234) );
  XOR U3179 ( .A(n3236), .B(n3237), .Z(n3228) );
  AND U3180 ( .A(n138), .B(n3227), .Z(n3237) );
  XNOR U3181 ( .A(n3238), .B(n3225), .Z(n3227) );
  XOR U3182 ( .A(n3239), .B(n3240), .Z(n3225) );
  AND U3183 ( .A(n162), .B(n3241), .Z(n3240) );
  IV U3184 ( .A(n3236), .Z(n3238) );
  XOR U3185 ( .A(n3242), .B(n3243), .Z(n3236) );
  AND U3186 ( .A(n146), .B(n3235), .Z(n3243) );
  XNOR U3187 ( .A(n3233), .B(n3242), .Z(n3235) );
  XNOR U3188 ( .A(n3244), .B(n3245), .Z(n3233) );
  AND U3189 ( .A(n150), .B(n3246), .Z(n3245) );
  XOR U3190 ( .A(p_input[55]), .B(n3244), .Z(n3246) );
  XNOR U3191 ( .A(n3247), .B(n3248), .Z(n3244) );
  AND U3192 ( .A(n154), .B(n3249), .Z(n3248) );
  XOR U3193 ( .A(n3250), .B(n3251), .Z(n3242) );
  AND U3194 ( .A(n158), .B(n3241), .Z(n3251) );
  XNOR U3195 ( .A(n3252), .B(n3239), .Z(n3241) );
  XOR U3196 ( .A(n3253), .B(n3254), .Z(n3239) );
  AND U3197 ( .A(n181), .B(n3255), .Z(n3254) );
  IV U3198 ( .A(n3250), .Z(n3252) );
  XOR U3199 ( .A(n3256), .B(n3257), .Z(n3250) );
  AND U3200 ( .A(n165), .B(n3249), .Z(n3257) );
  XNOR U3201 ( .A(n3247), .B(n3256), .Z(n3249) );
  XNOR U3202 ( .A(n3258), .B(n3259), .Z(n3247) );
  AND U3203 ( .A(n169), .B(n3260), .Z(n3259) );
  XOR U3204 ( .A(p_input[87]), .B(n3258), .Z(n3260) );
  XNOR U3205 ( .A(n3261), .B(n3262), .Z(n3258) );
  AND U3206 ( .A(n173), .B(n3263), .Z(n3262) );
  XOR U3207 ( .A(n3264), .B(n3265), .Z(n3256) );
  AND U3208 ( .A(n177), .B(n3255), .Z(n3265) );
  XNOR U3209 ( .A(n3266), .B(n3253), .Z(n3255) );
  XOR U3210 ( .A(n3267), .B(n3268), .Z(n3253) );
  AND U3211 ( .A(n200), .B(n3269), .Z(n3268) );
  IV U3212 ( .A(n3264), .Z(n3266) );
  XOR U3213 ( .A(n3270), .B(n3271), .Z(n3264) );
  AND U3214 ( .A(n184), .B(n3263), .Z(n3271) );
  XNOR U3215 ( .A(n3261), .B(n3270), .Z(n3263) );
  XNOR U3216 ( .A(n3272), .B(n3273), .Z(n3261) );
  AND U3217 ( .A(n188), .B(n3274), .Z(n3273) );
  XOR U3218 ( .A(p_input[119]), .B(n3272), .Z(n3274) );
  XNOR U3219 ( .A(n3275), .B(n3276), .Z(n3272) );
  AND U3220 ( .A(n192), .B(n3277), .Z(n3276) );
  XOR U3221 ( .A(n3278), .B(n3279), .Z(n3270) );
  AND U3222 ( .A(n196), .B(n3269), .Z(n3279) );
  XNOR U3223 ( .A(n3280), .B(n3267), .Z(n3269) );
  XOR U3224 ( .A(n3281), .B(n3282), .Z(n3267) );
  AND U3225 ( .A(n219), .B(n3283), .Z(n3282) );
  IV U3226 ( .A(n3278), .Z(n3280) );
  XOR U3227 ( .A(n3284), .B(n3285), .Z(n3278) );
  AND U3228 ( .A(n203), .B(n3277), .Z(n3285) );
  XNOR U3229 ( .A(n3275), .B(n3284), .Z(n3277) );
  XNOR U3230 ( .A(n3286), .B(n3287), .Z(n3275) );
  AND U3231 ( .A(n207), .B(n3288), .Z(n3287) );
  XOR U3232 ( .A(p_input[151]), .B(n3286), .Z(n3288) );
  XNOR U3233 ( .A(n3289), .B(n3290), .Z(n3286) );
  AND U3234 ( .A(n211), .B(n3291), .Z(n3290) );
  XOR U3235 ( .A(n3292), .B(n3293), .Z(n3284) );
  AND U3236 ( .A(n215), .B(n3283), .Z(n3293) );
  XNOR U3237 ( .A(n3294), .B(n3281), .Z(n3283) );
  XOR U3238 ( .A(n3295), .B(n3296), .Z(n3281) );
  AND U3239 ( .A(n238), .B(n3297), .Z(n3296) );
  IV U3240 ( .A(n3292), .Z(n3294) );
  XOR U3241 ( .A(n3298), .B(n3299), .Z(n3292) );
  AND U3242 ( .A(n222), .B(n3291), .Z(n3299) );
  XNOR U3243 ( .A(n3289), .B(n3298), .Z(n3291) );
  XNOR U3244 ( .A(n3300), .B(n3301), .Z(n3289) );
  AND U3245 ( .A(n226), .B(n3302), .Z(n3301) );
  XOR U3246 ( .A(p_input[183]), .B(n3300), .Z(n3302) );
  XNOR U3247 ( .A(n3303), .B(n3304), .Z(n3300) );
  AND U3248 ( .A(n230), .B(n3305), .Z(n3304) );
  XOR U3249 ( .A(n3306), .B(n3307), .Z(n3298) );
  AND U3250 ( .A(n234), .B(n3297), .Z(n3307) );
  XNOR U3251 ( .A(n3308), .B(n3295), .Z(n3297) );
  XOR U3252 ( .A(n3309), .B(n3310), .Z(n3295) );
  AND U3253 ( .A(n257), .B(n3311), .Z(n3310) );
  IV U3254 ( .A(n3306), .Z(n3308) );
  XOR U3255 ( .A(n3312), .B(n3313), .Z(n3306) );
  AND U3256 ( .A(n241), .B(n3305), .Z(n3313) );
  XNOR U3257 ( .A(n3303), .B(n3312), .Z(n3305) );
  XNOR U3258 ( .A(n3314), .B(n3315), .Z(n3303) );
  AND U3259 ( .A(n245), .B(n3316), .Z(n3315) );
  XOR U3260 ( .A(p_input[215]), .B(n3314), .Z(n3316) );
  XNOR U3261 ( .A(n3317), .B(n3318), .Z(n3314) );
  AND U3262 ( .A(n249), .B(n3319), .Z(n3318) );
  XOR U3263 ( .A(n3320), .B(n3321), .Z(n3312) );
  AND U3264 ( .A(n253), .B(n3311), .Z(n3321) );
  XNOR U3265 ( .A(n3322), .B(n3309), .Z(n3311) );
  XOR U3266 ( .A(n3323), .B(n3324), .Z(n3309) );
  AND U3267 ( .A(n276), .B(n3325), .Z(n3324) );
  IV U3268 ( .A(n3320), .Z(n3322) );
  XOR U3269 ( .A(n3326), .B(n3327), .Z(n3320) );
  AND U3270 ( .A(n260), .B(n3319), .Z(n3327) );
  XNOR U3271 ( .A(n3317), .B(n3326), .Z(n3319) );
  XNOR U3272 ( .A(n3328), .B(n3329), .Z(n3317) );
  AND U3273 ( .A(n264), .B(n3330), .Z(n3329) );
  XOR U3274 ( .A(p_input[247]), .B(n3328), .Z(n3330) );
  XNOR U3275 ( .A(n3331), .B(n3332), .Z(n3328) );
  AND U3276 ( .A(n268), .B(n3333), .Z(n3332) );
  XOR U3277 ( .A(n3334), .B(n3335), .Z(n3326) );
  AND U3278 ( .A(n272), .B(n3325), .Z(n3335) );
  XNOR U3279 ( .A(n3336), .B(n3323), .Z(n3325) );
  XOR U3280 ( .A(n3337), .B(n3338), .Z(n3323) );
  AND U3281 ( .A(n295), .B(n3339), .Z(n3338) );
  IV U3282 ( .A(n3334), .Z(n3336) );
  XOR U3283 ( .A(n3340), .B(n3341), .Z(n3334) );
  AND U3284 ( .A(n279), .B(n3333), .Z(n3341) );
  XNOR U3285 ( .A(n3331), .B(n3340), .Z(n3333) );
  XNOR U3286 ( .A(n3342), .B(n3343), .Z(n3331) );
  AND U3287 ( .A(n283), .B(n3344), .Z(n3343) );
  XOR U3288 ( .A(p_input[279]), .B(n3342), .Z(n3344) );
  XNOR U3289 ( .A(n3345), .B(n3346), .Z(n3342) );
  AND U3290 ( .A(n287), .B(n3347), .Z(n3346) );
  XOR U3291 ( .A(n3348), .B(n3349), .Z(n3340) );
  AND U3292 ( .A(n291), .B(n3339), .Z(n3349) );
  XNOR U3293 ( .A(n3350), .B(n3337), .Z(n3339) );
  XOR U3294 ( .A(n3351), .B(n3352), .Z(n3337) );
  AND U3295 ( .A(n314), .B(n3353), .Z(n3352) );
  IV U3296 ( .A(n3348), .Z(n3350) );
  XOR U3297 ( .A(n3354), .B(n3355), .Z(n3348) );
  AND U3298 ( .A(n298), .B(n3347), .Z(n3355) );
  XNOR U3299 ( .A(n3345), .B(n3354), .Z(n3347) );
  XNOR U3300 ( .A(n3356), .B(n3357), .Z(n3345) );
  AND U3301 ( .A(n302), .B(n3358), .Z(n3357) );
  XOR U3302 ( .A(p_input[311]), .B(n3356), .Z(n3358) );
  XNOR U3303 ( .A(n3359), .B(n3360), .Z(n3356) );
  AND U3304 ( .A(n306), .B(n3361), .Z(n3360) );
  XOR U3305 ( .A(n3362), .B(n3363), .Z(n3354) );
  AND U3306 ( .A(n310), .B(n3353), .Z(n3363) );
  XNOR U3307 ( .A(n3364), .B(n3351), .Z(n3353) );
  XOR U3308 ( .A(n3365), .B(n3366), .Z(n3351) );
  AND U3309 ( .A(n333), .B(n3367), .Z(n3366) );
  IV U3310 ( .A(n3362), .Z(n3364) );
  XOR U3311 ( .A(n3368), .B(n3369), .Z(n3362) );
  AND U3312 ( .A(n317), .B(n3361), .Z(n3369) );
  XNOR U3313 ( .A(n3359), .B(n3368), .Z(n3361) );
  XNOR U3314 ( .A(n3370), .B(n3371), .Z(n3359) );
  AND U3315 ( .A(n321), .B(n3372), .Z(n3371) );
  XOR U3316 ( .A(p_input[343]), .B(n3370), .Z(n3372) );
  XNOR U3317 ( .A(n3373), .B(n3374), .Z(n3370) );
  AND U3318 ( .A(n325), .B(n3375), .Z(n3374) );
  XOR U3319 ( .A(n3376), .B(n3377), .Z(n3368) );
  AND U3320 ( .A(n329), .B(n3367), .Z(n3377) );
  XNOR U3321 ( .A(n3378), .B(n3365), .Z(n3367) );
  XOR U3322 ( .A(n3379), .B(n3380), .Z(n3365) );
  AND U3323 ( .A(n352), .B(n3381), .Z(n3380) );
  IV U3324 ( .A(n3376), .Z(n3378) );
  XOR U3325 ( .A(n3382), .B(n3383), .Z(n3376) );
  AND U3326 ( .A(n336), .B(n3375), .Z(n3383) );
  XNOR U3327 ( .A(n3373), .B(n3382), .Z(n3375) );
  XNOR U3328 ( .A(n3384), .B(n3385), .Z(n3373) );
  AND U3329 ( .A(n340), .B(n3386), .Z(n3385) );
  XOR U3330 ( .A(p_input[375]), .B(n3384), .Z(n3386) );
  XNOR U3331 ( .A(n3387), .B(n3388), .Z(n3384) );
  AND U3332 ( .A(n344), .B(n3389), .Z(n3388) );
  XOR U3333 ( .A(n3390), .B(n3391), .Z(n3382) );
  AND U3334 ( .A(n348), .B(n3381), .Z(n3391) );
  XNOR U3335 ( .A(n3392), .B(n3379), .Z(n3381) );
  XOR U3336 ( .A(n3393), .B(n3394), .Z(n3379) );
  AND U3337 ( .A(n370), .B(n3395), .Z(n3394) );
  IV U3338 ( .A(n3390), .Z(n3392) );
  XOR U3339 ( .A(n3396), .B(n3397), .Z(n3390) );
  AND U3340 ( .A(n355), .B(n3389), .Z(n3397) );
  XNOR U3341 ( .A(n3387), .B(n3396), .Z(n3389) );
  XNOR U3342 ( .A(n3398), .B(n3399), .Z(n3387) );
  AND U3343 ( .A(n359), .B(n3400), .Z(n3399) );
  XOR U3344 ( .A(p_input[407]), .B(n3398), .Z(n3400) );
  XOR U3345 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][23] ), .B(n3401), 
        .Z(n3398) );
  AND U3346 ( .A(n362), .B(n3402), .Z(n3401) );
  XOR U3347 ( .A(n3403), .B(n3404), .Z(n3396) );
  AND U3348 ( .A(n366), .B(n3395), .Z(n3404) );
  XNOR U3349 ( .A(n3405), .B(n3393), .Z(n3395) );
  XOR U3350 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n3406), .Z(n3393) );
  AND U3351 ( .A(n378), .B(n3407), .Z(n3406) );
  IV U3352 ( .A(n3403), .Z(n3405) );
  XOR U3353 ( .A(n3408), .B(n3409), .Z(n3403) );
  AND U3354 ( .A(n373), .B(n3402), .Z(n3409) );
  XOR U3355 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][23] ), .B(n3408), 
        .Z(n3402) );
  XOR U3356 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .B(n3410), 
        .Z(n3408) );
  AND U3357 ( .A(n375), .B(n3407), .Z(n3410) );
  XOR U3358 ( .A(n3411), .B(n3412), .Z(n3407) );
  IV U3359 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .Z(n3412) );
  IV U3360 ( .A(\knn_comb_/min_val_out[0][23] ), .Z(n3411) );
  XOR U3361 ( .A(n93), .B(n3413), .Z(o[22]) );
  AND U3362 ( .A(n122), .B(n3414), .Z(n93) );
  XOR U3363 ( .A(n94), .B(n3413), .Z(n3414) );
  XOR U3364 ( .A(n3415), .B(n3416), .Z(n3413) );
  AND U3365 ( .A(n142), .B(n3417), .Z(n3416) );
  XOR U3366 ( .A(n3418), .B(n23), .Z(n94) );
  AND U3367 ( .A(n125), .B(n3419), .Z(n23) );
  XOR U3368 ( .A(n24), .B(n3418), .Z(n3419) );
  XOR U3369 ( .A(n3420), .B(n3421), .Z(n24) );
  AND U3370 ( .A(n130), .B(n3422), .Z(n3421) );
  XOR U3371 ( .A(p_input[22]), .B(n3420), .Z(n3422) );
  XNOR U3372 ( .A(n3423), .B(n3424), .Z(n3420) );
  AND U3373 ( .A(n134), .B(n3425), .Z(n3424) );
  XOR U3374 ( .A(n3426), .B(n3427), .Z(n3418) );
  AND U3375 ( .A(n138), .B(n3417), .Z(n3427) );
  XNOR U3376 ( .A(n3428), .B(n3415), .Z(n3417) );
  XOR U3377 ( .A(n3429), .B(n3430), .Z(n3415) );
  AND U3378 ( .A(n162), .B(n3431), .Z(n3430) );
  IV U3379 ( .A(n3426), .Z(n3428) );
  XOR U3380 ( .A(n3432), .B(n3433), .Z(n3426) );
  AND U3381 ( .A(n146), .B(n3425), .Z(n3433) );
  XNOR U3382 ( .A(n3423), .B(n3432), .Z(n3425) );
  XNOR U3383 ( .A(n3434), .B(n3435), .Z(n3423) );
  AND U3384 ( .A(n150), .B(n3436), .Z(n3435) );
  XOR U3385 ( .A(p_input[54]), .B(n3434), .Z(n3436) );
  XNOR U3386 ( .A(n3437), .B(n3438), .Z(n3434) );
  AND U3387 ( .A(n154), .B(n3439), .Z(n3438) );
  XOR U3388 ( .A(n3440), .B(n3441), .Z(n3432) );
  AND U3389 ( .A(n158), .B(n3431), .Z(n3441) );
  XNOR U3390 ( .A(n3442), .B(n3429), .Z(n3431) );
  XOR U3391 ( .A(n3443), .B(n3444), .Z(n3429) );
  AND U3392 ( .A(n181), .B(n3445), .Z(n3444) );
  IV U3393 ( .A(n3440), .Z(n3442) );
  XOR U3394 ( .A(n3446), .B(n3447), .Z(n3440) );
  AND U3395 ( .A(n165), .B(n3439), .Z(n3447) );
  XNOR U3396 ( .A(n3437), .B(n3446), .Z(n3439) );
  XNOR U3397 ( .A(n3448), .B(n3449), .Z(n3437) );
  AND U3398 ( .A(n169), .B(n3450), .Z(n3449) );
  XOR U3399 ( .A(p_input[86]), .B(n3448), .Z(n3450) );
  XNOR U3400 ( .A(n3451), .B(n3452), .Z(n3448) );
  AND U3401 ( .A(n173), .B(n3453), .Z(n3452) );
  XOR U3402 ( .A(n3454), .B(n3455), .Z(n3446) );
  AND U3403 ( .A(n177), .B(n3445), .Z(n3455) );
  XNOR U3404 ( .A(n3456), .B(n3443), .Z(n3445) );
  XOR U3405 ( .A(n3457), .B(n3458), .Z(n3443) );
  AND U3406 ( .A(n200), .B(n3459), .Z(n3458) );
  IV U3407 ( .A(n3454), .Z(n3456) );
  XOR U3408 ( .A(n3460), .B(n3461), .Z(n3454) );
  AND U3409 ( .A(n184), .B(n3453), .Z(n3461) );
  XNOR U3410 ( .A(n3451), .B(n3460), .Z(n3453) );
  XNOR U3411 ( .A(n3462), .B(n3463), .Z(n3451) );
  AND U3412 ( .A(n188), .B(n3464), .Z(n3463) );
  XOR U3413 ( .A(p_input[118]), .B(n3462), .Z(n3464) );
  XNOR U3414 ( .A(n3465), .B(n3466), .Z(n3462) );
  AND U3415 ( .A(n192), .B(n3467), .Z(n3466) );
  XOR U3416 ( .A(n3468), .B(n3469), .Z(n3460) );
  AND U3417 ( .A(n196), .B(n3459), .Z(n3469) );
  XNOR U3418 ( .A(n3470), .B(n3457), .Z(n3459) );
  XOR U3419 ( .A(n3471), .B(n3472), .Z(n3457) );
  AND U3420 ( .A(n219), .B(n3473), .Z(n3472) );
  IV U3421 ( .A(n3468), .Z(n3470) );
  XOR U3422 ( .A(n3474), .B(n3475), .Z(n3468) );
  AND U3423 ( .A(n203), .B(n3467), .Z(n3475) );
  XNOR U3424 ( .A(n3465), .B(n3474), .Z(n3467) );
  XNOR U3425 ( .A(n3476), .B(n3477), .Z(n3465) );
  AND U3426 ( .A(n207), .B(n3478), .Z(n3477) );
  XOR U3427 ( .A(p_input[150]), .B(n3476), .Z(n3478) );
  XNOR U3428 ( .A(n3479), .B(n3480), .Z(n3476) );
  AND U3429 ( .A(n211), .B(n3481), .Z(n3480) );
  XOR U3430 ( .A(n3482), .B(n3483), .Z(n3474) );
  AND U3431 ( .A(n215), .B(n3473), .Z(n3483) );
  XNOR U3432 ( .A(n3484), .B(n3471), .Z(n3473) );
  XOR U3433 ( .A(n3485), .B(n3486), .Z(n3471) );
  AND U3434 ( .A(n238), .B(n3487), .Z(n3486) );
  IV U3435 ( .A(n3482), .Z(n3484) );
  XOR U3436 ( .A(n3488), .B(n3489), .Z(n3482) );
  AND U3437 ( .A(n222), .B(n3481), .Z(n3489) );
  XNOR U3438 ( .A(n3479), .B(n3488), .Z(n3481) );
  XNOR U3439 ( .A(n3490), .B(n3491), .Z(n3479) );
  AND U3440 ( .A(n226), .B(n3492), .Z(n3491) );
  XOR U3441 ( .A(p_input[182]), .B(n3490), .Z(n3492) );
  XNOR U3442 ( .A(n3493), .B(n3494), .Z(n3490) );
  AND U3443 ( .A(n230), .B(n3495), .Z(n3494) );
  XOR U3444 ( .A(n3496), .B(n3497), .Z(n3488) );
  AND U3445 ( .A(n234), .B(n3487), .Z(n3497) );
  XNOR U3446 ( .A(n3498), .B(n3485), .Z(n3487) );
  XOR U3447 ( .A(n3499), .B(n3500), .Z(n3485) );
  AND U3448 ( .A(n257), .B(n3501), .Z(n3500) );
  IV U3449 ( .A(n3496), .Z(n3498) );
  XOR U3450 ( .A(n3502), .B(n3503), .Z(n3496) );
  AND U3451 ( .A(n241), .B(n3495), .Z(n3503) );
  XNOR U3452 ( .A(n3493), .B(n3502), .Z(n3495) );
  XNOR U3453 ( .A(n3504), .B(n3505), .Z(n3493) );
  AND U3454 ( .A(n245), .B(n3506), .Z(n3505) );
  XOR U3455 ( .A(p_input[214]), .B(n3504), .Z(n3506) );
  XNOR U3456 ( .A(n3507), .B(n3508), .Z(n3504) );
  AND U3457 ( .A(n249), .B(n3509), .Z(n3508) );
  XOR U3458 ( .A(n3510), .B(n3511), .Z(n3502) );
  AND U3459 ( .A(n253), .B(n3501), .Z(n3511) );
  XNOR U3460 ( .A(n3512), .B(n3499), .Z(n3501) );
  XOR U3461 ( .A(n3513), .B(n3514), .Z(n3499) );
  AND U3462 ( .A(n276), .B(n3515), .Z(n3514) );
  IV U3463 ( .A(n3510), .Z(n3512) );
  XOR U3464 ( .A(n3516), .B(n3517), .Z(n3510) );
  AND U3465 ( .A(n260), .B(n3509), .Z(n3517) );
  XNOR U3466 ( .A(n3507), .B(n3516), .Z(n3509) );
  XNOR U3467 ( .A(n3518), .B(n3519), .Z(n3507) );
  AND U3468 ( .A(n264), .B(n3520), .Z(n3519) );
  XOR U3469 ( .A(p_input[246]), .B(n3518), .Z(n3520) );
  XNOR U3470 ( .A(n3521), .B(n3522), .Z(n3518) );
  AND U3471 ( .A(n268), .B(n3523), .Z(n3522) );
  XOR U3472 ( .A(n3524), .B(n3525), .Z(n3516) );
  AND U3473 ( .A(n272), .B(n3515), .Z(n3525) );
  XNOR U3474 ( .A(n3526), .B(n3513), .Z(n3515) );
  XOR U3475 ( .A(n3527), .B(n3528), .Z(n3513) );
  AND U3476 ( .A(n295), .B(n3529), .Z(n3528) );
  IV U3477 ( .A(n3524), .Z(n3526) );
  XOR U3478 ( .A(n3530), .B(n3531), .Z(n3524) );
  AND U3479 ( .A(n279), .B(n3523), .Z(n3531) );
  XNOR U3480 ( .A(n3521), .B(n3530), .Z(n3523) );
  XNOR U3481 ( .A(n3532), .B(n3533), .Z(n3521) );
  AND U3482 ( .A(n283), .B(n3534), .Z(n3533) );
  XOR U3483 ( .A(p_input[278]), .B(n3532), .Z(n3534) );
  XNOR U3484 ( .A(n3535), .B(n3536), .Z(n3532) );
  AND U3485 ( .A(n287), .B(n3537), .Z(n3536) );
  XOR U3486 ( .A(n3538), .B(n3539), .Z(n3530) );
  AND U3487 ( .A(n291), .B(n3529), .Z(n3539) );
  XNOR U3488 ( .A(n3540), .B(n3527), .Z(n3529) );
  XOR U3489 ( .A(n3541), .B(n3542), .Z(n3527) );
  AND U3490 ( .A(n314), .B(n3543), .Z(n3542) );
  IV U3491 ( .A(n3538), .Z(n3540) );
  XOR U3492 ( .A(n3544), .B(n3545), .Z(n3538) );
  AND U3493 ( .A(n298), .B(n3537), .Z(n3545) );
  XNOR U3494 ( .A(n3535), .B(n3544), .Z(n3537) );
  XNOR U3495 ( .A(n3546), .B(n3547), .Z(n3535) );
  AND U3496 ( .A(n302), .B(n3548), .Z(n3547) );
  XOR U3497 ( .A(p_input[310]), .B(n3546), .Z(n3548) );
  XNOR U3498 ( .A(n3549), .B(n3550), .Z(n3546) );
  AND U3499 ( .A(n306), .B(n3551), .Z(n3550) );
  XOR U3500 ( .A(n3552), .B(n3553), .Z(n3544) );
  AND U3501 ( .A(n310), .B(n3543), .Z(n3553) );
  XNOR U3502 ( .A(n3554), .B(n3541), .Z(n3543) );
  XOR U3503 ( .A(n3555), .B(n3556), .Z(n3541) );
  AND U3504 ( .A(n333), .B(n3557), .Z(n3556) );
  IV U3505 ( .A(n3552), .Z(n3554) );
  XOR U3506 ( .A(n3558), .B(n3559), .Z(n3552) );
  AND U3507 ( .A(n317), .B(n3551), .Z(n3559) );
  XNOR U3508 ( .A(n3549), .B(n3558), .Z(n3551) );
  XNOR U3509 ( .A(n3560), .B(n3561), .Z(n3549) );
  AND U3510 ( .A(n321), .B(n3562), .Z(n3561) );
  XOR U3511 ( .A(p_input[342]), .B(n3560), .Z(n3562) );
  XNOR U3512 ( .A(n3563), .B(n3564), .Z(n3560) );
  AND U3513 ( .A(n325), .B(n3565), .Z(n3564) );
  XOR U3514 ( .A(n3566), .B(n3567), .Z(n3558) );
  AND U3515 ( .A(n329), .B(n3557), .Z(n3567) );
  XNOR U3516 ( .A(n3568), .B(n3555), .Z(n3557) );
  XOR U3517 ( .A(n3569), .B(n3570), .Z(n3555) );
  AND U3518 ( .A(n352), .B(n3571), .Z(n3570) );
  IV U3519 ( .A(n3566), .Z(n3568) );
  XOR U3520 ( .A(n3572), .B(n3573), .Z(n3566) );
  AND U3521 ( .A(n336), .B(n3565), .Z(n3573) );
  XNOR U3522 ( .A(n3563), .B(n3572), .Z(n3565) );
  XNOR U3523 ( .A(n3574), .B(n3575), .Z(n3563) );
  AND U3524 ( .A(n340), .B(n3576), .Z(n3575) );
  XOR U3525 ( .A(p_input[374]), .B(n3574), .Z(n3576) );
  XNOR U3526 ( .A(n3577), .B(n3578), .Z(n3574) );
  AND U3527 ( .A(n344), .B(n3579), .Z(n3578) );
  XOR U3528 ( .A(n3580), .B(n3581), .Z(n3572) );
  AND U3529 ( .A(n348), .B(n3571), .Z(n3581) );
  XNOR U3530 ( .A(n3582), .B(n3569), .Z(n3571) );
  XOR U3531 ( .A(n3583), .B(n3584), .Z(n3569) );
  AND U3532 ( .A(n370), .B(n3585), .Z(n3584) );
  IV U3533 ( .A(n3580), .Z(n3582) );
  XOR U3534 ( .A(n3586), .B(n3587), .Z(n3580) );
  AND U3535 ( .A(n355), .B(n3579), .Z(n3587) );
  XNOR U3536 ( .A(n3577), .B(n3586), .Z(n3579) );
  XNOR U3537 ( .A(n3588), .B(n3589), .Z(n3577) );
  AND U3538 ( .A(n359), .B(n3590), .Z(n3589) );
  XOR U3539 ( .A(p_input[406]), .B(n3588), .Z(n3590) );
  XOR U3540 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][22] ), .B(n3591), 
        .Z(n3588) );
  AND U3541 ( .A(n362), .B(n3592), .Z(n3591) );
  XOR U3542 ( .A(n3593), .B(n3594), .Z(n3586) );
  AND U3543 ( .A(n366), .B(n3585), .Z(n3594) );
  XNOR U3544 ( .A(n3595), .B(n3583), .Z(n3585) );
  XOR U3545 ( .A(\knn_comb_/min_val_out[0][22] ), .B(n3596), .Z(n3583) );
  AND U3546 ( .A(n378), .B(n3597), .Z(n3596) );
  IV U3547 ( .A(n3593), .Z(n3595) );
  XOR U3548 ( .A(n3598), .B(n3599), .Z(n3593) );
  AND U3549 ( .A(n373), .B(n3592), .Z(n3599) );
  XOR U3550 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][22] ), .B(n3598), 
        .Z(n3592) );
  XOR U3551 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .B(n3600), 
        .Z(n3598) );
  AND U3552 ( .A(n375), .B(n3597), .Z(n3600) );
  XOR U3553 ( .A(\knn_comb_/min_val_out[0][22] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .Z(n3597) );
  XOR U3554 ( .A(n95), .B(n3601), .Z(o[21]) );
  AND U3555 ( .A(n122), .B(n3602), .Z(n95) );
  XOR U3556 ( .A(n96), .B(n3601), .Z(n3602) );
  XOR U3557 ( .A(n3603), .B(n3604), .Z(n3601) );
  AND U3558 ( .A(n142), .B(n3605), .Z(n3604) );
  XOR U3559 ( .A(n3606), .B(n25), .Z(n96) );
  AND U3560 ( .A(n125), .B(n3607), .Z(n25) );
  XOR U3561 ( .A(n26), .B(n3606), .Z(n3607) );
  XOR U3562 ( .A(n3608), .B(n3609), .Z(n26) );
  AND U3563 ( .A(n130), .B(n3610), .Z(n3609) );
  XOR U3564 ( .A(p_input[21]), .B(n3608), .Z(n3610) );
  XNOR U3565 ( .A(n3611), .B(n3612), .Z(n3608) );
  AND U3566 ( .A(n134), .B(n3613), .Z(n3612) );
  XOR U3567 ( .A(n3614), .B(n3615), .Z(n3606) );
  AND U3568 ( .A(n138), .B(n3605), .Z(n3615) );
  XNOR U3569 ( .A(n3616), .B(n3603), .Z(n3605) );
  XOR U3570 ( .A(n3617), .B(n3618), .Z(n3603) );
  AND U3571 ( .A(n162), .B(n3619), .Z(n3618) );
  IV U3572 ( .A(n3614), .Z(n3616) );
  XOR U3573 ( .A(n3620), .B(n3621), .Z(n3614) );
  AND U3574 ( .A(n146), .B(n3613), .Z(n3621) );
  XNOR U3575 ( .A(n3611), .B(n3620), .Z(n3613) );
  XNOR U3576 ( .A(n3622), .B(n3623), .Z(n3611) );
  AND U3577 ( .A(n150), .B(n3624), .Z(n3623) );
  XOR U3578 ( .A(p_input[53]), .B(n3622), .Z(n3624) );
  XNOR U3579 ( .A(n3625), .B(n3626), .Z(n3622) );
  AND U3580 ( .A(n154), .B(n3627), .Z(n3626) );
  XOR U3581 ( .A(n3628), .B(n3629), .Z(n3620) );
  AND U3582 ( .A(n158), .B(n3619), .Z(n3629) );
  XNOR U3583 ( .A(n3630), .B(n3617), .Z(n3619) );
  XOR U3584 ( .A(n3631), .B(n3632), .Z(n3617) );
  AND U3585 ( .A(n181), .B(n3633), .Z(n3632) );
  IV U3586 ( .A(n3628), .Z(n3630) );
  XOR U3587 ( .A(n3634), .B(n3635), .Z(n3628) );
  AND U3588 ( .A(n165), .B(n3627), .Z(n3635) );
  XNOR U3589 ( .A(n3625), .B(n3634), .Z(n3627) );
  XNOR U3590 ( .A(n3636), .B(n3637), .Z(n3625) );
  AND U3591 ( .A(n169), .B(n3638), .Z(n3637) );
  XOR U3592 ( .A(p_input[85]), .B(n3636), .Z(n3638) );
  XNOR U3593 ( .A(n3639), .B(n3640), .Z(n3636) );
  AND U3594 ( .A(n173), .B(n3641), .Z(n3640) );
  XOR U3595 ( .A(n3642), .B(n3643), .Z(n3634) );
  AND U3596 ( .A(n177), .B(n3633), .Z(n3643) );
  XNOR U3597 ( .A(n3644), .B(n3631), .Z(n3633) );
  XOR U3598 ( .A(n3645), .B(n3646), .Z(n3631) );
  AND U3599 ( .A(n200), .B(n3647), .Z(n3646) );
  IV U3600 ( .A(n3642), .Z(n3644) );
  XOR U3601 ( .A(n3648), .B(n3649), .Z(n3642) );
  AND U3602 ( .A(n184), .B(n3641), .Z(n3649) );
  XNOR U3603 ( .A(n3639), .B(n3648), .Z(n3641) );
  XNOR U3604 ( .A(n3650), .B(n3651), .Z(n3639) );
  AND U3605 ( .A(n188), .B(n3652), .Z(n3651) );
  XOR U3606 ( .A(p_input[117]), .B(n3650), .Z(n3652) );
  XNOR U3607 ( .A(n3653), .B(n3654), .Z(n3650) );
  AND U3608 ( .A(n192), .B(n3655), .Z(n3654) );
  XOR U3609 ( .A(n3656), .B(n3657), .Z(n3648) );
  AND U3610 ( .A(n196), .B(n3647), .Z(n3657) );
  XNOR U3611 ( .A(n3658), .B(n3645), .Z(n3647) );
  XOR U3612 ( .A(n3659), .B(n3660), .Z(n3645) );
  AND U3613 ( .A(n219), .B(n3661), .Z(n3660) );
  IV U3614 ( .A(n3656), .Z(n3658) );
  XOR U3615 ( .A(n3662), .B(n3663), .Z(n3656) );
  AND U3616 ( .A(n203), .B(n3655), .Z(n3663) );
  XNOR U3617 ( .A(n3653), .B(n3662), .Z(n3655) );
  XNOR U3618 ( .A(n3664), .B(n3665), .Z(n3653) );
  AND U3619 ( .A(n207), .B(n3666), .Z(n3665) );
  XOR U3620 ( .A(p_input[149]), .B(n3664), .Z(n3666) );
  XNOR U3621 ( .A(n3667), .B(n3668), .Z(n3664) );
  AND U3622 ( .A(n211), .B(n3669), .Z(n3668) );
  XOR U3623 ( .A(n3670), .B(n3671), .Z(n3662) );
  AND U3624 ( .A(n215), .B(n3661), .Z(n3671) );
  XNOR U3625 ( .A(n3672), .B(n3659), .Z(n3661) );
  XOR U3626 ( .A(n3673), .B(n3674), .Z(n3659) );
  AND U3627 ( .A(n238), .B(n3675), .Z(n3674) );
  IV U3628 ( .A(n3670), .Z(n3672) );
  XOR U3629 ( .A(n3676), .B(n3677), .Z(n3670) );
  AND U3630 ( .A(n222), .B(n3669), .Z(n3677) );
  XNOR U3631 ( .A(n3667), .B(n3676), .Z(n3669) );
  XNOR U3632 ( .A(n3678), .B(n3679), .Z(n3667) );
  AND U3633 ( .A(n226), .B(n3680), .Z(n3679) );
  XOR U3634 ( .A(p_input[181]), .B(n3678), .Z(n3680) );
  XNOR U3635 ( .A(n3681), .B(n3682), .Z(n3678) );
  AND U3636 ( .A(n230), .B(n3683), .Z(n3682) );
  XOR U3637 ( .A(n3684), .B(n3685), .Z(n3676) );
  AND U3638 ( .A(n234), .B(n3675), .Z(n3685) );
  XNOR U3639 ( .A(n3686), .B(n3673), .Z(n3675) );
  XOR U3640 ( .A(n3687), .B(n3688), .Z(n3673) );
  AND U3641 ( .A(n257), .B(n3689), .Z(n3688) );
  IV U3642 ( .A(n3684), .Z(n3686) );
  XOR U3643 ( .A(n3690), .B(n3691), .Z(n3684) );
  AND U3644 ( .A(n241), .B(n3683), .Z(n3691) );
  XNOR U3645 ( .A(n3681), .B(n3690), .Z(n3683) );
  XNOR U3646 ( .A(n3692), .B(n3693), .Z(n3681) );
  AND U3647 ( .A(n245), .B(n3694), .Z(n3693) );
  XOR U3648 ( .A(p_input[213]), .B(n3692), .Z(n3694) );
  XNOR U3649 ( .A(n3695), .B(n3696), .Z(n3692) );
  AND U3650 ( .A(n249), .B(n3697), .Z(n3696) );
  XOR U3651 ( .A(n3698), .B(n3699), .Z(n3690) );
  AND U3652 ( .A(n253), .B(n3689), .Z(n3699) );
  XNOR U3653 ( .A(n3700), .B(n3687), .Z(n3689) );
  XOR U3654 ( .A(n3701), .B(n3702), .Z(n3687) );
  AND U3655 ( .A(n276), .B(n3703), .Z(n3702) );
  IV U3656 ( .A(n3698), .Z(n3700) );
  XOR U3657 ( .A(n3704), .B(n3705), .Z(n3698) );
  AND U3658 ( .A(n260), .B(n3697), .Z(n3705) );
  XNOR U3659 ( .A(n3695), .B(n3704), .Z(n3697) );
  XNOR U3660 ( .A(n3706), .B(n3707), .Z(n3695) );
  AND U3661 ( .A(n264), .B(n3708), .Z(n3707) );
  XOR U3662 ( .A(p_input[245]), .B(n3706), .Z(n3708) );
  XNOR U3663 ( .A(n3709), .B(n3710), .Z(n3706) );
  AND U3664 ( .A(n268), .B(n3711), .Z(n3710) );
  XOR U3665 ( .A(n3712), .B(n3713), .Z(n3704) );
  AND U3666 ( .A(n272), .B(n3703), .Z(n3713) );
  XNOR U3667 ( .A(n3714), .B(n3701), .Z(n3703) );
  XOR U3668 ( .A(n3715), .B(n3716), .Z(n3701) );
  AND U3669 ( .A(n295), .B(n3717), .Z(n3716) );
  IV U3670 ( .A(n3712), .Z(n3714) );
  XOR U3671 ( .A(n3718), .B(n3719), .Z(n3712) );
  AND U3672 ( .A(n279), .B(n3711), .Z(n3719) );
  XNOR U3673 ( .A(n3709), .B(n3718), .Z(n3711) );
  XNOR U3674 ( .A(n3720), .B(n3721), .Z(n3709) );
  AND U3675 ( .A(n283), .B(n3722), .Z(n3721) );
  XOR U3676 ( .A(p_input[277]), .B(n3720), .Z(n3722) );
  XNOR U3677 ( .A(n3723), .B(n3724), .Z(n3720) );
  AND U3678 ( .A(n287), .B(n3725), .Z(n3724) );
  XOR U3679 ( .A(n3726), .B(n3727), .Z(n3718) );
  AND U3680 ( .A(n291), .B(n3717), .Z(n3727) );
  XNOR U3681 ( .A(n3728), .B(n3715), .Z(n3717) );
  XOR U3682 ( .A(n3729), .B(n3730), .Z(n3715) );
  AND U3683 ( .A(n314), .B(n3731), .Z(n3730) );
  IV U3684 ( .A(n3726), .Z(n3728) );
  XOR U3685 ( .A(n3732), .B(n3733), .Z(n3726) );
  AND U3686 ( .A(n298), .B(n3725), .Z(n3733) );
  XNOR U3687 ( .A(n3723), .B(n3732), .Z(n3725) );
  XNOR U3688 ( .A(n3734), .B(n3735), .Z(n3723) );
  AND U3689 ( .A(n302), .B(n3736), .Z(n3735) );
  XOR U3690 ( .A(p_input[309]), .B(n3734), .Z(n3736) );
  XNOR U3691 ( .A(n3737), .B(n3738), .Z(n3734) );
  AND U3692 ( .A(n306), .B(n3739), .Z(n3738) );
  XOR U3693 ( .A(n3740), .B(n3741), .Z(n3732) );
  AND U3694 ( .A(n310), .B(n3731), .Z(n3741) );
  XNOR U3695 ( .A(n3742), .B(n3729), .Z(n3731) );
  XOR U3696 ( .A(n3743), .B(n3744), .Z(n3729) );
  AND U3697 ( .A(n333), .B(n3745), .Z(n3744) );
  IV U3698 ( .A(n3740), .Z(n3742) );
  XOR U3699 ( .A(n3746), .B(n3747), .Z(n3740) );
  AND U3700 ( .A(n317), .B(n3739), .Z(n3747) );
  XNOR U3701 ( .A(n3737), .B(n3746), .Z(n3739) );
  XNOR U3702 ( .A(n3748), .B(n3749), .Z(n3737) );
  AND U3703 ( .A(n321), .B(n3750), .Z(n3749) );
  XOR U3704 ( .A(p_input[341]), .B(n3748), .Z(n3750) );
  XNOR U3705 ( .A(n3751), .B(n3752), .Z(n3748) );
  AND U3706 ( .A(n325), .B(n3753), .Z(n3752) );
  XOR U3707 ( .A(n3754), .B(n3755), .Z(n3746) );
  AND U3708 ( .A(n329), .B(n3745), .Z(n3755) );
  XNOR U3709 ( .A(n3756), .B(n3743), .Z(n3745) );
  XOR U3710 ( .A(n3757), .B(n3758), .Z(n3743) );
  AND U3711 ( .A(n352), .B(n3759), .Z(n3758) );
  IV U3712 ( .A(n3754), .Z(n3756) );
  XOR U3713 ( .A(n3760), .B(n3761), .Z(n3754) );
  AND U3714 ( .A(n336), .B(n3753), .Z(n3761) );
  XNOR U3715 ( .A(n3751), .B(n3760), .Z(n3753) );
  XNOR U3716 ( .A(n3762), .B(n3763), .Z(n3751) );
  AND U3717 ( .A(n340), .B(n3764), .Z(n3763) );
  XOR U3718 ( .A(p_input[373]), .B(n3762), .Z(n3764) );
  XNOR U3719 ( .A(n3765), .B(n3766), .Z(n3762) );
  AND U3720 ( .A(n344), .B(n3767), .Z(n3766) );
  XOR U3721 ( .A(n3768), .B(n3769), .Z(n3760) );
  AND U3722 ( .A(n348), .B(n3759), .Z(n3769) );
  XNOR U3723 ( .A(n3770), .B(n3757), .Z(n3759) );
  XOR U3724 ( .A(n3771), .B(n3772), .Z(n3757) );
  AND U3725 ( .A(n370), .B(n3773), .Z(n3772) );
  IV U3726 ( .A(n3768), .Z(n3770) );
  XOR U3727 ( .A(n3774), .B(n3775), .Z(n3768) );
  AND U3728 ( .A(n355), .B(n3767), .Z(n3775) );
  XNOR U3729 ( .A(n3765), .B(n3774), .Z(n3767) );
  XNOR U3730 ( .A(n3776), .B(n3777), .Z(n3765) );
  AND U3731 ( .A(n359), .B(n3778), .Z(n3777) );
  XOR U3732 ( .A(p_input[405]), .B(n3776), .Z(n3778) );
  XOR U3733 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][21] ), .B(n3779), 
        .Z(n3776) );
  AND U3734 ( .A(n362), .B(n3780), .Z(n3779) );
  XOR U3735 ( .A(n3781), .B(n3782), .Z(n3774) );
  AND U3736 ( .A(n366), .B(n3773), .Z(n3782) );
  XNOR U3737 ( .A(n3783), .B(n3771), .Z(n3773) );
  XOR U3738 ( .A(\knn_comb_/min_val_out[0][21] ), .B(n3784), .Z(n3771) );
  AND U3739 ( .A(n378), .B(n3785), .Z(n3784) );
  IV U3740 ( .A(n3781), .Z(n3783) );
  XOR U3741 ( .A(n3786), .B(n3787), .Z(n3781) );
  AND U3742 ( .A(n373), .B(n3780), .Z(n3787) );
  XOR U3743 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][21] ), .B(n3786), 
        .Z(n3780) );
  XOR U3744 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .B(n3788), 
        .Z(n3786) );
  AND U3745 ( .A(n375), .B(n3785), .Z(n3788) );
  XOR U3746 ( .A(\knn_comb_/min_val_out[0][21] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .Z(n3785) );
  XOR U3747 ( .A(n97), .B(n3789), .Z(o[20]) );
  AND U3748 ( .A(n122), .B(n3790), .Z(n97) );
  XOR U3749 ( .A(n98), .B(n3789), .Z(n3790) );
  XOR U3750 ( .A(n3791), .B(n3792), .Z(n3789) );
  AND U3751 ( .A(n142), .B(n3793), .Z(n3792) );
  XOR U3752 ( .A(n3794), .B(n27), .Z(n98) );
  AND U3753 ( .A(n125), .B(n3795), .Z(n27) );
  XOR U3754 ( .A(n28), .B(n3794), .Z(n3795) );
  XOR U3755 ( .A(n3796), .B(n3797), .Z(n28) );
  AND U3756 ( .A(n130), .B(n3798), .Z(n3797) );
  XOR U3757 ( .A(p_input[20]), .B(n3796), .Z(n3798) );
  XNOR U3758 ( .A(n3799), .B(n3800), .Z(n3796) );
  AND U3759 ( .A(n134), .B(n3801), .Z(n3800) );
  XOR U3760 ( .A(n3802), .B(n3803), .Z(n3794) );
  AND U3761 ( .A(n138), .B(n3793), .Z(n3803) );
  XNOR U3762 ( .A(n3804), .B(n3791), .Z(n3793) );
  XOR U3763 ( .A(n3805), .B(n3806), .Z(n3791) );
  AND U3764 ( .A(n162), .B(n3807), .Z(n3806) );
  IV U3765 ( .A(n3802), .Z(n3804) );
  XOR U3766 ( .A(n3808), .B(n3809), .Z(n3802) );
  AND U3767 ( .A(n146), .B(n3801), .Z(n3809) );
  XNOR U3768 ( .A(n3799), .B(n3808), .Z(n3801) );
  XNOR U3769 ( .A(n3810), .B(n3811), .Z(n3799) );
  AND U3770 ( .A(n150), .B(n3812), .Z(n3811) );
  XOR U3771 ( .A(p_input[52]), .B(n3810), .Z(n3812) );
  XNOR U3772 ( .A(n3813), .B(n3814), .Z(n3810) );
  AND U3773 ( .A(n154), .B(n3815), .Z(n3814) );
  XOR U3774 ( .A(n3816), .B(n3817), .Z(n3808) );
  AND U3775 ( .A(n158), .B(n3807), .Z(n3817) );
  XNOR U3776 ( .A(n3818), .B(n3805), .Z(n3807) );
  XOR U3777 ( .A(n3819), .B(n3820), .Z(n3805) );
  AND U3778 ( .A(n181), .B(n3821), .Z(n3820) );
  IV U3779 ( .A(n3816), .Z(n3818) );
  XOR U3780 ( .A(n3822), .B(n3823), .Z(n3816) );
  AND U3781 ( .A(n165), .B(n3815), .Z(n3823) );
  XNOR U3782 ( .A(n3813), .B(n3822), .Z(n3815) );
  XNOR U3783 ( .A(n3824), .B(n3825), .Z(n3813) );
  AND U3784 ( .A(n169), .B(n3826), .Z(n3825) );
  XOR U3785 ( .A(p_input[84]), .B(n3824), .Z(n3826) );
  XNOR U3786 ( .A(n3827), .B(n3828), .Z(n3824) );
  AND U3787 ( .A(n173), .B(n3829), .Z(n3828) );
  XOR U3788 ( .A(n3830), .B(n3831), .Z(n3822) );
  AND U3789 ( .A(n177), .B(n3821), .Z(n3831) );
  XNOR U3790 ( .A(n3832), .B(n3819), .Z(n3821) );
  XOR U3791 ( .A(n3833), .B(n3834), .Z(n3819) );
  AND U3792 ( .A(n200), .B(n3835), .Z(n3834) );
  IV U3793 ( .A(n3830), .Z(n3832) );
  XOR U3794 ( .A(n3836), .B(n3837), .Z(n3830) );
  AND U3795 ( .A(n184), .B(n3829), .Z(n3837) );
  XNOR U3796 ( .A(n3827), .B(n3836), .Z(n3829) );
  XNOR U3797 ( .A(n3838), .B(n3839), .Z(n3827) );
  AND U3798 ( .A(n188), .B(n3840), .Z(n3839) );
  XOR U3799 ( .A(p_input[116]), .B(n3838), .Z(n3840) );
  XNOR U3800 ( .A(n3841), .B(n3842), .Z(n3838) );
  AND U3801 ( .A(n192), .B(n3843), .Z(n3842) );
  XOR U3802 ( .A(n3844), .B(n3845), .Z(n3836) );
  AND U3803 ( .A(n196), .B(n3835), .Z(n3845) );
  XNOR U3804 ( .A(n3846), .B(n3833), .Z(n3835) );
  XOR U3805 ( .A(n3847), .B(n3848), .Z(n3833) );
  AND U3806 ( .A(n219), .B(n3849), .Z(n3848) );
  IV U3807 ( .A(n3844), .Z(n3846) );
  XOR U3808 ( .A(n3850), .B(n3851), .Z(n3844) );
  AND U3809 ( .A(n203), .B(n3843), .Z(n3851) );
  XNOR U3810 ( .A(n3841), .B(n3850), .Z(n3843) );
  XNOR U3811 ( .A(n3852), .B(n3853), .Z(n3841) );
  AND U3812 ( .A(n207), .B(n3854), .Z(n3853) );
  XOR U3813 ( .A(p_input[148]), .B(n3852), .Z(n3854) );
  XNOR U3814 ( .A(n3855), .B(n3856), .Z(n3852) );
  AND U3815 ( .A(n211), .B(n3857), .Z(n3856) );
  XOR U3816 ( .A(n3858), .B(n3859), .Z(n3850) );
  AND U3817 ( .A(n215), .B(n3849), .Z(n3859) );
  XNOR U3818 ( .A(n3860), .B(n3847), .Z(n3849) );
  XOR U3819 ( .A(n3861), .B(n3862), .Z(n3847) );
  AND U3820 ( .A(n238), .B(n3863), .Z(n3862) );
  IV U3821 ( .A(n3858), .Z(n3860) );
  XOR U3822 ( .A(n3864), .B(n3865), .Z(n3858) );
  AND U3823 ( .A(n222), .B(n3857), .Z(n3865) );
  XNOR U3824 ( .A(n3855), .B(n3864), .Z(n3857) );
  XNOR U3825 ( .A(n3866), .B(n3867), .Z(n3855) );
  AND U3826 ( .A(n226), .B(n3868), .Z(n3867) );
  XOR U3827 ( .A(p_input[180]), .B(n3866), .Z(n3868) );
  XNOR U3828 ( .A(n3869), .B(n3870), .Z(n3866) );
  AND U3829 ( .A(n230), .B(n3871), .Z(n3870) );
  XOR U3830 ( .A(n3872), .B(n3873), .Z(n3864) );
  AND U3831 ( .A(n234), .B(n3863), .Z(n3873) );
  XNOR U3832 ( .A(n3874), .B(n3861), .Z(n3863) );
  XOR U3833 ( .A(n3875), .B(n3876), .Z(n3861) );
  AND U3834 ( .A(n257), .B(n3877), .Z(n3876) );
  IV U3835 ( .A(n3872), .Z(n3874) );
  XOR U3836 ( .A(n3878), .B(n3879), .Z(n3872) );
  AND U3837 ( .A(n241), .B(n3871), .Z(n3879) );
  XNOR U3838 ( .A(n3869), .B(n3878), .Z(n3871) );
  XNOR U3839 ( .A(n3880), .B(n3881), .Z(n3869) );
  AND U3840 ( .A(n245), .B(n3882), .Z(n3881) );
  XOR U3841 ( .A(p_input[212]), .B(n3880), .Z(n3882) );
  XNOR U3842 ( .A(n3883), .B(n3884), .Z(n3880) );
  AND U3843 ( .A(n249), .B(n3885), .Z(n3884) );
  XOR U3844 ( .A(n3886), .B(n3887), .Z(n3878) );
  AND U3845 ( .A(n253), .B(n3877), .Z(n3887) );
  XNOR U3846 ( .A(n3888), .B(n3875), .Z(n3877) );
  XOR U3847 ( .A(n3889), .B(n3890), .Z(n3875) );
  AND U3848 ( .A(n276), .B(n3891), .Z(n3890) );
  IV U3849 ( .A(n3886), .Z(n3888) );
  XOR U3850 ( .A(n3892), .B(n3893), .Z(n3886) );
  AND U3851 ( .A(n260), .B(n3885), .Z(n3893) );
  XNOR U3852 ( .A(n3883), .B(n3892), .Z(n3885) );
  XNOR U3853 ( .A(n3894), .B(n3895), .Z(n3883) );
  AND U3854 ( .A(n264), .B(n3896), .Z(n3895) );
  XOR U3855 ( .A(p_input[244]), .B(n3894), .Z(n3896) );
  XNOR U3856 ( .A(n3897), .B(n3898), .Z(n3894) );
  AND U3857 ( .A(n268), .B(n3899), .Z(n3898) );
  XOR U3858 ( .A(n3900), .B(n3901), .Z(n3892) );
  AND U3859 ( .A(n272), .B(n3891), .Z(n3901) );
  XNOR U3860 ( .A(n3902), .B(n3889), .Z(n3891) );
  XOR U3861 ( .A(n3903), .B(n3904), .Z(n3889) );
  AND U3862 ( .A(n295), .B(n3905), .Z(n3904) );
  IV U3863 ( .A(n3900), .Z(n3902) );
  XOR U3864 ( .A(n3906), .B(n3907), .Z(n3900) );
  AND U3865 ( .A(n279), .B(n3899), .Z(n3907) );
  XNOR U3866 ( .A(n3897), .B(n3906), .Z(n3899) );
  XNOR U3867 ( .A(n3908), .B(n3909), .Z(n3897) );
  AND U3868 ( .A(n283), .B(n3910), .Z(n3909) );
  XOR U3869 ( .A(p_input[276]), .B(n3908), .Z(n3910) );
  XNOR U3870 ( .A(n3911), .B(n3912), .Z(n3908) );
  AND U3871 ( .A(n287), .B(n3913), .Z(n3912) );
  XOR U3872 ( .A(n3914), .B(n3915), .Z(n3906) );
  AND U3873 ( .A(n291), .B(n3905), .Z(n3915) );
  XNOR U3874 ( .A(n3916), .B(n3903), .Z(n3905) );
  XOR U3875 ( .A(n3917), .B(n3918), .Z(n3903) );
  AND U3876 ( .A(n314), .B(n3919), .Z(n3918) );
  IV U3877 ( .A(n3914), .Z(n3916) );
  XOR U3878 ( .A(n3920), .B(n3921), .Z(n3914) );
  AND U3879 ( .A(n298), .B(n3913), .Z(n3921) );
  XNOR U3880 ( .A(n3911), .B(n3920), .Z(n3913) );
  XNOR U3881 ( .A(n3922), .B(n3923), .Z(n3911) );
  AND U3882 ( .A(n302), .B(n3924), .Z(n3923) );
  XOR U3883 ( .A(p_input[308]), .B(n3922), .Z(n3924) );
  XNOR U3884 ( .A(n3925), .B(n3926), .Z(n3922) );
  AND U3885 ( .A(n306), .B(n3927), .Z(n3926) );
  XOR U3886 ( .A(n3928), .B(n3929), .Z(n3920) );
  AND U3887 ( .A(n310), .B(n3919), .Z(n3929) );
  XNOR U3888 ( .A(n3930), .B(n3917), .Z(n3919) );
  XOR U3889 ( .A(n3931), .B(n3932), .Z(n3917) );
  AND U3890 ( .A(n333), .B(n3933), .Z(n3932) );
  IV U3891 ( .A(n3928), .Z(n3930) );
  XOR U3892 ( .A(n3934), .B(n3935), .Z(n3928) );
  AND U3893 ( .A(n317), .B(n3927), .Z(n3935) );
  XNOR U3894 ( .A(n3925), .B(n3934), .Z(n3927) );
  XNOR U3895 ( .A(n3936), .B(n3937), .Z(n3925) );
  AND U3896 ( .A(n321), .B(n3938), .Z(n3937) );
  XOR U3897 ( .A(p_input[340]), .B(n3936), .Z(n3938) );
  XNOR U3898 ( .A(n3939), .B(n3940), .Z(n3936) );
  AND U3899 ( .A(n325), .B(n3941), .Z(n3940) );
  XOR U3900 ( .A(n3942), .B(n3943), .Z(n3934) );
  AND U3901 ( .A(n329), .B(n3933), .Z(n3943) );
  XNOR U3902 ( .A(n3944), .B(n3931), .Z(n3933) );
  XOR U3903 ( .A(n3945), .B(n3946), .Z(n3931) );
  AND U3904 ( .A(n352), .B(n3947), .Z(n3946) );
  IV U3905 ( .A(n3942), .Z(n3944) );
  XOR U3906 ( .A(n3948), .B(n3949), .Z(n3942) );
  AND U3907 ( .A(n336), .B(n3941), .Z(n3949) );
  XNOR U3908 ( .A(n3939), .B(n3948), .Z(n3941) );
  XNOR U3909 ( .A(n3950), .B(n3951), .Z(n3939) );
  AND U3910 ( .A(n340), .B(n3952), .Z(n3951) );
  XOR U3911 ( .A(p_input[372]), .B(n3950), .Z(n3952) );
  XNOR U3912 ( .A(n3953), .B(n3954), .Z(n3950) );
  AND U3913 ( .A(n344), .B(n3955), .Z(n3954) );
  XOR U3914 ( .A(n3956), .B(n3957), .Z(n3948) );
  AND U3915 ( .A(n348), .B(n3947), .Z(n3957) );
  XNOR U3916 ( .A(n3958), .B(n3945), .Z(n3947) );
  XOR U3917 ( .A(n3959), .B(n3960), .Z(n3945) );
  AND U3918 ( .A(n370), .B(n3961), .Z(n3960) );
  IV U3919 ( .A(n3956), .Z(n3958) );
  XOR U3920 ( .A(n3962), .B(n3963), .Z(n3956) );
  AND U3921 ( .A(n355), .B(n3955), .Z(n3963) );
  XNOR U3922 ( .A(n3953), .B(n3962), .Z(n3955) );
  XNOR U3923 ( .A(n3964), .B(n3965), .Z(n3953) );
  AND U3924 ( .A(n359), .B(n3966), .Z(n3965) );
  XOR U3925 ( .A(p_input[404]), .B(n3964), .Z(n3966) );
  XOR U3926 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][20] ), .B(n3967), 
        .Z(n3964) );
  AND U3927 ( .A(n362), .B(n3968), .Z(n3967) );
  XOR U3928 ( .A(n3969), .B(n3970), .Z(n3962) );
  AND U3929 ( .A(n366), .B(n3961), .Z(n3970) );
  XNOR U3930 ( .A(n3971), .B(n3959), .Z(n3961) );
  XOR U3931 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n3972), .Z(n3959) );
  AND U3932 ( .A(n378), .B(n3973), .Z(n3972) );
  IV U3933 ( .A(n3969), .Z(n3971) );
  XOR U3934 ( .A(n3974), .B(n3975), .Z(n3969) );
  AND U3935 ( .A(n373), .B(n3968), .Z(n3975) );
  XOR U3936 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][20] ), .B(n3974), 
        .Z(n3968) );
  XOR U3937 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .B(n3976), 
        .Z(n3974) );
  AND U3938 ( .A(n375), .B(n3973), .Z(n3976) );
  XOR U3939 ( .A(n3977), .B(n3978), .Z(n3973) );
  IV U3940 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .Z(n3978) );
  IV U3941 ( .A(\knn_comb_/min_val_out[0][20] ), .Z(n3977) );
  XOR U3942 ( .A(n1521), .B(n3979), .Z(o[1]) );
  AND U3943 ( .A(n122), .B(n3980), .Z(n1521) );
  XOR U3944 ( .A(n1522), .B(n3979), .Z(n3980) );
  XOR U3945 ( .A(n3981), .B(n3982), .Z(n3979) );
  AND U3946 ( .A(n142), .B(n3983), .Z(n3982) );
  XOR U3947 ( .A(n3984), .B(n69), .Z(n1522) );
  AND U3948 ( .A(n125), .B(n3985), .Z(n69) );
  XOR U3949 ( .A(n70), .B(n3984), .Z(n3985) );
  XOR U3950 ( .A(n3986), .B(n3987), .Z(n70) );
  AND U3951 ( .A(n130), .B(n3988), .Z(n3987) );
  XOR U3952 ( .A(p_input[1]), .B(n3986), .Z(n3988) );
  XNOR U3953 ( .A(n3989), .B(n3990), .Z(n3986) );
  AND U3954 ( .A(n134), .B(n3991), .Z(n3990) );
  XOR U3955 ( .A(n3992), .B(n3993), .Z(n3984) );
  AND U3956 ( .A(n138), .B(n3983), .Z(n3993) );
  XNOR U3957 ( .A(n3994), .B(n3981), .Z(n3983) );
  XOR U3958 ( .A(n3995), .B(n3996), .Z(n3981) );
  AND U3959 ( .A(n162), .B(n3997), .Z(n3996) );
  IV U3960 ( .A(n3992), .Z(n3994) );
  XOR U3961 ( .A(n3998), .B(n3999), .Z(n3992) );
  AND U3962 ( .A(n146), .B(n3991), .Z(n3999) );
  XNOR U3963 ( .A(n3989), .B(n3998), .Z(n3991) );
  XNOR U3964 ( .A(n4000), .B(n4001), .Z(n3989) );
  AND U3965 ( .A(n150), .B(n4002), .Z(n4001) );
  XOR U3966 ( .A(p_input[33]), .B(n4000), .Z(n4002) );
  XNOR U3967 ( .A(n4003), .B(n4004), .Z(n4000) );
  AND U3968 ( .A(n154), .B(n4005), .Z(n4004) );
  XOR U3969 ( .A(n4006), .B(n4007), .Z(n3998) );
  AND U3970 ( .A(n158), .B(n3997), .Z(n4007) );
  XNOR U3971 ( .A(n4008), .B(n3995), .Z(n3997) );
  XOR U3972 ( .A(n4009), .B(n4010), .Z(n3995) );
  AND U3973 ( .A(n181), .B(n4011), .Z(n4010) );
  IV U3974 ( .A(n4006), .Z(n4008) );
  XOR U3975 ( .A(n4012), .B(n4013), .Z(n4006) );
  AND U3976 ( .A(n165), .B(n4005), .Z(n4013) );
  XNOR U3977 ( .A(n4003), .B(n4012), .Z(n4005) );
  XNOR U3978 ( .A(n4014), .B(n4015), .Z(n4003) );
  AND U3979 ( .A(n169), .B(n4016), .Z(n4015) );
  XOR U3980 ( .A(p_input[65]), .B(n4014), .Z(n4016) );
  XNOR U3981 ( .A(n4017), .B(n4018), .Z(n4014) );
  AND U3982 ( .A(n173), .B(n4019), .Z(n4018) );
  XOR U3983 ( .A(n4020), .B(n4021), .Z(n4012) );
  AND U3984 ( .A(n177), .B(n4011), .Z(n4021) );
  XNOR U3985 ( .A(n4022), .B(n4009), .Z(n4011) );
  XOR U3986 ( .A(n4023), .B(n4024), .Z(n4009) );
  AND U3987 ( .A(n200), .B(n4025), .Z(n4024) );
  IV U3988 ( .A(n4020), .Z(n4022) );
  XOR U3989 ( .A(n4026), .B(n4027), .Z(n4020) );
  AND U3990 ( .A(n184), .B(n4019), .Z(n4027) );
  XNOR U3991 ( .A(n4017), .B(n4026), .Z(n4019) );
  XNOR U3992 ( .A(n4028), .B(n4029), .Z(n4017) );
  AND U3993 ( .A(n188), .B(n4030), .Z(n4029) );
  XOR U3994 ( .A(p_input[97]), .B(n4028), .Z(n4030) );
  XNOR U3995 ( .A(n4031), .B(n4032), .Z(n4028) );
  AND U3996 ( .A(n192), .B(n4033), .Z(n4032) );
  XOR U3997 ( .A(n4034), .B(n4035), .Z(n4026) );
  AND U3998 ( .A(n196), .B(n4025), .Z(n4035) );
  XNOR U3999 ( .A(n4036), .B(n4023), .Z(n4025) );
  XOR U4000 ( .A(n4037), .B(n4038), .Z(n4023) );
  AND U4001 ( .A(n219), .B(n4039), .Z(n4038) );
  IV U4002 ( .A(n4034), .Z(n4036) );
  XOR U4003 ( .A(n4040), .B(n4041), .Z(n4034) );
  AND U4004 ( .A(n203), .B(n4033), .Z(n4041) );
  XNOR U4005 ( .A(n4031), .B(n4040), .Z(n4033) );
  XNOR U4006 ( .A(n4042), .B(n4043), .Z(n4031) );
  AND U4007 ( .A(n207), .B(n4044), .Z(n4043) );
  XOR U4008 ( .A(p_input[129]), .B(n4042), .Z(n4044) );
  XNOR U4009 ( .A(n4045), .B(n4046), .Z(n4042) );
  AND U4010 ( .A(n211), .B(n4047), .Z(n4046) );
  XOR U4011 ( .A(n4048), .B(n4049), .Z(n4040) );
  AND U4012 ( .A(n215), .B(n4039), .Z(n4049) );
  XNOR U4013 ( .A(n4050), .B(n4037), .Z(n4039) );
  XOR U4014 ( .A(n4051), .B(n4052), .Z(n4037) );
  AND U4015 ( .A(n238), .B(n4053), .Z(n4052) );
  IV U4016 ( .A(n4048), .Z(n4050) );
  XOR U4017 ( .A(n4054), .B(n4055), .Z(n4048) );
  AND U4018 ( .A(n222), .B(n4047), .Z(n4055) );
  XNOR U4019 ( .A(n4045), .B(n4054), .Z(n4047) );
  XNOR U4020 ( .A(n4056), .B(n4057), .Z(n4045) );
  AND U4021 ( .A(n226), .B(n4058), .Z(n4057) );
  XOR U4022 ( .A(p_input[161]), .B(n4056), .Z(n4058) );
  XNOR U4023 ( .A(n4059), .B(n4060), .Z(n4056) );
  AND U4024 ( .A(n230), .B(n4061), .Z(n4060) );
  XOR U4025 ( .A(n4062), .B(n4063), .Z(n4054) );
  AND U4026 ( .A(n234), .B(n4053), .Z(n4063) );
  XNOR U4027 ( .A(n4064), .B(n4051), .Z(n4053) );
  XOR U4028 ( .A(n4065), .B(n4066), .Z(n4051) );
  AND U4029 ( .A(n257), .B(n4067), .Z(n4066) );
  IV U4030 ( .A(n4062), .Z(n4064) );
  XOR U4031 ( .A(n4068), .B(n4069), .Z(n4062) );
  AND U4032 ( .A(n241), .B(n4061), .Z(n4069) );
  XNOR U4033 ( .A(n4059), .B(n4068), .Z(n4061) );
  XNOR U4034 ( .A(n4070), .B(n4071), .Z(n4059) );
  AND U4035 ( .A(n245), .B(n4072), .Z(n4071) );
  XOR U4036 ( .A(p_input[193]), .B(n4070), .Z(n4072) );
  XNOR U4037 ( .A(n4073), .B(n4074), .Z(n4070) );
  AND U4038 ( .A(n249), .B(n4075), .Z(n4074) );
  XOR U4039 ( .A(n4076), .B(n4077), .Z(n4068) );
  AND U4040 ( .A(n253), .B(n4067), .Z(n4077) );
  XNOR U4041 ( .A(n4078), .B(n4065), .Z(n4067) );
  XOR U4042 ( .A(n4079), .B(n4080), .Z(n4065) );
  AND U4043 ( .A(n276), .B(n4081), .Z(n4080) );
  IV U4044 ( .A(n4076), .Z(n4078) );
  XOR U4045 ( .A(n4082), .B(n4083), .Z(n4076) );
  AND U4046 ( .A(n260), .B(n4075), .Z(n4083) );
  XNOR U4047 ( .A(n4073), .B(n4082), .Z(n4075) );
  XNOR U4048 ( .A(n4084), .B(n4085), .Z(n4073) );
  AND U4049 ( .A(n264), .B(n4086), .Z(n4085) );
  XOR U4050 ( .A(p_input[225]), .B(n4084), .Z(n4086) );
  XNOR U4051 ( .A(n4087), .B(n4088), .Z(n4084) );
  AND U4052 ( .A(n268), .B(n4089), .Z(n4088) );
  XOR U4053 ( .A(n4090), .B(n4091), .Z(n4082) );
  AND U4054 ( .A(n272), .B(n4081), .Z(n4091) );
  XNOR U4055 ( .A(n4092), .B(n4079), .Z(n4081) );
  XOR U4056 ( .A(n4093), .B(n4094), .Z(n4079) );
  AND U4057 ( .A(n295), .B(n4095), .Z(n4094) );
  IV U4058 ( .A(n4090), .Z(n4092) );
  XOR U4059 ( .A(n4096), .B(n4097), .Z(n4090) );
  AND U4060 ( .A(n279), .B(n4089), .Z(n4097) );
  XNOR U4061 ( .A(n4087), .B(n4096), .Z(n4089) );
  XNOR U4062 ( .A(n4098), .B(n4099), .Z(n4087) );
  AND U4063 ( .A(n283), .B(n4100), .Z(n4099) );
  XOR U4064 ( .A(p_input[257]), .B(n4098), .Z(n4100) );
  XNOR U4065 ( .A(n4101), .B(n4102), .Z(n4098) );
  AND U4066 ( .A(n287), .B(n4103), .Z(n4102) );
  XOR U4067 ( .A(n4104), .B(n4105), .Z(n4096) );
  AND U4068 ( .A(n291), .B(n4095), .Z(n4105) );
  XNOR U4069 ( .A(n4106), .B(n4093), .Z(n4095) );
  XOR U4070 ( .A(n4107), .B(n4108), .Z(n4093) );
  AND U4071 ( .A(n314), .B(n4109), .Z(n4108) );
  IV U4072 ( .A(n4104), .Z(n4106) );
  XOR U4073 ( .A(n4110), .B(n4111), .Z(n4104) );
  AND U4074 ( .A(n298), .B(n4103), .Z(n4111) );
  XNOR U4075 ( .A(n4101), .B(n4110), .Z(n4103) );
  XNOR U4076 ( .A(n4112), .B(n4113), .Z(n4101) );
  AND U4077 ( .A(n302), .B(n4114), .Z(n4113) );
  XOR U4078 ( .A(p_input[289]), .B(n4112), .Z(n4114) );
  XNOR U4079 ( .A(n4115), .B(n4116), .Z(n4112) );
  AND U4080 ( .A(n306), .B(n4117), .Z(n4116) );
  XOR U4081 ( .A(n4118), .B(n4119), .Z(n4110) );
  AND U4082 ( .A(n310), .B(n4109), .Z(n4119) );
  XNOR U4083 ( .A(n4120), .B(n4107), .Z(n4109) );
  XOR U4084 ( .A(n4121), .B(n4122), .Z(n4107) );
  AND U4085 ( .A(n333), .B(n4123), .Z(n4122) );
  IV U4086 ( .A(n4118), .Z(n4120) );
  XOR U4087 ( .A(n4124), .B(n4125), .Z(n4118) );
  AND U4088 ( .A(n317), .B(n4117), .Z(n4125) );
  XNOR U4089 ( .A(n4115), .B(n4124), .Z(n4117) );
  XNOR U4090 ( .A(n4126), .B(n4127), .Z(n4115) );
  AND U4091 ( .A(n321), .B(n4128), .Z(n4127) );
  XOR U4092 ( .A(p_input[321]), .B(n4126), .Z(n4128) );
  XNOR U4093 ( .A(n4129), .B(n4130), .Z(n4126) );
  AND U4094 ( .A(n325), .B(n4131), .Z(n4130) );
  XOR U4095 ( .A(n4132), .B(n4133), .Z(n4124) );
  AND U4096 ( .A(n329), .B(n4123), .Z(n4133) );
  XNOR U4097 ( .A(n4134), .B(n4121), .Z(n4123) );
  XOR U4098 ( .A(n4135), .B(n4136), .Z(n4121) );
  AND U4099 ( .A(n352), .B(n4137), .Z(n4136) );
  IV U4100 ( .A(n4132), .Z(n4134) );
  XOR U4101 ( .A(n4138), .B(n4139), .Z(n4132) );
  AND U4102 ( .A(n336), .B(n4131), .Z(n4139) );
  XNOR U4103 ( .A(n4129), .B(n4138), .Z(n4131) );
  XNOR U4104 ( .A(n4140), .B(n4141), .Z(n4129) );
  AND U4105 ( .A(n340), .B(n4142), .Z(n4141) );
  XOR U4106 ( .A(p_input[353]), .B(n4140), .Z(n4142) );
  XNOR U4107 ( .A(n4143), .B(n4144), .Z(n4140) );
  AND U4108 ( .A(n344), .B(n4145), .Z(n4144) );
  XOR U4109 ( .A(n4146), .B(n4147), .Z(n4138) );
  AND U4110 ( .A(n348), .B(n4137), .Z(n4147) );
  XNOR U4111 ( .A(n4148), .B(n4135), .Z(n4137) );
  XOR U4112 ( .A(n4149), .B(n4150), .Z(n4135) );
  AND U4113 ( .A(n370), .B(n4151), .Z(n4150) );
  IV U4114 ( .A(n4146), .Z(n4148) );
  XOR U4115 ( .A(n4152), .B(n4153), .Z(n4146) );
  AND U4116 ( .A(n355), .B(n4145), .Z(n4153) );
  XNOR U4117 ( .A(n4143), .B(n4152), .Z(n4145) );
  XNOR U4118 ( .A(n4154), .B(n4155), .Z(n4143) );
  AND U4119 ( .A(n359), .B(n4156), .Z(n4155) );
  XOR U4120 ( .A(p_input[385]), .B(n4154), .Z(n4156) );
  XOR U4121 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n4157), 
        .Z(n4154) );
  AND U4122 ( .A(n362), .B(n4158), .Z(n4157) );
  XOR U4123 ( .A(n4159), .B(n4160), .Z(n4152) );
  AND U4124 ( .A(n366), .B(n4151), .Z(n4160) );
  XNOR U4125 ( .A(n4161), .B(n4149), .Z(n4151) );
  XOR U4126 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n4162), .Z(n4149) );
  AND U4127 ( .A(n378), .B(n4163), .Z(n4162) );
  IV U4128 ( .A(n4159), .Z(n4161) );
  XOR U4129 ( .A(n4164), .B(n4165), .Z(n4159) );
  AND U4130 ( .A(n373), .B(n4158), .Z(n4165) );
  XOR U4131 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n4164), 
        .Z(n4158) );
  XOR U4132 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(n4166), 
        .Z(n4164) );
  AND U4133 ( .A(n375), .B(n4163), .Z(n4166) );
  XOR U4134 ( .A(\knn_comb_/min_val_out[0][1] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .Z(n4163) );
  XOR U4135 ( .A(n99), .B(n4167), .Z(o[19]) );
  AND U4136 ( .A(n122), .B(n4168), .Z(n99) );
  XOR U4137 ( .A(n100), .B(n4167), .Z(n4168) );
  XOR U4138 ( .A(n4169), .B(n4170), .Z(n4167) );
  AND U4139 ( .A(n142), .B(n4171), .Z(n4170) );
  XOR U4140 ( .A(n4172), .B(n29), .Z(n100) );
  AND U4141 ( .A(n125), .B(n4173), .Z(n29) );
  XOR U4142 ( .A(n30), .B(n4172), .Z(n4173) );
  XOR U4143 ( .A(n4174), .B(n4175), .Z(n30) );
  AND U4144 ( .A(n130), .B(n4176), .Z(n4175) );
  XOR U4145 ( .A(p_input[19]), .B(n4174), .Z(n4176) );
  XNOR U4146 ( .A(n4177), .B(n4178), .Z(n4174) );
  AND U4147 ( .A(n134), .B(n4179), .Z(n4178) );
  XOR U4148 ( .A(n4180), .B(n4181), .Z(n4172) );
  AND U4149 ( .A(n138), .B(n4171), .Z(n4181) );
  XNOR U4150 ( .A(n4182), .B(n4169), .Z(n4171) );
  XOR U4151 ( .A(n4183), .B(n4184), .Z(n4169) );
  AND U4152 ( .A(n162), .B(n4185), .Z(n4184) );
  IV U4153 ( .A(n4180), .Z(n4182) );
  XOR U4154 ( .A(n4186), .B(n4187), .Z(n4180) );
  AND U4155 ( .A(n146), .B(n4179), .Z(n4187) );
  XNOR U4156 ( .A(n4177), .B(n4186), .Z(n4179) );
  XNOR U4157 ( .A(n4188), .B(n4189), .Z(n4177) );
  AND U4158 ( .A(n150), .B(n4190), .Z(n4189) );
  XOR U4159 ( .A(p_input[51]), .B(n4188), .Z(n4190) );
  XNOR U4160 ( .A(n4191), .B(n4192), .Z(n4188) );
  AND U4161 ( .A(n154), .B(n4193), .Z(n4192) );
  XOR U4162 ( .A(n4194), .B(n4195), .Z(n4186) );
  AND U4163 ( .A(n158), .B(n4185), .Z(n4195) );
  XNOR U4164 ( .A(n4196), .B(n4183), .Z(n4185) );
  XOR U4165 ( .A(n4197), .B(n4198), .Z(n4183) );
  AND U4166 ( .A(n181), .B(n4199), .Z(n4198) );
  IV U4167 ( .A(n4194), .Z(n4196) );
  XOR U4168 ( .A(n4200), .B(n4201), .Z(n4194) );
  AND U4169 ( .A(n165), .B(n4193), .Z(n4201) );
  XNOR U4170 ( .A(n4191), .B(n4200), .Z(n4193) );
  XNOR U4171 ( .A(n4202), .B(n4203), .Z(n4191) );
  AND U4172 ( .A(n169), .B(n4204), .Z(n4203) );
  XOR U4173 ( .A(p_input[83]), .B(n4202), .Z(n4204) );
  XNOR U4174 ( .A(n4205), .B(n4206), .Z(n4202) );
  AND U4175 ( .A(n173), .B(n4207), .Z(n4206) );
  XOR U4176 ( .A(n4208), .B(n4209), .Z(n4200) );
  AND U4177 ( .A(n177), .B(n4199), .Z(n4209) );
  XNOR U4178 ( .A(n4210), .B(n4197), .Z(n4199) );
  XOR U4179 ( .A(n4211), .B(n4212), .Z(n4197) );
  AND U4180 ( .A(n200), .B(n4213), .Z(n4212) );
  IV U4181 ( .A(n4208), .Z(n4210) );
  XOR U4182 ( .A(n4214), .B(n4215), .Z(n4208) );
  AND U4183 ( .A(n184), .B(n4207), .Z(n4215) );
  XNOR U4184 ( .A(n4205), .B(n4214), .Z(n4207) );
  XNOR U4185 ( .A(n4216), .B(n4217), .Z(n4205) );
  AND U4186 ( .A(n188), .B(n4218), .Z(n4217) );
  XOR U4187 ( .A(p_input[115]), .B(n4216), .Z(n4218) );
  XNOR U4188 ( .A(n4219), .B(n4220), .Z(n4216) );
  AND U4189 ( .A(n192), .B(n4221), .Z(n4220) );
  XOR U4190 ( .A(n4222), .B(n4223), .Z(n4214) );
  AND U4191 ( .A(n196), .B(n4213), .Z(n4223) );
  XNOR U4192 ( .A(n4224), .B(n4211), .Z(n4213) );
  XOR U4193 ( .A(n4225), .B(n4226), .Z(n4211) );
  AND U4194 ( .A(n219), .B(n4227), .Z(n4226) );
  IV U4195 ( .A(n4222), .Z(n4224) );
  XOR U4196 ( .A(n4228), .B(n4229), .Z(n4222) );
  AND U4197 ( .A(n203), .B(n4221), .Z(n4229) );
  XNOR U4198 ( .A(n4219), .B(n4228), .Z(n4221) );
  XNOR U4199 ( .A(n4230), .B(n4231), .Z(n4219) );
  AND U4200 ( .A(n207), .B(n4232), .Z(n4231) );
  XOR U4201 ( .A(p_input[147]), .B(n4230), .Z(n4232) );
  XNOR U4202 ( .A(n4233), .B(n4234), .Z(n4230) );
  AND U4203 ( .A(n211), .B(n4235), .Z(n4234) );
  XOR U4204 ( .A(n4236), .B(n4237), .Z(n4228) );
  AND U4205 ( .A(n215), .B(n4227), .Z(n4237) );
  XNOR U4206 ( .A(n4238), .B(n4225), .Z(n4227) );
  XOR U4207 ( .A(n4239), .B(n4240), .Z(n4225) );
  AND U4208 ( .A(n238), .B(n4241), .Z(n4240) );
  IV U4209 ( .A(n4236), .Z(n4238) );
  XOR U4210 ( .A(n4242), .B(n4243), .Z(n4236) );
  AND U4211 ( .A(n222), .B(n4235), .Z(n4243) );
  XNOR U4212 ( .A(n4233), .B(n4242), .Z(n4235) );
  XNOR U4213 ( .A(n4244), .B(n4245), .Z(n4233) );
  AND U4214 ( .A(n226), .B(n4246), .Z(n4245) );
  XOR U4215 ( .A(p_input[179]), .B(n4244), .Z(n4246) );
  XNOR U4216 ( .A(n4247), .B(n4248), .Z(n4244) );
  AND U4217 ( .A(n230), .B(n4249), .Z(n4248) );
  XOR U4218 ( .A(n4250), .B(n4251), .Z(n4242) );
  AND U4219 ( .A(n234), .B(n4241), .Z(n4251) );
  XNOR U4220 ( .A(n4252), .B(n4239), .Z(n4241) );
  XOR U4221 ( .A(n4253), .B(n4254), .Z(n4239) );
  AND U4222 ( .A(n257), .B(n4255), .Z(n4254) );
  IV U4223 ( .A(n4250), .Z(n4252) );
  XOR U4224 ( .A(n4256), .B(n4257), .Z(n4250) );
  AND U4225 ( .A(n241), .B(n4249), .Z(n4257) );
  XNOR U4226 ( .A(n4247), .B(n4256), .Z(n4249) );
  XNOR U4227 ( .A(n4258), .B(n4259), .Z(n4247) );
  AND U4228 ( .A(n245), .B(n4260), .Z(n4259) );
  XOR U4229 ( .A(p_input[211]), .B(n4258), .Z(n4260) );
  XNOR U4230 ( .A(n4261), .B(n4262), .Z(n4258) );
  AND U4231 ( .A(n249), .B(n4263), .Z(n4262) );
  XOR U4232 ( .A(n4264), .B(n4265), .Z(n4256) );
  AND U4233 ( .A(n253), .B(n4255), .Z(n4265) );
  XNOR U4234 ( .A(n4266), .B(n4253), .Z(n4255) );
  XOR U4235 ( .A(n4267), .B(n4268), .Z(n4253) );
  AND U4236 ( .A(n276), .B(n4269), .Z(n4268) );
  IV U4237 ( .A(n4264), .Z(n4266) );
  XOR U4238 ( .A(n4270), .B(n4271), .Z(n4264) );
  AND U4239 ( .A(n260), .B(n4263), .Z(n4271) );
  XNOR U4240 ( .A(n4261), .B(n4270), .Z(n4263) );
  XNOR U4241 ( .A(n4272), .B(n4273), .Z(n4261) );
  AND U4242 ( .A(n264), .B(n4274), .Z(n4273) );
  XOR U4243 ( .A(p_input[243]), .B(n4272), .Z(n4274) );
  XNOR U4244 ( .A(n4275), .B(n4276), .Z(n4272) );
  AND U4245 ( .A(n268), .B(n4277), .Z(n4276) );
  XOR U4246 ( .A(n4278), .B(n4279), .Z(n4270) );
  AND U4247 ( .A(n272), .B(n4269), .Z(n4279) );
  XNOR U4248 ( .A(n4280), .B(n4267), .Z(n4269) );
  XOR U4249 ( .A(n4281), .B(n4282), .Z(n4267) );
  AND U4250 ( .A(n295), .B(n4283), .Z(n4282) );
  IV U4251 ( .A(n4278), .Z(n4280) );
  XOR U4252 ( .A(n4284), .B(n4285), .Z(n4278) );
  AND U4253 ( .A(n279), .B(n4277), .Z(n4285) );
  XNOR U4254 ( .A(n4275), .B(n4284), .Z(n4277) );
  XNOR U4255 ( .A(n4286), .B(n4287), .Z(n4275) );
  AND U4256 ( .A(n283), .B(n4288), .Z(n4287) );
  XOR U4257 ( .A(p_input[275]), .B(n4286), .Z(n4288) );
  XNOR U4258 ( .A(n4289), .B(n4290), .Z(n4286) );
  AND U4259 ( .A(n287), .B(n4291), .Z(n4290) );
  XOR U4260 ( .A(n4292), .B(n4293), .Z(n4284) );
  AND U4261 ( .A(n291), .B(n4283), .Z(n4293) );
  XNOR U4262 ( .A(n4294), .B(n4281), .Z(n4283) );
  XOR U4263 ( .A(n4295), .B(n4296), .Z(n4281) );
  AND U4264 ( .A(n314), .B(n4297), .Z(n4296) );
  IV U4265 ( .A(n4292), .Z(n4294) );
  XOR U4266 ( .A(n4298), .B(n4299), .Z(n4292) );
  AND U4267 ( .A(n298), .B(n4291), .Z(n4299) );
  XNOR U4268 ( .A(n4289), .B(n4298), .Z(n4291) );
  XNOR U4269 ( .A(n4300), .B(n4301), .Z(n4289) );
  AND U4270 ( .A(n302), .B(n4302), .Z(n4301) );
  XOR U4271 ( .A(p_input[307]), .B(n4300), .Z(n4302) );
  XNOR U4272 ( .A(n4303), .B(n4304), .Z(n4300) );
  AND U4273 ( .A(n306), .B(n4305), .Z(n4304) );
  XOR U4274 ( .A(n4306), .B(n4307), .Z(n4298) );
  AND U4275 ( .A(n310), .B(n4297), .Z(n4307) );
  XNOR U4276 ( .A(n4308), .B(n4295), .Z(n4297) );
  XOR U4277 ( .A(n4309), .B(n4310), .Z(n4295) );
  AND U4278 ( .A(n333), .B(n4311), .Z(n4310) );
  IV U4279 ( .A(n4306), .Z(n4308) );
  XOR U4280 ( .A(n4312), .B(n4313), .Z(n4306) );
  AND U4281 ( .A(n317), .B(n4305), .Z(n4313) );
  XNOR U4282 ( .A(n4303), .B(n4312), .Z(n4305) );
  XNOR U4283 ( .A(n4314), .B(n4315), .Z(n4303) );
  AND U4284 ( .A(n321), .B(n4316), .Z(n4315) );
  XOR U4285 ( .A(p_input[339]), .B(n4314), .Z(n4316) );
  XNOR U4286 ( .A(n4317), .B(n4318), .Z(n4314) );
  AND U4287 ( .A(n325), .B(n4319), .Z(n4318) );
  XOR U4288 ( .A(n4320), .B(n4321), .Z(n4312) );
  AND U4289 ( .A(n329), .B(n4311), .Z(n4321) );
  XNOR U4290 ( .A(n4322), .B(n4309), .Z(n4311) );
  XOR U4291 ( .A(n4323), .B(n4324), .Z(n4309) );
  AND U4292 ( .A(n352), .B(n4325), .Z(n4324) );
  IV U4293 ( .A(n4320), .Z(n4322) );
  XOR U4294 ( .A(n4326), .B(n4327), .Z(n4320) );
  AND U4295 ( .A(n336), .B(n4319), .Z(n4327) );
  XNOR U4296 ( .A(n4317), .B(n4326), .Z(n4319) );
  XNOR U4297 ( .A(n4328), .B(n4329), .Z(n4317) );
  AND U4298 ( .A(n340), .B(n4330), .Z(n4329) );
  XOR U4299 ( .A(p_input[371]), .B(n4328), .Z(n4330) );
  XNOR U4300 ( .A(n4331), .B(n4332), .Z(n4328) );
  AND U4301 ( .A(n344), .B(n4333), .Z(n4332) );
  XOR U4302 ( .A(n4334), .B(n4335), .Z(n4326) );
  AND U4303 ( .A(n348), .B(n4325), .Z(n4335) );
  XNOR U4304 ( .A(n4336), .B(n4323), .Z(n4325) );
  XOR U4305 ( .A(n4337), .B(n4338), .Z(n4323) );
  AND U4306 ( .A(n370), .B(n4339), .Z(n4338) );
  IV U4307 ( .A(n4334), .Z(n4336) );
  XOR U4308 ( .A(n4340), .B(n4341), .Z(n4334) );
  AND U4309 ( .A(n355), .B(n4333), .Z(n4341) );
  XNOR U4310 ( .A(n4331), .B(n4340), .Z(n4333) );
  XNOR U4311 ( .A(n4342), .B(n4343), .Z(n4331) );
  AND U4312 ( .A(n359), .B(n4344), .Z(n4343) );
  XOR U4313 ( .A(p_input[403]), .B(n4342), .Z(n4344) );
  XOR U4314 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][19] ), .B(n4345), 
        .Z(n4342) );
  AND U4315 ( .A(n362), .B(n4346), .Z(n4345) );
  XOR U4316 ( .A(n4347), .B(n4348), .Z(n4340) );
  AND U4317 ( .A(n366), .B(n4339), .Z(n4348) );
  XNOR U4318 ( .A(n4349), .B(n4337), .Z(n4339) );
  XOR U4319 ( .A(\knn_comb_/min_val_out[0][19] ), .B(n4350), .Z(n4337) );
  AND U4320 ( .A(n378), .B(n4351), .Z(n4350) );
  IV U4321 ( .A(n4347), .Z(n4349) );
  XOR U4322 ( .A(n4352), .B(n4353), .Z(n4347) );
  AND U4323 ( .A(n373), .B(n4346), .Z(n4353) );
  XOR U4324 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][19] ), .B(n4352), 
        .Z(n4346) );
  XOR U4325 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .B(n4354), 
        .Z(n4352) );
  AND U4326 ( .A(n375), .B(n4351), .Z(n4354) );
  XOR U4327 ( .A(\knn_comb_/min_val_out[0][19] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .Z(n4351) );
  XOR U4328 ( .A(n101), .B(n4355), .Z(o[18]) );
  AND U4329 ( .A(n122), .B(n4356), .Z(n101) );
  XOR U4330 ( .A(n102), .B(n4355), .Z(n4356) );
  XOR U4331 ( .A(n4357), .B(n4358), .Z(n4355) );
  AND U4332 ( .A(n142), .B(n4359), .Z(n4358) );
  XOR U4333 ( .A(n4360), .B(n31), .Z(n102) );
  AND U4334 ( .A(n125), .B(n4361), .Z(n31) );
  XOR U4335 ( .A(n32), .B(n4360), .Z(n4361) );
  XOR U4336 ( .A(n4362), .B(n4363), .Z(n32) );
  AND U4337 ( .A(n130), .B(n4364), .Z(n4363) );
  XOR U4338 ( .A(p_input[18]), .B(n4362), .Z(n4364) );
  XNOR U4339 ( .A(n4365), .B(n4366), .Z(n4362) );
  AND U4340 ( .A(n134), .B(n4367), .Z(n4366) );
  XOR U4341 ( .A(n4368), .B(n4369), .Z(n4360) );
  AND U4342 ( .A(n138), .B(n4359), .Z(n4369) );
  XNOR U4343 ( .A(n4370), .B(n4357), .Z(n4359) );
  XOR U4344 ( .A(n4371), .B(n4372), .Z(n4357) );
  AND U4345 ( .A(n162), .B(n4373), .Z(n4372) );
  IV U4346 ( .A(n4368), .Z(n4370) );
  XOR U4347 ( .A(n4374), .B(n4375), .Z(n4368) );
  AND U4348 ( .A(n146), .B(n4367), .Z(n4375) );
  XNOR U4349 ( .A(n4365), .B(n4374), .Z(n4367) );
  XNOR U4350 ( .A(n4376), .B(n4377), .Z(n4365) );
  AND U4351 ( .A(n150), .B(n4378), .Z(n4377) );
  XOR U4352 ( .A(p_input[50]), .B(n4376), .Z(n4378) );
  XNOR U4353 ( .A(n4379), .B(n4380), .Z(n4376) );
  AND U4354 ( .A(n154), .B(n4381), .Z(n4380) );
  XOR U4355 ( .A(n4382), .B(n4383), .Z(n4374) );
  AND U4356 ( .A(n158), .B(n4373), .Z(n4383) );
  XNOR U4357 ( .A(n4384), .B(n4371), .Z(n4373) );
  XOR U4358 ( .A(n4385), .B(n4386), .Z(n4371) );
  AND U4359 ( .A(n181), .B(n4387), .Z(n4386) );
  IV U4360 ( .A(n4382), .Z(n4384) );
  XOR U4361 ( .A(n4388), .B(n4389), .Z(n4382) );
  AND U4362 ( .A(n165), .B(n4381), .Z(n4389) );
  XNOR U4363 ( .A(n4379), .B(n4388), .Z(n4381) );
  XNOR U4364 ( .A(n4390), .B(n4391), .Z(n4379) );
  AND U4365 ( .A(n169), .B(n4392), .Z(n4391) );
  XOR U4366 ( .A(p_input[82]), .B(n4390), .Z(n4392) );
  XNOR U4367 ( .A(n4393), .B(n4394), .Z(n4390) );
  AND U4368 ( .A(n173), .B(n4395), .Z(n4394) );
  XOR U4369 ( .A(n4396), .B(n4397), .Z(n4388) );
  AND U4370 ( .A(n177), .B(n4387), .Z(n4397) );
  XNOR U4371 ( .A(n4398), .B(n4385), .Z(n4387) );
  XOR U4372 ( .A(n4399), .B(n4400), .Z(n4385) );
  AND U4373 ( .A(n200), .B(n4401), .Z(n4400) );
  IV U4374 ( .A(n4396), .Z(n4398) );
  XOR U4375 ( .A(n4402), .B(n4403), .Z(n4396) );
  AND U4376 ( .A(n184), .B(n4395), .Z(n4403) );
  XNOR U4377 ( .A(n4393), .B(n4402), .Z(n4395) );
  XNOR U4378 ( .A(n4404), .B(n4405), .Z(n4393) );
  AND U4379 ( .A(n188), .B(n4406), .Z(n4405) );
  XOR U4380 ( .A(p_input[114]), .B(n4404), .Z(n4406) );
  XNOR U4381 ( .A(n4407), .B(n4408), .Z(n4404) );
  AND U4382 ( .A(n192), .B(n4409), .Z(n4408) );
  XOR U4383 ( .A(n4410), .B(n4411), .Z(n4402) );
  AND U4384 ( .A(n196), .B(n4401), .Z(n4411) );
  XNOR U4385 ( .A(n4412), .B(n4399), .Z(n4401) );
  XOR U4386 ( .A(n4413), .B(n4414), .Z(n4399) );
  AND U4387 ( .A(n219), .B(n4415), .Z(n4414) );
  IV U4388 ( .A(n4410), .Z(n4412) );
  XOR U4389 ( .A(n4416), .B(n4417), .Z(n4410) );
  AND U4390 ( .A(n203), .B(n4409), .Z(n4417) );
  XNOR U4391 ( .A(n4407), .B(n4416), .Z(n4409) );
  XNOR U4392 ( .A(n4418), .B(n4419), .Z(n4407) );
  AND U4393 ( .A(n207), .B(n4420), .Z(n4419) );
  XOR U4394 ( .A(p_input[146]), .B(n4418), .Z(n4420) );
  XNOR U4395 ( .A(n4421), .B(n4422), .Z(n4418) );
  AND U4396 ( .A(n211), .B(n4423), .Z(n4422) );
  XOR U4397 ( .A(n4424), .B(n4425), .Z(n4416) );
  AND U4398 ( .A(n215), .B(n4415), .Z(n4425) );
  XNOR U4399 ( .A(n4426), .B(n4413), .Z(n4415) );
  XOR U4400 ( .A(n4427), .B(n4428), .Z(n4413) );
  AND U4401 ( .A(n238), .B(n4429), .Z(n4428) );
  IV U4402 ( .A(n4424), .Z(n4426) );
  XOR U4403 ( .A(n4430), .B(n4431), .Z(n4424) );
  AND U4404 ( .A(n222), .B(n4423), .Z(n4431) );
  XNOR U4405 ( .A(n4421), .B(n4430), .Z(n4423) );
  XNOR U4406 ( .A(n4432), .B(n4433), .Z(n4421) );
  AND U4407 ( .A(n226), .B(n4434), .Z(n4433) );
  XOR U4408 ( .A(p_input[178]), .B(n4432), .Z(n4434) );
  XNOR U4409 ( .A(n4435), .B(n4436), .Z(n4432) );
  AND U4410 ( .A(n230), .B(n4437), .Z(n4436) );
  XOR U4411 ( .A(n4438), .B(n4439), .Z(n4430) );
  AND U4412 ( .A(n234), .B(n4429), .Z(n4439) );
  XNOR U4413 ( .A(n4440), .B(n4427), .Z(n4429) );
  XOR U4414 ( .A(n4441), .B(n4442), .Z(n4427) );
  AND U4415 ( .A(n257), .B(n4443), .Z(n4442) );
  IV U4416 ( .A(n4438), .Z(n4440) );
  XOR U4417 ( .A(n4444), .B(n4445), .Z(n4438) );
  AND U4418 ( .A(n241), .B(n4437), .Z(n4445) );
  XNOR U4419 ( .A(n4435), .B(n4444), .Z(n4437) );
  XNOR U4420 ( .A(n4446), .B(n4447), .Z(n4435) );
  AND U4421 ( .A(n245), .B(n4448), .Z(n4447) );
  XOR U4422 ( .A(p_input[210]), .B(n4446), .Z(n4448) );
  XNOR U4423 ( .A(n4449), .B(n4450), .Z(n4446) );
  AND U4424 ( .A(n249), .B(n4451), .Z(n4450) );
  XOR U4425 ( .A(n4452), .B(n4453), .Z(n4444) );
  AND U4426 ( .A(n253), .B(n4443), .Z(n4453) );
  XNOR U4427 ( .A(n4454), .B(n4441), .Z(n4443) );
  XOR U4428 ( .A(n4455), .B(n4456), .Z(n4441) );
  AND U4429 ( .A(n276), .B(n4457), .Z(n4456) );
  IV U4430 ( .A(n4452), .Z(n4454) );
  XOR U4431 ( .A(n4458), .B(n4459), .Z(n4452) );
  AND U4432 ( .A(n260), .B(n4451), .Z(n4459) );
  XNOR U4433 ( .A(n4449), .B(n4458), .Z(n4451) );
  XNOR U4434 ( .A(n4460), .B(n4461), .Z(n4449) );
  AND U4435 ( .A(n264), .B(n4462), .Z(n4461) );
  XOR U4436 ( .A(p_input[242]), .B(n4460), .Z(n4462) );
  XNOR U4437 ( .A(n4463), .B(n4464), .Z(n4460) );
  AND U4438 ( .A(n268), .B(n4465), .Z(n4464) );
  XOR U4439 ( .A(n4466), .B(n4467), .Z(n4458) );
  AND U4440 ( .A(n272), .B(n4457), .Z(n4467) );
  XNOR U4441 ( .A(n4468), .B(n4455), .Z(n4457) );
  XOR U4442 ( .A(n4469), .B(n4470), .Z(n4455) );
  AND U4443 ( .A(n295), .B(n4471), .Z(n4470) );
  IV U4444 ( .A(n4466), .Z(n4468) );
  XOR U4445 ( .A(n4472), .B(n4473), .Z(n4466) );
  AND U4446 ( .A(n279), .B(n4465), .Z(n4473) );
  XNOR U4447 ( .A(n4463), .B(n4472), .Z(n4465) );
  XNOR U4448 ( .A(n4474), .B(n4475), .Z(n4463) );
  AND U4449 ( .A(n283), .B(n4476), .Z(n4475) );
  XOR U4450 ( .A(p_input[274]), .B(n4474), .Z(n4476) );
  XNOR U4451 ( .A(n4477), .B(n4478), .Z(n4474) );
  AND U4452 ( .A(n287), .B(n4479), .Z(n4478) );
  XOR U4453 ( .A(n4480), .B(n4481), .Z(n4472) );
  AND U4454 ( .A(n291), .B(n4471), .Z(n4481) );
  XNOR U4455 ( .A(n4482), .B(n4469), .Z(n4471) );
  XOR U4456 ( .A(n4483), .B(n4484), .Z(n4469) );
  AND U4457 ( .A(n314), .B(n4485), .Z(n4484) );
  IV U4458 ( .A(n4480), .Z(n4482) );
  XOR U4459 ( .A(n4486), .B(n4487), .Z(n4480) );
  AND U4460 ( .A(n298), .B(n4479), .Z(n4487) );
  XNOR U4461 ( .A(n4477), .B(n4486), .Z(n4479) );
  XNOR U4462 ( .A(n4488), .B(n4489), .Z(n4477) );
  AND U4463 ( .A(n302), .B(n4490), .Z(n4489) );
  XOR U4464 ( .A(p_input[306]), .B(n4488), .Z(n4490) );
  XNOR U4465 ( .A(n4491), .B(n4492), .Z(n4488) );
  AND U4466 ( .A(n306), .B(n4493), .Z(n4492) );
  XOR U4467 ( .A(n4494), .B(n4495), .Z(n4486) );
  AND U4468 ( .A(n310), .B(n4485), .Z(n4495) );
  XNOR U4469 ( .A(n4496), .B(n4483), .Z(n4485) );
  XOR U4470 ( .A(n4497), .B(n4498), .Z(n4483) );
  AND U4471 ( .A(n333), .B(n4499), .Z(n4498) );
  IV U4472 ( .A(n4494), .Z(n4496) );
  XOR U4473 ( .A(n4500), .B(n4501), .Z(n4494) );
  AND U4474 ( .A(n317), .B(n4493), .Z(n4501) );
  XNOR U4475 ( .A(n4491), .B(n4500), .Z(n4493) );
  XNOR U4476 ( .A(n4502), .B(n4503), .Z(n4491) );
  AND U4477 ( .A(n321), .B(n4504), .Z(n4503) );
  XOR U4478 ( .A(p_input[338]), .B(n4502), .Z(n4504) );
  XNOR U4479 ( .A(n4505), .B(n4506), .Z(n4502) );
  AND U4480 ( .A(n325), .B(n4507), .Z(n4506) );
  XOR U4481 ( .A(n4508), .B(n4509), .Z(n4500) );
  AND U4482 ( .A(n329), .B(n4499), .Z(n4509) );
  XNOR U4483 ( .A(n4510), .B(n4497), .Z(n4499) );
  XOR U4484 ( .A(n4511), .B(n4512), .Z(n4497) );
  AND U4485 ( .A(n352), .B(n4513), .Z(n4512) );
  IV U4486 ( .A(n4508), .Z(n4510) );
  XOR U4487 ( .A(n4514), .B(n4515), .Z(n4508) );
  AND U4488 ( .A(n336), .B(n4507), .Z(n4515) );
  XNOR U4489 ( .A(n4505), .B(n4514), .Z(n4507) );
  XNOR U4490 ( .A(n4516), .B(n4517), .Z(n4505) );
  AND U4491 ( .A(n340), .B(n4518), .Z(n4517) );
  XOR U4492 ( .A(p_input[370]), .B(n4516), .Z(n4518) );
  XNOR U4493 ( .A(n4519), .B(n4520), .Z(n4516) );
  AND U4494 ( .A(n344), .B(n4521), .Z(n4520) );
  XOR U4495 ( .A(n4522), .B(n4523), .Z(n4514) );
  AND U4496 ( .A(n348), .B(n4513), .Z(n4523) );
  XNOR U4497 ( .A(n4524), .B(n4511), .Z(n4513) );
  XOR U4498 ( .A(n4525), .B(n4526), .Z(n4511) );
  AND U4499 ( .A(n370), .B(n4527), .Z(n4526) );
  IV U4500 ( .A(n4522), .Z(n4524) );
  XOR U4501 ( .A(n4528), .B(n4529), .Z(n4522) );
  AND U4502 ( .A(n355), .B(n4521), .Z(n4529) );
  XNOR U4503 ( .A(n4519), .B(n4528), .Z(n4521) );
  XNOR U4504 ( .A(n4530), .B(n4531), .Z(n4519) );
  AND U4505 ( .A(n359), .B(n4532), .Z(n4531) );
  XOR U4506 ( .A(p_input[402]), .B(n4530), .Z(n4532) );
  XOR U4507 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][18] ), .B(n4533), 
        .Z(n4530) );
  AND U4508 ( .A(n362), .B(n4534), .Z(n4533) );
  XOR U4509 ( .A(n4535), .B(n4536), .Z(n4528) );
  AND U4510 ( .A(n366), .B(n4527), .Z(n4536) );
  XNOR U4511 ( .A(n4537), .B(n4525), .Z(n4527) );
  XOR U4512 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n4538), .Z(n4525) );
  AND U4513 ( .A(n378), .B(n4539), .Z(n4538) );
  IV U4514 ( .A(n4535), .Z(n4537) );
  XOR U4515 ( .A(n4540), .B(n4541), .Z(n4535) );
  AND U4516 ( .A(n373), .B(n4534), .Z(n4541) );
  XOR U4517 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][18] ), .B(n4540), 
        .Z(n4534) );
  XOR U4518 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .B(n4542), 
        .Z(n4540) );
  AND U4519 ( .A(n375), .B(n4539), .Z(n4542) );
  XOR U4520 ( .A(\knn_comb_/min_val_out[0][18] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .Z(n4539) );
  XOR U4521 ( .A(n105), .B(n4543), .Z(o[17]) );
  AND U4522 ( .A(n122), .B(n4544), .Z(n105) );
  XOR U4523 ( .A(n106), .B(n4543), .Z(n4544) );
  XOR U4524 ( .A(n4545), .B(n4546), .Z(n4543) );
  AND U4525 ( .A(n142), .B(n4547), .Z(n4546) );
  XOR U4526 ( .A(n4548), .B(n33), .Z(n106) );
  AND U4527 ( .A(n125), .B(n4549), .Z(n33) );
  XOR U4528 ( .A(n34), .B(n4548), .Z(n4549) );
  XOR U4529 ( .A(n4550), .B(n4551), .Z(n34) );
  AND U4530 ( .A(n130), .B(n4552), .Z(n4551) );
  XOR U4531 ( .A(p_input[17]), .B(n4550), .Z(n4552) );
  XNOR U4532 ( .A(n4553), .B(n4554), .Z(n4550) );
  AND U4533 ( .A(n134), .B(n4555), .Z(n4554) );
  XOR U4534 ( .A(n4556), .B(n4557), .Z(n4548) );
  AND U4535 ( .A(n138), .B(n4547), .Z(n4557) );
  XNOR U4536 ( .A(n4558), .B(n4545), .Z(n4547) );
  XOR U4537 ( .A(n4559), .B(n4560), .Z(n4545) );
  AND U4538 ( .A(n162), .B(n4561), .Z(n4560) );
  IV U4539 ( .A(n4556), .Z(n4558) );
  XOR U4540 ( .A(n4562), .B(n4563), .Z(n4556) );
  AND U4541 ( .A(n146), .B(n4555), .Z(n4563) );
  XNOR U4542 ( .A(n4553), .B(n4562), .Z(n4555) );
  XNOR U4543 ( .A(n4564), .B(n4565), .Z(n4553) );
  AND U4544 ( .A(n150), .B(n4566), .Z(n4565) );
  XOR U4545 ( .A(p_input[49]), .B(n4564), .Z(n4566) );
  XNOR U4546 ( .A(n4567), .B(n4568), .Z(n4564) );
  AND U4547 ( .A(n154), .B(n4569), .Z(n4568) );
  XOR U4548 ( .A(n4570), .B(n4571), .Z(n4562) );
  AND U4549 ( .A(n158), .B(n4561), .Z(n4571) );
  XNOR U4550 ( .A(n4572), .B(n4559), .Z(n4561) );
  XOR U4551 ( .A(n4573), .B(n4574), .Z(n4559) );
  AND U4552 ( .A(n181), .B(n4575), .Z(n4574) );
  IV U4553 ( .A(n4570), .Z(n4572) );
  XOR U4554 ( .A(n4576), .B(n4577), .Z(n4570) );
  AND U4555 ( .A(n165), .B(n4569), .Z(n4577) );
  XNOR U4556 ( .A(n4567), .B(n4576), .Z(n4569) );
  XNOR U4557 ( .A(n4578), .B(n4579), .Z(n4567) );
  AND U4558 ( .A(n169), .B(n4580), .Z(n4579) );
  XOR U4559 ( .A(p_input[81]), .B(n4578), .Z(n4580) );
  XNOR U4560 ( .A(n4581), .B(n4582), .Z(n4578) );
  AND U4561 ( .A(n173), .B(n4583), .Z(n4582) );
  XOR U4562 ( .A(n4584), .B(n4585), .Z(n4576) );
  AND U4563 ( .A(n177), .B(n4575), .Z(n4585) );
  XNOR U4564 ( .A(n4586), .B(n4573), .Z(n4575) );
  XOR U4565 ( .A(n4587), .B(n4588), .Z(n4573) );
  AND U4566 ( .A(n200), .B(n4589), .Z(n4588) );
  IV U4567 ( .A(n4584), .Z(n4586) );
  XOR U4568 ( .A(n4590), .B(n4591), .Z(n4584) );
  AND U4569 ( .A(n184), .B(n4583), .Z(n4591) );
  XNOR U4570 ( .A(n4581), .B(n4590), .Z(n4583) );
  XNOR U4571 ( .A(n4592), .B(n4593), .Z(n4581) );
  AND U4572 ( .A(n188), .B(n4594), .Z(n4593) );
  XOR U4573 ( .A(p_input[113]), .B(n4592), .Z(n4594) );
  XNOR U4574 ( .A(n4595), .B(n4596), .Z(n4592) );
  AND U4575 ( .A(n192), .B(n4597), .Z(n4596) );
  XOR U4576 ( .A(n4598), .B(n4599), .Z(n4590) );
  AND U4577 ( .A(n196), .B(n4589), .Z(n4599) );
  XNOR U4578 ( .A(n4600), .B(n4587), .Z(n4589) );
  XOR U4579 ( .A(n4601), .B(n4602), .Z(n4587) );
  AND U4580 ( .A(n219), .B(n4603), .Z(n4602) );
  IV U4581 ( .A(n4598), .Z(n4600) );
  XOR U4582 ( .A(n4604), .B(n4605), .Z(n4598) );
  AND U4583 ( .A(n203), .B(n4597), .Z(n4605) );
  XNOR U4584 ( .A(n4595), .B(n4604), .Z(n4597) );
  XNOR U4585 ( .A(n4606), .B(n4607), .Z(n4595) );
  AND U4586 ( .A(n207), .B(n4608), .Z(n4607) );
  XOR U4587 ( .A(p_input[145]), .B(n4606), .Z(n4608) );
  XNOR U4588 ( .A(n4609), .B(n4610), .Z(n4606) );
  AND U4589 ( .A(n211), .B(n4611), .Z(n4610) );
  XOR U4590 ( .A(n4612), .B(n4613), .Z(n4604) );
  AND U4591 ( .A(n215), .B(n4603), .Z(n4613) );
  XNOR U4592 ( .A(n4614), .B(n4601), .Z(n4603) );
  XOR U4593 ( .A(n4615), .B(n4616), .Z(n4601) );
  AND U4594 ( .A(n238), .B(n4617), .Z(n4616) );
  IV U4595 ( .A(n4612), .Z(n4614) );
  XOR U4596 ( .A(n4618), .B(n4619), .Z(n4612) );
  AND U4597 ( .A(n222), .B(n4611), .Z(n4619) );
  XNOR U4598 ( .A(n4609), .B(n4618), .Z(n4611) );
  XNOR U4599 ( .A(n4620), .B(n4621), .Z(n4609) );
  AND U4600 ( .A(n226), .B(n4622), .Z(n4621) );
  XOR U4601 ( .A(p_input[177]), .B(n4620), .Z(n4622) );
  XNOR U4602 ( .A(n4623), .B(n4624), .Z(n4620) );
  AND U4603 ( .A(n230), .B(n4625), .Z(n4624) );
  XOR U4604 ( .A(n4626), .B(n4627), .Z(n4618) );
  AND U4605 ( .A(n234), .B(n4617), .Z(n4627) );
  XNOR U4606 ( .A(n4628), .B(n4615), .Z(n4617) );
  XOR U4607 ( .A(n4629), .B(n4630), .Z(n4615) );
  AND U4608 ( .A(n257), .B(n4631), .Z(n4630) );
  IV U4609 ( .A(n4626), .Z(n4628) );
  XOR U4610 ( .A(n4632), .B(n4633), .Z(n4626) );
  AND U4611 ( .A(n241), .B(n4625), .Z(n4633) );
  XNOR U4612 ( .A(n4623), .B(n4632), .Z(n4625) );
  XNOR U4613 ( .A(n4634), .B(n4635), .Z(n4623) );
  AND U4614 ( .A(n245), .B(n4636), .Z(n4635) );
  XOR U4615 ( .A(p_input[209]), .B(n4634), .Z(n4636) );
  XNOR U4616 ( .A(n4637), .B(n4638), .Z(n4634) );
  AND U4617 ( .A(n249), .B(n4639), .Z(n4638) );
  XOR U4618 ( .A(n4640), .B(n4641), .Z(n4632) );
  AND U4619 ( .A(n253), .B(n4631), .Z(n4641) );
  XNOR U4620 ( .A(n4642), .B(n4629), .Z(n4631) );
  XOR U4621 ( .A(n4643), .B(n4644), .Z(n4629) );
  AND U4622 ( .A(n276), .B(n4645), .Z(n4644) );
  IV U4623 ( .A(n4640), .Z(n4642) );
  XOR U4624 ( .A(n4646), .B(n4647), .Z(n4640) );
  AND U4625 ( .A(n260), .B(n4639), .Z(n4647) );
  XNOR U4626 ( .A(n4637), .B(n4646), .Z(n4639) );
  XNOR U4627 ( .A(n4648), .B(n4649), .Z(n4637) );
  AND U4628 ( .A(n264), .B(n4650), .Z(n4649) );
  XOR U4629 ( .A(p_input[241]), .B(n4648), .Z(n4650) );
  XNOR U4630 ( .A(n4651), .B(n4652), .Z(n4648) );
  AND U4631 ( .A(n268), .B(n4653), .Z(n4652) );
  XOR U4632 ( .A(n4654), .B(n4655), .Z(n4646) );
  AND U4633 ( .A(n272), .B(n4645), .Z(n4655) );
  XNOR U4634 ( .A(n4656), .B(n4643), .Z(n4645) );
  XOR U4635 ( .A(n4657), .B(n4658), .Z(n4643) );
  AND U4636 ( .A(n295), .B(n4659), .Z(n4658) );
  IV U4637 ( .A(n4654), .Z(n4656) );
  XOR U4638 ( .A(n4660), .B(n4661), .Z(n4654) );
  AND U4639 ( .A(n279), .B(n4653), .Z(n4661) );
  XNOR U4640 ( .A(n4651), .B(n4660), .Z(n4653) );
  XNOR U4641 ( .A(n4662), .B(n4663), .Z(n4651) );
  AND U4642 ( .A(n283), .B(n4664), .Z(n4663) );
  XOR U4643 ( .A(p_input[273]), .B(n4662), .Z(n4664) );
  XNOR U4644 ( .A(n4665), .B(n4666), .Z(n4662) );
  AND U4645 ( .A(n287), .B(n4667), .Z(n4666) );
  XOR U4646 ( .A(n4668), .B(n4669), .Z(n4660) );
  AND U4647 ( .A(n291), .B(n4659), .Z(n4669) );
  XNOR U4648 ( .A(n4670), .B(n4657), .Z(n4659) );
  XOR U4649 ( .A(n4671), .B(n4672), .Z(n4657) );
  AND U4650 ( .A(n314), .B(n4673), .Z(n4672) );
  IV U4651 ( .A(n4668), .Z(n4670) );
  XOR U4652 ( .A(n4674), .B(n4675), .Z(n4668) );
  AND U4653 ( .A(n298), .B(n4667), .Z(n4675) );
  XNOR U4654 ( .A(n4665), .B(n4674), .Z(n4667) );
  XNOR U4655 ( .A(n4676), .B(n4677), .Z(n4665) );
  AND U4656 ( .A(n302), .B(n4678), .Z(n4677) );
  XOR U4657 ( .A(p_input[305]), .B(n4676), .Z(n4678) );
  XNOR U4658 ( .A(n4679), .B(n4680), .Z(n4676) );
  AND U4659 ( .A(n306), .B(n4681), .Z(n4680) );
  XOR U4660 ( .A(n4682), .B(n4683), .Z(n4674) );
  AND U4661 ( .A(n310), .B(n4673), .Z(n4683) );
  XNOR U4662 ( .A(n4684), .B(n4671), .Z(n4673) );
  XOR U4663 ( .A(n4685), .B(n4686), .Z(n4671) );
  AND U4664 ( .A(n333), .B(n4687), .Z(n4686) );
  IV U4665 ( .A(n4682), .Z(n4684) );
  XOR U4666 ( .A(n4688), .B(n4689), .Z(n4682) );
  AND U4667 ( .A(n317), .B(n4681), .Z(n4689) );
  XNOR U4668 ( .A(n4679), .B(n4688), .Z(n4681) );
  XNOR U4669 ( .A(n4690), .B(n4691), .Z(n4679) );
  AND U4670 ( .A(n321), .B(n4692), .Z(n4691) );
  XOR U4671 ( .A(p_input[337]), .B(n4690), .Z(n4692) );
  XNOR U4672 ( .A(n4693), .B(n4694), .Z(n4690) );
  AND U4673 ( .A(n325), .B(n4695), .Z(n4694) );
  XOR U4674 ( .A(n4696), .B(n4697), .Z(n4688) );
  AND U4675 ( .A(n329), .B(n4687), .Z(n4697) );
  XNOR U4676 ( .A(n4698), .B(n4685), .Z(n4687) );
  XOR U4677 ( .A(n4699), .B(n4700), .Z(n4685) );
  AND U4678 ( .A(n352), .B(n4701), .Z(n4700) );
  IV U4679 ( .A(n4696), .Z(n4698) );
  XOR U4680 ( .A(n4702), .B(n4703), .Z(n4696) );
  AND U4681 ( .A(n336), .B(n4695), .Z(n4703) );
  XNOR U4682 ( .A(n4693), .B(n4702), .Z(n4695) );
  XNOR U4683 ( .A(n4704), .B(n4705), .Z(n4693) );
  AND U4684 ( .A(n340), .B(n4706), .Z(n4705) );
  XOR U4685 ( .A(p_input[369]), .B(n4704), .Z(n4706) );
  XNOR U4686 ( .A(n4707), .B(n4708), .Z(n4704) );
  AND U4687 ( .A(n344), .B(n4709), .Z(n4708) );
  XOR U4688 ( .A(n4710), .B(n4711), .Z(n4702) );
  AND U4689 ( .A(n348), .B(n4701), .Z(n4711) );
  XNOR U4690 ( .A(n4712), .B(n4699), .Z(n4701) );
  XOR U4691 ( .A(n4713), .B(n4714), .Z(n4699) );
  AND U4692 ( .A(n370), .B(n4715), .Z(n4714) );
  IV U4693 ( .A(n4710), .Z(n4712) );
  XOR U4694 ( .A(n4716), .B(n4717), .Z(n4710) );
  AND U4695 ( .A(n355), .B(n4709), .Z(n4717) );
  XNOR U4696 ( .A(n4707), .B(n4716), .Z(n4709) );
  XNOR U4697 ( .A(n4718), .B(n4719), .Z(n4707) );
  AND U4698 ( .A(n359), .B(n4720), .Z(n4719) );
  XOR U4699 ( .A(p_input[401]), .B(n4718), .Z(n4720) );
  XOR U4700 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][17] ), .B(n4721), 
        .Z(n4718) );
  AND U4701 ( .A(n362), .B(n4722), .Z(n4721) );
  XOR U4702 ( .A(n4723), .B(n4724), .Z(n4716) );
  AND U4703 ( .A(n366), .B(n4715), .Z(n4724) );
  XNOR U4704 ( .A(n4725), .B(n4713), .Z(n4715) );
  XOR U4705 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n4726), .Z(n4713) );
  AND U4706 ( .A(n378), .B(n4727), .Z(n4726) );
  IV U4707 ( .A(n4723), .Z(n4725) );
  XOR U4708 ( .A(n4728), .B(n4729), .Z(n4723) );
  AND U4709 ( .A(n373), .B(n4722), .Z(n4729) );
  XOR U4710 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][17] ), .B(n4728), 
        .Z(n4722) );
  XOR U4711 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .B(n4730), 
        .Z(n4728) );
  AND U4712 ( .A(n375), .B(n4727), .Z(n4730) );
  XOR U4713 ( .A(\knn_comb_/min_val_out[0][17] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .Z(n4727) );
  XOR U4714 ( .A(n107), .B(n4731), .Z(o[16]) );
  AND U4715 ( .A(n122), .B(n4732), .Z(n107) );
  XOR U4716 ( .A(n108), .B(n4731), .Z(n4732) );
  XOR U4717 ( .A(n4733), .B(n4734), .Z(n4731) );
  AND U4718 ( .A(n142), .B(n4735), .Z(n4734) );
  XOR U4719 ( .A(n4736), .B(n35), .Z(n108) );
  AND U4720 ( .A(n125), .B(n4737), .Z(n35) );
  XOR U4721 ( .A(n36), .B(n4736), .Z(n4737) );
  XOR U4722 ( .A(n4738), .B(n4739), .Z(n36) );
  AND U4723 ( .A(n130), .B(n4740), .Z(n4739) );
  XOR U4724 ( .A(p_input[16]), .B(n4738), .Z(n4740) );
  XNOR U4725 ( .A(n4741), .B(n4742), .Z(n4738) );
  AND U4726 ( .A(n134), .B(n4743), .Z(n4742) );
  XOR U4727 ( .A(n4744), .B(n4745), .Z(n4736) );
  AND U4728 ( .A(n138), .B(n4735), .Z(n4745) );
  XNOR U4729 ( .A(n4746), .B(n4733), .Z(n4735) );
  XOR U4730 ( .A(n4747), .B(n4748), .Z(n4733) );
  AND U4731 ( .A(n162), .B(n4749), .Z(n4748) );
  IV U4732 ( .A(n4744), .Z(n4746) );
  XOR U4733 ( .A(n4750), .B(n4751), .Z(n4744) );
  AND U4734 ( .A(n146), .B(n4743), .Z(n4751) );
  XNOR U4735 ( .A(n4741), .B(n4750), .Z(n4743) );
  XNOR U4736 ( .A(n4752), .B(n4753), .Z(n4741) );
  AND U4737 ( .A(n150), .B(n4754), .Z(n4753) );
  XOR U4738 ( .A(p_input[48]), .B(n4752), .Z(n4754) );
  XNOR U4739 ( .A(n4755), .B(n4756), .Z(n4752) );
  AND U4740 ( .A(n154), .B(n4757), .Z(n4756) );
  XOR U4741 ( .A(n4758), .B(n4759), .Z(n4750) );
  AND U4742 ( .A(n158), .B(n4749), .Z(n4759) );
  XNOR U4743 ( .A(n4760), .B(n4747), .Z(n4749) );
  XOR U4744 ( .A(n4761), .B(n4762), .Z(n4747) );
  AND U4745 ( .A(n181), .B(n4763), .Z(n4762) );
  IV U4746 ( .A(n4758), .Z(n4760) );
  XOR U4747 ( .A(n4764), .B(n4765), .Z(n4758) );
  AND U4748 ( .A(n165), .B(n4757), .Z(n4765) );
  XNOR U4749 ( .A(n4755), .B(n4764), .Z(n4757) );
  XNOR U4750 ( .A(n4766), .B(n4767), .Z(n4755) );
  AND U4751 ( .A(n169), .B(n4768), .Z(n4767) );
  XOR U4752 ( .A(p_input[80]), .B(n4766), .Z(n4768) );
  XNOR U4753 ( .A(n4769), .B(n4770), .Z(n4766) );
  AND U4754 ( .A(n173), .B(n4771), .Z(n4770) );
  XOR U4755 ( .A(n4772), .B(n4773), .Z(n4764) );
  AND U4756 ( .A(n177), .B(n4763), .Z(n4773) );
  XNOR U4757 ( .A(n4774), .B(n4761), .Z(n4763) );
  XOR U4758 ( .A(n4775), .B(n4776), .Z(n4761) );
  AND U4759 ( .A(n200), .B(n4777), .Z(n4776) );
  IV U4760 ( .A(n4772), .Z(n4774) );
  XOR U4761 ( .A(n4778), .B(n4779), .Z(n4772) );
  AND U4762 ( .A(n184), .B(n4771), .Z(n4779) );
  XNOR U4763 ( .A(n4769), .B(n4778), .Z(n4771) );
  XNOR U4764 ( .A(n4780), .B(n4781), .Z(n4769) );
  AND U4765 ( .A(n188), .B(n4782), .Z(n4781) );
  XOR U4766 ( .A(p_input[112]), .B(n4780), .Z(n4782) );
  XNOR U4767 ( .A(n4783), .B(n4784), .Z(n4780) );
  AND U4768 ( .A(n192), .B(n4785), .Z(n4784) );
  XOR U4769 ( .A(n4786), .B(n4787), .Z(n4778) );
  AND U4770 ( .A(n196), .B(n4777), .Z(n4787) );
  XNOR U4771 ( .A(n4788), .B(n4775), .Z(n4777) );
  XOR U4772 ( .A(n4789), .B(n4790), .Z(n4775) );
  AND U4773 ( .A(n219), .B(n4791), .Z(n4790) );
  IV U4774 ( .A(n4786), .Z(n4788) );
  XOR U4775 ( .A(n4792), .B(n4793), .Z(n4786) );
  AND U4776 ( .A(n203), .B(n4785), .Z(n4793) );
  XNOR U4777 ( .A(n4783), .B(n4792), .Z(n4785) );
  XNOR U4778 ( .A(n4794), .B(n4795), .Z(n4783) );
  AND U4779 ( .A(n207), .B(n4796), .Z(n4795) );
  XOR U4780 ( .A(p_input[144]), .B(n4794), .Z(n4796) );
  XNOR U4781 ( .A(n4797), .B(n4798), .Z(n4794) );
  AND U4782 ( .A(n211), .B(n4799), .Z(n4798) );
  XOR U4783 ( .A(n4800), .B(n4801), .Z(n4792) );
  AND U4784 ( .A(n215), .B(n4791), .Z(n4801) );
  XNOR U4785 ( .A(n4802), .B(n4789), .Z(n4791) );
  XOR U4786 ( .A(n4803), .B(n4804), .Z(n4789) );
  AND U4787 ( .A(n238), .B(n4805), .Z(n4804) );
  IV U4788 ( .A(n4800), .Z(n4802) );
  XOR U4789 ( .A(n4806), .B(n4807), .Z(n4800) );
  AND U4790 ( .A(n222), .B(n4799), .Z(n4807) );
  XNOR U4791 ( .A(n4797), .B(n4806), .Z(n4799) );
  XNOR U4792 ( .A(n4808), .B(n4809), .Z(n4797) );
  AND U4793 ( .A(n226), .B(n4810), .Z(n4809) );
  XOR U4794 ( .A(p_input[176]), .B(n4808), .Z(n4810) );
  XNOR U4795 ( .A(n4811), .B(n4812), .Z(n4808) );
  AND U4796 ( .A(n230), .B(n4813), .Z(n4812) );
  XOR U4797 ( .A(n4814), .B(n4815), .Z(n4806) );
  AND U4798 ( .A(n234), .B(n4805), .Z(n4815) );
  XNOR U4799 ( .A(n4816), .B(n4803), .Z(n4805) );
  XOR U4800 ( .A(n4817), .B(n4818), .Z(n4803) );
  AND U4801 ( .A(n257), .B(n4819), .Z(n4818) );
  IV U4802 ( .A(n4814), .Z(n4816) );
  XOR U4803 ( .A(n4820), .B(n4821), .Z(n4814) );
  AND U4804 ( .A(n241), .B(n4813), .Z(n4821) );
  XNOR U4805 ( .A(n4811), .B(n4820), .Z(n4813) );
  XNOR U4806 ( .A(n4822), .B(n4823), .Z(n4811) );
  AND U4807 ( .A(n245), .B(n4824), .Z(n4823) );
  XOR U4808 ( .A(p_input[208]), .B(n4822), .Z(n4824) );
  XNOR U4809 ( .A(n4825), .B(n4826), .Z(n4822) );
  AND U4810 ( .A(n249), .B(n4827), .Z(n4826) );
  XOR U4811 ( .A(n4828), .B(n4829), .Z(n4820) );
  AND U4812 ( .A(n253), .B(n4819), .Z(n4829) );
  XNOR U4813 ( .A(n4830), .B(n4817), .Z(n4819) );
  XOR U4814 ( .A(n4831), .B(n4832), .Z(n4817) );
  AND U4815 ( .A(n276), .B(n4833), .Z(n4832) );
  IV U4816 ( .A(n4828), .Z(n4830) );
  XOR U4817 ( .A(n4834), .B(n4835), .Z(n4828) );
  AND U4818 ( .A(n260), .B(n4827), .Z(n4835) );
  XNOR U4819 ( .A(n4825), .B(n4834), .Z(n4827) );
  XNOR U4820 ( .A(n4836), .B(n4837), .Z(n4825) );
  AND U4821 ( .A(n264), .B(n4838), .Z(n4837) );
  XOR U4822 ( .A(p_input[240]), .B(n4836), .Z(n4838) );
  XNOR U4823 ( .A(n4839), .B(n4840), .Z(n4836) );
  AND U4824 ( .A(n268), .B(n4841), .Z(n4840) );
  XOR U4825 ( .A(n4842), .B(n4843), .Z(n4834) );
  AND U4826 ( .A(n272), .B(n4833), .Z(n4843) );
  XNOR U4827 ( .A(n4844), .B(n4831), .Z(n4833) );
  XOR U4828 ( .A(n4845), .B(n4846), .Z(n4831) );
  AND U4829 ( .A(n295), .B(n4847), .Z(n4846) );
  IV U4830 ( .A(n4842), .Z(n4844) );
  XOR U4831 ( .A(n4848), .B(n4849), .Z(n4842) );
  AND U4832 ( .A(n279), .B(n4841), .Z(n4849) );
  XNOR U4833 ( .A(n4839), .B(n4848), .Z(n4841) );
  XNOR U4834 ( .A(n4850), .B(n4851), .Z(n4839) );
  AND U4835 ( .A(n283), .B(n4852), .Z(n4851) );
  XOR U4836 ( .A(p_input[272]), .B(n4850), .Z(n4852) );
  XNOR U4837 ( .A(n4853), .B(n4854), .Z(n4850) );
  AND U4838 ( .A(n287), .B(n4855), .Z(n4854) );
  XOR U4839 ( .A(n4856), .B(n4857), .Z(n4848) );
  AND U4840 ( .A(n291), .B(n4847), .Z(n4857) );
  XNOR U4841 ( .A(n4858), .B(n4845), .Z(n4847) );
  XOR U4842 ( .A(n4859), .B(n4860), .Z(n4845) );
  AND U4843 ( .A(n314), .B(n4861), .Z(n4860) );
  IV U4844 ( .A(n4856), .Z(n4858) );
  XOR U4845 ( .A(n4862), .B(n4863), .Z(n4856) );
  AND U4846 ( .A(n298), .B(n4855), .Z(n4863) );
  XNOR U4847 ( .A(n4853), .B(n4862), .Z(n4855) );
  XNOR U4848 ( .A(n4864), .B(n4865), .Z(n4853) );
  AND U4849 ( .A(n302), .B(n4866), .Z(n4865) );
  XOR U4850 ( .A(p_input[304]), .B(n4864), .Z(n4866) );
  XNOR U4851 ( .A(n4867), .B(n4868), .Z(n4864) );
  AND U4852 ( .A(n306), .B(n4869), .Z(n4868) );
  XOR U4853 ( .A(n4870), .B(n4871), .Z(n4862) );
  AND U4854 ( .A(n310), .B(n4861), .Z(n4871) );
  XNOR U4855 ( .A(n4872), .B(n4859), .Z(n4861) );
  XOR U4856 ( .A(n4873), .B(n4874), .Z(n4859) );
  AND U4857 ( .A(n333), .B(n4875), .Z(n4874) );
  IV U4858 ( .A(n4870), .Z(n4872) );
  XOR U4859 ( .A(n4876), .B(n4877), .Z(n4870) );
  AND U4860 ( .A(n317), .B(n4869), .Z(n4877) );
  XNOR U4861 ( .A(n4867), .B(n4876), .Z(n4869) );
  XNOR U4862 ( .A(n4878), .B(n4879), .Z(n4867) );
  AND U4863 ( .A(n321), .B(n4880), .Z(n4879) );
  XOR U4864 ( .A(p_input[336]), .B(n4878), .Z(n4880) );
  XNOR U4865 ( .A(n4881), .B(n4882), .Z(n4878) );
  AND U4866 ( .A(n325), .B(n4883), .Z(n4882) );
  XOR U4867 ( .A(n4884), .B(n4885), .Z(n4876) );
  AND U4868 ( .A(n329), .B(n4875), .Z(n4885) );
  XNOR U4869 ( .A(n4886), .B(n4873), .Z(n4875) );
  XOR U4870 ( .A(n4887), .B(n4888), .Z(n4873) );
  AND U4871 ( .A(n352), .B(n4889), .Z(n4888) );
  IV U4872 ( .A(n4884), .Z(n4886) );
  XOR U4873 ( .A(n4890), .B(n4891), .Z(n4884) );
  AND U4874 ( .A(n336), .B(n4883), .Z(n4891) );
  XNOR U4875 ( .A(n4881), .B(n4890), .Z(n4883) );
  XNOR U4876 ( .A(n4892), .B(n4893), .Z(n4881) );
  AND U4877 ( .A(n340), .B(n4894), .Z(n4893) );
  XOR U4878 ( .A(p_input[368]), .B(n4892), .Z(n4894) );
  XNOR U4879 ( .A(n4895), .B(n4896), .Z(n4892) );
  AND U4880 ( .A(n344), .B(n4897), .Z(n4896) );
  XOR U4881 ( .A(n4898), .B(n4899), .Z(n4890) );
  AND U4882 ( .A(n348), .B(n4889), .Z(n4899) );
  XNOR U4883 ( .A(n4900), .B(n4887), .Z(n4889) );
  XOR U4884 ( .A(n4901), .B(n4902), .Z(n4887) );
  AND U4885 ( .A(n370), .B(n4903), .Z(n4902) );
  IV U4886 ( .A(n4898), .Z(n4900) );
  XOR U4887 ( .A(n4904), .B(n4905), .Z(n4898) );
  AND U4888 ( .A(n355), .B(n4897), .Z(n4905) );
  XNOR U4889 ( .A(n4895), .B(n4904), .Z(n4897) );
  XNOR U4890 ( .A(n4906), .B(n4907), .Z(n4895) );
  AND U4891 ( .A(n359), .B(n4908), .Z(n4907) );
  XOR U4892 ( .A(p_input[400]), .B(n4906), .Z(n4908) );
  XOR U4893 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][16] ), .B(n4909), 
        .Z(n4906) );
  AND U4894 ( .A(n362), .B(n4910), .Z(n4909) );
  XOR U4895 ( .A(n4911), .B(n4912), .Z(n4904) );
  AND U4896 ( .A(n366), .B(n4903), .Z(n4912) );
  XNOR U4897 ( .A(n4913), .B(n4901), .Z(n4903) );
  XOR U4898 ( .A(\knn_comb_/min_val_out[0][16] ), .B(n4914), .Z(n4901) );
  AND U4899 ( .A(n378), .B(n4915), .Z(n4914) );
  IV U4900 ( .A(n4911), .Z(n4913) );
  XOR U4901 ( .A(n4916), .B(n4917), .Z(n4911) );
  AND U4902 ( .A(n373), .B(n4910), .Z(n4917) );
  XOR U4903 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][16] ), .B(n4916), 
        .Z(n4910) );
  XOR U4904 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .B(n4918), 
        .Z(n4916) );
  AND U4905 ( .A(n375), .B(n4915), .Z(n4918) );
  XOR U4906 ( .A(n4919), .B(n4920), .Z(n4915) );
  IV U4907 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .Z(n4920) );
  IV U4908 ( .A(\knn_comb_/min_val_out[0][16] ), .Z(n4919) );
  XOR U4909 ( .A(n109), .B(n4921), .Z(o[15]) );
  AND U4910 ( .A(n122), .B(n4922), .Z(n109) );
  XOR U4911 ( .A(n110), .B(n4921), .Z(n4922) );
  XOR U4912 ( .A(n4923), .B(n4924), .Z(n4921) );
  AND U4913 ( .A(n142), .B(n4925), .Z(n4924) );
  XOR U4914 ( .A(n4926), .B(n39), .Z(n110) );
  AND U4915 ( .A(n125), .B(n4927), .Z(n39) );
  XOR U4916 ( .A(n40), .B(n4926), .Z(n4927) );
  XOR U4917 ( .A(n4928), .B(n4929), .Z(n40) );
  AND U4918 ( .A(n130), .B(n4930), .Z(n4929) );
  XOR U4919 ( .A(p_input[15]), .B(n4928), .Z(n4930) );
  XNOR U4920 ( .A(n4931), .B(n4932), .Z(n4928) );
  AND U4921 ( .A(n134), .B(n4933), .Z(n4932) );
  XOR U4922 ( .A(n4934), .B(n4935), .Z(n4926) );
  AND U4923 ( .A(n138), .B(n4925), .Z(n4935) );
  XNOR U4924 ( .A(n4936), .B(n4923), .Z(n4925) );
  XOR U4925 ( .A(n4937), .B(n4938), .Z(n4923) );
  AND U4926 ( .A(n162), .B(n4939), .Z(n4938) );
  IV U4927 ( .A(n4934), .Z(n4936) );
  XOR U4928 ( .A(n4940), .B(n4941), .Z(n4934) );
  AND U4929 ( .A(n146), .B(n4933), .Z(n4941) );
  XNOR U4930 ( .A(n4931), .B(n4940), .Z(n4933) );
  XNOR U4931 ( .A(n4942), .B(n4943), .Z(n4931) );
  AND U4932 ( .A(n150), .B(n4944), .Z(n4943) );
  XOR U4933 ( .A(p_input[47]), .B(n4942), .Z(n4944) );
  XNOR U4934 ( .A(n4945), .B(n4946), .Z(n4942) );
  AND U4935 ( .A(n154), .B(n4947), .Z(n4946) );
  XOR U4936 ( .A(n4948), .B(n4949), .Z(n4940) );
  AND U4937 ( .A(n158), .B(n4939), .Z(n4949) );
  XNOR U4938 ( .A(n4950), .B(n4937), .Z(n4939) );
  XOR U4939 ( .A(n4951), .B(n4952), .Z(n4937) );
  AND U4940 ( .A(n181), .B(n4953), .Z(n4952) );
  IV U4941 ( .A(n4948), .Z(n4950) );
  XOR U4942 ( .A(n4954), .B(n4955), .Z(n4948) );
  AND U4943 ( .A(n165), .B(n4947), .Z(n4955) );
  XNOR U4944 ( .A(n4945), .B(n4954), .Z(n4947) );
  XNOR U4945 ( .A(n4956), .B(n4957), .Z(n4945) );
  AND U4946 ( .A(n169), .B(n4958), .Z(n4957) );
  XOR U4947 ( .A(p_input[79]), .B(n4956), .Z(n4958) );
  XNOR U4948 ( .A(n4959), .B(n4960), .Z(n4956) );
  AND U4949 ( .A(n173), .B(n4961), .Z(n4960) );
  XOR U4950 ( .A(n4962), .B(n4963), .Z(n4954) );
  AND U4951 ( .A(n177), .B(n4953), .Z(n4963) );
  XNOR U4952 ( .A(n4964), .B(n4951), .Z(n4953) );
  XOR U4953 ( .A(n4965), .B(n4966), .Z(n4951) );
  AND U4954 ( .A(n200), .B(n4967), .Z(n4966) );
  IV U4955 ( .A(n4962), .Z(n4964) );
  XOR U4956 ( .A(n4968), .B(n4969), .Z(n4962) );
  AND U4957 ( .A(n184), .B(n4961), .Z(n4969) );
  XNOR U4958 ( .A(n4959), .B(n4968), .Z(n4961) );
  XNOR U4959 ( .A(n4970), .B(n4971), .Z(n4959) );
  AND U4960 ( .A(n188), .B(n4972), .Z(n4971) );
  XOR U4961 ( .A(p_input[111]), .B(n4970), .Z(n4972) );
  XNOR U4962 ( .A(n4973), .B(n4974), .Z(n4970) );
  AND U4963 ( .A(n192), .B(n4975), .Z(n4974) );
  XOR U4964 ( .A(n4976), .B(n4977), .Z(n4968) );
  AND U4965 ( .A(n196), .B(n4967), .Z(n4977) );
  XNOR U4966 ( .A(n4978), .B(n4965), .Z(n4967) );
  XOR U4967 ( .A(n4979), .B(n4980), .Z(n4965) );
  AND U4968 ( .A(n219), .B(n4981), .Z(n4980) );
  IV U4969 ( .A(n4976), .Z(n4978) );
  XOR U4970 ( .A(n4982), .B(n4983), .Z(n4976) );
  AND U4971 ( .A(n203), .B(n4975), .Z(n4983) );
  XNOR U4972 ( .A(n4973), .B(n4982), .Z(n4975) );
  XNOR U4973 ( .A(n4984), .B(n4985), .Z(n4973) );
  AND U4974 ( .A(n207), .B(n4986), .Z(n4985) );
  XOR U4975 ( .A(p_input[143]), .B(n4984), .Z(n4986) );
  XNOR U4976 ( .A(n4987), .B(n4988), .Z(n4984) );
  AND U4977 ( .A(n211), .B(n4989), .Z(n4988) );
  XOR U4978 ( .A(n4990), .B(n4991), .Z(n4982) );
  AND U4979 ( .A(n215), .B(n4981), .Z(n4991) );
  XNOR U4980 ( .A(n4992), .B(n4979), .Z(n4981) );
  XOR U4981 ( .A(n4993), .B(n4994), .Z(n4979) );
  AND U4982 ( .A(n238), .B(n4995), .Z(n4994) );
  IV U4983 ( .A(n4990), .Z(n4992) );
  XOR U4984 ( .A(n4996), .B(n4997), .Z(n4990) );
  AND U4985 ( .A(n222), .B(n4989), .Z(n4997) );
  XNOR U4986 ( .A(n4987), .B(n4996), .Z(n4989) );
  XNOR U4987 ( .A(n4998), .B(n4999), .Z(n4987) );
  AND U4988 ( .A(n226), .B(n5000), .Z(n4999) );
  XOR U4989 ( .A(p_input[175]), .B(n4998), .Z(n5000) );
  XNOR U4990 ( .A(n5001), .B(n5002), .Z(n4998) );
  AND U4991 ( .A(n230), .B(n5003), .Z(n5002) );
  XOR U4992 ( .A(n5004), .B(n5005), .Z(n4996) );
  AND U4993 ( .A(n234), .B(n4995), .Z(n5005) );
  XNOR U4994 ( .A(n5006), .B(n4993), .Z(n4995) );
  XOR U4995 ( .A(n5007), .B(n5008), .Z(n4993) );
  AND U4996 ( .A(n257), .B(n5009), .Z(n5008) );
  IV U4997 ( .A(n5004), .Z(n5006) );
  XOR U4998 ( .A(n5010), .B(n5011), .Z(n5004) );
  AND U4999 ( .A(n241), .B(n5003), .Z(n5011) );
  XNOR U5000 ( .A(n5001), .B(n5010), .Z(n5003) );
  XNOR U5001 ( .A(n5012), .B(n5013), .Z(n5001) );
  AND U5002 ( .A(n245), .B(n5014), .Z(n5013) );
  XOR U5003 ( .A(p_input[207]), .B(n5012), .Z(n5014) );
  XNOR U5004 ( .A(n5015), .B(n5016), .Z(n5012) );
  AND U5005 ( .A(n249), .B(n5017), .Z(n5016) );
  XOR U5006 ( .A(n5018), .B(n5019), .Z(n5010) );
  AND U5007 ( .A(n253), .B(n5009), .Z(n5019) );
  XNOR U5008 ( .A(n5020), .B(n5007), .Z(n5009) );
  XOR U5009 ( .A(n5021), .B(n5022), .Z(n5007) );
  AND U5010 ( .A(n276), .B(n5023), .Z(n5022) );
  IV U5011 ( .A(n5018), .Z(n5020) );
  XOR U5012 ( .A(n5024), .B(n5025), .Z(n5018) );
  AND U5013 ( .A(n260), .B(n5017), .Z(n5025) );
  XNOR U5014 ( .A(n5015), .B(n5024), .Z(n5017) );
  XNOR U5015 ( .A(n5026), .B(n5027), .Z(n5015) );
  AND U5016 ( .A(n264), .B(n5028), .Z(n5027) );
  XOR U5017 ( .A(p_input[239]), .B(n5026), .Z(n5028) );
  XNOR U5018 ( .A(n5029), .B(n5030), .Z(n5026) );
  AND U5019 ( .A(n268), .B(n5031), .Z(n5030) );
  XOR U5020 ( .A(n5032), .B(n5033), .Z(n5024) );
  AND U5021 ( .A(n272), .B(n5023), .Z(n5033) );
  XNOR U5022 ( .A(n5034), .B(n5021), .Z(n5023) );
  XOR U5023 ( .A(n5035), .B(n5036), .Z(n5021) );
  AND U5024 ( .A(n295), .B(n5037), .Z(n5036) );
  IV U5025 ( .A(n5032), .Z(n5034) );
  XOR U5026 ( .A(n5038), .B(n5039), .Z(n5032) );
  AND U5027 ( .A(n279), .B(n5031), .Z(n5039) );
  XNOR U5028 ( .A(n5029), .B(n5038), .Z(n5031) );
  XNOR U5029 ( .A(n5040), .B(n5041), .Z(n5029) );
  AND U5030 ( .A(n283), .B(n5042), .Z(n5041) );
  XOR U5031 ( .A(p_input[271]), .B(n5040), .Z(n5042) );
  XNOR U5032 ( .A(n5043), .B(n5044), .Z(n5040) );
  AND U5033 ( .A(n287), .B(n5045), .Z(n5044) );
  XOR U5034 ( .A(n5046), .B(n5047), .Z(n5038) );
  AND U5035 ( .A(n291), .B(n5037), .Z(n5047) );
  XNOR U5036 ( .A(n5048), .B(n5035), .Z(n5037) );
  XOR U5037 ( .A(n5049), .B(n5050), .Z(n5035) );
  AND U5038 ( .A(n314), .B(n5051), .Z(n5050) );
  IV U5039 ( .A(n5046), .Z(n5048) );
  XOR U5040 ( .A(n5052), .B(n5053), .Z(n5046) );
  AND U5041 ( .A(n298), .B(n5045), .Z(n5053) );
  XNOR U5042 ( .A(n5043), .B(n5052), .Z(n5045) );
  XNOR U5043 ( .A(n5054), .B(n5055), .Z(n5043) );
  AND U5044 ( .A(n302), .B(n5056), .Z(n5055) );
  XOR U5045 ( .A(p_input[303]), .B(n5054), .Z(n5056) );
  XNOR U5046 ( .A(n5057), .B(n5058), .Z(n5054) );
  AND U5047 ( .A(n306), .B(n5059), .Z(n5058) );
  XOR U5048 ( .A(n5060), .B(n5061), .Z(n5052) );
  AND U5049 ( .A(n310), .B(n5051), .Z(n5061) );
  XNOR U5050 ( .A(n5062), .B(n5049), .Z(n5051) );
  XOR U5051 ( .A(n5063), .B(n5064), .Z(n5049) );
  AND U5052 ( .A(n333), .B(n5065), .Z(n5064) );
  IV U5053 ( .A(n5060), .Z(n5062) );
  XOR U5054 ( .A(n5066), .B(n5067), .Z(n5060) );
  AND U5055 ( .A(n317), .B(n5059), .Z(n5067) );
  XNOR U5056 ( .A(n5057), .B(n5066), .Z(n5059) );
  XNOR U5057 ( .A(n5068), .B(n5069), .Z(n5057) );
  AND U5058 ( .A(n321), .B(n5070), .Z(n5069) );
  XOR U5059 ( .A(p_input[335]), .B(n5068), .Z(n5070) );
  XNOR U5060 ( .A(n5071), .B(n5072), .Z(n5068) );
  AND U5061 ( .A(n325), .B(n5073), .Z(n5072) );
  XOR U5062 ( .A(n5074), .B(n5075), .Z(n5066) );
  AND U5063 ( .A(n329), .B(n5065), .Z(n5075) );
  XNOR U5064 ( .A(n5076), .B(n5063), .Z(n5065) );
  XOR U5065 ( .A(n5077), .B(n5078), .Z(n5063) );
  AND U5066 ( .A(n352), .B(n5079), .Z(n5078) );
  IV U5067 ( .A(n5074), .Z(n5076) );
  XOR U5068 ( .A(n5080), .B(n5081), .Z(n5074) );
  AND U5069 ( .A(n336), .B(n5073), .Z(n5081) );
  XNOR U5070 ( .A(n5071), .B(n5080), .Z(n5073) );
  XNOR U5071 ( .A(n5082), .B(n5083), .Z(n5071) );
  AND U5072 ( .A(n340), .B(n5084), .Z(n5083) );
  XOR U5073 ( .A(p_input[367]), .B(n5082), .Z(n5084) );
  XNOR U5074 ( .A(n5085), .B(n5086), .Z(n5082) );
  AND U5075 ( .A(n344), .B(n5087), .Z(n5086) );
  XOR U5076 ( .A(n5088), .B(n5089), .Z(n5080) );
  AND U5077 ( .A(n348), .B(n5079), .Z(n5089) );
  XNOR U5078 ( .A(n5090), .B(n5077), .Z(n5079) );
  XOR U5079 ( .A(n5091), .B(n5092), .Z(n5077) );
  AND U5080 ( .A(n370), .B(n5093), .Z(n5092) );
  IV U5081 ( .A(n5088), .Z(n5090) );
  XOR U5082 ( .A(n5094), .B(n5095), .Z(n5088) );
  AND U5083 ( .A(n355), .B(n5087), .Z(n5095) );
  XNOR U5084 ( .A(n5085), .B(n5094), .Z(n5087) );
  XNOR U5085 ( .A(n5096), .B(n5097), .Z(n5085) );
  AND U5086 ( .A(n359), .B(n5098), .Z(n5097) );
  XOR U5087 ( .A(p_input[399]), .B(n5096), .Z(n5098) );
  XOR U5088 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n5099), 
        .Z(n5096) );
  AND U5089 ( .A(n362), .B(n5100), .Z(n5099) );
  XOR U5090 ( .A(n5101), .B(n5102), .Z(n5094) );
  AND U5091 ( .A(n366), .B(n5093), .Z(n5102) );
  XNOR U5092 ( .A(n5103), .B(n5091), .Z(n5093) );
  XOR U5093 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n5104), .Z(n5091) );
  AND U5094 ( .A(n378), .B(n5105), .Z(n5104) );
  IV U5095 ( .A(n5101), .Z(n5103) );
  XOR U5096 ( .A(n5106), .B(n5107), .Z(n5101) );
  AND U5097 ( .A(n373), .B(n5100), .Z(n5107) );
  XOR U5098 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n5106), 
        .Z(n5100) );
  XOR U5099 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(n5108), 
        .Z(n5106) );
  AND U5100 ( .A(n375), .B(n5105), .Z(n5108) );
  XOR U5101 ( .A(n5109), .B(n5110), .Z(n5105) );
  IV U5102 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .Z(n5110) );
  IV U5103 ( .A(\knn_comb_/min_val_out[0][15] ), .Z(n5109) );
  XOR U5104 ( .A(n111), .B(n5111), .Z(o[14]) );
  AND U5105 ( .A(n122), .B(n5112), .Z(n111) );
  XOR U5106 ( .A(n112), .B(n5111), .Z(n5112) );
  XOR U5107 ( .A(n5113), .B(n5114), .Z(n5111) );
  AND U5108 ( .A(n142), .B(n5115), .Z(n5114) );
  XOR U5109 ( .A(n5116), .B(n41), .Z(n112) );
  AND U5110 ( .A(n125), .B(n5117), .Z(n41) );
  XOR U5111 ( .A(n42), .B(n5116), .Z(n5117) );
  XOR U5112 ( .A(n5118), .B(n5119), .Z(n42) );
  AND U5113 ( .A(n130), .B(n5120), .Z(n5119) );
  XOR U5114 ( .A(p_input[14]), .B(n5118), .Z(n5120) );
  XNOR U5115 ( .A(n5121), .B(n5122), .Z(n5118) );
  AND U5116 ( .A(n134), .B(n5123), .Z(n5122) );
  XOR U5117 ( .A(n5124), .B(n5125), .Z(n5116) );
  AND U5118 ( .A(n138), .B(n5115), .Z(n5125) );
  XNOR U5119 ( .A(n5126), .B(n5113), .Z(n5115) );
  XOR U5120 ( .A(n5127), .B(n5128), .Z(n5113) );
  AND U5121 ( .A(n162), .B(n5129), .Z(n5128) );
  IV U5122 ( .A(n5124), .Z(n5126) );
  XOR U5123 ( .A(n5130), .B(n5131), .Z(n5124) );
  AND U5124 ( .A(n146), .B(n5123), .Z(n5131) );
  XNOR U5125 ( .A(n5121), .B(n5130), .Z(n5123) );
  XNOR U5126 ( .A(n5132), .B(n5133), .Z(n5121) );
  AND U5127 ( .A(n150), .B(n5134), .Z(n5133) );
  XOR U5128 ( .A(p_input[46]), .B(n5132), .Z(n5134) );
  XNOR U5129 ( .A(n5135), .B(n5136), .Z(n5132) );
  AND U5130 ( .A(n154), .B(n5137), .Z(n5136) );
  XOR U5131 ( .A(n5138), .B(n5139), .Z(n5130) );
  AND U5132 ( .A(n158), .B(n5129), .Z(n5139) );
  XNOR U5133 ( .A(n5140), .B(n5127), .Z(n5129) );
  XOR U5134 ( .A(n5141), .B(n5142), .Z(n5127) );
  AND U5135 ( .A(n181), .B(n5143), .Z(n5142) );
  IV U5136 ( .A(n5138), .Z(n5140) );
  XOR U5137 ( .A(n5144), .B(n5145), .Z(n5138) );
  AND U5138 ( .A(n165), .B(n5137), .Z(n5145) );
  XNOR U5139 ( .A(n5135), .B(n5144), .Z(n5137) );
  XNOR U5140 ( .A(n5146), .B(n5147), .Z(n5135) );
  AND U5141 ( .A(n169), .B(n5148), .Z(n5147) );
  XOR U5142 ( .A(p_input[78]), .B(n5146), .Z(n5148) );
  XNOR U5143 ( .A(n5149), .B(n5150), .Z(n5146) );
  AND U5144 ( .A(n173), .B(n5151), .Z(n5150) );
  XOR U5145 ( .A(n5152), .B(n5153), .Z(n5144) );
  AND U5146 ( .A(n177), .B(n5143), .Z(n5153) );
  XNOR U5147 ( .A(n5154), .B(n5141), .Z(n5143) );
  XOR U5148 ( .A(n5155), .B(n5156), .Z(n5141) );
  AND U5149 ( .A(n200), .B(n5157), .Z(n5156) );
  IV U5150 ( .A(n5152), .Z(n5154) );
  XOR U5151 ( .A(n5158), .B(n5159), .Z(n5152) );
  AND U5152 ( .A(n184), .B(n5151), .Z(n5159) );
  XNOR U5153 ( .A(n5149), .B(n5158), .Z(n5151) );
  XNOR U5154 ( .A(n5160), .B(n5161), .Z(n5149) );
  AND U5155 ( .A(n188), .B(n5162), .Z(n5161) );
  XOR U5156 ( .A(p_input[110]), .B(n5160), .Z(n5162) );
  XNOR U5157 ( .A(n5163), .B(n5164), .Z(n5160) );
  AND U5158 ( .A(n192), .B(n5165), .Z(n5164) );
  XOR U5159 ( .A(n5166), .B(n5167), .Z(n5158) );
  AND U5160 ( .A(n196), .B(n5157), .Z(n5167) );
  XNOR U5161 ( .A(n5168), .B(n5155), .Z(n5157) );
  XOR U5162 ( .A(n5169), .B(n5170), .Z(n5155) );
  AND U5163 ( .A(n219), .B(n5171), .Z(n5170) );
  IV U5164 ( .A(n5166), .Z(n5168) );
  XOR U5165 ( .A(n5172), .B(n5173), .Z(n5166) );
  AND U5166 ( .A(n203), .B(n5165), .Z(n5173) );
  XNOR U5167 ( .A(n5163), .B(n5172), .Z(n5165) );
  XNOR U5168 ( .A(n5174), .B(n5175), .Z(n5163) );
  AND U5169 ( .A(n207), .B(n5176), .Z(n5175) );
  XOR U5170 ( .A(p_input[142]), .B(n5174), .Z(n5176) );
  XNOR U5171 ( .A(n5177), .B(n5178), .Z(n5174) );
  AND U5172 ( .A(n211), .B(n5179), .Z(n5178) );
  XOR U5173 ( .A(n5180), .B(n5181), .Z(n5172) );
  AND U5174 ( .A(n215), .B(n5171), .Z(n5181) );
  XNOR U5175 ( .A(n5182), .B(n5169), .Z(n5171) );
  XOR U5176 ( .A(n5183), .B(n5184), .Z(n5169) );
  AND U5177 ( .A(n238), .B(n5185), .Z(n5184) );
  IV U5178 ( .A(n5180), .Z(n5182) );
  XOR U5179 ( .A(n5186), .B(n5187), .Z(n5180) );
  AND U5180 ( .A(n222), .B(n5179), .Z(n5187) );
  XNOR U5181 ( .A(n5177), .B(n5186), .Z(n5179) );
  XNOR U5182 ( .A(n5188), .B(n5189), .Z(n5177) );
  AND U5183 ( .A(n226), .B(n5190), .Z(n5189) );
  XOR U5184 ( .A(p_input[174]), .B(n5188), .Z(n5190) );
  XNOR U5185 ( .A(n5191), .B(n5192), .Z(n5188) );
  AND U5186 ( .A(n230), .B(n5193), .Z(n5192) );
  XOR U5187 ( .A(n5194), .B(n5195), .Z(n5186) );
  AND U5188 ( .A(n234), .B(n5185), .Z(n5195) );
  XNOR U5189 ( .A(n5196), .B(n5183), .Z(n5185) );
  XOR U5190 ( .A(n5197), .B(n5198), .Z(n5183) );
  AND U5191 ( .A(n257), .B(n5199), .Z(n5198) );
  IV U5192 ( .A(n5194), .Z(n5196) );
  XOR U5193 ( .A(n5200), .B(n5201), .Z(n5194) );
  AND U5194 ( .A(n241), .B(n5193), .Z(n5201) );
  XNOR U5195 ( .A(n5191), .B(n5200), .Z(n5193) );
  XNOR U5196 ( .A(n5202), .B(n5203), .Z(n5191) );
  AND U5197 ( .A(n245), .B(n5204), .Z(n5203) );
  XOR U5198 ( .A(p_input[206]), .B(n5202), .Z(n5204) );
  XNOR U5199 ( .A(n5205), .B(n5206), .Z(n5202) );
  AND U5200 ( .A(n249), .B(n5207), .Z(n5206) );
  XOR U5201 ( .A(n5208), .B(n5209), .Z(n5200) );
  AND U5202 ( .A(n253), .B(n5199), .Z(n5209) );
  XNOR U5203 ( .A(n5210), .B(n5197), .Z(n5199) );
  XOR U5204 ( .A(n5211), .B(n5212), .Z(n5197) );
  AND U5205 ( .A(n276), .B(n5213), .Z(n5212) );
  IV U5206 ( .A(n5208), .Z(n5210) );
  XOR U5207 ( .A(n5214), .B(n5215), .Z(n5208) );
  AND U5208 ( .A(n260), .B(n5207), .Z(n5215) );
  XNOR U5209 ( .A(n5205), .B(n5214), .Z(n5207) );
  XNOR U5210 ( .A(n5216), .B(n5217), .Z(n5205) );
  AND U5211 ( .A(n264), .B(n5218), .Z(n5217) );
  XOR U5212 ( .A(p_input[238]), .B(n5216), .Z(n5218) );
  XNOR U5213 ( .A(n5219), .B(n5220), .Z(n5216) );
  AND U5214 ( .A(n268), .B(n5221), .Z(n5220) );
  XOR U5215 ( .A(n5222), .B(n5223), .Z(n5214) );
  AND U5216 ( .A(n272), .B(n5213), .Z(n5223) );
  XNOR U5217 ( .A(n5224), .B(n5211), .Z(n5213) );
  XOR U5218 ( .A(n5225), .B(n5226), .Z(n5211) );
  AND U5219 ( .A(n295), .B(n5227), .Z(n5226) );
  IV U5220 ( .A(n5222), .Z(n5224) );
  XOR U5221 ( .A(n5228), .B(n5229), .Z(n5222) );
  AND U5222 ( .A(n279), .B(n5221), .Z(n5229) );
  XNOR U5223 ( .A(n5219), .B(n5228), .Z(n5221) );
  XNOR U5224 ( .A(n5230), .B(n5231), .Z(n5219) );
  AND U5225 ( .A(n283), .B(n5232), .Z(n5231) );
  XOR U5226 ( .A(p_input[270]), .B(n5230), .Z(n5232) );
  XNOR U5227 ( .A(n5233), .B(n5234), .Z(n5230) );
  AND U5228 ( .A(n287), .B(n5235), .Z(n5234) );
  XOR U5229 ( .A(n5236), .B(n5237), .Z(n5228) );
  AND U5230 ( .A(n291), .B(n5227), .Z(n5237) );
  XNOR U5231 ( .A(n5238), .B(n5225), .Z(n5227) );
  XOR U5232 ( .A(n5239), .B(n5240), .Z(n5225) );
  AND U5233 ( .A(n314), .B(n5241), .Z(n5240) );
  IV U5234 ( .A(n5236), .Z(n5238) );
  XOR U5235 ( .A(n5242), .B(n5243), .Z(n5236) );
  AND U5236 ( .A(n298), .B(n5235), .Z(n5243) );
  XNOR U5237 ( .A(n5233), .B(n5242), .Z(n5235) );
  XNOR U5238 ( .A(n5244), .B(n5245), .Z(n5233) );
  AND U5239 ( .A(n302), .B(n5246), .Z(n5245) );
  XOR U5240 ( .A(p_input[302]), .B(n5244), .Z(n5246) );
  XNOR U5241 ( .A(n5247), .B(n5248), .Z(n5244) );
  AND U5242 ( .A(n306), .B(n5249), .Z(n5248) );
  XOR U5243 ( .A(n5250), .B(n5251), .Z(n5242) );
  AND U5244 ( .A(n310), .B(n5241), .Z(n5251) );
  XNOR U5245 ( .A(n5252), .B(n5239), .Z(n5241) );
  XOR U5246 ( .A(n5253), .B(n5254), .Z(n5239) );
  AND U5247 ( .A(n333), .B(n5255), .Z(n5254) );
  IV U5248 ( .A(n5250), .Z(n5252) );
  XOR U5249 ( .A(n5256), .B(n5257), .Z(n5250) );
  AND U5250 ( .A(n317), .B(n5249), .Z(n5257) );
  XNOR U5251 ( .A(n5247), .B(n5256), .Z(n5249) );
  XNOR U5252 ( .A(n5258), .B(n5259), .Z(n5247) );
  AND U5253 ( .A(n321), .B(n5260), .Z(n5259) );
  XOR U5254 ( .A(p_input[334]), .B(n5258), .Z(n5260) );
  XNOR U5255 ( .A(n5261), .B(n5262), .Z(n5258) );
  AND U5256 ( .A(n325), .B(n5263), .Z(n5262) );
  XOR U5257 ( .A(n5264), .B(n5265), .Z(n5256) );
  AND U5258 ( .A(n329), .B(n5255), .Z(n5265) );
  XNOR U5259 ( .A(n5266), .B(n5253), .Z(n5255) );
  XOR U5260 ( .A(n5267), .B(n5268), .Z(n5253) );
  AND U5261 ( .A(n352), .B(n5269), .Z(n5268) );
  IV U5262 ( .A(n5264), .Z(n5266) );
  XOR U5263 ( .A(n5270), .B(n5271), .Z(n5264) );
  AND U5264 ( .A(n336), .B(n5263), .Z(n5271) );
  XNOR U5265 ( .A(n5261), .B(n5270), .Z(n5263) );
  XNOR U5266 ( .A(n5272), .B(n5273), .Z(n5261) );
  AND U5267 ( .A(n340), .B(n5274), .Z(n5273) );
  XOR U5268 ( .A(p_input[366]), .B(n5272), .Z(n5274) );
  XNOR U5269 ( .A(n5275), .B(n5276), .Z(n5272) );
  AND U5270 ( .A(n344), .B(n5277), .Z(n5276) );
  XOR U5271 ( .A(n5278), .B(n5279), .Z(n5270) );
  AND U5272 ( .A(n348), .B(n5269), .Z(n5279) );
  XNOR U5273 ( .A(n5280), .B(n5267), .Z(n5269) );
  XOR U5274 ( .A(n5281), .B(n5282), .Z(n5267) );
  AND U5275 ( .A(n370), .B(n5283), .Z(n5282) );
  IV U5276 ( .A(n5278), .Z(n5280) );
  XOR U5277 ( .A(n5284), .B(n5285), .Z(n5278) );
  AND U5278 ( .A(n355), .B(n5277), .Z(n5285) );
  XNOR U5279 ( .A(n5275), .B(n5284), .Z(n5277) );
  XNOR U5280 ( .A(n5286), .B(n5287), .Z(n5275) );
  AND U5281 ( .A(n359), .B(n5288), .Z(n5287) );
  XOR U5282 ( .A(p_input[398]), .B(n5286), .Z(n5288) );
  XOR U5283 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n5289), 
        .Z(n5286) );
  AND U5284 ( .A(n362), .B(n5290), .Z(n5289) );
  XOR U5285 ( .A(n5291), .B(n5292), .Z(n5284) );
  AND U5286 ( .A(n366), .B(n5283), .Z(n5292) );
  XNOR U5287 ( .A(n5293), .B(n5281), .Z(n5283) );
  XOR U5288 ( .A(\knn_comb_/min_val_out[0][14] ), .B(n5294), .Z(n5281) );
  AND U5289 ( .A(n378), .B(n5295), .Z(n5294) );
  IV U5290 ( .A(n5291), .Z(n5293) );
  XOR U5291 ( .A(n5296), .B(n5297), .Z(n5291) );
  AND U5292 ( .A(n373), .B(n5290), .Z(n5297) );
  XOR U5293 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(n5296), 
        .Z(n5290) );
  XOR U5294 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(n5298), 
        .Z(n5296) );
  AND U5295 ( .A(n375), .B(n5295), .Z(n5298) );
  XOR U5296 ( .A(\knn_comb_/min_val_out[0][14] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .Z(n5295) );
  XOR U5297 ( .A(n113), .B(n5299), .Z(o[13]) );
  AND U5298 ( .A(n122), .B(n5300), .Z(n113) );
  XOR U5299 ( .A(n114), .B(n5299), .Z(n5300) );
  XOR U5300 ( .A(n5301), .B(n5302), .Z(n5299) );
  AND U5301 ( .A(n142), .B(n5303), .Z(n5302) );
  XOR U5302 ( .A(n5304), .B(n43), .Z(n114) );
  AND U5303 ( .A(n125), .B(n5305), .Z(n43) );
  XOR U5304 ( .A(n44), .B(n5304), .Z(n5305) );
  XOR U5305 ( .A(n5306), .B(n5307), .Z(n44) );
  AND U5306 ( .A(n130), .B(n5308), .Z(n5307) );
  XOR U5307 ( .A(p_input[13]), .B(n5306), .Z(n5308) );
  XNOR U5308 ( .A(n5309), .B(n5310), .Z(n5306) );
  AND U5309 ( .A(n134), .B(n5311), .Z(n5310) );
  XOR U5310 ( .A(n5312), .B(n5313), .Z(n5304) );
  AND U5311 ( .A(n138), .B(n5303), .Z(n5313) );
  XNOR U5312 ( .A(n5314), .B(n5301), .Z(n5303) );
  XOR U5313 ( .A(n5315), .B(n5316), .Z(n5301) );
  AND U5314 ( .A(n162), .B(n5317), .Z(n5316) );
  IV U5315 ( .A(n5312), .Z(n5314) );
  XOR U5316 ( .A(n5318), .B(n5319), .Z(n5312) );
  AND U5317 ( .A(n146), .B(n5311), .Z(n5319) );
  XNOR U5318 ( .A(n5309), .B(n5318), .Z(n5311) );
  XNOR U5319 ( .A(n5320), .B(n5321), .Z(n5309) );
  AND U5320 ( .A(n150), .B(n5322), .Z(n5321) );
  XOR U5321 ( .A(p_input[45]), .B(n5320), .Z(n5322) );
  XNOR U5322 ( .A(n5323), .B(n5324), .Z(n5320) );
  AND U5323 ( .A(n154), .B(n5325), .Z(n5324) );
  XOR U5324 ( .A(n5326), .B(n5327), .Z(n5318) );
  AND U5325 ( .A(n158), .B(n5317), .Z(n5327) );
  XNOR U5326 ( .A(n5328), .B(n5315), .Z(n5317) );
  XOR U5327 ( .A(n5329), .B(n5330), .Z(n5315) );
  AND U5328 ( .A(n181), .B(n5331), .Z(n5330) );
  IV U5329 ( .A(n5326), .Z(n5328) );
  XOR U5330 ( .A(n5332), .B(n5333), .Z(n5326) );
  AND U5331 ( .A(n165), .B(n5325), .Z(n5333) );
  XNOR U5332 ( .A(n5323), .B(n5332), .Z(n5325) );
  XNOR U5333 ( .A(n5334), .B(n5335), .Z(n5323) );
  AND U5334 ( .A(n169), .B(n5336), .Z(n5335) );
  XOR U5335 ( .A(p_input[77]), .B(n5334), .Z(n5336) );
  XNOR U5336 ( .A(n5337), .B(n5338), .Z(n5334) );
  AND U5337 ( .A(n173), .B(n5339), .Z(n5338) );
  XOR U5338 ( .A(n5340), .B(n5341), .Z(n5332) );
  AND U5339 ( .A(n177), .B(n5331), .Z(n5341) );
  XNOR U5340 ( .A(n5342), .B(n5329), .Z(n5331) );
  XOR U5341 ( .A(n5343), .B(n5344), .Z(n5329) );
  AND U5342 ( .A(n200), .B(n5345), .Z(n5344) );
  IV U5343 ( .A(n5340), .Z(n5342) );
  XOR U5344 ( .A(n5346), .B(n5347), .Z(n5340) );
  AND U5345 ( .A(n184), .B(n5339), .Z(n5347) );
  XNOR U5346 ( .A(n5337), .B(n5346), .Z(n5339) );
  XNOR U5347 ( .A(n5348), .B(n5349), .Z(n5337) );
  AND U5348 ( .A(n188), .B(n5350), .Z(n5349) );
  XOR U5349 ( .A(p_input[109]), .B(n5348), .Z(n5350) );
  XNOR U5350 ( .A(n5351), .B(n5352), .Z(n5348) );
  AND U5351 ( .A(n192), .B(n5353), .Z(n5352) );
  XOR U5352 ( .A(n5354), .B(n5355), .Z(n5346) );
  AND U5353 ( .A(n196), .B(n5345), .Z(n5355) );
  XNOR U5354 ( .A(n5356), .B(n5343), .Z(n5345) );
  XOR U5355 ( .A(n5357), .B(n5358), .Z(n5343) );
  AND U5356 ( .A(n219), .B(n5359), .Z(n5358) );
  IV U5357 ( .A(n5354), .Z(n5356) );
  XOR U5358 ( .A(n5360), .B(n5361), .Z(n5354) );
  AND U5359 ( .A(n203), .B(n5353), .Z(n5361) );
  XNOR U5360 ( .A(n5351), .B(n5360), .Z(n5353) );
  XNOR U5361 ( .A(n5362), .B(n5363), .Z(n5351) );
  AND U5362 ( .A(n207), .B(n5364), .Z(n5363) );
  XOR U5363 ( .A(p_input[141]), .B(n5362), .Z(n5364) );
  XNOR U5364 ( .A(n5365), .B(n5366), .Z(n5362) );
  AND U5365 ( .A(n211), .B(n5367), .Z(n5366) );
  XOR U5366 ( .A(n5368), .B(n5369), .Z(n5360) );
  AND U5367 ( .A(n215), .B(n5359), .Z(n5369) );
  XNOR U5368 ( .A(n5370), .B(n5357), .Z(n5359) );
  XOR U5369 ( .A(n5371), .B(n5372), .Z(n5357) );
  AND U5370 ( .A(n238), .B(n5373), .Z(n5372) );
  IV U5371 ( .A(n5368), .Z(n5370) );
  XOR U5372 ( .A(n5374), .B(n5375), .Z(n5368) );
  AND U5373 ( .A(n222), .B(n5367), .Z(n5375) );
  XNOR U5374 ( .A(n5365), .B(n5374), .Z(n5367) );
  XNOR U5375 ( .A(n5376), .B(n5377), .Z(n5365) );
  AND U5376 ( .A(n226), .B(n5378), .Z(n5377) );
  XOR U5377 ( .A(p_input[173]), .B(n5376), .Z(n5378) );
  XNOR U5378 ( .A(n5379), .B(n5380), .Z(n5376) );
  AND U5379 ( .A(n230), .B(n5381), .Z(n5380) );
  XOR U5380 ( .A(n5382), .B(n5383), .Z(n5374) );
  AND U5381 ( .A(n234), .B(n5373), .Z(n5383) );
  XNOR U5382 ( .A(n5384), .B(n5371), .Z(n5373) );
  XOR U5383 ( .A(n5385), .B(n5386), .Z(n5371) );
  AND U5384 ( .A(n257), .B(n5387), .Z(n5386) );
  IV U5385 ( .A(n5382), .Z(n5384) );
  XOR U5386 ( .A(n5388), .B(n5389), .Z(n5382) );
  AND U5387 ( .A(n241), .B(n5381), .Z(n5389) );
  XNOR U5388 ( .A(n5379), .B(n5388), .Z(n5381) );
  XNOR U5389 ( .A(n5390), .B(n5391), .Z(n5379) );
  AND U5390 ( .A(n245), .B(n5392), .Z(n5391) );
  XOR U5391 ( .A(p_input[205]), .B(n5390), .Z(n5392) );
  XNOR U5392 ( .A(n5393), .B(n5394), .Z(n5390) );
  AND U5393 ( .A(n249), .B(n5395), .Z(n5394) );
  XOR U5394 ( .A(n5396), .B(n5397), .Z(n5388) );
  AND U5395 ( .A(n253), .B(n5387), .Z(n5397) );
  XNOR U5396 ( .A(n5398), .B(n5385), .Z(n5387) );
  XOR U5397 ( .A(n5399), .B(n5400), .Z(n5385) );
  AND U5398 ( .A(n276), .B(n5401), .Z(n5400) );
  IV U5399 ( .A(n5396), .Z(n5398) );
  XOR U5400 ( .A(n5402), .B(n5403), .Z(n5396) );
  AND U5401 ( .A(n260), .B(n5395), .Z(n5403) );
  XNOR U5402 ( .A(n5393), .B(n5402), .Z(n5395) );
  XNOR U5403 ( .A(n5404), .B(n5405), .Z(n5393) );
  AND U5404 ( .A(n264), .B(n5406), .Z(n5405) );
  XOR U5405 ( .A(p_input[237]), .B(n5404), .Z(n5406) );
  XNOR U5406 ( .A(n5407), .B(n5408), .Z(n5404) );
  AND U5407 ( .A(n268), .B(n5409), .Z(n5408) );
  XOR U5408 ( .A(n5410), .B(n5411), .Z(n5402) );
  AND U5409 ( .A(n272), .B(n5401), .Z(n5411) );
  XNOR U5410 ( .A(n5412), .B(n5399), .Z(n5401) );
  XOR U5411 ( .A(n5413), .B(n5414), .Z(n5399) );
  AND U5412 ( .A(n295), .B(n5415), .Z(n5414) );
  IV U5413 ( .A(n5410), .Z(n5412) );
  XOR U5414 ( .A(n5416), .B(n5417), .Z(n5410) );
  AND U5415 ( .A(n279), .B(n5409), .Z(n5417) );
  XNOR U5416 ( .A(n5407), .B(n5416), .Z(n5409) );
  XNOR U5417 ( .A(n5418), .B(n5419), .Z(n5407) );
  AND U5418 ( .A(n283), .B(n5420), .Z(n5419) );
  XOR U5419 ( .A(p_input[269]), .B(n5418), .Z(n5420) );
  XNOR U5420 ( .A(n5421), .B(n5422), .Z(n5418) );
  AND U5421 ( .A(n287), .B(n5423), .Z(n5422) );
  XOR U5422 ( .A(n5424), .B(n5425), .Z(n5416) );
  AND U5423 ( .A(n291), .B(n5415), .Z(n5425) );
  XNOR U5424 ( .A(n5426), .B(n5413), .Z(n5415) );
  XOR U5425 ( .A(n5427), .B(n5428), .Z(n5413) );
  AND U5426 ( .A(n314), .B(n5429), .Z(n5428) );
  IV U5427 ( .A(n5424), .Z(n5426) );
  XOR U5428 ( .A(n5430), .B(n5431), .Z(n5424) );
  AND U5429 ( .A(n298), .B(n5423), .Z(n5431) );
  XNOR U5430 ( .A(n5421), .B(n5430), .Z(n5423) );
  XNOR U5431 ( .A(n5432), .B(n5433), .Z(n5421) );
  AND U5432 ( .A(n302), .B(n5434), .Z(n5433) );
  XOR U5433 ( .A(p_input[301]), .B(n5432), .Z(n5434) );
  XNOR U5434 ( .A(n5435), .B(n5436), .Z(n5432) );
  AND U5435 ( .A(n306), .B(n5437), .Z(n5436) );
  XOR U5436 ( .A(n5438), .B(n5439), .Z(n5430) );
  AND U5437 ( .A(n310), .B(n5429), .Z(n5439) );
  XNOR U5438 ( .A(n5440), .B(n5427), .Z(n5429) );
  XOR U5439 ( .A(n5441), .B(n5442), .Z(n5427) );
  AND U5440 ( .A(n333), .B(n5443), .Z(n5442) );
  IV U5441 ( .A(n5438), .Z(n5440) );
  XOR U5442 ( .A(n5444), .B(n5445), .Z(n5438) );
  AND U5443 ( .A(n317), .B(n5437), .Z(n5445) );
  XNOR U5444 ( .A(n5435), .B(n5444), .Z(n5437) );
  XNOR U5445 ( .A(n5446), .B(n5447), .Z(n5435) );
  AND U5446 ( .A(n321), .B(n5448), .Z(n5447) );
  XOR U5447 ( .A(p_input[333]), .B(n5446), .Z(n5448) );
  XNOR U5448 ( .A(n5449), .B(n5450), .Z(n5446) );
  AND U5449 ( .A(n325), .B(n5451), .Z(n5450) );
  XOR U5450 ( .A(n5452), .B(n5453), .Z(n5444) );
  AND U5451 ( .A(n329), .B(n5443), .Z(n5453) );
  XNOR U5452 ( .A(n5454), .B(n5441), .Z(n5443) );
  XOR U5453 ( .A(n5455), .B(n5456), .Z(n5441) );
  AND U5454 ( .A(n352), .B(n5457), .Z(n5456) );
  IV U5455 ( .A(n5452), .Z(n5454) );
  XOR U5456 ( .A(n5458), .B(n5459), .Z(n5452) );
  AND U5457 ( .A(n336), .B(n5451), .Z(n5459) );
  XNOR U5458 ( .A(n5449), .B(n5458), .Z(n5451) );
  XNOR U5459 ( .A(n5460), .B(n5461), .Z(n5449) );
  AND U5460 ( .A(n340), .B(n5462), .Z(n5461) );
  XOR U5461 ( .A(p_input[365]), .B(n5460), .Z(n5462) );
  XNOR U5462 ( .A(n5463), .B(n5464), .Z(n5460) );
  AND U5463 ( .A(n344), .B(n5465), .Z(n5464) );
  XOR U5464 ( .A(n5466), .B(n5467), .Z(n5458) );
  AND U5465 ( .A(n348), .B(n5457), .Z(n5467) );
  XNOR U5466 ( .A(n5468), .B(n5455), .Z(n5457) );
  XOR U5467 ( .A(n5469), .B(n5470), .Z(n5455) );
  AND U5468 ( .A(n370), .B(n5471), .Z(n5470) );
  IV U5469 ( .A(n5466), .Z(n5468) );
  XOR U5470 ( .A(n5472), .B(n5473), .Z(n5466) );
  AND U5471 ( .A(n355), .B(n5465), .Z(n5473) );
  XNOR U5472 ( .A(n5463), .B(n5472), .Z(n5465) );
  XNOR U5473 ( .A(n5474), .B(n5475), .Z(n5463) );
  AND U5474 ( .A(n359), .B(n5476), .Z(n5475) );
  XOR U5475 ( .A(p_input[397]), .B(n5474), .Z(n5476) );
  XOR U5476 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(n5477), 
        .Z(n5474) );
  AND U5477 ( .A(n362), .B(n5478), .Z(n5477) );
  XOR U5478 ( .A(n5479), .B(n5480), .Z(n5472) );
  AND U5479 ( .A(n366), .B(n5471), .Z(n5480) );
  XNOR U5480 ( .A(n5481), .B(n5469), .Z(n5471) );
  XOR U5481 ( .A(\knn_comb_/min_val_out[0][13] ), .B(n5482), .Z(n5469) );
  AND U5482 ( .A(n378), .B(n5483), .Z(n5482) );
  IV U5483 ( .A(n5479), .Z(n5481) );
  XOR U5484 ( .A(n5484), .B(n5485), .Z(n5479) );
  AND U5485 ( .A(n373), .B(n5478), .Z(n5485) );
  XOR U5486 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(n5484), 
        .Z(n5478) );
  XOR U5487 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(n5486), 
        .Z(n5484) );
  AND U5488 ( .A(n375), .B(n5483), .Z(n5486) );
  XOR U5489 ( .A(\knn_comb_/min_val_out[0][13] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .Z(n5483) );
  XOR U5490 ( .A(n115), .B(n5487), .Z(o[12]) );
  AND U5491 ( .A(n122), .B(n5488), .Z(n115) );
  XOR U5492 ( .A(n116), .B(n5487), .Z(n5488) );
  XOR U5493 ( .A(n5489), .B(n5490), .Z(n5487) );
  AND U5494 ( .A(n142), .B(n5491), .Z(n5490) );
  XOR U5495 ( .A(n5492), .B(n45), .Z(n116) );
  AND U5496 ( .A(n125), .B(n5493), .Z(n45) );
  XOR U5497 ( .A(n46), .B(n5492), .Z(n5493) );
  XOR U5498 ( .A(n5494), .B(n5495), .Z(n46) );
  AND U5499 ( .A(n130), .B(n5496), .Z(n5495) );
  XOR U5500 ( .A(p_input[12]), .B(n5494), .Z(n5496) );
  XNOR U5501 ( .A(n5497), .B(n5498), .Z(n5494) );
  AND U5502 ( .A(n134), .B(n5499), .Z(n5498) );
  XOR U5503 ( .A(n5500), .B(n5501), .Z(n5492) );
  AND U5504 ( .A(n138), .B(n5491), .Z(n5501) );
  XNOR U5505 ( .A(n5502), .B(n5489), .Z(n5491) );
  XOR U5506 ( .A(n5503), .B(n5504), .Z(n5489) );
  AND U5507 ( .A(n162), .B(n5505), .Z(n5504) );
  IV U5508 ( .A(n5500), .Z(n5502) );
  XOR U5509 ( .A(n5506), .B(n5507), .Z(n5500) );
  AND U5510 ( .A(n146), .B(n5499), .Z(n5507) );
  XNOR U5511 ( .A(n5497), .B(n5506), .Z(n5499) );
  XNOR U5512 ( .A(n5508), .B(n5509), .Z(n5497) );
  AND U5513 ( .A(n150), .B(n5510), .Z(n5509) );
  XOR U5514 ( .A(p_input[44]), .B(n5508), .Z(n5510) );
  XNOR U5515 ( .A(n5511), .B(n5512), .Z(n5508) );
  AND U5516 ( .A(n154), .B(n5513), .Z(n5512) );
  XOR U5517 ( .A(n5514), .B(n5515), .Z(n5506) );
  AND U5518 ( .A(n158), .B(n5505), .Z(n5515) );
  XNOR U5519 ( .A(n5516), .B(n5503), .Z(n5505) );
  XOR U5520 ( .A(n5517), .B(n5518), .Z(n5503) );
  AND U5521 ( .A(n181), .B(n5519), .Z(n5518) );
  IV U5522 ( .A(n5514), .Z(n5516) );
  XOR U5523 ( .A(n5520), .B(n5521), .Z(n5514) );
  AND U5524 ( .A(n165), .B(n5513), .Z(n5521) );
  XNOR U5525 ( .A(n5511), .B(n5520), .Z(n5513) );
  XNOR U5526 ( .A(n5522), .B(n5523), .Z(n5511) );
  AND U5527 ( .A(n169), .B(n5524), .Z(n5523) );
  XOR U5528 ( .A(p_input[76]), .B(n5522), .Z(n5524) );
  XNOR U5529 ( .A(n5525), .B(n5526), .Z(n5522) );
  AND U5530 ( .A(n173), .B(n5527), .Z(n5526) );
  XOR U5531 ( .A(n5528), .B(n5529), .Z(n5520) );
  AND U5532 ( .A(n177), .B(n5519), .Z(n5529) );
  XNOR U5533 ( .A(n5530), .B(n5517), .Z(n5519) );
  XOR U5534 ( .A(n5531), .B(n5532), .Z(n5517) );
  AND U5535 ( .A(n200), .B(n5533), .Z(n5532) );
  IV U5536 ( .A(n5528), .Z(n5530) );
  XOR U5537 ( .A(n5534), .B(n5535), .Z(n5528) );
  AND U5538 ( .A(n184), .B(n5527), .Z(n5535) );
  XNOR U5539 ( .A(n5525), .B(n5534), .Z(n5527) );
  XNOR U5540 ( .A(n5536), .B(n5537), .Z(n5525) );
  AND U5541 ( .A(n188), .B(n5538), .Z(n5537) );
  XOR U5542 ( .A(p_input[108]), .B(n5536), .Z(n5538) );
  XNOR U5543 ( .A(n5539), .B(n5540), .Z(n5536) );
  AND U5544 ( .A(n192), .B(n5541), .Z(n5540) );
  XOR U5545 ( .A(n5542), .B(n5543), .Z(n5534) );
  AND U5546 ( .A(n196), .B(n5533), .Z(n5543) );
  XNOR U5547 ( .A(n5544), .B(n5531), .Z(n5533) );
  XOR U5548 ( .A(n5545), .B(n5546), .Z(n5531) );
  AND U5549 ( .A(n219), .B(n5547), .Z(n5546) );
  IV U5550 ( .A(n5542), .Z(n5544) );
  XOR U5551 ( .A(n5548), .B(n5549), .Z(n5542) );
  AND U5552 ( .A(n203), .B(n5541), .Z(n5549) );
  XNOR U5553 ( .A(n5539), .B(n5548), .Z(n5541) );
  XNOR U5554 ( .A(n5550), .B(n5551), .Z(n5539) );
  AND U5555 ( .A(n207), .B(n5552), .Z(n5551) );
  XOR U5556 ( .A(p_input[140]), .B(n5550), .Z(n5552) );
  XNOR U5557 ( .A(n5553), .B(n5554), .Z(n5550) );
  AND U5558 ( .A(n211), .B(n5555), .Z(n5554) );
  XOR U5559 ( .A(n5556), .B(n5557), .Z(n5548) );
  AND U5560 ( .A(n215), .B(n5547), .Z(n5557) );
  XNOR U5561 ( .A(n5558), .B(n5545), .Z(n5547) );
  XOR U5562 ( .A(n5559), .B(n5560), .Z(n5545) );
  AND U5563 ( .A(n238), .B(n5561), .Z(n5560) );
  IV U5564 ( .A(n5556), .Z(n5558) );
  XOR U5565 ( .A(n5562), .B(n5563), .Z(n5556) );
  AND U5566 ( .A(n222), .B(n5555), .Z(n5563) );
  XNOR U5567 ( .A(n5553), .B(n5562), .Z(n5555) );
  XNOR U5568 ( .A(n5564), .B(n5565), .Z(n5553) );
  AND U5569 ( .A(n226), .B(n5566), .Z(n5565) );
  XOR U5570 ( .A(p_input[172]), .B(n5564), .Z(n5566) );
  XNOR U5571 ( .A(n5567), .B(n5568), .Z(n5564) );
  AND U5572 ( .A(n230), .B(n5569), .Z(n5568) );
  XOR U5573 ( .A(n5570), .B(n5571), .Z(n5562) );
  AND U5574 ( .A(n234), .B(n5561), .Z(n5571) );
  XNOR U5575 ( .A(n5572), .B(n5559), .Z(n5561) );
  XOR U5576 ( .A(n5573), .B(n5574), .Z(n5559) );
  AND U5577 ( .A(n257), .B(n5575), .Z(n5574) );
  IV U5578 ( .A(n5570), .Z(n5572) );
  XOR U5579 ( .A(n5576), .B(n5577), .Z(n5570) );
  AND U5580 ( .A(n241), .B(n5569), .Z(n5577) );
  XNOR U5581 ( .A(n5567), .B(n5576), .Z(n5569) );
  XNOR U5582 ( .A(n5578), .B(n5579), .Z(n5567) );
  AND U5583 ( .A(n245), .B(n5580), .Z(n5579) );
  XOR U5584 ( .A(p_input[204]), .B(n5578), .Z(n5580) );
  XNOR U5585 ( .A(n5581), .B(n5582), .Z(n5578) );
  AND U5586 ( .A(n249), .B(n5583), .Z(n5582) );
  XOR U5587 ( .A(n5584), .B(n5585), .Z(n5576) );
  AND U5588 ( .A(n253), .B(n5575), .Z(n5585) );
  XNOR U5589 ( .A(n5586), .B(n5573), .Z(n5575) );
  XOR U5590 ( .A(n5587), .B(n5588), .Z(n5573) );
  AND U5591 ( .A(n276), .B(n5589), .Z(n5588) );
  IV U5592 ( .A(n5584), .Z(n5586) );
  XOR U5593 ( .A(n5590), .B(n5591), .Z(n5584) );
  AND U5594 ( .A(n260), .B(n5583), .Z(n5591) );
  XNOR U5595 ( .A(n5581), .B(n5590), .Z(n5583) );
  XNOR U5596 ( .A(n5592), .B(n5593), .Z(n5581) );
  AND U5597 ( .A(n264), .B(n5594), .Z(n5593) );
  XOR U5598 ( .A(p_input[236]), .B(n5592), .Z(n5594) );
  XNOR U5599 ( .A(n5595), .B(n5596), .Z(n5592) );
  AND U5600 ( .A(n268), .B(n5597), .Z(n5596) );
  XOR U5601 ( .A(n5598), .B(n5599), .Z(n5590) );
  AND U5602 ( .A(n272), .B(n5589), .Z(n5599) );
  XNOR U5603 ( .A(n5600), .B(n5587), .Z(n5589) );
  XOR U5604 ( .A(n5601), .B(n5602), .Z(n5587) );
  AND U5605 ( .A(n295), .B(n5603), .Z(n5602) );
  IV U5606 ( .A(n5598), .Z(n5600) );
  XOR U5607 ( .A(n5604), .B(n5605), .Z(n5598) );
  AND U5608 ( .A(n279), .B(n5597), .Z(n5605) );
  XNOR U5609 ( .A(n5595), .B(n5604), .Z(n5597) );
  XNOR U5610 ( .A(n5606), .B(n5607), .Z(n5595) );
  AND U5611 ( .A(n283), .B(n5608), .Z(n5607) );
  XOR U5612 ( .A(p_input[268]), .B(n5606), .Z(n5608) );
  XNOR U5613 ( .A(n5609), .B(n5610), .Z(n5606) );
  AND U5614 ( .A(n287), .B(n5611), .Z(n5610) );
  XOR U5615 ( .A(n5612), .B(n5613), .Z(n5604) );
  AND U5616 ( .A(n291), .B(n5603), .Z(n5613) );
  XNOR U5617 ( .A(n5614), .B(n5601), .Z(n5603) );
  XOR U5618 ( .A(n5615), .B(n5616), .Z(n5601) );
  AND U5619 ( .A(n314), .B(n5617), .Z(n5616) );
  IV U5620 ( .A(n5612), .Z(n5614) );
  XOR U5621 ( .A(n5618), .B(n5619), .Z(n5612) );
  AND U5622 ( .A(n298), .B(n5611), .Z(n5619) );
  XNOR U5623 ( .A(n5609), .B(n5618), .Z(n5611) );
  XNOR U5624 ( .A(n5620), .B(n5621), .Z(n5609) );
  AND U5625 ( .A(n302), .B(n5622), .Z(n5621) );
  XOR U5626 ( .A(p_input[300]), .B(n5620), .Z(n5622) );
  XNOR U5627 ( .A(n5623), .B(n5624), .Z(n5620) );
  AND U5628 ( .A(n306), .B(n5625), .Z(n5624) );
  XOR U5629 ( .A(n5626), .B(n5627), .Z(n5618) );
  AND U5630 ( .A(n310), .B(n5617), .Z(n5627) );
  XNOR U5631 ( .A(n5628), .B(n5615), .Z(n5617) );
  XOR U5632 ( .A(n5629), .B(n5630), .Z(n5615) );
  AND U5633 ( .A(n333), .B(n5631), .Z(n5630) );
  IV U5634 ( .A(n5626), .Z(n5628) );
  XOR U5635 ( .A(n5632), .B(n5633), .Z(n5626) );
  AND U5636 ( .A(n317), .B(n5625), .Z(n5633) );
  XNOR U5637 ( .A(n5623), .B(n5632), .Z(n5625) );
  XNOR U5638 ( .A(n5634), .B(n5635), .Z(n5623) );
  AND U5639 ( .A(n321), .B(n5636), .Z(n5635) );
  XOR U5640 ( .A(p_input[332]), .B(n5634), .Z(n5636) );
  XNOR U5641 ( .A(n5637), .B(n5638), .Z(n5634) );
  AND U5642 ( .A(n325), .B(n5639), .Z(n5638) );
  XOR U5643 ( .A(n5640), .B(n5641), .Z(n5632) );
  AND U5644 ( .A(n329), .B(n5631), .Z(n5641) );
  XNOR U5645 ( .A(n5642), .B(n5629), .Z(n5631) );
  XOR U5646 ( .A(n5643), .B(n5644), .Z(n5629) );
  AND U5647 ( .A(n352), .B(n5645), .Z(n5644) );
  IV U5648 ( .A(n5640), .Z(n5642) );
  XOR U5649 ( .A(n5646), .B(n5647), .Z(n5640) );
  AND U5650 ( .A(n336), .B(n5639), .Z(n5647) );
  XNOR U5651 ( .A(n5637), .B(n5646), .Z(n5639) );
  XNOR U5652 ( .A(n5648), .B(n5649), .Z(n5637) );
  AND U5653 ( .A(n340), .B(n5650), .Z(n5649) );
  XOR U5654 ( .A(p_input[364]), .B(n5648), .Z(n5650) );
  XNOR U5655 ( .A(n5651), .B(n5652), .Z(n5648) );
  AND U5656 ( .A(n344), .B(n5653), .Z(n5652) );
  XOR U5657 ( .A(n5654), .B(n5655), .Z(n5646) );
  AND U5658 ( .A(n348), .B(n5645), .Z(n5655) );
  XNOR U5659 ( .A(n5656), .B(n5643), .Z(n5645) );
  XOR U5660 ( .A(n5657), .B(n5658), .Z(n5643) );
  AND U5661 ( .A(n370), .B(n5659), .Z(n5658) );
  IV U5662 ( .A(n5654), .Z(n5656) );
  XOR U5663 ( .A(n5660), .B(n5661), .Z(n5654) );
  AND U5664 ( .A(n355), .B(n5653), .Z(n5661) );
  XNOR U5665 ( .A(n5651), .B(n5660), .Z(n5653) );
  XNOR U5666 ( .A(n5662), .B(n5663), .Z(n5651) );
  AND U5667 ( .A(n359), .B(n5664), .Z(n5663) );
  XOR U5668 ( .A(p_input[396]), .B(n5662), .Z(n5664) );
  XOR U5669 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n5665), 
        .Z(n5662) );
  AND U5670 ( .A(n362), .B(n5666), .Z(n5665) );
  XOR U5671 ( .A(n5667), .B(n5668), .Z(n5660) );
  AND U5672 ( .A(n366), .B(n5659), .Z(n5668) );
  XNOR U5673 ( .A(n5669), .B(n5657), .Z(n5659) );
  XOR U5674 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n5670), .Z(n5657) );
  AND U5675 ( .A(n378), .B(n5671), .Z(n5670) );
  IV U5676 ( .A(n5667), .Z(n5669) );
  XOR U5677 ( .A(n5672), .B(n5673), .Z(n5667) );
  AND U5678 ( .A(n373), .B(n5666), .Z(n5673) );
  XOR U5679 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n5672), 
        .Z(n5666) );
  XOR U5680 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(n5674), 
        .Z(n5672) );
  AND U5681 ( .A(n375), .B(n5671), .Z(n5674) );
  XOR U5682 ( .A(n5675), .B(n5676), .Z(n5671) );
  IV U5683 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .Z(n5676) );
  IV U5684 ( .A(\knn_comb_/min_val_out[0][12] ), .Z(n5675) );
  XOR U5685 ( .A(n117), .B(n5677), .Z(o[11]) );
  AND U5686 ( .A(n122), .B(n5678), .Z(n117) );
  XOR U5687 ( .A(n118), .B(n5677), .Z(n5678) );
  XOR U5688 ( .A(n5679), .B(n5680), .Z(n5677) );
  AND U5689 ( .A(n142), .B(n5681), .Z(n5680) );
  XOR U5690 ( .A(n5682), .B(n47), .Z(n118) );
  AND U5691 ( .A(n125), .B(n5683), .Z(n47) );
  XOR U5692 ( .A(n48), .B(n5682), .Z(n5683) );
  XOR U5693 ( .A(n5684), .B(n5685), .Z(n48) );
  AND U5694 ( .A(n130), .B(n5686), .Z(n5685) );
  XOR U5695 ( .A(p_input[11]), .B(n5684), .Z(n5686) );
  XNOR U5696 ( .A(n5687), .B(n5688), .Z(n5684) );
  AND U5697 ( .A(n134), .B(n5689), .Z(n5688) );
  XOR U5698 ( .A(n5690), .B(n5691), .Z(n5682) );
  AND U5699 ( .A(n138), .B(n5681), .Z(n5691) );
  XNOR U5700 ( .A(n5692), .B(n5679), .Z(n5681) );
  XOR U5701 ( .A(n5693), .B(n5694), .Z(n5679) );
  AND U5702 ( .A(n162), .B(n5695), .Z(n5694) );
  IV U5703 ( .A(n5690), .Z(n5692) );
  XOR U5704 ( .A(n5696), .B(n5697), .Z(n5690) );
  AND U5705 ( .A(n146), .B(n5689), .Z(n5697) );
  XNOR U5706 ( .A(n5687), .B(n5696), .Z(n5689) );
  XNOR U5707 ( .A(n5698), .B(n5699), .Z(n5687) );
  AND U5708 ( .A(n150), .B(n5700), .Z(n5699) );
  XOR U5709 ( .A(p_input[43]), .B(n5698), .Z(n5700) );
  XNOR U5710 ( .A(n5701), .B(n5702), .Z(n5698) );
  AND U5711 ( .A(n154), .B(n5703), .Z(n5702) );
  XOR U5712 ( .A(n5704), .B(n5705), .Z(n5696) );
  AND U5713 ( .A(n158), .B(n5695), .Z(n5705) );
  XNOR U5714 ( .A(n5706), .B(n5693), .Z(n5695) );
  XOR U5715 ( .A(n5707), .B(n5708), .Z(n5693) );
  AND U5716 ( .A(n181), .B(n5709), .Z(n5708) );
  IV U5717 ( .A(n5704), .Z(n5706) );
  XOR U5718 ( .A(n5710), .B(n5711), .Z(n5704) );
  AND U5719 ( .A(n165), .B(n5703), .Z(n5711) );
  XNOR U5720 ( .A(n5701), .B(n5710), .Z(n5703) );
  XNOR U5721 ( .A(n5712), .B(n5713), .Z(n5701) );
  AND U5722 ( .A(n169), .B(n5714), .Z(n5713) );
  XOR U5723 ( .A(p_input[75]), .B(n5712), .Z(n5714) );
  XNOR U5724 ( .A(n5715), .B(n5716), .Z(n5712) );
  AND U5725 ( .A(n173), .B(n5717), .Z(n5716) );
  XOR U5726 ( .A(n5718), .B(n5719), .Z(n5710) );
  AND U5727 ( .A(n177), .B(n5709), .Z(n5719) );
  XNOR U5728 ( .A(n5720), .B(n5707), .Z(n5709) );
  XOR U5729 ( .A(n5721), .B(n5722), .Z(n5707) );
  AND U5730 ( .A(n200), .B(n5723), .Z(n5722) );
  IV U5731 ( .A(n5718), .Z(n5720) );
  XOR U5732 ( .A(n5724), .B(n5725), .Z(n5718) );
  AND U5733 ( .A(n184), .B(n5717), .Z(n5725) );
  XNOR U5734 ( .A(n5715), .B(n5724), .Z(n5717) );
  XNOR U5735 ( .A(n5726), .B(n5727), .Z(n5715) );
  AND U5736 ( .A(n188), .B(n5728), .Z(n5727) );
  XOR U5737 ( .A(p_input[107]), .B(n5726), .Z(n5728) );
  XNOR U5738 ( .A(n5729), .B(n5730), .Z(n5726) );
  AND U5739 ( .A(n192), .B(n5731), .Z(n5730) );
  XOR U5740 ( .A(n5732), .B(n5733), .Z(n5724) );
  AND U5741 ( .A(n196), .B(n5723), .Z(n5733) );
  XNOR U5742 ( .A(n5734), .B(n5721), .Z(n5723) );
  XOR U5743 ( .A(n5735), .B(n5736), .Z(n5721) );
  AND U5744 ( .A(n219), .B(n5737), .Z(n5736) );
  IV U5745 ( .A(n5732), .Z(n5734) );
  XOR U5746 ( .A(n5738), .B(n5739), .Z(n5732) );
  AND U5747 ( .A(n203), .B(n5731), .Z(n5739) );
  XNOR U5748 ( .A(n5729), .B(n5738), .Z(n5731) );
  XNOR U5749 ( .A(n5740), .B(n5741), .Z(n5729) );
  AND U5750 ( .A(n207), .B(n5742), .Z(n5741) );
  XOR U5751 ( .A(p_input[139]), .B(n5740), .Z(n5742) );
  XNOR U5752 ( .A(n5743), .B(n5744), .Z(n5740) );
  AND U5753 ( .A(n211), .B(n5745), .Z(n5744) );
  XOR U5754 ( .A(n5746), .B(n5747), .Z(n5738) );
  AND U5755 ( .A(n215), .B(n5737), .Z(n5747) );
  XNOR U5756 ( .A(n5748), .B(n5735), .Z(n5737) );
  XOR U5757 ( .A(n5749), .B(n5750), .Z(n5735) );
  AND U5758 ( .A(n238), .B(n5751), .Z(n5750) );
  IV U5759 ( .A(n5746), .Z(n5748) );
  XOR U5760 ( .A(n5752), .B(n5753), .Z(n5746) );
  AND U5761 ( .A(n222), .B(n5745), .Z(n5753) );
  XNOR U5762 ( .A(n5743), .B(n5752), .Z(n5745) );
  XNOR U5763 ( .A(n5754), .B(n5755), .Z(n5743) );
  AND U5764 ( .A(n226), .B(n5756), .Z(n5755) );
  XOR U5765 ( .A(p_input[171]), .B(n5754), .Z(n5756) );
  XNOR U5766 ( .A(n5757), .B(n5758), .Z(n5754) );
  AND U5767 ( .A(n230), .B(n5759), .Z(n5758) );
  XOR U5768 ( .A(n5760), .B(n5761), .Z(n5752) );
  AND U5769 ( .A(n234), .B(n5751), .Z(n5761) );
  XNOR U5770 ( .A(n5762), .B(n5749), .Z(n5751) );
  XOR U5771 ( .A(n5763), .B(n5764), .Z(n5749) );
  AND U5772 ( .A(n257), .B(n5765), .Z(n5764) );
  IV U5773 ( .A(n5760), .Z(n5762) );
  XOR U5774 ( .A(n5766), .B(n5767), .Z(n5760) );
  AND U5775 ( .A(n241), .B(n5759), .Z(n5767) );
  XNOR U5776 ( .A(n5757), .B(n5766), .Z(n5759) );
  XNOR U5777 ( .A(n5768), .B(n5769), .Z(n5757) );
  AND U5778 ( .A(n245), .B(n5770), .Z(n5769) );
  XOR U5779 ( .A(p_input[203]), .B(n5768), .Z(n5770) );
  XNOR U5780 ( .A(n5771), .B(n5772), .Z(n5768) );
  AND U5781 ( .A(n249), .B(n5773), .Z(n5772) );
  XOR U5782 ( .A(n5774), .B(n5775), .Z(n5766) );
  AND U5783 ( .A(n253), .B(n5765), .Z(n5775) );
  XNOR U5784 ( .A(n5776), .B(n5763), .Z(n5765) );
  XOR U5785 ( .A(n5777), .B(n5778), .Z(n5763) );
  AND U5786 ( .A(n276), .B(n5779), .Z(n5778) );
  IV U5787 ( .A(n5774), .Z(n5776) );
  XOR U5788 ( .A(n5780), .B(n5781), .Z(n5774) );
  AND U5789 ( .A(n260), .B(n5773), .Z(n5781) );
  XNOR U5790 ( .A(n5771), .B(n5780), .Z(n5773) );
  XNOR U5791 ( .A(n5782), .B(n5783), .Z(n5771) );
  AND U5792 ( .A(n264), .B(n5784), .Z(n5783) );
  XOR U5793 ( .A(p_input[235]), .B(n5782), .Z(n5784) );
  XNOR U5794 ( .A(n5785), .B(n5786), .Z(n5782) );
  AND U5795 ( .A(n268), .B(n5787), .Z(n5786) );
  XOR U5796 ( .A(n5788), .B(n5789), .Z(n5780) );
  AND U5797 ( .A(n272), .B(n5779), .Z(n5789) );
  XNOR U5798 ( .A(n5790), .B(n5777), .Z(n5779) );
  XOR U5799 ( .A(n5791), .B(n5792), .Z(n5777) );
  AND U5800 ( .A(n295), .B(n5793), .Z(n5792) );
  IV U5801 ( .A(n5788), .Z(n5790) );
  XOR U5802 ( .A(n5794), .B(n5795), .Z(n5788) );
  AND U5803 ( .A(n279), .B(n5787), .Z(n5795) );
  XNOR U5804 ( .A(n5785), .B(n5794), .Z(n5787) );
  XNOR U5805 ( .A(n5796), .B(n5797), .Z(n5785) );
  AND U5806 ( .A(n283), .B(n5798), .Z(n5797) );
  XOR U5807 ( .A(p_input[267]), .B(n5796), .Z(n5798) );
  XNOR U5808 ( .A(n5799), .B(n5800), .Z(n5796) );
  AND U5809 ( .A(n287), .B(n5801), .Z(n5800) );
  XOR U5810 ( .A(n5802), .B(n5803), .Z(n5794) );
  AND U5811 ( .A(n291), .B(n5793), .Z(n5803) );
  XNOR U5812 ( .A(n5804), .B(n5791), .Z(n5793) );
  XOR U5813 ( .A(n5805), .B(n5806), .Z(n5791) );
  AND U5814 ( .A(n314), .B(n5807), .Z(n5806) );
  IV U5815 ( .A(n5802), .Z(n5804) );
  XOR U5816 ( .A(n5808), .B(n5809), .Z(n5802) );
  AND U5817 ( .A(n298), .B(n5801), .Z(n5809) );
  XNOR U5818 ( .A(n5799), .B(n5808), .Z(n5801) );
  XNOR U5819 ( .A(n5810), .B(n5811), .Z(n5799) );
  AND U5820 ( .A(n302), .B(n5812), .Z(n5811) );
  XOR U5821 ( .A(p_input[299]), .B(n5810), .Z(n5812) );
  XNOR U5822 ( .A(n5813), .B(n5814), .Z(n5810) );
  AND U5823 ( .A(n306), .B(n5815), .Z(n5814) );
  XOR U5824 ( .A(n5816), .B(n5817), .Z(n5808) );
  AND U5825 ( .A(n310), .B(n5807), .Z(n5817) );
  XNOR U5826 ( .A(n5818), .B(n5805), .Z(n5807) );
  XOR U5827 ( .A(n5819), .B(n5820), .Z(n5805) );
  AND U5828 ( .A(n333), .B(n5821), .Z(n5820) );
  IV U5829 ( .A(n5816), .Z(n5818) );
  XOR U5830 ( .A(n5822), .B(n5823), .Z(n5816) );
  AND U5831 ( .A(n317), .B(n5815), .Z(n5823) );
  XNOR U5832 ( .A(n5813), .B(n5822), .Z(n5815) );
  XNOR U5833 ( .A(n5824), .B(n5825), .Z(n5813) );
  AND U5834 ( .A(n321), .B(n5826), .Z(n5825) );
  XOR U5835 ( .A(p_input[331]), .B(n5824), .Z(n5826) );
  XNOR U5836 ( .A(n5827), .B(n5828), .Z(n5824) );
  AND U5837 ( .A(n325), .B(n5829), .Z(n5828) );
  XOR U5838 ( .A(n5830), .B(n5831), .Z(n5822) );
  AND U5839 ( .A(n329), .B(n5821), .Z(n5831) );
  XNOR U5840 ( .A(n5832), .B(n5819), .Z(n5821) );
  XOR U5841 ( .A(n5833), .B(n5834), .Z(n5819) );
  AND U5842 ( .A(n352), .B(n5835), .Z(n5834) );
  IV U5843 ( .A(n5830), .Z(n5832) );
  XOR U5844 ( .A(n5836), .B(n5837), .Z(n5830) );
  AND U5845 ( .A(n336), .B(n5829), .Z(n5837) );
  XNOR U5846 ( .A(n5827), .B(n5836), .Z(n5829) );
  XNOR U5847 ( .A(n5838), .B(n5839), .Z(n5827) );
  AND U5848 ( .A(n340), .B(n5840), .Z(n5839) );
  XOR U5849 ( .A(p_input[363]), .B(n5838), .Z(n5840) );
  XNOR U5850 ( .A(n5841), .B(n5842), .Z(n5838) );
  AND U5851 ( .A(n344), .B(n5843), .Z(n5842) );
  XOR U5852 ( .A(n5844), .B(n5845), .Z(n5836) );
  AND U5853 ( .A(n348), .B(n5835), .Z(n5845) );
  XNOR U5854 ( .A(n5846), .B(n5833), .Z(n5835) );
  XOR U5855 ( .A(n5847), .B(n5848), .Z(n5833) );
  AND U5856 ( .A(n370), .B(n5849), .Z(n5848) );
  IV U5857 ( .A(n5844), .Z(n5846) );
  XOR U5858 ( .A(n5850), .B(n5851), .Z(n5844) );
  AND U5859 ( .A(n355), .B(n5843), .Z(n5851) );
  XNOR U5860 ( .A(n5841), .B(n5850), .Z(n5843) );
  XNOR U5861 ( .A(n5852), .B(n5853), .Z(n5841) );
  AND U5862 ( .A(n359), .B(n5854), .Z(n5853) );
  XOR U5863 ( .A(p_input[395]), .B(n5852), .Z(n5854) );
  XOR U5864 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n5855), 
        .Z(n5852) );
  AND U5865 ( .A(n362), .B(n5856), .Z(n5855) );
  XOR U5866 ( .A(n5857), .B(n5858), .Z(n5850) );
  AND U5867 ( .A(n366), .B(n5849), .Z(n5858) );
  XNOR U5868 ( .A(n5859), .B(n5847), .Z(n5849) );
  XOR U5869 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n5860), .Z(n5847) );
  AND U5870 ( .A(n378), .B(n5861), .Z(n5860) );
  IV U5871 ( .A(n5857), .Z(n5859) );
  XOR U5872 ( .A(n5862), .B(n5863), .Z(n5857) );
  AND U5873 ( .A(n373), .B(n5856), .Z(n5863) );
  XOR U5874 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n5862), 
        .Z(n5856) );
  XOR U5875 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n5864), 
        .Z(n5862) );
  AND U5876 ( .A(n375), .B(n5861), .Z(n5864) );
  XOR U5877 ( .A(\knn_comb_/min_val_out[0][11] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .Z(n5861) );
  XOR U5878 ( .A(n119), .B(n5865), .Z(o[10]) );
  AND U5879 ( .A(n122), .B(n5866), .Z(n119) );
  XOR U5880 ( .A(n120), .B(n5865), .Z(n5866) );
  XOR U5881 ( .A(n5867), .B(n5868), .Z(n5865) );
  AND U5882 ( .A(n142), .B(n5869), .Z(n5868) );
  XOR U5883 ( .A(n5870), .B(n49), .Z(n120) );
  AND U5884 ( .A(n125), .B(n5871), .Z(n49) );
  XOR U5885 ( .A(n50), .B(n5870), .Z(n5871) );
  XOR U5886 ( .A(n5872), .B(n5873), .Z(n50) );
  AND U5887 ( .A(n130), .B(n5874), .Z(n5873) );
  XOR U5888 ( .A(p_input[10]), .B(n5872), .Z(n5874) );
  XNOR U5889 ( .A(n5875), .B(n5876), .Z(n5872) );
  AND U5890 ( .A(n134), .B(n5877), .Z(n5876) );
  XOR U5891 ( .A(n5878), .B(n5879), .Z(n5870) );
  AND U5892 ( .A(n138), .B(n5869), .Z(n5879) );
  XNOR U5893 ( .A(n5880), .B(n5867), .Z(n5869) );
  XOR U5894 ( .A(n5881), .B(n5882), .Z(n5867) );
  AND U5895 ( .A(n162), .B(n5883), .Z(n5882) );
  IV U5896 ( .A(n5878), .Z(n5880) );
  XOR U5897 ( .A(n5884), .B(n5885), .Z(n5878) );
  AND U5898 ( .A(n146), .B(n5877), .Z(n5885) );
  XNOR U5899 ( .A(n5875), .B(n5884), .Z(n5877) );
  XNOR U5900 ( .A(n5886), .B(n5887), .Z(n5875) );
  AND U5901 ( .A(n150), .B(n5888), .Z(n5887) );
  XOR U5902 ( .A(p_input[42]), .B(n5886), .Z(n5888) );
  XNOR U5903 ( .A(n5889), .B(n5890), .Z(n5886) );
  AND U5904 ( .A(n154), .B(n5891), .Z(n5890) );
  XOR U5905 ( .A(n5892), .B(n5893), .Z(n5884) );
  AND U5906 ( .A(n158), .B(n5883), .Z(n5893) );
  XNOR U5907 ( .A(n5894), .B(n5881), .Z(n5883) );
  XOR U5908 ( .A(n5895), .B(n5896), .Z(n5881) );
  AND U5909 ( .A(n181), .B(n5897), .Z(n5896) );
  IV U5910 ( .A(n5892), .Z(n5894) );
  XOR U5911 ( .A(n5898), .B(n5899), .Z(n5892) );
  AND U5912 ( .A(n165), .B(n5891), .Z(n5899) );
  XNOR U5913 ( .A(n5889), .B(n5898), .Z(n5891) );
  XNOR U5914 ( .A(n5900), .B(n5901), .Z(n5889) );
  AND U5915 ( .A(n169), .B(n5902), .Z(n5901) );
  XOR U5916 ( .A(p_input[74]), .B(n5900), .Z(n5902) );
  XNOR U5917 ( .A(n5903), .B(n5904), .Z(n5900) );
  AND U5918 ( .A(n173), .B(n5905), .Z(n5904) );
  XOR U5919 ( .A(n5906), .B(n5907), .Z(n5898) );
  AND U5920 ( .A(n177), .B(n5897), .Z(n5907) );
  XNOR U5921 ( .A(n5908), .B(n5895), .Z(n5897) );
  XOR U5922 ( .A(n5909), .B(n5910), .Z(n5895) );
  AND U5923 ( .A(n200), .B(n5911), .Z(n5910) );
  IV U5924 ( .A(n5906), .Z(n5908) );
  XOR U5925 ( .A(n5912), .B(n5913), .Z(n5906) );
  AND U5926 ( .A(n184), .B(n5905), .Z(n5913) );
  XNOR U5927 ( .A(n5903), .B(n5912), .Z(n5905) );
  XNOR U5928 ( .A(n5914), .B(n5915), .Z(n5903) );
  AND U5929 ( .A(n188), .B(n5916), .Z(n5915) );
  XOR U5930 ( .A(p_input[106]), .B(n5914), .Z(n5916) );
  XNOR U5931 ( .A(n5917), .B(n5918), .Z(n5914) );
  AND U5932 ( .A(n192), .B(n5919), .Z(n5918) );
  XOR U5933 ( .A(n5920), .B(n5921), .Z(n5912) );
  AND U5934 ( .A(n196), .B(n5911), .Z(n5921) );
  XNOR U5935 ( .A(n5922), .B(n5909), .Z(n5911) );
  XOR U5936 ( .A(n5923), .B(n5924), .Z(n5909) );
  AND U5937 ( .A(n219), .B(n5925), .Z(n5924) );
  IV U5938 ( .A(n5920), .Z(n5922) );
  XOR U5939 ( .A(n5926), .B(n5927), .Z(n5920) );
  AND U5940 ( .A(n203), .B(n5919), .Z(n5927) );
  XNOR U5941 ( .A(n5917), .B(n5926), .Z(n5919) );
  XNOR U5942 ( .A(n5928), .B(n5929), .Z(n5917) );
  AND U5943 ( .A(n207), .B(n5930), .Z(n5929) );
  XOR U5944 ( .A(p_input[138]), .B(n5928), .Z(n5930) );
  XNOR U5945 ( .A(n5931), .B(n5932), .Z(n5928) );
  AND U5946 ( .A(n211), .B(n5933), .Z(n5932) );
  XOR U5947 ( .A(n5934), .B(n5935), .Z(n5926) );
  AND U5948 ( .A(n215), .B(n5925), .Z(n5935) );
  XNOR U5949 ( .A(n5936), .B(n5923), .Z(n5925) );
  XOR U5950 ( .A(n5937), .B(n5938), .Z(n5923) );
  AND U5951 ( .A(n238), .B(n5939), .Z(n5938) );
  IV U5952 ( .A(n5934), .Z(n5936) );
  XOR U5953 ( .A(n5940), .B(n5941), .Z(n5934) );
  AND U5954 ( .A(n222), .B(n5933), .Z(n5941) );
  XNOR U5955 ( .A(n5931), .B(n5940), .Z(n5933) );
  XNOR U5956 ( .A(n5942), .B(n5943), .Z(n5931) );
  AND U5957 ( .A(n226), .B(n5944), .Z(n5943) );
  XOR U5958 ( .A(p_input[170]), .B(n5942), .Z(n5944) );
  XNOR U5959 ( .A(n5945), .B(n5946), .Z(n5942) );
  AND U5960 ( .A(n230), .B(n5947), .Z(n5946) );
  XOR U5961 ( .A(n5948), .B(n5949), .Z(n5940) );
  AND U5962 ( .A(n234), .B(n5939), .Z(n5949) );
  XNOR U5963 ( .A(n5950), .B(n5937), .Z(n5939) );
  XOR U5964 ( .A(n5951), .B(n5952), .Z(n5937) );
  AND U5965 ( .A(n257), .B(n5953), .Z(n5952) );
  IV U5966 ( .A(n5948), .Z(n5950) );
  XOR U5967 ( .A(n5954), .B(n5955), .Z(n5948) );
  AND U5968 ( .A(n241), .B(n5947), .Z(n5955) );
  XNOR U5969 ( .A(n5945), .B(n5954), .Z(n5947) );
  XNOR U5970 ( .A(n5956), .B(n5957), .Z(n5945) );
  AND U5971 ( .A(n245), .B(n5958), .Z(n5957) );
  XOR U5972 ( .A(p_input[202]), .B(n5956), .Z(n5958) );
  XNOR U5973 ( .A(n5959), .B(n5960), .Z(n5956) );
  AND U5974 ( .A(n249), .B(n5961), .Z(n5960) );
  XOR U5975 ( .A(n5962), .B(n5963), .Z(n5954) );
  AND U5976 ( .A(n253), .B(n5953), .Z(n5963) );
  XNOR U5977 ( .A(n5964), .B(n5951), .Z(n5953) );
  XOR U5978 ( .A(n5965), .B(n5966), .Z(n5951) );
  AND U5979 ( .A(n276), .B(n5967), .Z(n5966) );
  IV U5980 ( .A(n5962), .Z(n5964) );
  XOR U5981 ( .A(n5968), .B(n5969), .Z(n5962) );
  AND U5982 ( .A(n260), .B(n5961), .Z(n5969) );
  XNOR U5983 ( .A(n5959), .B(n5968), .Z(n5961) );
  XNOR U5984 ( .A(n5970), .B(n5971), .Z(n5959) );
  AND U5985 ( .A(n264), .B(n5972), .Z(n5971) );
  XOR U5986 ( .A(p_input[234]), .B(n5970), .Z(n5972) );
  XNOR U5987 ( .A(n5973), .B(n5974), .Z(n5970) );
  AND U5988 ( .A(n268), .B(n5975), .Z(n5974) );
  XOR U5989 ( .A(n5976), .B(n5977), .Z(n5968) );
  AND U5990 ( .A(n272), .B(n5967), .Z(n5977) );
  XNOR U5991 ( .A(n5978), .B(n5965), .Z(n5967) );
  XOR U5992 ( .A(n5979), .B(n5980), .Z(n5965) );
  AND U5993 ( .A(n295), .B(n5981), .Z(n5980) );
  IV U5994 ( .A(n5976), .Z(n5978) );
  XOR U5995 ( .A(n5982), .B(n5983), .Z(n5976) );
  AND U5996 ( .A(n279), .B(n5975), .Z(n5983) );
  XNOR U5997 ( .A(n5973), .B(n5982), .Z(n5975) );
  XNOR U5998 ( .A(n5984), .B(n5985), .Z(n5973) );
  AND U5999 ( .A(n283), .B(n5986), .Z(n5985) );
  XOR U6000 ( .A(p_input[266]), .B(n5984), .Z(n5986) );
  XNOR U6001 ( .A(n5987), .B(n5988), .Z(n5984) );
  AND U6002 ( .A(n287), .B(n5989), .Z(n5988) );
  XOR U6003 ( .A(n5990), .B(n5991), .Z(n5982) );
  AND U6004 ( .A(n291), .B(n5981), .Z(n5991) );
  XNOR U6005 ( .A(n5992), .B(n5979), .Z(n5981) );
  XOR U6006 ( .A(n5993), .B(n5994), .Z(n5979) );
  AND U6007 ( .A(n314), .B(n5995), .Z(n5994) );
  IV U6008 ( .A(n5990), .Z(n5992) );
  XOR U6009 ( .A(n5996), .B(n5997), .Z(n5990) );
  AND U6010 ( .A(n298), .B(n5989), .Z(n5997) );
  XNOR U6011 ( .A(n5987), .B(n5996), .Z(n5989) );
  XNOR U6012 ( .A(n5998), .B(n5999), .Z(n5987) );
  AND U6013 ( .A(n302), .B(n6000), .Z(n5999) );
  XOR U6014 ( .A(p_input[298]), .B(n5998), .Z(n6000) );
  XNOR U6015 ( .A(n6001), .B(n6002), .Z(n5998) );
  AND U6016 ( .A(n306), .B(n6003), .Z(n6002) );
  XOR U6017 ( .A(n6004), .B(n6005), .Z(n5996) );
  AND U6018 ( .A(n310), .B(n5995), .Z(n6005) );
  XNOR U6019 ( .A(n6006), .B(n5993), .Z(n5995) );
  XOR U6020 ( .A(n6007), .B(n6008), .Z(n5993) );
  AND U6021 ( .A(n333), .B(n6009), .Z(n6008) );
  IV U6022 ( .A(n6004), .Z(n6006) );
  XOR U6023 ( .A(n6010), .B(n6011), .Z(n6004) );
  AND U6024 ( .A(n317), .B(n6003), .Z(n6011) );
  XNOR U6025 ( .A(n6001), .B(n6010), .Z(n6003) );
  XNOR U6026 ( .A(n6012), .B(n6013), .Z(n6001) );
  AND U6027 ( .A(n321), .B(n6014), .Z(n6013) );
  XOR U6028 ( .A(p_input[330]), .B(n6012), .Z(n6014) );
  XNOR U6029 ( .A(n6015), .B(n6016), .Z(n6012) );
  AND U6030 ( .A(n325), .B(n6017), .Z(n6016) );
  XOR U6031 ( .A(n6018), .B(n6019), .Z(n6010) );
  AND U6032 ( .A(n329), .B(n6009), .Z(n6019) );
  XNOR U6033 ( .A(n6020), .B(n6007), .Z(n6009) );
  XOR U6034 ( .A(n6021), .B(n6022), .Z(n6007) );
  AND U6035 ( .A(n352), .B(n6023), .Z(n6022) );
  IV U6036 ( .A(n6018), .Z(n6020) );
  XOR U6037 ( .A(n6024), .B(n6025), .Z(n6018) );
  AND U6038 ( .A(n336), .B(n6017), .Z(n6025) );
  XNOR U6039 ( .A(n6015), .B(n6024), .Z(n6017) );
  XNOR U6040 ( .A(n6026), .B(n6027), .Z(n6015) );
  AND U6041 ( .A(n340), .B(n6028), .Z(n6027) );
  XOR U6042 ( .A(p_input[362]), .B(n6026), .Z(n6028) );
  XNOR U6043 ( .A(n6029), .B(n6030), .Z(n6026) );
  AND U6044 ( .A(n344), .B(n6031), .Z(n6030) );
  XOR U6045 ( .A(n6032), .B(n6033), .Z(n6024) );
  AND U6046 ( .A(n348), .B(n6023), .Z(n6033) );
  XNOR U6047 ( .A(n6034), .B(n6021), .Z(n6023) );
  XOR U6048 ( .A(n6035), .B(n6036), .Z(n6021) );
  AND U6049 ( .A(n370), .B(n6037), .Z(n6036) );
  IV U6050 ( .A(n6032), .Z(n6034) );
  XOR U6051 ( .A(n6038), .B(n6039), .Z(n6032) );
  AND U6052 ( .A(n355), .B(n6031), .Z(n6039) );
  XNOR U6053 ( .A(n6029), .B(n6038), .Z(n6031) );
  XNOR U6054 ( .A(n6040), .B(n6041), .Z(n6029) );
  AND U6055 ( .A(n359), .B(n6042), .Z(n6041) );
  XOR U6056 ( .A(p_input[394]), .B(n6040), .Z(n6042) );
  XOR U6057 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n6043), 
        .Z(n6040) );
  AND U6058 ( .A(n362), .B(n6044), .Z(n6043) );
  XOR U6059 ( .A(n6045), .B(n6046), .Z(n6038) );
  AND U6060 ( .A(n366), .B(n6037), .Z(n6046) );
  XNOR U6061 ( .A(n6047), .B(n6035), .Z(n6037) );
  XOR U6062 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n6048), .Z(n6035) );
  AND U6063 ( .A(n378), .B(n6049), .Z(n6048) );
  IV U6064 ( .A(n6045), .Z(n6047) );
  XOR U6065 ( .A(n6050), .B(n6051), .Z(n6045) );
  AND U6066 ( .A(n373), .B(n6044), .Z(n6051) );
  XOR U6067 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n6050), 
        .Z(n6044) );
  XOR U6068 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(n6052), 
        .Z(n6050) );
  AND U6069 ( .A(n375), .B(n6049), .Z(n6052) );
  XOR U6070 ( .A(\knn_comb_/min_val_out[0][10] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .Z(n6049) );
  XOR U6071 ( .A(n1523), .B(n6053), .Z(o[0]) );
  AND U6072 ( .A(n122), .B(n6054), .Z(n1523) );
  XOR U6073 ( .A(n1524), .B(n6053), .Z(n6054) );
  XOR U6074 ( .A(n6055), .B(n6056), .Z(n6053) );
  AND U6075 ( .A(n142), .B(n6057), .Z(n6056) );
  XOR U6076 ( .A(n6058), .B(n71), .Z(n1524) );
  AND U6077 ( .A(n125), .B(n6059), .Z(n71) );
  XOR U6078 ( .A(n72), .B(n6058), .Z(n6059) );
  XOR U6079 ( .A(n6060), .B(n6061), .Z(n72) );
  AND U6080 ( .A(n130), .B(n6062), .Z(n6061) );
  XOR U6081 ( .A(p_input[0]), .B(n6060), .Z(n6062) );
  XNOR U6082 ( .A(n6063), .B(n6064), .Z(n6060) );
  AND U6083 ( .A(n134), .B(n6065), .Z(n6064) );
  XOR U6084 ( .A(n6066), .B(n6067), .Z(n6058) );
  AND U6085 ( .A(n138), .B(n6057), .Z(n6067) );
  XNOR U6086 ( .A(n6068), .B(n6055), .Z(n6057) );
  XOR U6087 ( .A(n6069), .B(n6070), .Z(n6055) );
  AND U6088 ( .A(n162), .B(n6071), .Z(n6070) );
  IV U6089 ( .A(n6066), .Z(n6068) );
  XOR U6090 ( .A(n6072), .B(n6073), .Z(n6066) );
  AND U6091 ( .A(n146), .B(n6065), .Z(n6073) );
  XNOR U6092 ( .A(n6063), .B(n6072), .Z(n6065) );
  XNOR U6093 ( .A(n6074), .B(n6075), .Z(n6063) );
  AND U6094 ( .A(n150), .B(n6076), .Z(n6075) );
  XOR U6095 ( .A(p_input[32]), .B(n6074), .Z(n6076) );
  XNOR U6096 ( .A(n6077), .B(n6078), .Z(n6074) );
  AND U6097 ( .A(n154), .B(n6079), .Z(n6078) );
  XOR U6098 ( .A(n6080), .B(n6081), .Z(n6072) );
  AND U6099 ( .A(n158), .B(n6071), .Z(n6081) );
  XNOR U6100 ( .A(n6082), .B(n6069), .Z(n6071) );
  XOR U6101 ( .A(n6083), .B(n6084), .Z(n6069) );
  AND U6102 ( .A(n181), .B(n6085), .Z(n6084) );
  IV U6103 ( .A(n6080), .Z(n6082) );
  XOR U6104 ( .A(n6086), .B(n6087), .Z(n6080) );
  AND U6105 ( .A(n165), .B(n6079), .Z(n6087) );
  XNOR U6106 ( .A(n6077), .B(n6086), .Z(n6079) );
  XNOR U6107 ( .A(n6088), .B(n6089), .Z(n6077) );
  AND U6108 ( .A(n169), .B(n6090), .Z(n6089) );
  XOR U6109 ( .A(p_input[64]), .B(n6088), .Z(n6090) );
  XNOR U6110 ( .A(n6091), .B(n6092), .Z(n6088) );
  AND U6111 ( .A(n173), .B(n6093), .Z(n6092) );
  XOR U6112 ( .A(n6094), .B(n6095), .Z(n6086) );
  AND U6113 ( .A(n177), .B(n6085), .Z(n6095) );
  XNOR U6114 ( .A(n6096), .B(n6083), .Z(n6085) );
  XOR U6115 ( .A(n6097), .B(n6098), .Z(n6083) );
  AND U6116 ( .A(n200), .B(n6099), .Z(n6098) );
  IV U6117 ( .A(n6094), .Z(n6096) );
  XOR U6118 ( .A(n6100), .B(n6101), .Z(n6094) );
  AND U6119 ( .A(n184), .B(n6093), .Z(n6101) );
  XNOR U6120 ( .A(n6091), .B(n6100), .Z(n6093) );
  XNOR U6121 ( .A(n6102), .B(n6103), .Z(n6091) );
  AND U6122 ( .A(n188), .B(n6104), .Z(n6103) );
  XOR U6123 ( .A(p_input[96]), .B(n6102), .Z(n6104) );
  XNOR U6124 ( .A(n6105), .B(n6106), .Z(n6102) );
  AND U6125 ( .A(n192), .B(n6107), .Z(n6106) );
  XOR U6126 ( .A(n6108), .B(n6109), .Z(n6100) );
  AND U6127 ( .A(n196), .B(n6099), .Z(n6109) );
  XNOR U6128 ( .A(n6110), .B(n6097), .Z(n6099) );
  XOR U6129 ( .A(n6111), .B(n6112), .Z(n6097) );
  AND U6130 ( .A(n219), .B(n6113), .Z(n6112) );
  IV U6131 ( .A(n6108), .Z(n6110) );
  XOR U6132 ( .A(n6114), .B(n6115), .Z(n6108) );
  AND U6133 ( .A(n203), .B(n6107), .Z(n6115) );
  XNOR U6134 ( .A(n6105), .B(n6114), .Z(n6107) );
  XNOR U6135 ( .A(n6116), .B(n6117), .Z(n6105) );
  AND U6136 ( .A(n207), .B(n6118), .Z(n6117) );
  XOR U6137 ( .A(p_input[128]), .B(n6116), .Z(n6118) );
  XNOR U6138 ( .A(n6119), .B(n6120), .Z(n6116) );
  AND U6139 ( .A(n211), .B(n6121), .Z(n6120) );
  XOR U6140 ( .A(n6122), .B(n6123), .Z(n6114) );
  AND U6141 ( .A(n215), .B(n6113), .Z(n6123) );
  XNOR U6142 ( .A(n6124), .B(n6111), .Z(n6113) );
  XOR U6143 ( .A(n6125), .B(n6126), .Z(n6111) );
  AND U6144 ( .A(n238), .B(n6127), .Z(n6126) );
  IV U6145 ( .A(n6122), .Z(n6124) );
  XOR U6146 ( .A(n6128), .B(n6129), .Z(n6122) );
  AND U6147 ( .A(n222), .B(n6121), .Z(n6129) );
  XNOR U6148 ( .A(n6119), .B(n6128), .Z(n6121) );
  XNOR U6149 ( .A(n6130), .B(n6131), .Z(n6119) );
  AND U6150 ( .A(n226), .B(n6132), .Z(n6131) );
  XOR U6151 ( .A(p_input[160]), .B(n6130), .Z(n6132) );
  XNOR U6152 ( .A(n6133), .B(n6134), .Z(n6130) );
  AND U6153 ( .A(n230), .B(n6135), .Z(n6134) );
  XOR U6154 ( .A(n6136), .B(n6137), .Z(n6128) );
  AND U6155 ( .A(n234), .B(n6127), .Z(n6137) );
  XNOR U6156 ( .A(n6138), .B(n6125), .Z(n6127) );
  XOR U6157 ( .A(n6139), .B(n6140), .Z(n6125) );
  AND U6158 ( .A(n257), .B(n6141), .Z(n6140) );
  IV U6159 ( .A(n6136), .Z(n6138) );
  XOR U6160 ( .A(n6142), .B(n6143), .Z(n6136) );
  AND U6161 ( .A(n241), .B(n6135), .Z(n6143) );
  XNOR U6162 ( .A(n6133), .B(n6142), .Z(n6135) );
  XNOR U6163 ( .A(n6144), .B(n6145), .Z(n6133) );
  AND U6164 ( .A(n245), .B(n6146), .Z(n6145) );
  XOR U6165 ( .A(p_input[192]), .B(n6144), .Z(n6146) );
  XNOR U6166 ( .A(n6147), .B(n6148), .Z(n6144) );
  AND U6167 ( .A(n249), .B(n6149), .Z(n6148) );
  XOR U6168 ( .A(n6150), .B(n6151), .Z(n6142) );
  AND U6169 ( .A(n253), .B(n6141), .Z(n6151) );
  XNOR U6170 ( .A(n6152), .B(n6139), .Z(n6141) );
  XOR U6171 ( .A(n6153), .B(n6154), .Z(n6139) );
  AND U6172 ( .A(n276), .B(n6155), .Z(n6154) );
  IV U6173 ( .A(n6150), .Z(n6152) );
  XOR U6174 ( .A(n6156), .B(n6157), .Z(n6150) );
  AND U6175 ( .A(n260), .B(n6149), .Z(n6157) );
  XNOR U6176 ( .A(n6147), .B(n6156), .Z(n6149) );
  XNOR U6177 ( .A(n6158), .B(n6159), .Z(n6147) );
  AND U6178 ( .A(n264), .B(n6160), .Z(n6159) );
  XOR U6179 ( .A(p_input[224]), .B(n6158), .Z(n6160) );
  XNOR U6180 ( .A(n6161), .B(n6162), .Z(n6158) );
  AND U6181 ( .A(n268), .B(n6163), .Z(n6162) );
  XOR U6182 ( .A(n6164), .B(n6165), .Z(n6156) );
  AND U6183 ( .A(n272), .B(n6155), .Z(n6165) );
  XNOR U6184 ( .A(n6166), .B(n6153), .Z(n6155) );
  XOR U6185 ( .A(n6167), .B(n6168), .Z(n6153) );
  AND U6186 ( .A(n295), .B(n6169), .Z(n6168) );
  IV U6187 ( .A(n6164), .Z(n6166) );
  XOR U6188 ( .A(n6170), .B(n6171), .Z(n6164) );
  AND U6189 ( .A(n279), .B(n6163), .Z(n6171) );
  XNOR U6190 ( .A(n6161), .B(n6170), .Z(n6163) );
  XNOR U6191 ( .A(n6172), .B(n6173), .Z(n6161) );
  AND U6192 ( .A(n283), .B(n6174), .Z(n6173) );
  XOR U6193 ( .A(p_input[256]), .B(n6172), .Z(n6174) );
  XNOR U6194 ( .A(n6175), .B(n6176), .Z(n6172) );
  AND U6195 ( .A(n287), .B(n6177), .Z(n6176) );
  XOR U6196 ( .A(n6178), .B(n6179), .Z(n6170) );
  AND U6197 ( .A(n291), .B(n6169), .Z(n6179) );
  XNOR U6198 ( .A(n6180), .B(n6167), .Z(n6169) );
  XOR U6199 ( .A(n6181), .B(n6182), .Z(n6167) );
  AND U6200 ( .A(n314), .B(n6183), .Z(n6182) );
  IV U6201 ( .A(n6178), .Z(n6180) );
  XOR U6202 ( .A(n6184), .B(n6185), .Z(n6178) );
  AND U6203 ( .A(n298), .B(n6177), .Z(n6185) );
  XNOR U6204 ( .A(n6175), .B(n6184), .Z(n6177) );
  XNOR U6205 ( .A(n6186), .B(n6187), .Z(n6175) );
  AND U6206 ( .A(n302), .B(n6188), .Z(n6187) );
  XOR U6207 ( .A(p_input[288]), .B(n6186), .Z(n6188) );
  XNOR U6208 ( .A(n6189), .B(n6190), .Z(n6186) );
  AND U6209 ( .A(n306), .B(n6191), .Z(n6190) );
  XOR U6210 ( .A(n6192), .B(n6193), .Z(n6184) );
  AND U6211 ( .A(n310), .B(n6183), .Z(n6193) );
  XNOR U6212 ( .A(n6194), .B(n6181), .Z(n6183) );
  XOR U6213 ( .A(n6195), .B(n6196), .Z(n6181) );
  AND U6214 ( .A(n333), .B(n6197), .Z(n6196) );
  IV U6215 ( .A(n6192), .Z(n6194) );
  XOR U6216 ( .A(n6198), .B(n6199), .Z(n6192) );
  AND U6217 ( .A(n317), .B(n6191), .Z(n6199) );
  XNOR U6218 ( .A(n6189), .B(n6198), .Z(n6191) );
  XNOR U6219 ( .A(n6200), .B(n6201), .Z(n6189) );
  AND U6220 ( .A(n321), .B(n6202), .Z(n6201) );
  XOR U6221 ( .A(p_input[320]), .B(n6200), .Z(n6202) );
  XNOR U6222 ( .A(n6203), .B(n6204), .Z(n6200) );
  AND U6223 ( .A(n325), .B(n6205), .Z(n6204) );
  XOR U6224 ( .A(n6206), .B(n6207), .Z(n6198) );
  AND U6225 ( .A(n329), .B(n6197), .Z(n6207) );
  XNOR U6226 ( .A(n6208), .B(n6195), .Z(n6197) );
  XOR U6227 ( .A(n6209), .B(n6210), .Z(n6195) );
  AND U6228 ( .A(n352), .B(n6211), .Z(n6210) );
  IV U6229 ( .A(n6206), .Z(n6208) );
  XOR U6230 ( .A(n6212), .B(n6213), .Z(n6206) );
  AND U6231 ( .A(n336), .B(n6205), .Z(n6213) );
  XNOR U6232 ( .A(n6203), .B(n6212), .Z(n6205) );
  XNOR U6233 ( .A(n6214), .B(n6215), .Z(n6203) );
  AND U6234 ( .A(n340), .B(n6216), .Z(n6215) );
  XOR U6235 ( .A(p_input[352]), .B(n6214), .Z(n6216) );
  XNOR U6236 ( .A(n6217), .B(n6218), .Z(n6214) );
  AND U6237 ( .A(n344), .B(n6219), .Z(n6218) );
  XOR U6238 ( .A(n6220), .B(n6221), .Z(n6212) );
  AND U6239 ( .A(n348), .B(n6211), .Z(n6221) );
  XNOR U6240 ( .A(n6222), .B(n6209), .Z(n6211) );
  XOR U6241 ( .A(n6223), .B(n6224), .Z(n6209) );
  AND U6242 ( .A(n370), .B(n6225), .Z(n6224) );
  IV U6243 ( .A(n6220), .Z(n6222) );
  XOR U6244 ( .A(n6226), .B(n6227), .Z(n6220) );
  AND U6245 ( .A(n355), .B(n6219), .Z(n6227) );
  XNOR U6246 ( .A(n6217), .B(n6226), .Z(n6219) );
  XNOR U6247 ( .A(n6228), .B(n6229), .Z(n6217) );
  AND U6248 ( .A(n359), .B(n6230), .Z(n6229) );
  XOR U6249 ( .A(p_input[384]), .B(n6228), .Z(n6230) );
  XOR U6250 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(n6231), 
        .Z(n6228) );
  AND U6251 ( .A(n362), .B(n6232), .Z(n6231) );
  XOR U6252 ( .A(n6233), .B(n6234), .Z(n6226) );
  AND U6253 ( .A(n366), .B(n6225), .Z(n6234) );
  XNOR U6254 ( .A(n6235), .B(n6223), .Z(n6225) );
  XOR U6255 ( .A(\knn_comb_/min_val_out[0][0] ), .B(n6236), .Z(n6223) );
  AND U6256 ( .A(n378), .B(n6237), .Z(n6236) );
  IV U6257 ( .A(n6233), .Z(n6235) );
  XOR U6258 ( .A(n6238), .B(n6239), .Z(n6233) );
  AND U6259 ( .A(n373), .B(n6232), .Z(n6239) );
  XOR U6260 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(n6238), 
        .Z(n6232) );
  XOR U6261 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(n6240), 
        .Z(n6238) );
  AND U6262 ( .A(n375), .B(n6237), .Z(n6240) );
  XOR U6263 ( .A(\knn_comb_/min_val_out[0][0] ), .B(
        \knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .Z(n6237) );
  XNOR U6264 ( .A(n6241), .B(n6242), .Z(n122) );
  AND U6265 ( .A(n6243), .B(n6244), .Z(n6242) );
  XNOR U6266 ( .A(n6241), .B(n6245), .Z(n6244) );
  XOR U6267 ( .A(n6246), .B(n6247), .Z(n6245) );
  AND U6268 ( .A(n125), .B(n6248), .Z(n6247) );
  XNOR U6269 ( .A(n6246), .B(n6249), .Z(n6248) );
  IV U6270 ( .A(n6250), .Z(n6246) );
  XNOR U6271 ( .A(n6241), .B(n6251), .Z(n6243) );
  XOR U6272 ( .A(n6252), .B(n6253), .Z(n6251) );
  AND U6273 ( .A(n142), .B(n6254), .Z(n6253) );
  XOR U6274 ( .A(n6255), .B(n6256), .Z(n6241) );
  AND U6275 ( .A(n6257), .B(n6258), .Z(n6256) );
  XOR U6276 ( .A(n6259), .B(n6255), .Z(n6258) );
  XNOR U6277 ( .A(n6260), .B(n6261), .Z(n6259) );
  AND U6278 ( .A(n125), .B(n6262), .Z(n6261) );
  XNOR U6279 ( .A(n6263), .B(n6260), .Z(n6262) );
  XNOR U6280 ( .A(n6255), .B(n6264), .Z(n6257) );
  XOR U6281 ( .A(n6265), .B(n6266), .Z(n6264) );
  AND U6282 ( .A(n142), .B(n6267), .Z(n6266) );
  XOR U6283 ( .A(n6268), .B(n6269), .Z(n6255) );
  AND U6284 ( .A(n6270), .B(n6271), .Z(n6269) );
  XOR U6285 ( .A(n6272), .B(n6268), .Z(n6271) );
  XNOR U6286 ( .A(n6273), .B(n6274), .Z(n6272) );
  AND U6287 ( .A(n125), .B(n6275), .Z(n6274) );
  XNOR U6288 ( .A(n6276), .B(n6273), .Z(n6275) );
  XNOR U6289 ( .A(n6268), .B(n6277), .Z(n6270) );
  XOR U6290 ( .A(n6278), .B(n6279), .Z(n6277) );
  AND U6291 ( .A(n142), .B(n6280), .Z(n6279) );
  XOR U6292 ( .A(n6281), .B(n6282), .Z(n6268) );
  AND U6293 ( .A(n6283), .B(n6284), .Z(n6282) );
  XOR U6294 ( .A(n6285), .B(n6281), .Z(n6284) );
  XNOR U6295 ( .A(n6286), .B(n6287), .Z(n6285) );
  AND U6296 ( .A(n125), .B(n6288), .Z(n6287) );
  XNOR U6297 ( .A(n6289), .B(n6286), .Z(n6288) );
  XNOR U6298 ( .A(n6281), .B(n6290), .Z(n6283) );
  XOR U6299 ( .A(n6291), .B(n6292), .Z(n6290) );
  AND U6300 ( .A(n142), .B(n6293), .Z(n6292) );
  XOR U6301 ( .A(n6294), .B(n6295), .Z(n6281) );
  AND U6302 ( .A(n6296), .B(n6297), .Z(n6295) );
  XOR U6303 ( .A(n6294), .B(n6298), .Z(n6297) );
  XOR U6304 ( .A(n6299), .B(n6300), .Z(n6298) );
  AND U6305 ( .A(n125), .B(n6301), .Z(n6300) );
  XOR U6306 ( .A(n6302), .B(n6299), .Z(n6301) );
  XNOR U6307 ( .A(n6303), .B(n6294), .Z(n6296) );
  XNOR U6308 ( .A(n6304), .B(n6305), .Z(n6303) );
  AND U6309 ( .A(n142), .B(n6306), .Z(n6305) );
  AND U6310 ( .A(n6307), .B(n6308), .Z(n6294) );
  XNOR U6311 ( .A(n6309), .B(n6310), .Z(n6308) );
  AND U6312 ( .A(n125), .B(n6311), .Z(n6310) );
  XNOR U6313 ( .A(n6312), .B(n6309), .Z(n6311) );
  XNOR U6314 ( .A(n6313), .B(n6314), .Z(n125) );
  AND U6315 ( .A(n6315), .B(n6316), .Z(n6314) );
  XOR U6316 ( .A(n6249), .B(n6313), .Z(n6316) );
  XOR U6317 ( .A(n6317), .B(n6318), .Z(n6249) );
  AND U6318 ( .A(n130), .B(n6319), .Z(n6318) );
  XOR U6319 ( .A(n6320), .B(n6317), .Z(n6319) );
  XNOR U6320 ( .A(n6250), .B(n6313), .Z(n6315) );
  XOR U6321 ( .A(n6321), .B(n6322), .Z(n6250) );
  AND U6322 ( .A(n138), .B(n6254), .Z(n6322) );
  XOR U6323 ( .A(n6252), .B(n6321), .Z(n6254) );
  XOR U6324 ( .A(n6323), .B(n6324), .Z(n6313) );
  AND U6325 ( .A(n6325), .B(n6326), .Z(n6324) );
  XOR U6326 ( .A(n6263), .B(n6323), .Z(n6326) );
  XOR U6327 ( .A(n6327), .B(n6328), .Z(n6263) );
  AND U6328 ( .A(n130), .B(n6329), .Z(n6328) );
  XOR U6329 ( .A(n6330), .B(n6327), .Z(n6329) );
  XOR U6330 ( .A(n6323), .B(n6260), .Z(n6325) );
  XOR U6331 ( .A(n6331), .B(n6332), .Z(n6260) );
  AND U6332 ( .A(n138), .B(n6267), .Z(n6332) );
  XOR U6333 ( .A(n6331), .B(n6333), .Z(n6267) );
  XOR U6334 ( .A(n6334), .B(n6335), .Z(n6323) );
  AND U6335 ( .A(n6336), .B(n6337), .Z(n6335) );
  XOR U6336 ( .A(n6276), .B(n6334), .Z(n6337) );
  XOR U6337 ( .A(n6338), .B(n6339), .Z(n6276) );
  AND U6338 ( .A(n130), .B(n6340), .Z(n6339) );
  XNOR U6339 ( .A(n6341), .B(n6338), .Z(n6340) );
  XOR U6340 ( .A(n6334), .B(n6273), .Z(n6336) );
  XOR U6341 ( .A(n6342), .B(n6343), .Z(n6273) );
  AND U6342 ( .A(n138), .B(n6280), .Z(n6343) );
  XOR U6343 ( .A(n6342), .B(n6344), .Z(n6280) );
  XOR U6344 ( .A(n6345), .B(n6346), .Z(n6334) );
  AND U6345 ( .A(n6347), .B(n6348), .Z(n6346) );
  XOR U6346 ( .A(n6289), .B(n6345), .Z(n6348) );
  XOR U6347 ( .A(n6349), .B(n6350), .Z(n6289) );
  AND U6348 ( .A(n130), .B(n6351), .Z(n6350) );
  XOR U6349 ( .A(n6352), .B(n6349), .Z(n6351) );
  XOR U6350 ( .A(n6345), .B(n6286), .Z(n6347) );
  XOR U6351 ( .A(n6353), .B(n6354), .Z(n6286) );
  AND U6352 ( .A(n138), .B(n6293), .Z(n6354) );
  XOR U6353 ( .A(n6353), .B(n6355), .Z(n6293) );
  XOR U6354 ( .A(n6356), .B(n6357), .Z(n6345) );
  AND U6355 ( .A(n6358), .B(n6359), .Z(n6357) );
  XOR U6356 ( .A(n6356), .B(n6302), .Z(n6359) );
  XOR U6357 ( .A(n6360), .B(n6361), .Z(n6302) );
  AND U6358 ( .A(n130), .B(n6362), .Z(n6361) );
  XNOR U6359 ( .A(n6363), .B(n6360), .Z(n6362) );
  XNOR U6360 ( .A(n6299), .B(n6356), .Z(n6358) );
  XNOR U6361 ( .A(n6364), .B(n6365), .Z(n6299) );
  AND U6362 ( .A(n138), .B(n6306), .Z(n6365) );
  XOR U6363 ( .A(n6364), .B(n6304), .Z(n6306) );
  AND U6364 ( .A(n6309), .B(n6312), .Z(n6356) );
  XOR U6365 ( .A(n6366), .B(n6367), .Z(n6312) );
  AND U6366 ( .A(n130), .B(n6368), .Z(n6367) );
  XNOR U6367 ( .A(n6369), .B(n6370), .Z(n6368) );
  XNOR U6368 ( .A(n6371), .B(n6372), .Z(n130) );
  AND U6369 ( .A(n6373), .B(n6374), .Z(n6372) );
  XOR U6370 ( .A(n6320), .B(n6371), .Z(n6374) );
  AND U6371 ( .A(n6375), .B(n6376), .Z(n6320) );
  XNOR U6372 ( .A(n6317), .B(n6371), .Z(n6373) );
  XNOR U6373 ( .A(n6377), .B(n6378), .Z(n6317) );
  AND U6374 ( .A(n134), .B(n6379), .Z(n6378) );
  XNOR U6375 ( .A(n6380), .B(n6381), .Z(n6379) );
  XOR U6376 ( .A(n6382), .B(n6383), .Z(n6371) );
  AND U6377 ( .A(n6384), .B(n6385), .Z(n6383) );
  XNOR U6378 ( .A(n6382), .B(n6375), .Z(n6385) );
  IV U6379 ( .A(n6330), .Z(n6375) );
  XOR U6380 ( .A(n6386), .B(n6387), .Z(n6330) );
  XOR U6381 ( .A(n6388), .B(n6376), .Z(n6387) );
  AND U6382 ( .A(n6341), .B(n6389), .Z(n6376) );
  AND U6383 ( .A(n6390), .B(n6391), .Z(n6388) );
  XOR U6384 ( .A(n6392), .B(n6386), .Z(n6390) );
  XNOR U6385 ( .A(n6327), .B(n6382), .Z(n6384) );
  XNOR U6386 ( .A(n6393), .B(n6394), .Z(n6327) );
  AND U6387 ( .A(n134), .B(n6395), .Z(n6394) );
  XNOR U6388 ( .A(n6396), .B(n6397), .Z(n6395) );
  XOR U6389 ( .A(n6398), .B(n6399), .Z(n6382) );
  AND U6390 ( .A(n6400), .B(n6401), .Z(n6399) );
  XNOR U6391 ( .A(n6398), .B(n6341), .Z(n6401) );
  XOR U6392 ( .A(n6402), .B(n6391), .Z(n6341) );
  XNOR U6393 ( .A(n6403), .B(n6386), .Z(n6391) );
  XOR U6394 ( .A(n6404), .B(n6405), .Z(n6386) );
  AND U6395 ( .A(n6406), .B(n6407), .Z(n6405) );
  XOR U6396 ( .A(n6408), .B(n6404), .Z(n6406) );
  XNOR U6397 ( .A(n6409), .B(n6410), .Z(n6403) );
  AND U6398 ( .A(n6411), .B(n6412), .Z(n6410) );
  XOR U6399 ( .A(n6409), .B(n6413), .Z(n6411) );
  XNOR U6400 ( .A(n6392), .B(n6389), .Z(n6402) );
  AND U6401 ( .A(n6414), .B(n6415), .Z(n6389) );
  XOR U6402 ( .A(n6416), .B(n6417), .Z(n6392) );
  AND U6403 ( .A(n6418), .B(n6419), .Z(n6417) );
  XOR U6404 ( .A(n6416), .B(n6420), .Z(n6418) );
  XNOR U6405 ( .A(n6338), .B(n6398), .Z(n6400) );
  XNOR U6406 ( .A(n6421), .B(n6422), .Z(n6338) );
  AND U6407 ( .A(n134), .B(n6423), .Z(n6422) );
  XNOR U6408 ( .A(n6424), .B(n6425), .Z(n6423) );
  XOR U6409 ( .A(n6426), .B(n6427), .Z(n6398) );
  AND U6410 ( .A(n6428), .B(n6429), .Z(n6427) );
  XNOR U6411 ( .A(n6426), .B(n6414), .Z(n6429) );
  IV U6412 ( .A(n6352), .Z(n6414) );
  XNOR U6413 ( .A(n6430), .B(n6407), .Z(n6352) );
  XNOR U6414 ( .A(n6431), .B(n6413), .Z(n6407) );
  XOR U6415 ( .A(n6432), .B(n6433), .Z(n6413) );
  AND U6416 ( .A(n6434), .B(n6435), .Z(n6433) );
  XOR U6417 ( .A(n6432), .B(n6436), .Z(n6434) );
  XNOR U6418 ( .A(n6412), .B(n6404), .Z(n6431) );
  XOR U6419 ( .A(n6437), .B(n6438), .Z(n6404) );
  AND U6420 ( .A(n6439), .B(n6440), .Z(n6438) );
  XNOR U6421 ( .A(n6441), .B(n6437), .Z(n6439) );
  XNOR U6422 ( .A(n6442), .B(n6409), .Z(n6412) );
  XOR U6423 ( .A(n6443), .B(n6444), .Z(n6409) );
  AND U6424 ( .A(n6445), .B(n6446), .Z(n6444) );
  XOR U6425 ( .A(n6443), .B(n6447), .Z(n6445) );
  XNOR U6426 ( .A(n6448), .B(n6449), .Z(n6442) );
  AND U6427 ( .A(n6450), .B(n6451), .Z(n6449) );
  XNOR U6428 ( .A(n6448), .B(n6452), .Z(n6450) );
  XNOR U6429 ( .A(n6408), .B(n6415), .Z(n6430) );
  AND U6430 ( .A(n6363), .B(n6453), .Z(n6415) );
  XOR U6431 ( .A(n6420), .B(n6419), .Z(n6408) );
  XNOR U6432 ( .A(n6454), .B(n6416), .Z(n6419) );
  XOR U6433 ( .A(n6455), .B(n6456), .Z(n6416) );
  AND U6434 ( .A(n6457), .B(n6458), .Z(n6456) );
  XOR U6435 ( .A(n6455), .B(n6459), .Z(n6457) );
  XNOR U6436 ( .A(n6460), .B(n6461), .Z(n6454) );
  AND U6437 ( .A(n6462), .B(n6463), .Z(n6461) );
  XOR U6438 ( .A(n6460), .B(n6464), .Z(n6462) );
  XOR U6439 ( .A(n6465), .B(n6466), .Z(n6420) );
  AND U6440 ( .A(n6467), .B(n6468), .Z(n6466) );
  XOR U6441 ( .A(n6465), .B(n6469), .Z(n6467) );
  XNOR U6442 ( .A(n6349), .B(n6426), .Z(n6428) );
  XNOR U6443 ( .A(n6470), .B(n6471), .Z(n6349) );
  AND U6444 ( .A(n134), .B(n6472), .Z(n6471) );
  XNOR U6445 ( .A(n6473), .B(n6474), .Z(n6472) );
  XOR U6446 ( .A(n6475), .B(n6476), .Z(n6426) );
  AND U6447 ( .A(n6477), .B(n6478), .Z(n6476) );
  XNOR U6448 ( .A(n6475), .B(n6363), .Z(n6478) );
  XOR U6449 ( .A(n6479), .B(n6440), .Z(n6363) );
  XNOR U6450 ( .A(n6480), .B(n6447), .Z(n6440) );
  XOR U6451 ( .A(n6436), .B(n6435), .Z(n6447) );
  XNOR U6452 ( .A(n6481), .B(n6432), .Z(n6435) );
  XOR U6453 ( .A(n6482), .B(n6483), .Z(n6432) );
  AND U6454 ( .A(n6484), .B(n6485), .Z(n6483) );
  XNOR U6455 ( .A(n6486), .B(n6487), .Z(n6484) );
  IV U6456 ( .A(n6482), .Z(n6486) );
  XNOR U6457 ( .A(n6488), .B(n6489), .Z(n6481) );
  NOR U6458 ( .A(n6490), .B(n6491), .Z(n6489) );
  XNOR U6459 ( .A(n6488), .B(n6492), .Z(n6490) );
  XOR U6460 ( .A(n6493), .B(n6494), .Z(n6436) );
  NOR U6461 ( .A(n6495), .B(n6496), .Z(n6494) );
  XNOR U6462 ( .A(n6493), .B(n6497), .Z(n6495) );
  XNOR U6463 ( .A(n6446), .B(n6437), .Z(n6480) );
  XOR U6464 ( .A(n6498), .B(n6499), .Z(n6437) );
  AND U6465 ( .A(n6500), .B(n6501), .Z(n6499) );
  XOR U6466 ( .A(n6498), .B(n6502), .Z(n6500) );
  XOR U6467 ( .A(n6503), .B(n6452), .Z(n6446) );
  XOR U6468 ( .A(n6504), .B(n6505), .Z(n6452) );
  NOR U6469 ( .A(n6506), .B(n6507), .Z(n6505) );
  XOR U6470 ( .A(n6504), .B(n6508), .Z(n6506) );
  XNOR U6471 ( .A(n6451), .B(n6443), .Z(n6503) );
  XOR U6472 ( .A(n6509), .B(n6510), .Z(n6443) );
  AND U6473 ( .A(n6511), .B(n6512), .Z(n6510) );
  XOR U6474 ( .A(n6509), .B(n6513), .Z(n6511) );
  XNOR U6475 ( .A(n6514), .B(n6448), .Z(n6451) );
  XOR U6476 ( .A(n6515), .B(n6516), .Z(n6448) );
  AND U6477 ( .A(n6517), .B(n6518), .Z(n6516) );
  XNOR U6478 ( .A(n6519), .B(n6520), .Z(n6517) );
  IV U6479 ( .A(n6515), .Z(n6519) );
  XNOR U6480 ( .A(n6521), .B(n6522), .Z(n6514) );
  NOR U6481 ( .A(n6523), .B(n6524), .Z(n6522) );
  XNOR U6482 ( .A(n6521), .B(n6525), .Z(n6523) );
  XOR U6483 ( .A(n6441), .B(n6453), .Z(n6479) );
  NOR U6484 ( .A(n6369), .B(n6526), .Z(n6453) );
  XNOR U6485 ( .A(n6459), .B(n6458), .Z(n6441) );
  XNOR U6486 ( .A(n6527), .B(n6464), .Z(n6458) );
  XNOR U6487 ( .A(n6528), .B(n6529), .Z(n6464) );
  NOR U6488 ( .A(n6530), .B(n6531), .Z(n6529) );
  XOR U6489 ( .A(n6528), .B(n6532), .Z(n6530) );
  XNOR U6490 ( .A(n6463), .B(n6455), .Z(n6527) );
  XOR U6491 ( .A(n6533), .B(n6534), .Z(n6455) );
  AND U6492 ( .A(n6535), .B(n6536), .Z(n6534) );
  XNOR U6493 ( .A(n6533), .B(n6537), .Z(n6535) );
  XNOR U6494 ( .A(n6538), .B(n6460), .Z(n6463) );
  XOR U6495 ( .A(n6539), .B(n6540), .Z(n6460) );
  AND U6496 ( .A(n6541), .B(n6542), .Z(n6540) );
  XNOR U6497 ( .A(n6543), .B(n6544), .Z(n6541) );
  IV U6498 ( .A(n6539), .Z(n6543) );
  XNOR U6499 ( .A(n6545), .B(n6546), .Z(n6538) );
  NOR U6500 ( .A(n6547), .B(n6548), .Z(n6546) );
  XNOR U6501 ( .A(n6545), .B(n6549), .Z(n6547) );
  XOR U6502 ( .A(n6469), .B(n6468), .Z(n6459) );
  XNOR U6503 ( .A(n6550), .B(n6465), .Z(n6468) );
  XOR U6504 ( .A(n6551), .B(n6552), .Z(n6465) );
  AND U6505 ( .A(n6553), .B(n6554), .Z(n6552) );
  XNOR U6506 ( .A(n6555), .B(n6556), .Z(n6553) );
  IV U6507 ( .A(n6551), .Z(n6555) );
  XNOR U6508 ( .A(n6557), .B(n6558), .Z(n6550) );
  NOR U6509 ( .A(n6559), .B(n6560), .Z(n6558) );
  XNOR U6510 ( .A(n6557), .B(n6561), .Z(n6559) );
  XOR U6511 ( .A(n6562), .B(n6563), .Z(n6469) );
  NOR U6512 ( .A(n6564), .B(n6565), .Z(n6563) );
  XNOR U6513 ( .A(n6562), .B(n6566), .Z(n6564) );
  XNOR U6514 ( .A(n6360), .B(n6475), .Z(n6477) );
  XNOR U6515 ( .A(n6567), .B(n6568), .Z(n6360) );
  AND U6516 ( .A(n134), .B(n6569), .Z(n6568) );
  XNOR U6517 ( .A(n6570), .B(n6571), .Z(n6569) );
  AND U6518 ( .A(n6370), .B(n6369), .Z(n6475) );
  XOR U6519 ( .A(n6572), .B(n6526), .Z(n6369) );
  XNOR U6520 ( .A(p_input[0]), .B(p_input[512]), .Z(n6526) );
  XNOR U6521 ( .A(n6502), .B(n6501), .Z(n6572) );
  XNOR U6522 ( .A(n6573), .B(n6513), .Z(n6501) );
  XOR U6523 ( .A(n6487), .B(n6485), .Z(n6513) );
  XNOR U6524 ( .A(n6574), .B(n6492), .Z(n6485) );
  XOR U6525 ( .A(p_input[24]), .B(p_input[536]), .Z(n6492) );
  XOR U6526 ( .A(n6482), .B(n6491), .Z(n6574) );
  XOR U6527 ( .A(n6575), .B(n6488), .Z(n6491) );
  XOR U6528 ( .A(p_input[22]), .B(p_input[534]), .Z(n6488) );
  XOR U6529 ( .A(p_input[23]), .B(n6576), .Z(n6575) );
  XOR U6530 ( .A(p_input[18]), .B(p_input[530]), .Z(n6482) );
  XNOR U6531 ( .A(n6497), .B(n6496), .Z(n6487) );
  XOR U6532 ( .A(n6577), .B(n6493), .Z(n6496) );
  XOR U6533 ( .A(p_input[19]), .B(p_input[531]), .Z(n6493) );
  XOR U6534 ( .A(p_input[20]), .B(n6578), .Z(n6577) );
  XOR U6535 ( .A(p_input[21]), .B(p_input[533]), .Z(n6497) );
  XOR U6536 ( .A(n6512), .B(n6579), .Z(n6573) );
  IV U6537 ( .A(n6498), .Z(n6579) );
  XOR U6538 ( .A(p_input[1]), .B(p_input[513]), .Z(n6498) );
  XNOR U6539 ( .A(n6580), .B(n6520), .Z(n6512) );
  XNOR U6540 ( .A(n6508), .B(n6507), .Z(n6520) );
  XNOR U6541 ( .A(n6581), .B(n6504), .Z(n6507) );
  XNOR U6542 ( .A(p_input[26]), .B(p_input[538]), .Z(n6504) );
  XOR U6543 ( .A(p_input[27]), .B(n6582), .Z(n6581) );
  XOR U6544 ( .A(p_input[28]), .B(p_input[540]), .Z(n6508) );
  XOR U6545 ( .A(n6518), .B(n6583), .Z(n6580) );
  IV U6546 ( .A(n6509), .Z(n6583) );
  XOR U6547 ( .A(p_input[17]), .B(p_input[529]), .Z(n6509) );
  XNOR U6548 ( .A(n6584), .B(n6525), .Z(n6518) );
  XNOR U6549 ( .A(p_input[31]), .B(n6585), .Z(n6525) );
  XOR U6550 ( .A(n6515), .B(n6524), .Z(n6584) );
  XOR U6551 ( .A(n6586), .B(n6521), .Z(n6524) );
  XOR U6552 ( .A(p_input[29]), .B(p_input[541]), .Z(n6521) );
  XOR U6553 ( .A(p_input[30]), .B(n6587), .Z(n6586) );
  XOR U6554 ( .A(p_input[25]), .B(p_input[537]), .Z(n6515) );
  XNOR U6555 ( .A(n6537), .B(n6536), .Z(n6502) );
  XNOR U6556 ( .A(n6588), .B(n6544), .Z(n6536) );
  XNOR U6557 ( .A(n6532), .B(n6531), .Z(n6544) );
  XNOR U6558 ( .A(n6589), .B(n6528), .Z(n6531) );
  XNOR U6559 ( .A(p_input[11]), .B(p_input[523]), .Z(n6528) );
  XOR U6560 ( .A(p_input[12]), .B(n6590), .Z(n6589) );
  XOR U6561 ( .A(p_input[13]), .B(p_input[525]), .Z(n6532) );
  XOR U6562 ( .A(n6542), .B(n6591), .Z(n6588) );
  IV U6563 ( .A(n6533), .Z(n6591) );
  XOR U6564 ( .A(p_input[2]), .B(p_input[514]), .Z(n6533) );
  XNOR U6565 ( .A(n6592), .B(n6549), .Z(n6542) );
  XNOR U6566 ( .A(p_input[16]), .B(n6593), .Z(n6549) );
  XOR U6567 ( .A(n6539), .B(n6548), .Z(n6592) );
  XOR U6568 ( .A(n6594), .B(n6545), .Z(n6548) );
  XOR U6569 ( .A(p_input[14]), .B(p_input[526]), .Z(n6545) );
  XOR U6570 ( .A(p_input[15]), .B(n6595), .Z(n6594) );
  XOR U6571 ( .A(p_input[10]), .B(p_input[522]), .Z(n6539) );
  XNOR U6572 ( .A(n6556), .B(n6554), .Z(n6537) );
  XNOR U6573 ( .A(n6596), .B(n6561), .Z(n6554) );
  XOR U6574 ( .A(p_input[521]), .B(p_input[9]), .Z(n6561) );
  XOR U6575 ( .A(n6551), .B(n6560), .Z(n6596) );
  XOR U6576 ( .A(n6597), .B(n6557), .Z(n6560) );
  XOR U6577 ( .A(p_input[519]), .B(p_input[7]), .Z(n6557) );
  XNOR U6578 ( .A(p_input[520]), .B(p_input[8]), .Z(n6597) );
  XOR U6579 ( .A(p_input[3]), .B(p_input[515]), .Z(n6551) );
  XNOR U6580 ( .A(n6566), .B(n6565), .Z(n6556) );
  XOR U6581 ( .A(n6598), .B(n6562), .Z(n6565) );
  XOR U6582 ( .A(p_input[4]), .B(p_input[516]), .Z(n6562) );
  XNOR U6583 ( .A(p_input[517]), .B(p_input[5]), .Z(n6598) );
  XOR U6584 ( .A(p_input[518]), .B(p_input[6]), .Z(n6566) );
  IV U6585 ( .A(n6366), .Z(n6370) );
  XOR U6586 ( .A(n6599), .B(n6600), .Z(n6366) );
  AND U6587 ( .A(n134), .B(n6601), .Z(n6600) );
  XNOR U6588 ( .A(n6602), .B(n6603), .Z(n134) );
  AND U6589 ( .A(n6604), .B(n6605), .Z(n6603) );
  XOR U6590 ( .A(n6381), .B(n6602), .Z(n6605) );
  XNOR U6591 ( .A(n6606), .B(n6602), .Z(n6604) );
  XOR U6592 ( .A(n6607), .B(n6608), .Z(n6602) );
  AND U6593 ( .A(n6609), .B(n6610), .Z(n6608) );
  XOR U6594 ( .A(n6396), .B(n6607), .Z(n6610) );
  XOR U6595 ( .A(n6607), .B(n6397), .Z(n6609) );
  XOR U6596 ( .A(n6611), .B(n6612), .Z(n6607) );
  AND U6597 ( .A(n6613), .B(n6614), .Z(n6612) );
  XOR U6598 ( .A(n6424), .B(n6611), .Z(n6614) );
  XOR U6599 ( .A(n6611), .B(n6425), .Z(n6613) );
  XOR U6600 ( .A(n6615), .B(n6616), .Z(n6611) );
  AND U6601 ( .A(n6617), .B(n6618), .Z(n6616) );
  XOR U6602 ( .A(n6473), .B(n6615), .Z(n6618) );
  XOR U6603 ( .A(n6615), .B(n6474), .Z(n6617) );
  XOR U6604 ( .A(n6619), .B(n6620), .Z(n6615) );
  AND U6605 ( .A(n6621), .B(n6622), .Z(n6620) );
  XOR U6606 ( .A(n6619), .B(n6570), .Z(n6622) );
  XNOR U6607 ( .A(n6623), .B(n6624), .Z(n6309) );
  AND U6608 ( .A(n138), .B(n6625), .Z(n6624) );
  XNOR U6609 ( .A(n6626), .B(n6627), .Z(n138) );
  AND U6610 ( .A(n6628), .B(n6629), .Z(n6627) );
  XOR U6611 ( .A(n6626), .B(n6321), .Z(n6629) );
  XNOR U6612 ( .A(n6626), .B(n6252), .Z(n6628) );
  XOR U6613 ( .A(n6630), .B(n6631), .Z(n6626) );
  AND U6614 ( .A(n6632), .B(n6633), .Z(n6631) );
  XNOR U6615 ( .A(n6331), .B(n6630), .Z(n6633) );
  XOR U6616 ( .A(n6630), .B(n6333), .Z(n6632) );
  XOR U6617 ( .A(n6634), .B(n6635), .Z(n6630) );
  AND U6618 ( .A(n6636), .B(n6637), .Z(n6635) );
  XNOR U6619 ( .A(n6342), .B(n6634), .Z(n6637) );
  XOR U6620 ( .A(n6634), .B(n6344), .Z(n6636) );
  IV U6621 ( .A(n6278), .Z(n6344) );
  XOR U6622 ( .A(n6638), .B(n6639), .Z(n6634) );
  AND U6623 ( .A(n6640), .B(n6641), .Z(n6639) );
  XOR U6624 ( .A(n6638), .B(n6355), .Z(n6640) );
  XOR U6625 ( .A(n6642), .B(n6643), .Z(n6307) );
  AND U6626 ( .A(n142), .B(n6625), .Z(n6643) );
  XNOR U6627 ( .A(n6623), .B(n6642), .Z(n6625) );
  XNOR U6628 ( .A(n6644), .B(n6645), .Z(n142) );
  AND U6629 ( .A(n6646), .B(n6647), .Z(n6645) );
  XNOR U6630 ( .A(n6648), .B(n6644), .Z(n6647) );
  IV U6631 ( .A(n6321), .Z(n6648) );
  XOR U6632 ( .A(n6606), .B(n6649), .Z(n6321) );
  AND U6633 ( .A(n146), .B(n6650), .Z(n6649) );
  XOR U6634 ( .A(n6380), .B(n6377), .Z(n6650) );
  IV U6635 ( .A(n6606), .Z(n6380) );
  XNOR U6636 ( .A(n6252), .B(n6644), .Z(n6646) );
  XOR U6637 ( .A(n6651), .B(n6652), .Z(n6252) );
  AND U6638 ( .A(n162), .B(n6653), .Z(n6652) );
  XOR U6639 ( .A(n6654), .B(n6655), .Z(n6644) );
  AND U6640 ( .A(n6656), .B(n6657), .Z(n6655) );
  XNOR U6641 ( .A(n6654), .B(n6331), .Z(n6657) );
  XOR U6642 ( .A(n6397), .B(n6658), .Z(n6331) );
  AND U6643 ( .A(n146), .B(n6659), .Z(n6658) );
  XOR U6644 ( .A(n6393), .B(n6397), .Z(n6659) );
  XNOR U6645 ( .A(n6265), .B(n6654), .Z(n6656) );
  IV U6646 ( .A(n6333), .Z(n6265) );
  XOR U6647 ( .A(n6660), .B(n6661), .Z(n6333) );
  AND U6648 ( .A(n162), .B(n6662), .Z(n6661) );
  XOR U6649 ( .A(n6663), .B(n6664), .Z(n6654) );
  AND U6650 ( .A(n6665), .B(n6666), .Z(n6664) );
  XNOR U6651 ( .A(n6663), .B(n6342), .Z(n6666) );
  XOR U6652 ( .A(n6425), .B(n6667), .Z(n6342) );
  AND U6653 ( .A(n146), .B(n6668), .Z(n6667) );
  XOR U6654 ( .A(n6421), .B(n6425), .Z(n6668) );
  XNOR U6655 ( .A(n6278), .B(n6663), .Z(n6665) );
  XNOR U6656 ( .A(n6669), .B(n6670), .Z(n6278) );
  AND U6657 ( .A(n162), .B(n6671), .Z(n6670) );
  XOR U6658 ( .A(n6638), .B(n6672), .Z(n6663) );
  AND U6659 ( .A(n6673), .B(n6641), .Z(n6672) );
  XNOR U6660 ( .A(n6353), .B(n6638), .Z(n6641) );
  XOR U6661 ( .A(n6474), .B(n6674), .Z(n6353) );
  AND U6662 ( .A(n146), .B(n6675), .Z(n6674) );
  XOR U6663 ( .A(n6470), .B(n6474), .Z(n6675) );
  XNOR U6664 ( .A(n6291), .B(n6638), .Z(n6673) );
  IV U6665 ( .A(n6355), .Z(n6291) );
  XOR U6666 ( .A(n6676), .B(n6677), .Z(n6355) );
  AND U6667 ( .A(n162), .B(n6678), .Z(n6677) );
  XOR U6668 ( .A(n6679), .B(n6680), .Z(n6638) );
  AND U6669 ( .A(n6681), .B(n6682), .Z(n6680) );
  XNOR U6670 ( .A(n6679), .B(n6364), .Z(n6682) );
  XOR U6671 ( .A(n6571), .B(n6683), .Z(n6364) );
  AND U6672 ( .A(n146), .B(n6684), .Z(n6683) );
  XOR U6673 ( .A(n6567), .B(n6571), .Z(n6684) );
  XNOR U6674 ( .A(n6685), .B(n6679), .Z(n6681) );
  IV U6675 ( .A(n6304), .Z(n6685) );
  XOR U6676 ( .A(n6686), .B(n6687), .Z(n6304) );
  AND U6677 ( .A(n162), .B(n6688), .Z(n6687) );
  AND U6678 ( .A(n6642), .B(n6623), .Z(n6679) );
  XNOR U6679 ( .A(n6689), .B(n6690), .Z(n6623) );
  AND U6680 ( .A(n146), .B(n6601), .Z(n6690) );
  XNOR U6681 ( .A(n6599), .B(n6689), .Z(n6601) );
  XNOR U6682 ( .A(n6691), .B(n6692), .Z(n146) );
  AND U6683 ( .A(n6693), .B(n6694), .Z(n6692) );
  XNOR U6684 ( .A(n6691), .B(n6377), .Z(n6694) );
  IV U6685 ( .A(n6381), .Z(n6377) );
  XOR U6686 ( .A(n6695), .B(n6696), .Z(n6381) );
  AND U6687 ( .A(n150), .B(n6697), .Z(n6696) );
  XOR U6688 ( .A(n6698), .B(n6695), .Z(n6697) );
  XNOR U6689 ( .A(n6691), .B(n6606), .Z(n6693) );
  XOR U6690 ( .A(n6699), .B(n6700), .Z(n6606) );
  AND U6691 ( .A(n158), .B(n6653), .Z(n6700) );
  XOR U6692 ( .A(n6651), .B(n6699), .Z(n6653) );
  XOR U6693 ( .A(n6701), .B(n6702), .Z(n6691) );
  AND U6694 ( .A(n6703), .B(n6704), .Z(n6702) );
  XNOR U6695 ( .A(n6701), .B(n6393), .Z(n6704) );
  IV U6696 ( .A(n6396), .Z(n6393) );
  XOR U6697 ( .A(n6705), .B(n6706), .Z(n6396) );
  AND U6698 ( .A(n150), .B(n6707), .Z(n6706) );
  XOR U6699 ( .A(n6708), .B(n6705), .Z(n6707) );
  XOR U6700 ( .A(n6397), .B(n6701), .Z(n6703) );
  XOR U6701 ( .A(n6709), .B(n6710), .Z(n6397) );
  AND U6702 ( .A(n158), .B(n6662), .Z(n6710) );
  XOR U6703 ( .A(n6709), .B(n6660), .Z(n6662) );
  XOR U6704 ( .A(n6711), .B(n6712), .Z(n6701) );
  AND U6705 ( .A(n6713), .B(n6714), .Z(n6712) );
  XNOR U6706 ( .A(n6711), .B(n6421), .Z(n6714) );
  IV U6707 ( .A(n6424), .Z(n6421) );
  XOR U6708 ( .A(n6715), .B(n6716), .Z(n6424) );
  AND U6709 ( .A(n150), .B(n6717), .Z(n6716) );
  XNOR U6710 ( .A(n6718), .B(n6715), .Z(n6717) );
  XOR U6711 ( .A(n6425), .B(n6711), .Z(n6713) );
  XOR U6712 ( .A(n6719), .B(n6720), .Z(n6425) );
  AND U6713 ( .A(n158), .B(n6671), .Z(n6720) );
  XOR U6714 ( .A(n6719), .B(n6669), .Z(n6671) );
  XOR U6715 ( .A(n6721), .B(n6722), .Z(n6711) );
  AND U6716 ( .A(n6723), .B(n6724), .Z(n6722) );
  XNOR U6717 ( .A(n6721), .B(n6470), .Z(n6724) );
  IV U6718 ( .A(n6473), .Z(n6470) );
  XOR U6719 ( .A(n6725), .B(n6726), .Z(n6473) );
  AND U6720 ( .A(n150), .B(n6727), .Z(n6726) );
  XOR U6721 ( .A(n6728), .B(n6725), .Z(n6727) );
  XOR U6722 ( .A(n6474), .B(n6721), .Z(n6723) );
  XOR U6723 ( .A(n6729), .B(n6730), .Z(n6474) );
  AND U6724 ( .A(n158), .B(n6678), .Z(n6730) );
  XOR U6725 ( .A(n6729), .B(n6676), .Z(n6678) );
  XOR U6726 ( .A(n6619), .B(n6731), .Z(n6721) );
  AND U6727 ( .A(n6621), .B(n6732), .Z(n6731) );
  XNOR U6728 ( .A(n6619), .B(n6567), .Z(n6732) );
  IV U6729 ( .A(n6570), .Z(n6567) );
  XOR U6730 ( .A(n6733), .B(n6734), .Z(n6570) );
  AND U6731 ( .A(n150), .B(n6735), .Z(n6734) );
  XNOR U6732 ( .A(n6736), .B(n6733), .Z(n6735) );
  XOR U6733 ( .A(n6571), .B(n6619), .Z(n6621) );
  XOR U6734 ( .A(n6737), .B(n6738), .Z(n6571) );
  AND U6735 ( .A(n158), .B(n6688), .Z(n6738) );
  XOR U6736 ( .A(n6737), .B(n6686), .Z(n6688) );
  AND U6737 ( .A(n6689), .B(n6599), .Z(n6619) );
  XNOR U6738 ( .A(n6739), .B(n6740), .Z(n6599) );
  AND U6739 ( .A(n150), .B(n6741), .Z(n6740) );
  XNOR U6740 ( .A(n6742), .B(n6739), .Z(n6741) );
  XNOR U6741 ( .A(n6743), .B(n6744), .Z(n150) );
  AND U6742 ( .A(n6745), .B(n6746), .Z(n6744) );
  XOR U6743 ( .A(n6698), .B(n6743), .Z(n6746) );
  AND U6744 ( .A(n6747), .B(n6748), .Z(n6698) );
  XNOR U6745 ( .A(n6695), .B(n6743), .Z(n6745) );
  XNOR U6746 ( .A(n6749), .B(n6750), .Z(n6695) );
  AND U6747 ( .A(n154), .B(n6751), .Z(n6750) );
  XNOR U6748 ( .A(n6752), .B(n6753), .Z(n6751) );
  XOR U6749 ( .A(n6754), .B(n6755), .Z(n6743) );
  AND U6750 ( .A(n6756), .B(n6757), .Z(n6755) );
  XNOR U6751 ( .A(n6754), .B(n6747), .Z(n6757) );
  IV U6752 ( .A(n6708), .Z(n6747) );
  XOR U6753 ( .A(n6758), .B(n6759), .Z(n6708) );
  XOR U6754 ( .A(n6760), .B(n6748), .Z(n6759) );
  AND U6755 ( .A(n6718), .B(n6761), .Z(n6748) );
  AND U6756 ( .A(n6762), .B(n6763), .Z(n6760) );
  XOR U6757 ( .A(n6764), .B(n6758), .Z(n6762) );
  XNOR U6758 ( .A(n6705), .B(n6754), .Z(n6756) );
  XNOR U6759 ( .A(n6765), .B(n6766), .Z(n6705) );
  AND U6760 ( .A(n154), .B(n6767), .Z(n6766) );
  XNOR U6761 ( .A(n6768), .B(n6769), .Z(n6767) );
  XOR U6762 ( .A(n6770), .B(n6771), .Z(n6754) );
  AND U6763 ( .A(n6772), .B(n6773), .Z(n6771) );
  XNOR U6764 ( .A(n6770), .B(n6718), .Z(n6773) );
  XOR U6765 ( .A(n6774), .B(n6763), .Z(n6718) );
  XNOR U6766 ( .A(n6775), .B(n6758), .Z(n6763) );
  XOR U6767 ( .A(n6776), .B(n6777), .Z(n6758) );
  AND U6768 ( .A(n6778), .B(n6779), .Z(n6777) );
  XOR U6769 ( .A(n6780), .B(n6776), .Z(n6778) );
  XNOR U6770 ( .A(n6781), .B(n6782), .Z(n6775) );
  AND U6771 ( .A(n6783), .B(n6784), .Z(n6782) );
  XOR U6772 ( .A(n6781), .B(n6785), .Z(n6783) );
  XNOR U6773 ( .A(n6764), .B(n6761), .Z(n6774) );
  AND U6774 ( .A(n6786), .B(n6787), .Z(n6761) );
  XOR U6775 ( .A(n6788), .B(n6789), .Z(n6764) );
  AND U6776 ( .A(n6790), .B(n6791), .Z(n6789) );
  XOR U6777 ( .A(n6788), .B(n6792), .Z(n6790) );
  XNOR U6778 ( .A(n6715), .B(n6770), .Z(n6772) );
  XNOR U6779 ( .A(n6793), .B(n6794), .Z(n6715) );
  AND U6780 ( .A(n154), .B(n6795), .Z(n6794) );
  XNOR U6781 ( .A(n6796), .B(n6797), .Z(n6795) );
  XOR U6782 ( .A(n6798), .B(n6799), .Z(n6770) );
  AND U6783 ( .A(n6800), .B(n6801), .Z(n6799) );
  XNOR U6784 ( .A(n6798), .B(n6786), .Z(n6801) );
  IV U6785 ( .A(n6728), .Z(n6786) );
  XNOR U6786 ( .A(n6802), .B(n6779), .Z(n6728) );
  XNOR U6787 ( .A(n6803), .B(n6785), .Z(n6779) );
  XOR U6788 ( .A(n6804), .B(n6805), .Z(n6785) );
  AND U6789 ( .A(n6806), .B(n6807), .Z(n6805) );
  XOR U6790 ( .A(n6804), .B(n6808), .Z(n6806) );
  XNOR U6791 ( .A(n6784), .B(n6776), .Z(n6803) );
  XOR U6792 ( .A(n6809), .B(n6810), .Z(n6776) );
  AND U6793 ( .A(n6811), .B(n6812), .Z(n6810) );
  XNOR U6794 ( .A(n6813), .B(n6809), .Z(n6811) );
  XNOR U6795 ( .A(n6814), .B(n6781), .Z(n6784) );
  XOR U6796 ( .A(n6815), .B(n6816), .Z(n6781) );
  AND U6797 ( .A(n6817), .B(n6818), .Z(n6816) );
  XOR U6798 ( .A(n6815), .B(n6819), .Z(n6817) );
  XNOR U6799 ( .A(n6820), .B(n6821), .Z(n6814) );
  AND U6800 ( .A(n6822), .B(n6823), .Z(n6821) );
  XNOR U6801 ( .A(n6820), .B(n6824), .Z(n6822) );
  XNOR U6802 ( .A(n6780), .B(n6787), .Z(n6802) );
  AND U6803 ( .A(n6736), .B(n6825), .Z(n6787) );
  XOR U6804 ( .A(n6792), .B(n6791), .Z(n6780) );
  XNOR U6805 ( .A(n6826), .B(n6788), .Z(n6791) );
  XOR U6806 ( .A(n6827), .B(n6828), .Z(n6788) );
  AND U6807 ( .A(n6829), .B(n6830), .Z(n6828) );
  XOR U6808 ( .A(n6827), .B(n6831), .Z(n6829) );
  XNOR U6809 ( .A(n6832), .B(n6833), .Z(n6826) );
  AND U6810 ( .A(n6834), .B(n6835), .Z(n6833) );
  XOR U6811 ( .A(n6832), .B(n6836), .Z(n6834) );
  XOR U6812 ( .A(n6837), .B(n6838), .Z(n6792) );
  AND U6813 ( .A(n6839), .B(n6840), .Z(n6838) );
  XOR U6814 ( .A(n6837), .B(n6841), .Z(n6839) );
  XNOR U6815 ( .A(n6725), .B(n6798), .Z(n6800) );
  XNOR U6816 ( .A(n6842), .B(n6843), .Z(n6725) );
  AND U6817 ( .A(n154), .B(n6844), .Z(n6843) );
  XNOR U6818 ( .A(n6845), .B(n6846), .Z(n6844) );
  XOR U6819 ( .A(n6847), .B(n6848), .Z(n6798) );
  AND U6820 ( .A(n6849), .B(n6850), .Z(n6848) );
  XNOR U6821 ( .A(n6847), .B(n6736), .Z(n6850) );
  XOR U6822 ( .A(n6851), .B(n6812), .Z(n6736) );
  XNOR U6823 ( .A(n6852), .B(n6819), .Z(n6812) );
  XOR U6824 ( .A(n6808), .B(n6807), .Z(n6819) );
  XNOR U6825 ( .A(n6853), .B(n6804), .Z(n6807) );
  XOR U6826 ( .A(n6854), .B(n6855), .Z(n6804) );
  AND U6827 ( .A(n6856), .B(n6857), .Z(n6855) );
  XNOR U6828 ( .A(n6858), .B(n6859), .Z(n6856) );
  IV U6829 ( .A(n6854), .Z(n6858) );
  XNOR U6830 ( .A(n6860), .B(n6861), .Z(n6853) );
  NOR U6831 ( .A(n6862), .B(n6863), .Z(n6861) );
  XNOR U6832 ( .A(n6860), .B(n6864), .Z(n6862) );
  XOR U6833 ( .A(n6865), .B(n6866), .Z(n6808) );
  NOR U6834 ( .A(n6867), .B(n6868), .Z(n6866) );
  XNOR U6835 ( .A(n6865), .B(n6869), .Z(n6867) );
  XNOR U6836 ( .A(n6818), .B(n6809), .Z(n6852) );
  XOR U6837 ( .A(n6870), .B(n6871), .Z(n6809) );
  NOR U6838 ( .A(n6872), .B(n6873), .Z(n6871) );
  XOR U6839 ( .A(n6874), .B(n6875), .Z(n6872) );
  XOR U6840 ( .A(n6876), .B(n6824), .Z(n6818) );
  XNOR U6841 ( .A(n6877), .B(n6878), .Z(n6824) );
  NOR U6842 ( .A(n6879), .B(n6880), .Z(n6878) );
  XNOR U6843 ( .A(n6877), .B(n6881), .Z(n6879) );
  XNOR U6844 ( .A(n6823), .B(n6815), .Z(n6876) );
  XOR U6845 ( .A(n6882), .B(n6883), .Z(n6815) );
  AND U6846 ( .A(n6884), .B(n6885), .Z(n6883) );
  XOR U6847 ( .A(n6882), .B(n6886), .Z(n6884) );
  XNOR U6848 ( .A(n6887), .B(n6820), .Z(n6823) );
  XOR U6849 ( .A(n6888), .B(n6889), .Z(n6820) );
  AND U6850 ( .A(n6890), .B(n6891), .Z(n6889) );
  XOR U6851 ( .A(n6888), .B(n6892), .Z(n6890) );
  XNOR U6852 ( .A(n6893), .B(n6894), .Z(n6887) );
  NOR U6853 ( .A(n6895), .B(n6896), .Z(n6894) );
  XOR U6854 ( .A(n6893), .B(n6897), .Z(n6895) );
  XOR U6855 ( .A(n6813), .B(n6825), .Z(n6851) );
  NOR U6856 ( .A(n6742), .B(n6898), .Z(n6825) );
  XNOR U6857 ( .A(n6831), .B(n6830), .Z(n6813) );
  XNOR U6858 ( .A(n6899), .B(n6836), .Z(n6830) );
  XNOR U6859 ( .A(n6900), .B(n6901), .Z(n6836) );
  NOR U6860 ( .A(n6902), .B(n6903), .Z(n6901) );
  XOR U6861 ( .A(n6900), .B(n6904), .Z(n6902) );
  XNOR U6862 ( .A(n6835), .B(n6827), .Z(n6899) );
  XOR U6863 ( .A(n6905), .B(n6906), .Z(n6827) );
  AND U6864 ( .A(n6907), .B(n6908), .Z(n6906) );
  XOR U6865 ( .A(n6905), .B(n6909), .Z(n6907) );
  XNOR U6866 ( .A(n6910), .B(n6832), .Z(n6835) );
  XOR U6867 ( .A(n6911), .B(n6912), .Z(n6832) );
  AND U6868 ( .A(n6913), .B(n6914), .Z(n6912) );
  XNOR U6869 ( .A(n6915), .B(n6916), .Z(n6913) );
  IV U6870 ( .A(n6911), .Z(n6915) );
  XNOR U6871 ( .A(n6917), .B(n6918), .Z(n6910) );
  NOR U6872 ( .A(n6919), .B(n6920), .Z(n6918) );
  XNOR U6873 ( .A(n6917), .B(n6921), .Z(n6919) );
  XOR U6874 ( .A(n6841), .B(n6840), .Z(n6831) );
  XNOR U6875 ( .A(n6922), .B(n6837), .Z(n6840) );
  XOR U6876 ( .A(n6923), .B(n6924), .Z(n6837) );
  AND U6877 ( .A(n6925), .B(n6926), .Z(n6924) );
  XNOR U6878 ( .A(n6927), .B(n6928), .Z(n6925) );
  IV U6879 ( .A(n6923), .Z(n6927) );
  XNOR U6880 ( .A(n6929), .B(n6930), .Z(n6922) );
  NOR U6881 ( .A(n6931), .B(n6932), .Z(n6930) );
  XNOR U6882 ( .A(n6929), .B(n6933), .Z(n6931) );
  XOR U6883 ( .A(n6934), .B(n6935), .Z(n6841) );
  NOR U6884 ( .A(n6936), .B(n6937), .Z(n6935) );
  XNOR U6885 ( .A(n6934), .B(n6938), .Z(n6936) );
  XNOR U6886 ( .A(n6733), .B(n6847), .Z(n6849) );
  XNOR U6887 ( .A(n6939), .B(n6940), .Z(n6733) );
  AND U6888 ( .A(n154), .B(n6941), .Z(n6940) );
  XNOR U6889 ( .A(n6942), .B(n6943), .Z(n6941) );
  AND U6890 ( .A(n6739), .B(n6742), .Z(n6847) );
  XOR U6891 ( .A(n6944), .B(n6898), .Z(n6742) );
  XNOR U6892 ( .A(p_input[32]), .B(p_input[512]), .Z(n6898) );
  XOR U6893 ( .A(n6875), .B(n6873), .Z(n6944) );
  XOR U6894 ( .A(n6945), .B(n6886), .Z(n6873) );
  XOR U6895 ( .A(n6859), .B(n6857), .Z(n6886) );
  XNOR U6896 ( .A(n6946), .B(n6864), .Z(n6857) );
  XOR U6897 ( .A(p_input[536]), .B(p_input[56]), .Z(n6864) );
  XOR U6898 ( .A(n6854), .B(n6863), .Z(n6946) );
  XOR U6899 ( .A(n6947), .B(n6860), .Z(n6863) );
  XOR U6900 ( .A(p_input[534]), .B(p_input[54]), .Z(n6860) );
  XNOR U6901 ( .A(p_input[535]), .B(p_input[55]), .Z(n6947) );
  XOR U6902 ( .A(p_input[50]), .B(p_input[530]), .Z(n6854) );
  XNOR U6903 ( .A(n6869), .B(n6868), .Z(n6859) );
  XOR U6904 ( .A(n6948), .B(n6865), .Z(n6868) );
  XOR U6905 ( .A(p_input[51]), .B(p_input[531]), .Z(n6865) );
  XOR U6906 ( .A(p_input[52]), .B(n6578), .Z(n6948) );
  XOR U6907 ( .A(p_input[533]), .B(p_input[53]), .Z(n6869) );
  XOR U6908 ( .A(n6885), .B(n6874), .Z(n6945) );
  IV U6909 ( .A(n6870), .Z(n6874) );
  XOR U6910 ( .A(p_input[33]), .B(p_input[513]), .Z(n6870) );
  XNOR U6911 ( .A(n6949), .B(n6892), .Z(n6885) );
  XNOR U6912 ( .A(n6881), .B(n6880), .Z(n6892) );
  XOR U6913 ( .A(n6950), .B(n6877), .Z(n6880) );
  XNOR U6914 ( .A(n6951), .B(p_input[58]), .Z(n6877) );
  XNOR U6915 ( .A(p_input[539]), .B(p_input[59]), .Z(n6950) );
  XOR U6916 ( .A(p_input[540]), .B(p_input[60]), .Z(n6881) );
  XOR U6917 ( .A(n6891), .B(n6952), .Z(n6949) );
  IV U6918 ( .A(n6882), .Z(n6952) );
  XOR U6919 ( .A(p_input[49]), .B(p_input[529]), .Z(n6882) );
  XOR U6920 ( .A(n6953), .B(n6897), .Z(n6891) );
  XNOR U6921 ( .A(p_input[543]), .B(p_input[63]), .Z(n6897) );
  XOR U6922 ( .A(n6888), .B(n6896), .Z(n6953) );
  XOR U6923 ( .A(n6954), .B(n6893), .Z(n6896) );
  XOR U6924 ( .A(p_input[541]), .B(p_input[61]), .Z(n6893) );
  XNOR U6925 ( .A(p_input[542]), .B(p_input[62]), .Z(n6954) );
  XNOR U6926 ( .A(n6955), .B(p_input[57]), .Z(n6888) );
  XOR U6927 ( .A(n6909), .B(n6908), .Z(n6875) );
  XNOR U6928 ( .A(n6956), .B(n6916), .Z(n6908) );
  XNOR U6929 ( .A(n6904), .B(n6903), .Z(n6916) );
  XNOR U6930 ( .A(n6957), .B(n6900), .Z(n6903) );
  XNOR U6931 ( .A(p_input[43]), .B(p_input[523]), .Z(n6900) );
  XOR U6932 ( .A(p_input[44]), .B(n6590), .Z(n6957) );
  XOR U6933 ( .A(p_input[45]), .B(p_input[525]), .Z(n6904) );
  XOR U6934 ( .A(n6914), .B(n6958), .Z(n6956) );
  IV U6935 ( .A(n6905), .Z(n6958) );
  XOR U6936 ( .A(p_input[34]), .B(p_input[514]), .Z(n6905) );
  XNOR U6937 ( .A(n6959), .B(n6921), .Z(n6914) );
  XNOR U6938 ( .A(p_input[48]), .B(n6593), .Z(n6921) );
  XOR U6939 ( .A(n6911), .B(n6920), .Z(n6959) );
  XOR U6940 ( .A(n6960), .B(n6917), .Z(n6920) );
  XOR U6941 ( .A(p_input[46]), .B(p_input[526]), .Z(n6917) );
  XOR U6942 ( .A(p_input[47]), .B(n6595), .Z(n6960) );
  XOR U6943 ( .A(p_input[42]), .B(p_input[522]), .Z(n6911) );
  XOR U6944 ( .A(n6928), .B(n6926), .Z(n6909) );
  XNOR U6945 ( .A(n6961), .B(n6933), .Z(n6926) );
  XOR U6946 ( .A(p_input[41]), .B(p_input[521]), .Z(n6933) );
  XOR U6947 ( .A(n6923), .B(n6932), .Z(n6961) );
  XOR U6948 ( .A(n6962), .B(n6929), .Z(n6932) );
  XOR U6949 ( .A(p_input[39]), .B(p_input[519]), .Z(n6929) );
  XOR U6950 ( .A(p_input[40]), .B(n6963), .Z(n6962) );
  XOR U6951 ( .A(p_input[35]), .B(p_input[515]), .Z(n6923) );
  XNOR U6952 ( .A(n6938), .B(n6937), .Z(n6928) );
  XOR U6953 ( .A(n6964), .B(n6934), .Z(n6937) );
  XOR U6954 ( .A(p_input[36]), .B(p_input[516]), .Z(n6934) );
  XOR U6955 ( .A(p_input[37]), .B(n6965), .Z(n6964) );
  XOR U6956 ( .A(p_input[38]), .B(p_input[518]), .Z(n6938) );
  XNOR U6957 ( .A(n6966), .B(n6967), .Z(n6739) );
  AND U6958 ( .A(n154), .B(n6968), .Z(n6967) );
  XNOR U6959 ( .A(n6969), .B(n6970), .Z(n154) );
  AND U6960 ( .A(n6971), .B(n6972), .Z(n6970) );
  XOR U6961 ( .A(n6753), .B(n6969), .Z(n6972) );
  XNOR U6962 ( .A(n6973), .B(n6969), .Z(n6971) );
  XOR U6963 ( .A(n6974), .B(n6975), .Z(n6969) );
  AND U6964 ( .A(n6976), .B(n6977), .Z(n6975) );
  XOR U6965 ( .A(n6768), .B(n6974), .Z(n6977) );
  XOR U6966 ( .A(n6974), .B(n6769), .Z(n6976) );
  XOR U6967 ( .A(n6978), .B(n6979), .Z(n6974) );
  AND U6968 ( .A(n6980), .B(n6981), .Z(n6979) );
  XOR U6969 ( .A(n6796), .B(n6978), .Z(n6981) );
  XOR U6970 ( .A(n6978), .B(n6797), .Z(n6980) );
  XOR U6971 ( .A(n6982), .B(n6983), .Z(n6978) );
  AND U6972 ( .A(n6984), .B(n6985), .Z(n6983) );
  XOR U6973 ( .A(n6845), .B(n6982), .Z(n6985) );
  XOR U6974 ( .A(n6982), .B(n6846), .Z(n6984) );
  XOR U6975 ( .A(n6986), .B(n6987), .Z(n6982) );
  AND U6976 ( .A(n6988), .B(n6989), .Z(n6987) );
  XOR U6977 ( .A(n6986), .B(n6942), .Z(n6989) );
  XNOR U6978 ( .A(n6990), .B(n6991), .Z(n6689) );
  AND U6979 ( .A(n158), .B(n6992), .Z(n6991) );
  XNOR U6980 ( .A(n6993), .B(n6994), .Z(n158) );
  AND U6981 ( .A(n6995), .B(n6996), .Z(n6994) );
  XOR U6982 ( .A(n6993), .B(n6699), .Z(n6996) );
  XNOR U6983 ( .A(n6993), .B(n6651), .Z(n6995) );
  XOR U6984 ( .A(n6997), .B(n6998), .Z(n6993) );
  AND U6985 ( .A(n6999), .B(n7000), .Z(n6998) );
  XNOR U6986 ( .A(n6709), .B(n6997), .Z(n7000) );
  XOR U6987 ( .A(n6997), .B(n6660), .Z(n6999) );
  XOR U6988 ( .A(n7001), .B(n7002), .Z(n6997) );
  AND U6989 ( .A(n7003), .B(n7004), .Z(n7002) );
  XNOR U6990 ( .A(n6719), .B(n7001), .Z(n7004) );
  XOR U6991 ( .A(n7001), .B(n6669), .Z(n7003) );
  XOR U6992 ( .A(n7005), .B(n7006), .Z(n7001) );
  AND U6993 ( .A(n7007), .B(n7008), .Z(n7006) );
  XOR U6994 ( .A(n7005), .B(n6676), .Z(n7007) );
  XOR U6995 ( .A(n7009), .B(n7010), .Z(n6642) );
  AND U6996 ( .A(n162), .B(n6992), .Z(n7010) );
  XNOR U6997 ( .A(n6990), .B(n7009), .Z(n6992) );
  XNOR U6998 ( .A(n7011), .B(n7012), .Z(n162) );
  AND U6999 ( .A(n7013), .B(n7014), .Z(n7012) );
  XNOR U7000 ( .A(n7015), .B(n7011), .Z(n7014) );
  IV U7001 ( .A(n6699), .Z(n7015) );
  XOR U7002 ( .A(n6973), .B(n7016), .Z(n6699) );
  AND U7003 ( .A(n165), .B(n7017), .Z(n7016) );
  XOR U7004 ( .A(n6752), .B(n6749), .Z(n7017) );
  IV U7005 ( .A(n6973), .Z(n6752) );
  XNOR U7006 ( .A(n6651), .B(n7011), .Z(n7013) );
  XOR U7007 ( .A(n7018), .B(n7019), .Z(n6651) );
  AND U7008 ( .A(n181), .B(n7020), .Z(n7019) );
  XOR U7009 ( .A(n7021), .B(n7022), .Z(n7011) );
  AND U7010 ( .A(n7023), .B(n7024), .Z(n7022) );
  XNOR U7011 ( .A(n7021), .B(n6709), .Z(n7024) );
  XOR U7012 ( .A(n6769), .B(n7025), .Z(n6709) );
  AND U7013 ( .A(n165), .B(n7026), .Z(n7025) );
  XOR U7014 ( .A(n6765), .B(n6769), .Z(n7026) );
  XNOR U7015 ( .A(n7027), .B(n7021), .Z(n7023) );
  IV U7016 ( .A(n6660), .Z(n7027) );
  XOR U7017 ( .A(n7028), .B(n7029), .Z(n6660) );
  AND U7018 ( .A(n181), .B(n7030), .Z(n7029) );
  XOR U7019 ( .A(n7031), .B(n7032), .Z(n7021) );
  AND U7020 ( .A(n7033), .B(n7034), .Z(n7032) );
  XNOR U7021 ( .A(n7031), .B(n6719), .Z(n7034) );
  XOR U7022 ( .A(n6797), .B(n7035), .Z(n6719) );
  AND U7023 ( .A(n165), .B(n7036), .Z(n7035) );
  XOR U7024 ( .A(n6793), .B(n6797), .Z(n7036) );
  XOR U7025 ( .A(n6669), .B(n7031), .Z(n7033) );
  XOR U7026 ( .A(n7037), .B(n7038), .Z(n6669) );
  AND U7027 ( .A(n181), .B(n7039), .Z(n7038) );
  XOR U7028 ( .A(n7005), .B(n7040), .Z(n7031) );
  AND U7029 ( .A(n7041), .B(n7008), .Z(n7040) );
  XNOR U7030 ( .A(n6729), .B(n7005), .Z(n7008) );
  XOR U7031 ( .A(n6846), .B(n7042), .Z(n6729) );
  AND U7032 ( .A(n165), .B(n7043), .Z(n7042) );
  XOR U7033 ( .A(n6842), .B(n6846), .Z(n7043) );
  XNOR U7034 ( .A(n7044), .B(n7005), .Z(n7041) );
  IV U7035 ( .A(n6676), .Z(n7044) );
  XOR U7036 ( .A(n7045), .B(n7046), .Z(n6676) );
  AND U7037 ( .A(n181), .B(n7047), .Z(n7046) );
  XOR U7038 ( .A(n7048), .B(n7049), .Z(n7005) );
  AND U7039 ( .A(n7050), .B(n7051), .Z(n7049) );
  XNOR U7040 ( .A(n7048), .B(n6737), .Z(n7051) );
  XOR U7041 ( .A(n6943), .B(n7052), .Z(n6737) );
  AND U7042 ( .A(n165), .B(n7053), .Z(n7052) );
  XOR U7043 ( .A(n6939), .B(n6943), .Z(n7053) );
  XNOR U7044 ( .A(n7054), .B(n7048), .Z(n7050) );
  IV U7045 ( .A(n6686), .Z(n7054) );
  XOR U7046 ( .A(n7055), .B(n7056), .Z(n6686) );
  AND U7047 ( .A(n181), .B(n7057), .Z(n7056) );
  AND U7048 ( .A(n7009), .B(n6990), .Z(n7048) );
  XNOR U7049 ( .A(n7058), .B(n7059), .Z(n6990) );
  AND U7050 ( .A(n165), .B(n6968), .Z(n7059) );
  XNOR U7051 ( .A(n6966), .B(n7058), .Z(n6968) );
  XNOR U7052 ( .A(n7060), .B(n7061), .Z(n165) );
  AND U7053 ( .A(n7062), .B(n7063), .Z(n7061) );
  XNOR U7054 ( .A(n7060), .B(n6749), .Z(n7063) );
  IV U7055 ( .A(n6753), .Z(n6749) );
  XOR U7056 ( .A(n7064), .B(n7065), .Z(n6753) );
  AND U7057 ( .A(n169), .B(n7066), .Z(n7065) );
  XOR U7058 ( .A(n7067), .B(n7064), .Z(n7066) );
  XNOR U7059 ( .A(n7060), .B(n6973), .Z(n7062) );
  XOR U7060 ( .A(n7068), .B(n7069), .Z(n6973) );
  AND U7061 ( .A(n177), .B(n7020), .Z(n7069) );
  XOR U7062 ( .A(n7018), .B(n7068), .Z(n7020) );
  XOR U7063 ( .A(n7070), .B(n7071), .Z(n7060) );
  AND U7064 ( .A(n7072), .B(n7073), .Z(n7071) );
  XNOR U7065 ( .A(n7070), .B(n6765), .Z(n7073) );
  IV U7066 ( .A(n6768), .Z(n6765) );
  XOR U7067 ( .A(n7074), .B(n7075), .Z(n6768) );
  AND U7068 ( .A(n169), .B(n7076), .Z(n7075) );
  XOR U7069 ( .A(n7077), .B(n7074), .Z(n7076) );
  XOR U7070 ( .A(n6769), .B(n7070), .Z(n7072) );
  XOR U7071 ( .A(n7078), .B(n7079), .Z(n6769) );
  AND U7072 ( .A(n177), .B(n7030), .Z(n7079) );
  XOR U7073 ( .A(n7078), .B(n7028), .Z(n7030) );
  XOR U7074 ( .A(n7080), .B(n7081), .Z(n7070) );
  AND U7075 ( .A(n7082), .B(n7083), .Z(n7081) );
  XNOR U7076 ( .A(n7080), .B(n6793), .Z(n7083) );
  IV U7077 ( .A(n6796), .Z(n6793) );
  XOR U7078 ( .A(n7084), .B(n7085), .Z(n6796) );
  AND U7079 ( .A(n169), .B(n7086), .Z(n7085) );
  XNOR U7080 ( .A(n7087), .B(n7084), .Z(n7086) );
  XOR U7081 ( .A(n6797), .B(n7080), .Z(n7082) );
  XOR U7082 ( .A(n7088), .B(n7089), .Z(n6797) );
  AND U7083 ( .A(n177), .B(n7039), .Z(n7089) );
  XOR U7084 ( .A(n7088), .B(n7037), .Z(n7039) );
  XOR U7085 ( .A(n7090), .B(n7091), .Z(n7080) );
  AND U7086 ( .A(n7092), .B(n7093), .Z(n7091) );
  XNOR U7087 ( .A(n7090), .B(n6842), .Z(n7093) );
  IV U7088 ( .A(n6845), .Z(n6842) );
  XOR U7089 ( .A(n7094), .B(n7095), .Z(n6845) );
  AND U7090 ( .A(n169), .B(n7096), .Z(n7095) );
  XOR U7091 ( .A(n7097), .B(n7094), .Z(n7096) );
  XOR U7092 ( .A(n6846), .B(n7090), .Z(n7092) );
  XOR U7093 ( .A(n7098), .B(n7099), .Z(n6846) );
  AND U7094 ( .A(n177), .B(n7047), .Z(n7099) );
  XOR U7095 ( .A(n7098), .B(n7045), .Z(n7047) );
  XOR U7096 ( .A(n6986), .B(n7100), .Z(n7090) );
  AND U7097 ( .A(n6988), .B(n7101), .Z(n7100) );
  XNOR U7098 ( .A(n6986), .B(n6939), .Z(n7101) );
  IV U7099 ( .A(n6942), .Z(n6939) );
  XOR U7100 ( .A(n7102), .B(n7103), .Z(n6942) );
  AND U7101 ( .A(n169), .B(n7104), .Z(n7103) );
  XNOR U7102 ( .A(n7105), .B(n7102), .Z(n7104) );
  XOR U7103 ( .A(n6943), .B(n6986), .Z(n6988) );
  XOR U7104 ( .A(n7106), .B(n7107), .Z(n6943) );
  AND U7105 ( .A(n177), .B(n7057), .Z(n7107) );
  XOR U7106 ( .A(n7106), .B(n7055), .Z(n7057) );
  AND U7107 ( .A(n7058), .B(n6966), .Z(n6986) );
  XNOR U7108 ( .A(n7108), .B(n7109), .Z(n6966) );
  AND U7109 ( .A(n169), .B(n7110), .Z(n7109) );
  XNOR U7110 ( .A(n7111), .B(n7108), .Z(n7110) );
  XNOR U7111 ( .A(n7112), .B(n7113), .Z(n169) );
  AND U7112 ( .A(n7114), .B(n7115), .Z(n7113) );
  XOR U7113 ( .A(n7067), .B(n7112), .Z(n7115) );
  AND U7114 ( .A(n7116), .B(n7117), .Z(n7067) );
  XNOR U7115 ( .A(n7064), .B(n7112), .Z(n7114) );
  XNOR U7116 ( .A(n7118), .B(n7119), .Z(n7064) );
  AND U7117 ( .A(n173), .B(n7120), .Z(n7119) );
  XNOR U7118 ( .A(n7121), .B(n7122), .Z(n7120) );
  XOR U7119 ( .A(n7123), .B(n7124), .Z(n7112) );
  AND U7120 ( .A(n7125), .B(n7126), .Z(n7124) );
  XNOR U7121 ( .A(n7123), .B(n7116), .Z(n7126) );
  IV U7122 ( .A(n7077), .Z(n7116) );
  XOR U7123 ( .A(n7127), .B(n7128), .Z(n7077) );
  XOR U7124 ( .A(n7129), .B(n7117), .Z(n7128) );
  AND U7125 ( .A(n7087), .B(n7130), .Z(n7117) );
  AND U7126 ( .A(n7131), .B(n7132), .Z(n7129) );
  XOR U7127 ( .A(n7133), .B(n7127), .Z(n7131) );
  XNOR U7128 ( .A(n7074), .B(n7123), .Z(n7125) );
  XNOR U7129 ( .A(n7134), .B(n7135), .Z(n7074) );
  AND U7130 ( .A(n173), .B(n7136), .Z(n7135) );
  XNOR U7131 ( .A(n7137), .B(n7138), .Z(n7136) );
  XOR U7132 ( .A(n7139), .B(n7140), .Z(n7123) );
  AND U7133 ( .A(n7141), .B(n7142), .Z(n7140) );
  XNOR U7134 ( .A(n7139), .B(n7087), .Z(n7142) );
  XOR U7135 ( .A(n7143), .B(n7132), .Z(n7087) );
  XNOR U7136 ( .A(n7144), .B(n7127), .Z(n7132) );
  XOR U7137 ( .A(n7145), .B(n7146), .Z(n7127) );
  AND U7138 ( .A(n7147), .B(n7148), .Z(n7146) );
  XOR U7139 ( .A(n7149), .B(n7145), .Z(n7147) );
  XNOR U7140 ( .A(n7150), .B(n7151), .Z(n7144) );
  AND U7141 ( .A(n7152), .B(n7153), .Z(n7151) );
  XOR U7142 ( .A(n7150), .B(n7154), .Z(n7152) );
  XNOR U7143 ( .A(n7133), .B(n7130), .Z(n7143) );
  AND U7144 ( .A(n7155), .B(n7156), .Z(n7130) );
  XOR U7145 ( .A(n7157), .B(n7158), .Z(n7133) );
  AND U7146 ( .A(n7159), .B(n7160), .Z(n7158) );
  XOR U7147 ( .A(n7157), .B(n7161), .Z(n7159) );
  XNOR U7148 ( .A(n7084), .B(n7139), .Z(n7141) );
  XNOR U7149 ( .A(n7162), .B(n7163), .Z(n7084) );
  AND U7150 ( .A(n173), .B(n7164), .Z(n7163) );
  XNOR U7151 ( .A(n7165), .B(n7166), .Z(n7164) );
  XOR U7152 ( .A(n7167), .B(n7168), .Z(n7139) );
  AND U7153 ( .A(n7169), .B(n7170), .Z(n7168) );
  XNOR U7154 ( .A(n7167), .B(n7155), .Z(n7170) );
  IV U7155 ( .A(n7097), .Z(n7155) );
  XNOR U7156 ( .A(n7171), .B(n7148), .Z(n7097) );
  XNOR U7157 ( .A(n7172), .B(n7154), .Z(n7148) );
  XOR U7158 ( .A(n7173), .B(n7174), .Z(n7154) );
  AND U7159 ( .A(n7175), .B(n7176), .Z(n7174) );
  XOR U7160 ( .A(n7173), .B(n7177), .Z(n7175) );
  XNOR U7161 ( .A(n7153), .B(n7145), .Z(n7172) );
  XOR U7162 ( .A(n7178), .B(n7179), .Z(n7145) );
  AND U7163 ( .A(n7180), .B(n7181), .Z(n7179) );
  XNOR U7164 ( .A(n7182), .B(n7178), .Z(n7180) );
  XNOR U7165 ( .A(n7183), .B(n7150), .Z(n7153) );
  XOR U7166 ( .A(n7184), .B(n7185), .Z(n7150) );
  AND U7167 ( .A(n7186), .B(n7187), .Z(n7185) );
  XOR U7168 ( .A(n7184), .B(n7188), .Z(n7186) );
  XNOR U7169 ( .A(n7189), .B(n7190), .Z(n7183) );
  AND U7170 ( .A(n7191), .B(n7192), .Z(n7190) );
  XNOR U7171 ( .A(n7189), .B(n7193), .Z(n7191) );
  XNOR U7172 ( .A(n7149), .B(n7156), .Z(n7171) );
  AND U7173 ( .A(n7105), .B(n7194), .Z(n7156) );
  XOR U7174 ( .A(n7161), .B(n7160), .Z(n7149) );
  XNOR U7175 ( .A(n7195), .B(n7157), .Z(n7160) );
  XOR U7176 ( .A(n7196), .B(n7197), .Z(n7157) );
  AND U7177 ( .A(n7198), .B(n7199), .Z(n7197) );
  XOR U7178 ( .A(n7196), .B(n7200), .Z(n7198) );
  XNOR U7179 ( .A(n7201), .B(n7202), .Z(n7195) );
  AND U7180 ( .A(n7203), .B(n7204), .Z(n7202) );
  XOR U7181 ( .A(n7201), .B(n7205), .Z(n7203) );
  XOR U7182 ( .A(n7206), .B(n7207), .Z(n7161) );
  AND U7183 ( .A(n7208), .B(n7209), .Z(n7207) );
  XOR U7184 ( .A(n7206), .B(n7210), .Z(n7208) );
  XNOR U7185 ( .A(n7094), .B(n7167), .Z(n7169) );
  XNOR U7186 ( .A(n7211), .B(n7212), .Z(n7094) );
  AND U7187 ( .A(n173), .B(n7213), .Z(n7212) );
  XNOR U7188 ( .A(n7214), .B(n7215), .Z(n7213) );
  XOR U7189 ( .A(n7216), .B(n7217), .Z(n7167) );
  AND U7190 ( .A(n7218), .B(n7219), .Z(n7217) );
  XNOR U7191 ( .A(n7216), .B(n7105), .Z(n7219) );
  XOR U7192 ( .A(n7220), .B(n7181), .Z(n7105) );
  XNOR U7193 ( .A(n7221), .B(n7188), .Z(n7181) );
  XOR U7194 ( .A(n7177), .B(n7176), .Z(n7188) );
  XNOR U7195 ( .A(n7222), .B(n7173), .Z(n7176) );
  XOR U7196 ( .A(n7223), .B(n7224), .Z(n7173) );
  AND U7197 ( .A(n7225), .B(n7226), .Z(n7224) );
  XOR U7198 ( .A(n7223), .B(n7227), .Z(n7225) );
  XNOR U7199 ( .A(n7228), .B(n7229), .Z(n7222) );
  NOR U7200 ( .A(n7230), .B(n7231), .Z(n7229) );
  XNOR U7201 ( .A(n7228), .B(n7232), .Z(n7230) );
  XOR U7202 ( .A(n7233), .B(n7234), .Z(n7177) );
  NOR U7203 ( .A(n7235), .B(n7236), .Z(n7234) );
  XNOR U7204 ( .A(n7233), .B(n7237), .Z(n7235) );
  XNOR U7205 ( .A(n7187), .B(n7178), .Z(n7221) );
  XOR U7206 ( .A(n7238), .B(n7239), .Z(n7178) );
  NOR U7207 ( .A(n7240), .B(n7241), .Z(n7239) );
  XNOR U7208 ( .A(n7238), .B(n7242), .Z(n7240) );
  XOR U7209 ( .A(n7243), .B(n7193), .Z(n7187) );
  XNOR U7210 ( .A(n7244), .B(n7245), .Z(n7193) );
  NOR U7211 ( .A(n7246), .B(n7247), .Z(n7245) );
  XNOR U7212 ( .A(n7244), .B(n7248), .Z(n7246) );
  XNOR U7213 ( .A(n7192), .B(n7184), .Z(n7243) );
  XOR U7214 ( .A(n7249), .B(n7250), .Z(n7184) );
  AND U7215 ( .A(n7251), .B(n7252), .Z(n7250) );
  XOR U7216 ( .A(n7249), .B(n7253), .Z(n7251) );
  XNOR U7217 ( .A(n7254), .B(n7189), .Z(n7192) );
  XOR U7218 ( .A(n7255), .B(n7256), .Z(n7189) );
  AND U7219 ( .A(n7257), .B(n7258), .Z(n7256) );
  XOR U7220 ( .A(n7255), .B(n7259), .Z(n7257) );
  XNOR U7221 ( .A(n7260), .B(n7261), .Z(n7254) );
  NOR U7222 ( .A(n7262), .B(n7263), .Z(n7261) );
  XOR U7223 ( .A(n7260), .B(n7264), .Z(n7262) );
  XOR U7224 ( .A(n7182), .B(n7194), .Z(n7220) );
  NOR U7225 ( .A(n7111), .B(n7265), .Z(n7194) );
  XNOR U7226 ( .A(n7200), .B(n7199), .Z(n7182) );
  XNOR U7227 ( .A(n7266), .B(n7205), .Z(n7199) );
  XOR U7228 ( .A(n7267), .B(n7268), .Z(n7205) );
  NOR U7229 ( .A(n7269), .B(n7270), .Z(n7268) );
  XNOR U7230 ( .A(n7267), .B(n7271), .Z(n7269) );
  XNOR U7231 ( .A(n7204), .B(n7196), .Z(n7266) );
  XOR U7232 ( .A(n7272), .B(n7273), .Z(n7196) );
  AND U7233 ( .A(n7274), .B(n7275), .Z(n7273) );
  XNOR U7234 ( .A(n7272), .B(n7276), .Z(n7274) );
  XNOR U7235 ( .A(n7277), .B(n7201), .Z(n7204) );
  XOR U7236 ( .A(n7278), .B(n7279), .Z(n7201) );
  AND U7237 ( .A(n7280), .B(n7281), .Z(n7279) );
  XOR U7238 ( .A(n7278), .B(n7282), .Z(n7280) );
  XNOR U7239 ( .A(n7283), .B(n7284), .Z(n7277) );
  NOR U7240 ( .A(n7285), .B(n7286), .Z(n7284) );
  XOR U7241 ( .A(n7283), .B(n7287), .Z(n7285) );
  XOR U7242 ( .A(n7210), .B(n7209), .Z(n7200) );
  XNOR U7243 ( .A(n7288), .B(n7206), .Z(n7209) );
  XOR U7244 ( .A(n7289), .B(n7290), .Z(n7206) );
  AND U7245 ( .A(n7291), .B(n7292), .Z(n7290) );
  XOR U7246 ( .A(n7289), .B(n7293), .Z(n7291) );
  XNOR U7247 ( .A(n7294), .B(n7295), .Z(n7288) );
  NOR U7248 ( .A(n7296), .B(n7297), .Z(n7295) );
  XNOR U7249 ( .A(n7294), .B(n7298), .Z(n7296) );
  XOR U7250 ( .A(n7299), .B(n7300), .Z(n7210) );
  NOR U7251 ( .A(n7301), .B(n7302), .Z(n7300) );
  XNOR U7252 ( .A(n7299), .B(n7303), .Z(n7301) );
  XNOR U7253 ( .A(n7102), .B(n7216), .Z(n7218) );
  XNOR U7254 ( .A(n7304), .B(n7305), .Z(n7102) );
  AND U7255 ( .A(n173), .B(n7306), .Z(n7305) );
  XNOR U7256 ( .A(n7307), .B(n7308), .Z(n7306) );
  AND U7257 ( .A(n7108), .B(n7111), .Z(n7216) );
  XOR U7258 ( .A(n7309), .B(n7265), .Z(n7111) );
  XNOR U7259 ( .A(p_input[512]), .B(p_input[64]), .Z(n7265) );
  XOR U7260 ( .A(n7242), .B(n7241), .Z(n7309) );
  XOR U7261 ( .A(n7310), .B(n7253), .Z(n7241) );
  XOR U7262 ( .A(n7227), .B(n7226), .Z(n7253) );
  XNOR U7263 ( .A(n7311), .B(n7232), .Z(n7226) );
  XOR U7264 ( .A(p_input[536]), .B(p_input[88]), .Z(n7232) );
  XOR U7265 ( .A(n7223), .B(n7231), .Z(n7311) );
  XOR U7266 ( .A(n7312), .B(n7228), .Z(n7231) );
  XOR U7267 ( .A(p_input[534]), .B(p_input[86]), .Z(n7228) );
  XNOR U7268 ( .A(p_input[535]), .B(p_input[87]), .Z(n7312) );
  XNOR U7269 ( .A(n7313), .B(p_input[82]), .Z(n7223) );
  XNOR U7270 ( .A(n7237), .B(n7236), .Z(n7227) );
  XOR U7271 ( .A(n7314), .B(n7233), .Z(n7236) );
  XOR U7272 ( .A(p_input[531]), .B(p_input[83]), .Z(n7233) );
  XNOR U7273 ( .A(p_input[532]), .B(p_input[84]), .Z(n7314) );
  XOR U7274 ( .A(p_input[533]), .B(p_input[85]), .Z(n7237) );
  XNOR U7275 ( .A(n7252), .B(n7238), .Z(n7310) );
  XNOR U7276 ( .A(n7315), .B(p_input[65]), .Z(n7238) );
  XNOR U7277 ( .A(n7316), .B(n7259), .Z(n7252) );
  XNOR U7278 ( .A(n7248), .B(n7247), .Z(n7259) );
  XOR U7279 ( .A(n7317), .B(n7244), .Z(n7247) );
  XNOR U7280 ( .A(n6951), .B(p_input[90]), .Z(n7244) );
  XNOR U7281 ( .A(p_input[539]), .B(p_input[91]), .Z(n7317) );
  XOR U7282 ( .A(p_input[540]), .B(p_input[92]), .Z(n7248) );
  XNOR U7283 ( .A(n7258), .B(n7249), .Z(n7316) );
  XNOR U7284 ( .A(n7318), .B(p_input[81]), .Z(n7249) );
  XOR U7285 ( .A(n7319), .B(n7264), .Z(n7258) );
  XNOR U7286 ( .A(p_input[543]), .B(p_input[95]), .Z(n7264) );
  XOR U7287 ( .A(n7255), .B(n7263), .Z(n7319) );
  XOR U7288 ( .A(n7320), .B(n7260), .Z(n7263) );
  XOR U7289 ( .A(p_input[541]), .B(p_input[93]), .Z(n7260) );
  XNOR U7290 ( .A(p_input[542]), .B(p_input[94]), .Z(n7320) );
  XNOR U7291 ( .A(n6955), .B(p_input[89]), .Z(n7255) );
  XNOR U7292 ( .A(n7276), .B(n7275), .Z(n7242) );
  XNOR U7293 ( .A(n7321), .B(n7282), .Z(n7275) );
  XNOR U7294 ( .A(n7271), .B(n7270), .Z(n7282) );
  XOR U7295 ( .A(n7322), .B(n7267), .Z(n7270) );
  XNOR U7296 ( .A(n7323), .B(p_input[75]), .Z(n7267) );
  XNOR U7297 ( .A(p_input[524]), .B(p_input[76]), .Z(n7322) );
  XOR U7298 ( .A(p_input[525]), .B(p_input[77]), .Z(n7271) );
  XNOR U7299 ( .A(n7281), .B(n7272), .Z(n7321) );
  XNOR U7300 ( .A(n7324), .B(p_input[66]), .Z(n7272) );
  XOR U7301 ( .A(n7325), .B(n7287), .Z(n7281) );
  XNOR U7302 ( .A(p_input[528]), .B(p_input[80]), .Z(n7287) );
  XOR U7303 ( .A(n7278), .B(n7286), .Z(n7325) );
  XOR U7304 ( .A(n7326), .B(n7283), .Z(n7286) );
  XOR U7305 ( .A(p_input[526]), .B(p_input[78]), .Z(n7283) );
  XNOR U7306 ( .A(p_input[527]), .B(p_input[79]), .Z(n7326) );
  XNOR U7307 ( .A(n7327), .B(p_input[74]), .Z(n7278) );
  XNOR U7308 ( .A(n7293), .B(n7292), .Z(n7276) );
  XNOR U7309 ( .A(n7328), .B(n7298), .Z(n7292) );
  XOR U7310 ( .A(p_input[521]), .B(p_input[73]), .Z(n7298) );
  XOR U7311 ( .A(n7289), .B(n7297), .Z(n7328) );
  XOR U7312 ( .A(n7329), .B(n7294), .Z(n7297) );
  XOR U7313 ( .A(p_input[519]), .B(p_input[71]), .Z(n7294) );
  XNOR U7314 ( .A(p_input[520]), .B(p_input[72]), .Z(n7329) );
  XNOR U7315 ( .A(n7330), .B(p_input[67]), .Z(n7289) );
  XNOR U7316 ( .A(n7303), .B(n7302), .Z(n7293) );
  XOR U7317 ( .A(n7331), .B(n7299), .Z(n7302) );
  XOR U7318 ( .A(p_input[516]), .B(p_input[68]), .Z(n7299) );
  XNOR U7319 ( .A(p_input[517]), .B(p_input[69]), .Z(n7331) );
  XOR U7320 ( .A(p_input[518]), .B(p_input[70]), .Z(n7303) );
  XNOR U7321 ( .A(n7332), .B(n7333), .Z(n7108) );
  AND U7322 ( .A(n173), .B(n7334), .Z(n7333) );
  XNOR U7323 ( .A(n7335), .B(n7336), .Z(n173) );
  AND U7324 ( .A(n7337), .B(n7338), .Z(n7336) );
  XOR U7325 ( .A(n7122), .B(n7335), .Z(n7338) );
  XNOR U7326 ( .A(n7339), .B(n7335), .Z(n7337) );
  XOR U7327 ( .A(n7340), .B(n7341), .Z(n7335) );
  AND U7328 ( .A(n7342), .B(n7343), .Z(n7341) );
  XOR U7329 ( .A(n7137), .B(n7340), .Z(n7343) );
  XOR U7330 ( .A(n7340), .B(n7138), .Z(n7342) );
  XOR U7331 ( .A(n7344), .B(n7345), .Z(n7340) );
  AND U7332 ( .A(n7346), .B(n7347), .Z(n7345) );
  XOR U7333 ( .A(n7165), .B(n7344), .Z(n7347) );
  XOR U7334 ( .A(n7344), .B(n7166), .Z(n7346) );
  XOR U7335 ( .A(n7348), .B(n7349), .Z(n7344) );
  AND U7336 ( .A(n7350), .B(n7351), .Z(n7349) );
  XOR U7337 ( .A(n7214), .B(n7348), .Z(n7351) );
  XOR U7338 ( .A(n7348), .B(n7215), .Z(n7350) );
  XOR U7339 ( .A(n7352), .B(n7353), .Z(n7348) );
  AND U7340 ( .A(n7354), .B(n7355), .Z(n7353) );
  XOR U7341 ( .A(n7352), .B(n7307), .Z(n7355) );
  XNOR U7342 ( .A(n7356), .B(n7357), .Z(n7058) );
  AND U7343 ( .A(n177), .B(n7358), .Z(n7357) );
  XNOR U7344 ( .A(n7359), .B(n7360), .Z(n177) );
  AND U7345 ( .A(n7361), .B(n7362), .Z(n7360) );
  XOR U7346 ( .A(n7359), .B(n7068), .Z(n7362) );
  XNOR U7347 ( .A(n7359), .B(n7018), .Z(n7361) );
  XOR U7348 ( .A(n7363), .B(n7364), .Z(n7359) );
  AND U7349 ( .A(n7365), .B(n7366), .Z(n7364) );
  XNOR U7350 ( .A(n7078), .B(n7363), .Z(n7366) );
  XOR U7351 ( .A(n7363), .B(n7028), .Z(n7365) );
  XOR U7352 ( .A(n7367), .B(n7368), .Z(n7363) );
  AND U7353 ( .A(n7369), .B(n7370), .Z(n7368) );
  XNOR U7354 ( .A(n7088), .B(n7367), .Z(n7370) );
  XOR U7355 ( .A(n7367), .B(n7037), .Z(n7369) );
  XOR U7356 ( .A(n7371), .B(n7372), .Z(n7367) );
  AND U7357 ( .A(n7373), .B(n7374), .Z(n7372) );
  XOR U7358 ( .A(n7371), .B(n7045), .Z(n7373) );
  XOR U7359 ( .A(n7375), .B(n7376), .Z(n7009) );
  AND U7360 ( .A(n181), .B(n7358), .Z(n7376) );
  XNOR U7361 ( .A(n7356), .B(n7375), .Z(n7358) );
  XNOR U7362 ( .A(n7377), .B(n7378), .Z(n181) );
  AND U7363 ( .A(n7379), .B(n7380), .Z(n7378) );
  XNOR U7364 ( .A(n7381), .B(n7377), .Z(n7380) );
  IV U7365 ( .A(n7068), .Z(n7381) );
  XOR U7366 ( .A(n7339), .B(n7382), .Z(n7068) );
  AND U7367 ( .A(n184), .B(n7383), .Z(n7382) );
  XOR U7368 ( .A(n7121), .B(n7118), .Z(n7383) );
  IV U7369 ( .A(n7339), .Z(n7121) );
  XNOR U7370 ( .A(n7018), .B(n7377), .Z(n7379) );
  XOR U7371 ( .A(n7384), .B(n7385), .Z(n7018) );
  AND U7372 ( .A(n200), .B(n7386), .Z(n7385) );
  XOR U7373 ( .A(n7387), .B(n7388), .Z(n7377) );
  AND U7374 ( .A(n7389), .B(n7390), .Z(n7388) );
  XNOR U7375 ( .A(n7387), .B(n7078), .Z(n7390) );
  XOR U7376 ( .A(n7138), .B(n7391), .Z(n7078) );
  AND U7377 ( .A(n184), .B(n7392), .Z(n7391) );
  XOR U7378 ( .A(n7134), .B(n7138), .Z(n7392) );
  XNOR U7379 ( .A(n7393), .B(n7387), .Z(n7389) );
  IV U7380 ( .A(n7028), .Z(n7393) );
  XOR U7381 ( .A(n7394), .B(n7395), .Z(n7028) );
  AND U7382 ( .A(n200), .B(n7396), .Z(n7395) );
  XOR U7383 ( .A(n7397), .B(n7398), .Z(n7387) );
  AND U7384 ( .A(n7399), .B(n7400), .Z(n7398) );
  XNOR U7385 ( .A(n7397), .B(n7088), .Z(n7400) );
  XOR U7386 ( .A(n7166), .B(n7401), .Z(n7088) );
  AND U7387 ( .A(n184), .B(n7402), .Z(n7401) );
  XOR U7388 ( .A(n7162), .B(n7166), .Z(n7402) );
  XOR U7389 ( .A(n7037), .B(n7397), .Z(n7399) );
  XOR U7390 ( .A(n7403), .B(n7404), .Z(n7037) );
  AND U7391 ( .A(n200), .B(n7405), .Z(n7404) );
  XOR U7392 ( .A(n7371), .B(n7406), .Z(n7397) );
  AND U7393 ( .A(n7407), .B(n7374), .Z(n7406) );
  XNOR U7394 ( .A(n7098), .B(n7371), .Z(n7374) );
  XOR U7395 ( .A(n7215), .B(n7408), .Z(n7098) );
  AND U7396 ( .A(n184), .B(n7409), .Z(n7408) );
  XOR U7397 ( .A(n7211), .B(n7215), .Z(n7409) );
  XNOR U7398 ( .A(n7410), .B(n7371), .Z(n7407) );
  IV U7399 ( .A(n7045), .Z(n7410) );
  XOR U7400 ( .A(n7411), .B(n7412), .Z(n7045) );
  AND U7401 ( .A(n200), .B(n7413), .Z(n7412) );
  XOR U7402 ( .A(n7414), .B(n7415), .Z(n7371) );
  AND U7403 ( .A(n7416), .B(n7417), .Z(n7415) );
  XNOR U7404 ( .A(n7414), .B(n7106), .Z(n7417) );
  XOR U7405 ( .A(n7308), .B(n7418), .Z(n7106) );
  AND U7406 ( .A(n184), .B(n7419), .Z(n7418) );
  XOR U7407 ( .A(n7304), .B(n7308), .Z(n7419) );
  XNOR U7408 ( .A(n7420), .B(n7414), .Z(n7416) );
  IV U7409 ( .A(n7055), .Z(n7420) );
  XOR U7410 ( .A(n7421), .B(n7422), .Z(n7055) );
  AND U7411 ( .A(n200), .B(n7423), .Z(n7422) );
  AND U7412 ( .A(n7375), .B(n7356), .Z(n7414) );
  XNOR U7413 ( .A(n7424), .B(n7425), .Z(n7356) );
  AND U7414 ( .A(n184), .B(n7334), .Z(n7425) );
  XNOR U7415 ( .A(n7332), .B(n7424), .Z(n7334) );
  XNOR U7416 ( .A(n7426), .B(n7427), .Z(n184) );
  AND U7417 ( .A(n7428), .B(n7429), .Z(n7427) );
  XNOR U7418 ( .A(n7426), .B(n7118), .Z(n7429) );
  IV U7419 ( .A(n7122), .Z(n7118) );
  XOR U7420 ( .A(n7430), .B(n7431), .Z(n7122) );
  AND U7421 ( .A(n188), .B(n7432), .Z(n7431) );
  XOR U7422 ( .A(n7433), .B(n7430), .Z(n7432) );
  XNOR U7423 ( .A(n7426), .B(n7339), .Z(n7428) );
  XOR U7424 ( .A(n7434), .B(n7435), .Z(n7339) );
  AND U7425 ( .A(n196), .B(n7386), .Z(n7435) );
  XOR U7426 ( .A(n7384), .B(n7434), .Z(n7386) );
  XOR U7427 ( .A(n7436), .B(n7437), .Z(n7426) );
  AND U7428 ( .A(n7438), .B(n7439), .Z(n7437) );
  XNOR U7429 ( .A(n7436), .B(n7134), .Z(n7439) );
  IV U7430 ( .A(n7137), .Z(n7134) );
  XOR U7431 ( .A(n7440), .B(n7441), .Z(n7137) );
  AND U7432 ( .A(n188), .B(n7442), .Z(n7441) );
  XOR U7433 ( .A(n7443), .B(n7440), .Z(n7442) );
  XOR U7434 ( .A(n7138), .B(n7436), .Z(n7438) );
  XOR U7435 ( .A(n7444), .B(n7445), .Z(n7138) );
  AND U7436 ( .A(n196), .B(n7396), .Z(n7445) );
  XOR U7437 ( .A(n7444), .B(n7394), .Z(n7396) );
  XOR U7438 ( .A(n7446), .B(n7447), .Z(n7436) );
  AND U7439 ( .A(n7448), .B(n7449), .Z(n7447) );
  XNOR U7440 ( .A(n7446), .B(n7162), .Z(n7449) );
  IV U7441 ( .A(n7165), .Z(n7162) );
  XOR U7442 ( .A(n7450), .B(n7451), .Z(n7165) );
  AND U7443 ( .A(n188), .B(n7452), .Z(n7451) );
  XNOR U7444 ( .A(n7453), .B(n7450), .Z(n7452) );
  XOR U7445 ( .A(n7166), .B(n7446), .Z(n7448) );
  XOR U7446 ( .A(n7454), .B(n7455), .Z(n7166) );
  AND U7447 ( .A(n196), .B(n7405), .Z(n7455) );
  XOR U7448 ( .A(n7454), .B(n7403), .Z(n7405) );
  XOR U7449 ( .A(n7456), .B(n7457), .Z(n7446) );
  AND U7450 ( .A(n7458), .B(n7459), .Z(n7457) );
  XNOR U7451 ( .A(n7456), .B(n7211), .Z(n7459) );
  IV U7452 ( .A(n7214), .Z(n7211) );
  XOR U7453 ( .A(n7460), .B(n7461), .Z(n7214) );
  AND U7454 ( .A(n188), .B(n7462), .Z(n7461) );
  XOR U7455 ( .A(n7463), .B(n7460), .Z(n7462) );
  XOR U7456 ( .A(n7215), .B(n7456), .Z(n7458) );
  XOR U7457 ( .A(n7464), .B(n7465), .Z(n7215) );
  AND U7458 ( .A(n196), .B(n7413), .Z(n7465) );
  XOR U7459 ( .A(n7464), .B(n7411), .Z(n7413) );
  XOR U7460 ( .A(n7352), .B(n7466), .Z(n7456) );
  AND U7461 ( .A(n7354), .B(n7467), .Z(n7466) );
  XNOR U7462 ( .A(n7352), .B(n7304), .Z(n7467) );
  IV U7463 ( .A(n7307), .Z(n7304) );
  XOR U7464 ( .A(n7468), .B(n7469), .Z(n7307) );
  AND U7465 ( .A(n188), .B(n7470), .Z(n7469) );
  XNOR U7466 ( .A(n7471), .B(n7468), .Z(n7470) );
  XOR U7467 ( .A(n7308), .B(n7352), .Z(n7354) );
  XOR U7468 ( .A(n7472), .B(n7473), .Z(n7308) );
  AND U7469 ( .A(n196), .B(n7423), .Z(n7473) );
  XOR U7470 ( .A(n7472), .B(n7421), .Z(n7423) );
  AND U7471 ( .A(n7424), .B(n7332), .Z(n7352) );
  XNOR U7472 ( .A(n7474), .B(n7475), .Z(n7332) );
  AND U7473 ( .A(n188), .B(n7476), .Z(n7475) );
  XNOR U7474 ( .A(n7477), .B(n7474), .Z(n7476) );
  XNOR U7475 ( .A(n7478), .B(n7479), .Z(n188) );
  AND U7476 ( .A(n7480), .B(n7481), .Z(n7479) );
  XOR U7477 ( .A(n7433), .B(n7478), .Z(n7481) );
  AND U7478 ( .A(n7482), .B(n7483), .Z(n7433) );
  XNOR U7479 ( .A(n7430), .B(n7478), .Z(n7480) );
  XNOR U7480 ( .A(n7484), .B(n7485), .Z(n7430) );
  AND U7481 ( .A(n192), .B(n7486), .Z(n7485) );
  XNOR U7482 ( .A(n7487), .B(n7488), .Z(n7486) );
  XOR U7483 ( .A(n7489), .B(n7490), .Z(n7478) );
  AND U7484 ( .A(n7491), .B(n7492), .Z(n7490) );
  XNOR U7485 ( .A(n7489), .B(n7482), .Z(n7492) );
  IV U7486 ( .A(n7443), .Z(n7482) );
  XOR U7487 ( .A(n7493), .B(n7494), .Z(n7443) );
  XOR U7488 ( .A(n7495), .B(n7483), .Z(n7494) );
  AND U7489 ( .A(n7453), .B(n7496), .Z(n7483) );
  AND U7490 ( .A(n7497), .B(n7498), .Z(n7495) );
  XOR U7491 ( .A(n7499), .B(n7493), .Z(n7497) );
  XNOR U7492 ( .A(n7440), .B(n7489), .Z(n7491) );
  XNOR U7493 ( .A(n7500), .B(n7501), .Z(n7440) );
  AND U7494 ( .A(n192), .B(n7502), .Z(n7501) );
  XNOR U7495 ( .A(n7503), .B(n7504), .Z(n7502) );
  XOR U7496 ( .A(n7505), .B(n7506), .Z(n7489) );
  AND U7497 ( .A(n7507), .B(n7508), .Z(n7506) );
  XNOR U7498 ( .A(n7505), .B(n7453), .Z(n7508) );
  XOR U7499 ( .A(n7509), .B(n7498), .Z(n7453) );
  XNOR U7500 ( .A(n7510), .B(n7493), .Z(n7498) );
  XOR U7501 ( .A(n7511), .B(n7512), .Z(n7493) );
  AND U7502 ( .A(n7513), .B(n7514), .Z(n7512) );
  XOR U7503 ( .A(n7515), .B(n7511), .Z(n7513) );
  XNOR U7504 ( .A(n7516), .B(n7517), .Z(n7510) );
  AND U7505 ( .A(n7518), .B(n7519), .Z(n7517) );
  XOR U7506 ( .A(n7516), .B(n7520), .Z(n7518) );
  XNOR U7507 ( .A(n7499), .B(n7496), .Z(n7509) );
  AND U7508 ( .A(n7521), .B(n7522), .Z(n7496) );
  XOR U7509 ( .A(n7523), .B(n7524), .Z(n7499) );
  AND U7510 ( .A(n7525), .B(n7526), .Z(n7524) );
  XOR U7511 ( .A(n7523), .B(n7527), .Z(n7525) );
  XNOR U7512 ( .A(n7450), .B(n7505), .Z(n7507) );
  XNOR U7513 ( .A(n7528), .B(n7529), .Z(n7450) );
  AND U7514 ( .A(n192), .B(n7530), .Z(n7529) );
  XNOR U7515 ( .A(n7531), .B(n7532), .Z(n7530) );
  XOR U7516 ( .A(n7533), .B(n7534), .Z(n7505) );
  AND U7517 ( .A(n7535), .B(n7536), .Z(n7534) );
  XNOR U7518 ( .A(n7533), .B(n7521), .Z(n7536) );
  IV U7519 ( .A(n7463), .Z(n7521) );
  XNOR U7520 ( .A(n7537), .B(n7514), .Z(n7463) );
  XNOR U7521 ( .A(n7538), .B(n7520), .Z(n7514) );
  XOR U7522 ( .A(n7539), .B(n7540), .Z(n7520) );
  AND U7523 ( .A(n7541), .B(n7542), .Z(n7540) );
  XOR U7524 ( .A(n7539), .B(n7543), .Z(n7541) );
  XNOR U7525 ( .A(n7519), .B(n7511), .Z(n7538) );
  XOR U7526 ( .A(n7544), .B(n7545), .Z(n7511) );
  AND U7527 ( .A(n7546), .B(n7547), .Z(n7545) );
  XNOR U7528 ( .A(n7548), .B(n7544), .Z(n7546) );
  XNOR U7529 ( .A(n7549), .B(n7516), .Z(n7519) );
  XOR U7530 ( .A(n7550), .B(n7551), .Z(n7516) );
  AND U7531 ( .A(n7552), .B(n7553), .Z(n7551) );
  XOR U7532 ( .A(n7550), .B(n7554), .Z(n7552) );
  XNOR U7533 ( .A(n7555), .B(n7556), .Z(n7549) );
  AND U7534 ( .A(n7557), .B(n7558), .Z(n7556) );
  XNOR U7535 ( .A(n7555), .B(n7559), .Z(n7557) );
  XNOR U7536 ( .A(n7515), .B(n7522), .Z(n7537) );
  AND U7537 ( .A(n7471), .B(n7560), .Z(n7522) );
  XOR U7538 ( .A(n7527), .B(n7526), .Z(n7515) );
  XNOR U7539 ( .A(n7561), .B(n7523), .Z(n7526) );
  XOR U7540 ( .A(n7562), .B(n7563), .Z(n7523) );
  AND U7541 ( .A(n7564), .B(n7565), .Z(n7563) );
  XOR U7542 ( .A(n7562), .B(n7566), .Z(n7564) );
  XNOR U7543 ( .A(n7567), .B(n7568), .Z(n7561) );
  AND U7544 ( .A(n7569), .B(n7570), .Z(n7568) );
  XOR U7545 ( .A(n7567), .B(n7571), .Z(n7569) );
  XOR U7546 ( .A(n7572), .B(n7573), .Z(n7527) );
  AND U7547 ( .A(n7574), .B(n7575), .Z(n7573) );
  XOR U7548 ( .A(n7572), .B(n7576), .Z(n7574) );
  XNOR U7549 ( .A(n7460), .B(n7533), .Z(n7535) );
  XNOR U7550 ( .A(n7577), .B(n7578), .Z(n7460) );
  AND U7551 ( .A(n192), .B(n7579), .Z(n7578) );
  XNOR U7552 ( .A(n7580), .B(n7581), .Z(n7579) );
  XOR U7553 ( .A(n7582), .B(n7583), .Z(n7533) );
  AND U7554 ( .A(n7584), .B(n7585), .Z(n7583) );
  XNOR U7555 ( .A(n7582), .B(n7471), .Z(n7585) );
  XOR U7556 ( .A(n7586), .B(n7547), .Z(n7471) );
  XNOR U7557 ( .A(n7587), .B(n7554), .Z(n7547) );
  XOR U7558 ( .A(n7543), .B(n7542), .Z(n7554) );
  XNOR U7559 ( .A(n7588), .B(n7539), .Z(n7542) );
  XOR U7560 ( .A(n7589), .B(n7590), .Z(n7539) );
  AND U7561 ( .A(n7591), .B(n7592), .Z(n7590) );
  XNOR U7562 ( .A(n7593), .B(n7594), .Z(n7591) );
  IV U7563 ( .A(n7589), .Z(n7593) );
  XNOR U7564 ( .A(n7595), .B(n7596), .Z(n7588) );
  NOR U7565 ( .A(n7597), .B(n7598), .Z(n7596) );
  XNOR U7566 ( .A(n7595), .B(n7599), .Z(n7597) );
  XOR U7567 ( .A(n7600), .B(n7601), .Z(n7543) );
  NOR U7568 ( .A(n7602), .B(n7603), .Z(n7601) );
  XNOR U7569 ( .A(n7600), .B(n7604), .Z(n7602) );
  XNOR U7570 ( .A(n7553), .B(n7544), .Z(n7587) );
  XOR U7571 ( .A(n7605), .B(n7606), .Z(n7544) );
  AND U7572 ( .A(n7607), .B(n7608), .Z(n7606) );
  XOR U7573 ( .A(n7605), .B(n7609), .Z(n7607) );
  XOR U7574 ( .A(n7610), .B(n7559), .Z(n7553) );
  XOR U7575 ( .A(n7611), .B(n7612), .Z(n7559) );
  NOR U7576 ( .A(n7613), .B(n7614), .Z(n7612) );
  XOR U7577 ( .A(n7611), .B(n7615), .Z(n7613) );
  XNOR U7578 ( .A(n7558), .B(n7550), .Z(n7610) );
  XOR U7579 ( .A(n7616), .B(n7617), .Z(n7550) );
  AND U7580 ( .A(n7618), .B(n7619), .Z(n7617) );
  XOR U7581 ( .A(n7616), .B(n7620), .Z(n7618) );
  XNOR U7582 ( .A(n7621), .B(n7555), .Z(n7558) );
  XOR U7583 ( .A(n7622), .B(n7623), .Z(n7555) );
  AND U7584 ( .A(n7624), .B(n7625), .Z(n7623) );
  XNOR U7585 ( .A(n7626), .B(n7627), .Z(n7624) );
  IV U7586 ( .A(n7622), .Z(n7626) );
  XNOR U7587 ( .A(n7628), .B(n7629), .Z(n7621) );
  NOR U7588 ( .A(n7630), .B(n7631), .Z(n7629) );
  XNOR U7589 ( .A(n7628), .B(n7632), .Z(n7630) );
  XOR U7590 ( .A(n7548), .B(n7560), .Z(n7586) );
  NOR U7591 ( .A(n7477), .B(n7633), .Z(n7560) );
  XNOR U7592 ( .A(n7566), .B(n7565), .Z(n7548) );
  XNOR U7593 ( .A(n7634), .B(n7571), .Z(n7565) );
  XNOR U7594 ( .A(n7635), .B(n7636), .Z(n7571) );
  NOR U7595 ( .A(n7637), .B(n7638), .Z(n7636) );
  XOR U7596 ( .A(n7635), .B(n7639), .Z(n7637) );
  XNOR U7597 ( .A(n7570), .B(n7562), .Z(n7634) );
  XOR U7598 ( .A(n7640), .B(n7641), .Z(n7562) );
  AND U7599 ( .A(n7642), .B(n7643), .Z(n7641) );
  XOR U7600 ( .A(n7640), .B(n7644), .Z(n7642) );
  XNOR U7601 ( .A(n7645), .B(n7567), .Z(n7570) );
  XOR U7602 ( .A(n7646), .B(n7647), .Z(n7567) );
  AND U7603 ( .A(n7648), .B(n7649), .Z(n7647) );
  XNOR U7604 ( .A(n7650), .B(n7651), .Z(n7648) );
  IV U7605 ( .A(n7646), .Z(n7650) );
  XNOR U7606 ( .A(n7652), .B(n7653), .Z(n7645) );
  NOR U7607 ( .A(n7654), .B(n7655), .Z(n7653) );
  XNOR U7608 ( .A(n7652), .B(n7656), .Z(n7654) );
  XOR U7609 ( .A(n7576), .B(n7575), .Z(n7566) );
  XNOR U7610 ( .A(n7657), .B(n7572), .Z(n7575) );
  XOR U7611 ( .A(n7658), .B(n7659), .Z(n7572) );
  AND U7612 ( .A(n7660), .B(n7661), .Z(n7659) );
  XOR U7613 ( .A(n7658), .B(n7662), .Z(n7660) );
  XNOR U7614 ( .A(n7663), .B(n7664), .Z(n7657) );
  NOR U7615 ( .A(n7665), .B(n7666), .Z(n7664) );
  XNOR U7616 ( .A(n7663), .B(n7667), .Z(n7665) );
  XOR U7617 ( .A(n7668), .B(n7669), .Z(n7576) );
  NOR U7618 ( .A(n7670), .B(n7671), .Z(n7669) );
  XNOR U7619 ( .A(n7668), .B(n7672), .Z(n7670) );
  XNOR U7620 ( .A(n7468), .B(n7582), .Z(n7584) );
  XNOR U7621 ( .A(n7673), .B(n7674), .Z(n7468) );
  AND U7622 ( .A(n192), .B(n7675), .Z(n7674) );
  XNOR U7623 ( .A(n7676), .B(n7677), .Z(n7675) );
  AND U7624 ( .A(n7474), .B(n7477), .Z(n7582) );
  XOR U7625 ( .A(n7678), .B(n7633), .Z(n7477) );
  XNOR U7626 ( .A(p_input[512]), .B(p_input[96]), .Z(n7633) );
  XNOR U7627 ( .A(n7609), .B(n7608), .Z(n7678) );
  XNOR U7628 ( .A(n7679), .B(n7620), .Z(n7608) );
  XOR U7629 ( .A(n7594), .B(n7592), .Z(n7620) );
  XNOR U7630 ( .A(n7680), .B(n7599), .Z(n7592) );
  XOR U7631 ( .A(p_input[120]), .B(p_input[536]), .Z(n7599) );
  XOR U7632 ( .A(n7589), .B(n7598), .Z(n7680) );
  XOR U7633 ( .A(n7681), .B(n7595), .Z(n7598) );
  XOR U7634 ( .A(p_input[118]), .B(p_input[534]), .Z(n7595) );
  XOR U7635 ( .A(p_input[119]), .B(n6576), .Z(n7681) );
  XOR U7636 ( .A(p_input[114]), .B(p_input[530]), .Z(n7589) );
  XNOR U7637 ( .A(n7604), .B(n7603), .Z(n7594) );
  XOR U7638 ( .A(n7682), .B(n7600), .Z(n7603) );
  XOR U7639 ( .A(p_input[115]), .B(p_input[531]), .Z(n7600) );
  XOR U7640 ( .A(p_input[116]), .B(n6578), .Z(n7682) );
  XOR U7641 ( .A(p_input[117]), .B(p_input[533]), .Z(n7604) );
  XNOR U7642 ( .A(n7619), .B(n7605), .Z(n7679) );
  XNOR U7643 ( .A(n7315), .B(p_input[97]), .Z(n7605) );
  XNOR U7644 ( .A(n7683), .B(n7627), .Z(n7619) );
  XNOR U7645 ( .A(n7615), .B(n7614), .Z(n7627) );
  XNOR U7646 ( .A(n7684), .B(n7611), .Z(n7614) );
  XNOR U7647 ( .A(p_input[122]), .B(p_input[538]), .Z(n7611) );
  XOR U7648 ( .A(p_input[123]), .B(n6582), .Z(n7684) );
  XOR U7649 ( .A(p_input[124]), .B(p_input[540]), .Z(n7615) );
  XOR U7650 ( .A(n7625), .B(n7685), .Z(n7683) );
  IV U7651 ( .A(n7616), .Z(n7685) );
  XOR U7652 ( .A(p_input[113]), .B(p_input[529]), .Z(n7616) );
  XNOR U7653 ( .A(n7686), .B(n7632), .Z(n7625) );
  XNOR U7654 ( .A(p_input[127]), .B(n6585), .Z(n7632) );
  XOR U7655 ( .A(n7622), .B(n7631), .Z(n7686) );
  XOR U7656 ( .A(n7687), .B(n7628), .Z(n7631) );
  XOR U7657 ( .A(p_input[125]), .B(p_input[541]), .Z(n7628) );
  XOR U7658 ( .A(p_input[126]), .B(n6587), .Z(n7687) );
  XOR U7659 ( .A(p_input[121]), .B(p_input[537]), .Z(n7622) );
  XOR U7660 ( .A(n7644), .B(n7643), .Z(n7609) );
  XNOR U7661 ( .A(n7688), .B(n7651), .Z(n7643) );
  XNOR U7662 ( .A(n7639), .B(n7638), .Z(n7651) );
  XNOR U7663 ( .A(n7689), .B(n7635), .Z(n7638) );
  XNOR U7664 ( .A(p_input[107]), .B(p_input[523]), .Z(n7635) );
  XOR U7665 ( .A(p_input[108]), .B(n6590), .Z(n7689) );
  XOR U7666 ( .A(p_input[109]), .B(p_input[525]), .Z(n7639) );
  XNOR U7667 ( .A(n7649), .B(n7640), .Z(n7688) );
  XNOR U7668 ( .A(n7324), .B(p_input[98]), .Z(n7640) );
  XNOR U7669 ( .A(n7690), .B(n7656), .Z(n7649) );
  XNOR U7670 ( .A(p_input[112]), .B(n6593), .Z(n7656) );
  XOR U7671 ( .A(n7646), .B(n7655), .Z(n7690) );
  XOR U7672 ( .A(n7691), .B(n7652), .Z(n7655) );
  XOR U7673 ( .A(p_input[110]), .B(p_input[526]), .Z(n7652) );
  XOR U7674 ( .A(p_input[111]), .B(n6595), .Z(n7691) );
  XOR U7675 ( .A(p_input[106]), .B(p_input[522]), .Z(n7646) );
  XOR U7676 ( .A(n7662), .B(n7661), .Z(n7644) );
  XNOR U7677 ( .A(n7692), .B(n7667), .Z(n7661) );
  XOR U7678 ( .A(p_input[105]), .B(p_input[521]), .Z(n7667) );
  XOR U7679 ( .A(n7658), .B(n7666), .Z(n7692) );
  XOR U7680 ( .A(n7693), .B(n7663), .Z(n7666) );
  XOR U7681 ( .A(p_input[103]), .B(p_input[519]), .Z(n7663) );
  XOR U7682 ( .A(p_input[104]), .B(n6963), .Z(n7693) );
  XNOR U7683 ( .A(n7330), .B(p_input[99]), .Z(n7658) );
  XNOR U7684 ( .A(n7672), .B(n7671), .Z(n7662) );
  XOR U7685 ( .A(n7694), .B(n7668), .Z(n7671) );
  XOR U7686 ( .A(p_input[100]), .B(p_input[516]), .Z(n7668) );
  XOR U7687 ( .A(p_input[101]), .B(n6965), .Z(n7694) );
  XOR U7688 ( .A(p_input[102]), .B(p_input[518]), .Z(n7672) );
  XNOR U7689 ( .A(n7695), .B(n7696), .Z(n7474) );
  AND U7690 ( .A(n192), .B(n7697), .Z(n7696) );
  XNOR U7691 ( .A(n7698), .B(n7699), .Z(n192) );
  AND U7692 ( .A(n7700), .B(n7701), .Z(n7699) );
  XOR U7693 ( .A(n7488), .B(n7698), .Z(n7701) );
  XNOR U7694 ( .A(n7702), .B(n7698), .Z(n7700) );
  XOR U7695 ( .A(n7703), .B(n7704), .Z(n7698) );
  AND U7696 ( .A(n7705), .B(n7706), .Z(n7704) );
  XOR U7697 ( .A(n7503), .B(n7703), .Z(n7706) );
  XOR U7698 ( .A(n7703), .B(n7504), .Z(n7705) );
  XOR U7699 ( .A(n7707), .B(n7708), .Z(n7703) );
  AND U7700 ( .A(n7709), .B(n7710), .Z(n7708) );
  XOR U7701 ( .A(n7531), .B(n7707), .Z(n7710) );
  XOR U7702 ( .A(n7707), .B(n7532), .Z(n7709) );
  XOR U7703 ( .A(n7711), .B(n7712), .Z(n7707) );
  AND U7704 ( .A(n7713), .B(n7714), .Z(n7712) );
  XOR U7705 ( .A(n7580), .B(n7711), .Z(n7714) );
  XOR U7706 ( .A(n7711), .B(n7581), .Z(n7713) );
  XOR U7707 ( .A(n7715), .B(n7716), .Z(n7711) );
  AND U7708 ( .A(n7717), .B(n7718), .Z(n7716) );
  XOR U7709 ( .A(n7715), .B(n7676), .Z(n7718) );
  XNOR U7710 ( .A(n7719), .B(n7720), .Z(n7424) );
  AND U7711 ( .A(n196), .B(n7721), .Z(n7720) );
  XNOR U7712 ( .A(n7722), .B(n7723), .Z(n196) );
  AND U7713 ( .A(n7724), .B(n7725), .Z(n7723) );
  XOR U7714 ( .A(n7722), .B(n7434), .Z(n7725) );
  XNOR U7715 ( .A(n7722), .B(n7384), .Z(n7724) );
  XOR U7716 ( .A(n7726), .B(n7727), .Z(n7722) );
  AND U7717 ( .A(n7728), .B(n7729), .Z(n7727) );
  XNOR U7718 ( .A(n7444), .B(n7726), .Z(n7729) );
  XOR U7719 ( .A(n7726), .B(n7394), .Z(n7728) );
  XOR U7720 ( .A(n7730), .B(n7731), .Z(n7726) );
  AND U7721 ( .A(n7732), .B(n7733), .Z(n7731) );
  XNOR U7722 ( .A(n7454), .B(n7730), .Z(n7733) );
  XOR U7723 ( .A(n7730), .B(n7403), .Z(n7732) );
  XOR U7724 ( .A(n7734), .B(n7735), .Z(n7730) );
  AND U7725 ( .A(n7736), .B(n7737), .Z(n7735) );
  XOR U7726 ( .A(n7734), .B(n7411), .Z(n7736) );
  XOR U7727 ( .A(n7738), .B(n7739), .Z(n7375) );
  AND U7728 ( .A(n200), .B(n7721), .Z(n7739) );
  XNOR U7729 ( .A(n7719), .B(n7738), .Z(n7721) );
  XNOR U7730 ( .A(n7740), .B(n7741), .Z(n200) );
  AND U7731 ( .A(n7742), .B(n7743), .Z(n7741) );
  XNOR U7732 ( .A(n7744), .B(n7740), .Z(n7743) );
  IV U7733 ( .A(n7434), .Z(n7744) );
  XOR U7734 ( .A(n7702), .B(n7745), .Z(n7434) );
  AND U7735 ( .A(n203), .B(n7746), .Z(n7745) );
  XOR U7736 ( .A(n7487), .B(n7484), .Z(n7746) );
  IV U7737 ( .A(n7702), .Z(n7487) );
  XNOR U7738 ( .A(n7384), .B(n7740), .Z(n7742) );
  XOR U7739 ( .A(n7747), .B(n7748), .Z(n7384) );
  AND U7740 ( .A(n219), .B(n7749), .Z(n7748) );
  XOR U7741 ( .A(n7750), .B(n7751), .Z(n7740) );
  AND U7742 ( .A(n7752), .B(n7753), .Z(n7751) );
  XNOR U7743 ( .A(n7750), .B(n7444), .Z(n7753) );
  XOR U7744 ( .A(n7504), .B(n7754), .Z(n7444) );
  AND U7745 ( .A(n203), .B(n7755), .Z(n7754) );
  XOR U7746 ( .A(n7500), .B(n7504), .Z(n7755) );
  XNOR U7747 ( .A(n7756), .B(n7750), .Z(n7752) );
  IV U7748 ( .A(n7394), .Z(n7756) );
  XOR U7749 ( .A(n7757), .B(n7758), .Z(n7394) );
  AND U7750 ( .A(n219), .B(n7759), .Z(n7758) );
  XOR U7751 ( .A(n7760), .B(n7761), .Z(n7750) );
  AND U7752 ( .A(n7762), .B(n7763), .Z(n7761) );
  XNOR U7753 ( .A(n7760), .B(n7454), .Z(n7763) );
  XOR U7754 ( .A(n7532), .B(n7764), .Z(n7454) );
  AND U7755 ( .A(n203), .B(n7765), .Z(n7764) );
  XOR U7756 ( .A(n7528), .B(n7532), .Z(n7765) );
  XOR U7757 ( .A(n7403), .B(n7760), .Z(n7762) );
  XOR U7758 ( .A(n7766), .B(n7767), .Z(n7403) );
  AND U7759 ( .A(n219), .B(n7768), .Z(n7767) );
  XOR U7760 ( .A(n7734), .B(n7769), .Z(n7760) );
  AND U7761 ( .A(n7770), .B(n7737), .Z(n7769) );
  XNOR U7762 ( .A(n7464), .B(n7734), .Z(n7737) );
  XOR U7763 ( .A(n7581), .B(n7771), .Z(n7464) );
  AND U7764 ( .A(n203), .B(n7772), .Z(n7771) );
  XOR U7765 ( .A(n7577), .B(n7581), .Z(n7772) );
  XNOR U7766 ( .A(n7773), .B(n7734), .Z(n7770) );
  IV U7767 ( .A(n7411), .Z(n7773) );
  XOR U7768 ( .A(n7774), .B(n7775), .Z(n7411) );
  AND U7769 ( .A(n219), .B(n7776), .Z(n7775) );
  XOR U7770 ( .A(n7777), .B(n7778), .Z(n7734) );
  AND U7771 ( .A(n7779), .B(n7780), .Z(n7778) );
  XNOR U7772 ( .A(n7777), .B(n7472), .Z(n7780) );
  XOR U7773 ( .A(n7677), .B(n7781), .Z(n7472) );
  AND U7774 ( .A(n203), .B(n7782), .Z(n7781) );
  XOR U7775 ( .A(n7673), .B(n7677), .Z(n7782) );
  XNOR U7776 ( .A(n7783), .B(n7777), .Z(n7779) );
  IV U7777 ( .A(n7421), .Z(n7783) );
  XOR U7778 ( .A(n7784), .B(n7785), .Z(n7421) );
  AND U7779 ( .A(n219), .B(n7786), .Z(n7785) );
  AND U7780 ( .A(n7738), .B(n7719), .Z(n7777) );
  XNOR U7781 ( .A(n7787), .B(n7788), .Z(n7719) );
  AND U7782 ( .A(n203), .B(n7697), .Z(n7788) );
  XNOR U7783 ( .A(n7695), .B(n7787), .Z(n7697) );
  XNOR U7784 ( .A(n7789), .B(n7790), .Z(n203) );
  AND U7785 ( .A(n7791), .B(n7792), .Z(n7790) );
  XNOR U7786 ( .A(n7789), .B(n7484), .Z(n7792) );
  IV U7787 ( .A(n7488), .Z(n7484) );
  XOR U7788 ( .A(n7793), .B(n7794), .Z(n7488) );
  AND U7789 ( .A(n207), .B(n7795), .Z(n7794) );
  XOR U7790 ( .A(n7796), .B(n7793), .Z(n7795) );
  XNOR U7791 ( .A(n7789), .B(n7702), .Z(n7791) );
  XOR U7792 ( .A(n7797), .B(n7798), .Z(n7702) );
  AND U7793 ( .A(n215), .B(n7749), .Z(n7798) );
  XOR U7794 ( .A(n7747), .B(n7797), .Z(n7749) );
  XOR U7795 ( .A(n7799), .B(n7800), .Z(n7789) );
  AND U7796 ( .A(n7801), .B(n7802), .Z(n7800) );
  XNOR U7797 ( .A(n7799), .B(n7500), .Z(n7802) );
  IV U7798 ( .A(n7503), .Z(n7500) );
  XOR U7799 ( .A(n7803), .B(n7804), .Z(n7503) );
  AND U7800 ( .A(n207), .B(n7805), .Z(n7804) );
  XOR U7801 ( .A(n7806), .B(n7803), .Z(n7805) );
  XOR U7802 ( .A(n7504), .B(n7799), .Z(n7801) );
  XOR U7803 ( .A(n7807), .B(n7808), .Z(n7504) );
  AND U7804 ( .A(n215), .B(n7759), .Z(n7808) );
  XOR U7805 ( .A(n7807), .B(n7757), .Z(n7759) );
  XOR U7806 ( .A(n7809), .B(n7810), .Z(n7799) );
  AND U7807 ( .A(n7811), .B(n7812), .Z(n7810) );
  XNOR U7808 ( .A(n7809), .B(n7528), .Z(n7812) );
  IV U7809 ( .A(n7531), .Z(n7528) );
  XOR U7810 ( .A(n7813), .B(n7814), .Z(n7531) );
  AND U7811 ( .A(n207), .B(n7815), .Z(n7814) );
  XNOR U7812 ( .A(n7816), .B(n7813), .Z(n7815) );
  XOR U7813 ( .A(n7532), .B(n7809), .Z(n7811) );
  XOR U7814 ( .A(n7817), .B(n7818), .Z(n7532) );
  AND U7815 ( .A(n215), .B(n7768), .Z(n7818) );
  XOR U7816 ( .A(n7817), .B(n7766), .Z(n7768) );
  XOR U7817 ( .A(n7819), .B(n7820), .Z(n7809) );
  AND U7818 ( .A(n7821), .B(n7822), .Z(n7820) );
  XNOR U7819 ( .A(n7819), .B(n7577), .Z(n7822) );
  IV U7820 ( .A(n7580), .Z(n7577) );
  XOR U7821 ( .A(n7823), .B(n7824), .Z(n7580) );
  AND U7822 ( .A(n207), .B(n7825), .Z(n7824) );
  XOR U7823 ( .A(n7826), .B(n7823), .Z(n7825) );
  XOR U7824 ( .A(n7581), .B(n7819), .Z(n7821) );
  XOR U7825 ( .A(n7827), .B(n7828), .Z(n7581) );
  AND U7826 ( .A(n215), .B(n7776), .Z(n7828) );
  XOR U7827 ( .A(n7827), .B(n7774), .Z(n7776) );
  XOR U7828 ( .A(n7715), .B(n7829), .Z(n7819) );
  AND U7829 ( .A(n7717), .B(n7830), .Z(n7829) );
  XNOR U7830 ( .A(n7715), .B(n7673), .Z(n7830) );
  IV U7831 ( .A(n7676), .Z(n7673) );
  XOR U7832 ( .A(n7831), .B(n7832), .Z(n7676) );
  AND U7833 ( .A(n207), .B(n7833), .Z(n7832) );
  XNOR U7834 ( .A(n7834), .B(n7831), .Z(n7833) );
  XOR U7835 ( .A(n7677), .B(n7715), .Z(n7717) );
  XOR U7836 ( .A(n7835), .B(n7836), .Z(n7677) );
  AND U7837 ( .A(n215), .B(n7786), .Z(n7836) );
  XOR U7838 ( .A(n7835), .B(n7784), .Z(n7786) );
  AND U7839 ( .A(n7787), .B(n7695), .Z(n7715) );
  XNOR U7840 ( .A(n7837), .B(n7838), .Z(n7695) );
  AND U7841 ( .A(n207), .B(n7839), .Z(n7838) );
  XNOR U7842 ( .A(n7840), .B(n7837), .Z(n7839) );
  XNOR U7843 ( .A(n7841), .B(n7842), .Z(n207) );
  AND U7844 ( .A(n7843), .B(n7844), .Z(n7842) );
  XOR U7845 ( .A(n7796), .B(n7841), .Z(n7844) );
  AND U7846 ( .A(n7845), .B(n7846), .Z(n7796) );
  XNOR U7847 ( .A(n7793), .B(n7841), .Z(n7843) );
  XNOR U7848 ( .A(n7847), .B(n7848), .Z(n7793) );
  AND U7849 ( .A(n211), .B(n7849), .Z(n7848) );
  XNOR U7850 ( .A(n7850), .B(n7851), .Z(n7849) );
  XOR U7851 ( .A(n7852), .B(n7853), .Z(n7841) );
  AND U7852 ( .A(n7854), .B(n7855), .Z(n7853) );
  XNOR U7853 ( .A(n7852), .B(n7845), .Z(n7855) );
  IV U7854 ( .A(n7806), .Z(n7845) );
  XOR U7855 ( .A(n7856), .B(n7857), .Z(n7806) );
  XOR U7856 ( .A(n7858), .B(n7846), .Z(n7857) );
  AND U7857 ( .A(n7816), .B(n7859), .Z(n7846) );
  AND U7858 ( .A(n7860), .B(n7861), .Z(n7858) );
  XOR U7859 ( .A(n7862), .B(n7856), .Z(n7860) );
  XNOR U7860 ( .A(n7803), .B(n7852), .Z(n7854) );
  XNOR U7861 ( .A(n7863), .B(n7864), .Z(n7803) );
  AND U7862 ( .A(n211), .B(n7865), .Z(n7864) );
  XNOR U7863 ( .A(n7866), .B(n7867), .Z(n7865) );
  XOR U7864 ( .A(n7868), .B(n7869), .Z(n7852) );
  AND U7865 ( .A(n7870), .B(n7871), .Z(n7869) );
  XNOR U7866 ( .A(n7868), .B(n7816), .Z(n7871) );
  XOR U7867 ( .A(n7872), .B(n7861), .Z(n7816) );
  XNOR U7868 ( .A(n7873), .B(n7856), .Z(n7861) );
  XOR U7869 ( .A(n7874), .B(n7875), .Z(n7856) );
  AND U7870 ( .A(n7876), .B(n7877), .Z(n7875) );
  XOR U7871 ( .A(n7878), .B(n7874), .Z(n7876) );
  XNOR U7872 ( .A(n7879), .B(n7880), .Z(n7873) );
  AND U7873 ( .A(n7881), .B(n7882), .Z(n7880) );
  XOR U7874 ( .A(n7879), .B(n7883), .Z(n7881) );
  XNOR U7875 ( .A(n7862), .B(n7859), .Z(n7872) );
  AND U7876 ( .A(n7884), .B(n7885), .Z(n7859) );
  XOR U7877 ( .A(n7886), .B(n7887), .Z(n7862) );
  AND U7878 ( .A(n7888), .B(n7889), .Z(n7887) );
  XOR U7879 ( .A(n7886), .B(n7890), .Z(n7888) );
  XNOR U7880 ( .A(n7813), .B(n7868), .Z(n7870) );
  XNOR U7881 ( .A(n7891), .B(n7892), .Z(n7813) );
  AND U7882 ( .A(n211), .B(n7893), .Z(n7892) );
  XNOR U7883 ( .A(n7894), .B(n7895), .Z(n7893) );
  XOR U7884 ( .A(n7896), .B(n7897), .Z(n7868) );
  AND U7885 ( .A(n7898), .B(n7899), .Z(n7897) );
  XNOR U7886 ( .A(n7896), .B(n7884), .Z(n7899) );
  IV U7887 ( .A(n7826), .Z(n7884) );
  XNOR U7888 ( .A(n7900), .B(n7877), .Z(n7826) );
  XNOR U7889 ( .A(n7901), .B(n7883), .Z(n7877) );
  XOR U7890 ( .A(n7902), .B(n7903), .Z(n7883) );
  AND U7891 ( .A(n7904), .B(n7905), .Z(n7903) );
  XOR U7892 ( .A(n7902), .B(n7906), .Z(n7904) );
  XNOR U7893 ( .A(n7882), .B(n7874), .Z(n7901) );
  XOR U7894 ( .A(n7907), .B(n7908), .Z(n7874) );
  AND U7895 ( .A(n7909), .B(n7910), .Z(n7908) );
  XNOR U7896 ( .A(n7911), .B(n7907), .Z(n7909) );
  XNOR U7897 ( .A(n7912), .B(n7879), .Z(n7882) );
  XOR U7898 ( .A(n7913), .B(n7914), .Z(n7879) );
  AND U7899 ( .A(n7915), .B(n7916), .Z(n7914) );
  XOR U7900 ( .A(n7913), .B(n7917), .Z(n7915) );
  XNOR U7901 ( .A(n7918), .B(n7919), .Z(n7912) );
  AND U7902 ( .A(n7920), .B(n7921), .Z(n7919) );
  XNOR U7903 ( .A(n7918), .B(n7922), .Z(n7920) );
  XNOR U7904 ( .A(n7878), .B(n7885), .Z(n7900) );
  AND U7905 ( .A(n7834), .B(n7923), .Z(n7885) );
  XOR U7906 ( .A(n7890), .B(n7889), .Z(n7878) );
  XNOR U7907 ( .A(n7924), .B(n7886), .Z(n7889) );
  XOR U7908 ( .A(n7925), .B(n7926), .Z(n7886) );
  AND U7909 ( .A(n7927), .B(n7928), .Z(n7926) );
  XOR U7910 ( .A(n7925), .B(n7929), .Z(n7927) );
  XNOR U7911 ( .A(n7930), .B(n7931), .Z(n7924) );
  AND U7912 ( .A(n7932), .B(n7933), .Z(n7931) );
  XOR U7913 ( .A(n7930), .B(n7934), .Z(n7932) );
  XOR U7914 ( .A(n7935), .B(n7936), .Z(n7890) );
  AND U7915 ( .A(n7937), .B(n7938), .Z(n7936) );
  XOR U7916 ( .A(n7935), .B(n7939), .Z(n7937) );
  XNOR U7917 ( .A(n7823), .B(n7896), .Z(n7898) );
  XNOR U7918 ( .A(n7940), .B(n7941), .Z(n7823) );
  AND U7919 ( .A(n211), .B(n7942), .Z(n7941) );
  XNOR U7920 ( .A(n7943), .B(n7944), .Z(n7942) );
  XOR U7921 ( .A(n7945), .B(n7946), .Z(n7896) );
  AND U7922 ( .A(n7947), .B(n7948), .Z(n7946) );
  XNOR U7923 ( .A(n7945), .B(n7834), .Z(n7948) );
  XOR U7924 ( .A(n7949), .B(n7910), .Z(n7834) );
  XNOR U7925 ( .A(n7950), .B(n7917), .Z(n7910) );
  XOR U7926 ( .A(n7906), .B(n7905), .Z(n7917) );
  XNOR U7927 ( .A(n7951), .B(n7902), .Z(n7905) );
  XOR U7928 ( .A(n7952), .B(n7953), .Z(n7902) );
  AND U7929 ( .A(n7954), .B(n7955), .Z(n7953) );
  XNOR U7930 ( .A(n7956), .B(n7957), .Z(n7954) );
  IV U7931 ( .A(n7952), .Z(n7956) );
  XNOR U7932 ( .A(n7958), .B(n7959), .Z(n7951) );
  NOR U7933 ( .A(n7960), .B(n7961), .Z(n7959) );
  XNOR U7934 ( .A(n7958), .B(n7962), .Z(n7960) );
  XOR U7935 ( .A(n7963), .B(n7964), .Z(n7906) );
  NOR U7936 ( .A(n7965), .B(n7966), .Z(n7964) );
  XNOR U7937 ( .A(n7963), .B(n7967), .Z(n7965) );
  XNOR U7938 ( .A(n7916), .B(n7907), .Z(n7950) );
  XOR U7939 ( .A(n7968), .B(n7969), .Z(n7907) );
  AND U7940 ( .A(n7970), .B(n7971), .Z(n7969) );
  XOR U7941 ( .A(n7968), .B(n7972), .Z(n7970) );
  XOR U7942 ( .A(n7973), .B(n7922), .Z(n7916) );
  XOR U7943 ( .A(n7974), .B(n7975), .Z(n7922) );
  NOR U7944 ( .A(n7976), .B(n7977), .Z(n7975) );
  XOR U7945 ( .A(n7974), .B(n7978), .Z(n7976) );
  XNOR U7946 ( .A(n7921), .B(n7913), .Z(n7973) );
  XOR U7947 ( .A(n7979), .B(n7980), .Z(n7913) );
  AND U7948 ( .A(n7981), .B(n7982), .Z(n7980) );
  XOR U7949 ( .A(n7979), .B(n7983), .Z(n7981) );
  XNOR U7950 ( .A(n7984), .B(n7918), .Z(n7921) );
  XOR U7951 ( .A(n7985), .B(n7986), .Z(n7918) );
  AND U7952 ( .A(n7987), .B(n7988), .Z(n7986) );
  XNOR U7953 ( .A(n7989), .B(n7990), .Z(n7987) );
  IV U7954 ( .A(n7985), .Z(n7989) );
  XNOR U7955 ( .A(n7991), .B(n7992), .Z(n7984) );
  NOR U7956 ( .A(n7993), .B(n7994), .Z(n7992) );
  XNOR U7957 ( .A(n7991), .B(n7995), .Z(n7993) );
  XOR U7958 ( .A(n7911), .B(n7923), .Z(n7949) );
  NOR U7959 ( .A(n7840), .B(n7996), .Z(n7923) );
  XNOR U7960 ( .A(n7929), .B(n7928), .Z(n7911) );
  XNOR U7961 ( .A(n7997), .B(n7934), .Z(n7928) );
  XNOR U7962 ( .A(n7998), .B(n7999), .Z(n7934) );
  NOR U7963 ( .A(n8000), .B(n8001), .Z(n7999) );
  XOR U7964 ( .A(n7998), .B(n8002), .Z(n8000) );
  XNOR U7965 ( .A(n7933), .B(n7925), .Z(n7997) );
  XOR U7966 ( .A(n8003), .B(n8004), .Z(n7925) );
  AND U7967 ( .A(n8005), .B(n8006), .Z(n8004) );
  XOR U7968 ( .A(n8003), .B(n8007), .Z(n8005) );
  XNOR U7969 ( .A(n8008), .B(n7930), .Z(n7933) );
  XOR U7970 ( .A(n8009), .B(n8010), .Z(n7930) );
  AND U7971 ( .A(n8011), .B(n8012), .Z(n8010) );
  XNOR U7972 ( .A(n8013), .B(n8014), .Z(n8011) );
  IV U7973 ( .A(n8009), .Z(n8013) );
  XNOR U7974 ( .A(n8015), .B(n8016), .Z(n8008) );
  NOR U7975 ( .A(n8017), .B(n8018), .Z(n8016) );
  XNOR U7976 ( .A(n8015), .B(n8019), .Z(n8017) );
  XOR U7977 ( .A(n7939), .B(n7938), .Z(n7929) );
  XNOR U7978 ( .A(n8020), .B(n7935), .Z(n7938) );
  XOR U7979 ( .A(n8021), .B(n8022), .Z(n7935) );
  AND U7980 ( .A(n8023), .B(n8024), .Z(n8022) );
  XNOR U7981 ( .A(n8025), .B(n8026), .Z(n8023) );
  IV U7982 ( .A(n8021), .Z(n8025) );
  XNOR U7983 ( .A(n8027), .B(n8028), .Z(n8020) );
  NOR U7984 ( .A(n8029), .B(n8030), .Z(n8028) );
  XNOR U7985 ( .A(n8027), .B(n8031), .Z(n8029) );
  XOR U7986 ( .A(n8032), .B(n8033), .Z(n7939) );
  NOR U7987 ( .A(n8034), .B(n8035), .Z(n8033) );
  XNOR U7988 ( .A(n8032), .B(n8036), .Z(n8034) );
  XNOR U7989 ( .A(n7831), .B(n7945), .Z(n7947) );
  XNOR U7990 ( .A(n8037), .B(n8038), .Z(n7831) );
  AND U7991 ( .A(n211), .B(n8039), .Z(n8038) );
  XNOR U7992 ( .A(n8040), .B(n8041), .Z(n8039) );
  AND U7993 ( .A(n7837), .B(n7840), .Z(n7945) );
  XOR U7994 ( .A(n8042), .B(n7996), .Z(n7840) );
  XNOR U7995 ( .A(p_input[128]), .B(p_input[512]), .Z(n7996) );
  XNOR U7996 ( .A(n7972), .B(n7971), .Z(n8042) );
  XNOR U7997 ( .A(n8043), .B(n7983), .Z(n7971) );
  XOR U7998 ( .A(n7957), .B(n7955), .Z(n7983) );
  XNOR U7999 ( .A(n8044), .B(n7962), .Z(n7955) );
  XOR U8000 ( .A(p_input[152]), .B(p_input[536]), .Z(n7962) );
  XOR U8001 ( .A(n7952), .B(n7961), .Z(n8044) );
  XOR U8002 ( .A(n8045), .B(n7958), .Z(n7961) );
  XOR U8003 ( .A(p_input[150]), .B(p_input[534]), .Z(n7958) );
  XOR U8004 ( .A(p_input[151]), .B(n6576), .Z(n8045) );
  XOR U8005 ( .A(p_input[146]), .B(p_input[530]), .Z(n7952) );
  XNOR U8006 ( .A(n7967), .B(n7966), .Z(n7957) );
  XOR U8007 ( .A(n8046), .B(n7963), .Z(n7966) );
  XOR U8008 ( .A(p_input[147]), .B(p_input[531]), .Z(n7963) );
  XOR U8009 ( .A(p_input[148]), .B(n6578), .Z(n8046) );
  XOR U8010 ( .A(p_input[149]), .B(p_input[533]), .Z(n7967) );
  XOR U8011 ( .A(n7982), .B(n8047), .Z(n8043) );
  IV U8012 ( .A(n7968), .Z(n8047) );
  XOR U8013 ( .A(p_input[129]), .B(p_input[513]), .Z(n7968) );
  XNOR U8014 ( .A(n8048), .B(n7990), .Z(n7982) );
  XNOR U8015 ( .A(n7978), .B(n7977), .Z(n7990) );
  XNOR U8016 ( .A(n8049), .B(n7974), .Z(n7977) );
  XNOR U8017 ( .A(p_input[154]), .B(p_input[538]), .Z(n7974) );
  XOR U8018 ( .A(p_input[155]), .B(n6582), .Z(n8049) );
  XOR U8019 ( .A(p_input[156]), .B(p_input[540]), .Z(n7978) );
  XOR U8020 ( .A(n7988), .B(n8050), .Z(n8048) );
  IV U8021 ( .A(n7979), .Z(n8050) );
  XOR U8022 ( .A(p_input[145]), .B(p_input[529]), .Z(n7979) );
  XNOR U8023 ( .A(n8051), .B(n7995), .Z(n7988) );
  XNOR U8024 ( .A(p_input[159]), .B(n6585), .Z(n7995) );
  XOR U8025 ( .A(n7985), .B(n7994), .Z(n8051) );
  XOR U8026 ( .A(n8052), .B(n7991), .Z(n7994) );
  XOR U8027 ( .A(p_input[157]), .B(p_input[541]), .Z(n7991) );
  XOR U8028 ( .A(p_input[158]), .B(n6587), .Z(n8052) );
  XOR U8029 ( .A(p_input[153]), .B(p_input[537]), .Z(n7985) );
  XOR U8030 ( .A(n8007), .B(n8006), .Z(n7972) );
  XNOR U8031 ( .A(n8053), .B(n8014), .Z(n8006) );
  XNOR U8032 ( .A(n8002), .B(n8001), .Z(n8014) );
  XNOR U8033 ( .A(n8054), .B(n7998), .Z(n8001) );
  XNOR U8034 ( .A(p_input[139]), .B(p_input[523]), .Z(n7998) );
  XOR U8035 ( .A(p_input[140]), .B(n6590), .Z(n8054) );
  XOR U8036 ( .A(p_input[141]), .B(p_input[525]), .Z(n8002) );
  XOR U8037 ( .A(n8012), .B(n8055), .Z(n8053) );
  IV U8038 ( .A(n8003), .Z(n8055) );
  XOR U8039 ( .A(p_input[130]), .B(p_input[514]), .Z(n8003) );
  XNOR U8040 ( .A(n8056), .B(n8019), .Z(n8012) );
  XNOR U8041 ( .A(p_input[144]), .B(n6593), .Z(n8019) );
  XOR U8042 ( .A(n8009), .B(n8018), .Z(n8056) );
  XOR U8043 ( .A(n8057), .B(n8015), .Z(n8018) );
  XOR U8044 ( .A(p_input[142]), .B(p_input[526]), .Z(n8015) );
  XOR U8045 ( .A(p_input[143]), .B(n6595), .Z(n8057) );
  XOR U8046 ( .A(p_input[138]), .B(p_input[522]), .Z(n8009) );
  XOR U8047 ( .A(n8026), .B(n8024), .Z(n8007) );
  XNOR U8048 ( .A(n8058), .B(n8031), .Z(n8024) );
  XOR U8049 ( .A(p_input[137]), .B(p_input[521]), .Z(n8031) );
  XOR U8050 ( .A(n8021), .B(n8030), .Z(n8058) );
  XOR U8051 ( .A(n8059), .B(n8027), .Z(n8030) );
  XOR U8052 ( .A(p_input[135]), .B(p_input[519]), .Z(n8027) );
  XOR U8053 ( .A(p_input[136]), .B(n6963), .Z(n8059) );
  XOR U8054 ( .A(p_input[131]), .B(p_input[515]), .Z(n8021) );
  XNOR U8055 ( .A(n8036), .B(n8035), .Z(n8026) );
  XOR U8056 ( .A(n8060), .B(n8032), .Z(n8035) );
  XOR U8057 ( .A(p_input[132]), .B(p_input[516]), .Z(n8032) );
  XOR U8058 ( .A(p_input[133]), .B(n6965), .Z(n8060) );
  XOR U8059 ( .A(p_input[134]), .B(p_input[518]), .Z(n8036) );
  XNOR U8060 ( .A(n8061), .B(n8062), .Z(n7837) );
  AND U8061 ( .A(n211), .B(n8063), .Z(n8062) );
  XNOR U8062 ( .A(n8064), .B(n8065), .Z(n211) );
  AND U8063 ( .A(n8066), .B(n8067), .Z(n8065) );
  XOR U8064 ( .A(n7851), .B(n8064), .Z(n8067) );
  XNOR U8065 ( .A(n8068), .B(n8064), .Z(n8066) );
  XOR U8066 ( .A(n8069), .B(n8070), .Z(n8064) );
  AND U8067 ( .A(n8071), .B(n8072), .Z(n8070) );
  XOR U8068 ( .A(n7866), .B(n8069), .Z(n8072) );
  XOR U8069 ( .A(n8069), .B(n7867), .Z(n8071) );
  XOR U8070 ( .A(n8073), .B(n8074), .Z(n8069) );
  AND U8071 ( .A(n8075), .B(n8076), .Z(n8074) );
  XOR U8072 ( .A(n7894), .B(n8073), .Z(n8076) );
  XOR U8073 ( .A(n8073), .B(n7895), .Z(n8075) );
  XOR U8074 ( .A(n8077), .B(n8078), .Z(n8073) );
  AND U8075 ( .A(n8079), .B(n8080), .Z(n8078) );
  XOR U8076 ( .A(n7943), .B(n8077), .Z(n8080) );
  XOR U8077 ( .A(n8077), .B(n7944), .Z(n8079) );
  XOR U8078 ( .A(n8081), .B(n8082), .Z(n8077) );
  AND U8079 ( .A(n8083), .B(n8084), .Z(n8082) );
  XOR U8080 ( .A(n8081), .B(n8040), .Z(n8084) );
  XNOR U8081 ( .A(n8085), .B(n8086), .Z(n7787) );
  AND U8082 ( .A(n215), .B(n8087), .Z(n8086) );
  XNOR U8083 ( .A(n8088), .B(n8089), .Z(n215) );
  AND U8084 ( .A(n8090), .B(n8091), .Z(n8089) );
  XOR U8085 ( .A(n8088), .B(n7797), .Z(n8091) );
  XNOR U8086 ( .A(n8088), .B(n7747), .Z(n8090) );
  XOR U8087 ( .A(n8092), .B(n8093), .Z(n8088) );
  AND U8088 ( .A(n8094), .B(n8095), .Z(n8093) );
  XNOR U8089 ( .A(n7807), .B(n8092), .Z(n8095) );
  XOR U8090 ( .A(n8092), .B(n7757), .Z(n8094) );
  XOR U8091 ( .A(n8096), .B(n8097), .Z(n8092) );
  AND U8092 ( .A(n8098), .B(n8099), .Z(n8097) );
  XNOR U8093 ( .A(n7817), .B(n8096), .Z(n8099) );
  XOR U8094 ( .A(n8096), .B(n7766), .Z(n8098) );
  XOR U8095 ( .A(n8100), .B(n8101), .Z(n8096) );
  AND U8096 ( .A(n8102), .B(n8103), .Z(n8101) );
  XOR U8097 ( .A(n8100), .B(n7774), .Z(n8102) );
  XOR U8098 ( .A(n8104), .B(n8105), .Z(n7738) );
  AND U8099 ( .A(n219), .B(n8087), .Z(n8105) );
  XNOR U8100 ( .A(n8085), .B(n8104), .Z(n8087) );
  XNOR U8101 ( .A(n8106), .B(n8107), .Z(n219) );
  AND U8102 ( .A(n8108), .B(n8109), .Z(n8107) );
  XNOR U8103 ( .A(n8110), .B(n8106), .Z(n8109) );
  IV U8104 ( .A(n7797), .Z(n8110) );
  XOR U8105 ( .A(n8068), .B(n8111), .Z(n7797) );
  AND U8106 ( .A(n222), .B(n8112), .Z(n8111) );
  XOR U8107 ( .A(n7850), .B(n7847), .Z(n8112) );
  IV U8108 ( .A(n8068), .Z(n7850) );
  XNOR U8109 ( .A(n7747), .B(n8106), .Z(n8108) );
  XOR U8110 ( .A(n8113), .B(n8114), .Z(n7747) );
  AND U8111 ( .A(n238), .B(n8115), .Z(n8114) );
  XOR U8112 ( .A(n8116), .B(n8117), .Z(n8106) );
  AND U8113 ( .A(n8118), .B(n8119), .Z(n8117) );
  XNOR U8114 ( .A(n8116), .B(n7807), .Z(n8119) );
  XOR U8115 ( .A(n7867), .B(n8120), .Z(n7807) );
  AND U8116 ( .A(n222), .B(n8121), .Z(n8120) );
  XOR U8117 ( .A(n7863), .B(n7867), .Z(n8121) );
  XNOR U8118 ( .A(n8122), .B(n8116), .Z(n8118) );
  IV U8119 ( .A(n7757), .Z(n8122) );
  XOR U8120 ( .A(n8123), .B(n8124), .Z(n7757) );
  AND U8121 ( .A(n238), .B(n8125), .Z(n8124) );
  XOR U8122 ( .A(n8126), .B(n8127), .Z(n8116) );
  AND U8123 ( .A(n8128), .B(n8129), .Z(n8127) );
  XNOR U8124 ( .A(n8126), .B(n7817), .Z(n8129) );
  XOR U8125 ( .A(n7895), .B(n8130), .Z(n7817) );
  AND U8126 ( .A(n222), .B(n8131), .Z(n8130) );
  XOR U8127 ( .A(n7891), .B(n7895), .Z(n8131) );
  XOR U8128 ( .A(n7766), .B(n8126), .Z(n8128) );
  XOR U8129 ( .A(n8132), .B(n8133), .Z(n7766) );
  AND U8130 ( .A(n238), .B(n8134), .Z(n8133) );
  XOR U8131 ( .A(n8100), .B(n8135), .Z(n8126) );
  AND U8132 ( .A(n8136), .B(n8103), .Z(n8135) );
  XNOR U8133 ( .A(n7827), .B(n8100), .Z(n8103) );
  XOR U8134 ( .A(n7944), .B(n8137), .Z(n7827) );
  AND U8135 ( .A(n222), .B(n8138), .Z(n8137) );
  XOR U8136 ( .A(n7940), .B(n7944), .Z(n8138) );
  XNOR U8137 ( .A(n8139), .B(n8100), .Z(n8136) );
  IV U8138 ( .A(n7774), .Z(n8139) );
  XOR U8139 ( .A(n8140), .B(n8141), .Z(n7774) );
  AND U8140 ( .A(n238), .B(n8142), .Z(n8141) );
  XOR U8141 ( .A(n8143), .B(n8144), .Z(n8100) );
  AND U8142 ( .A(n8145), .B(n8146), .Z(n8144) );
  XNOR U8143 ( .A(n8143), .B(n7835), .Z(n8146) );
  XOR U8144 ( .A(n8041), .B(n8147), .Z(n7835) );
  AND U8145 ( .A(n222), .B(n8148), .Z(n8147) );
  XOR U8146 ( .A(n8037), .B(n8041), .Z(n8148) );
  XNOR U8147 ( .A(n8149), .B(n8143), .Z(n8145) );
  IV U8148 ( .A(n7784), .Z(n8149) );
  XOR U8149 ( .A(n8150), .B(n8151), .Z(n7784) );
  AND U8150 ( .A(n238), .B(n8152), .Z(n8151) );
  AND U8151 ( .A(n8104), .B(n8085), .Z(n8143) );
  XNOR U8152 ( .A(n8153), .B(n8154), .Z(n8085) );
  AND U8153 ( .A(n222), .B(n8063), .Z(n8154) );
  XNOR U8154 ( .A(n8061), .B(n8153), .Z(n8063) );
  XNOR U8155 ( .A(n8155), .B(n8156), .Z(n222) );
  AND U8156 ( .A(n8157), .B(n8158), .Z(n8156) );
  XNOR U8157 ( .A(n8155), .B(n7847), .Z(n8158) );
  IV U8158 ( .A(n7851), .Z(n7847) );
  XOR U8159 ( .A(n8159), .B(n8160), .Z(n7851) );
  AND U8160 ( .A(n226), .B(n8161), .Z(n8160) );
  XOR U8161 ( .A(n8162), .B(n8159), .Z(n8161) );
  XNOR U8162 ( .A(n8155), .B(n8068), .Z(n8157) );
  XOR U8163 ( .A(n8163), .B(n8164), .Z(n8068) );
  AND U8164 ( .A(n234), .B(n8115), .Z(n8164) );
  XOR U8165 ( .A(n8113), .B(n8163), .Z(n8115) );
  XOR U8166 ( .A(n8165), .B(n8166), .Z(n8155) );
  AND U8167 ( .A(n8167), .B(n8168), .Z(n8166) );
  XNOR U8168 ( .A(n8165), .B(n7863), .Z(n8168) );
  IV U8169 ( .A(n7866), .Z(n7863) );
  XOR U8170 ( .A(n8169), .B(n8170), .Z(n7866) );
  AND U8171 ( .A(n226), .B(n8171), .Z(n8170) );
  XOR U8172 ( .A(n8172), .B(n8169), .Z(n8171) );
  XOR U8173 ( .A(n7867), .B(n8165), .Z(n8167) );
  XOR U8174 ( .A(n8173), .B(n8174), .Z(n7867) );
  AND U8175 ( .A(n234), .B(n8125), .Z(n8174) );
  XOR U8176 ( .A(n8173), .B(n8123), .Z(n8125) );
  XOR U8177 ( .A(n8175), .B(n8176), .Z(n8165) );
  AND U8178 ( .A(n8177), .B(n8178), .Z(n8176) );
  XNOR U8179 ( .A(n8175), .B(n7891), .Z(n8178) );
  IV U8180 ( .A(n7894), .Z(n7891) );
  XOR U8181 ( .A(n8179), .B(n8180), .Z(n7894) );
  AND U8182 ( .A(n226), .B(n8181), .Z(n8180) );
  XNOR U8183 ( .A(n8182), .B(n8179), .Z(n8181) );
  XOR U8184 ( .A(n7895), .B(n8175), .Z(n8177) );
  XOR U8185 ( .A(n8183), .B(n8184), .Z(n7895) );
  AND U8186 ( .A(n234), .B(n8134), .Z(n8184) );
  XOR U8187 ( .A(n8183), .B(n8132), .Z(n8134) );
  XOR U8188 ( .A(n8185), .B(n8186), .Z(n8175) );
  AND U8189 ( .A(n8187), .B(n8188), .Z(n8186) );
  XNOR U8190 ( .A(n8185), .B(n7940), .Z(n8188) );
  IV U8191 ( .A(n7943), .Z(n7940) );
  XOR U8192 ( .A(n8189), .B(n8190), .Z(n7943) );
  AND U8193 ( .A(n226), .B(n8191), .Z(n8190) );
  XOR U8194 ( .A(n8192), .B(n8189), .Z(n8191) );
  XOR U8195 ( .A(n7944), .B(n8185), .Z(n8187) );
  XOR U8196 ( .A(n8193), .B(n8194), .Z(n7944) );
  AND U8197 ( .A(n234), .B(n8142), .Z(n8194) );
  XOR U8198 ( .A(n8193), .B(n8140), .Z(n8142) );
  XOR U8199 ( .A(n8081), .B(n8195), .Z(n8185) );
  AND U8200 ( .A(n8083), .B(n8196), .Z(n8195) );
  XNOR U8201 ( .A(n8081), .B(n8037), .Z(n8196) );
  IV U8202 ( .A(n8040), .Z(n8037) );
  XOR U8203 ( .A(n8197), .B(n8198), .Z(n8040) );
  AND U8204 ( .A(n226), .B(n8199), .Z(n8198) );
  XNOR U8205 ( .A(n8200), .B(n8197), .Z(n8199) );
  XOR U8206 ( .A(n8041), .B(n8081), .Z(n8083) );
  XOR U8207 ( .A(n8201), .B(n8202), .Z(n8041) );
  AND U8208 ( .A(n234), .B(n8152), .Z(n8202) );
  XOR U8209 ( .A(n8201), .B(n8150), .Z(n8152) );
  AND U8210 ( .A(n8153), .B(n8061), .Z(n8081) );
  XNOR U8211 ( .A(n8203), .B(n8204), .Z(n8061) );
  AND U8212 ( .A(n226), .B(n8205), .Z(n8204) );
  XNOR U8213 ( .A(n8206), .B(n8203), .Z(n8205) );
  XNOR U8214 ( .A(n8207), .B(n8208), .Z(n226) );
  AND U8215 ( .A(n8209), .B(n8210), .Z(n8208) );
  XOR U8216 ( .A(n8162), .B(n8207), .Z(n8210) );
  AND U8217 ( .A(n8211), .B(n8212), .Z(n8162) );
  XNOR U8218 ( .A(n8159), .B(n8207), .Z(n8209) );
  XNOR U8219 ( .A(n8213), .B(n8214), .Z(n8159) );
  AND U8220 ( .A(n230), .B(n8215), .Z(n8214) );
  XNOR U8221 ( .A(n8216), .B(n8217), .Z(n8215) );
  XOR U8222 ( .A(n8218), .B(n8219), .Z(n8207) );
  AND U8223 ( .A(n8220), .B(n8221), .Z(n8219) );
  XNOR U8224 ( .A(n8218), .B(n8211), .Z(n8221) );
  IV U8225 ( .A(n8172), .Z(n8211) );
  XOR U8226 ( .A(n8222), .B(n8223), .Z(n8172) );
  XOR U8227 ( .A(n8224), .B(n8212), .Z(n8223) );
  AND U8228 ( .A(n8182), .B(n8225), .Z(n8212) );
  AND U8229 ( .A(n8226), .B(n8227), .Z(n8224) );
  XOR U8230 ( .A(n8228), .B(n8222), .Z(n8226) );
  XNOR U8231 ( .A(n8169), .B(n8218), .Z(n8220) );
  XNOR U8232 ( .A(n8229), .B(n8230), .Z(n8169) );
  AND U8233 ( .A(n230), .B(n8231), .Z(n8230) );
  XNOR U8234 ( .A(n8232), .B(n8233), .Z(n8231) );
  XOR U8235 ( .A(n8234), .B(n8235), .Z(n8218) );
  AND U8236 ( .A(n8236), .B(n8237), .Z(n8235) );
  XNOR U8237 ( .A(n8234), .B(n8182), .Z(n8237) );
  XOR U8238 ( .A(n8238), .B(n8227), .Z(n8182) );
  XNOR U8239 ( .A(n8239), .B(n8222), .Z(n8227) );
  XOR U8240 ( .A(n8240), .B(n8241), .Z(n8222) );
  AND U8241 ( .A(n8242), .B(n8243), .Z(n8241) );
  XOR U8242 ( .A(n8244), .B(n8240), .Z(n8242) );
  XNOR U8243 ( .A(n8245), .B(n8246), .Z(n8239) );
  AND U8244 ( .A(n8247), .B(n8248), .Z(n8246) );
  XOR U8245 ( .A(n8245), .B(n8249), .Z(n8247) );
  XNOR U8246 ( .A(n8228), .B(n8225), .Z(n8238) );
  AND U8247 ( .A(n8250), .B(n8251), .Z(n8225) );
  XOR U8248 ( .A(n8252), .B(n8253), .Z(n8228) );
  AND U8249 ( .A(n8254), .B(n8255), .Z(n8253) );
  XOR U8250 ( .A(n8252), .B(n8256), .Z(n8254) );
  XNOR U8251 ( .A(n8179), .B(n8234), .Z(n8236) );
  XNOR U8252 ( .A(n8257), .B(n8258), .Z(n8179) );
  AND U8253 ( .A(n230), .B(n8259), .Z(n8258) );
  XNOR U8254 ( .A(n8260), .B(n8261), .Z(n8259) );
  XOR U8255 ( .A(n8262), .B(n8263), .Z(n8234) );
  AND U8256 ( .A(n8264), .B(n8265), .Z(n8263) );
  XNOR U8257 ( .A(n8262), .B(n8250), .Z(n8265) );
  IV U8258 ( .A(n8192), .Z(n8250) );
  XNOR U8259 ( .A(n8266), .B(n8243), .Z(n8192) );
  XNOR U8260 ( .A(n8267), .B(n8249), .Z(n8243) );
  XOR U8261 ( .A(n8268), .B(n8269), .Z(n8249) );
  AND U8262 ( .A(n8270), .B(n8271), .Z(n8269) );
  XOR U8263 ( .A(n8268), .B(n8272), .Z(n8270) );
  XNOR U8264 ( .A(n8248), .B(n8240), .Z(n8267) );
  XOR U8265 ( .A(n8273), .B(n8274), .Z(n8240) );
  AND U8266 ( .A(n8275), .B(n8276), .Z(n8274) );
  XNOR U8267 ( .A(n8277), .B(n8273), .Z(n8275) );
  XNOR U8268 ( .A(n8278), .B(n8245), .Z(n8248) );
  XOR U8269 ( .A(n8279), .B(n8280), .Z(n8245) );
  AND U8270 ( .A(n8281), .B(n8282), .Z(n8280) );
  XOR U8271 ( .A(n8279), .B(n8283), .Z(n8281) );
  XNOR U8272 ( .A(n8284), .B(n8285), .Z(n8278) );
  AND U8273 ( .A(n8286), .B(n8287), .Z(n8285) );
  XNOR U8274 ( .A(n8284), .B(n8288), .Z(n8286) );
  XNOR U8275 ( .A(n8244), .B(n8251), .Z(n8266) );
  AND U8276 ( .A(n8200), .B(n8289), .Z(n8251) );
  XOR U8277 ( .A(n8256), .B(n8255), .Z(n8244) );
  XNOR U8278 ( .A(n8290), .B(n8252), .Z(n8255) );
  XOR U8279 ( .A(n8291), .B(n8292), .Z(n8252) );
  AND U8280 ( .A(n8293), .B(n8294), .Z(n8292) );
  XOR U8281 ( .A(n8291), .B(n8295), .Z(n8293) );
  XNOR U8282 ( .A(n8296), .B(n8297), .Z(n8290) );
  AND U8283 ( .A(n8298), .B(n8299), .Z(n8297) );
  XOR U8284 ( .A(n8296), .B(n8300), .Z(n8298) );
  XOR U8285 ( .A(n8301), .B(n8302), .Z(n8256) );
  AND U8286 ( .A(n8303), .B(n8304), .Z(n8302) );
  XOR U8287 ( .A(n8301), .B(n8305), .Z(n8303) );
  XNOR U8288 ( .A(n8189), .B(n8262), .Z(n8264) );
  XNOR U8289 ( .A(n8306), .B(n8307), .Z(n8189) );
  AND U8290 ( .A(n230), .B(n8308), .Z(n8307) );
  XNOR U8291 ( .A(n8309), .B(n8310), .Z(n8308) );
  XOR U8292 ( .A(n8311), .B(n8312), .Z(n8262) );
  AND U8293 ( .A(n8313), .B(n8314), .Z(n8312) );
  XNOR U8294 ( .A(n8311), .B(n8200), .Z(n8314) );
  XOR U8295 ( .A(n8315), .B(n8276), .Z(n8200) );
  XNOR U8296 ( .A(n8316), .B(n8283), .Z(n8276) );
  XOR U8297 ( .A(n8272), .B(n8271), .Z(n8283) );
  XNOR U8298 ( .A(n8317), .B(n8268), .Z(n8271) );
  XOR U8299 ( .A(n8318), .B(n8319), .Z(n8268) );
  AND U8300 ( .A(n8320), .B(n8321), .Z(n8319) );
  XNOR U8301 ( .A(n8322), .B(n8323), .Z(n8320) );
  IV U8302 ( .A(n8318), .Z(n8322) );
  XNOR U8303 ( .A(n8324), .B(n8325), .Z(n8317) );
  NOR U8304 ( .A(n8326), .B(n8327), .Z(n8325) );
  XNOR U8305 ( .A(n8324), .B(n8328), .Z(n8326) );
  XOR U8306 ( .A(n8329), .B(n8330), .Z(n8272) );
  NOR U8307 ( .A(n8331), .B(n8332), .Z(n8330) );
  XNOR U8308 ( .A(n8329), .B(n8333), .Z(n8331) );
  XNOR U8309 ( .A(n8282), .B(n8273), .Z(n8316) );
  XOR U8310 ( .A(n8334), .B(n8335), .Z(n8273) );
  AND U8311 ( .A(n8336), .B(n8337), .Z(n8335) );
  XOR U8312 ( .A(n8334), .B(n8338), .Z(n8336) );
  XOR U8313 ( .A(n8339), .B(n8288), .Z(n8282) );
  XOR U8314 ( .A(n8340), .B(n8341), .Z(n8288) );
  NOR U8315 ( .A(n8342), .B(n8343), .Z(n8341) );
  XOR U8316 ( .A(n8340), .B(n8344), .Z(n8342) );
  XNOR U8317 ( .A(n8287), .B(n8279), .Z(n8339) );
  XOR U8318 ( .A(n8345), .B(n8346), .Z(n8279) );
  AND U8319 ( .A(n8347), .B(n8348), .Z(n8346) );
  XOR U8320 ( .A(n8345), .B(n8349), .Z(n8347) );
  XNOR U8321 ( .A(n8350), .B(n8284), .Z(n8287) );
  XOR U8322 ( .A(n8351), .B(n8352), .Z(n8284) );
  AND U8323 ( .A(n8353), .B(n8354), .Z(n8352) );
  XNOR U8324 ( .A(n8355), .B(n8356), .Z(n8353) );
  IV U8325 ( .A(n8351), .Z(n8355) );
  XNOR U8326 ( .A(n8357), .B(n8358), .Z(n8350) );
  NOR U8327 ( .A(n8359), .B(n8360), .Z(n8358) );
  XNOR U8328 ( .A(n8357), .B(n8361), .Z(n8359) );
  XOR U8329 ( .A(n8277), .B(n8289), .Z(n8315) );
  NOR U8330 ( .A(n8206), .B(n8362), .Z(n8289) );
  XNOR U8331 ( .A(n8295), .B(n8294), .Z(n8277) );
  XNOR U8332 ( .A(n8363), .B(n8300), .Z(n8294) );
  XNOR U8333 ( .A(n8364), .B(n8365), .Z(n8300) );
  NOR U8334 ( .A(n8366), .B(n8367), .Z(n8365) );
  XOR U8335 ( .A(n8364), .B(n8368), .Z(n8366) );
  XNOR U8336 ( .A(n8299), .B(n8291), .Z(n8363) );
  XOR U8337 ( .A(n8369), .B(n8370), .Z(n8291) );
  AND U8338 ( .A(n8371), .B(n8372), .Z(n8370) );
  XOR U8339 ( .A(n8369), .B(n8373), .Z(n8371) );
  XNOR U8340 ( .A(n8374), .B(n8296), .Z(n8299) );
  XOR U8341 ( .A(n8375), .B(n8376), .Z(n8296) );
  AND U8342 ( .A(n8377), .B(n8378), .Z(n8376) );
  XNOR U8343 ( .A(n8379), .B(n8380), .Z(n8377) );
  IV U8344 ( .A(n8375), .Z(n8379) );
  XNOR U8345 ( .A(n8381), .B(n8382), .Z(n8374) );
  NOR U8346 ( .A(n8383), .B(n8384), .Z(n8382) );
  XNOR U8347 ( .A(n8381), .B(n8385), .Z(n8383) );
  XOR U8348 ( .A(n8305), .B(n8304), .Z(n8295) );
  XNOR U8349 ( .A(n8386), .B(n8301), .Z(n8304) );
  XOR U8350 ( .A(n8387), .B(n8388), .Z(n8301) );
  AND U8351 ( .A(n8389), .B(n8390), .Z(n8388) );
  XNOR U8352 ( .A(n8391), .B(n8392), .Z(n8389) );
  IV U8353 ( .A(n8387), .Z(n8391) );
  XNOR U8354 ( .A(n8393), .B(n8394), .Z(n8386) );
  NOR U8355 ( .A(n8395), .B(n8396), .Z(n8394) );
  XNOR U8356 ( .A(n8393), .B(n8397), .Z(n8395) );
  XOR U8357 ( .A(n8398), .B(n8399), .Z(n8305) );
  NOR U8358 ( .A(n8400), .B(n8401), .Z(n8399) );
  XNOR U8359 ( .A(n8398), .B(n8402), .Z(n8400) );
  XNOR U8360 ( .A(n8197), .B(n8311), .Z(n8313) );
  XNOR U8361 ( .A(n8403), .B(n8404), .Z(n8197) );
  AND U8362 ( .A(n230), .B(n8405), .Z(n8404) );
  XNOR U8363 ( .A(n8406), .B(n8407), .Z(n8405) );
  AND U8364 ( .A(n8203), .B(n8206), .Z(n8311) );
  XOR U8365 ( .A(n8408), .B(n8362), .Z(n8206) );
  XNOR U8366 ( .A(p_input[160]), .B(p_input[512]), .Z(n8362) );
  XNOR U8367 ( .A(n8338), .B(n8337), .Z(n8408) );
  XNOR U8368 ( .A(n8409), .B(n8349), .Z(n8337) );
  XOR U8369 ( .A(n8323), .B(n8321), .Z(n8349) );
  XNOR U8370 ( .A(n8410), .B(n8328), .Z(n8321) );
  XOR U8371 ( .A(p_input[184]), .B(p_input[536]), .Z(n8328) );
  XOR U8372 ( .A(n8318), .B(n8327), .Z(n8410) );
  XOR U8373 ( .A(n8411), .B(n8324), .Z(n8327) );
  XOR U8374 ( .A(p_input[182]), .B(p_input[534]), .Z(n8324) );
  XOR U8375 ( .A(p_input[183]), .B(n6576), .Z(n8411) );
  XOR U8376 ( .A(p_input[178]), .B(p_input[530]), .Z(n8318) );
  XNOR U8377 ( .A(n8333), .B(n8332), .Z(n8323) );
  XOR U8378 ( .A(n8412), .B(n8329), .Z(n8332) );
  XOR U8379 ( .A(p_input[179]), .B(p_input[531]), .Z(n8329) );
  XOR U8380 ( .A(p_input[180]), .B(n6578), .Z(n8412) );
  XOR U8381 ( .A(p_input[181]), .B(p_input[533]), .Z(n8333) );
  XOR U8382 ( .A(n8348), .B(n8413), .Z(n8409) );
  IV U8383 ( .A(n8334), .Z(n8413) );
  XOR U8384 ( .A(p_input[161]), .B(p_input[513]), .Z(n8334) );
  XNOR U8385 ( .A(n8414), .B(n8356), .Z(n8348) );
  XNOR U8386 ( .A(n8344), .B(n8343), .Z(n8356) );
  XNOR U8387 ( .A(n8415), .B(n8340), .Z(n8343) );
  XNOR U8388 ( .A(p_input[186]), .B(p_input[538]), .Z(n8340) );
  XOR U8389 ( .A(p_input[187]), .B(n6582), .Z(n8415) );
  XOR U8390 ( .A(p_input[188]), .B(p_input[540]), .Z(n8344) );
  XOR U8391 ( .A(n8354), .B(n8416), .Z(n8414) );
  IV U8392 ( .A(n8345), .Z(n8416) );
  XOR U8393 ( .A(p_input[177]), .B(p_input[529]), .Z(n8345) );
  XNOR U8394 ( .A(n8417), .B(n8361), .Z(n8354) );
  XNOR U8395 ( .A(p_input[191]), .B(n6585), .Z(n8361) );
  XOR U8396 ( .A(n8351), .B(n8360), .Z(n8417) );
  XOR U8397 ( .A(n8418), .B(n8357), .Z(n8360) );
  XOR U8398 ( .A(p_input[189]), .B(p_input[541]), .Z(n8357) );
  XOR U8399 ( .A(p_input[190]), .B(n6587), .Z(n8418) );
  XOR U8400 ( .A(p_input[185]), .B(p_input[537]), .Z(n8351) );
  XOR U8401 ( .A(n8373), .B(n8372), .Z(n8338) );
  XNOR U8402 ( .A(n8419), .B(n8380), .Z(n8372) );
  XNOR U8403 ( .A(n8368), .B(n8367), .Z(n8380) );
  XNOR U8404 ( .A(n8420), .B(n8364), .Z(n8367) );
  XNOR U8405 ( .A(p_input[171]), .B(p_input[523]), .Z(n8364) );
  XOR U8406 ( .A(p_input[172]), .B(n6590), .Z(n8420) );
  XOR U8407 ( .A(p_input[173]), .B(p_input[525]), .Z(n8368) );
  XOR U8408 ( .A(n8378), .B(n8421), .Z(n8419) );
  IV U8409 ( .A(n8369), .Z(n8421) );
  XOR U8410 ( .A(p_input[162]), .B(p_input[514]), .Z(n8369) );
  XNOR U8411 ( .A(n8422), .B(n8385), .Z(n8378) );
  XNOR U8412 ( .A(p_input[176]), .B(n6593), .Z(n8385) );
  XOR U8413 ( .A(n8375), .B(n8384), .Z(n8422) );
  XOR U8414 ( .A(n8423), .B(n8381), .Z(n8384) );
  XOR U8415 ( .A(p_input[174]), .B(p_input[526]), .Z(n8381) );
  XOR U8416 ( .A(p_input[175]), .B(n6595), .Z(n8423) );
  XOR U8417 ( .A(p_input[170]), .B(p_input[522]), .Z(n8375) );
  XOR U8418 ( .A(n8392), .B(n8390), .Z(n8373) );
  XNOR U8419 ( .A(n8424), .B(n8397), .Z(n8390) );
  XOR U8420 ( .A(p_input[169]), .B(p_input[521]), .Z(n8397) );
  XOR U8421 ( .A(n8387), .B(n8396), .Z(n8424) );
  XOR U8422 ( .A(n8425), .B(n8393), .Z(n8396) );
  XOR U8423 ( .A(p_input[167]), .B(p_input[519]), .Z(n8393) );
  XOR U8424 ( .A(p_input[168]), .B(n6963), .Z(n8425) );
  XOR U8425 ( .A(p_input[163]), .B(p_input[515]), .Z(n8387) );
  XNOR U8426 ( .A(n8402), .B(n8401), .Z(n8392) );
  XOR U8427 ( .A(n8426), .B(n8398), .Z(n8401) );
  XOR U8428 ( .A(p_input[164]), .B(p_input[516]), .Z(n8398) );
  XOR U8429 ( .A(p_input[165]), .B(n6965), .Z(n8426) );
  XOR U8430 ( .A(p_input[166]), .B(p_input[518]), .Z(n8402) );
  XNOR U8431 ( .A(n8427), .B(n8428), .Z(n8203) );
  AND U8432 ( .A(n230), .B(n8429), .Z(n8428) );
  XNOR U8433 ( .A(n8430), .B(n8431), .Z(n230) );
  AND U8434 ( .A(n8432), .B(n8433), .Z(n8431) );
  XOR U8435 ( .A(n8217), .B(n8430), .Z(n8433) );
  XNOR U8436 ( .A(n8434), .B(n8430), .Z(n8432) );
  XOR U8437 ( .A(n8435), .B(n8436), .Z(n8430) );
  AND U8438 ( .A(n8437), .B(n8438), .Z(n8436) );
  XOR U8439 ( .A(n8232), .B(n8435), .Z(n8438) );
  XOR U8440 ( .A(n8435), .B(n8233), .Z(n8437) );
  XOR U8441 ( .A(n8439), .B(n8440), .Z(n8435) );
  AND U8442 ( .A(n8441), .B(n8442), .Z(n8440) );
  XOR U8443 ( .A(n8260), .B(n8439), .Z(n8442) );
  XOR U8444 ( .A(n8439), .B(n8261), .Z(n8441) );
  XOR U8445 ( .A(n8443), .B(n8444), .Z(n8439) );
  AND U8446 ( .A(n8445), .B(n8446), .Z(n8444) );
  XOR U8447 ( .A(n8309), .B(n8443), .Z(n8446) );
  XOR U8448 ( .A(n8443), .B(n8310), .Z(n8445) );
  XOR U8449 ( .A(n8447), .B(n8448), .Z(n8443) );
  AND U8450 ( .A(n8449), .B(n8450), .Z(n8448) );
  XOR U8451 ( .A(n8447), .B(n8406), .Z(n8450) );
  XNOR U8452 ( .A(n8451), .B(n8452), .Z(n8153) );
  AND U8453 ( .A(n234), .B(n8453), .Z(n8452) );
  XNOR U8454 ( .A(n8454), .B(n8455), .Z(n234) );
  AND U8455 ( .A(n8456), .B(n8457), .Z(n8455) );
  XOR U8456 ( .A(n8454), .B(n8163), .Z(n8457) );
  XNOR U8457 ( .A(n8454), .B(n8113), .Z(n8456) );
  XOR U8458 ( .A(n8458), .B(n8459), .Z(n8454) );
  AND U8459 ( .A(n8460), .B(n8461), .Z(n8459) );
  XNOR U8460 ( .A(n8173), .B(n8458), .Z(n8461) );
  XOR U8461 ( .A(n8458), .B(n8123), .Z(n8460) );
  XOR U8462 ( .A(n8462), .B(n8463), .Z(n8458) );
  AND U8463 ( .A(n8464), .B(n8465), .Z(n8463) );
  XNOR U8464 ( .A(n8183), .B(n8462), .Z(n8465) );
  XOR U8465 ( .A(n8462), .B(n8132), .Z(n8464) );
  XOR U8466 ( .A(n8466), .B(n8467), .Z(n8462) );
  AND U8467 ( .A(n8468), .B(n8469), .Z(n8467) );
  XOR U8468 ( .A(n8466), .B(n8140), .Z(n8468) );
  XOR U8469 ( .A(n8470), .B(n8471), .Z(n8104) );
  AND U8470 ( .A(n238), .B(n8453), .Z(n8471) );
  XNOR U8471 ( .A(n8451), .B(n8470), .Z(n8453) );
  XNOR U8472 ( .A(n8472), .B(n8473), .Z(n238) );
  AND U8473 ( .A(n8474), .B(n8475), .Z(n8473) );
  XNOR U8474 ( .A(n8476), .B(n8472), .Z(n8475) );
  IV U8475 ( .A(n8163), .Z(n8476) );
  XOR U8476 ( .A(n8434), .B(n8477), .Z(n8163) );
  AND U8477 ( .A(n241), .B(n8478), .Z(n8477) );
  XOR U8478 ( .A(n8216), .B(n8213), .Z(n8478) );
  IV U8479 ( .A(n8434), .Z(n8216) );
  XNOR U8480 ( .A(n8113), .B(n8472), .Z(n8474) );
  XOR U8481 ( .A(n8479), .B(n8480), .Z(n8113) );
  AND U8482 ( .A(n257), .B(n8481), .Z(n8480) );
  XOR U8483 ( .A(n8482), .B(n8483), .Z(n8472) );
  AND U8484 ( .A(n8484), .B(n8485), .Z(n8483) );
  XNOR U8485 ( .A(n8482), .B(n8173), .Z(n8485) );
  XOR U8486 ( .A(n8233), .B(n8486), .Z(n8173) );
  AND U8487 ( .A(n241), .B(n8487), .Z(n8486) );
  XOR U8488 ( .A(n8229), .B(n8233), .Z(n8487) );
  XNOR U8489 ( .A(n8488), .B(n8482), .Z(n8484) );
  IV U8490 ( .A(n8123), .Z(n8488) );
  XOR U8491 ( .A(n8489), .B(n8490), .Z(n8123) );
  AND U8492 ( .A(n257), .B(n8491), .Z(n8490) );
  XOR U8493 ( .A(n8492), .B(n8493), .Z(n8482) );
  AND U8494 ( .A(n8494), .B(n8495), .Z(n8493) );
  XNOR U8495 ( .A(n8492), .B(n8183), .Z(n8495) );
  XOR U8496 ( .A(n8261), .B(n8496), .Z(n8183) );
  AND U8497 ( .A(n241), .B(n8497), .Z(n8496) );
  XOR U8498 ( .A(n8257), .B(n8261), .Z(n8497) );
  XOR U8499 ( .A(n8132), .B(n8492), .Z(n8494) );
  XOR U8500 ( .A(n8498), .B(n8499), .Z(n8132) );
  AND U8501 ( .A(n257), .B(n8500), .Z(n8499) );
  XOR U8502 ( .A(n8466), .B(n8501), .Z(n8492) );
  AND U8503 ( .A(n8502), .B(n8469), .Z(n8501) );
  XNOR U8504 ( .A(n8193), .B(n8466), .Z(n8469) );
  XOR U8505 ( .A(n8310), .B(n8503), .Z(n8193) );
  AND U8506 ( .A(n241), .B(n8504), .Z(n8503) );
  XOR U8507 ( .A(n8306), .B(n8310), .Z(n8504) );
  XNOR U8508 ( .A(n8505), .B(n8466), .Z(n8502) );
  IV U8509 ( .A(n8140), .Z(n8505) );
  XOR U8510 ( .A(n8506), .B(n8507), .Z(n8140) );
  AND U8511 ( .A(n257), .B(n8508), .Z(n8507) );
  XOR U8512 ( .A(n8509), .B(n8510), .Z(n8466) );
  AND U8513 ( .A(n8511), .B(n8512), .Z(n8510) );
  XNOR U8514 ( .A(n8509), .B(n8201), .Z(n8512) );
  XOR U8515 ( .A(n8407), .B(n8513), .Z(n8201) );
  AND U8516 ( .A(n241), .B(n8514), .Z(n8513) );
  XOR U8517 ( .A(n8403), .B(n8407), .Z(n8514) );
  XNOR U8518 ( .A(n8515), .B(n8509), .Z(n8511) );
  IV U8519 ( .A(n8150), .Z(n8515) );
  XOR U8520 ( .A(n8516), .B(n8517), .Z(n8150) );
  AND U8521 ( .A(n257), .B(n8518), .Z(n8517) );
  AND U8522 ( .A(n8470), .B(n8451), .Z(n8509) );
  XNOR U8523 ( .A(n8519), .B(n8520), .Z(n8451) );
  AND U8524 ( .A(n241), .B(n8429), .Z(n8520) );
  XNOR U8525 ( .A(n8427), .B(n8519), .Z(n8429) );
  XNOR U8526 ( .A(n8521), .B(n8522), .Z(n241) );
  AND U8527 ( .A(n8523), .B(n8524), .Z(n8522) );
  XNOR U8528 ( .A(n8521), .B(n8213), .Z(n8524) );
  IV U8529 ( .A(n8217), .Z(n8213) );
  XOR U8530 ( .A(n8525), .B(n8526), .Z(n8217) );
  AND U8531 ( .A(n245), .B(n8527), .Z(n8526) );
  XOR U8532 ( .A(n8528), .B(n8525), .Z(n8527) );
  XNOR U8533 ( .A(n8521), .B(n8434), .Z(n8523) );
  XOR U8534 ( .A(n8529), .B(n8530), .Z(n8434) );
  AND U8535 ( .A(n253), .B(n8481), .Z(n8530) );
  XOR U8536 ( .A(n8479), .B(n8529), .Z(n8481) );
  XOR U8537 ( .A(n8531), .B(n8532), .Z(n8521) );
  AND U8538 ( .A(n8533), .B(n8534), .Z(n8532) );
  XNOR U8539 ( .A(n8531), .B(n8229), .Z(n8534) );
  IV U8540 ( .A(n8232), .Z(n8229) );
  XOR U8541 ( .A(n8535), .B(n8536), .Z(n8232) );
  AND U8542 ( .A(n245), .B(n8537), .Z(n8536) );
  XOR U8543 ( .A(n8538), .B(n8535), .Z(n8537) );
  XOR U8544 ( .A(n8233), .B(n8531), .Z(n8533) );
  XOR U8545 ( .A(n8539), .B(n8540), .Z(n8233) );
  AND U8546 ( .A(n253), .B(n8491), .Z(n8540) );
  XOR U8547 ( .A(n8539), .B(n8489), .Z(n8491) );
  XOR U8548 ( .A(n8541), .B(n8542), .Z(n8531) );
  AND U8549 ( .A(n8543), .B(n8544), .Z(n8542) );
  XNOR U8550 ( .A(n8541), .B(n8257), .Z(n8544) );
  IV U8551 ( .A(n8260), .Z(n8257) );
  XOR U8552 ( .A(n8545), .B(n8546), .Z(n8260) );
  AND U8553 ( .A(n245), .B(n8547), .Z(n8546) );
  XNOR U8554 ( .A(n8548), .B(n8545), .Z(n8547) );
  XOR U8555 ( .A(n8261), .B(n8541), .Z(n8543) );
  XOR U8556 ( .A(n8549), .B(n8550), .Z(n8261) );
  AND U8557 ( .A(n253), .B(n8500), .Z(n8550) );
  XOR U8558 ( .A(n8549), .B(n8498), .Z(n8500) );
  XOR U8559 ( .A(n8551), .B(n8552), .Z(n8541) );
  AND U8560 ( .A(n8553), .B(n8554), .Z(n8552) );
  XNOR U8561 ( .A(n8551), .B(n8306), .Z(n8554) );
  IV U8562 ( .A(n8309), .Z(n8306) );
  XOR U8563 ( .A(n8555), .B(n8556), .Z(n8309) );
  AND U8564 ( .A(n245), .B(n8557), .Z(n8556) );
  XOR U8565 ( .A(n8558), .B(n8555), .Z(n8557) );
  XOR U8566 ( .A(n8310), .B(n8551), .Z(n8553) );
  XOR U8567 ( .A(n8559), .B(n8560), .Z(n8310) );
  AND U8568 ( .A(n253), .B(n8508), .Z(n8560) );
  XOR U8569 ( .A(n8559), .B(n8506), .Z(n8508) );
  XOR U8570 ( .A(n8447), .B(n8561), .Z(n8551) );
  AND U8571 ( .A(n8449), .B(n8562), .Z(n8561) );
  XNOR U8572 ( .A(n8447), .B(n8403), .Z(n8562) );
  IV U8573 ( .A(n8406), .Z(n8403) );
  XOR U8574 ( .A(n8563), .B(n8564), .Z(n8406) );
  AND U8575 ( .A(n245), .B(n8565), .Z(n8564) );
  XNOR U8576 ( .A(n8566), .B(n8563), .Z(n8565) );
  XOR U8577 ( .A(n8407), .B(n8447), .Z(n8449) );
  XOR U8578 ( .A(n8567), .B(n8568), .Z(n8407) );
  AND U8579 ( .A(n253), .B(n8518), .Z(n8568) );
  XOR U8580 ( .A(n8567), .B(n8516), .Z(n8518) );
  AND U8581 ( .A(n8519), .B(n8427), .Z(n8447) );
  XNOR U8582 ( .A(n8569), .B(n8570), .Z(n8427) );
  AND U8583 ( .A(n245), .B(n8571), .Z(n8570) );
  XNOR U8584 ( .A(n8572), .B(n8569), .Z(n8571) );
  XNOR U8585 ( .A(n8573), .B(n8574), .Z(n245) );
  AND U8586 ( .A(n8575), .B(n8576), .Z(n8574) );
  XOR U8587 ( .A(n8528), .B(n8573), .Z(n8576) );
  AND U8588 ( .A(n8577), .B(n8578), .Z(n8528) );
  XNOR U8589 ( .A(n8525), .B(n8573), .Z(n8575) );
  XNOR U8590 ( .A(n8579), .B(n8580), .Z(n8525) );
  AND U8591 ( .A(n249), .B(n8581), .Z(n8580) );
  XNOR U8592 ( .A(n8582), .B(n8583), .Z(n8581) );
  XOR U8593 ( .A(n8584), .B(n8585), .Z(n8573) );
  AND U8594 ( .A(n8586), .B(n8587), .Z(n8585) );
  XNOR U8595 ( .A(n8584), .B(n8577), .Z(n8587) );
  IV U8596 ( .A(n8538), .Z(n8577) );
  XOR U8597 ( .A(n8588), .B(n8589), .Z(n8538) );
  XOR U8598 ( .A(n8590), .B(n8578), .Z(n8589) );
  AND U8599 ( .A(n8548), .B(n8591), .Z(n8578) );
  AND U8600 ( .A(n8592), .B(n8593), .Z(n8590) );
  XOR U8601 ( .A(n8594), .B(n8588), .Z(n8592) );
  XNOR U8602 ( .A(n8535), .B(n8584), .Z(n8586) );
  XNOR U8603 ( .A(n8595), .B(n8596), .Z(n8535) );
  AND U8604 ( .A(n249), .B(n8597), .Z(n8596) );
  XNOR U8605 ( .A(n8598), .B(n8599), .Z(n8597) );
  XOR U8606 ( .A(n8600), .B(n8601), .Z(n8584) );
  AND U8607 ( .A(n8602), .B(n8603), .Z(n8601) );
  XNOR U8608 ( .A(n8600), .B(n8548), .Z(n8603) );
  XOR U8609 ( .A(n8604), .B(n8593), .Z(n8548) );
  XNOR U8610 ( .A(n8605), .B(n8588), .Z(n8593) );
  XOR U8611 ( .A(n8606), .B(n8607), .Z(n8588) );
  AND U8612 ( .A(n8608), .B(n8609), .Z(n8607) );
  XOR U8613 ( .A(n8610), .B(n8606), .Z(n8608) );
  XNOR U8614 ( .A(n8611), .B(n8612), .Z(n8605) );
  AND U8615 ( .A(n8613), .B(n8614), .Z(n8612) );
  XOR U8616 ( .A(n8611), .B(n8615), .Z(n8613) );
  XNOR U8617 ( .A(n8594), .B(n8591), .Z(n8604) );
  AND U8618 ( .A(n8616), .B(n8617), .Z(n8591) );
  XOR U8619 ( .A(n8618), .B(n8619), .Z(n8594) );
  AND U8620 ( .A(n8620), .B(n8621), .Z(n8619) );
  XOR U8621 ( .A(n8618), .B(n8622), .Z(n8620) );
  XNOR U8622 ( .A(n8545), .B(n8600), .Z(n8602) );
  XNOR U8623 ( .A(n8623), .B(n8624), .Z(n8545) );
  AND U8624 ( .A(n249), .B(n8625), .Z(n8624) );
  XNOR U8625 ( .A(n8626), .B(n8627), .Z(n8625) );
  XOR U8626 ( .A(n8628), .B(n8629), .Z(n8600) );
  AND U8627 ( .A(n8630), .B(n8631), .Z(n8629) );
  XNOR U8628 ( .A(n8628), .B(n8616), .Z(n8631) );
  IV U8629 ( .A(n8558), .Z(n8616) );
  XNOR U8630 ( .A(n8632), .B(n8609), .Z(n8558) );
  XNOR U8631 ( .A(n8633), .B(n8615), .Z(n8609) );
  XOR U8632 ( .A(n8634), .B(n8635), .Z(n8615) );
  AND U8633 ( .A(n8636), .B(n8637), .Z(n8635) );
  XOR U8634 ( .A(n8634), .B(n8638), .Z(n8636) );
  XNOR U8635 ( .A(n8614), .B(n8606), .Z(n8633) );
  XOR U8636 ( .A(n8639), .B(n8640), .Z(n8606) );
  AND U8637 ( .A(n8641), .B(n8642), .Z(n8640) );
  XNOR U8638 ( .A(n8643), .B(n8639), .Z(n8641) );
  XNOR U8639 ( .A(n8644), .B(n8611), .Z(n8614) );
  XOR U8640 ( .A(n8645), .B(n8646), .Z(n8611) );
  AND U8641 ( .A(n8647), .B(n8648), .Z(n8646) );
  XOR U8642 ( .A(n8645), .B(n8649), .Z(n8647) );
  XNOR U8643 ( .A(n8650), .B(n8651), .Z(n8644) );
  AND U8644 ( .A(n8652), .B(n8653), .Z(n8651) );
  XNOR U8645 ( .A(n8650), .B(n8654), .Z(n8652) );
  XNOR U8646 ( .A(n8610), .B(n8617), .Z(n8632) );
  AND U8647 ( .A(n8566), .B(n8655), .Z(n8617) );
  XOR U8648 ( .A(n8622), .B(n8621), .Z(n8610) );
  XNOR U8649 ( .A(n8656), .B(n8618), .Z(n8621) );
  XOR U8650 ( .A(n8657), .B(n8658), .Z(n8618) );
  AND U8651 ( .A(n8659), .B(n8660), .Z(n8658) );
  XOR U8652 ( .A(n8657), .B(n8661), .Z(n8659) );
  XNOR U8653 ( .A(n8662), .B(n8663), .Z(n8656) );
  AND U8654 ( .A(n8664), .B(n8665), .Z(n8663) );
  XOR U8655 ( .A(n8662), .B(n8666), .Z(n8664) );
  XOR U8656 ( .A(n8667), .B(n8668), .Z(n8622) );
  AND U8657 ( .A(n8669), .B(n8670), .Z(n8668) );
  XOR U8658 ( .A(n8667), .B(n8671), .Z(n8669) );
  XNOR U8659 ( .A(n8555), .B(n8628), .Z(n8630) );
  XNOR U8660 ( .A(n8672), .B(n8673), .Z(n8555) );
  AND U8661 ( .A(n249), .B(n8674), .Z(n8673) );
  XNOR U8662 ( .A(n8675), .B(n8676), .Z(n8674) );
  XOR U8663 ( .A(n8677), .B(n8678), .Z(n8628) );
  AND U8664 ( .A(n8679), .B(n8680), .Z(n8678) );
  XNOR U8665 ( .A(n8677), .B(n8566), .Z(n8680) );
  XOR U8666 ( .A(n8681), .B(n8642), .Z(n8566) );
  XNOR U8667 ( .A(n8682), .B(n8649), .Z(n8642) );
  XOR U8668 ( .A(n8638), .B(n8637), .Z(n8649) );
  XNOR U8669 ( .A(n8683), .B(n8634), .Z(n8637) );
  XOR U8670 ( .A(n8684), .B(n8685), .Z(n8634) );
  AND U8671 ( .A(n8686), .B(n8687), .Z(n8685) );
  XNOR U8672 ( .A(n8688), .B(n8689), .Z(n8686) );
  IV U8673 ( .A(n8684), .Z(n8688) );
  XNOR U8674 ( .A(n8690), .B(n8691), .Z(n8683) );
  NOR U8675 ( .A(n8692), .B(n8693), .Z(n8691) );
  XNOR U8676 ( .A(n8690), .B(n8694), .Z(n8692) );
  XOR U8677 ( .A(n8695), .B(n8696), .Z(n8638) );
  NOR U8678 ( .A(n8697), .B(n8698), .Z(n8696) );
  XNOR U8679 ( .A(n8695), .B(n8699), .Z(n8697) );
  XNOR U8680 ( .A(n8648), .B(n8639), .Z(n8682) );
  XOR U8681 ( .A(n8700), .B(n8701), .Z(n8639) );
  AND U8682 ( .A(n8702), .B(n8703), .Z(n8701) );
  XOR U8683 ( .A(n8700), .B(n8704), .Z(n8702) );
  XOR U8684 ( .A(n8705), .B(n8654), .Z(n8648) );
  XOR U8685 ( .A(n8706), .B(n8707), .Z(n8654) );
  NOR U8686 ( .A(n8708), .B(n8709), .Z(n8707) );
  XOR U8687 ( .A(n8706), .B(n8710), .Z(n8708) );
  XNOR U8688 ( .A(n8653), .B(n8645), .Z(n8705) );
  XOR U8689 ( .A(n8711), .B(n8712), .Z(n8645) );
  AND U8690 ( .A(n8713), .B(n8714), .Z(n8712) );
  XOR U8691 ( .A(n8711), .B(n8715), .Z(n8713) );
  XNOR U8692 ( .A(n8716), .B(n8650), .Z(n8653) );
  XOR U8693 ( .A(n8717), .B(n8718), .Z(n8650) );
  AND U8694 ( .A(n8719), .B(n8720), .Z(n8718) );
  XNOR U8695 ( .A(n8721), .B(n8722), .Z(n8719) );
  IV U8696 ( .A(n8717), .Z(n8721) );
  XNOR U8697 ( .A(n8723), .B(n8724), .Z(n8716) );
  NOR U8698 ( .A(n8725), .B(n8726), .Z(n8724) );
  XNOR U8699 ( .A(n8723), .B(n8727), .Z(n8725) );
  XOR U8700 ( .A(n8643), .B(n8655), .Z(n8681) );
  NOR U8701 ( .A(n8572), .B(n8728), .Z(n8655) );
  XNOR U8702 ( .A(n8661), .B(n8660), .Z(n8643) );
  XNOR U8703 ( .A(n8729), .B(n8666), .Z(n8660) );
  XNOR U8704 ( .A(n8730), .B(n8731), .Z(n8666) );
  NOR U8705 ( .A(n8732), .B(n8733), .Z(n8731) );
  XOR U8706 ( .A(n8730), .B(n8734), .Z(n8732) );
  XNOR U8707 ( .A(n8665), .B(n8657), .Z(n8729) );
  XOR U8708 ( .A(n8735), .B(n8736), .Z(n8657) );
  AND U8709 ( .A(n8737), .B(n8738), .Z(n8736) );
  XOR U8710 ( .A(n8735), .B(n8739), .Z(n8737) );
  XNOR U8711 ( .A(n8740), .B(n8662), .Z(n8665) );
  XOR U8712 ( .A(n8741), .B(n8742), .Z(n8662) );
  AND U8713 ( .A(n8743), .B(n8744), .Z(n8742) );
  XNOR U8714 ( .A(n8745), .B(n8746), .Z(n8743) );
  IV U8715 ( .A(n8741), .Z(n8745) );
  XNOR U8716 ( .A(n8747), .B(n8748), .Z(n8740) );
  NOR U8717 ( .A(n8749), .B(n8750), .Z(n8748) );
  XNOR U8718 ( .A(n8747), .B(n8751), .Z(n8749) );
  XOR U8719 ( .A(n8671), .B(n8670), .Z(n8661) );
  XNOR U8720 ( .A(n8752), .B(n8667), .Z(n8670) );
  XOR U8721 ( .A(n8753), .B(n8754), .Z(n8667) );
  AND U8722 ( .A(n8755), .B(n8756), .Z(n8754) );
  XNOR U8723 ( .A(n8757), .B(n8758), .Z(n8755) );
  IV U8724 ( .A(n8753), .Z(n8757) );
  XNOR U8725 ( .A(n8759), .B(n8760), .Z(n8752) );
  NOR U8726 ( .A(n8761), .B(n8762), .Z(n8760) );
  XNOR U8727 ( .A(n8759), .B(n8763), .Z(n8761) );
  XOR U8728 ( .A(n8764), .B(n8765), .Z(n8671) );
  NOR U8729 ( .A(n8766), .B(n8767), .Z(n8765) );
  XNOR U8730 ( .A(n8764), .B(n8768), .Z(n8766) );
  XNOR U8731 ( .A(n8563), .B(n8677), .Z(n8679) );
  XNOR U8732 ( .A(n8769), .B(n8770), .Z(n8563) );
  AND U8733 ( .A(n249), .B(n8771), .Z(n8770) );
  XNOR U8734 ( .A(n8772), .B(n8773), .Z(n8771) );
  AND U8735 ( .A(n8569), .B(n8572), .Z(n8677) );
  XOR U8736 ( .A(n8774), .B(n8728), .Z(n8572) );
  XNOR U8737 ( .A(p_input[192]), .B(p_input[512]), .Z(n8728) );
  XNOR U8738 ( .A(n8704), .B(n8703), .Z(n8774) );
  XNOR U8739 ( .A(n8775), .B(n8715), .Z(n8703) );
  XOR U8740 ( .A(n8689), .B(n8687), .Z(n8715) );
  XNOR U8741 ( .A(n8776), .B(n8694), .Z(n8687) );
  XOR U8742 ( .A(p_input[216]), .B(p_input[536]), .Z(n8694) );
  XOR U8743 ( .A(n8684), .B(n8693), .Z(n8776) );
  XOR U8744 ( .A(n8777), .B(n8690), .Z(n8693) );
  XOR U8745 ( .A(p_input[214]), .B(p_input[534]), .Z(n8690) );
  XOR U8746 ( .A(p_input[215]), .B(n6576), .Z(n8777) );
  XOR U8747 ( .A(p_input[210]), .B(p_input[530]), .Z(n8684) );
  XNOR U8748 ( .A(n8699), .B(n8698), .Z(n8689) );
  XOR U8749 ( .A(n8778), .B(n8695), .Z(n8698) );
  XOR U8750 ( .A(p_input[211]), .B(p_input[531]), .Z(n8695) );
  XOR U8751 ( .A(p_input[212]), .B(n6578), .Z(n8778) );
  XOR U8752 ( .A(p_input[213]), .B(p_input[533]), .Z(n8699) );
  XOR U8753 ( .A(n8714), .B(n8779), .Z(n8775) );
  IV U8754 ( .A(n8700), .Z(n8779) );
  XOR U8755 ( .A(p_input[193]), .B(p_input[513]), .Z(n8700) );
  XNOR U8756 ( .A(n8780), .B(n8722), .Z(n8714) );
  XNOR U8757 ( .A(n8710), .B(n8709), .Z(n8722) );
  XNOR U8758 ( .A(n8781), .B(n8706), .Z(n8709) );
  XNOR U8759 ( .A(p_input[218]), .B(p_input[538]), .Z(n8706) );
  XOR U8760 ( .A(p_input[219]), .B(n6582), .Z(n8781) );
  XOR U8761 ( .A(p_input[220]), .B(p_input[540]), .Z(n8710) );
  XOR U8762 ( .A(n8720), .B(n8782), .Z(n8780) );
  IV U8763 ( .A(n8711), .Z(n8782) );
  XOR U8764 ( .A(p_input[209]), .B(p_input[529]), .Z(n8711) );
  XNOR U8765 ( .A(n8783), .B(n8727), .Z(n8720) );
  XNOR U8766 ( .A(p_input[223]), .B(n6585), .Z(n8727) );
  XOR U8767 ( .A(n8717), .B(n8726), .Z(n8783) );
  XOR U8768 ( .A(n8784), .B(n8723), .Z(n8726) );
  XOR U8769 ( .A(p_input[221]), .B(p_input[541]), .Z(n8723) );
  XOR U8770 ( .A(p_input[222]), .B(n6587), .Z(n8784) );
  XOR U8771 ( .A(p_input[217]), .B(p_input[537]), .Z(n8717) );
  XOR U8772 ( .A(n8739), .B(n8738), .Z(n8704) );
  XNOR U8773 ( .A(n8785), .B(n8746), .Z(n8738) );
  XNOR U8774 ( .A(n8734), .B(n8733), .Z(n8746) );
  XNOR U8775 ( .A(n8786), .B(n8730), .Z(n8733) );
  XNOR U8776 ( .A(p_input[203]), .B(p_input[523]), .Z(n8730) );
  XOR U8777 ( .A(p_input[204]), .B(n6590), .Z(n8786) );
  XOR U8778 ( .A(p_input[205]), .B(p_input[525]), .Z(n8734) );
  XOR U8779 ( .A(n8744), .B(n8787), .Z(n8785) );
  IV U8780 ( .A(n8735), .Z(n8787) );
  XOR U8781 ( .A(p_input[194]), .B(p_input[514]), .Z(n8735) );
  XNOR U8782 ( .A(n8788), .B(n8751), .Z(n8744) );
  XNOR U8783 ( .A(p_input[208]), .B(n6593), .Z(n8751) );
  XOR U8784 ( .A(n8741), .B(n8750), .Z(n8788) );
  XOR U8785 ( .A(n8789), .B(n8747), .Z(n8750) );
  XOR U8786 ( .A(p_input[206]), .B(p_input[526]), .Z(n8747) );
  XOR U8787 ( .A(p_input[207]), .B(n6595), .Z(n8789) );
  XOR U8788 ( .A(p_input[202]), .B(p_input[522]), .Z(n8741) );
  XOR U8789 ( .A(n8758), .B(n8756), .Z(n8739) );
  XNOR U8790 ( .A(n8790), .B(n8763), .Z(n8756) );
  XOR U8791 ( .A(p_input[201]), .B(p_input[521]), .Z(n8763) );
  XOR U8792 ( .A(n8753), .B(n8762), .Z(n8790) );
  XOR U8793 ( .A(n8791), .B(n8759), .Z(n8762) );
  XOR U8794 ( .A(p_input[199]), .B(p_input[519]), .Z(n8759) );
  XOR U8795 ( .A(p_input[200]), .B(n6963), .Z(n8791) );
  XOR U8796 ( .A(p_input[195]), .B(p_input[515]), .Z(n8753) );
  XNOR U8797 ( .A(n8768), .B(n8767), .Z(n8758) );
  XOR U8798 ( .A(n8792), .B(n8764), .Z(n8767) );
  XOR U8799 ( .A(p_input[196]), .B(p_input[516]), .Z(n8764) );
  XOR U8800 ( .A(p_input[197]), .B(n6965), .Z(n8792) );
  XOR U8801 ( .A(p_input[198]), .B(p_input[518]), .Z(n8768) );
  XNOR U8802 ( .A(n8793), .B(n8794), .Z(n8569) );
  AND U8803 ( .A(n249), .B(n8795), .Z(n8794) );
  XNOR U8804 ( .A(n8796), .B(n8797), .Z(n249) );
  AND U8805 ( .A(n8798), .B(n8799), .Z(n8797) );
  XOR U8806 ( .A(n8583), .B(n8796), .Z(n8799) );
  XNOR U8807 ( .A(n8800), .B(n8796), .Z(n8798) );
  XOR U8808 ( .A(n8801), .B(n8802), .Z(n8796) );
  AND U8809 ( .A(n8803), .B(n8804), .Z(n8802) );
  XOR U8810 ( .A(n8598), .B(n8801), .Z(n8804) );
  XOR U8811 ( .A(n8801), .B(n8599), .Z(n8803) );
  XOR U8812 ( .A(n8805), .B(n8806), .Z(n8801) );
  AND U8813 ( .A(n8807), .B(n8808), .Z(n8806) );
  XOR U8814 ( .A(n8626), .B(n8805), .Z(n8808) );
  XOR U8815 ( .A(n8805), .B(n8627), .Z(n8807) );
  XOR U8816 ( .A(n8809), .B(n8810), .Z(n8805) );
  AND U8817 ( .A(n8811), .B(n8812), .Z(n8810) );
  XOR U8818 ( .A(n8675), .B(n8809), .Z(n8812) );
  XOR U8819 ( .A(n8809), .B(n8676), .Z(n8811) );
  XOR U8820 ( .A(n8813), .B(n8814), .Z(n8809) );
  AND U8821 ( .A(n8815), .B(n8816), .Z(n8814) );
  XOR U8822 ( .A(n8813), .B(n8772), .Z(n8816) );
  XNOR U8823 ( .A(n8817), .B(n8818), .Z(n8519) );
  AND U8824 ( .A(n253), .B(n8819), .Z(n8818) );
  XNOR U8825 ( .A(n8820), .B(n8821), .Z(n253) );
  AND U8826 ( .A(n8822), .B(n8823), .Z(n8821) );
  XOR U8827 ( .A(n8820), .B(n8529), .Z(n8823) );
  XNOR U8828 ( .A(n8820), .B(n8479), .Z(n8822) );
  XOR U8829 ( .A(n8824), .B(n8825), .Z(n8820) );
  AND U8830 ( .A(n8826), .B(n8827), .Z(n8825) );
  XNOR U8831 ( .A(n8539), .B(n8824), .Z(n8827) );
  XOR U8832 ( .A(n8824), .B(n8489), .Z(n8826) );
  XOR U8833 ( .A(n8828), .B(n8829), .Z(n8824) );
  AND U8834 ( .A(n8830), .B(n8831), .Z(n8829) );
  XNOR U8835 ( .A(n8549), .B(n8828), .Z(n8831) );
  XOR U8836 ( .A(n8828), .B(n8498), .Z(n8830) );
  XOR U8837 ( .A(n8832), .B(n8833), .Z(n8828) );
  AND U8838 ( .A(n8834), .B(n8835), .Z(n8833) );
  XOR U8839 ( .A(n8832), .B(n8506), .Z(n8834) );
  XOR U8840 ( .A(n8836), .B(n8837), .Z(n8470) );
  AND U8841 ( .A(n257), .B(n8819), .Z(n8837) );
  XNOR U8842 ( .A(n8817), .B(n8836), .Z(n8819) );
  XNOR U8843 ( .A(n8838), .B(n8839), .Z(n257) );
  AND U8844 ( .A(n8840), .B(n8841), .Z(n8839) );
  XNOR U8845 ( .A(n8842), .B(n8838), .Z(n8841) );
  IV U8846 ( .A(n8529), .Z(n8842) );
  XOR U8847 ( .A(n8800), .B(n8843), .Z(n8529) );
  AND U8848 ( .A(n260), .B(n8844), .Z(n8843) );
  XOR U8849 ( .A(n8582), .B(n8579), .Z(n8844) );
  IV U8850 ( .A(n8800), .Z(n8582) );
  XNOR U8851 ( .A(n8479), .B(n8838), .Z(n8840) );
  XOR U8852 ( .A(n8845), .B(n8846), .Z(n8479) );
  AND U8853 ( .A(n276), .B(n8847), .Z(n8846) );
  XOR U8854 ( .A(n8848), .B(n8849), .Z(n8838) );
  AND U8855 ( .A(n8850), .B(n8851), .Z(n8849) );
  XNOR U8856 ( .A(n8848), .B(n8539), .Z(n8851) );
  XOR U8857 ( .A(n8599), .B(n8852), .Z(n8539) );
  AND U8858 ( .A(n260), .B(n8853), .Z(n8852) );
  XOR U8859 ( .A(n8595), .B(n8599), .Z(n8853) );
  XNOR U8860 ( .A(n8854), .B(n8848), .Z(n8850) );
  IV U8861 ( .A(n8489), .Z(n8854) );
  XOR U8862 ( .A(n8855), .B(n8856), .Z(n8489) );
  AND U8863 ( .A(n276), .B(n8857), .Z(n8856) );
  XOR U8864 ( .A(n8858), .B(n8859), .Z(n8848) );
  AND U8865 ( .A(n8860), .B(n8861), .Z(n8859) );
  XNOR U8866 ( .A(n8858), .B(n8549), .Z(n8861) );
  XOR U8867 ( .A(n8627), .B(n8862), .Z(n8549) );
  AND U8868 ( .A(n260), .B(n8863), .Z(n8862) );
  XOR U8869 ( .A(n8623), .B(n8627), .Z(n8863) );
  XOR U8870 ( .A(n8498), .B(n8858), .Z(n8860) );
  XOR U8871 ( .A(n8864), .B(n8865), .Z(n8498) );
  AND U8872 ( .A(n276), .B(n8866), .Z(n8865) );
  XOR U8873 ( .A(n8832), .B(n8867), .Z(n8858) );
  AND U8874 ( .A(n8868), .B(n8835), .Z(n8867) );
  XNOR U8875 ( .A(n8559), .B(n8832), .Z(n8835) );
  XOR U8876 ( .A(n8676), .B(n8869), .Z(n8559) );
  AND U8877 ( .A(n260), .B(n8870), .Z(n8869) );
  XOR U8878 ( .A(n8672), .B(n8676), .Z(n8870) );
  XNOR U8879 ( .A(n8871), .B(n8832), .Z(n8868) );
  IV U8880 ( .A(n8506), .Z(n8871) );
  XOR U8881 ( .A(n8872), .B(n8873), .Z(n8506) );
  AND U8882 ( .A(n276), .B(n8874), .Z(n8873) );
  XOR U8883 ( .A(n8875), .B(n8876), .Z(n8832) );
  AND U8884 ( .A(n8877), .B(n8878), .Z(n8876) );
  XNOR U8885 ( .A(n8875), .B(n8567), .Z(n8878) );
  XOR U8886 ( .A(n8773), .B(n8879), .Z(n8567) );
  AND U8887 ( .A(n260), .B(n8880), .Z(n8879) );
  XOR U8888 ( .A(n8769), .B(n8773), .Z(n8880) );
  XNOR U8889 ( .A(n8881), .B(n8875), .Z(n8877) );
  IV U8890 ( .A(n8516), .Z(n8881) );
  XOR U8891 ( .A(n8882), .B(n8883), .Z(n8516) );
  AND U8892 ( .A(n276), .B(n8884), .Z(n8883) );
  AND U8893 ( .A(n8836), .B(n8817), .Z(n8875) );
  XNOR U8894 ( .A(n8885), .B(n8886), .Z(n8817) );
  AND U8895 ( .A(n260), .B(n8795), .Z(n8886) );
  XNOR U8896 ( .A(n8793), .B(n8885), .Z(n8795) );
  XNOR U8897 ( .A(n8887), .B(n8888), .Z(n260) );
  AND U8898 ( .A(n8889), .B(n8890), .Z(n8888) );
  XNOR U8899 ( .A(n8887), .B(n8579), .Z(n8890) );
  IV U8900 ( .A(n8583), .Z(n8579) );
  XOR U8901 ( .A(n8891), .B(n8892), .Z(n8583) );
  AND U8902 ( .A(n264), .B(n8893), .Z(n8892) );
  XOR U8903 ( .A(n8894), .B(n8891), .Z(n8893) );
  XNOR U8904 ( .A(n8887), .B(n8800), .Z(n8889) );
  XOR U8905 ( .A(n8895), .B(n8896), .Z(n8800) );
  AND U8906 ( .A(n272), .B(n8847), .Z(n8896) );
  XOR U8907 ( .A(n8845), .B(n8895), .Z(n8847) );
  XOR U8908 ( .A(n8897), .B(n8898), .Z(n8887) );
  AND U8909 ( .A(n8899), .B(n8900), .Z(n8898) );
  XNOR U8910 ( .A(n8897), .B(n8595), .Z(n8900) );
  IV U8911 ( .A(n8598), .Z(n8595) );
  XOR U8912 ( .A(n8901), .B(n8902), .Z(n8598) );
  AND U8913 ( .A(n264), .B(n8903), .Z(n8902) );
  XOR U8914 ( .A(n8904), .B(n8901), .Z(n8903) );
  XOR U8915 ( .A(n8599), .B(n8897), .Z(n8899) );
  XOR U8916 ( .A(n8905), .B(n8906), .Z(n8599) );
  AND U8917 ( .A(n272), .B(n8857), .Z(n8906) );
  XOR U8918 ( .A(n8905), .B(n8855), .Z(n8857) );
  XOR U8919 ( .A(n8907), .B(n8908), .Z(n8897) );
  AND U8920 ( .A(n8909), .B(n8910), .Z(n8908) );
  XNOR U8921 ( .A(n8907), .B(n8623), .Z(n8910) );
  IV U8922 ( .A(n8626), .Z(n8623) );
  XOR U8923 ( .A(n8911), .B(n8912), .Z(n8626) );
  AND U8924 ( .A(n264), .B(n8913), .Z(n8912) );
  XNOR U8925 ( .A(n8914), .B(n8911), .Z(n8913) );
  XOR U8926 ( .A(n8627), .B(n8907), .Z(n8909) );
  XOR U8927 ( .A(n8915), .B(n8916), .Z(n8627) );
  AND U8928 ( .A(n272), .B(n8866), .Z(n8916) );
  XOR U8929 ( .A(n8915), .B(n8864), .Z(n8866) );
  XOR U8930 ( .A(n8917), .B(n8918), .Z(n8907) );
  AND U8931 ( .A(n8919), .B(n8920), .Z(n8918) );
  XNOR U8932 ( .A(n8917), .B(n8672), .Z(n8920) );
  IV U8933 ( .A(n8675), .Z(n8672) );
  XOR U8934 ( .A(n8921), .B(n8922), .Z(n8675) );
  AND U8935 ( .A(n264), .B(n8923), .Z(n8922) );
  XOR U8936 ( .A(n8924), .B(n8921), .Z(n8923) );
  XOR U8937 ( .A(n8676), .B(n8917), .Z(n8919) );
  XOR U8938 ( .A(n8925), .B(n8926), .Z(n8676) );
  AND U8939 ( .A(n272), .B(n8874), .Z(n8926) );
  XOR U8940 ( .A(n8925), .B(n8872), .Z(n8874) );
  XOR U8941 ( .A(n8813), .B(n8927), .Z(n8917) );
  AND U8942 ( .A(n8815), .B(n8928), .Z(n8927) );
  XNOR U8943 ( .A(n8813), .B(n8769), .Z(n8928) );
  IV U8944 ( .A(n8772), .Z(n8769) );
  XOR U8945 ( .A(n8929), .B(n8930), .Z(n8772) );
  AND U8946 ( .A(n264), .B(n8931), .Z(n8930) );
  XNOR U8947 ( .A(n8932), .B(n8929), .Z(n8931) );
  XOR U8948 ( .A(n8773), .B(n8813), .Z(n8815) );
  XOR U8949 ( .A(n8933), .B(n8934), .Z(n8773) );
  AND U8950 ( .A(n272), .B(n8884), .Z(n8934) );
  XOR U8951 ( .A(n8933), .B(n8882), .Z(n8884) );
  AND U8952 ( .A(n8885), .B(n8793), .Z(n8813) );
  XNOR U8953 ( .A(n8935), .B(n8936), .Z(n8793) );
  AND U8954 ( .A(n264), .B(n8937), .Z(n8936) );
  XNOR U8955 ( .A(n8938), .B(n8935), .Z(n8937) );
  XNOR U8956 ( .A(n8939), .B(n8940), .Z(n264) );
  AND U8957 ( .A(n8941), .B(n8942), .Z(n8940) );
  XOR U8958 ( .A(n8894), .B(n8939), .Z(n8942) );
  AND U8959 ( .A(n8943), .B(n8944), .Z(n8894) );
  XNOR U8960 ( .A(n8891), .B(n8939), .Z(n8941) );
  XNOR U8961 ( .A(n8945), .B(n8946), .Z(n8891) );
  AND U8962 ( .A(n268), .B(n8947), .Z(n8946) );
  XNOR U8963 ( .A(n8948), .B(n8949), .Z(n8947) );
  XOR U8964 ( .A(n8950), .B(n8951), .Z(n8939) );
  AND U8965 ( .A(n8952), .B(n8953), .Z(n8951) );
  XNOR U8966 ( .A(n8950), .B(n8943), .Z(n8953) );
  IV U8967 ( .A(n8904), .Z(n8943) );
  XOR U8968 ( .A(n8954), .B(n8955), .Z(n8904) );
  XOR U8969 ( .A(n8956), .B(n8944), .Z(n8955) );
  AND U8970 ( .A(n8914), .B(n8957), .Z(n8944) );
  AND U8971 ( .A(n8958), .B(n8959), .Z(n8956) );
  XOR U8972 ( .A(n8960), .B(n8954), .Z(n8958) );
  XNOR U8973 ( .A(n8901), .B(n8950), .Z(n8952) );
  XNOR U8974 ( .A(n8961), .B(n8962), .Z(n8901) );
  AND U8975 ( .A(n268), .B(n8963), .Z(n8962) );
  XNOR U8976 ( .A(n8964), .B(n8965), .Z(n8963) );
  XOR U8977 ( .A(n8966), .B(n8967), .Z(n8950) );
  AND U8978 ( .A(n8968), .B(n8969), .Z(n8967) );
  XNOR U8979 ( .A(n8966), .B(n8914), .Z(n8969) );
  XOR U8980 ( .A(n8970), .B(n8959), .Z(n8914) );
  XNOR U8981 ( .A(n8971), .B(n8954), .Z(n8959) );
  XOR U8982 ( .A(n8972), .B(n8973), .Z(n8954) );
  AND U8983 ( .A(n8974), .B(n8975), .Z(n8973) );
  XOR U8984 ( .A(n8976), .B(n8972), .Z(n8974) );
  XNOR U8985 ( .A(n8977), .B(n8978), .Z(n8971) );
  AND U8986 ( .A(n8979), .B(n8980), .Z(n8978) );
  XOR U8987 ( .A(n8977), .B(n8981), .Z(n8979) );
  XNOR U8988 ( .A(n8960), .B(n8957), .Z(n8970) );
  AND U8989 ( .A(n8982), .B(n8983), .Z(n8957) );
  XOR U8990 ( .A(n8984), .B(n8985), .Z(n8960) );
  AND U8991 ( .A(n8986), .B(n8987), .Z(n8985) );
  XOR U8992 ( .A(n8984), .B(n8988), .Z(n8986) );
  XNOR U8993 ( .A(n8911), .B(n8966), .Z(n8968) );
  XNOR U8994 ( .A(n8989), .B(n8990), .Z(n8911) );
  AND U8995 ( .A(n268), .B(n8991), .Z(n8990) );
  XNOR U8996 ( .A(n8992), .B(n8993), .Z(n8991) );
  XOR U8997 ( .A(n8994), .B(n8995), .Z(n8966) );
  AND U8998 ( .A(n8996), .B(n8997), .Z(n8995) );
  XNOR U8999 ( .A(n8994), .B(n8982), .Z(n8997) );
  IV U9000 ( .A(n8924), .Z(n8982) );
  XNOR U9001 ( .A(n8998), .B(n8975), .Z(n8924) );
  XNOR U9002 ( .A(n8999), .B(n8981), .Z(n8975) );
  XOR U9003 ( .A(n9000), .B(n9001), .Z(n8981) );
  AND U9004 ( .A(n9002), .B(n9003), .Z(n9001) );
  XOR U9005 ( .A(n9000), .B(n9004), .Z(n9002) );
  XNOR U9006 ( .A(n8980), .B(n8972), .Z(n8999) );
  XOR U9007 ( .A(n9005), .B(n9006), .Z(n8972) );
  AND U9008 ( .A(n9007), .B(n9008), .Z(n9006) );
  XNOR U9009 ( .A(n9009), .B(n9005), .Z(n9007) );
  XNOR U9010 ( .A(n9010), .B(n8977), .Z(n8980) );
  XOR U9011 ( .A(n9011), .B(n9012), .Z(n8977) );
  AND U9012 ( .A(n9013), .B(n9014), .Z(n9012) );
  XOR U9013 ( .A(n9011), .B(n9015), .Z(n9013) );
  XNOR U9014 ( .A(n9016), .B(n9017), .Z(n9010) );
  AND U9015 ( .A(n9018), .B(n9019), .Z(n9017) );
  XNOR U9016 ( .A(n9016), .B(n9020), .Z(n9018) );
  XNOR U9017 ( .A(n8976), .B(n8983), .Z(n8998) );
  AND U9018 ( .A(n8932), .B(n9021), .Z(n8983) );
  XOR U9019 ( .A(n8988), .B(n8987), .Z(n8976) );
  XNOR U9020 ( .A(n9022), .B(n8984), .Z(n8987) );
  XOR U9021 ( .A(n9023), .B(n9024), .Z(n8984) );
  AND U9022 ( .A(n9025), .B(n9026), .Z(n9024) );
  XOR U9023 ( .A(n9023), .B(n9027), .Z(n9025) );
  XNOR U9024 ( .A(n9028), .B(n9029), .Z(n9022) );
  AND U9025 ( .A(n9030), .B(n9031), .Z(n9029) );
  XOR U9026 ( .A(n9028), .B(n9032), .Z(n9030) );
  XOR U9027 ( .A(n9033), .B(n9034), .Z(n8988) );
  AND U9028 ( .A(n9035), .B(n9036), .Z(n9034) );
  XOR U9029 ( .A(n9033), .B(n9037), .Z(n9035) );
  XNOR U9030 ( .A(n8921), .B(n8994), .Z(n8996) );
  XNOR U9031 ( .A(n9038), .B(n9039), .Z(n8921) );
  AND U9032 ( .A(n268), .B(n9040), .Z(n9039) );
  XNOR U9033 ( .A(n9041), .B(n9042), .Z(n9040) );
  XOR U9034 ( .A(n9043), .B(n9044), .Z(n8994) );
  AND U9035 ( .A(n9045), .B(n9046), .Z(n9044) );
  XNOR U9036 ( .A(n9043), .B(n8932), .Z(n9046) );
  XOR U9037 ( .A(n9047), .B(n9008), .Z(n8932) );
  XNOR U9038 ( .A(n9048), .B(n9015), .Z(n9008) );
  XOR U9039 ( .A(n9004), .B(n9003), .Z(n9015) );
  XNOR U9040 ( .A(n9049), .B(n9000), .Z(n9003) );
  XOR U9041 ( .A(n9050), .B(n9051), .Z(n9000) );
  AND U9042 ( .A(n9052), .B(n9053), .Z(n9051) );
  XNOR U9043 ( .A(n9054), .B(n9055), .Z(n9052) );
  IV U9044 ( .A(n9050), .Z(n9054) );
  XNOR U9045 ( .A(n9056), .B(n9057), .Z(n9049) );
  NOR U9046 ( .A(n9058), .B(n9059), .Z(n9057) );
  XNOR U9047 ( .A(n9056), .B(n9060), .Z(n9058) );
  XOR U9048 ( .A(n9061), .B(n9062), .Z(n9004) );
  NOR U9049 ( .A(n9063), .B(n9064), .Z(n9062) );
  XNOR U9050 ( .A(n9061), .B(n9065), .Z(n9063) );
  XNOR U9051 ( .A(n9014), .B(n9005), .Z(n9048) );
  XOR U9052 ( .A(n9066), .B(n9067), .Z(n9005) );
  AND U9053 ( .A(n9068), .B(n9069), .Z(n9067) );
  XOR U9054 ( .A(n9066), .B(n9070), .Z(n9068) );
  XOR U9055 ( .A(n9071), .B(n9020), .Z(n9014) );
  XOR U9056 ( .A(n9072), .B(n9073), .Z(n9020) );
  NOR U9057 ( .A(n9074), .B(n9075), .Z(n9073) );
  XOR U9058 ( .A(n9072), .B(n9076), .Z(n9074) );
  XNOR U9059 ( .A(n9019), .B(n9011), .Z(n9071) );
  XOR U9060 ( .A(n9077), .B(n9078), .Z(n9011) );
  AND U9061 ( .A(n9079), .B(n9080), .Z(n9078) );
  XOR U9062 ( .A(n9077), .B(n9081), .Z(n9079) );
  XNOR U9063 ( .A(n9082), .B(n9016), .Z(n9019) );
  XOR U9064 ( .A(n9083), .B(n9084), .Z(n9016) );
  AND U9065 ( .A(n9085), .B(n9086), .Z(n9084) );
  XNOR U9066 ( .A(n9087), .B(n9088), .Z(n9085) );
  IV U9067 ( .A(n9083), .Z(n9087) );
  XNOR U9068 ( .A(n9089), .B(n9090), .Z(n9082) );
  NOR U9069 ( .A(n9091), .B(n9092), .Z(n9090) );
  XNOR U9070 ( .A(n9089), .B(n9093), .Z(n9091) );
  XOR U9071 ( .A(n9009), .B(n9021), .Z(n9047) );
  NOR U9072 ( .A(n8938), .B(n9094), .Z(n9021) );
  XNOR U9073 ( .A(n9027), .B(n9026), .Z(n9009) );
  XNOR U9074 ( .A(n9095), .B(n9032), .Z(n9026) );
  XNOR U9075 ( .A(n9096), .B(n9097), .Z(n9032) );
  NOR U9076 ( .A(n9098), .B(n9099), .Z(n9097) );
  XOR U9077 ( .A(n9096), .B(n9100), .Z(n9098) );
  XNOR U9078 ( .A(n9031), .B(n9023), .Z(n9095) );
  XOR U9079 ( .A(n9101), .B(n9102), .Z(n9023) );
  AND U9080 ( .A(n9103), .B(n9104), .Z(n9102) );
  XOR U9081 ( .A(n9101), .B(n9105), .Z(n9103) );
  XNOR U9082 ( .A(n9106), .B(n9028), .Z(n9031) );
  XOR U9083 ( .A(n9107), .B(n9108), .Z(n9028) );
  AND U9084 ( .A(n9109), .B(n9110), .Z(n9108) );
  XNOR U9085 ( .A(n9111), .B(n9112), .Z(n9109) );
  IV U9086 ( .A(n9107), .Z(n9111) );
  XNOR U9087 ( .A(n9113), .B(n9114), .Z(n9106) );
  NOR U9088 ( .A(n9115), .B(n9116), .Z(n9114) );
  XNOR U9089 ( .A(n9113), .B(n9117), .Z(n9115) );
  XOR U9090 ( .A(n9037), .B(n9036), .Z(n9027) );
  XNOR U9091 ( .A(n9118), .B(n9033), .Z(n9036) );
  XOR U9092 ( .A(n9119), .B(n9120), .Z(n9033) );
  AND U9093 ( .A(n9121), .B(n9122), .Z(n9120) );
  XNOR U9094 ( .A(n9123), .B(n9124), .Z(n9121) );
  IV U9095 ( .A(n9119), .Z(n9123) );
  XNOR U9096 ( .A(n9125), .B(n9126), .Z(n9118) );
  NOR U9097 ( .A(n9127), .B(n9128), .Z(n9126) );
  XNOR U9098 ( .A(n9125), .B(n9129), .Z(n9127) );
  XOR U9099 ( .A(n9130), .B(n9131), .Z(n9037) );
  NOR U9100 ( .A(n9132), .B(n9133), .Z(n9131) );
  XNOR U9101 ( .A(n9130), .B(n9134), .Z(n9132) );
  XNOR U9102 ( .A(n8929), .B(n9043), .Z(n9045) );
  XNOR U9103 ( .A(n9135), .B(n9136), .Z(n8929) );
  AND U9104 ( .A(n268), .B(n9137), .Z(n9136) );
  XNOR U9105 ( .A(n9138), .B(n9139), .Z(n9137) );
  AND U9106 ( .A(n8935), .B(n8938), .Z(n9043) );
  XOR U9107 ( .A(n9140), .B(n9094), .Z(n8938) );
  XNOR U9108 ( .A(p_input[224]), .B(p_input[512]), .Z(n9094) );
  XNOR U9109 ( .A(n9070), .B(n9069), .Z(n9140) );
  XNOR U9110 ( .A(n9141), .B(n9081), .Z(n9069) );
  XOR U9111 ( .A(n9055), .B(n9053), .Z(n9081) );
  XNOR U9112 ( .A(n9142), .B(n9060), .Z(n9053) );
  XOR U9113 ( .A(p_input[248]), .B(p_input[536]), .Z(n9060) );
  XOR U9114 ( .A(n9050), .B(n9059), .Z(n9142) );
  XOR U9115 ( .A(n9143), .B(n9056), .Z(n9059) );
  XOR U9116 ( .A(p_input[246]), .B(p_input[534]), .Z(n9056) );
  XOR U9117 ( .A(p_input[247]), .B(n6576), .Z(n9143) );
  XOR U9118 ( .A(p_input[242]), .B(p_input[530]), .Z(n9050) );
  XNOR U9119 ( .A(n9065), .B(n9064), .Z(n9055) );
  XOR U9120 ( .A(n9144), .B(n9061), .Z(n9064) );
  XOR U9121 ( .A(p_input[243]), .B(p_input[531]), .Z(n9061) );
  XOR U9122 ( .A(p_input[244]), .B(n6578), .Z(n9144) );
  XOR U9123 ( .A(p_input[245]), .B(p_input[533]), .Z(n9065) );
  XOR U9124 ( .A(n9080), .B(n9145), .Z(n9141) );
  IV U9125 ( .A(n9066), .Z(n9145) );
  XOR U9126 ( .A(p_input[225]), .B(p_input[513]), .Z(n9066) );
  XNOR U9127 ( .A(n9146), .B(n9088), .Z(n9080) );
  XNOR U9128 ( .A(n9076), .B(n9075), .Z(n9088) );
  XNOR U9129 ( .A(n9147), .B(n9072), .Z(n9075) );
  XNOR U9130 ( .A(p_input[250]), .B(p_input[538]), .Z(n9072) );
  XOR U9131 ( .A(p_input[251]), .B(n6582), .Z(n9147) );
  XOR U9132 ( .A(p_input[252]), .B(p_input[540]), .Z(n9076) );
  XOR U9133 ( .A(n9086), .B(n9148), .Z(n9146) );
  IV U9134 ( .A(n9077), .Z(n9148) );
  XOR U9135 ( .A(p_input[241]), .B(p_input[529]), .Z(n9077) );
  XNOR U9136 ( .A(n9149), .B(n9093), .Z(n9086) );
  XNOR U9137 ( .A(p_input[255]), .B(n6585), .Z(n9093) );
  XOR U9138 ( .A(n9083), .B(n9092), .Z(n9149) );
  XOR U9139 ( .A(n9150), .B(n9089), .Z(n9092) );
  XOR U9140 ( .A(p_input[253]), .B(p_input[541]), .Z(n9089) );
  XOR U9141 ( .A(p_input[254]), .B(n6587), .Z(n9150) );
  XOR U9142 ( .A(p_input[249]), .B(p_input[537]), .Z(n9083) );
  XOR U9143 ( .A(n9105), .B(n9104), .Z(n9070) );
  XNOR U9144 ( .A(n9151), .B(n9112), .Z(n9104) );
  XNOR U9145 ( .A(n9100), .B(n9099), .Z(n9112) );
  XNOR U9146 ( .A(n9152), .B(n9096), .Z(n9099) );
  XNOR U9147 ( .A(p_input[235]), .B(p_input[523]), .Z(n9096) );
  XOR U9148 ( .A(p_input[236]), .B(n6590), .Z(n9152) );
  XOR U9149 ( .A(p_input[237]), .B(p_input[525]), .Z(n9100) );
  XOR U9150 ( .A(n9110), .B(n9153), .Z(n9151) );
  IV U9151 ( .A(n9101), .Z(n9153) );
  XOR U9152 ( .A(p_input[226]), .B(p_input[514]), .Z(n9101) );
  XNOR U9153 ( .A(n9154), .B(n9117), .Z(n9110) );
  XNOR U9154 ( .A(p_input[240]), .B(n6593), .Z(n9117) );
  XOR U9155 ( .A(n9107), .B(n9116), .Z(n9154) );
  XOR U9156 ( .A(n9155), .B(n9113), .Z(n9116) );
  XOR U9157 ( .A(p_input[238]), .B(p_input[526]), .Z(n9113) );
  XOR U9158 ( .A(p_input[239]), .B(n6595), .Z(n9155) );
  XOR U9159 ( .A(p_input[234]), .B(p_input[522]), .Z(n9107) );
  XOR U9160 ( .A(n9124), .B(n9122), .Z(n9105) );
  XNOR U9161 ( .A(n9156), .B(n9129), .Z(n9122) );
  XOR U9162 ( .A(p_input[233]), .B(p_input[521]), .Z(n9129) );
  XOR U9163 ( .A(n9119), .B(n9128), .Z(n9156) );
  XOR U9164 ( .A(n9157), .B(n9125), .Z(n9128) );
  XOR U9165 ( .A(p_input[231]), .B(p_input[519]), .Z(n9125) );
  XOR U9166 ( .A(p_input[232]), .B(n6963), .Z(n9157) );
  XOR U9167 ( .A(p_input[227]), .B(p_input[515]), .Z(n9119) );
  XNOR U9168 ( .A(n9134), .B(n9133), .Z(n9124) );
  XOR U9169 ( .A(n9158), .B(n9130), .Z(n9133) );
  XOR U9170 ( .A(p_input[228]), .B(p_input[516]), .Z(n9130) );
  XOR U9171 ( .A(p_input[229]), .B(n6965), .Z(n9158) );
  XOR U9172 ( .A(p_input[230]), .B(p_input[518]), .Z(n9134) );
  XNOR U9173 ( .A(n9159), .B(n9160), .Z(n8935) );
  AND U9174 ( .A(n268), .B(n9161), .Z(n9160) );
  XNOR U9175 ( .A(n9162), .B(n9163), .Z(n268) );
  AND U9176 ( .A(n9164), .B(n9165), .Z(n9163) );
  XOR U9177 ( .A(n8949), .B(n9162), .Z(n9165) );
  XNOR U9178 ( .A(n9166), .B(n9162), .Z(n9164) );
  XOR U9179 ( .A(n9167), .B(n9168), .Z(n9162) );
  AND U9180 ( .A(n9169), .B(n9170), .Z(n9168) );
  XOR U9181 ( .A(n8964), .B(n9167), .Z(n9170) );
  XOR U9182 ( .A(n9167), .B(n8965), .Z(n9169) );
  XOR U9183 ( .A(n9171), .B(n9172), .Z(n9167) );
  AND U9184 ( .A(n9173), .B(n9174), .Z(n9172) );
  XOR U9185 ( .A(n8992), .B(n9171), .Z(n9174) );
  XOR U9186 ( .A(n9171), .B(n8993), .Z(n9173) );
  XOR U9187 ( .A(n9175), .B(n9176), .Z(n9171) );
  AND U9188 ( .A(n9177), .B(n9178), .Z(n9176) );
  XOR U9189 ( .A(n9041), .B(n9175), .Z(n9178) );
  XOR U9190 ( .A(n9175), .B(n9042), .Z(n9177) );
  XOR U9191 ( .A(n9179), .B(n9180), .Z(n9175) );
  AND U9192 ( .A(n9181), .B(n9182), .Z(n9180) );
  XOR U9193 ( .A(n9179), .B(n9138), .Z(n9182) );
  XNOR U9194 ( .A(n9183), .B(n9184), .Z(n8885) );
  AND U9195 ( .A(n272), .B(n9185), .Z(n9184) );
  XNOR U9196 ( .A(n9186), .B(n9187), .Z(n272) );
  AND U9197 ( .A(n9188), .B(n9189), .Z(n9187) );
  XOR U9198 ( .A(n9186), .B(n8895), .Z(n9189) );
  XNOR U9199 ( .A(n9186), .B(n8845), .Z(n9188) );
  XOR U9200 ( .A(n9190), .B(n9191), .Z(n9186) );
  AND U9201 ( .A(n9192), .B(n9193), .Z(n9191) );
  XNOR U9202 ( .A(n8905), .B(n9190), .Z(n9193) );
  XOR U9203 ( .A(n9190), .B(n8855), .Z(n9192) );
  XOR U9204 ( .A(n9194), .B(n9195), .Z(n9190) );
  AND U9205 ( .A(n9196), .B(n9197), .Z(n9195) );
  XNOR U9206 ( .A(n8915), .B(n9194), .Z(n9197) );
  XOR U9207 ( .A(n9194), .B(n8864), .Z(n9196) );
  XOR U9208 ( .A(n9198), .B(n9199), .Z(n9194) );
  AND U9209 ( .A(n9200), .B(n9201), .Z(n9199) );
  XOR U9210 ( .A(n9198), .B(n8872), .Z(n9200) );
  XOR U9211 ( .A(n9202), .B(n9203), .Z(n8836) );
  AND U9212 ( .A(n276), .B(n9185), .Z(n9203) );
  XNOR U9213 ( .A(n9183), .B(n9202), .Z(n9185) );
  XNOR U9214 ( .A(n9204), .B(n9205), .Z(n276) );
  AND U9215 ( .A(n9206), .B(n9207), .Z(n9205) );
  XNOR U9216 ( .A(n9208), .B(n9204), .Z(n9207) );
  IV U9217 ( .A(n8895), .Z(n9208) );
  XOR U9218 ( .A(n9166), .B(n9209), .Z(n8895) );
  AND U9219 ( .A(n279), .B(n9210), .Z(n9209) );
  XOR U9220 ( .A(n8948), .B(n8945), .Z(n9210) );
  IV U9221 ( .A(n9166), .Z(n8948) );
  XNOR U9222 ( .A(n8845), .B(n9204), .Z(n9206) );
  XOR U9223 ( .A(n9211), .B(n9212), .Z(n8845) );
  AND U9224 ( .A(n295), .B(n9213), .Z(n9212) );
  XOR U9225 ( .A(n9214), .B(n9215), .Z(n9204) );
  AND U9226 ( .A(n9216), .B(n9217), .Z(n9215) );
  XNOR U9227 ( .A(n9214), .B(n8905), .Z(n9217) );
  XOR U9228 ( .A(n8965), .B(n9218), .Z(n8905) );
  AND U9229 ( .A(n279), .B(n9219), .Z(n9218) );
  XOR U9230 ( .A(n8961), .B(n8965), .Z(n9219) );
  XNOR U9231 ( .A(n9220), .B(n9214), .Z(n9216) );
  IV U9232 ( .A(n8855), .Z(n9220) );
  XOR U9233 ( .A(n9221), .B(n9222), .Z(n8855) );
  AND U9234 ( .A(n295), .B(n9223), .Z(n9222) );
  XOR U9235 ( .A(n9224), .B(n9225), .Z(n9214) );
  AND U9236 ( .A(n9226), .B(n9227), .Z(n9225) );
  XNOR U9237 ( .A(n9224), .B(n8915), .Z(n9227) );
  XOR U9238 ( .A(n8993), .B(n9228), .Z(n8915) );
  AND U9239 ( .A(n279), .B(n9229), .Z(n9228) );
  XOR U9240 ( .A(n8989), .B(n8993), .Z(n9229) );
  XOR U9241 ( .A(n8864), .B(n9224), .Z(n9226) );
  XOR U9242 ( .A(n9230), .B(n9231), .Z(n8864) );
  AND U9243 ( .A(n295), .B(n9232), .Z(n9231) );
  XOR U9244 ( .A(n9198), .B(n9233), .Z(n9224) );
  AND U9245 ( .A(n9234), .B(n9201), .Z(n9233) );
  XNOR U9246 ( .A(n8925), .B(n9198), .Z(n9201) );
  XOR U9247 ( .A(n9042), .B(n9235), .Z(n8925) );
  AND U9248 ( .A(n279), .B(n9236), .Z(n9235) );
  XOR U9249 ( .A(n9038), .B(n9042), .Z(n9236) );
  XNOR U9250 ( .A(n9237), .B(n9198), .Z(n9234) );
  IV U9251 ( .A(n8872), .Z(n9237) );
  XOR U9252 ( .A(n9238), .B(n9239), .Z(n8872) );
  AND U9253 ( .A(n295), .B(n9240), .Z(n9239) );
  XOR U9254 ( .A(n9241), .B(n9242), .Z(n9198) );
  AND U9255 ( .A(n9243), .B(n9244), .Z(n9242) );
  XNOR U9256 ( .A(n9241), .B(n8933), .Z(n9244) );
  XOR U9257 ( .A(n9139), .B(n9245), .Z(n8933) );
  AND U9258 ( .A(n279), .B(n9246), .Z(n9245) );
  XOR U9259 ( .A(n9135), .B(n9139), .Z(n9246) );
  XNOR U9260 ( .A(n9247), .B(n9241), .Z(n9243) );
  IV U9261 ( .A(n8882), .Z(n9247) );
  XOR U9262 ( .A(n9248), .B(n9249), .Z(n8882) );
  AND U9263 ( .A(n295), .B(n9250), .Z(n9249) );
  AND U9264 ( .A(n9202), .B(n9183), .Z(n9241) );
  XNOR U9265 ( .A(n9251), .B(n9252), .Z(n9183) );
  AND U9266 ( .A(n279), .B(n9161), .Z(n9252) );
  XNOR U9267 ( .A(n9159), .B(n9251), .Z(n9161) );
  XNOR U9268 ( .A(n9253), .B(n9254), .Z(n279) );
  AND U9269 ( .A(n9255), .B(n9256), .Z(n9254) );
  XNOR U9270 ( .A(n9253), .B(n8945), .Z(n9256) );
  IV U9271 ( .A(n8949), .Z(n8945) );
  XOR U9272 ( .A(n9257), .B(n9258), .Z(n8949) );
  AND U9273 ( .A(n283), .B(n9259), .Z(n9258) );
  XOR U9274 ( .A(n9260), .B(n9257), .Z(n9259) );
  XNOR U9275 ( .A(n9253), .B(n9166), .Z(n9255) );
  XOR U9276 ( .A(n9261), .B(n9262), .Z(n9166) );
  AND U9277 ( .A(n291), .B(n9213), .Z(n9262) );
  XOR U9278 ( .A(n9211), .B(n9261), .Z(n9213) );
  XOR U9279 ( .A(n9263), .B(n9264), .Z(n9253) );
  AND U9280 ( .A(n9265), .B(n9266), .Z(n9264) );
  XNOR U9281 ( .A(n9263), .B(n8961), .Z(n9266) );
  IV U9282 ( .A(n8964), .Z(n8961) );
  XOR U9283 ( .A(n9267), .B(n9268), .Z(n8964) );
  AND U9284 ( .A(n283), .B(n9269), .Z(n9268) );
  XOR U9285 ( .A(n9270), .B(n9267), .Z(n9269) );
  XOR U9286 ( .A(n8965), .B(n9263), .Z(n9265) );
  XOR U9287 ( .A(n9271), .B(n9272), .Z(n8965) );
  AND U9288 ( .A(n291), .B(n9223), .Z(n9272) );
  XOR U9289 ( .A(n9271), .B(n9221), .Z(n9223) );
  XOR U9290 ( .A(n9273), .B(n9274), .Z(n9263) );
  AND U9291 ( .A(n9275), .B(n9276), .Z(n9274) );
  XNOR U9292 ( .A(n9273), .B(n8989), .Z(n9276) );
  IV U9293 ( .A(n8992), .Z(n8989) );
  XOR U9294 ( .A(n9277), .B(n9278), .Z(n8992) );
  AND U9295 ( .A(n283), .B(n9279), .Z(n9278) );
  XNOR U9296 ( .A(n9280), .B(n9277), .Z(n9279) );
  XOR U9297 ( .A(n8993), .B(n9273), .Z(n9275) );
  XOR U9298 ( .A(n9281), .B(n9282), .Z(n8993) );
  AND U9299 ( .A(n291), .B(n9232), .Z(n9282) );
  XOR U9300 ( .A(n9281), .B(n9230), .Z(n9232) );
  XOR U9301 ( .A(n9283), .B(n9284), .Z(n9273) );
  AND U9302 ( .A(n9285), .B(n9286), .Z(n9284) );
  XNOR U9303 ( .A(n9283), .B(n9038), .Z(n9286) );
  IV U9304 ( .A(n9041), .Z(n9038) );
  XOR U9305 ( .A(n9287), .B(n9288), .Z(n9041) );
  AND U9306 ( .A(n283), .B(n9289), .Z(n9288) );
  XOR U9307 ( .A(n9290), .B(n9287), .Z(n9289) );
  XOR U9308 ( .A(n9042), .B(n9283), .Z(n9285) );
  XOR U9309 ( .A(n9291), .B(n9292), .Z(n9042) );
  AND U9310 ( .A(n291), .B(n9240), .Z(n9292) );
  XOR U9311 ( .A(n9291), .B(n9238), .Z(n9240) );
  XOR U9312 ( .A(n9179), .B(n9293), .Z(n9283) );
  AND U9313 ( .A(n9181), .B(n9294), .Z(n9293) );
  XNOR U9314 ( .A(n9179), .B(n9135), .Z(n9294) );
  IV U9315 ( .A(n9138), .Z(n9135) );
  XOR U9316 ( .A(n9295), .B(n9296), .Z(n9138) );
  AND U9317 ( .A(n283), .B(n9297), .Z(n9296) );
  XNOR U9318 ( .A(n9298), .B(n9295), .Z(n9297) );
  XOR U9319 ( .A(n9139), .B(n9179), .Z(n9181) );
  XOR U9320 ( .A(n9299), .B(n9300), .Z(n9139) );
  AND U9321 ( .A(n291), .B(n9250), .Z(n9300) );
  XOR U9322 ( .A(n9299), .B(n9248), .Z(n9250) );
  AND U9323 ( .A(n9251), .B(n9159), .Z(n9179) );
  XNOR U9324 ( .A(n9301), .B(n9302), .Z(n9159) );
  AND U9325 ( .A(n283), .B(n9303), .Z(n9302) );
  XNOR U9326 ( .A(n9304), .B(n9301), .Z(n9303) );
  XNOR U9327 ( .A(n9305), .B(n9306), .Z(n283) );
  AND U9328 ( .A(n9307), .B(n9308), .Z(n9306) );
  XOR U9329 ( .A(n9260), .B(n9305), .Z(n9308) );
  AND U9330 ( .A(n9309), .B(n9310), .Z(n9260) );
  XNOR U9331 ( .A(n9257), .B(n9305), .Z(n9307) );
  XNOR U9332 ( .A(n9311), .B(n9312), .Z(n9257) );
  AND U9333 ( .A(n287), .B(n9313), .Z(n9312) );
  XNOR U9334 ( .A(n9314), .B(n9315), .Z(n9313) );
  XOR U9335 ( .A(n9316), .B(n9317), .Z(n9305) );
  AND U9336 ( .A(n9318), .B(n9319), .Z(n9317) );
  XNOR U9337 ( .A(n9316), .B(n9309), .Z(n9319) );
  IV U9338 ( .A(n9270), .Z(n9309) );
  XOR U9339 ( .A(n9320), .B(n9321), .Z(n9270) );
  XOR U9340 ( .A(n9322), .B(n9310), .Z(n9321) );
  AND U9341 ( .A(n9280), .B(n9323), .Z(n9310) );
  AND U9342 ( .A(n9324), .B(n9325), .Z(n9322) );
  XOR U9343 ( .A(n9326), .B(n9320), .Z(n9324) );
  XNOR U9344 ( .A(n9267), .B(n9316), .Z(n9318) );
  XNOR U9345 ( .A(n9327), .B(n9328), .Z(n9267) );
  AND U9346 ( .A(n287), .B(n9329), .Z(n9328) );
  XNOR U9347 ( .A(n9330), .B(n9331), .Z(n9329) );
  XOR U9348 ( .A(n9332), .B(n9333), .Z(n9316) );
  AND U9349 ( .A(n9334), .B(n9335), .Z(n9333) );
  XNOR U9350 ( .A(n9332), .B(n9280), .Z(n9335) );
  XOR U9351 ( .A(n9336), .B(n9325), .Z(n9280) );
  XNOR U9352 ( .A(n9337), .B(n9320), .Z(n9325) );
  XOR U9353 ( .A(n9338), .B(n9339), .Z(n9320) );
  AND U9354 ( .A(n9340), .B(n9341), .Z(n9339) );
  XOR U9355 ( .A(n9342), .B(n9338), .Z(n9340) );
  XNOR U9356 ( .A(n9343), .B(n9344), .Z(n9337) );
  AND U9357 ( .A(n9345), .B(n9346), .Z(n9344) );
  XOR U9358 ( .A(n9343), .B(n9347), .Z(n9345) );
  XNOR U9359 ( .A(n9326), .B(n9323), .Z(n9336) );
  AND U9360 ( .A(n9348), .B(n9349), .Z(n9323) );
  XOR U9361 ( .A(n9350), .B(n9351), .Z(n9326) );
  AND U9362 ( .A(n9352), .B(n9353), .Z(n9351) );
  XOR U9363 ( .A(n9350), .B(n9354), .Z(n9352) );
  XNOR U9364 ( .A(n9277), .B(n9332), .Z(n9334) );
  XNOR U9365 ( .A(n9355), .B(n9356), .Z(n9277) );
  AND U9366 ( .A(n287), .B(n9357), .Z(n9356) );
  XNOR U9367 ( .A(n9358), .B(n9359), .Z(n9357) );
  XOR U9368 ( .A(n9360), .B(n9361), .Z(n9332) );
  AND U9369 ( .A(n9362), .B(n9363), .Z(n9361) );
  XNOR U9370 ( .A(n9360), .B(n9348), .Z(n9363) );
  IV U9371 ( .A(n9290), .Z(n9348) );
  XNOR U9372 ( .A(n9364), .B(n9341), .Z(n9290) );
  XNOR U9373 ( .A(n9365), .B(n9347), .Z(n9341) );
  XOR U9374 ( .A(n9366), .B(n9367), .Z(n9347) );
  AND U9375 ( .A(n9368), .B(n9369), .Z(n9367) );
  XOR U9376 ( .A(n9366), .B(n9370), .Z(n9368) );
  XNOR U9377 ( .A(n9346), .B(n9338), .Z(n9365) );
  XOR U9378 ( .A(n9371), .B(n9372), .Z(n9338) );
  AND U9379 ( .A(n9373), .B(n9374), .Z(n9372) );
  XNOR U9380 ( .A(n9375), .B(n9371), .Z(n9373) );
  XNOR U9381 ( .A(n9376), .B(n9343), .Z(n9346) );
  XOR U9382 ( .A(n9377), .B(n9378), .Z(n9343) );
  AND U9383 ( .A(n9379), .B(n9380), .Z(n9378) );
  XOR U9384 ( .A(n9377), .B(n9381), .Z(n9379) );
  XNOR U9385 ( .A(n9382), .B(n9383), .Z(n9376) );
  AND U9386 ( .A(n9384), .B(n9385), .Z(n9383) );
  XNOR U9387 ( .A(n9382), .B(n9386), .Z(n9384) );
  XNOR U9388 ( .A(n9342), .B(n9349), .Z(n9364) );
  AND U9389 ( .A(n9298), .B(n9387), .Z(n9349) );
  XOR U9390 ( .A(n9354), .B(n9353), .Z(n9342) );
  XNOR U9391 ( .A(n9388), .B(n9350), .Z(n9353) );
  XOR U9392 ( .A(n9389), .B(n9390), .Z(n9350) );
  AND U9393 ( .A(n9391), .B(n9392), .Z(n9390) );
  XOR U9394 ( .A(n9389), .B(n9393), .Z(n9391) );
  XNOR U9395 ( .A(n9394), .B(n9395), .Z(n9388) );
  AND U9396 ( .A(n9396), .B(n9397), .Z(n9395) );
  XOR U9397 ( .A(n9394), .B(n9398), .Z(n9396) );
  XOR U9398 ( .A(n9399), .B(n9400), .Z(n9354) );
  AND U9399 ( .A(n9401), .B(n9402), .Z(n9400) );
  XOR U9400 ( .A(n9399), .B(n9403), .Z(n9401) );
  XNOR U9401 ( .A(n9287), .B(n9360), .Z(n9362) );
  XNOR U9402 ( .A(n9404), .B(n9405), .Z(n9287) );
  AND U9403 ( .A(n287), .B(n9406), .Z(n9405) );
  XNOR U9404 ( .A(n9407), .B(n9408), .Z(n9406) );
  XOR U9405 ( .A(n9409), .B(n9410), .Z(n9360) );
  AND U9406 ( .A(n9411), .B(n9412), .Z(n9410) );
  XNOR U9407 ( .A(n9409), .B(n9298), .Z(n9412) );
  XOR U9408 ( .A(n9413), .B(n9374), .Z(n9298) );
  XNOR U9409 ( .A(n9414), .B(n9381), .Z(n9374) );
  XOR U9410 ( .A(n9370), .B(n9369), .Z(n9381) );
  XNOR U9411 ( .A(n9415), .B(n9366), .Z(n9369) );
  XOR U9412 ( .A(n9416), .B(n9417), .Z(n9366) );
  AND U9413 ( .A(n9418), .B(n9419), .Z(n9417) );
  XNOR U9414 ( .A(n9420), .B(n9421), .Z(n9418) );
  IV U9415 ( .A(n9416), .Z(n9420) );
  XNOR U9416 ( .A(n9422), .B(n9423), .Z(n9415) );
  NOR U9417 ( .A(n9424), .B(n9425), .Z(n9423) );
  XNOR U9418 ( .A(n9422), .B(n9426), .Z(n9424) );
  XOR U9419 ( .A(n9427), .B(n9428), .Z(n9370) );
  NOR U9420 ( .A(n9429), .B(n9430), .Z(n9428) );
  XNOR U9421 ( .A(n9427), .B(n9431), .Z(n9429) );
  XNOR U9422 ( .A(n9380), .B(n9371), .Z(n9414) );
  XOR U9423 ( .A(n9432), .B(n9433), .Z(n9371) );
  AND U9424 ( .A(n9434), .B(n9435), .Z(n9433) );
  XOR U9425 ( .A(n9432), .B(n9436), .Z(n9434) );
  XOR U9426 ( .A(n9437), .B(n9386), .Z(n9380) );
  XOR U9427 ( .A(n9438), .B(n9439), .Z(n9386) );
  NOR U9428 ( .A(n9440), .B(n9441), .Z(n9439) );
  XOR U9429 ( .A(n9438), .B(n9442), .Z(n9440) );
  XNOR U9430 ( .A(n9385), .B(n9377), .Z(n9437) );
  XOR U9431 ( .A(n9443), .B(n9444), .Z(n9377) );
  AND U9432 ( .A(n9445), .B(n9446), .Z(n9444) );
  XOR U9433 ( .A(n9443), .B(n9447), .Z(n9445) );
  XNOR U9434 ( .A(n9448), .B(n9382), .Z(n9385) );
  XOR U9435 ( .A(n9449), .B(n9450), .Z(n9382) );
  AND U9436 ( .A(n9451), .B(n9452), .Z(n9450) );
  XNOR U9437 ( .A(n9453), .B(n9454), .Z(n9451) );
  IV U9438 ( .A(n9449), .Z(n9453) );
  XNOR U9439 ( .A(n9455), .B(n9456), .Z(n9448) );
  NOR U9440 ( .A(n9457), .B(n9458), .Z(n9456) );
  XNOR U9441 ( .A(n9455), .B(n9459), .Z(n9457) );
  XOR U9442 ( .A(n9375), .B(n9387), .Z(n9413) );
  NOR U9443 ( .A(n9304), .B(n9460), .Z(n9387) );
  XNOR U9444 ( .A(n9393), .B(n9392), .Z(n9375) );
  XNOR U9445 ( .A(n9461), .B(n9398), .Z(n9392) );
  XNOR U9446 ( .A(n9462), .B(n9463), .Z(n9398) );
  NOR U9447 ( .A(n9464), .B(n9465), .Z(n9463) );
  XOR U9448 ( .A(n9462), .B(n9466), .Z(n9464) );
  XNOR U9449 ( .A(n9397), .B(n9389), .Z(n9461) );
  XOR U9450 ( .A(n9467), .B(n9468), .Z(n9389) );
  AND U9451 ( .A(n9469), .B(n9470), .Z(n9468) );
  XOR U9452 ( .A(n9467), .B(n9471), .Z(n9469) );
  XNOR U9453 ( .A(n9472), .B(n9394), .Z(n9397) );
  XOR U9454 ( .A(n9473), .B(n9474), .Z(n9394) );
  AND U9455 ( .A(n9475), .B(n9476), .Z(n9474) );
  XNOR U9456 ( .A(n9477), .B(n9478), .Z(n9475) );
  IV U9457 ( .A(n9473), .Z(n9477) );
  XNOR U9458 ( .A(n9479), .B(n9480), .Z(n9472) );
  NOR U9459 ( .A(n9481), .B(n9482), .Z(n9480) );
  XNOR U9460 ( .A(n9479), .B(n9483), .Z(n9481) );
  XOR U9461 ( .A(n9403), .B(n9402), .Z(n9393) );
  XNOR U9462 ( .A(n9484), .B(n9399), .Z(n9402) );
  XOR U9463 ( .A(n9485), .B(n9486), .Z(n9399) );
  AND U9464 ( .A(n9487), .B(n9488), .Z(n9486) );
  XNOR U9465 ( .A(n9489), .B(n9490), .Z(n9487) );
  IV U9466 ( .A(n9485), .Z(n9489) );
  XNOR U9467 ( .A(n9491), .B(n9492), .Z(n9484) );
  NOR U9468 ( .A(n9493), .B(n9494), .Z(n9492) );
  XNOR U9469 ( .A(n9491), .B(n9495), .Z(n9493) );
  XOR U9470 ( .A(n9496), .B(n9497), .Z(n9403) );
  NOR U9471 ( .A(n9498), .B(n9499), .Z(n9497) );
  XNOR U9472 ( .A(n9496), .B(n9500), .Z(n9498) );
  XNOR U9473 ( .A(n9295), .B(n9409), .Z(n9411) );
  XNOR U9474 ( .A(n9501), .B(n9502), .Z(n9295) );
  AND U9475 ( .A(n287), .B(n9503), .Z(n9502) );
  XNOR U9476 ( .A(n9504), .B(n9505), .Z(n9503) );
  AND U9477 ( .A(n9301), .B(n9304), .Z(n9409) );
  XOR U9478 ( .A(n9506), .B(n9460), .Z(n9304) );
  XNOR U9479 ( .A(p_input[256]), .B(p_input[512]), .Z(n9460) );
  XNOR U9480 ( .A(n9436), .B(n9435), .Z(n9506) );
  XNOR U9481 ( .A(n9507), .B(n9447), .Z(n9435) );
  XOR U9482 ( .A(n9421), .B(n9419), .Z(n9447) );
  XNOR U9483 ( .A(n9508), .B(n9426), .Z(n9419) );
  XOR U9484 ( .A(p_input[280]), .B(p_input[536]), .Z(n9426) );
  XOR U9485 ( .A(n9416), .B(n9425), .Z(n9508) );
  XOR U9486 ( .A(n9509), .B(n9422), .Z(n9425) );
  XOR U9487 ( .A(p_input[278]), .B(p_input[534]), .Z(n9422) );
  XOR U9488 ( .A(p_input[279]), .B(n6576), .Z(n9509) );
  XOR U9489 ( .A(p_input[274]), .B(p_input[530]), .Z(n9416) );
  XNOR U9490 ( .A(n9431), .B(n9430), .Z(n9421) );
  XOR U9491 ( .A(n9510), .B(n9427), .Z(n9430) );
  XOR U9492 ( .A(p_input[275]), .B(p_input[531]), .Z(n9427) );
  XOR U9493 ( .A(p_input[276]), .B(n6578), .Z(n9510) );
  XOR U9494 ( .A(p_input[277]), .B(p_input[533]), .Z(n9431) );
  XOR U9495 ( .A(n9446), .B(n9511), .Z(n9507) );
  IV U9496 ( .A(n9432), .Z(n9511) );
  XOR U9497 ( .A(p_input[257]), .B(p_input[513]), .Z(n9432) );
  XNOR U9498 ( .A(n9512), .B(n9454), .Z(n9446) );
  XNOR U9499 ( .A(n9442), .B(n9441), .Z(n9454) );
  XNOR U9500 ( .A(n9513), .B(n9438), .Z(n9441) );
  XNOR U9501 ( .A(p_input[282]), .B(p_input[538]), .Z(n9438) );
  XOR U9502 ( .A(p_input[283]), .B(n6582), .Z(n9513) );
  XOR U9503 ( .A(p_input[284]), .B(p_input[540]), .Z(n9442) );
  XOR U9504 ( .A(n9452), .B(n9514), .Z(n9512) );
  IV U9505 ( .A(n9443), .Z(n9514) );
  XOR U9506 ( .A(p_input[273]), .B(p_input[529]), .Z(n9443) );
  XNOR U9507 ( .A(n9515), .B(n9459), .Z(n9452) );
  XNOR U9508 ( .A(p_input[287]), .B(n6585), .Z(n9459) );
  XOR U9509 ( .A(n9449), .B(n9458), .Z(n9515) );
  XOR U9510 ( .A(n9516), .B(n9455), .Z(n9458) );
  XOR U9511 ( .A(p_input[285]), .B(p_input[541]), .Z(n9455) );
  XOR U9512 ( .A(p_input[286]), .B(n6587), .Z(n9516) );
  XOR U9513 ( .A(p_input[281]), .B(p_input[537]), .Z(n9449) );
  XOR U9514 ( .A(n9471), .B(n9470), .Z(n9436) );
  XNOR U9515 ( .A(n9517), .B(n9478), .Z(n9470) );
  XNOR U9516 ( .A(n9466), .B(n9465), .Z(n9478) );
  XNOR U9517 ( .A(n9518), .B(n9462), .Z(n9465) );
  XNOR U9518 ( .A(p_input[267]), .B(p_input[523]), .Z(n9462) );
  XOR U9519 ( .A(p_input[268]), .B(n6590), .Z(n9518) );
  XOR U9520 ( .A(p_input[269]), .B(p_input[525]), .Z(n9466) );
  XOR U9521 ( .A(n9476), .B(n9519), .Z(n9517) );
  IV U9522 ( .A(n9467), .Z(n9519) );
  XOR U9523 ( .A(p_input[258]), .B(p_input[514]), .Z(n9467) );
  XNOR U9524 ( .A(n9520), .B(n9483), .Z(n9476) );
  XNOR U9525 ( .A(p_input[272]), .B(n6593), .Z(n9483) );
  XOR U9526 ( .A(n9473), .B(n9482), .Z(n9520) );
  XOR U9527 ( .A(n9521), .B(n9479), .Z(n9482) );
  XOR U9528 ( .A(p_input[270]), .B(p_input[526]), .Z(n9479) );
  XOR U9529 ( .A(p_input[271]), .B(n6595), .Z(n9521) );
  XOR U9530 ( .A(p_input[266]), .B(p_input[522]), .Z(n9473) );
  XOR U9531 ( .A(n9490), .B(n9488), .Z(n9471) );
  XNOR U9532 ( .A(n9522), .B(n9495), .Z(n9488) );
  XOR U9533 ( .A(p_input[265]), .B(p_input[521]), .Z(n9495) );
  XOR U9534 ( .A(n9485), .B(n9494), .Z(n9522) );
  XOR U9535 ( .A(n9523), .B(n9491), .Z(n9494) );
  XOR U9536 ( .A(p_input[263]), .B(p_input[519]), .Z(n9491) );
  XOR U9537 ( .A(p_input[264]), .B(n6963), .Z(n9523) );
  XOR U9538 ( .A(p_input[259]), .B(p_input[515]), .Z(n9485) );
  XNOR U9539 ( .A(n9500), .B(n9499), .Z(n9490) );
  XOR U9540 ( .A(n9524), .B(n9496), .Z(n9499) );
  XOR U9541 ( .A(p_input[260]), .B(p_input[516]), .Z(n9496) );
  XOR U9542 ( .A(p_input[261]), .B(n6965), .Z(n9524) );
  XOR U9543 ( .A(p_input[262]), .B(p_input[518]), .Z(n9500) );
  XNOR U9544 ( .A(n9525), .B(n9526), .Z(n9301) );
  AND U9545 ( .A(n287), .B(n9527), .Z(n9526) );
  XNOR U9546 ( .A(n9528), .B(n9529), .Z(n287) );
  AND U9547 ( .A(n9530), .B(n9531), .Z(n9529) );
  XOR U9548 ( .A(n9315), .B(n9528), .Z(n9531) );
  XNOR U9549 ( .A(n9532), .B(n9528), .Z(n9530) );
  XOR U9550 ( .A(n9533), .B(n9534), .Z(n9528) );
  AND U9551 ( .A(n9535), .B(n9536), .Z(n9534) );
  XOR U9552 ( .A(n9330), .B(n9533), .Z(n9536) );
  XOR U9553 ( .A(n9533), .B(n9331), .Z(n9535) );
  XOR U9554 ( .A(n9537), .B(n9538), .Z(n9533) );
  AND U9555 ( .A(n9539), .B(n9540), .Z(n9538) );
  XOR U9556 ( .A(n9358), .B(n9537), .Z(n9540) );
  XOR U9557 ( .A(n9537), .B(n9359), .Z(n9539) );
  XOR U9558 ( .A(n9541), .B(n9542), .Z(n9537) );
  AND U9559 ( .A(n9543), .B(n9544), .Z(n9542) );
  XOR U9560 ( .A(n9407), .B(n9541), .Z(n9544) );
  XOR U9561 ( .A(n9541), .B(n9408), .Z(n9543) );
  XOR U9562 ( .A(n9545), .B(n9546), .Z(n9541) );
  AND U9563 ( .A(n9547), .B(n9548), .Z(n9546) );
  XOR U9564 ( .A(n9545), .B(n9504), .Z(n9548) );
  XNOR U9565 ( .A(n9549), .B(n9550), .Z(n9251) );
  AND U9566 ( .A(n291), .B(n9551), .Z(n9550) );
  XNOR U9567 ( .A(n9552), .B(n9553), .Z(n291) );
  AND U9568 ( .A(n9554), .B(n9555), .Z(n9553) );
  XOR U9569 ( .A(n9552), .B(n9261), .Z(n9555) );
  XNOR U9570 ( .A(n9552), .B(n9211), .Z(n9554) );
  XOR U9571 ( .A(n9556), .B(n9557), .Z(n9552) );
  AND U9572 ( .A(n9558), .B(n9559), .Z(n9557) );
  XNOR U9573 ( .A(n9271), .B(n9556), .Z(n9559) );
  XOR U9574 ( .A(n9556), .B(n9221), .Z(n9558) );
  XOR U9575 ( .A(n9560), .B(n9561), .Z(n9556) );
  AND U9576 ( .A(n9562), .B(n9563), .Z(n9561) );
  XNOR U9577 ( .A(n9281), .B(n9560), .Z(n9563) );
  XOR U9578 ( .A(n9560), .B(n9230), .Z(n9562) );
  XOR U9579 ( .A(n9564), .B(n9565), .Z(n9560) );
  AND U9580 ( .A(n9566), .B(n9567), .Z(n9565) );
  XOR U9581 ( .A(n9564), .B(n9238), .Z(n9566) );
  XOR U9582 ( .A(n9568), .B(n9569), .Z(n9202) );
  AND U9583 ( .A(n295), .B(n9551), .Z(n9569) );
  XNOR U9584 ( .A(n9549), .B(n9568), .Z(n9551) );
  XNOR U9585 ( .A(n9570), .B(n9571), .Z(n295) );
  AND U9586 ( .A(n9572), .B(n9573), .Z(n9571) );
  XNOR U9587 ( .A(n9574), .B(n9570), .Z(n9573) );
  IV U9588 ( .A(n9261), .Z(n9574) );
  XOR U9589 ( .A(n9532), .B(n9575), .Z(n9261) );
  AND U9590 ( .A(n298), .B(n9576), .Z(n9575) );
  XOR U9591 ( .A(n9314), .B(n9311), .Z(n9576) );
  XNOR U9592 ( .A(n9211), .B(n9570), .Z(n9572) );
  XNOR U9593 ( .A(n9577), .B(n9578), .Z(n9211) );
  AND U9594 ( .A(n314), .B(n9579), .Z(n9578) );
  XNOR U9595 ( .A(n9580), .B(n9581), .Z(n9579) );
  XOR U9596 ( .A(n9582), .B(n9583), .Z(n9570) );
  AND U9597 ( .A(n9584), .B(n9585), .Z(n9583) );
  XNOR U9598 ( .A(n9582), .B(n9271), .Z(n9585) );
  XOR U9599 ( .A(n9331), .B(n9586), .Z(n9271) );
  AND U9600 ( .A(n298), .B(n9587), .Z(n9586) );
  XOR U9601 ( .A(n9327), .B(n9331), .Z(n9587) );
  XNOR U9602 ( .A(n9588), .B(n9582), .Z(n9584) );
  IV U9603 ( .A(n9221), .Z(n9588) );
  XOR U9604 ( .A(n9589), .B(n9590), .Z(n9221) );
  AND U9605 ( .A(n314), .B(n9591), .Z(n9590) );
  XOR U9606 ( .A(n9592), .B(n9593), .Z(n9582) );
  AND U9607 ( .A(n9594), .B(n9595), .Z(n9593) );
  XNOR U9608 ( .A(n9592), .B(n9281), .Z(n9595) );
  XOR U9609 ( .A(n9359), .B(n9596), .Z(n9281) );
  AND U9610 ( .A(n298), .B(n9597), .Z(n9596) );
  XOR U9611 ( .A(n9355), .B(n9359), .Z(n9597) );
  XOR U9612 ( .A(n9230), .B(n9592), .Z(n9594) );
  XOR U9613 ( .A(n9598), .B(n9599), .Z(n9230) );
  AND U9614 ( .A(n314), .B(n9600), .Z(n9599) );
  XOR U9615 ( .A(n9564), .B(n9601), .Z(n9592) );
  AND U9616 ( .A(n9602), .B(n9567), .Z(n9601) );
  XNOR U9617 ( .A(n9291), .B(n9564), .Z(n9567) );
  XOR U9618 ( .A(n9408), .B(n9603), .Z(n9291) );
  AND U9619 ( .A(n298), .B(n9604), .Z(n9603) );
  XOR U9620 ( .A(n9404), .B(n9408), .Z(n9604) );
  XNOR U9621 ( .A(n9605), .B(n9564), .Z(n9602) );
  IV U9622 ( .A(n9238), .Z(n9605) );
  XOR U9623 ( .A(n9606), .B(n9607), .Z(n9238) );
  AND U9624 ( .A(n314), .B(n9608), .Z(n9607) );
  XOR U9625 ( .A(n9609), .B(n9610), .Z(n9564) );
  AND U9626 ( .A(n9611), .B(n9612), .Z(n9610) );
  XNOR U9627 ( .A(n9609), .B(n9299), .Z(n9612) );
  XOR U9628 ( .A(n9505), .B(n9613), .Z(n9299) );
  AND U9629 ( .A(n298), .B(n9614), .Z(n9613) );
  XOR U9630 ( .A(n9501), .B(n9505), .Z(n9614) );
  XNOR U9631 ( .A(n9615), .B(n9609), .Z(n9611) );
  IV U9632 ( .A(n9248), .Z(n9615) );
  XOR U9633 ( .A(n9616), .B(n9617), .Z(n9248) );
  AND U9634 ( .A(n314), .B(n9618), .Z(n9617) );
  AND U9635 ( .A(n9568), .B(n9549), .Z(n9609) );
  XNOR U9636 ( .A(n9619), .B(n9620), .Z(n9549) );
  AND U9637 ( .A(n298), .B(n9527), .Z(n9620) );
  XNOR U9638 ( .A(n9525), .B(n9619), .Z(n9527) );
  XNOR U9639 ( .A(n9621), .B(n9622), .Z(n298) );
  AND U9640 ( .A(n9623), .B(n9624), .Z(n9622) );
  XNOR U9641 ( .A(n9621), .B(n9311), .Z(n9624) );
  IV U9642 ( .A(n9315), .Z(n9311) );
  XOR U9643 ( .A(n9625), .B(n9626), .Z(n9315) );
  AND U9644 ( .A(n302), .B(n9627), .Z(n9626) );
  XOR U9645 ( .A(n9628), .B(n9625), .Z(n9627) );
  XNOR U9646 ( .A(n9621), .B(n9532), .Z(n9623) );
  IV U9647 ( .A(n9314), .Z(n9532) );
  XOR U9648 ( .A(n9580), .B(n9629), .Z(n9314) );
  AND U9649 ( .A(n310), .B(n9630), .Z(n9629) );
  XOR U9650 ( .A(n9580), .B(n9577), .Z(n9630) );
  XOR U9651 ( .A(n9631), .B(n9632), .Z(n9621) );
  AND U9652 ( .A(n9633), .B(n9634), .Z(n9632) );
  XNOR U9653 ( .A(n9631), .B(n9327), .Z(n9634) );
  IV U9654 ( .A(n9330), .Z(n9327) );
  XOR U9655 ( .A(n9635), .B(n9636), .Z(n9330) );
  AND U9656 ( .A(n302), .B(n9637), .Z(n9636) );
  XOR U9657 ( .A(n9638), .B(n9635), .Z(n9637) );
  XOR U9658 ( .A(n9331), .B(n9631), .Z(n9633) );
  XOR U9659 ( .A(n9639), .B(n9640), .Z(n9331) );
  AND U9660 ( .A(n310), .B(n9591), .Z(n9640) );
  XOR U9661 ( .A(n9639), .B(n9589), .Z(n9591) );
  XOR U9662 ( .A(n9641), .B(n9642), .Z(n9631) );
  AND U9663 ( .A(n9643), .B(n9644), .Z(n9642) );
  XNOR U9664 ( .A(n9641), .B(n9355), .Z(n9644) );
  IV U9665 ( .A(n9358), .Z(n9355) );
  XOR U9666 ( .A(n9645), .B(n9646), .Z(n9358) );
  AND U9667 ( .A(n302), .B(n9647), .Z(n9646) );
  XNOR U9668 ( .A(n9648), .B(n9645), .Z(n9647) );
  XOR U9669 ( .A(n9359), .B(n9641), .Z(n9643) );
  XOR U9670 ( .A(n9649), .B(n9650), .Z(n9359) );
  AND U9671 ( .A(n310), .B(n9600), .Z(n9650) );
  XOR U9672 ( .A(n9649), .B(n9598), .Z(n9600) );
  XOR U9673 ( .A(n9651), .B(n9652), .Z(n9641) );
  AND U9674 ( .A(n9653), .B(n9654), .Z(n9652) );
  XNOR U9675 ( .A(n9651), .B(n9404), .Z(n9654) );
  IV U9676 ( .A(n9407), .Z(n9404) );
  XOR U9677 ( .A(n9655), .B(n9656), .Z(n9407) );
  AND U9678 ( .A(n302), .B(n9657), .Z(n9656) );
  XOR U9679 ( .A(n9658), .B(n9655), .Z(n9657) );
  XOR U9680 ( .A(n9408), .B(n9651), .Z(n9653) );
  XOR U9681 ( .A(n9659), .B(n9660), .Z(n9408) );
  AND U9682 ( .A(n310), .B(n9608), .Z(n9660) );
  XOR U9683 ( .A(n9659), .B(n9606), .Z(n9608) );
  XOR U9684 ( .A(n9545), .B(n9661), .Z(n9651) );
  AND U9685 ( .A(n9547), .B(n9662), .Z(n9661) );
  XNOR U9686 ( .A(n9545), .B(n9501), .Z(n9662) );
  IV U9687 ( .A(n9504), .Z(n9501) );
  XOR U9688 ( .A(n9663), .B(n9664), .Z(n9504) );
  AND U9689 ( .A(n302), .B(n9665), .Z(n9664) );
  XNOR U9690 ( .A(n9666), .B(n9663), .Z(n9665) );
  XOR U9691 ( .A(n9505), .B(n9545), .Z(n9547) );
  XOR U9692 ( .A(n9667), .B(n9668), .Z(n9505) );
  AND U9693 ( .A(n310), .B(n9618), .Z(n9668) );
  XOR U9694 ( .A(n9667), .B(n9616), .Z(n9618) );
  AND U9695 ( .A(n9619), .B(n9525), .Z(n9545) );
  XNOR U9696 ( .A(n9669), .B(n9670), .Z(n9525) );
  AND U9697 ( .A(n302), .B(n9671), .Z(n9670) );
  XNOR U9698 ( .A(n9672), .B(n9669), .Z(n9671) );
  XNOR U9699 ( .A(n9673), .B(n9674), .Z(n302) );
  AND U9700 ( .A(n9675), .B(n9676), .Z(n9674) );
  XOR U9701 ( .A(n9628), .B(n9673), .Z(n9676) );
  AND U9702 ( .A(n9677), .B(n9678), .Z(n9628) );
  XNOR U9703 ( .A(n9625), .B(n9673), .Z(n9675) );
  XNOR U9704 ( .A(n9679), .B(n9680), .Z(n9625) );
  AND U9705 ( .A(n9681), .B(n306), .Z(n9680) );
  XOR U9706 ( .A(n9682), .B(n9683), .Z(n9673) );
  AND U9707 ( .A(n9684), .B(n9685), .Z(n9683) );
  XNOR U9708 ( .A(n9682), .B(n9677), .Z(n9685) );
  IV U9709 ( .A(n9638), .Z(n9677) );
  XOR U9710 ( .A(n9686), .B(n9687), .Z(n9638) );
  XOR U9711 ( .A(n9688), .B(n9678), .Z(n9687) );
  AND U9712 ( .A(n9648), .B(n9689), .Z(n9678) );
  AND U9713 ( .A(n9690), .B(n9691), .Z(n9688) );
  XOR U9714 ( .A(n9692), .B(n9686), .Z(n9690) );
  XNOR U9715 ( .A(n9635), .B(n9682), .Z(n9684) );
  XNOR U9716 ( .A(n9693), .B(n9694), .Z(n9635) );
  AND U9717 ( .A(n306), .B(n9695), .Z(n9694) );
  XNOR U9718 ( .A(n9696), .B(n9697), .Z(n9695) );
  XOR U9719 ( .A(n9698), .B(n9699), .Z(n9682) );
  AND U9720 ( .A(n9700), .B(n9701), .Z(n9699) );
  XNOR U9721 ( .A(n9698), .B(n9648), .Z(n9701) );
  XOR U9722 ( .A(n9702), .B(n9691), .Z(n9648) );
  XNOR U9723 ( .A(n9703), .B(n9686), .Z(n9691) );
  XOR U9724 ( .A(n9704), .B(n9705), .Z(n9686) );
  AND U9725 ( .A(n9706), .B(n9707), .Z(n9705) );
  XOR U9726 ( .A(n9708), .B(n9704), .Z(n9706) );
  XNOR U9727 ( .A(n9709), .B(n9710), .Z(n9703) );
  AND U9728 ( .A(n9711), .B(n9712), .Z(n9710) );
  XOR U9729 ( .A(n9709), .B(n9713), .Z(n9711) );
  XNOR U9730 ( .A(n9692), .B(n9689), .Z(n9702) );
  AND U9731 ( .A(n9714), .B(n9715), .Z(n9689) );
  XOR U9732 ( .A(n9716), .B(n9717), .Z(n9692) );
  AND U9733 ( .A(n9718), .B(n9719), .Z(n9717) );
  XOR U9734 ( .A(n9716), .B(n9720), .Z(n9718) );
  XNOR U9735 ( .A(n9645), .B(n9698), .Z(n9700) );
  XNOR U9736 ( .A(n9721), .B(n9722), .Z(n9645) );
  AND U9737 ( .A(n306), .B(n9723), .Z(n9722) );
  XNOR U9738 ( .A(n9724), .B(n9725), .Z(n9723) );
  XOR U9739 ( .A(n9726), .B(n9727), .Z(n9698) );
  AND U9740 ( .A(n9728), .B(n9729), .Z(n9727) );
  XNOR U9741 ( .A(n9726), .B(n9714), .Z(n9729) );
  IV U9742 ( .A(n9658), .Z(n9714) );
  XNOR U9743 ( .A(n9730), .B(n9707), .Z(n9658) );
  XNOR U9744 ( .A(n9731), .B(n9713), .Z(n9707) );
  XOR U9745 ( .A(n9732), .B(n9733), .Z(n9713) );
  AND U9746 ( .A(n9734), .B(n9735), .Z(n9733) );
  XOR U9747 ( .A(n9732), .B(n9736), .Z(n9734) );
  XNOR U9748 ( .A(n9712), .B(n9704), .Z(n9731) );
  XOR U9749 ( .A(n9737), .B(n9738), .Z(n9704) );
  AND U9750 ( .A(n9739), .B(n9740), .Z(n9738) );
  XNOR U9751 ( .A(n9741), .B(n9737), .Z(n9739) );
  XNOR U9752 ( .A(n9742), .B(n9709), .Z(n9712) );
  XOR U9753 ( .A(n9743), .B(n9744), .Z(n9709) );
  AND U9754 ( .A(n9745), .B(n9746), .Z(n9744) );
  XOR U9755 ( .A(n9743), .B(n9747), .Z(n9745) );
  XNOR U9756 ( .A(n9748), .B(n9749), .Z(n9742) );
  AND U9757 ( .A(n9750), .B(n9751), .Z(n9749) );
  XNOR U9758 ( .A(n9748), .B(n9752), .Z(n9750) );
  XNOR U9759 ( .A(n9708), .B(n9715), .Z(n9730) );
  AND U9760 ( .A(n9666), .B(n9753), .Z(n9715) );
  XOR U9761 ( .A(n9720), .B(n9719), .Z(n9708) );
  XNOR U9762 ( .A(n9754), .B(n9716), .Z(n9719) );
  XOR U9763 ( .A(n9755), .B(n9756), .Z(n9716) );
  AND U9764 ( .A(n9757), .B(n9758), .Z(n9756) );
  XOR U9765 ( .A(n9755), .B(n9759), .Z(n9757) );
  XNOR U9766 ( .A(n9760), .B(n9761), .Z(n9754) );
  AND U9767 ( .A(n9762), .B(n9763), .Z(n9761) );
  XOR U9768 ( .A(n9760), .B(n9764), .Z(n9762) );
  XOR U9769 ( .A(n9765), .B(n9766), .Z(n9720) );
  AND U9770 ( .A(n9767), .B(n9768), .Z(n9766) );
  XOR U9771 ( .A(n9765), .B(n9769), .Z(n9767) );
  XNOR U9772 ( .A(n9655), .B(n9726), .Z(n9728) );
  XNOR U9773 ( .A(n9770), .B(n9771), .Z(n9655) );
  AND U9774 ( .A(n306), .B(n9772), .Z(n9771) );
  XNOR U9775 ( .A(n9773), .B(n9774), .Z(n9772) );
  XOR U9776 ( .A(n9775), .B(n9776), .Z(n9726) );
  AND U9777 ( .A(n9777), .B(n9778), .Z(n9776) );
  XNOR U9778 ( .A(n9775), .B(n9666), .Z(n9778) );
  XOR U9779 ( .A(n9779), .B(n9740), .Z(n9666) );
  XNOR U9780 ( .A(n9780), .B(n9747), .Z(n9740) );
  XOR U9781 ( .A(n9736), .B(n9735), .Z(n9747) );
  XNOR U9782 ( .A(n9781), .B(n9732), .Z(n9735) );
  XOR U9783 ( .A(n9782), .B(n9783), .Z(n9732) );
  AND U9784 ( .A(n9784), .B(n9785), .Z(n9783) );
  XNOR U9785 ( .A(n9786), .B(n9787), .Z(n9784) );
  IV U9786 ( .A(n9782), .Z(n9786) );
  XNOR U9787 ( .A(n9788), .B(n9789), .Z(n9781) );
  NOR U9788 ( .A(n9790), .B(n9791), .Z(n9789) );
  XNOR U9789 ( .A(n9788), .B(n9792), .Z(n9790) );
  XOR U9790 ( .A(n9793), .B(n9794), .Z(n9736) );
  NOR U9791 ( .A(n9795), .B(n9796), .Z(n9794) );
  XNOR U9792 ( .A(n9793), .B(n9797), .Z(n9795) );
  XNOR U9793 ( .A(n9746), .B(n9737), .Z(n9780) );
  XOR U9794 ( .A(n9798), .B(n9799), .Z(n9737) );
  AND U9795 ( .A(n9800), .B(n9801), .Z(n9799) );
  XOR U9796 ( .A(n9798), .B(n9802), .Z(n9800) );
  XOR U9797 ( .A(n9803), .B(n9752), .Z(n9746) );
  XOR U9798 ( .A(n9804), .B(n9805), .Z(n9752) );
  NOR U9799 ( .A(n9806), .B(n9807), .Z(n9805) );
  XOR U9800 ( .A(n9804), .B(n9808), .Z(n9806) );
  XNOR U9801 ( .A(n9751), .B(n9743), .Z(n9803) );
  XOR U9802 ( .A(n9809), .B(n9810), .Z(n9743) );
  AND U9803 ( .A(n9811), .B(n9812), .Z(n9810) );
  XOR U9804 ( .A(n9809), .B(n9813), .Z(n9811) );
  XNOR U9805 ( .A(n9814), .B(n9748), .Z(n9751) );
  XOR U9806 ( .A(n9815), .B(n9816), .Z(n9748) );
  AND U9807 ( .A(n9817), .B(n9818), .Z(n9816) );
  XNOR U9808 ( .A(n9819), .B(n9820), .Z(n9817) );
  IV U9809 ( .A(n9815), .Z(n9819) );
  XNOR U9810 ( .A(n9821), .B(n9822), .Z(n9814) );
  NOR U9811 ( .A(n9823), .B(n9824), .Z(n9822) );
  XNOR U9812 ( .A(n9821), .B(n9825), .Z(n9823) );
  XOR U9813 ( .A(n9741), .B(n9753), .Z(n9779) );
  NOR U9814 ( .A(n9672), .B(n9826), .Z(n9753) );
  XNOR U9815 ( .A(n9759), .B(n9758), .Z(n9741) );
  XNOR U9816 ( .A(n9827), .B(n9764), .Z(n9758) );
  XNOR U9817 ( .A(n9828), .B(n9829), .Z(n9764) );
  NOR U9818 ( .A(n9830), .B(n9831), .Z(n9829) );
  XOR U9819 ( .A(n9828), .B(n9832), .Z(n9830) );
  XNOR U9820 ( .A(n9763), .B(n9755), .Z(n9827) );
  XOR U9821 ( .A(n9833), .B(n9834), .Z(n9755) );
  AND U9822 ( .A(n9835), .B(n9836), .Z(n9834) );
  XOR U9823 ( .A(n9833), .B(n9837), .Z(n9835) );
  XNOR U9824 ( .A(n9838), .B(n9760), .Z(n9763) );
  XOR U9825 ( .A(n9839), .B(n9840), .Z(n9760) );
  AND U9826 ( .A(n9841), .B(n9842), .Z(n9840) );
  XNOR U9827 ( .A(n9843), .B(n9844), .Z(n9841) );
  IV U9828 ( .A(n9839), .Z(n9843) );
  XNOR U9829 ( .A(n9845), .B(n9846), .Z(n9838) );
  NOR U9830 ( .A(n9847), .B(n9848), .Z(n9846) );
  XNOR U9831 ( .A(n9845), .B(n9849), .Z(n9847) );
  XOR U9832 ( .A(n9769), .B(n9768), .Z(n9759) );
  XNOR U9833 ( .A(n9850), .B(n9765), .Z(n9768) );
  XOR U9834 ( .A(n9851), .B(n9852), .Z(n9765) );
  AND U9835 ( .A(n9853), .B(n9854), .Z(n9852) );
  XNOR U9836 ( .A(n9855), .B(n9856), .Z(n9853) );
  IV U9837 ( .A(n9851), .Z(n9855) );
  XNOR U9838 ( .A(n9857), .B(n9858), .Z(n9850) );
  NOR U9839 ( .A(n9859), .B(n9860), .Z(n9858) );
  XNOR U9840 ( .A(n9857), .B(n9861), .Z(n9859) );
  XOR U9841 ( .A(n9862), .B(n9863), .Z(n9769) );
  NOR U9842 ( .A(n9864), .B(n9865), .Z(n9863) );
  XNOR U9843 ( .A(n9862), .B(n9866), .Z(n9864) );
  XNOR U9844 ( .A(n9663), .B(n9775), .Z(n9777) );
  XNOR U9845 ( .A(n9867), .B(n9868), .Z(n9663) );
  AND U9846 ( .A(n306), .B(n9869), .Z(n9868) );
  XNOR U9847 ( .A(n9870), .B(n9871), .Z(n9869) );
  AND U9848 ( .A(n9669), .B(n9672), .Z(n9775) );
  XOR U9849 ( .A(n9872), .B(n9826), .Z(n9672) );
  XNOR U9850 ( .A(p_input[288]), .B(p_input[512]), .Z(n9826) );
  XNOR U9851 ( .A(n9802), .B(n9801), .Z(n9872) );
  XNOR U9852 ( .A(n9873), .B(n9813), .Z(n9801) );
  XOR U9853 ( .A(n9787), .B(n9785), .Z(n9813) );
  XNOR U9854 ( .A(n9874), .B(n9792), .Z(n9785) );
  XOR U9855 ( .A(p_input[312]), .B(p_input[536]), .Z(n9792) );
  XOR U9856 ( .A(n9782), .B(n9791), .Z(n9874) );
  XOR U9857 ( .A(n9875), .B(n9788), .Z(n9791) );
  XOR U9858 ( .A(p_input[310]), .B(p_input[534]), .Z(n9788) );
  XOR U9859 ( .A(p_input[311]), .B(n6576), .Z(n9875) );
  XOR U9860 ( .A(p_input[306]), .B(p_input[530]), .Z(n9782) );
  XNOR U9861 ( .A(n9797), .B(n9796), .Z(n9787) );
  XOR U9862 ( .A(n9876), .B(n9793), .Z(n9796) );
  XOR U9863 ( .A(p_input[307]), .B(p_input[531]), .Z(n9793) );
  XOR U9864 ( .A(p_input[308]), .B(n6578), .Z(n9876) );
  XOR U9865 ( .A(p_input[309]), .B(p_input[533]), .Z(n9797) );
  XOR U9866 ( .A(n9812), .B(n9877), .Z(n9873) );
  IV U9867 ( .A(n9798), .Z(n9877) );
  XOR U9868 ( .A(p_input[289]), .B(p_input[513]), .Z(n9798) );
  XNOR U9869 ( .A(n9878), .B(n9820), .Z(n9812) );
  XNOR U9870 ( .A(n9808), .B(n9807), .Z(n9820) );
  XNOR U9871 ( .A(n9879), .B(n9804), .Z(n9807) );
  XNOR U9872 ( .A(p_input[314]), .B(p_input[538]), .Z(n9804) );
  XOR U9873 ( .A(p_input[315]), .B(n6582), .Z(n9879) );
  XOR U9874 ( .A(p_input[316]), .B(p_input[540]), .Z(n9808) );
  XOR U9875 ( .A(n9818), .B(n9880), .Z(n9878) );
  IV U9876 ( .A(n9809), .Z(n9880) );
  XOR U9877 ( .A(p_input[305]), .B(p_input[529]), .Z(n9809) );
  XNOR U9878 ( .A(n9881), .B(n9825), .Z(n9818) );
  XNOR U9879 ( .A(p_input[319]), .B(n6585), .Z(n9825) );
  XOR U9880 ( .A(n9815), .B(n9824), .Z(n9881) );
  XOR U9881 ( .A(n9882), .B(n9821), .Z(n9824) );
  XOR U9882 ( .A(p_input[317]), .B(p_input[541]), .Z(n9821) );
  XOR U9883 ( .A(p_input[318]), .B(n6587), .Z(n9882) );
  XOR U9884 ( .A(p_input[313]), .B(p_input[537]), .Z(n9815) );
  XOR U9885 ( .A(n9837), .B(n9836), .Z(n9802) );
  XNOR U9886 ( .A(n9883), .B(n9844), .Z(n9836) );
  XNOR U9887 ( .A(n9832), .B(n9831), .Z(n9844) );
  XNOR U9888 ( .A(n9884), .B(n9828), .Z(n9831) );
  XNOR U9889 ( .A(p_input[299]), .B(p_input[523]), .Z(n9828) );
  XOR U9890 ( .A(p_input[300]), .B(n6590), .Z(n9884) );
  XOR U9891 ( .A(p_input[301]), .B(p_input[525]), .Z(n9832) );
  XOR U9892 ( .A(n9842), .B(n9885), .Z(n9883) );
  IV U9893 ( .A(n9833), .Z(n9885) );
  XOR U9894 ( .A(p_input[290]), .B(p_input[514]), .Z(n9833) );
  XNOR U9895 ( .A(n9886), .B(n9849), .Z(n9842) );
  XNOR U9896 ( .A(p_input[304]), .B(n6593), .Z(n9849) );
  XOR U9897 ( .A(n9839), .B(n9848), .Z(n9886) );
  XOR U9898 ( .A(n9887), .B(n9845), .Z(n9848) );
  XOR U9899 ( .A(p_input[302]), .B(p_input[526]), .Z(n9845) );
  XOR U9900 ( .A(p_input[303]), .B(n6595), .Z(n9887) );
  XOR U9901 ( .A(p_input[298]), .B(p_input[522]), .Z(n9839) );
  XOR U9902 ( .A(n9856), .B(n9854), .Z(n9837) );
  XNOR U9903 ( .A(n9888), .B(n9861), .Z(n9854) );
  XOR U9904 ( .A(p_input[297]), .B(p_input[521]), .Z(n9861) );
  XOR U9905 ( .A(n9851), .B(n9860), .Z(n9888) );
  XOR U9906 ( .A(n9889), .B(n9857), .Z(n9860) );
  XOR U9907 ( .A(p_input[295]), .B(p_input[519]), .Z(n9857) );
  XOR U9908 ( .A(p_input[296]), .B(n6963), .Z(n9889) );
  XOR U9909 ( .A(p_input[291]), .B(p_input[515]), .Z(n9851) );
  XNOR U9910 ( .A(n9866), .B(n9865), .Z(n9856) );
  XOR U9911 ( .A(n9890), .B(n9862), .Z(n9865) );
  XOR U9912 ( .A(p_input[292]), .B(p_input[516]), .Z(n9862) );
  XOR U9913 ( .A(p_input[293]), .B(n6965), .Z(n9890) );
  XOR U9914 ( .A(p_input[294]), .B(p_input[518]), .Z(n9866) );
  XNOR U9915 ( .A(n9891), .B(n9892), .Z(n9669) );
  AND U9916 ( .A(n306), .B(n9893), .Z(n9892) );
  XNOR U9917 ( .A(n9894), .B(n9895), .Z(n306) );
  NOR U9918 ( .A(n9896), .B(n9897), .Z(n9895) );
  XNOR U9919 ( .A(n9898), .B(n9899), .Z(n9897) );
  AND U9920 ( .A(n9898), .B(n9679), .Z(n9896) );
  IV U9921 ( .A(n9894), .Z(n9898) );
  XOR U9922 ( .A(n9900), .B(n9901), .Z(n9894) );
  AND U9923 ( .A(n9902), .B(n9903), .Z(n9901) );
  XOR U9924 ( .A(n9696), .B(n9900), .Z(n9903) );
  XOR U9925 ( .A(n9900), .B(n9697), .Z(n9902) );
  XOR U9926 ( .A(n9904), .B(n9905), .Z(n9900) );
  AND U9927 ( .A(n9906), .B(n9907), .Z(n9905) );
  XOR U9928 ( .A(n9724), .B(n9904), .Z(n9907) );
  XOR U9929 ( .A(n9904), .B(n9725), .Z(n9906) );
  XOR U9930 ( .A(n9908), .B(n9909), .Z(n9904) );
  AND U9931 ( .A(n9910), .B(n9911), .Z(n9909) );
  XOR U9932 ( .A(n9773), .B(n9908), .Z(n9911) );
  XOR U9933 ( .A(n9908), .B(n9774), .Z(n9910) );
  XOR U9934 ( .A(n9912), .B(n9913), .Z(n9908) );
  AND U9935 ( .A(n9914), .B(n9915), .Z(n9913) );
  XOR U9936 ( .A(n9912), .B(n9870), .Z(n9915) );
  XNOR U9937 ( .A(n9916), .B(n9917), .Z(n9619) );
  AND U9938 ( .A(n310), .B(n9918), .Z(n9917) );
  XNOR U9939 ( .A(n9919), .B(n9920), .Z(n310) );
  AND U9940 ( .A(n9921), .B(n9922), .Z(n9920) );
  XNOR U9941 ( .A(n9919), .B(n9580), .Z(n9922) );
  XOR U9942 ( .A(n9919), .B(n9577), .Z(n9921) );
  XOR U9943 ( .A(n9923), .B(n9924), .Z(n9919) );
  AND U9944 ( .A(n9925), .B(n9926), .Z(n9924) );
  XNOR U9945 ( .A(n9639), .B(n9923), .Z(n9926) );
  XOR U9946 ( .A(n9923), .B(n9589), .Z(n9925) );
  XOR U9947 ( .A(n9927), .B(n9928), .Z(n9923) );
  AND U9948 ( .A(n9929), .B(n9930), .Z(n9928) );
  XNOR U9949 ( .A(n9649), .B(n9927), .Z(n9930) );
  XOR U9950 ( .A(n9927), .B(n9598), .Z(n9929) );
  XOR U9951 ( .A(n9931), .B(n9932), .Z(n9927) );
  AND U9952 ( .A(n9933), .B(n9934), .Z(n9932) );
  XOR U9953 ( .A(n9931), .B(n9606), .Z(n9933) );
  XOR U9954 ( .A(n9935), .B(n9936), .Z(n9568) );
  AND U9955 ( .A(n314), .B(n9918), .Z(n9936) );
  XNOR U9956 ( .A(n9916), .B(n9935), .Z(n9918) );
  XNOR U9957 ( .A(n9937), .B(n9938), .Z(n314) );
  AND U9958 ( .A(n9939), .B(n9940), .Z(n9938) );
  XNOR U9959 ( .A(n9580), .B(n9937), .Z(n9940) );
  XNOR U9960 ( .A(n9899), .B(n9941), .Z(n9580) );
  AND U9961 ( .A(n9681), .B(n317), .Z(n9941) );
  NOR U9962 ( .A(n9942), .B(n9943), .Z(n9681) );
  XOR U9963 ( .A(n9937), .B(n9577), .Z(n9939) );
  IV U9964 ( .A(n9581), .Z(n9577) );
  AND U9965 ( .A(n9944), .B(n9945), .Z(n9581) );
  XOR U9966 ( .A(n9946), .B(n9947), .Z(n9937) );
  AND U9967 ( .A(n9948), .B(n9949), .Z(n9947) );
  XNOR U9968 ( .A(n9946), .B(n9639), .Z(n9949) );
  XOR U9969 ( .A(n9697), .B(n9950), .Z(n9639) );
  AND U9970 ( .A(n317), .B(n9951), .Z(n9950) );
  XOR U9971 ( .A(n9693), .B(n9697), .Z(n9951) );
  XNOR U9972 ( .A(n9952), .B(n9946), .Z(n9948) );
  IV U9973 ( .A(n9589), .Z(n9952) );
  XOR U9974 ( .A(n9953), .B(n9954), .Z(n9589) );
  AND U9975 ( .A(n333), .B(n9955), .Z(n9954) );
  XOR U9976 ( .A(n9956), .B(n9957), .Z(n9946) );
  AND U9977 ( .A(n9958), .B(n9959), .Z(n9957) );
  XNOR U9978 ( .A(n9956), .B(n9649), .Z(n9959) );
  XOR U9979 ( .A(n9725), .B(n9960), .Z(n9649) );
  AND U9980 ( .A(n317), .B(n9961), .Z(n9960) );
  XOR U9981 ( .A(n9721), .B(n9725), .Z(n9961) );
  XOR U9982 ( .A(n9598), .B(n9956), .Z(n9958) );
  XOR U9983 ( .A(n9962), .B(n9963), .Z(n9598) );
  AND U9984 ( .A(n333), .B(n9964), .Z(n9963) );
  XOR U9985 ( .A(n9931), .B(n9965), .Z(n9956) );
  AND U9986 ( .A(n9966), .B(n9934), .Z(n9965) );
  XNOR U9987 ( .A(n9659), .B(n9931), .Z(n9934) );
  XOR U9988 ( .A(n9774), .B(n9967), .Z(n9659) );
  AND U9989 ( .A(n317), .B(n9968), .Z(n9967) );
  XOR U9990 ( .A(n9770), .B(n9774), .Z(n9968) );
  XNOR U9991 ( .A(n9969), .B(n9931), .Z(n9966) );
  IV U9992 ( .A(n9606), .Z(n9969) );
  XOR U9993 ( .A(n9970), .B(n9971), .Z(n9606) );
  AND U9994 ( .A(n333), .B(n9972), .Z(n9971) );
  XOR U9995 ( .A(n9973), .B(n9974), .Z(n9931) );
  AND U9996 ( .A(n9975), .B(n9976), .Z(n9974) );
  XNOR U9997 ( .A(n9973), .B(n9667), .Z(n9976) );
  XOR U9998 ( .A(n9871), .B(n9977), .Z(n9667) );
  AND U9999 ( .A(n317), .B(n9978), .Z(n9977) );
  XOR U10000 ( .A(n9867), .B(n9871), .Z(n9978) );
  XNOR U10001 ( .A(n9979), .B(n9973), .Z(n9975) );
  IV U10002 ( .A(n9616), .Z(n9979) );
  XOR U10003 ( .A(n9980), .B(n9981), .Z(n9616) );
  AND U10004 ( .A(n333), .B(n9982), .Z(n9981) );
  AND U10005 ( .A(n9935), .B(n9916), .Z(n9973) );
  XNOR U10006 ( .A(n9983), .B(n9984), .Z(n9916) );
  AND U10007 ( .A(n317), .B(n9893), .Z(n9984) );
  XNOR U10008 ( .A(n9891), .B(n9983), .Z(n9893) );
  XNOR U10009 ( .A(n9985), .B(n9986), .Z(n317) );
  NOR U10010 ( .A(n9987), .B(n9988), .Z(n9986) );
  XNOR U10011 ( .A(n9989), .B(n9899), .Z(n9988) );
  IV U10012 ( .A(n9943), .Z(n9899) );
  NOR U10013 ( .A(n9944), .B(n9945), .Z(n9943) );
  AND U10014 ( .A(n9989), .B(n9679), .Z(n9987) );
  IV U10015 ( .A(n9942), .Z(n9679) );
  AND U10016 ( .A(n9990), .B(n9991), .Z(n9942) );
  IV U10017 ( .A(n9992), .Z(n9990) );
  IV U10018 ( .A(n9985), .Z(n9989) );
  XOR U10019 ( .A(n9993), .B(n9994), .Z(n9985) );
  AND U10020 ( .A(n9995), .B(n9996), .Z(n9994) );
  XNOR U10021 ( .A(n9993), .B(n9693), .Z(n9996) );
  IV U10022 ( .A(n9696), .Z(n9693) );
  XOR U10023 ( .A(n9997), .B(n9998), .Z(n9696) );
  AND U10024 ( .A(n321), .B(n9999), .Z(n9998) );
  XOR U10025 ( .A(n10000), .B(n9997), .Z(n9999) );
  XOR U10026 ( .A(n9697), .B(n9993), .Z(n9995) );
  XOR U10027 ( .A(n10001), .B(n10002), .Z(n9697) );
  AND U10028 ( .A(n329), .B(n9955), .Z(n10002) );
  XOR U10029 ( .A(n10001), .B(n9953), .Z(n9955) );
  XOR U10030 ( .A(n10003), .B(n10004), .Z(n9993) );
  AND U10031 ( .A(n10005), .B(n10006), .Z(n10004) );
  XNOR U10032 ( .A(n10003), .B(n9721), .Z(n10006) );
  IV U10033 ( .A(n9724), .Z(n9721) );
  XOR U10034 ( .A(n10007), .B(n10008), .Z(n9724) );
  AND U10035 ( .A(n321), .B(n10009), .Z(n10008) );
  XNOR U10036 ( .A(n10010), .B(n10007), .Z(n10009) );
  XOR U10037 ( .A(n9725), .B(n10003), .Z(n10005) );
  XOR U10038 ( .A(n10011), .B(n10012), .Z(n9725) );
  AND U10039 ( .A(n329), .B(n9964), .Z(n10012) );
  XOR U10040 ( .A(n10011), .B(n9962), .Z(n9964) );
  XOR U10041 ( .A(n10013), .B(n10014), .Z(n10003) );
  AND U10042 ( .A(n10015), .B(n10016), .Z(n10014) );
  XNOR U10043 ( .A(n10013), .B(n9770), .Z(n10016) );
  IV U10044 ( .A(n9773), .Z(n9770) );
  XOR U10045 ( .A(n10017), .B(n10018), .Z(n9773) );
  AND U10046 ( .A(n321), .B(n10019), .Z(n10018) );
  XOR U10047 ( .A(n10020), .B(n10017), .Z(n10019) );
  XOR U10048 ( .A(n9774), .B(n10013), .Z(n10015) );
  XOR U10049 ( .A(n10021), .B(n10022), .Z(n9774) );
  AND U10050 ( .A(n329), .B(n9972), .Z(n10022) );
  XOR U10051 ( .A(n10021), .B(n9970), .Z(n9972) );
  XOR U10052 ( .A(n9912), .B(n10023), .Z(n10013) );
  AND U10053 ( .A(n9914), .B(n10024), .Z(n10023) );
  XNOR U10054 ( .A(n9912), .B(n9867), .Z(n10024) );
  IV U10055 ( .A(n9870), .Z(n9867) );
  XOR U10056 ( .A(n10025), .B(n10026), .Z(n9870) );
  AND U10057 ( .A(n321), .B(n10027), .Z(n10026) );
  XNOR U10058 ( .A(n10028), .B(n10025), .Z(n10027) );
  XOR U10059 ( .A(n9871), .B(n9912), .Z(n9914) );
  XOR U10060 ( .A(n10029), .B(n10030), .Z(n9871) );
  AND U10061 ( .A(n329), .B(n9982), .Z(n10030) );
  XOR U10062 ( .A(n10029), .B(n9980), .Z(n9982) );
  AND U10063 ( .A(n9983), .B(n9891), .Z(n9912) );
  XNOR U10064 ( .A(n10031), .B(n10032), .Z(n9891) );
  AND U10065 ( .A(n321), .B(n10033), .Z(n10032) );
  XNOR U10066 ( .A(n10034), .B(n10031), .Z(n10033) );
  XNOR U10067 ( .A(n10035), .B(n10036), .Z(n321) );
  NOR U10068 ( .A(n10037), .B(n10038), .Z(n10036) );
  XNOR U10069 ( .A(n10035), .B(n9992), .Z(n10038) );
  NOR U10070 ( .A(n10039), .B(n10040), .Z(n9992) );
  NOR U10071 ( .A(n10035), .B(n9991), .Z(n10037) );
  AND U10072 ( .A(n10041), .B(n10042), .Z(n9991) );
  XOR U10073 ( .A(n10043), .B(n10044), .Z(n10035) );
  AND U10074 ( .A(n10045), .B(n10046), .Z(n10044) );
  XNOR U10075 ( .A(n10043), .B(n10041), .Z(n10046) );
  IV U10076 ( .A(n10000), .Z(n10041) );
  XOR U10077 ( .A(n10047), .B(n10048), .Z(n10000) );
  XOR U10078 ( .A(n10049), .B(n10042), .Z(n10048) );
  AND U10079 ( .A(n10010), .B(n10050), .Z(n10042) );
  AND U10080 ( .A(n10051), .B(n10052), .Z(n10049) );
  XOR U10081 ( .A(n10053), .B(n10047), .Z(n10051) );
  XNOR U10082 ( .A(n9997), .B(n10043), .Z(n10045) );
  XNOR U10083 ( .A(n10054), .B(n10055), .Z(n9997) );
  AND U10084 ( .A(n325), .B(n10056), .Z(n10055) );
  XNOR U10085 ( .A(n10057), .B(n10058), .Z(n10056) );
  XOR U10086 ( .A(n10059), .B(n10060), .Z(n10043) );
  AND U10087 ( .A(n10061), .B(n10062), .Z(n10060) );
  XNOR U10088 ( .A(n10059), .B(n10010), .Z(n10062) );
  XOR U10089 ( .A(n10063), .B(n10052), .Z(n10010) );
  XNOR U10090 ( .A(n10064), .B(n10047), .Z(n10052) );
  XOR U10091 ( .A(n10065), .B(n10066), .Z(n10047) );
  AND U10092 ( .A(n10067), .B(n10068), .Z(n10066) );
  XOR U10093 ( .A(n10069), .B(n10065), .Z(n10067) );
  XNOR U10094 ( .A(n10070), .B(n10071), .Z(n10064) );
  AND U10095 ( .A(n10072), .B(n10073), .Z(n10071) );
  XOR U10096 ( .A(n10070), .B(n10074), .Z(n10072) );
  XNOR U10097 ( .A(n10053), .B(n10050), .Z(n10063) );
  AND U10098 ( .A(n10075), .B(n10076), .Z(n10050) );
  XOR U10099 ( .A(n10077), .B(n10078), .Z(n10053) );
  AND U10100 ( .A(n10079), .B(n10080), .Z(n10078) );
  XOR U10101 ( .A(n10077), .B(n10081), .Z(n10079) );
  XNOR U10102 ( .A(n10007), .B(n10059), .Z(n10061) );
  XNOR U10103 ( .A(n10082), .B(n10083), .Z(n10007) );
  AND U10104 ( .A(n325), .B(n10084), .Z(n10083) );
  XNOR U10105 ( .A(n10085), .B(n10086), .Z(n10084) );
  XOR U10106 ( .A(n10087), .B(n10088), .Z(n10059) );
  AND U10107 ( .A(n10089), .B(n10090), .Z(n10088) );
  XNOR U10108 ( .A(n10087), .B(n10075), .Z(n10090) );
  IV U10109 ( .A(n10020), .Z(n10075) );
  XNOR U10110 ( .A(n10091), .B(n10068), .Z(n10020) );
  XNOR U10111 ( .A(n10092), .B(n10074), .Z(n10068) );
  XOR U10112 ( .A(n10093), .B(n10094), .Z(n10074) );
  AND U10113 ( .A(n10095), .B(n10096), .Z(n10094) );
  XOR U10114 ( .A(n10093), .B(n10097), .Z(n10095) );
  XNOR U10115 ( .A(n10073), .B(n10065), .Z(n10092) );
  XOR U10116 ( .A(n10098), .B(n10099), .Z(n10065) );
  AND U10117 ( .A(n10100), .B(n10101), .Z(n10099) );
  XNOR U10118 ( .A(n10102), .B(n10098), .Z(n10100) );
  XNOR U10119 ( .A(n10103), .B(n10070), .Z(n10073) );
  XOR U10120 ( .A(n10104), .B(n10105), .Z(n10070) );
  AND U10121 ( .A(n10106), .B(n10107), .Z(n10105) );
  XOR U10122 ( .A(n10104), .B(n10108), .Z(n10106) );
  XNOR U10123 ( .A(n10109), .B(n10110), .Z(n10103) );
  AND U10124 ( .A(n10111), .B(n10112), .Z(n10110) );
  XNOR U10125 ( .A(n10109), .B(n10113), .Z(n10111) );
  XNOR U10126 ( .A(n10069), .B(n10076), .Z(n10091) );
  AND U10127 ( .A(n10028), .B(n10114), .Z(n10076) );
  XOR U10128 ( .A(n10081), .B(n10080), .Z(n10069) );
  XNOR U10129 ( .A(n10115), .B(n10077), .Z(n10080) );
  XOR U10130 ( .A(n10116), .B(n10117), .Z(n10077) );
  AND U10131 ( .A(n10118), .B(n10119), .Z(n10117) );
  XOR U10132 ( .A(n10116), .B(n10120), .Z(n10118) );
  XNOR U10133 ( .A(n10121), .B(n10122), .Z(n10115) );
  AND U10134 ( .A(n10123), .B(n10124), .Z(n10122) );
  XOR U10135 ( .A(n10121), .B(n10125), .Z(n10123) );
  XOR U10136 ( .A(n10126), .B(n10127), .Z(n10081) );
  AND U10137 ( .A(n10128), .B(n10129), .Z(n10127) );
  XOR U10138 ( .A(n10126), .B(n10130), .Z(n10128) );
  XNOR U10139 ( .A(n10017), .B(n10087), .Z(n10089) );
  XNOR U10140 ( .A(n10131), .B(n10132), .Z(n10017) );
  AND U10141 ( .A(n325), .B(n10133), .Z(n10132) );
  XNOR U10142 ( .A(n10134), .B(n10135), .Z(n10133) );
  XOR U10143 ( .A(n10136), .B(n10137), .Z(n10087) );
  AND U10144 ( .A(n10138), .B(n10139), .Z(n10137) );
  XNOR U10145 ( .A(n10136), .B(n10028), .Z(n10139) );
  XOR U10146 ( .A(n10140), .B(n10101), .Z(n10028) );
  XNOR U10147 ( .A(n10141), .B(n10108), .Z(n10101) );
  XOR U10148 ( .A(n10097), .B(n10096), .Z(n10108) );
  XNOR U10149 ( .A(n10142), .B(n10093), .Z(n10096) );
  XOR U10150 ( .A(n10143), .B(n10144), .Z(n10093) );
  AND U10151 ( .A(n10145), .B(n10146), .Z(n10144) );
  XNOR U10152 ( .A(n10147), .B(n10148), .Z(n10145) );
  IV U10153 ( .A(n10143), .Z(n10147) );
  XNOR U10154 ( .A(n10149), .B(n10150), .Z(n10142) );
  NOR U10155 ( .A(n10151), .B(n10152), .Z(n10150) );
  XNOR U10156 ( .A(n10149), .B(n10153), .Z(n10151) );
  XOR U10157 ( .A(n10154), .B(n10155), .Z(n10097) );
  NOR U10158 ( .A(n10156), .B(n10157), .Z(n10155) );
  XNOR U10159 ( .A(n10154), .B(n10158), .Z(n10156) );
  XNOR U10160 ( .A(n10107), .B(n10098), .Z(n10141) );
  XOR U10161 ( .A(n10159), .B(n10160), .Z(n10098) );
  AND U10162 ( .A(n10161), .B(n10162), .Z(n10160) );
  XOR U10163 ( .A(n10159), .B(n10163), .Z(n10161) );
  XOR U10164 ( .A(n10164), .B(n10113), .Z(n10107) );
  XOR U10165 ( .A(n10165), .B(n10166), .Z(n10113) );
  NOR U10166 ( .A(n10167), .B(n10168), .Z(n10166) );
  XOR U10167 ( .A(n10165), .B(n10169), .Z(n10167) );
  XNOR U10168 ( .A(n10112), .B(n10104), .Z(n10164) );
  XOR U10169 ( .A(n10170), .B(n10171), .Z(n10104) );
  AND U10170 ( .A(n10172), .B(n10173), .Z(n10171) );
  XOR U10171 ( .A(n10170), .B(n10174), .Z(n10172) );
  XNOR U10172 ( .A(n10175), .B(n10109), .Z(n10112) );
  XOR U10173 ( .A(n10176), .B(n10177), .Z(n10109) );
  AND U10174 ( .A(n10178), .B(n10179), .Z(n10177) );
  XNOR U10175 ( .A(n10180), .B(n10181), .Z(n10178) );
  IV U10176 ( .A(n10176), .Z(n10180) );
  XNOR U10177 ( .A(n10182), .B(n10183), .Z(n10175) );
  NOR U10178 ( .A(n10184), .B(n10185), .Z(n10183) );
  XNOR U10179 ( .A(n10182), .B(n10186), .Z(n10184) );
  XOR U10180 ( .A(n10102), .B(n10114), .Z(n10140) );
  NOR U10181 ( .A(n10034), .B(n10187), .Z(n10114) );
  XNOR U10182 ( .A(n10120), .B(n10119), .Z(n10102) );
  XNOR U10183 ( .A(n10188), .B(n10125), .Z(n10119) );
  XNOR U10184 ( .A(n10189), .B(n10190), .Z(n10125) );
  NOR U10185 ( .A(n10191), .B(n10192), .Z(n10190) );
  XOR U10186 ( .A(n10189), .B(n10193), .Z(n10191) );
  XNOR U10187 ( .A(n10124), .B(n10116), .Z(n10188) );
  XOR U10188 ( .A(n10194), .B(n10195), .Z(n10116) );
  AND U10189 ( .A(n10196), .B(n10197), .Z(n10195) );
  XOR U10190 ( .A(n10194), .B(n10198), .Z(n10196) );
  XNOR U10191 ( .A(n10199), .B(n10121), .Z(n10124) );
  XOR U10192 ( .A(n10200), .B(n10201), .Z(n10121) );
  AND U10193 ( .A(n10202), .B(n10203), .Z(n10201) );
  XNOR U10194 ( .A(n10204), .B(n10205), .Z(n10202) );
  IV U10195 ( .A(n10200), .Z(n10204) );
  XNOR U10196 ( .A(n10206), .B(n10207), .Z(n10199) );
  NOR U10197 ( .A(n10208), .B(n10209), .Z(n10207) );
  XNOR U10198 ( .A(n10206), .B(n10210), .Z(n10208) );
  XOR U10199 ( .A(n10130), .B(n10129), .Z(n10120) );
  XNOR U10200 ( .A(n10211), .B(n10126), .Z(n10129) );
  XOR U10201 ( .A(n10212), .B(n10213), .Z(n10126) );
  AND U10202 ( .A(n10214), .B(n10215), .Z(n10213) );
  XNOR U10203 ( .A(n10216), .B(n10217), .Z(n10214) );
  IV U10204 ( .A(n10212), .Z(n10216) );
  XNOR U10205 ( .A(n10218), .B(n10219), .Z(n10211) );
  NOR U10206 ( .A(n10220), .B(n10221), .Z(n10219) );
  XNOR U10207 ( .A(n10218), .B(n10222), .Z(n10220) );
  XOR U10208 ( .A(n10223), .B(n10224), .Z(n10130) );
  NOR U10209 ( .A(n10225), .B(n10226), .Z(n10224) );
  XNOR U10210 ( .A(n10223), .B(n10227), .Z(n10225) );
  XNOR U10211 ( .A(n10025), .B(n10136), .Z(n10138) );
  XNOR U10212 ( .A(n10228), .B(n10229), .Z(n10025) );
  AND U10213 ( .A(n325), .B(n10230), .Z(n10229) );
  XNOR U10214 ( .A(n10231), .B(n10232), .Z(n10230) );
  AND U10215 ( .A(n10031), .B(n10034), .Z(n10136) );
  XOR U10216 ( .A(n10233), .B(n10187), .Z(n10034) );
  XNOR U10217 ( .A(p_input[320]), .B(p_input[512]), .Z(n10187) );
  XNOR U10218 ( .A(n10163), .B(n10162), .Z(n10233) );
  XNOR U10219 ( .A(n10234), .B(n10174), .Z(n10162) );
  XOR U10220 ( .A(n10148), .B(n10146), .Z(n10174) );
  XNOR U10221 ( .A(n10235), .B(n10153), .Z(n10146) );
  XOR U10222 ( .A(p_input[344]), .B(p_input[536]), .Z(n10153) );
  XOR U10223 ( .A(n10143), .B(n10152), .Z(n10235) );
  XOR U10224 ( .A(n10236), .B(n10149), .Z(n10152) );
  XOR U10225 ( .A(p_input[342]), .B(p_input[534]), .Z(n10149) );
  XOR U10226 ( .A(p_input[343]), .B(n6576), .Z(n10236) );
  XOR U10227 ( .A(p_input[338]), .B(p_input[530]), .Z(n10143) );
  XNOR U10228 ( .A(n10158), .B(n10157), .Z(n10148) );
  XOR U10229 ( .A(n10237), .B(n10154), .Z(n10157) );
  XOR U10230 ( .A(p_input[339]), .B(p_input[531]), .Z(n10154) );
  XOR U10231 ( .A(p_input[340]), .B(n6578), .Z(n10237) );
  XOR U10232 ( .A(p_input[341]), .B(p_input[533]), .Z(n10158) );
  XOR U10233 ( .A(n10173), .B(n10238), .Z(n10234) );
  IV U10234 ( .A(n10159), .Z(n10238) );
  XOR U10235 ( .A(p_input[321]), .B(p_input[513]), .Z(n10159) );
  XNOR U10236 ( .A(n10239), .B(n10181), .Z(n10173) );
  XNOR U10237 ( .A(n10169), .B(n10168), .Z(n10181) );
  XNOR U10238 ( .A(n10240), .B(n10165), .Z(n10168) );
  XNOR U10239 ( .A(p_input[346]), .B(p_input[538]), .Z(n10165) );
  XOR U10240 ( .A(p_input[347]), .B(n6582), .Z(n10240) );
  XOR U10241 ( .A(p_input[348]), .B(p_input[540]), .Z(n10169) );
  XOR U10242 ( .A(n10179), .B(n10241), .Z(n10239) );
  IV U10243 ( .A(n10170), .Z(n10241) );
  XOR U10244 ( .A(p_input[337]), .B(p_input[529]), .Z(n10170) );
  XNOR U10245 ( .A(n10242), .B(n10186), .Z(n10179) );
  XNOR U10246 ( .A(p_input[351]), .B(n6585), .Z(n10186) );
  XOR U10247 ( .A(n10176), .B(n10185), .Z(n10242) );
  XOR U10248 ( .A(n10243), .B(n10182), .Z(n10185) );
  XOR U10249 ( .A(p_input[349]), .B(p_input[541]), .Z(n10182) );
  XOR U10250 ( .A(p_input[350]), .B(n6587), .Z(n10243) );
  XOR U10251 ( .A(p_input[345]), .B(p_input[537]), .Z(n10176) );
  XOR U10252 ( .A(n10198), .B(n10197), .Z(n10163) );
  XNOR U10253 ( .A(n10244), .B(n10205), .Z(n10197) );
  XNOR U10254 ( .A(n10193), .B(n10192), .Z(n10205) );
  XNOR U10255 ( .A(n10245), .B(n10189), .Z(n10192) );
  XNOR U10256 ( .A(p_input[331]), .B(p_input[523]), .Z(n10189) );
  XOR U10257 ( .A(p_input[332]), .B(n6590), .Z(n10245) );
  XOR U10258 ( .A(p_input[333]), .B(p_input[525]), .Z(n10193) );
  XOR U10259 ( .A(n10203), .B(n10246), .Z(n10244) );
  IV U10260 ( .A(n10194), .Z(n10246) );
  XOR U10261 ( .A(p_input[322]), .B(p_input[514]), .Z(n10194) );
  XNOR U10262 ( .A(n10247), .B(n10210), .Z(n10203) );
  XNOR U10263 ( .A(p_input[336]), .B(n6593), .Z(n10210) );
  XOR U10264 ( .A(n10200), .B(n10209), .Z(n10247) );
  XOR U10265 ( .A(n10248), .B(n10206), .Z(n10209) );
  XOR U10266 ( .A(p_input[334]), .B(p_input[526]), .Z(n10206) );
  XOR U10267 ( .A(p_input[335]), .B(n6595), .Z(n10248) );
  XOR U10268 ( .A(p_input[330]), .B(p_input[522]), .Z(n10200) );
  XOR U10269 ( .A(n10217), .B(n10215), .Z(n10198) );
  XNOR U10270 ( .A(n10249), .B(n10222), .Z(n10215) );
  XOR U10271 ( .A(p_input[329]), .B(p_input[521]), .Z(n10222) );
  XOR U10272 ( .A(n10212), .B(n10221), .Z(n10249) );
  XOR U10273 ( .A(n10250), .B(n10218), .Z(n10221) );
  XOR U10274 ( .A(p_input[327]), .B(p_input[519]), .Z(n10218) );
  XOR U10275 ( .A(p_input[328]), .B(n6963), .Z(n10250) );
  XOR U10276 ( .A(p_input[323]), .B(p_input[515]), .Z(n10212) );
  XNOR U10277 ( .A(n10227), .B(n10226), .Z(n10217) );
  XOR U10278 ( .A(n10251), .B(n10223), .Z(n10226) );
  XOR U10279 ( .A(p_input[324]), .B(p_input[516]), .Z(n10223) );
  XOR U10280 ( .A(p_input[325]), .B(n6965), .Z(n10251) );
  XOR U10281 ( .A(p_input[326]), .B(p_input[518]), .Z(n10227) );
  XNOR U10282 ( .A(n10252), .B(n10253), .Z(n10031) );
  AND U10283 ( .A(n325), .B(n10254), .Z(n10253) );
  XNOR U10284 ( .A(n10255), .B(n10256), .Z(n325) );
  NOR U10285 ( .A(n10257), .B(n10258), .Z(n10256) );
  XNOR U10286 ( .A(n10255), .B(n10259), .Z(n10258) );
  NOR U10287 ( .A(n10255), .B(n10040), .Z(n10257) );
  XOR U10288 ( .A(n10260), .B(n10261), .Z(n10255) );
  AND U10289 ( .A(n10262), .B(n10263), .Z(n10261) );
  XOR U10290 ( .A(n10057), .B(n10260), .Z(n10263) );
  XOR U10291 ( .A(n10260), .B(n10058), .Z(n10262) );
  XOR U10292 ( .A(n10264), .B(n10265), .Z(n10260) );
  AND U10293 ( .A(n10266), .B(n10267), .Z(n10265) );
  XOR U10294 ( .A(n10085), .B(n10264), .Z(n10267) );
  XOR U10295 ( .A(n10264), .B(n10086), .Z(n10266) );
  XOR U10296 ( .A(n10268), .B(n10269), .Z(n10264) );
  AND U10297 ( .A(n10270), .B(n10271), .Z(n10269) );
  XOR U10298 ( .A(n10134), .B(n10268), .Z(n10271) );
  XOR U10299 ( .A(n10268), .B(n10135), .Z(n10270) );
  XOR U10300 ( .A(n10272), .B(n10273), .Z(n10268) );
  AND U10301 ( .A(n10274), .B(n10275), .Z(n10273) );
  XOR U10302 ( .A(n10272), .B(n10231), .Z(n10275) );
  XNOR U10303 ( .A(n10276), .B(n10277), .Z(n9983) );
  AND U10304 ( .A(n329), .B(n10278), .Z(n10277) );
  XNOR U10305 ( .A(n10279), .B(n10280), .Z(n329) );
  NOR U10306 ( .A(n10281), .B(n10282), .Z(n10280) );
  XOR U10307 ( .A(n9945), .B(n10279), .Z(n10282) );
  NOR U10308 ( .A(n10279), .B(n9944), .Z(n10281) );
  XOR U10309 ( .A(n10283), .B(n10284), .Z(n10279) );
  AND U10310 ( .A(n10285), .B(n10286), .Z(n10284) );
  XNOR U10311 ( .A(n10001), .B(n10283), .Z(n10286) );
  XOR U10312 ( .A(n10283), .B(n9953), .Z(n10285) );
  XOR U10313 ( .A(n10287), .B(n10288), .Z(n10283) );
  AND U10314 ( .A(n10289), .B(n10290), .Z(n10288) );
  XNOR U10315 ( .A(n10011), .B(n10287), .Z(n10290) );
  XOR U10316 ( .A(n10287), .B(n9962), .Z(n10289) );
  XOR U10317 ( .A(n10291), .B(n10292), .Z(n10287) );
  AND U10318 ( .A(n10293), .B(n10294), .Z(n10292) );
  XOR U10319 ( .A(n10291), .B(n9970), .Z(n10293) );
  XOR U10320 ( .A(n10295), .B(n10296), .Z(n9935) );
  AND U10321 ( .A(n333), .B(n10278), .Z(n10296) );
  XNOR U10322 ( .A(n10276), .B(n10295), .Z(n10278) );
  XNOR U10323 ( .A(n10297), .B(n10298), .Z(n333) );
  NOR U10324 ( .A(n10299), .B(n10300), .Z(n10298) );
  XNOR U10325 ( .A(n9945), .B(n10301), .Z(n10300) );
  IV U10326 ( .A(n10297), .Z(n10301) );
  AND U10327 ( .A(n10302), .B(n10303), .Z(n9945) );
  NOR U10328 ( .A(n10297), .B(n9944), .Z(n10299) );
  AND U10329 ( .A(n10040), .B(n10039), .Z(n9944) );
  IV U10330 ( .A(n10259), .Z(n10039) );
  XOR U10331 ( .A(n10304), .B(n10305), .Z(n10297) );
  AND U10332 ( .A(n10306), .B(n10307), .Z(n10305) );
  XNOR U10333 ( .A(n10304), .B(n10001), .Z(n10307) );
  XOR U10334 ( .A(n10058), .B(n10308), .Z(n10001) );
  AND U10335 ( .A(n336), .B(n10309), .Z(n10308) );
  XOR U10336 ( .A(n10054), .B(n10058), .Z(n10309) );
  XNOR U10337 ( .A(n10310), .B(n10304), .Z(n10306) );
  IV U10338 ( .A(n9953), .Z(n10310) );
  XOR U10339 ( .A(n10311), .B(n10312), .Z(n9953) );
  AND U10340 ( .A(n352), .B(n10313), .Z(n10312) );
  XOR U10341 ( .A(n10314), .B(n10315), .Z(n10304) );
  AND U10342 ( .A(n10316), .B(n10317), .Z(n10315) );
  XNOR U10343 ( .A(n10314), .B(n10011), .Z(n10317) );
  XOR U10344 ( .A(n10086), .B(n10318), .Z(n10011) );
  AND U10345 ( .A(n336), .B(n10319), .Z(n10318) );
  XOR U10346 ( .A(n10082), .B(n10086), .Z(n10319) );
  XOR U10347 ( .A(n9962), .B(n10314), .Z(n10316) );
  XOR U10348 ( .A(n10320), .B(n10321), .Z(n9962) );
  AND U10349 ( .A(n352), .B(n10322), .Z(n10321) );
  XOR U10350 ( .A(n10291), .B(n10323), .Z(n10314) );
  AND U10351 ( .A(n10324), .B(n10294), .Z(n10323) );
  XNOR U10352 ( .A(n10021), .B(n10291), .Z(n10294) );
  XOR U10353 ( .A(n10135), .B(n10325), .Z(n10021) );
  AND U10354 ( .A(n336), .B(n10326), .Z(n10325) );
  XOR U10355 ( .A(n10131), .B(n10135), .Z(n10326) );
  XNOR U10356 ( .A(n10327), .B(n10291), .Z(n10324) );
  IV U10357 ( .A(n9970), .Z(n10327) );
  XOR U10358 ( .A(n10328), .B(n10329), .Z(n9970) );
  AND U10359 ( .A(n352), .B(n10330), .Z(n10329) );
  XOR U10360 ( .A(n10331), .B(n10332), .Z(n10291) );
  AND U10361 ( .A(n10333), .B(n10334), .Z(n10332) );
  XNOR U10362 ( .A(n10331), .B(n10029), .Z(n10334) );
  XOR U10363 ( .A(n10232), .B(n10335), .Z(n10029) );
  AND U10364 ( .A(n336), .B(n10336), .Z(n10335) );
  XOR U10365 ( .A(n10228), .B(n10232), .Z(n10336) );
  XNOR U10366 ( .A(n10337), .B(n10331), .Z(n10333) );
  IV U10367 ( .A(n9980), .Z(n10337) );
  XOR U10368 ( .A(n10338), .B(n10339), .Z(n9980) );
  AND U10369 ( .A(n352), .B(n10340), .Z(n10339) );
  AND U10370 ( .A(n10295), .B(n10276), .Z(n10331) );
  XNOR U10371 ( .A(n10341), .B(n10342), .Z(n10276) );
  AND U10372 ( .A(n336), .B(n10254), .Z(n10342) );
  XNOR U10373 ( .A(n10252), .B(n10341), .Z(n10254) );
  XNOR U10374 ( .A(n10343), .B(n10344), .Z(n336) );
  NOR U10375 ( .A(n10345), .B(n10346), .Z(n10344) );
  XNOR U10376 ( .A(n10343), .B(n10259), .Z(n10346) );
  NOR U10377 ( .A(n10302), .B(n10303), .Z(n10259) );
  NOR U10378 ( .A(n10343), .B(n10040), .Z(n10345) );
  AND U10379 ( .A(n10347), .B(n10348), .Z(n10040) );
  IV U10380 ( .A(n10349), .Z(n10347) );
  XOR U10381 ( .A(n10350), .B(n10351), .Z(n10343) );
  AND U10382 ( .A(n10352), .B(n10353), .Z(n10351) );
  XNOR U10383 ( .A(n10350), .B(n10054), .Z(n10353) );
  IV U10384 ( .A(n10057), .Z(n10054) );
  XOR U10385 ( .A(n10354), .B(n10355), .Z(n10057) );
  AND U10386 ( .A(n340), .B(n10356), .Z(n10355) );
  XOR U10387 ( .A(n10357), .B(n10354), .Z(n10356) );
  XOR U10388 ( .A(n10058), .B(n10350), .Z(n10352) );
  XOR U10389 ( .A(n10358), .B(n10359), .Z(n10058) );
  AND U10390 ( .A(n348), .B(n10313), .Z(n10359) );
  XOR U10391 ( .A(n10358), .B(n10311), .Z(n10313) );
  XOR U10392 ( .A(n10360), .B(n10361), .Z(n10350) );
  AND U10393 ( .A(n10362), .B(n10363), .Z(n10361) );
  XNOR U10394 ( .A(n10360), .B(n10082), .Z(n10363) );
  IV U10395 ( .A(n10085), .Z(n10082) );
  XOR U10396 ( .A(n10364), .B(n10365), .Z(n10085) );
  AND U10397 ( .A(n340), .B(n10366), .Z(n10365) );
  XNOR U10398 ( .A(n10367), .B(n10364), .Z(n10366) );
  XOR U10399 ( .A(n10086), .B(n10360), .Z(n10362) );
  XOR U10400 ( .A(n10368), .B(n10369), .Z(n10086) );
  AND U10401 ( .A(n348), .B(n10322), .Z(n10369) );
  XOR U10402 ( .A(n10368), .B(n10320), .Z(n10322) );
  XOR U10403 ( .A(n10370), .B(n10371), .Z(n10360) );
  AND U10404 ( .A(n10372), .B(n10373), .Z(n10371) );
  XNOR U10405 ( .A(n10370), .B(n10131), .Z(n10373) );
  IV U10406 ( .A(n10134), .Z(n10131) );
  XOR U10407 ( .A(n10374), .B(n10375), .Z(n10134) );
  AND U10408 ( .A(n340), .B(n10376), .Z(n10375) );
  XOR U10409 ( .A(n10377), .B(n10374), .Z(n10376) );
  XOR U10410 ( .A(n10135), .B(n10370), .Z(n10372) );
  XOR U10411 ( .A(n10378), .B(n10379), .Z(n10135) );
  AND U10412 ( .A(n348), .B(n10330), .Z(n10379) );
  XOR U10413 ( .A(n10378), .B(n10328), .Z(n10330) );
  XOR U10414 ( .A(n10272), .B(n10380), .Z(n10370) );
  AND U10415 ( .A(n10274), .B(n10381), .Z(n10380) );
  XNOR U10416 ( .A(n10272), .B(n10228), .Z(n10381) );
  IV U10417 ( .A(n10231), .Z(n10228) );
  XOR U10418 ( .A(n10382), .B(n10383), .Z(n10231) );
  AND U10419 ( .A(n340), .B(n10384), .Z(n10383) );
  XNOR U10420 ( .A(n10385), .B(n10382), .Z(n10384) );
  XOR U10421 ( .A(n10232), .B(n10272), .Z(n10274) );
  XOR U10422 ( .A(n10386), .B(n10387), .Z(n10232) );
  AND U10423 ( .A(n348), .B(n10340), .Z(n10387) );
  XOR U10424 ( .A(n10386), .B(n10338), .Z(n10340) );
  AND U10425 ( .A(n10341), .B(n10252), .Z(n10272) );
  XNOR U10426 ( .A(n10388), .B(n10389), .Z(n10252) );
  AND U10427 ( .A(n340), .B(n10390), .Z(n10389) );
  XNOR U10428 ( .A(n10391), .B(n10388), .Z(n10390) );
  XNOR U10429 ( .A(n10392), .B(n10393), .Z(n340) );
  NOR U10430 ( .A(n10394), .B(n10395), .Z(n10393) );
  XNOR U10431 ( .A(n10392), .B(n10349), .Z(n10395) );
  NOR U10432 ( .A(n10396), .B(n10397), .Z(n10349) );
  NOR U10433 ( .A(n10392), .B(n10348), .Z(n10394) );
  AND U10434 ( .A(n10398), .B(n10399), .Z(n10348) );
  XOR U10435 ( .A(n10400), .B(n10401), .Z(n10392) );
  AND U10436 ( .A(n10402), .B(n10403), .Z(n10401) );
  XNOR U10437 ( .A(n10400), .B(n10398), .Z(n10403) );
  IV U10438 ( .A(n10357), .Z(n10398) );
  XOR U10439 ( .A(n10404), .B(n10405), .Z(n10357) );
  XOR U10440 ( .A(n10406), .B(n10399), .Z(n10405) );
  AND U10441 ( .A(n10367), .B(n10407), .Z(n10399) );
  AND U10442 ( .A(n10408), .B(n10409), .Z(n10406) );
  XOR U10443 ( .A(n10410), .B(n10404), .Z(n10408) );
  XNOR U10444 ( .A(n10354), .B(n10400), .Z(n10402) );
  XNOR U10445 ( .A(n10411), .B(n10412), .Z(n10354) );
  AND U10446 ( .A(n344), .B(n10413), .Z(n10412) );
  XNOR U10447 ( .A(n10414), .B(n10415), .Z(n10413) );
  XOR U10448 ( .A(n10416), .B(n10417), .Z(n10400) );
  AND U10449 ( .A(n10418), .B(n10419), .Z(n10417) );
  XNOR U10450 ( .A(n10416), .B(n10367), .Z(n10419) );
  XOR U10451 ( .A(n10420), .B(n10409), .Z(n10367) );
  XNOR U10452 ( .A(n10421), .B(n10404), .Z(n10409) );
  XOR U10453 ( .A(n10422), .B(n10423), .Z(n10404) );
  AND U10454 ( .A(n10424), .B(n10425), .Z(n10423) );
  XOR U10455 ( .A(n10426), .B(n10422), .Z(n10424) );
  XNOR U10456 ( .A(n10427), .B(n10428), .Z(n10421) );
  AND U10457 ( .A(n10429), .B(n10430), .Z(n10428) );
  XOR U10458 ( .A(n10427), .B(n10431), .Z(n10429) );
  XNOR U10459 ( .A(n10410), .B(n10407), .Z(n10420) );
  AND U10460 ( .A(n10432), .B(n10433), .Z(n10407) );
  XOR U10461 ( .A(n10434), .B(n10435), .Z(n10410) );
  AND U10462 ( .A(n10436), .B(n10437), .Z(n10435) );
  XOR U10463 ( .A(n10434), .B(n10438), .Z(n10436) );
  XNOR U10464 ( .A(n10364), .B(n10416), .Z(n10418) );
  XNOR U10465 ( .A(n10439), .B(n10440), .Z(n10364) );
  AND U10466 ( .A(n344), .B(n10441), .Z(n10440) );
  XNOR U10467 ( .A(n10442), .B(n10443), .Z(n10441) );
  XOR U10468 ( .A(n10444), .B(n10445), .Z(n10416) );
  AND U10469 ( .A(n10446), .B(n10447), .Z(n10445) );
  XNOR U10470 ( .A(n10444), .B(n10432), .Z(n10447) );
  IV U10471 ( .A(n10377), .Z(n10432) );
  XNOR U10472 ( .A(n10448), .B(n10425), .Z(n10377) );
  XNOR U10473 ( .A(n10449), .B(n10431), .Z(n10425) );
  XOR U10474 ( .A(n10450), .B(n10451), .Z(n10431) );
  AND U10475 ( .A(n10452), .B(n10453), .Z(n10451) );
  XOR U10476 ( .A(n10450), .B(n10454), .Z(n10452) );
  XNOR U10477 ( .A(n10430), .B(n10422), .Z(n10449) );
  XOR U10478 ( .A(n10455), .B(n10456), .Z(n10422) );
  AND U10479 ( .A(n10457), .B(n10458), .Z(n10456) );
  XNOR U10480 ( .A(n10459), .B(n10455), .Z(n10457) );
  XNOR U10481 ( .A(n10460), .B(n10427), .Z(n10430) );
  XOR U10482 ( .A(n10461), .B(n10462), .Z(n10427) );
  AND U10483 ( .A(n10463), .B(n10464), .Z(n10462) );
  XOR U10484 ( .A(n10461), .B(n10465), .Z(n10463) );
  XNOR U10485 ( .A(n10466), .B(n10467), .Z(n10460) );
  AND U10486 ( .A(n10468), .B(n10469), .Z(n10467) );
  XNOR U10487 ( .A(n10466), .B(n10470), .Z(n10468) );
  XNOR U10488 ( .A(n10426), .B(n10433), .Z(n10448) );
  AND U10489 ( .A(n10385), .B(n10471), .Z(n10433) );
  XOR U10490 ( .A(n10438), .B(n10437), .Z(n10426) );
  XNOR U10491 ( .A(n10472), .B(n10434), .Z(n10437) );
  XOR U10492 ( .A(n10473), .B(n10474), .Z(n10434) );
  AND U10493 ( .A(n10475), .B(n10476), .Z(n10474) );
  XOR U10494 ( .A(n10473), .B(n10477), .Z(n10475) );
  XNOR U10495 ( .A(n10478), .B(n10479), .Z(n10472) );
  AND U10496 ( .A(n10480), .B(n10481), .Z(n10479) );
  XOR U10497 ( .A(n10478), .B(n10482), .Z(n10480) );
  XOR U10498 ( .A(n10483), .B(n10484), .Z(n10438) );
  AND U10499 ( .A(n10485), .B(n10486), .Z(n10484) );
  XOR U10500 ( .A(n10483), .B(n10487), .Z(n10485) );
  XNOR U10501 ( .A(n10374), .B(n10444), .Z(n10446) );
  XNOR U10502 ( .A(n10488), .B(n10489), .Z(n10374) );
  AND U10503 ( .A(n344), .B(n10490), .Z(n10489) );
  XNOR U10504 ( .A(n10491), .B(n10492), .Z(n10490) );
  XOR U10505 ( .A(n10493), .B(n10494), .Z(n10444) );
  AND U10506 ( .A(n10495), .B(n10496), .Z(n10494) );
  XNOR U10507 ( .A(n10493), .B(n10385), .Z(n10496) );
  XOR U10508 ( .A(n10497), .B(n10458), .Z(n10385) );
  XNOR U10509 ( .A(n10498), .B(n10465), .Z(n10458) );
  XOR U10510 ( .A(n10454), .B(n10453), .Z(n10465) );
  XNOR U10511 ( .A(n10499), .B(n10450), .Z(n10453) );
  XOR U10512 ( .A(n10500), .B(n10501), .Z(n10450) );
  AND U10513 ( .A(n10502), .B(n10503), .Z(n10501) );
  XNOR U10514 ( .A(n10504), .B(n10505), .Z(n10502) );
  IV U10515 ( .A(n10500), .Z(n10504) );
  XNOR U10516 ( .A(n10506), .B(n10507), .Z(n10499) );
  NOR U10517 ( .A(n10508), .B(n10509), .Z(n10507) );
  XNOR U10518 ( .A(n10506), .B(n10510), .Z(n10508) );
  XOR U10519 ( .A(n10511), .B(n10512), .Z(n10454) );
  NOR U10520 ( .A(n10513), .B(n10514), .Z(n10512) );
  XNOR U10521 ( .A(n10511), .B(n10515), .Z(n10513) );
  XNOR U10522 ( .A(n10464), .B(n10455), .Z(n10498) );
  XOR U10523 ( .A(n10516), .B(n10517), .Z(n10455) );
  AND U10524 ( .A(n10518), .B(n10519), .Z(n10517) );
  XOR U10525 ( .A(n10516), .B(n10520), .Z(n10518) );
  XOR U10526 ( .A(n10521), .B(n10470), .Z(n10464) );
  XOR U10527 ( .A(n10522), .B(n10523), .Z(n10470) );
  NOR U10528 ( .A(n10524), .B(n10525), .Z(n10523) );
  XOR U10529 ( .A(n10522), .B(n10526), .Z(n10524) );
  XNOR U10530 ( .A(n10469), .B(n10461), .Z(n10521) );
  XOR U10531 ( .A(n10527), .B(n10528), .Z(n10461) );
  AND U10532 ( .A(n10529), .B(n10530), .Z(n10528) );
  XOR U10533 ( .A(n10527), .B(n10531), .Z(n10529) );
  XNOR U10534 ( .A(n10532), .B(n10466), .Z(n10469) );
  XOR U10535 ( .A(n10533), .B(n10534), .Z(n10466) );
  AND U10536 ( .A(n10535), .B(n10536), .Z(n10534) );
  XNOR U10537 ( .A(n10537), .B(n10538), .Z(n10535) );
  IV U10538 ( .A(n10533), .Z(n10537) );
  XNOR U10539 ( .A(n10539), .B(n10540), .Z(n10532) );
  NOR U10540 ( .A(n10541), .B(n10542), .Z(n10540) );
  XNOR U10541 ( .A(n10539), .B(n10543), .Z(n10541) );
  XOR U10542 ( .A(n10459), .B(n10471), .Z(n10497) );
  NOR U10543 ( .A(n10391), .B(n10544), .Z(n10471) );
  XNOR U10544 ( .A(n10477), .B(n10476), .Z(n10459) );
  XNOR U10545 ( .A(n10545), .B(n10482), .Z(n10476) );
  XNOR U10546 ( .A(n10546), .B(n10547), .Z(n10482) );
  NOR U10547 ( .A(n10548), .B(n10549), .Z(n10547) );
  XOR U10548 ( .A(n10546), .B(n10550), .Z(n10548) );
  XNOR U10549 ( .A(n10481), .B(n10473), .Z(n10545) );
  XOR U10550 ( .A(n10551), .B(n10552), .Z(n10473) );
  AND U10551 ( .A(n10553), .B(n10554), .Z(n10552) );
  XOR U10552 ( .A(n10551), .B(n10555), .Z(n10553) );
  XNOR U10553 ( .A(n10556), .B(n10478), .Z(n10481) );
  XOR U10554 ( .A(n10557), .B(n10558), .Z(n10478) );
  AND U10555 ( .A(n10559), .B(n10560), .Z(n10558) );
  XNOR U10556 ( .A(n10561), .B(n10562), .Z(n10559) );
  IV U10557 ( .A(n10557), .Z(n10561) );
  XNOR U10558 ( .A(n10563), .B(n10564), .Z(n10556) );
  NOR U10559 ( .A(n10565), .B(n10566), .Z(n10564) );
  XNOR U10560 ( .A(n10563), .B(n10567), .Z(n10565) );
  XOR U10561 ( .A(n10487), .B(n10486), .Z(n10477) );
  XNOR U10562 ( .A(n10568), .B(n10483), .Z(n10486) );
  XOR U10563 ( .A(n10569), .B(n10570), .Z(n10483) );
  AND U10564 ( .A(n10571), .B(n10572), .Z(n10570) );
  XNOR U10565 ( .A(n10573), .B(n10574), .Z(n10571) );
  IV U10566 ( .A(n10569), .Z(n10573) );
  XNOR U10567 ( .A(n10575), .B(n10576), .Z(n10568) );
  NOR U10568 ( .A(n10577), .B(n10578), .Z(n10576) );
  XNOR U10569 ( .A(n10575), .B(n10579), .Z(n10577) );
  XOR U10570 ( .A(n10580), .B(n10581), .Z(n10487) );
  NOR U10571 ( .A(n10582), .B(n10583), .Z(n10581) );
  XNOR U10572 ( .A(n10580), .B(n10584), .Z(n10582) );
  XNOR U10573 ( .A(n10382), .B(n10493), .Z(n10495) );
  XNOR U10574 ( .A(n10585), .B(n10586), .Z(n10382) );
  AND U10575 ( .A(n344), .B(n10587), .Z(n10586) );
  XNOR U10576 ( .A(n10588), .B(n10589), .Z(n10587) );
  AND U10577 ( .A(n10388), .B(n10391), .Z(n10493) );
  XOR U10578 ( .A(n10590), .B(n10544), .Z(n10391) );
  XNOR U10579 ( .A(p_input[352]), .B(p_input[512]), .Z(n10544) );
  XNOR U10580 ( .A(n10520), .B(n10519), .Z(n10590) );
  XNOR U10581 ( .A(n10591), .B(n10531), .Z(n10519) );
  XOR U10582 ( .A(n10505), .B(n10503), .Z(n10531) );
  XNOR U10583 ( .A(n10592), .B(n10510), .Z(n10503) );
  XOR U10584 ( .A(p_input[376]), .B(p_input[536]), .Z(n10510) );
  XOR U10585 ( .A(n10500), .B(n10509), .Z(n10592) );
  XOR U10586 ( .A(n10593), .B(n10506), .Z(n10509) );
  XOR U10587 ( .A(p_input[374]), .B(p_input[534]), .Z(n10506) );
  XOR U10588 ( .A(p_input[375]), .B(n6576), .Z(n10593) );
  XOR U10589 ( .A(p_input[370]), .B(p_input[530]), .Z(n10500) );
  XNOR U10590 ( .A(n10515), .B(n10514), .Z(n10505) );
  XOR U10591 ( .A(n10594), .B(n10511), .Z(n10514) );
  XOR U10592 ( .A(p_input[371]), .B(p_input[531]), .Z(n10511) );
  XOR U10593 ( .A(p_input[372]), .B(n6578), .Z(n10594) );
  XOR U10594 ( .A(p_input[373]), .B(p_input[533]), .Z(n10515) );
  XOR U10595 ( .A(n10530), .B(n10595), .Z(n10591) );
  IV U10596 ( .A(n10516), .Z(n10595) );
  XOR U10597 ( .A(p_input[353]), .B(p_input[513]), .Z(n10516) );
  XNOR U10598 ( .A(n10596), .B(n10538), .Z(n10530) );
  XNOR U10599 ( .A(n10526), .B(n10525), .Z(n10538) );
  XNOR U10600 ( .A(n10597), .B(n10522), .Z(n10525) );
  XNOR U10601 ( .A(p_input[378]), .B(p_input[538]), .Z(n10522) );
  XOR U10602 ( .A(p_input[379]), .B(n6582), .Z(n10597) );
  XOR U10603 ( .A(p_input[380]), .B(p_input[540]), .Z(n10526) );
  XOR U10604 ( .A(n10536), .B(n10598), .Z(n10596) );
  IV U10605 ( .A(n10527), .Z(n10598) );
  XOR U10606 ( .A(p_input[369]), .B(p_input[529]), .Z(n10527) );
  XNOR U10607 ( .A(n10599), .B(n10543), .Z(n10536) );
  XNOR U10608 ( .A(p_input[383]), .B(n6585), .Z(n10543) );
  XOR U10609 ( .A(n10533), .B(n10542), .Z(n10599) );
  XOR U10610 ( .A(n10600), .B(n10539), .Z(n10542) );
  XOR U10611 ( .A(p_input[381]), .B(p_input[541]), .Z(n10539) );
  XOR U10612 ( .A(p_input[382]), .B(n6587), .Z(n10600) );
  XOR U10613 ( .A(p_input[377]), .B(p_input[537]), .Z(n10533) );
  XOR U10614 ( .A(n10555), .B(n10554), .Z(n10520) );
  XNOR U10615 ( .A(n10601), .B(n10562), .Z(n10554) );
  XNOR U10616 ( .A(n10550), .B(n10549), .Z(n10562) );
  XNOR U10617 ( .A(n10602), .B(n10546), .Z(n10549) );
  XNOR U10618 ( .A(p_input[363]), .B(p_input[523]), .Z(n10546) );
  XOR U10619 ( .A(p_input[364]), .B(n6590), .Z(n10602) );
  XOR U10620 ( .A(p_input[365]), .B(p_input[525]), .Z(n10550) );
  XOR U10621 ( .A(n10560), .B(n10603), .Z(n10601) );
  IV U10622 ( .A(n10551), .Z(n10603) );
  XOR U10623 ( .A(p_input[354]), .B(p_input[514]), .Z(n10551) );
  XNOR U10624 ( .A(n10604), .B(n10567), .Z(n10560) );
  XNOR U10625 ( .A(p_input[368]), .B(n6593), .Z(n10567) );
  XOR U10626 ( .A(n10557), .B(n10566), .Z(n10604) );
  XOR U10627 ( .A(n10605), .B(n10563), .Z(n10566) );
  XOR U10628 ( .A(p_input[366]), .B(p_input[526]), .Z(n10563) );
  XOR U10629 ( .A(p_input[367]), .B(n6595), .Z(n10605) );
  XOR U10630 ( .A(p_input[362]), .B(p_input[522]), .Z(n10557) );
  XOR U10631 ( .A(n10574), .B(n10572), .Z(n10555) );
  XNOR U10632 ( .A(n10606), .B(n10579), .Z(n10572) );
  XOR U10633 ( .A(p_input[361]), .B(p_input[521]), .Z(n10579) );
  XOR U10634 ( .A(n10569), .B(n10578), .Z(n10606) );
  XOR U10635 ( .A(n10607), .B(n10575), .Z(n10578) );
  XOR U10636 ( .A(p_input[359]), .B(p_input[519]), .Z(n10575) );
  XOR U10637 ( .A(p_input[360]), .B(n6963), .Z(n10607) );
  XOR U10638 ( .A(p_input[355]), .B(p_input[515]), .Z(n10569) );
  XNOR U10639 ( .A(n10584), .B(n10583), .Z(n10574) );
  XOR U10640 ( .A(n10608), .B(n10580), .Z(n10583) );
  XOR U10641 ( .A(p_input[356]), .B(p_input[516]), .Z(n10580) );
  XOR U10642 ( .A(p_input[357]), .B(n6965), .Z(n10608) );
  XOR U10643 ( .A(p_input[358]), .B(p_input[518]), .Z(n10584) );
  XNOR U10644 ( .A(n10609), .B(n10610), .Z(n10388) );
  AND U10645 ( .A(n344), .B(n10611), .Z(n10610) );
  XNOR U10646 ( .A(n10612), .B(n10613), .Z(n344) );
  NOR U10647 ( .A(n10614), .B(n10615), .Z(n10613) );
  XNOR U10648 ( .A(n10612), .B(n10616), .Z(n10615) );
  NOR U10649 ( .A(n10612), .B(n10397), .Z(n10614) );
  XOR U10650 ( .A(n10617), .B(n10618), .Z(n10612) );
  AND U10651 ( .A(n10619), .B(n10620), .Z(n10618) );
  XOR U10652 ( .A(n10414), .B(n10617), .Z(n10620) );
  XOR U10653 ( .A(n10617), .B(n10415), .Z(n10619) );
  XOR U10654 ( .A(n10621), .B(n10622), .Z(n10617) );
  AND U10655 ( .A(n10623), .B(n10624), .Z(n10622) );
  XOR U10656 ( .A(n10442), .B(n10621), .Z(n10624) );
  XOR U10657 ( .A(n10621), .B(n10443), .Z(n10623) );
  XOR U10658 ( .A(n10625), .B(n10626), .Z(n10621) );
  AND U10659 ( .A(n10627), .B(n10628), .Z(n10626) );
  XOR U10660 ( .A(n10491), .B(n10625), .Z(n10628) );
  XOR U10661 ( .A(n10625), .B(n10492), .Z(n10627) );
  XOR U10662 ( .A(n10629), .B(n10630), .Z(n10625) );
  AND U10663 ( .A(n10631), .B(n10632), .Z(n10630) );
  XOR U10664 ( .A(n10629), .B(n10588), .Z(n10632) );
  XNOR U10665 ( .A(n10633), .B(n10634), .Z(n10341) );
  AND U10666 ( .A(n348), .B(n10635), .Z(n10634) );
  XNOR U10667 ( .A(n10636), .B(n10637), .Z(n348) );
  NOR U10668 ( .A(n10638), .B(n10639), .Z(n10637) );
  XOR U10669 ( .A(n10303), .B(n10636), .Z(n10639) );
  NOR U10670 ( .A(n10636), .B(n10302), .Z(n10638) );
  XOR U10671 ( .A(n10640), .B(n10641), .Z(n10636) );
  AND U10672 ( .A(n10642), .B(n10643), .Z(n10641) );
  XNOR U10673 ( .A(n10358), .B(n10640), .Z(n10643) );
  XOR U10674 ( .A(n10640), .B(n10311), .Z(n10642) );
  XOR U10675 ( .A(n10644), .B(n10645), .Z(n10640) );
  AND U10676 ( .A(n10646), .B(n10647), .Z(n10645) );
  XNOR U10677 ( .A(n10368), .B(n10644), .Z(n10647) );
  XOR U10678 ( .A(n10644), .B(n10320), .Z(n10646) );
  XOR U10679 ( .A(n10648), .B(n10649), .Z(n10644) );
  AND U10680 ( .A(n10650), .B(n10651), .Z(n10649) );
  XOR U10681 ( .A(n10648), .B(n10328), .Z(n10650) );
  XOR U10682 ( .A(n10652), .B(n10653), .Z(n10295) );
  AND U10683 ( .A(n352), .B(n10635), .Z(n10653) );
  XNOR U10684 ( .A(n10633), .B(n10652), .Z(n10635) );
  XNOR U10685 ( .A(n10654), .B(n10655), .Z(n352) );
  NOR U10686 ( .A(n10656), .B(n10657), .Z(n10655) );
  XNOR U10687 ( .A(n10303), .B(n10658), .Z(n10657) );
  IV U10688 ( .A(n10654), .Z(n10658) );
  AND U10689 ( .A(n10659), .B(n10660), .Z(n10303) );
  NOR U10690 ( .A(n10654), .B(n10302), .Z(n10656) );
  AND U10691 ( .A(n10397), .B(n10396), .Z(n10302) );
  IV U10692 ( .A(n10616), .Z(n10396) );
  XOR U10693 ( .A(n10661), .B(n10662), .Z(n10654) );
  AND U10694 ( .A(n10663), .B(n10664), .Z(n10662) );
  XNOR U10695 ( .A(n10661), .B(n10358), .Z(n10664) );
  XOR U10696 ( .A(n10415), .B(n10665), .Z(n10358) );
  AND U10697 ( .A(n355), .B(n10666), .Z(n10665) );
  XOR U10698 ( .A(n10411), .B(n10415), .Z(n10666) );
  XNOR U10699 ( .A(n10667), .B(n10661), .Z(n10663) );
  IV U10700 ( .A(n10311), .Z(n10667) );
  XOR U10701 ( .A(n10668), .B(n10669), .Z(n10311) );
  AND U10702 ( .A(n370), .B(n10670), .Z(n10669) );
  XOR U10703 ( .A(n10671), .B(n10672), .Z(n10661) );
  AND U10704 ( .A(n10673), .B(n10674), .Z(n10672) );
  XNOR U10705 ( .A(n10671), .B(n10368), .Z(n10674) );
  XOR U10706 ( .A(n10443), .B(n10675), .Z(n10368) );
  AND U10707 ( .A(n355), .B(n10676), .Z(n10675) );
  XOR U10708 ( .A(n10439), .B(n10443), .Z(n10676) );
  XOR U10709 ( .A(n10320), .B(n10671), .Z(n10673) );
  XOR U10710 ( .A(n10677), .B(n10678), .Z(n10320) );
  AND U10711 ( .A(n370), .B(n10679), .Z(n10678) );
  XOR U10712 ( .A(n10648), .B(n10680), .Z(n10671) );
  AND U10713 ( .A(n10681), .B(n10651), .Z(n10680) );
  XNOR U10714 ( .A(n10378), .B(n10648), .Z(n10651) );
  XOR U10715 ( .A(n10492), .B(n10682), .Z(n10378) );
  AND U10716 ( .A(n355), .B(n10683), .Z(n10682) );
  XOR U10717 ( .A(n10488), .B(n10492), .Z(n10683) );
  XNOR U10718 ( .A(n10684), .B(n10648), .Z(n10681) );
  IV U10719 ( .A(n10328), .Z(n10684) );
  XOR U10720 ( .A(n10685), .B(n10686), .Z(n10328) );
  AND U10721 ( .A(n370), .B(n10687), .Z(n10686) );
  XOR U10722 ( .A(n10688), .B(n10689), .Z(n10648) );
  AND U10723 ( .A(n10690), .B(n10691), .Z(n10689) );
  XNOR U10724 ( .A(n10688), .B(n10386), .Z(n10691) );
  XOR U10725 ( .A(n10589), .B(n10692), .Z(n10386) );
  AND U10726 ( .A(n355), .B(n10693), .Z(n10692) );
  XOR U10727 ( .A(n10585), .B(n10589), .Z(n10693) );
  XNOR U10728 ( .A(n10694), .B(n10688), .Z(n10690) );
  IV U10729 ( .A(n10338), .Z(n10694) );
  XOR U10730 ( .A(n10695), .B(n10696), .Z(n10338) );
  AND U10731 ( .A(n370), .B(n10697), .Z(n10696) );
  AND U10732 ( .A(n10652), .B(n10633), .Z(n10688) );
  XNOR U10733 ( .A(n10698), .B(n10699), .Z(n10633) );
  AND U10734 ( .A(n355), .B(n10611), .Z(n10699) );
  XNOR U10735 ( .A(n10609), .B(n10698), .Z(n10611) );
  XNOR U10736 ( .A(n10700), .B(n10701), .Z(n355) );
  NOR U10737 ( .A(n10702), .B(n10703), .Z(n10701) );
  XNOR U10738 ( .A(n10700), .B(n10616), .Z(n10703) );
  NOR U10739 ( .A(n10659), .B(n10660), .Z(n10616) );
  NOR U10740 ( .A(n10700), .B(n10397), .Z(n10702) );
  AND U10741 ( .A(n10704), .B(n10705), .Z(n10397) );
  IV U10742 ( .A(n10706), .Z(n10704) );
  XOR U10743 ( .A(n10707), .B(n10708), .Z(n10700) );
  AND U10744 ( .A(n10709), .B(n10710), .Z(n10708) );
  XNOR U10745 ( .A(n10707), .B(n10411), .Z(n10710) );
  IV U10746 ( .A(n10414), .Z(n10411) );
  XOR U10747 ( .A(n10711), .B(n10712), .Z(n10414) );
  AND U10748 ( .A(n359), .B(n10713), .Z(n10712) );
  XOR U10749 ( .A(n10714), .B(n10711), .Z(n10713) );
  XOR U10750 ( .A(n10415), .B(n10707), .Z(n10709) );
  XOR U10751 ( .A(n10715), .B(n10716), .Z(n10415) );
  AND U10752 ( .A(n366), .B(n10670), .Z(n10716) );
  XOR U10753 ( .A(n10715), .B(n10668), .Z(n10670) );
  XOR U10754 ( .A(n10717), .B(n10718), .Z(n10707) );
  AND U10755 ( .A(n10719), .B(n10720), .Z(n10718) );
  XNOR U10756 ( .A(n10717), .B(n10439), .Z(n10720) );
  IV U10757 ( .A(n10442), .Z(n10439) );
  XOR U10758 ( .A(n10721), .B(n10722), .Z(n10442) );
  AND U10759 ( .A(n359), .B(n10723), .Z(n10722) );
  XNOR U10760 ( .A(n10724), .B(n10721), .Z(n10723) );
  XOR U10761 ( .A(n10443), .B(n10717), .Z(n10719) );
  XOR U10762 ( .A(n10725), .B(n10726), .Z(n10443) );
  AND U10763 ( .A(n366), .B(n10679), .Z(n10726) );
  XOR U10764 ( .A(n10725), .B(n10677), .Z(n10679) );
  XOR U10765 ( .A(n10727), .B(n10728), .Z(n10717) );
  AND U10766 ( .A(n10729), .B(n10730), .Z(n10728) );
  XNOR U10767 ( .A(n10727), .B(n10488), .Z(n10730) );
  IV U10768 ( .A(n10491), .Z(n10488) );
  XOR U10769 ( .A(n10731), .B(n10732), .Z(n10491) );
  AND U10770 ( .A(n359), .B(n10733), .Z(n10732) );
  XOR U10771 ( .A(n10734), .B(n10731), .Z(n10733) );
  XOR U10772 ( .A(n10492), .B(n10727), .Z(n10729) );
  XOR U10773 ( .A(n10735), .B(n10736), .Z(n10492) );
  AND U10774 ( .A(n366), .B(n10687), .Z(n10736) );
  XOR U10775 ( .A(n10735), .B(n10685), .Z(n10687) );
  XOR U10776 ( .A(n10629), .B(n10737), .Z(n10727) );
  AND U10777 ( .A(n10631), .B(n10738), .Z(n10737) );
  XNOR U10778 ( .A(n10629), .B(n10585), .Z(n10738) );
  IV U10779 ( .A(n10588), .Z(n10585) );
  XOR U10780 ( .A(n10739), .B(n10740), .Z(n10588) );
  AND U10781 ( .A(n359), .B(n10741), .Z(n10740) );
  XNOR U10782 ( .A(n10742), .B(n10739), .Z(n10741) );
  XOR U10783 ( .A(n10589), .B(n10629), .Z(n10631) );
  XOR U10784 ( .A(n10743), .B(n10744), .Z(n10589) );
  AND U10785 ( .A(n366), .B(n10697), .Z(n10744) );
  XOR U10786 ( .A(n10743), .B(n10695), .Z(n10697) );
  AND U10787 ( .A(n10698), .B(n10609), .Z(n10629) );
  XNOR U10788 ( .A(n10745), .B(n10746), .Z(n10609) );
  AND U10789 ( .A(n359), .B(n10747), .Z(n10746) );
  XNOR U10790 ( .A(n10748), .B(n10745), .Z(n10747) );
  XNOR U10791 ( .A(n10749), .B(n10750), .Z(n359) );
  NOR U10792 ( .A(n10751), .B(n10752), .Z(n10750) );
  XNOR U10793 ( .A(n10749), .B(n10706), .Z(n10752) );
  NOR U10794 ( .A(n10753), .B(n10754), .Z(n10706) );
  NOR U10795 ( .A(n10749), .B(n10705), .Z(n10751) );
  AND U10796 ( .A(n10755), .B(n10756), .Z(n10705) );
  XOR U10797 ( .A(n10757), .B(n10758), .Z(n10749) );
  AND U10798 ( .A(n10759), .B(n10760), .Z(n10758) );
  XNOR U10799 ( .A(n10757), .B(n10755), .Z(n10760) );
  IV U10800 ( .A(n10714), .Z(n10755) );
  XOR U10801 ( .A(n10761), .B(n10762), .Z(n10714) );
  XOR U10802 ( .A(n10763), .B(n10756), .Z(n10762) );
  AND U10803 ( .A(n10724), .B(n10764), .Z(n10756) );
  AND U10804 ( .A(n10765), .B(n10766), .Z(n10763) );
  XOR U10805 ( .A(n10767), .B(n10761), .Z(n10765) );
  XNOR U10806 ( .A(n10711), .B(n10757), .Z(n10759) );
  XNOR U10807 ( .A(n10768), .B(n10769), .Z(n10711) );
  AND U10808 ( .A(n362), .B(n10770), .Z(n10769) );
  XOR U10809 ( .A(n10771), .B(n10772), .Z(n10757) );
  AND U10810 ( .A(n10773), .B(n10774), .Z(n10772) );
  XNOR U10811 ( .A(n10771), .B(n10724), .Z(n10774) );
  XOR U10812 ( .A(n10775), .B(n10766), .Z(n10724) );
  XNOR U10813 ( .A(n10776), .B(n10761), .Z(n10766) );
  XOR U10814 ( .A(n10777), .B(n10778), .Z(n10761) );
  AND U10815 ( .A(n10779), .B(n10780), .Z(n10778) );
  XOR U10816 ( .A(n10781), .B(n10777), .Z(n10779) );
  XNOR U10817 ( .A(n10782), .B(n10783), .Z(n10776) );
  AND U10818 ( .A(n10784), .B(n10785), .Z(n10783) );
  XOR U10819 ( .A(n10782), .B(n10786), .Z(n10784) );
  XNOR U10820 ( .A(n10767), .B(n10764), .Z(n10775) );
  AND U10821 ( .A(n10787), .B(n10788), .Z(n10764) );
  XOR U10822 ( .A(n10789), .B(n10790), .Z(n10767) );
  AND U10823 ( .A(n10791), .B(n10792), .Z(n10790) );
  XOR U10824 ( .A(n10789), .B(n10793), .Z(n10791) );
  XNOR U10825 ( .A(n10721), .B(n10771), .Z(n10773) );
  XNOR U10826 ( .A(n10794), .B(n10795), .Z(n10721) );
  AND U10827 ( .A(n362), .B(n10796), .Z(n10795) );
  XOR U10828 ( .A(n10797), .B(n10798), .Z(n10771) );
  AND U10829 ( .A(n10799), .B(n10800), .Z(n10798) );
  XNOR U10830 ( .A(n10797), .B(n10787), .Z(n10800) );
  IV U10831 ( .A(n10734), .Z(n10787) );
  XNOR U10832 ( .A(n10801), .B(n10780), .Z(n10734) );
  XNOR U10833 ( .A(n10802), .B(n10786), .Z(n10780) );
  XOR U10834 ( .A(n10803), .B(n10804), .Z(n10786) );
  AND U10835 ( .A(n10805), .B(n10806), .Z(n10804) );
  XOR U10836 ( .A(n10803), .B(n10807), .Z(n10805) );
  XNOR U10837 ( .A(n10785), .B(n10777), .Z(n10802) );
  XOR U10838 ( .A(n10808), .B(n10809), .Z(n10777) );
  AND U10839 ( .A(n10810), .B(n10811), .Z(n10809) );
  XNOR U10840 ( .A(n10812), .B(n10808), .Z(n10810) );
  XNOR U10841 ( .A(n10813), .B(n10782), .Z(n10785) );
  XOR U10842 ( .A(n10814), .B(n10815), .Z(n10782) );
  AND U10843 ( .A(n10816), .B(n10817), .Z(n10815) );
  XOR U10844 ( .A(n10814), .B(n10818), .Z(n10816) );
  XNOR U10845 ( .A(n10819), .B(n10820), .Z(n10813) );
  AND U10846 ( .A(n10821), .B(n10822), .Z(n10820) );
  XNOR U10847 ( .A(n10819), .B(n10823), .Z(n10821) );
  XNOR U10848 ( .A(n10781), .B(n10788), .Z(n10801) );
  AND U10849 ( .A(n10742), .B(n10824), .Z(n10788) );
  XOR U10850 ( .A(n10793), .B(n10792), .Z(n10781) );
  XNOR U10851 ( .A(n10825), .B(n10789), .Z(n10792) );
  XOR U10852 ( .A(n10826), .B(n10827), .Z(n10789) );
  AND U10853 ( .A(n10828), .B(n10829), .Z(n10827) );
  XOR U10854 ( .A(n10826), .B(n10830), .Z(n10828) );
  XNOR U10855 ( .A(n10831), .B(n10832), .Z(n10825) );
  AND U10856 ( .A(n10833), .B(n10834), .Z(n10832) );
  XOR U10857 ( .A(n10831), .B(n10835), .Z(n10833) );
  XOR U10858 ( .A(n10836), .B(n10837), .Z(n10793) );
  AND U10859 ( .A(n10838), .B(n10839), .Z(n10837) );
  XOR U10860 ( .A(n10836), .B(n10840), .Z(n10838) );
  XNOR U10861 ( .A(n10731), .B(n10797), .Z(n10799) );
  XNOR U10862 ( .A(n10841), .B(n10842), .Z(n10731) );
  AND U10863 ( .A(n362), .B(n10843), .Z(n10842) );
  XNOR U10864 ( .A(n10844), .B(n10845), .Z(n10843) );
  XOR U10865 ( .A(n10846), .B(n10847), .Z(n10797) );
  AND U10866 ( .A(n10848), .B(n10849), .Z(n10847) );
  XNOR U10867 ( .A(n10846), .B(n10742), .Z(n10849) );
  XOR U10868 ( .A(n10850), .B(n10811), .Z(n10742) );
  XNOR U10869 ( .A(n10851), .B(n10818), .Z(n10811) );
  XOR U10870 ( .A(n10807), .B(n10806), .Z(n10818) );
  XNOR U10871 ( .A(n10852), .B(n10803), .Z(n10806) );
  XOR U10872 ( .A(n10853), .B(n10854), .Z(n10803) );
  AND U10873 ( .A(n10855), .B(n10856), .Z(n10854) );
  XNOR U10874 ( .A(n10857), .B(n10858), .Z(n10855) );
  IV U10875 ( .A(n10853), .Z(n10857) );
  XNOR U10876 ( .A(n10859), .B(n10860), .Z(n10852) );
  NOR U10877 ( .A(n10861), .B(n10862), .Z(n10860) );
  XNOR U10878 ( .A(n10859), .B(n10863), .Z(n10861) );
  XOR U10879 ( .A(n10864), .B(n10865), .Z(n10807) );
  NOR U10880 ( .A(n10866), .B(n10867), .Z(n10865) );
  XNOR U10881 ( .A(n10864), .B(n10868), .Z(n10866) );
  XNOR U10882 ( .A(n10817), .B(n10808), .Z(n10851) );
  XOR U10883 ( .A(n10869), .B(n10870), .Z(n10808) );
  AND U10884 ( .A(n10871), .B(n10872), .Z(n10870) );
  XOR U10885 ( .A(n10869), .B(n10873), .Z(n10871) );
  XOR U10886 ( .A(n10874), .B(n10823), .Z(n10817) );
  XOR U10887 ( .A(n10875), .B(n10876), .Z(n10823) );
  NOR U10888 ( .A(n10877), .B(n10878), .Z(n10876) );
  XOR U10889 ( .A(n10875), .B(n10879), .Z(n10877) );
  XNOR U10890 ( .A(n10822), .B(n10814), .Z(n10874) );
  XOR U10891 ( .A(n10880), .B(n10881), .Z(n10814) );
  AND U10892 ( .A(n10882), .B(n10883), .Z(n10881) );
  XOR U10893 ( .A(n10880), .B(n10884), .Z(n10882) );
  XNOR U10894 ( .A(n10885), .B(n10819), .Z(n10822) );
  XOR U10895 ( .A(n10886), .B(n10887), .Z(n10819) );
  AND U10896 ( .A(n10888), .B(n10889), .Z(n10887) );
  XNOR U10897 ( .A(n10890), .B(n10891), .Z(n10888) );
  IV U10898 ( .A(n10886), .Z(n10890) );
  XNOR U10899 ( .A(n10892), .B(n10893), .Z(n10885) );
  NOR U10900 ( .A(n10894), .B(n10895), .Z(n10893) );
  XNOR U10901 ( .A(n10892), .B(n10896), .Z(n10894) );
  XOR U10902 ( .A(n10812), .B(n10824), .Z(n10850) );
  NOR U10903 ( .A(n10748), .B(n10897), .Z(n10824) );
  XNOR U10904 ( .A(n10830), .B(n10829), .Z(n10812) );
  XNOR U10905 ( .A(n10898), .B(n10835), .Z(n10829) );
  XNOR U10906 ( .A(n10899), .B(n10900), .Z(n10835) );
  NOR U10907 ( .A(n10901), .B(n10902), .Z(n10900) );
  XOR U10908 ( .A(n10899), .B(n10903), .Z(n10901) );
  XNOR U10909 ( .A(n10834), .B(n10826), .Z(n10898) );
  XOR U10910 ( .A(n10904), .B(n10905), .Z(n10826) );
  AND U10911 ( .A(n10906), .B(n10907), .Z(n10905) );
  XOR U10912 ( .A(n10904), .B(n10908), .Z(n10906) );
  XNOR U10913 ( .A(n10909), .B(n10831), .Z(n10834) );
  XOR U10914 ( .A(n10910), .B(n10911), .Z(n10831) );
  AND U10915 ( .A(n10912), .B(n10913), .Z(n10911) );
  XNOR U10916 ( .A(n10914), .B(n10915), .Z(n10912) );
  IV U10917 ( .A(n10910), .Z(n10914) );
  XNOR U10918 ( .A(n10916), .B(n10917), .Z(n10909) );
  NOR U10919 ( .A(n10918), .B(n10919), .Z(n10917) );
  XNOR U10920 ( .A(n10916), .B(n10920), .Z(n10918) );
  XOR U10921 ( .A(n10840), .B(n10839), .Z(n10830) );
  XNOR U10922 ( .A(n10921), .B(n10836), .Z(n10839) );
  XOR U10923 ( .A(n10922), .B(n10923), .Z(n10836) );
  AND U10924 ( .A(n10924), .B(n10925), .Z(n10923) );
  XNOR U10925 ( .A(n10926), .B(n10927), .Z(n10924) );
  IV U10926 ( .A(n10922), .Z(n10926) );
  XNOR U10927 ( .A(n10928), .B(n10929), .Z(n10921) );
  NOR U10928 ( .A(n10930), .B(n10931), .Z(n10929) );
  XNOR U10929 ( .A(n10928), .B(n10932), .Z(n10930) );
  XOR U10930 ( .A(n10933), .B(n10934), .Z(n10840) );
  NOR U10931 ( .A(n10935), .B(n10936), .Z(n10934) );
  XNOR U10932 ( .A(n10933), .B(n10937), .Z(n10935) );
  XNOR U10933 ( .A(n10739), .B(n10846), .Z(n10848) );
  XNOR U10934 ( .A(n10938), .B(n10939), .Z(n10739) );
  AND U10935 ( .A(n362), .B(n10940), .Z(n10939) );
  AND U10936 ( .A(n10745), .B(n10748), .Z(n10846) );
  XOR U10937 ( .A(n10941), .B(n10897), .Z(n10748) );
  XNOR U10938 ( .A(p_input[384]), .B(p_input[512]), .Z(n10897) );
  XNOR U10939 ( .A(n10873), .B(n10872), .Z(n10941) );
  XNOR U10940 ( .A(n10942), .B(n10884), .Z(n10872) );
  XOR U10941 ( .A(n10858), .B(n10856), .Z(n10884) );
  XNOR U10942 ( .A(n10943), .B(n10863), .Z(n10856) );
  XOR U10943 ( .A(p_input[408]), .B(p_input[536]), .Z(n10863) );
  XOR U10944 ( .A(n10853), .B(n10862), .Z(n10943) );
  XOR U10945 ( .A(n10944), .B(n10859), .Z(n10862) );
  XOR U10946 ( .A(p_input[406]), .B(p_input[534]), .Z(n10859) );
  XOR U10947 ( .A(p_input[407]), .B(n6576), .Z(n10944) );
  XOR U10948 ( .A(p_input[402]), .B(p_input[530]), .Z(n10853) );
  XNOR U10949 ( .A(n10868), .B(n10867), .Z(n10858) );
  XOR U10950 ( .A(n10945), .B(n10864), .Z(n10867) );
  XOR U10951 ( .A(p_input[403]), .B(p_input[531]), .Z(n10864) );
  XOR U10952 ( .A(p_input[404]), .B(n6578), .Z(n10945) );
  XOR U10953 ( .A(p_input[405]), .B(p_input[533]), .Z(n10868) );
  XOR U10954 ( .A(n10883), .B(n10946), .Z(n10942) );
  IV U10955 ( .A(n10869), .Z(n10946) );
  XOR U10956 ( .A(p_input[385]), .B(p_input[513]), .Z(n10869) );
  XNOR U10957 ( .A(n10947), .B(n10891), .Z(n10883) );
  XNOR U10958 ( .A(n10879), .B(n10878), .Z(n10891) );
  XNOR U10959 ( .A(n10948), .B(n10875), .Z(n10878) );
  XNOR U10960 ( .A(p_input[410]), .B(p_input[538]), .Z(n10875) );
  XOR U10961 ( .A(p_input[411]), .B(n6582), .Z(n10948) );
  XOR U10962 ( .A(p_input[412]), .B(p_input[540]), .Z(n10879) );
  XOR U10963 ( .A(n10889), .B(n10949), .Z(n10947) );
  IV U10964 ( .A(n10880), .Z(n10949) );
  XOR U10965 ( .A(p_input[401]), .B(p_input[529]), .Z(n10880) );
  XNOR U10966 ( .A(n10950), .B(n10896), .Z(n10889) );
  XNOR U10967 ( .A(p_input[415]), .B(n6585), .Z(n10896) );
  IV U10968 ( .A(p_input[543]), .Z(n6585) );
  XOR U10969 ( .A(n10886), .B(n10895), .Z(n10950) );
  XOR U10970 ( .A(n10951), .B(n10892), .Z(n10895) );
  XOR U10971 ( .A(p_input[413]), .B(p_input[541]), .Z(n10892) );
  XOR U10972 ( .A(p_input[414]), .B(n6587), .Z(n10951) );
  XOR U10973 ( .A(p_input[409]), .B(p_input[537]), .Z(n10886) );
  XOR U10974 ( .A(n10908), .B(n10907), .Z(n10873) );
  XNOR U10975 ( .A(n10952), .B(n10915), .Z(n10907) );
  XNOR U10976 ( .A(n10903), .B(n10902), .Z(n10915) );
  XNOR U10977 ( .A(n10953), .B(n10899), .Z(n10902) );
  XNOR U10978 ( .A(p_input[395]), .B(p_input[523]), .Z(n10899) );
  XOR U10979 ( .A(p_input[396]), .B(n6590), .Z(n10953) );
  XOR U10980 ( .A(p_input[397]), .B(p_input[525]), .Z(n10903) );
  XOR U10981 ( .A(n10913), .B(n10954), .Z(n10952) );
  IV U10982 ( .A(n10904), .Z(n10954) );
  XOR U10983 ( .A(p_input[386]), .B(p_input[514]), .Z(n10904) );
  XNOR U10984 ( .A(n10955), .B(n10920), .Z(n10913) );
  XNOR U10985 ( .A(p_input[400]), .B(n6593), .Z(n10920) );
  IV U10986 ( .A(p_input[528]), .Z(n6593) );
  XOR U10987 ( .A(n10910), .B(n10919), .Z(n10955) );
  XOR U10988 ( .A(n10956), .B(n10916), .Z(n10919) );
  XOR U10989 ( .A(p_input[398]), .B(p_input[526]), .Z(n10916) );
  XOR U10990 ( .A(p_input[399]), .B(n6595), .Z(n10956) );
  XOR U10991 ( .A(p_input[394]), .B(p_input[522]), .Z(n10910) );
  XOR U10992 ( .A(n10927), .B(n10925), .Z(n10908) );
  XNOR U10993 ( .A(n10957), .B(n10932), .Z(n10925) );
  XOR U10994 ( .A(p_input[393]), .B(p_input[521]), .Z(n10932) );
  XOR U10995 ( .A(n10922), .B(n10931), .Z(n10957) );
  XOR U10996 ( .A(n10958), .B(n10928), .Z(n10931) );
  XOR U10997 ( .A(p_input[391]), .B(p_input[519]), .Z(n10928) );
  XOR U10998 ( .A(p_input[392]), .B(n6963), .Z(n10958) );
  XOR U10999 ( .A(p_input[387]), .B(p_input[515]), .Z(n10922) );
  XNOR U11000 ( .A(n10937), .B(n10936), .Z(n10927) );
  XOR U11001 ( .A(n10959), .B(n10933), .Z(n10936) );
  XOR U11002 ( .A(p_input[388]), .B(p_input[516]), .Z(n10933) );
  XOR U11003 ( .A(p_input[389]), .B(n6965), .Z(n10959) );
  XOR U11004 ( .A(p_input[390]), .B(p_input[518]), .Z(n10937) );
  XNOR U11005 ( .A(n10960), .B(n10961), .Z(n10745) );
  AND U11006 ( .A(n362), .B(n10962), .Z(n10961) );
  XNOR U11007 ( .A(n10963), .B(n10964), .Z(n362) );
  NOR U11008 ( .A(n10965), .B(n10966), .Z(n10964) );
  XOR U11009 ( .A(n10963), .B(n10753), .Z(n10966) );
  XNOR U11010 ( .A(n10967), .B(n10968), .Z(n10698) );
  AND U11011 ( .A(n366), .B(n10969), .Z(n10968) );
  XNOR U11012 ( .A(n10970), .B(n10971), .Z(n366) );
  NOR U11013 ( .A(n10972), .B(n10973), .Z(n10971) );
  XOR U11014 ( .A(n10660), .B(n10970), .Z(n10973) );
  NOR U11015 ( .A(n10970), .B(n10659), .Z(n10972) );
  XOR U11016 ( .A(n10974), .B(n10975), .Z(n10970) );
  AND U11017 ( .A(n10976), .B(n10977), .Z(n10975) );
  XNOR U11018 ( .A(n10715), .B(n10974), .Z(n10977) );
  XOR U11019 ( .A(n10974), .B(n10668), .Z(n10976) );
  XOR U11020 ( .A(n10978), .B(n10979), .Z(n10974) );
  AND U11021 ( .A(n10980), .B(n10981), .Z(n10979) );
  XNOR U11022 ( .A(n10725), .B(n10978), .Z(n10981) );
  XOR U11023 ( .A(n10978), .B(n10677), .Z(n10980) );
  XOR U11024 ( .A(n10982), .B(n10983), .Z(n10978) );
  AND U11025 ( .A(n10984), .B(n10985), .Z(n10983) );
  XOR U11026 ( .A(n10982), .B(n10685), .Z(n10984) );
  XOR U11027 ( .A(n10986), .B(n10987), .Z(n10652) );
  AND U11028 ( .A(n370), .B(n10969), .Z(n10987) );
  XNOR U11029 ( .A(n10967), .B(n10986), .Z(n10969) );
  XNOR U11030 ( .A(n10988), .B(n10989), .Z(n370) );
  NOR U11031 ( .A(n10990), .B(n10991), .Z(n10989) );
  XNOR U11032 ( .A(n10660), .B(n10992), .Z(n10991) );
  IV U11033 ( .A(n10988), .Z(n10992) );
  AND U11034 ( .A(n10993), .B(n10994), .Z(n10660) );
  NOR U11035 ( .A(n10988), .B(n10659), .Z(n10990) );
  AND U11036 ( .A(n10753), .B(n10754), .Z(n10659) );
  IV U11037 ( .A(n10995), .Z(n10753) );
  XOR U11038 ( .A(n10996), .B(n10997), .Z(n10988) );
  AND U11039 ( .A(n10998), .B(n10999), .Z(n10997) );
  XNOR U11040 ( .A(n10996), .B(n10715), .Z(n10999) );
  XOR U11041 ( .A(n11000), .B(n11001), .Z(n10715) );
  AND U11042 ( .A(n373), .B(n10770), .Z(n11001) );
  XOR U11043 ( .A(n10768), .B(n11000), .Z(n10770) );
  XNOR U11044 ( .A(n11002), .B(n10996), .Z(n10998) );
  IV U11045 ( .A(n10668), .Z(n11002) );
  XOR U11046 ( .A(n11003), .B(n11004), .Z(n10668) );
  AND U11047 ( .A(n378), .B(n11005), .Z(n11004) );
  XOR U11048 ( .A(n11006), .B(n11007), .Z(n10996) );
  AND U11049 ( .A(n11008), .B(n11009), .Z(n11007) );
  XNOR U11050 ( .A(n11006), .B(n10725), .Z(n11009) );
  XOR U11051 ( .A(n11010), .B(n11011), .Z(n10725) );
  AND U11052 ( .A(n373), .B(n10796), .Z(n11011) );
  XOR U11053 ( .A(n10794), .B(n11010), .Z(n10796) );
  XOR U11054 ( .A(n10677), .B(n11006), .Z(n11008) );
  XOR U11055 ( .A(n11012), .B(n11013), .Z(n10677) );
  AND U11056 ( .A(n378), .B(n11014), .Z(n11013) );
  XOR U11057 ( .A(n10982), .B(n11015), .Z(n11006) );
  AND U11058 ( .A(n11016), .B(n10985), .Z(n11015) );
  XNOR U11059 ( .A(n10735), .B(n10982), .Z(n10985) );
  XOR U11060 ( .A(n10845), .B(n11017), .Z(n10735) );
  AND U11061 ( .A(n373), .B(n11018), .Z(n11017) );
  XOR U11062 ( .A(n10841), .B(n10845), .Z(n11018) );
  XNOR U11063 ( .A(n11019), .B(n10982), .Z(n11016) );
  IV U11064 ( .A(n10685), .Z(n11019) );
  XOR U11065 ( .A(n11020), .B(n11021), .Z(n10685) );
  AND U11066 ( .A(n378), .B(n11022), .Z(n11021) );
  XOR U11067 ( .A(n11023), .B(n11024), .Z(n10982) );
  AND U11068 ( .A(n11025), .B(n11026), .Z(n11024) );
  XNOR U11069 ( .A(n11023), .B(n10743), .Z(n11026) );
  XNOR U11070 ( .A(n11027), .B(n11028), .Z(n10743) );
  AND U11071 ( .A(n373), .B(n10940), .Z(n11028) );
  XOR U11072 ( .A(n10938), .B(n11029), .Z(n10940) );
  IV U11073 ( .A(n11027), .Z(n11029) );
  XNOR U11074 ( .A(n11030), .B(n11023), .Z(n11025) );
  IV U11075 ( .A(n10695), .Z(n11030) );
  XOR U11076 ( .A(n11031), .B(n11032), .Z(n10695) );
  AND U11077 ( .A(n378), .B(n11033), .Z(n11032) );
  AND U11078 ( .A(n10986), .B(n10967), .Z(n11023) );
  XNOR U11079 ( .A(n11034), .B(n11035), .Z(n10967) );
  AND U11080 ( .A(n373), .B(n10962), .Z(n11035) );
  XOR U11081 ( .A(n11036), .B(n11034), .Z(n10962) );
  XNOR U11082 ( .A(n10963), .B(n11037), .Z(n373) );
  NOR U11083 ( .A(n10965), .B(n11038), .Z(n11037) );
  XNOR U11084 ( .A(n10963), .B(n10995), .Z(n11038) );
  NOR U11085 ( .A(n10993), .B(n10994), .Z(n10995) );
  NOR U11086 ( .A(n10963), .B(n10754), .Z(n10965) );
  AND U11087 ( .A(n10768), .B(n11039), .Z(n10754) );
  XOR U11088 ( .A(n11040), .B(n11041), .Z(n10963) );
  AND U11089 ( .A(n11042), .B(n11043), .Z(n11041) );
  XNOR U11090 ( .A(n10768), .B(n11040), .Z(n11043) );
  XNOR U11091 ( .A(n11044), .B(n11045), .Z(n10768) );
  XOR U11092 ( .A(n11046), .B(n11039), .Z(n11045) );
  AND U11093 ( .A(n10794), .B(n11047), .Z(n11039) );
  AND U11094 ( .A(n11048), .B(n11049), .Z(n11046) );
  XOR U11095 ( .A(n11050), .B(n11044), .Z(n11048) );
  XOR U11096 ( .A(n11040), .B(n11000), .Z(n11042) );
  XOR U11097 ( .A(n11051), .B(n11052), .Z(n11000) );
  AND U11098 ( .A(n375), .B(n11005), .Z(n11052) );
  XOR U11099 ( .A(n11051), .B(n11003), .Z(n11005) );
  XOR U11100 ( .A(n11053), .B(n11054), .Z(n11040) );
  AND U11101 ( .A(n11055), .B(n11056), .Z(n11054) );
  XNOR U11102 ( .A(n10794), .B(n11053), .Z(n11056) );
  XOR U11103 ( .A(n11057), .B(n11049), .Z(n10794) );
  XNOR U11104 ( .A(n11058), .B(n11044), .Z(n11049) );
  XOR U11105 ( .A(n11059), .B(n11060), .Z(n11044) );
  AND U11106 ( .A(n11061), .B(n11062), .Z(n11060) );
  XOR U11107 ( .A(n11063), .B(n11059), .Z(n11061) );
  XNOR U11108 ( .A(n11064), .B(n11065), .Z(n11058) );
  AND U11109 ( .A(n11066), .B(n11067), .Z(n11065) );
  XOR U11110 ( .A(n11064), .B(n11068), .Z(n11066) );
  XNOR U11111 ( .A(n11050), .B(n11047), .Z(n11057) );
  AND U11112 ( .A(n10841), .B(n11069), .Z(n11047) );
  XOR U11113 ( .A(n11070), .B(n11071), .Z(n11050) );
  AND U11114 ( .A(n11072), .B(n11073), .Z(n11071) );
  XOR U11115 ( .A(n11070), .B(n11074), .Z(n11072) );
  XOR U11116 ( .A(n11053), .B(n11010), .Z(n11055) );
  XOR U11117 ( .A(n11075), .B(n11076), .Z(n11010) );
  AND U11118 ( .A(n375), .B(n11014), .Z(n11076) );
  XOR U11119 ( .A(n11075), .B(n11012), .Z(n11014) );
  XOR U11120 ( .A(n11077), .B(n11078), .Z(n11053) );
  AND U11121 ( .A(n11079), .B(n11080), .Z(n11078) );
  XNOR U11122 ( .A(n10841), .B(n11077), .Z(n11080) );
  IV U11123 ( .A(n10844), .Z(n10841) );
  XNOR U11124 ( .A(n11081), .B(n11062), .Z(n10844) );
  XNOR U11125 ( .A(n11082), .B(n11068), .Z(n11062) );
  XOR U11126 ( .A(n11083), .B(n11084), .Z(n11068) );
  AND U11127 ( .A(n11085), .B(n11086), .Z(n11084) );
  XOR U11128 ( .A(n11083), .B(n11087), .Z(n11085) );
  XNOR U11129 ( .A(n11067), .B(n11059), .Z(n11082) );
  XOR U11130 ( .A(n11088), .B(n11089), .Z(n11059) );
  AND U11131 ( .A(n11090), .B(n11091), .Z(n11089) );
  XNOR U11132 ( .A(n11092), .B(n11088), .Z(n11090) );
  XNOR U11133 ( .A(n11093), .B(n11064), .Z(n11067) );
  XOR U11134 ( .A(n11094), .B(n11095), .Z(n11064) );
  AND U11135 ( .A(n11096), .B(n11097), .Z(n11095) );
  XOR U11136 ( .A(n11094), .B(n11098), .Z(n11096) );
  XNOR U11137 ( .A(n11099), .B(n11100), .Z(n11093) );
  AND U11138 ( .A(n11101), .B(n11102), .Z(n11100) );
  XNOR U11139 ( .A(n11099), .B(n11103), .Z(n11101) );
  XNOR U11140 ( .A(n11063), .B(n11069), .Z(n11081) );
  AND U11141 ( .A(n10938), .B(n11104), .Z(n11069) );
  XOR U11142 ( .A(n11074), .B(n11073), .Z(n11063) );
  XNOR U11143 ( .A(n11105), .B(n11070), .Z(n11073) );
  XOR U11144 ( .A(n11106), .B(n11107), .Z(n11070) );
  AND U11145 ( .A(n11108), .B(n11109), .Z(n11107) );
  XOR U11146 ( .A(n11106), .B(n11110), .Z(n11108) );
  XNOR U11147 ( .A(n11111), .B(n11112), .Z(n11105) );
  AND U11148 ( .A(n11113), .B(n11114), .Z(n11112) );
  XOR U11149 ( .A(n11111), .B(n11115), .Z(n11113) );
  XOR U11150 ( .A(n11116), .B(n11117), .Z(n11074) );
  AND U11151 ( .A(n11118), .B(n11119), .Z(n11117) );
  XOR U11152 ( .A(n11116), .B(n11120), .Z(n11118) );
  XOR U11153 ( .A(n11077), .B(n10845), .Z(n11079) );
  XOR U11154 ( .A(n11121), .B(n11122), .Z(n10845) );
  AND U11155 ( .A(n375), .B(n11022), .Z(n11122) );
  XOR U11156 ( .A(n11121), .B(n11020), .Z(n11022) );
  XOR U11157 ( .A(n11123), .B(n11124), .Z(n11077) );
  AND U11158 ( .A(n11125), .B(n11126), .Z(n11124) );
  XNOR U11159 ( .A(n11123), .B(n10938), .Z(n11126) );
  XOR U11160 ( .A(n11127), .B(n11091), .Z(n10938) );
  XNOR U11161 ( .A(n11128), .B(n11098), .Z(n11091) );
  XOR U11162 ( .A(n11087), .B(n11086), .Z(n11098) );
  XNOR U11163 ( .A(n11129), .B(n11083), .Z(n11086) );
  XOR U11164 ( .A(n11130), .B(n11131), .Z(n11083) );
  AND U11165 ( .A(n11132), .B(n11133), .Z(n11131) );
  XOR U11166 ( .A(n11130), .B(n11134), .Z(n11132) );
  XNOR U11167 ( .A(n11135), .B(n11136), .Z(n11129) );
  NOR U11168 ( .A(n11137), .B(n11138), .Z(n11136) );
  XNOR U11169 ( .A(n11135), .B(n11139), .Z(n11137) );
  XOR U11170 ( .A(n11140), .B(n11141), .Z(n11087) );
  NOR U11171 ( .A(n11142), .B(n11143), .Z(n11141) );
  XNOR U11172 ( .A(n11140), .B(n11144), .Z(n11142) );
  XNOR U11173 ( .A(n11097), .B(n11088), .Z(n11128) );
  XOR U11174 ( .A(n11145), .B(n11146), .Z(n11088) );
  NOR U11175 ( .A(n11147), .B(n11148), .Z(n11146) );
  XNOR U11176 ( .A(n11145), .B(n11149), .Z(n11147) );
  XOR U11177 ( .A(n11150), .B(n11103), .Z(n11097) );
  XNOR U11178 ( .A(n11151), .B(n11152), .Z(n11103) );
  NOR U11179 ( .A(n11153), .B(n11154), .Z(n11152) );
  XNOR U11180 ( .A(n11151), .B(n11155), .Z(n11153) );
  XNOR U11181 ( .A(n11102), .B(n11094), .Z(n11150) );
  XOR U11182 ( .A(n11156), .B(n11157), .Z(n11094) );
  AND U11183 ( .A(n11158), .B(n11159), .Z(n11157) );
  XOR U11184 ( .A(n11156), .B(n11160), .Z(n11158) );
  XNOR U11185 ( .A(n11161), .B(n11099), .Z(n11102) );
  XOR U11186 ( .A(n11162), .B(n11163), .Z(n11099) );
  AND U11187 ( .A(n11164), .B(n11165), .Z(n11163) );
  XOR U11188 ( .A(n11162), .B(n11166), .Z(n11164) );
  XNOR U11189 ( .A(n11167), .B(n11168), .Z(n11161) );
  NOR U11190 ( .A(n11169), .B(n11170), .Z(n11168) );
  XOR U11191 ( .A(n11167), .B(n11171), .Z(n11169) );
  XOR U11192 ( .A(n11092), .B(n11104), .Z(n11127) );
  AND U11193 ( .A(n11036), .B(n11172), .Z(n11104) );
  IV U11194 ( .A(n10960), .Z(n11036) );
  XNOR U11195 ( .A(n11110), .B(n11109), .Z(n11092) );
  XNOR U11196 ( .A(n11173), .B(n11115), .Z(n11109) );
  XOR U11197 ( .A(n11174), .B(n11175), .Z(n11115) );
  NOR U11198 ( .A(n11176), .B(n11177), .Z(n11175) );
  XNOR U11199 ( .A(n11174), .B(n11178), .Z(n11176) );
  XNOR U11200 ( .A(n11114), .B(n11106), .Z(n11173) );
  XOR U11201 ( .A(n11179), .B(n11180), .Z(n11106) );
  AND U11202 ( .A(n11181), .B(n11182), .Z(n11180) );
  XNOR U11203 ( .A(n11179), .B(n11183), .Z(n11181) );
  XNOR U11204 ( .A(n11184), .B(n11111), .Z(n11114) );
  XOR U11205 ( .A(n11185), .B(n11186), .Z(n11111) );
  AND U11206 ( .A(n11187), .B(n11188), .Z(n11186) );
  XOR U11207 ( .A(n11185), .B(n11189), .Z(n11187) );
  XNOR U11208 ( .A(n11190), .B(n11191), .Z(n11184) );
  NOR U11209 ( .A(n11192), .B(n11193), .Z(n11191) );
  XOR U11210 ( .A(n11190), .B(n11194), .Z(n11192) );
  XOR U11211 ( .A(n11120), .B(n11119), .Z(n11110) );
  XNOR U11212 ( .A(n11195), .B(n11116), .Z(n11119) );
  XOR U11213 ( .A(n11196), .B(n11197), .Z(n11116) );
  AND U11214 ( .A(n11198), .B(n11199), .Z(n11197) );
  XOR U11215 ( .A(n11196), .B(n11200), .Z(n11198) );
  XNOR U11216 ( .A(n11201), .B(n11202), .Z(n11195) );
  NOR U11217 ( .A(n11203), .B(n11204), .Z(n11202) );
  XNOR U11218 ( .A(n11201), .B(n11205), .Z(n11203) );
  XOR U11219 ( .A(n11206), .B(n11207), .Z(n11120) );
  NOR U11220 ( .A(n11208), .B(n11209), .Z(n11207) );
  XNOR U11221 ( .A(n11206), .B(n11210), .Z(n11208) );
  XNOR U11222 ( .A(n11027), .B(n11123), .Z(n11125) );
  XNOR U11223 ( .A(n11211), .B(n11212), .Z(n11027) );
  AND U11224 ( .A(n375), .B(n11033), .Z(n11212) );
  XOR U11225 ( .A(n11211), .B(n11031), .Z(n11033) );
  AND U11226 ( .A(n11034), .B(n10960), .Z(n11123) );
  XNOR U11227 ( .A(n11213), .B(n11172), .Z(n10960) );
  XOR U11228 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][0] ), .B(
        p_input[512]), .Z(n11172) );
  XOR U11229 ( .A(n11149), .B(n11148), .Z(n11213) );
  XOR U11230 ( .A(n11214), .B(n11160), .Z(n11148) );
  XOR U11231 ( .A(n11134), .B(n11133), .Z(n11160) );
  XNOR U11232 ( .A(n11215), .B(n11139), .Z(n11133) );
  XOR U11233 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][24] ), .B(
        p_input[536]), .Z(n11139) );
  XOR U11234 ( .A(n11130), .B(n11138), .Z(n11215) );
  XOR U11235 ( .A(n11216), .B(n11135), .Z(n11138) );
  XOR U11236 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][22] ), .B(
        p_input[534]), .Z(n11135) );
  XOR U11237 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][23] ), .B(n6576), 
        .Z(n11216) );
  XNOR U11238 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][18] ), .B(n7313), 
        .Z(n11130) );
  XNOR U11239 ( .A(n11144), .B(n11143), .Z(n11134) );
  XOR U11240 ( .A(n11217), .B(n11140), .Z(n11143) );
  XOR U11241 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][19] ), .B(
        p_input[531]), .Z(n11140) );
  XOR U11242 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][20] ), .B(n6578), 
        .Z(n11217) );
  XOR U11243 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][21] ), .B(
        p_input[533]), .Z(n11144) );
  XNOR U11244 ( .A(n11159), .B(n11145), .Z(n11214) );
  XNOR U11245 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][1] ), .B(n7315), 
        .Z(n11145) );
  XNOR U11246 ( .A(n11218), .B(n11166), .Z(n11159) );
  XNOR U11247 ( .A(n11155), .B(n11154), .Z(n11166) );
  XOR U11248 ( .A(n11219), .B(n11151), .Z(n11154) );
  XNOR U11249 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][26] ), .B(n6951), 
        .Z(n11151) );
  XOR U11250 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][27] ), .B(n6582), 
        .Z(n11219) );
  XOR U11251 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][28] ), .B(
        p_input[540]), .Z(n11155) );
  XNOR U11252 ( .A(n11165), .B(n11156), .Z(n11218) );
  XNOR U11253 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][17] ), .B(n7318), 
        .Z(n11156) );
  XOR U11254 ( .A(n11220), .B(n11171), .Z(n11165) );
  XNOR U11255 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][31] ), .B(
        p_input[543]), .Z(n11171) );
  XOR U11256 ( .A(n11162), .B(n11170), .Z(n11220) );
  XOR U11257 ( .A(n11221), .B(n11167), .Z(n11170) );
  XOR U11258 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][29] ), .B(
        p_input[541]), .Z(n11167) );
  XOR U11259 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][30] ), .B(n6587), 
        .Z(n11221) );
  XNOR U11260 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][25] ), .B(n6955), 
        .Z(n11162) );
  XNOR U11261 ( .A(n11183), .B(n11182), .Z(n11149) );
  XNOR U11262 ( .A(n11222), .B(n11189), .Z(n11182) );
  XNOR U11263 ( .A(n11178), .B(n11177), .Z(n11189) );
  XOR U11264 ( .A(n11223), .B(n11174), .Z(n11177) );
  XNOR U11265 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][11] ), .B(n7323), 
        .Z(n11174) );
  XOR U11266 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][12] ), .B(n6590), 
        .Z(n11223) );
  XOR U11267 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][13] ), .B(
        p_input[525]), .Z(n11178) );
  XNOR U11268 ( .A(n11188), .B(n11179), .Z(n11222) );
  XNOR U11269 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][2] ), .B(n7324), 
        .Z(n11179) );
  XOR U11270 ( .A(n11224), .B(n11194), .Z(n11188) );
  XNOR U11271 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][16] ), .B(
        p_input[528]), .Z(n11194) );
  XOR U11272 ( .A(n11185), .B(n11193), .Z(n11224) );
  XOR U11273 ( .A(n11225), .B(n11190), .Z(n11193) );
  XOR U11274 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][14] ), .B(
        p_input[526]), .Z(n11190) );
  XOR U11275 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][15] ), .B(n6595), 
        .Z(n11225) );
  XNOR U11276 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][10] ), .B(n7327), 
        .Z(n11185) );
  XNOR U11277 ( .A(n11200), .B(n11199), .Z(n11183) );
  XNOR U11278 ( .A(n11226), .B(n11205), .Z(n11199) );
  XOR U11279 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][9] ), .B(
        p_input[521]), .Z(n11205) );
  XOR U11280 ( .A(n11196), .B(n11204), .Z(n11226) );
  XOR U11281 ( .A(n11227), .B(n11201), .Z(n11204) );
  XOR U11282 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][7] ), .B(
        p_input[519]), .Z(n11201) );
  XOR U11283 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][8] ), .B(n6963), 
        .Z(n11227) );
  XNOR U11284 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][3] ), .B(n7330), 
        .Z(n11196) );
  XNOR U11285 ( .A(n11210), .B(n11209), .Z(n11200) );
  XOR U11286 ( .A(n11228), .B(n11206), .Z(n11209) );
  XOR U11287 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][4] ), .B(
        p_input[516]), .Z(n11206) );
  XOR U11288 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][5] ), .B(n6965), 
        .Z(n11228) );
  XOR U11289 ( .A(\knn_comb_/ASN_1[2].knn_/local_min_val[2][6] ), .B(
        p_input[518]), .Z(n11210) );
  XNOR U11290 ( .A(n11229), .B(n11230), .Z(n11034) );
  AND U11291 ( .A(n375), .B(n11231), .Z(n11230) );
  XNOR U11292 ( .A(n11232), .B(n11233), .Z(n375) );
  NOR U11293 ( .A(n11234), .B(n11235), .Z(n11233) );
  XOR U11294 ( .A(n10994), .B(n11232), .Z(n11235) );
  NOR U11295 ( .A(n11232), .B(n10993), .Z(n11234) );
  XOR U11296 ( .A(n11236), .B(n11237), .Z(n11232) );
  AND U11297 ( .A(n11238), .B(n11239), .Z(n11237) );
  XNOR U11298 ( .A(n11051), .B(n11236), .Z(n11239) );
  XOR U11299 ( .A(n11236), .B(n11003), .Z(n11238) );
  XOR U11300 ( .A(n11240), .B(n11241), .Z(n11236) );
  AND U11301 ( .A(n11242), .B(n11243), .Z(n11241) );
  XNOR U11302 ( .A(n11075), .B(n11240), .Z(n11243) );
  XOR U11303 ( .A(n11240), .B(n11012), .Z(n11242) );
  XOR U11304 ( .A(n11244), .B(n11245), .Z(n11240) );
  AND U11305 ( .A(n11246), .B(n11247), .Z(n11245) );
  XOR U11306 ( .A(n11244), .B(n11020), .Z(n11246) );
  XOR U11307 ( .A(n11248), .B(n11249), .Z(n10986) );
  AND U11308 ( .A(n378), .B(n11231), .Z(n11249) );
  XOR U11309 ( .A(n11250), .B(n11248), .Z(n11231) );
  XNOR U11310 ( .A(n11251), .B(n11252), .Z(n378) );
  NOR U11311 ( .A(n11253), .B(n11254), .Z(n11252) );
  XNOR U11312 ( .A(n10994), .B(n11255), .Z(n11254) );
  IV U11313 ( .A(n11251), .Z(n11255) );
  AND U11314 ( .A(n11003), .B(n11256), .Z(n10994) );
  NOR U11315 ( .A(n11251), .B(n10993), .Z(n11253) );
  AND U11316 ( .A(n11051), .B(n11257), .Z(n10993) );
  XOR U11317 ( .A(n11258), .B(n11259), .Z(n11251) );
  AND U11318 ( .A(n11260), .B(n11261), .Z(n11259) );
  XNOR U11319 ( .A(n11258), .B(n11051), .Z(n11261) );
  XNOR U11320 ( .A(n11262), .B(n11263), .Z(n11051) );
  XOR U11321 ( .A(n11264), .B(n11257), .Z(n11263) );
  AND U11322 ( .A(n11075), .B(n11265), .Z(n11257) );
  AND U11323 ( .A(n11266), .B(n11267), .Z(n11264) );
  XOR U11324 ( .A(n11268), .B(n11262), .Z(n11266) );
  XNOR U11325 ( .A(n11269), .B(n11258), .Z(n11260) );
  IV U11326 ( .A(n11003), .Z(n11269) );
  XNOR U11327 ( .A(n11270), .B(n11271), .Z(n11003) );
  XOR U11328 ( .A(n11272), .B(n11256), .Z(n11271) );
  AND U11329 ( .A(n11012), .B(n11273), .Z(n11256) );
  AND U11330 ( .A(n11274), .B(n11275), .Z(n11272) );
  XNOR U11331 ( .A(n11270), .B(n11276), .Z(n11274) );
  XOR U11332 ( .A(n11277), .B(n11278), .Z(n11258) );
  AND U11333 ( .A(n11279), .B(n11280), .Z(n11278) );
  XNOR U11334 ( .A(n11277), .B(n11075), .Z(n11280) );
  XOR U11335 ( .A(n11281), .B(n11267), .Z(n11075) );
  XNOR U11336 ( .A(n11282), .B(n11262), .Z(n11267) );
  XOR U11337 ( .A(n11283), .B(n11284), .Z(n11262) );
  AND U11338 ( .A(n11285), .B(n11286), .Z(n11284) );
  XOR U11339 ( .A(n11287), .B(n11283), .Z(n11285) );
  XNOR U11340 ( .A(n11288), .B(n11289), .Z(n11282) );
  AND U11341 ( .A(n11290), .B(n11291), .Z(n11289) );
  XOR U11342 ( .A(n11288), .B(n11292), .Z(n11290) );
  XNOR U11343 ( .A(n11268), .B(n11265), .Z(n11281) );
  AND U11344 ( .A(n11121), .B(n11293), .Z(n11265) );
  XOR U11345 ( .A(n11294), .B(n11295), .Z(n11268) );
  AND U11346 ( .A(n11296), .B(n11297), .Z(n11295) );
  XOR U11347 ( .A(n11294), .B(n11298), .Z(n11296) );
  XOR U11348 ( .A(n11012), .B(n11277), .Z(n11279) );
  XNOR U11349 ( .A(n11299), .B(n11276), .Z(n11012) );
  XNOR U11350 ( .A(n11300), .B(n11301), .Z(n11276) );
  AND U11351 ( .A(n11302), .B(n11303), .Z(n11301) );
  XOR U11352 ( .A(n11300), .B(n11304), .Z(n11302) );
  XNOR U11353 ( .A(n11275), .B(n11273), .Z(n11299) );
  AND U11354 ( .A(n11020), .B(n11305), .Z(n11273) );
  XNOR U11355 ( .A(n11306), .B(n11270), .Z(n11275) );
  XOR U11356 ( .A(n11307), .B(n11308), .Z(n11270) );
  AND U11357 ( .A(n11309), .B(n11310), .Z(n11308) );
  XOR U11358 ( .A(n11307), .B(n11311), .Z(n11309) );
  XNOR U11359 ( .A(n11312), .B(n11313), .Z(n11306) );
  AND U11360 ( .A(n11314), .B(n11315), .Z(n11313) );
  XNOR U11361 ( .A(n11312), .B(n11316), .Z(n11314) );
  XOR U11362 ( .A(n11244), .B(n11317), .Z(n11277) );
  AND U11363 ( .A(n11318), .B(n11247), .Z(n11317) );
  XNOR U11364 ( .A(n11121), .B(n11244), .Z(n11247) );
  XOR U11365 ( .A(n11319), .B(n11286), .Z(n11121) );
  XNOR U11366 ( .A(n11320), .B(n11292), .Z(n11286) );
  XOR U11367 ( .A(n11321), .B(n11322), .Z(n11292) );
  AND U11368 ( .A(n11323), .B(n11324), .Z(n11322) );
  XOR U11369 ( .A(n11321), .B(n11325), .Z(n11323) );
  XNOR U11370 ( .A(n11291), .B(n11283), .Z(n11320) );
  XOR U11371 ( .A(n11326), .B(n11327), .Z(n11283) );
  AND U11372 ( .A(n11328), .B(n11329), .Z(n11327) );
  XNOR U11373 ( .A(n11330), .B(n11326), .Z(n11328) );
  XNOR U11374 ( .A(n11331), .B(n11288), .Z(n11291) );
  XOR U11375 ( .A(n11332), .B(n11333), .Z(n11288) );
  AND U11376 ( .A(n11334), .B(n11335), .Z(n11333) );
  XOR U11377 ( .A(n11332), .B(n11336), .Z(n11334) );
  XNOR U11378 ( .A(n11337), .B(n11338), .Z(n11331) );
  AND U11379 ( .A(n11339), .B(n11340), .Z(n11338) );
  XNOR U11380 ( .A(n11337), .B(n11341), .Z(n11339) );
  XNOR U11381 ( .A(n11287), .B(n11293), .Z(n11319) );
  AND U11382 ( .A(n11211), .B(n11342), .Z(n11293) );
  XOR U11383 ( .A(n11298), .B(n11297), .Z(n11287) );
  XNOR U11384 ( .A(n11343), .B(n11294), .Z(n11297) );
  XOR U11385 ( .A(n11344), .B(n11345), .Z(n11294) );
  AND U11386 ( .A(n11346), .B(n11347), .Z(n11345) );
  XOR U11387 ( .A(n11344), .B(n11348), .Z(n11346) );
  XNOR U11388 ( .A(n11349), .B(n11350), .Z(n11343) );
  AND U11389 ( .A(n11351), .B(n11352), .Z(n11350) );
  XOR U11390 ( .A(n11349), .B(n11353), .Z(n11351) );
  XOR U11391 ( .A(n11354), .B(n11355), .Z(n11298) );
  AND U11392 ( .A(n11356), .B(n11357), .Z(n11355) );
  XOR U11393 ( .A(n11354), .B(n11358), .Z(n11356) );
  XNOR U11394 ( .A(n11359), .B(n11244), .Z(n11318) );
  IV U11395 ( .A(n11020), .Z(n11359) );
  XOR U11396 ( .A(n11360), .B(n11311), .Z(n11020) );
  XOR U11397 ( .A(n11304), .B(n11303), .Z(n11311) );
  XNOR U11398 ( .A(n11361), .B(n11300), .Z(n11303) );
  XOR U11399 ( .A(n11362), .B(n11363), .Z(n11300) );
  AND U11400 ( .A(n11364), .B(n11365), .Z(n11363) );
  XOR U11401 ( .A(n11362), .B(n11366), .Z(n11364) );
  XNOR U11402 ( .A(n11367), .B(n11368), .Z(n11361) );
  AND U11403 ( .A(n11369), .B(n11370), .Z(n11368) );
  XOR U11404 ( .A(n11367), .B(n11371), .Z(n11369) );
  XOR U11405 ( .A(n11372), .B(n11373), .Z(n11304) );
  AND U11406 ( .A(n11374), .B(n11375), .Z(n11373) );
  XOR U11407 ( .A(n11372), .B(n11376), .Z(n11374) );
  XNOR U11408 ( .A(n11310), .B(n11305), .Z(n11360) );
  AND U11409 ( .A(n11031), .B(n11377), .Z(n11305) );
  XOR U11410 ( .A(n11378), .B(n11316), .Z(n11310) );
  XNOR U11411 ( .A(n11379), .B(n11380), .Z(n11316) );
  AND U11412 ( .A(n11381), .B(n11382), .Z(n11380) );
  XOR U11413 ( .A(n11379), .B(n11383), .Z(n11381) );
  XNOR U11414 ( .A(n11315), .B(n11307), .Z(n11378) );
  XOR U11415 ( .A(n11384), .B(n11385), .Z(n11307) );
  AND U11416 ( .A(n11386), .B(n11387), .Z(n11385) );
  XOR U11417 ( .A(n11384), .B(n11388), .Z(n11386) );
  XNOR U11418 ( .A(n11389), .B(n11312), .Z(n11315) );
  XOR U11419 ( .A(n11390), .B(n11391), .Z(n11312) );
  AND U11420 ( .A(n11392), .B(n11393), .Z(n11391) );
  XOR U11421 ( .A(n11390), .B(n11394), .Z(n11392) );
  XNOR U11422 ( .A(n11395), .B(n11396), .Z(n11389) );
  AND U11423 ( .A(n11397), .B(n11398), .Z(n11396) );
  XNOR U11424 ( .A(n11395), .B(n11399), .Z(n11397) );
  XOR U11425 ( .A(n11400), .B(n11401), .Z(n11244) );
  AND U11426 ( .A(n11402), .B(n11403), .Z(n11401) );
  XNOR U11427 ( .A(n11400), .B(n11211), .Z(n11403) );
  XOR U11428 ( .A(n11404), .B(n11329), .Z(n11211) );
  XNOR U11429 ( .A(n11405), .B(n11336), .Z(n11329) );
  XOR U11430 ( .A(n11325), .B(n11324), .Z(n11336) );
  XNOR U11431 ( .A(n11406), .B(n11321), .Z(n11324) );
  XOR U11432 ( .A(n11407), .B(n11408), .Z(n11321) );
  AND U11433 ( .A(n11409), .B(n11410), .Z(n11408) );
  XOR U11434 ( .A(n11407), .B(n11411), .Z(n11409) );
  XNOR U11435 ( .A(n11412), .B(n11413), .Z(n11406) );
  NOR U11436 ( .A(n11414), .B(n11415), .Z(n11413) );
  XNOR U11437 ( .A(n11412), .B(n11416), .Z(n11414) );
  XOR U11438 ( .A(n11417), .B(n11418), .Z(n11325) );
  NOR U11439 ( .A(n11419), .B(n11420), .Z(n11418) );
  XNOR U11440 ( .A(n11417), .B(n11421), .Z(n11419) );
  XNOR U11441 ( .A(n11335), .B(n11326), .Z(n11405) );
  XOR U11442 ( .A(n11422), .B(n11423), .Z(n11326) );
  NOR U11443 ( .A(n11424), .B(n11425), .Z(n11423) );
  XNOR U11444 ( .A(n11422), .B(n11426), .Z(n11424) );
  XOR U11445 ( .A(n11427), .B(n11341), .Z(n11335) );
  XNOR U11446 ( .A(n11428), .B(n11429), .Z(n11341) );
  NOR U11447 ( .A(n11430), .B(n11431), .Z(n11429) );
  XNOR U11448 ( .A(n11428), .B(n11432), .Z(n11430) );
  XNOR U11449 ( .A(n11340), .B(n11332), .Z(n11427) );
  XOR U11450 ( .A(n11433), .B(n11434), .Z(n11332) );
  AND U11451 ( .A(n11435), .B(n11436), .Z(n11434) );
  XOR U11452 ( .A(n11433), .B(n11437), .Z(n11435) );
  XNOR U11453 ( .A(n11438), .B(n11337), .Z(n11340) );
  XOR U11454 ( .A(n11439), .B(n11440), .Z(n11337) );
  AND U11455 ( .A(n11441), .B(n11442), .Z(n11440) );
  XOR U11456 ( .A(n11439), .B(n11443), .Z(n11441) );
  XNOR U11457 ( .A(n11444), .B(n11445), .Z(n11438) );
  NOR U11458 ( .A(n11446), .B(n11447), .Z(n11445) );
  XOR U11459 ( .A(n11444), .B(n11448), .Z(n11446) );
  XOR U11460 ( .A(n11330), .B(n11342), .Z(n11404) );
  AND U11461 ( .A(n11250), .B(n11449), .Z(n11342) );
  IV U11462 ( .A(n11229), .Z(n11250) );
  XNOR U11463 ( .A(n11348), .B(n11347), .Z(n11330) );
  XNOR U11464 ( .A(n11450), .B(n11353), .Z(n11347) );
  XOR U11465 ( .A(n11451), .B(n11452), .Z(n11353) );
  NOR U11466 ( .A(n11453), .B(n11454), .Z(n11452) );
  XNOR U11467 ( .A(n11451), .B(n11455), .Z(n11453) );
  XNOR U11468 ( .A(n11352), .B(n11344), .Z(n11450) );
  XOR U11469 ( .A(n11456), .B(n11457), .Z(n11344) );
  AND U11470 ( .A(n11458), .B(n11459), .Z(n11457) );
  XNOR U11471 ( .A(n11456), .B(n11460), .Z(n11458) );
  XNOR U11472 ( .A(n11461), .B(n11349), .Z(n11352) );
  XOR U11473 ( .A(n11462), .B(n11463), .Z(n11349) );
  AND U11474 ( .A(n11464), .B(n11465), .Z(n11463) );
  XOR U11475 ( .A(n11462), .B(n11466), .Z(n11464) );
  XNOR U11476 ( .A(n11467), .B(n11468), .Z(n11461) );
  NOR U11477 ( .A(n11469), .B(n11470), .Z(n11468) );
  XOR U11478 ( .A(n11467), .B(n11471), .Z(n11469) );
  XOR U11479 ( .A(n11358), .B(n11357), .Z(n11348) );
  XNOR U11480 ( .A(n11472), .B(n11354), .Z(n11357) );
  XOR U11481 ( .A(n11473), .B(n11474), .Z(n11354) );
  AND U11482 ( .A(n11475), .B(n11476), .Z(n11474) );
  XOR U11483 ( .A(n11473), .B(n11477), .Z(n11475) );
  XNOR U11484 ( .A(n11478), .B(n11479), .Z(n11472) );
  NOR U11485 ( .A(n11480), .B(n11481), .Z(n11479) );
  XNOR U11486 ( .A(n11478), .B(n11482), .Z(n11480) );
  XOR U11487 ( .A(n11483), .B(n11484), .Z(n11358) );
  NOR U11488 ( .A(n11485), .B(n11486), .Z(n11484) );
  XNOR U11489 ( .A(n11483), .B(n11487), .Z(n11485) );
  XNOR U11490 ( .A(n11488), .B(n11400), .Z(n11402) );
  IV U11491 ( .A(n11031), .Z(n11488) );
  XOR U11492 ( .A(n11489), .B(n11388), .Z(n11031) );
  XOR U11493 ( .A(n11366), .B(n11365), .Z(n11388) );
  XNOR U11494 ( .A(n11490), .B(n11371), .Z(n11365) );
  XOR U11495 ( .A(n11491), .B(n11492), .Z(n11371) );
  NOR U11496 ( .A(n11493), .B(n11494), .Z(n11492) );
  XNOR U11497 ( .A(n11491), .B(n11495), .Z(n11493) );
  XNOR U11498 ( .A(n11370), .B(n11362), .Z(n11490) );
  XOR U11499 ( .A(n11496), .B(n11497), .Z(n11362) );
  AND U11500 ( .A(n11498), .B(n11499), .Z(n11497) );
  XNOR U11501 ( .A(n11496), .B(n11500), .Z(n11498) );
  XNOR U11502 ( .A(n11501), .B(n11367), .Z(n11370) );
  XOR U11503 ( .A(n11502), .B(n11503), .Z(n11367) );
  AND U11504 ( .A(n11504), .B(n11505), .Z(n11503) );
  XOR U11505 ( .A(n11502), .B(n11506), .Z(n11504) );
  XNOR U11506 ( .A(n11507), .B(n11508), .Z(n11501) );
  NOR U11507 ( .A(n11509), .B(n11510), .Z(n11508) );
  XOR U11508 ( .A(n11507), .B(n11511), .Z(n11509) );
  XOR U11509 ( .A(n11376), .B(n11375), .Z(n11366) );
  XNOR U11510 ( .A(n11512), .B(n11372), .Z(n11375) );
  XOR U11511 ( .A(n11513), .B(n11514), .Z(n11372) );
  AND U11512 ( .A(n11515), .B(n11516), .Z(n11514) );
  XOR U11513 ( .A(n11513), .B(n11517), .Z(n11515) );
  XNOR U11514 ( .A(n11518), .B(n11519), .Z(n11512) );
  NOR U11515 ( .A(n11520), .B(n11521), .Z(n11519) );
  XNOR U11516 ( .A(n11518), .B(n11522), .Z(n11520) );
  XOR U11517 ( .A(n11523), .B(n11524), .Z(n11376) );
  NOR U11518 ( .A(n11525), .B(n11526), .Z(n11524) );
  XNOR U11519 ( .A(n11523), .B(n11527), .Z(n11525) );
  XNOR U11520 ( .A(n11387), .B(n11377), .Z(n11489) );
  AND U11521 ( .A(n11248), .B(n11528), .Z(n11377) );
  XNOR U11522 ( .A(n11529), .B(n11394), .Z(n11387) );
  XOR U11523 ( .A(n11383), .B(n11382), .Z(n11394) );
  XNOR U11524 ( .A(n11530), .B(n11379), .Z(n11382) );
  XOR U11525 ( .A(n11531), .B(n11532), .Z(n11379) );
  AND U11526 ( .A(n11533), .B(n11534), .Z(n11532) );
  XOR U11527 ( .A(n11531), .B(n11535), .Z(n11533) );
  XNOR U11528 ( .A(n11536), .B(n11537), .Z(n11530) );
  NOR U11529 ( .A(n11538), .B(n11539), .Z(n11537) );
  XNOR U11530 ( .A(n11536), .B(n11540), .Z(n11538) );
  XOR U11531 ( .A(n11541), .B(n11542), .Z(n11383) );
  NOR U11532 ( .A(n11543), .B(n11544), .Z(n11542) );
  XNOR U11533 ( .A(n11541), .B(n11545), .Z(n11543) );
  XNOR U11534 ( .A(n11393), .B(n11384), .Z(n11529) );
  XOR U11535 ( .A(n11546), .B(n11547), .Z(n11384) );
  NOR U11536 ( .A(n11548), .B(n11549), .Z(n11547) );
  XNOR U11537 ( .A(n11546), .B(n11550), .Z(n11548) );
  XOR U11538 ( .A(n11551), .B(n11399), .Z(n11393) );
  XNOR U11539 ( .A(n11552), .B(n11553), .Z(n11399) );
  NOR U11540 ( .A(n11554), .B(n11555), .Z(n11553) );
  XNOR U11541 ( .A(n11552), .B(n11556), .Z(n11554) );
  XNOR U11542 ( .A(n11398), .B(n11390), .Z(n11551) );
  XOR U11543 ( .A(n11557), .B(n11558), .Z(n11390) );
  AND U11544 ( .A(n11559), .B(n11560), .Z(n11558) );
  XOR U11545 ( .A(n11557), .B(n11561), .Z(n11559) );
  XNOR U11546 ( .A(n11562), .B(n11395), .Z(n11398) );
  XOR U11547 ( .A(n11563), .B(n11564), .Z(n11395) );
  AND U11548 ( .A(n11565), .B(n11566), .Z(n11564) );
  XOR U11549 ( .A(n11563), .B(n11567), .Z(n11565) );
  XNOR U11550 ( .A(n11568), .B(n11569), .Z(n11562) );
  NOR U11551 ( .A(n11570), .B(n11571), .Z(n11569) );
  XOR U11552 ( .A(n11568), .B(n11572), .Z(n11570) );
  AND U11553 ( .A(n11248), .B(n11229), .Z(n11400) );
  XNOR U11554 ( .A(n11573), .B(n11449), .Z(n11229) );
  XOR U11555 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][0] ), .B(
        p_input[512]), .Z(n11449) );
  XOR U11556 ( .A(n11426), .B(n11425), .Z(n11573) );
  XOR U11557 ( .A(n11574), .B(n11437), .Z(n11425) );
  XOR U11558 ( .A(n11411), .B(n11410), .Z(n11437) );
  XNOR U11559 ( .A(n11575), .B(n11416), .Z(n11410) );
  XOR U11560 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][24] ), .B(
        p_input[536]), .Z(n11416) );
  XOR U11561 ( .A(n11407), .B(n11415), .Z(n11575) );
  XOR U11562 ( .A(n11576), .B(n11412), .Z(n11415) );
  XOR U11563 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][22] ), .B(
        p_input[534]), .Z(n11412) );
  XOR U11564 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][23] ), .B(n6576), 
        .Z(n11576) );
  XNOR U11565 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][18] ), .B(n7313), 
        .Z(n11407) );
  XNOR U11566 ( .A(n11421), .B(n11420), .Z(n11411) );
  XOR U11567 ( .A(n11577), .B(n11417), .Z(n11420) );
  XOR U11568 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][19] ), .B(
        p_input[531]), .Z(n11417) );
  XOR U11569 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][20] ), .B(n6578), 
        .Z(n11577) );
  XOR U11570 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][21] ), .B(
        p_input[533]), .Z(n11421) );
  XNOR U11571 ( .A(n11436), .B(n11422), .Z(n11574) );
  XNOR U11572 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][1] ), .B(n7315), 
        .Z(n11422) );
  XNOR U11573 ( .A(n11578), .B(n11443), .Z(n11436) );
  XNOR U11574 ( .A(n11432), .B(n11431), .Z(n11443) );
  XOR U11575 ( .A(n11579), .B(n11428), .Z(n11431) );
  XNOR U11576 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][26] ), .B(n6951), 
        .Z(n11428) );
  XOR U11577 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][27] ), .B(n6582), 
        .Z(n11579) );
  XOR U11578 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][28] ), .B(
        p_input[540]), .Z(n11432) );
  XNOR U11579 ( .A(n11442), .B(n11433), .Z(n11578) );
  XNOR U11580 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][17] ), .B(n7318), 
        .Z(n11433) );
  XOR U11581 ( .A(n11580), .B(n11448), .Z(n11442) );
  XNOR U11582 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][31] ), .B(
        p_input[543]), .Z(n11448) );
  XOR U11583 ( .A(n11439), .B(n11447), .Z(n11580) );
  XOR U11584 ( .A(n11581), .B(n11444), .Z(n11447) );
  XOR U11585 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][29] ), .B(
        p_input[541]), .Z(n11444) );
  XOR U11586 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][30] ), .B(n6587), 
        .Z(n11581) );
  XNOR U11587 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][25] ), .B(n6955), 
        .Z(n11439) );
  XNOR U11588 ( .A(n11460), .B(n11459), .Z(n11426) );
  XNOR U11589 ( .A(n11582), .B(n11466), .Z(n11459) );
  XNOR U11590 ( .A(n11455), .B(n11454), .Z(n11466) );
  XOR U11591 ( .A(n11583), .B(n11451), .Z(n11454) );
  XNOR U11592 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][11] ), .B(n7323), 
        .Z(n11451) );
  XOR U11593 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][12] ), .B(n6590), 
        .Z(n11583) );
  XOR U11594 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][13] ), .B(
        p_input[525]), .Z(n11455) );
  XNOR U11595 ( .A(n11465), .B(n11456), .Z(n11582) );
  XNOR U11596 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][2] ), .B(n7324), 
        .Z(n11456) );
  XOR U11597 ( .A(n11584), .B(n11471), .Z(n11465) );
  XNOR U11598 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][16] ), .B(
        p_input[528]), .Z(n11471) );
  XOR U11599 ( .A(n11462), .B(n11470), .Z(n11584) );
  XOR U11600 ( .A(n11585), .B(n11467), .Z(n11470) );
  XOR U11601 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][14] ), .B(
        p_input[526]), .Z(n11467) );
  XOR U11602 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][15] ), .B(n6595), 
        .Z(n11585) );
  XNOR U11603 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][10] ), .B(n7327), 
        .Z(n11462) );
  XNOR U11604 ( .A(n11477), .B(n11476), .Z(n11460) );
  XNOR U11605 ( .A(n11586), .B(n11482), .Z(n11476) );
  XNOR U11606 ( .A(n380), .B(p_input[521]), .Z(n11482) );
  IV U11607 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][9] ), .Z(n380) );
  XOR U11608 ( .A(n11473), .B(n11481), .Z(n11586) );
  XOR U11609 ( .A(n11587), .B(n11478), .Z(n11481) );
  XNOR U11610 ( .A(n764), .B(p_input[519]), .Z(n11478) );
  IV U11611 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][7] ), .Z(n764) );
  XOR U11612 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][8] ), .B(n6963), 
        .Z(n11587) );
  XNOR U11613 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][3] ), .B(n7330), 
        .Z(n11473) );
  XNOR U11614 ( .A(n11487), .B(n11486), .Z(n11477) );
  XOR U11615 ( .A(n11588), .B(n11483), .Z(n11486) );
  XOR U11616 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][4] ), .B(
        p_input[516]), .Z(n11483) );
  XOR U11617 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][5] ), .B(n6965), 
        .Z(n11588) );
  XOR U11618 ( .A(\knn_comb_/ASN_1[1].knn_/local_min_val[1][6] ), .B(
        p_input[518]), .Z(n11487) );
  XOR U11619 ( .A(n11589), .B(n11550), .Z(n11248) );
  XNOR U11620 ( .A(n11500), .B(n11499), .Z(n11550) );
  XNOR U11621 ( .A(n11590), .B(n11506), .Z(n11499) );
  XNOR U11622 ( .A(n11495), .B(n11494), .Z(n11506) );
  XOR U11623 ( .A(n11591), .B(n11491), .Z(n11494) );
  XNOR U11624 ( .A(\knn_comb_/min_val_out[0][11] ), .B(n7323), .Z(n11491) );
  IV U11625 ( .A(p_input[523]), .Z(n7323) );
  XOR U11626 ( .A(\knn_comb_/min_val_out[0][12] ), .B(n6590), .Z(n11591) );
  IV U11627 ( .A(p_input[524]), .Z(n6590) );
  XOR U11628 ( .A(\knn_comb_/min_val_out[0][13] ), .B(p_input[525]), .Z(n11495) );
  XNOR U11629 ( .A(n11505), .B(n11496), .Z(n11590) );
  XNOR U11630 ( .A(\knn_comb_/min_val_out[0][2] ), .B(n7324), .Z(n11496) );
  IV U11631 ( .A(p_input[514]), .Z(n7324) );
  XOR U11632 ( .A(n11592), .B(n11511), .Z(n11505) );
  XNOR U11633 ( .A(\knn_comb_/min_val_out[0][16] ), .B(p_input[528]), .Z(
        n11511) );
  XOR U11634 ( .A(n11502), .B(n11510), .Z(n11592) );
  XOR U11635 ( .A(n11593), .B(n11507), .Z(n11510) );
  XOR U11636 ( .A(\knn_comb_/min_val_out[0][14] ), .B(p_input[526]), .Z(n11507) );
  XOR U11637 ( .A(\knn_comb_/min_val_out[0][15] ), .B(n6595), .Z(n11593) );
  IV U11638 ( .A(p_input[527]), .Z(n6595) );
  XNOR U11639 ( .A(\knn_comb_/min_val_out[0][10] ), .B(n7327), .Z(n11502) );
  IV U11640 ( .A(p_input[522]), .Z(n7327) );
  XNOR U11641 ( .A(n11517), .B(n11516), .Z(n11500) );
  XNOR U11642 ( .A(n11594), .B(n11522), .Z(n11516) );
  XNOR U11643 ( .A(n379), .B(p_input[521]), .Z(n11522) );
  IV U11644 ( .A(\knn_comb_/min_val_out[0][9] ), .Z(n379) );
  XOR U11645 ( .A(n11513), .B(n11521), .Z(n11594) );
  XOR U11646 ( .A(n11595), .B(n11518), .Z(n11521) );
  XNOR U11647 ( .A(n763), .B(p_input[519]), .Z(n11518) );
  IV U11648 ( .A(\knn_comb_/min_val_out[0][7] ), .Z(n763) );
  XOR U11649 ( .A(\knn_comb_/min_val_out[0][8] ), .B(n6963), .Z(n11595) );
  IV U11650 ( .A(p_input[520]), .Z(n6963) );
  XNOR U11651 ( .A(\knn_comb_/min_val_out[0][3] ), .B(n7330), .Z(n11513) );
  IV U11652 ( .A(p_input[515]), .Z(n7330) );
  XNOR U11653 ( .A(n11527), .B(n11526), .Z(n11517) );
  XOR U11654 ( .A(n11596), .B(n11523), .Z(n11526) );
  XOR U11655 ( .A(\knn_comb_/min_val_out[0][4] ), .B(p_input[516]), .Z(n11523)
         );
  XOR U11656 ( .A(\knn_comb_/min_val_out[0][5] ), .B(n6965), .Z(n11596) );
  IV U11657 ( .A(p_input[517]), .Z(n6965) );
  XOR U11658 ( .A(\knn_comb_/min_val_out[0][6] ), .B(p_input[518]), .Z(n11527)
         );
  XOR U11659 ( .A(n11549), .B(n11528), .Z(n11589) );
  XOR U11660 ( .A(\knn_comb_/min_val_out[0][0] ), .B(p_input[512]), .Z(n11528)
         );
  XOR U11661 ( .A(n11597), .B(n11561), .Z(n11549) );
  XOR U11662 ( .A(n11535), .B(n11534), .Z(n11561) );
  XNOR U11663 ( .A(n11598), .B(n11540), .Z(n11534) );
  XOR U11664 ( .A(\knn_comb_/min_val_out[0][24] ), .B(p_input[536]), .Z(n11540) );
  XOR U11665 ( .A(n11531), .B(n11539), .Z(n11598) );
  XOR U11666 ( .A(n11599), .B(n11536), .Z(n11539) );
  XOR U11667 ( .A(\knn_comb_/min_val_out[0][22] ), .B(p_input[534]), .Z(n11536) );
  XOR U11668 ( .A(\knn_comb_/min_val_out[0][23] ), .B(n6576), .Z(n11599) );
  IV U11669 ( .A(p_input[535]), .Z(n6576) );
  XNOR U11670 ( .A(\knn_comb_/min_val_out[0][18] ), .B(n7313), .Z(n11531) );
  IV U11671 ( .A(p_input[530]), .Z(n7313) );
  XNOR U11672 ( .A(n11545), .B(n11544), .Z(n11535) );
  XOR U11673 ( .A(n11600), .B(n11541), .Z(n11544) );
  XOR U11674 ( .A(\knn_comb_/min_val_out[0][19] ), .B(p_input[531]), .Z(n11541) );
  XOR U11675 ( .A(\knn_comb_/min_val_out[0][20] ), .B(n6578), .Z(n11600) );
  IV U11676 ( .A(p_input[532]), .Z(n6578) );
  XOR U11677 ( .A(\knn_comb_/min_val_out[0][21] ), .B(p_input[533]), .Z(n11545) );
  XNOR U11678 ( .A(n11560), .B(n11546), .Z(n11597) );
  XNOR U11679 ( .A(\knn_comb_/min_val_out[0][1] ), .B(n7315), .Z(n11546) );
  IV U11680 ( .A(p_input[513]), .Z(n7315) );
  XNOR U11681 ( .A(n11601), .B(n11567), .Z(n11560) );
  XNOR U11682 ( .A(n11556), .B(n11555), .Z(n11567) );
  XOR U11683 ( .A(n11602), .B(n11552), .Z(n11555) );
  XNOR U11684 ( .A(\knn_comb_/min_val_out[0][26] ), .B(n6951), .Z(n11552) );
  IV U11685 ( .A(p_input[538]), .Z(n6951) );
  XOR U11686 ( .A(\knn_comb_/min_val_out[0][27] ), .B(n6582), .Z(n11602) );
  IV U11687 ( .A(p_input[539]), .Z(n6582) );
  XOR U11688 ( .A(\knn_comb_/min_val_out[0][28] ), .B(p_input[540]), .Z(n11556) );
  XNOR U11689 ( .A(n11566), .B(n11557), .Z(n11601) );
  XNOR U11690 ( .A(\knn_comb_/min_val_out[0][17] ), .B(n7318), .Z(n11557) );
  IV U11691 ( .A(p_input[529]), .Z(n7318) );
  XOR U11692 ( .A(n11603), .B(n11572), .Z(n11566) );
  XNOR U11693 ( .A(\knn_comb_/min_val_out[0][31] ), .B(p_input[543]), .Z(
        n11572) );
  XOR U11694 ( .A(n11563), .B(n11571), .Z(n11603) );
  XOR U11695 ( .A(n11604), .B(n11568), .Z(n11571) );
  XOR U11696 ( .A(\knn_comb_/min_val_out[0][29] ), .B(p_input[541]), .Z(n11568) );
  XOR U11697 ( .A(\knn_comb_/min_val_out[0][30] ), .B(n6587), .Z(n11604) );
  IV U11698 ( .A(p_input[542]), .Z(n6587) );
  XNOR U11699 ( .A(\knn_comb_/min_val_out[0][25] ), .B(n6955), .Z(n11563) );
  IV U11700 ( .A(p_input[537]), .Z(n6955) );
endmodule

